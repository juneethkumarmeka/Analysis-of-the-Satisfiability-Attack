module basic_2500_25000_3000_10_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_645,In_157);
nand U1 (N_1,In_867,In_2404);
or U2 (N_2,In_669,In_2054);
nor U3 (N_3,In_1189,In_1831);
or U4 (N_4,In_592,In_861);
nand U5 (N_5,In_182,In_1178);
or U6 (N_6,In_1557,In_2289);
nand U7 (N_7,In_1878,In_2471);
nand U8 (N_8,In_98,In_1773);
xor U9 (N_9,In_2055,In_1924);
nor U10 (N_10,In_1143,In_128);
or U11 (N_11,In_1346,In_943);
or U12 (N_12,In_1607,In_2195);
nand U13 (N_13,In_928,In_175);
nand U14 (N_14,In_2419,In_719);
nand U15 (N_15,In_1930,In_1414);
or U16 (N_16,In_1226,In_1903);
and U17 (N_17,In_268,In_1083);
nor U18 (N_18,In_1036,In_1888);
nand U19 (N_19,In_1141,In_264);
or U20 (N_20,In_2359,In_1181);
nand U21 (N_21,In_144,In_1644);
nand U22 (N_22,In_2433,In_2282);
or U23 (N_23,In_718,In_988);
nand U24 (N_24,In_2081,In_726);
or U25 (N_25,In_2337,In_2480);
or U26 (N_26,In_1906,In_292);
nand U27 (N_27,In_1138,In_1545);
nor U28 (N_28,In_1011,In_1761);
or U29 (N_29,In_2265,In_2116);
and U30 (N_30,In_1330,In_2018);
nand U31 (N_31,In_2271,In_1871);
or U32 (N_32,In_1328,In_1269);
and U33 (N_33,In_821,In_1240);
xnor U34 (N_34,In_2113,In_320);
nand U35 (N_35,In_1858,In_735);
or U36 (N_36,In_449,In_2462);
and U37 (N_37,In_1565,In_565);
nand U38 (N_38,In_1061,In_1837);
or U39 (N_39,In_2415,In_2365);
nand U40 (N_40,In_2343,In_627);
or U41 (N_41,In_1267,In_37);
nand U42 (N_42,In_2384,In_749);
nand U43 (N_43,In_906,In_2028);
and U44 (N_44,In_262,In_608);
nor U45 (N_45,In_319,In_2331);
xnor U46 (N_46,In_2021,In_2290);
and U47 (N_47,In_458,In_1253);
nand U48 (N_48,In_1881,In_1265);
or U49 (N_49,In_1772,In_945);
xor U50 (N_50,In_790,In_1437);
or U51 (N_51,In_1742,In_555);
nand U52 (N_52,In_2294,In_2315);
nand U53 (N_53,In_2225,In_1343);
and U54 (N_54,In_2106,In_2342);
and U55 (N_55,In_2196,In_2308);
nand U56 (N_56,In_1608,In_437);
xnor U57 (N_57,In_1818,In_1839);
xor U58 (N_58,In_934,In_2114);
or U59 (N_59,In_305,In_1869);
xnor U60 (N_60,In_1605,In_1922);
nand U61 (N_61,In_623,In_1499);
and U62 (N_62,In_1713,In_1337);
or U63 (N_63,In_1725,In_249);
or U64 (N_64,In_886,In_211);
and U65 (N_65,In_206,In_956);
or U66 (N_66,In_139,In_824);
or U67 (N_67,In_1769,In_465);
nand U68 (N_68,In_17,In_2256);
nand U69 (N_69,In_523,In_2060);
and U70 (N_70,In_926,In_579);
nand U71 (N_71,In_1600,In_2340);
nand U72 (N_72,In_279,In_542);
or U73 (N_73,In_2356,In_978);
or U74 (N_74,In_922,In_79);
and U75 (N_75,In_870,In_10);
or U76 (N_76,In_1179,In_130);
nand U77 (N_77,In_609,In_2170);
and U78 (N_78,In_2279,In_1079);
and U79 (N_79,In_1307,In_1099);
nor U80 (N_80,In_487,In_2352);
or U81 (N_81,In_2448,In_1085);
and U82 (N_82,In_1955,In_1052);
xor U83 (N_83,In_2067,In_509);
or U84 (N_84,In_911,In_1149);
nand U85 (N_85,In_2309,In_1554);
nor U86 (N_86,In_2453,In_2232);
and U87 (N_87,In_1126,In_1579);
nand U88 (N_88,In_1205,In_60);
and U89 (N_89,In_2373,In_2161);
and U90 (N_90,In_2201,In_962);
and U91 (N_91,In_2378,In_1984);
and U92 (N_92,In_1494,In_1689);
or U93 (N_93,In_2095,In_1824);
and U94 (N_94,In_226,In_161);
or U95 (N_95,In_1251,In_1191);
nor U96 (N_96,In_2082,In_2367);
or U97 (N_97,In_2094,In_1076);
and U98 (N_98,In_2413,In_877);
and U99 (N_99,In_1302,In_860);
nand U100 (N_100,In_1175,In_101);
nor U101 (N_101,In_1020,In_2389);
and U102 (N_102,In_1846,In_1314);
or U103 (N_103,In_622,In_1441);
and U104 (N_104,In_1650,In_2109);
nand U105 (N_105,In_1012,In_1326);
or U106 (N_106,In_2108,In_1788);
nand U107 (N_107,In_1505,In_1956);
and U108 (N_108,In_2068,In_242);
and U109 (N_109,In_2045,In_1610);
nand U110 (N_110,In_879,In_1192);
nand U111 (N_111,In_1682,In_952);
and U112 (N_112,In_941,In_479);
nor U113 (N_113,In_1901,In_2085);
nand U114 (N_114,In_740,In_6);
xnor U115 (N_115,In_2175,In_2385);
nand U116 (N_116,In_352,In_1047);
and U117 (N_117,In_1448,In_572);
or U118 (N_118,In_2303,In_1700);
xor U119 (N_119,In_2307,In_1528);
and U120 (N_120,In_968,In_1640);
and U121 (N_121,In_1213,In_1292);
and U122 (N_122,In_2463,In_1680);
nand U123 (N_123,In_142,In_1703);
nand U124 (N_124,In_1028,In_1458);
nand U125 (N_125,In_61,In_1690);
nand U126 (N_126,In_371,In_2469);
nor U127 (N_127,In_1926,In_2405);
or U128 (N_128,In_644,In_1928);
nor U129 (N_129,In_713,In_1790);
nand U130 (N_130,In_1540,In_2251);
nand U131 (N_131,In_2358,In_257);
or U132 (N_132,In_1524,In_250);
or U133 (N_133,In_2286,In_1355);
or U134 (N_134,In_2046,In_1856);
and U135 (N_135,In_2040,In_1870);
and U136 (N_136,In_778,In_2016);
nor U137 (N_137,In_1523,In_648);
and U138 (N_138,In_1646,In_1936);
xor U139 (N_139,In_1058,In_1407);
and U140 (N_140,In_2386,In_1370);
or U141 (N_141,In_413,In_984);
nand U142 (N_142,In_341,In_2066);
or U143 (N_143,In_1492,In_1546);
nand U144 (N_144,In_57,In_102);
nand U145 (N_145,In_875,In_436);
and U146 (N_146,In_1185,In_935);
xnor U147 (N_147,In_699,In_1342);
nor U148 (N_148,In_818,In_951);
and U149 (N_149,In_1549,In_1595);
nand U150 (N_150,In_854,In_183);
or U151 (N_151,In_1077,In_1351);
or U152 (N_152,In_1368,In_1257);
nand U153 (N_153,In_1807,In_1765);
xor U154 (N_154,In_2173,In_1110);
or U155 (N_155,In_460,In_727);
or U156 (N_156,In_1538,In_307);
nor U157 (N_157,In_480,In_7);
and U158 (N_158,In_2422,In_516);
or U159 (N_159,In_885,In_2211);
or U160 (N_160,In_425,In_363);
nor U161 (N_161,In_2276,In_2351);
and U162 (N_162,In_357,In_1197);
xor U163 (N_163,In_546,In_1551);
or U164 (N_164,In_1416,In_905);
nor U165 (N_165,In_99,In_184);
or U166 (N_166,In_1569,In_2150);
nor U167 (N_167,In_2270,In_1186);
and U168 (N_168,In_1025,In_800);
or U169 (N_169,In_1622,In_1805);
nand U170 (N_170,In_2187,In_167);
and U171 (N_171,In_1744,In_1793);
xor U172 (N_172,In_1239,In_300);
or U173 (N_173,In_400,In_725);
nand U174 (N_174,In_1043,In_2058);
nand U175 (N_175,In_317,In_2197);
nor U176 (N_176,In_1559,In_306);
xnor U177 (N_177,In_799,In_16);
or U178 (N_178,In_1714,In_692);
nand U179 (N_179,In_561,In_1335);
xor U180 (N_180,In_775,In_2119);
nand U181 (N_181,In_1300,In_2052);
xor U182 (N_182,In_1027,In_2362);
and U183 (N_183,In_1392,In_2442);
and U184 (N_184,In_414,In_1225);
nor U185 (N_185,In_596,In_49);
and U186 (N_186,In_486,In_1723);
and U187 (N_187,In_2032,In_2084);
xnor U188 (N_188,In_1276,In_1954);
nand U189 (N_189,In_366,In_930);
xor U190 (N_190,In_1578,In_2283);
nor U191 (N_191,In_1951,In_2247);
and U192 (N_192,In_1188,In_636);
xnor U193 (N_193,In_1850,In_393);
and U194 (N_194,In_2280,In_2498);
nor U195 (N_195,In_1223,In_1291);
nand U196 (N_196,In_443,In_360);
nand U197 (N_197,In_2379,In_1115);
nand U198 (N_198,In_214,In_24);
and U199 (N_199,In_798,In_859);
and U200 (N_200,In_668,In_2155);
or U201 (N_201,In_154,In_1660);
and U202 (N_202,In_2482,In_1763);
and U203 (N_203,In_1486,In_2138);
or U204 (N_204,In_331,In_2468);
and U205 (N_205,In_2380,In_2179);
nor U206 (N_206,In_981,In_1325);
or U207 (N_207,In_1344,In_839);
or U208 (N_208,In_782,In_25);
xnor U209 (N_209,In_971,In_630);
or U210 (N_210,In_403,In_2325);
nor U211 (N_211,In_567,In_328);
nand U212 (N_212,In_1566,In_1576);
nand U213 (N_213,In_2439,In_478);
xor U214 (N_214,In_667,In_963);
xor U215 (N_215,In_2222,In_1718);
and U216 (N_216,In_1720,In_1514);
nor U217 (N_217,In_993,In_1161);
nor U218 (N_218,In_41,In_601);
and U219 (N_219,In_1740,In_791);
nand U220 (N_220,In_1018,In_1567);
or U221 (N_221,In_1921,In_1460);
nor U222 (N_222,In_1998,In_1602);
or U223 (N_223,In_2117,In_1993);
nand U224 (N_224,In_68,In_767);
or U225 (N_225,In_633,In_1480);
and U226 (N_226,In_2131,In_260);
or U227 (N_227,In_619,In_1709);
or U228 (N_228,In_2355,In_841);
or U229 (N_229,In_1521,In_1203);
nand U230 (N_230,In_2485,In_1775);
nor U231 (N_231,In_698,In_1641);
xor U232 (N_232,In_180,In_624);
and U233 (N_233,In_634,In_1677);
xor U234 (N_234,In_1562,In_241);
or U235 (N_235,In_86,In_2295);
or U236 (N_236,In_876,In_1746);
and U237 (N_237,In_1541,In_1451);
xor U238 (N_238,In_2475,In_2377);
nand U239 (N_239,In_1748,In_852);
or U240 (N_240,In_2228,In_689);
nand U241 (N_241,In_477,In_646);
and U242 (N_242,In_2078,In_2091);
xor U243 (N_243,In_1481,In_2031);
and U244 (N_244,In_1676,In_140);
and U245 (N_245,In_1361,In_1367);
xnor U246 (N_246,In_238,In_2151);
xor U247 (N_247,In_2235,In_1943);
nand U248 (N_248,In_893,In_1041);
or U249 (N_249,In_1167,In_1753);
xor U250 (N_250,In_1310,In_1296);
nor U251 (N_251,In_571,In_2159);
or U252 (N_252,In_2072,In_398);
and U253 (N_253,In_2242,In_429);
nor U254 (N_254,In_408,In_1374);
nand U255 (N_255,In_2112,In_1611);
and U256 (N_256,In_2266,In_370);
nand U257 (N_257,In_2318,In_1639);
or U258 (N_258,In_2446,In_677);
or U259 (N_259,In_1652,In_2328);
and U260 (N_260,In_1661,In_2486);
nand U261 (N_261,In_783,In_1455);
nand U262 (N_262,In_1065,In_469);
nand U263 (N_263,In_1270,In_1679);
and U264 (N_264,In_954,In_1177);
or U265 (N_265,In_858,In_1909);
nand U266 (N_266,In_1667,In_1397);
nor U267 (N_267,In_2053,In_904);
nor U268 (N_268,In_2157,In_452);
xnor U269 (N_269,In_1316,In_552);
and U270 (N_270,In_2275,In_1379);
and U271 (N_271,In_1444,In_1996);
and U272 (N_272,In_846,In_549);
xor U273 (N_273,In_1030,In_1349);
nor U274 (N_274,In_35,In_2427);
nor U275 (N_275,In_1057,In_510);
nand U276 (N_276,In_751,In_2438);
nor U277 (N_277,In_1868,In_953);
nor U278 (N_278,In_58,In_1506);
nor U279 (N_279,In_1082,In_1393);
or U280 (N_280,In_1822,In_1697);
xnor U281 (N_281,In_2341,In_2437);
and U282 (N_282,In_817,In_64);
nand U283 (N_283,In_1983,In_2350);
and U284 (N_284,In_1208,In_686);
or U285 (N_285,In_433,In_1080);
nand U286 (N_286,In_2217,In_1732);
nor U287 (N_287,In_1518,In_2497);
nand U288 (N_288,In_13,In_2035);
nor U289 (N_289,In_382,In_1303);
nor U290 (N_290,In_942,In_1591);
nor U291 (N_291,In_1892,In_2057);
nand U292 (N_292,In_1716,In_1702);
and U293 (N_293,In_569,In_856);
or U294 (N_294,In_362,In_266);
nand U295 (N_295,In_2144,In_696);
or U296 (N_296,In_2069,In_1804);
or U297 (N_297,In_1931,In_2165);
and U298 (N_298,In_1802,In_333);
nand U299 (N_299,In_54,In_1467);
nor U300 (N_300,In_1979,In_1550);
nor U301 (N_301,In_421,In_2255);
or U302 (N_302,In_1814,In_1848);
xnor U303 (N_303,In_671,In_832);
nand U304 (N_304,In_2003,In_2076);
or U305 (N_305,In_2499,In_1133);
xnor U306 (N_306,In_695,In_1163);
nand U307 (N_307,In_1687,In_294);
nor U308 (N_308,In_2183,In_618);
or U309 (N_309,In_1162,In_1264);
or U310 (N_310,In_177,In_499);
nor U311 (N_311,In_1321,In_1948);
nand U312 (N_312,In_1332,In_743);
or U313 (N_313,In_1182,In_69);
and U314 (N_314,In_51,In_109);
and U315 (N_315,In_2220,In_375);
nand U316 (N_316,In_75,In_805);
or U317 (N_317,In_958,In_899);
nand U318 (N_318,In_1504,In_1781);
nor U319 (N_319,In_426,In_2444);
or U320 (N_320,In_2237,In_97);
nand U321 (N_321,In_896,In_271);
or U322 (N_322,In_1318,In_2403);
and U323 (N_323,In_2002,In_1598);
nor U324 (N_324,In_195,In_105);
and U325 (N_325,In_2477,In_597);
and U326 (N_326,In_1560,In_1568);
and U327 (N_327,In_2353,In_1920);
nand U328 (N_328,In_138,In_1176);
and U329 (N_329,In_2014,In_1095);
nor U330 (N_330,In_1299,In_1705);
nand U331 (N_331,In_197,In_297);
and U332 (N_332,In_1454,In_678);
nor U333 (N_333,In_253,In_1707);
or U334 (N_334,In_2322,In_1685);
nand U335 (N_335,In_1945,In_655);
nor U336 (N_336,In_525,In_1730);
or U337 (N_337,In_461,In_1840);
nor U338 (N_338,In_759,In_2388);
xnor U339 (N_339,In_715,In_77);
xor U340 (N_340,In_1678,In_1465);
xnor U341 (N_341,In_663,In_496);
nand U342 (N_342,In_1241,In_445);
nand U343 (N_343,In_766,In_658);
or U344 (N_344,In_1385,In_1366);
xor U345 (N_345,In_424,In_1760);
nor U346 (N_346,In_729,In_2145);
or U347 (N_347,In_2412,In_190);
nor U348 (N_348,In_309,In_794);
and U349 (N_349,In_121,In_1633);
nor U350 (N_350,In_2007,In_2411);
or U351 (N_351,In_1313,In_863);
nor U352 (N_352,In_342,In_2169);
nor U353 (N_353,In_1669,In_777);
nor U354 (N_354,In_924,In_1966);
nor U355 (N_355,In_2261,In_1311);
xnor U356 (N_356,In_474,In_1168);
nor U357 (N_357,In_450,In_558);
and U358 (N_358,In_526,In_2493);
or U359 (N_359,In_1803,In_1245);
or U360 (N_360,In_1075,In_194);
xnor U361 (N_361,In_638,In_2432);
or U362 (N_362,In_1575,In_148);
or U363 (N_363,In_2020,In_240);
or U364 (N_364,In_672,In_772);
or U365 (N_365,In_311,In_2314);
and U366 (N_366,In_216,In_1599);
and U367 (N_367,In_171,In_1919);
and U368 (N_368,In_2172,In_1396);
nor U369 (N_369,In_1672,In_2181);
or U370 (N_370,In_1668,In_1787);
nand U371 (N_371,In_2304,In_2042);
xor U372 (N_372,In_1195,In_1777);
nor U373 (N_373,In_570,In_227);
nand U374 (N_374,In_541,In_2260);
or U375 (N_375,In_534,In_2061);
nand U376 (N_376,In_593,In_1000);
nor U377 (N_377,In_1698,In_2296);
nand U378 (N_378,In_539,In_2186);
nor U379 (N_379,In_489,In_936);
nand U380 (N_380,In_302,In_2148);
nand U381 (N_381,In_908,In_1354);
or U382 (N_382,In_915,In_106);
xnor U383 (N_383,In_1,In_2125);
nor U384 (N_384,In_965,In_673);
nor U385 (N_385,In_2206,In_347);
or U386 (N_386,In_612,In_491);
and U387 (N_387,In_2000,In_234);
nand U388 (N_388,In_312,In_2123);
nand U389 (N_389,In_2402,In_1563);
and U390 (N_390,In_1784,In_1386);
nand U391 (N_391,In_372,In_18);
or U392 (N_392,In_276,In_1908);
or U393 (N_393,In_0,In_742);
or U394 (N_394,In_163,In_607);
nor U395 (N_395,In_236,In_2126);
or U396 (N_396,In_2259,In_1135);
nor U397 (N_397,In_1737,In_210);
nand U398 (N_398,In_625,In_2209);
or U399 (N_399,In_530,In_1169);
and U400 (N_400,In_1688,In_223);
and U401 (N_401,In_531,In_2115);
xor U402 (N_402,In_198,In_1778);
nand U403 (N_403,In_652,In_1498);
nor U404 (N_404,In_284,In_2167);
nor U405 (N_405,In_476,In_2346);
nor U406 (N_406,In_1063,In_215);
or U407 (N_407,In_1603,In_1046);
nor U408 (N_408,In_156,In_1529);
nand U409 (N_409,In_1066,In_2401);
xnor U410 (N_410,In_1235,In_1774);
nand U411 (N_411,In_844,In_917);
or U412 (N_412,In_1456,In_1522);
and U413 (N_413,In_15,In_1347);
nand U414 (N_414,In_2090,In_2387);
or U415 (N_415,In_34,In_1331);
nor U416 (N_416,In_120,In_641);
nor U417 (N_417,In_721,In_573);
xnor U418 (N_418,In_2435,In_162);
and U419 (N_419,In_1715,In_2335);
nand U420 (N_420,In_1902,In_127);
and U421 (N_421,In_131,In_595);
nor U422 (N_422,In_472,In_1665);
nor U423 (N_423,In_1937,In_1572);
nor U424 (N_424,In_1693,In_354);
nand U425 (N_425,In_1621,In_1584);
nor U426 (N_426,In_392,In_1874);
nand U427 (N_427,In_1972,In_475);
or U428 (N_428,In_1237,In_399);
or U429 (N_429,In_473,In_724);
or U430 (N_430,In_2461,In_882);
or U431 (N_431,In_2124,In_1153);
nor U432 (N_432,In_1333,In_902);
and U433 (N_433,In_3,In_1675);
nand U434 (N_434,In_43,In_1210);
and U435 (N_435,In_324,In_178);
xor U436 (N_436,In_674,In_462);
and U437 (N_437,In_1647,In_2224);
and U438 (N_438,In_1103,In_2354);
nand U439 (N_439,In_345,In_807);
xnor U440 (N_440,In_2417,In_961);
nor U441 (N_441,In_731,In_1638);
nand U442 (N_442,In_1116,In_2025);
or U443 (N_443,In_2110,In_969);
nand U444 (N_444,In_4,In_1320);
xor U445 (N_445,In_2381,In_1101);
nor U446 (N_446,In_851,In_568);
or U447 (N_447,In_1286,In_949);
and U448 (N_448,In_1403,In_1424);
and U449 (N_449,In_583,In_2193);
nand U450 (N_450,In_702,In_1446);
nor U451 (N_451,In_2202,In_2252);
nand U452 (N_452,In_2460,In_1425);
nor U453 (N_453,In_1277,In_1917);
xor U454 (N_454,In_1957,In_827);
or U455 (N_455,In_1691,In_803);
nor U456 (N_456,In_2357,In_470);
or U457 (N_457,In_997,In_1463);
and U458 (N_458,In_1755,In_932);
and U459 (N_459,In_2240,In_1613);
nand U460 (N_460,In_2476,In_385);
xnor U461 (N_461,In_2324,In_410);
nand U462 (N_462,In_816,In_1234);
and U463 (N_463,In_2277,In_22);
xor U464 (N_464,In_2496,In_1695);
nand U465 (N_465,In_1420,In_1604);
nand U466 (N_466,In_1671,In_2174);
and U467 (N_467,In_590,In_1329);
nor U468 (N_468,In_849,In_2249);
and U469 (N_469,In_787,In_979);
nand U470 (N_470,In_1373,In_1829);
xor U471 (N_471,In_1096,In_1847);
and U472 (N_472,In_872,In_145);
nor U473 (N_473,In_1068,In_1206);
or U474 (N_474,In_1734,In_258);
or U475 (N_475,In_205,In_213);
or U476 (N_476,In_1144,In_221);
or U477 (N_477,In_2473,In_517);
nor U478 (N_478,In_2214,In_2288);
nor U479 (N_479,In_1340,In_1490);
or U480 (N_480,In_2243,In_2374);
nand U481 (N_481,In_2063,In_1991);
nand U482 (N_482,In_84,In_927);
and U483 (N_483,In_514,In_432);
nor U484 (N_484,In_390,In_1973);
nand U485 (N_485,In_2323,In_451);
and U486 (N_486,In_1722,In_2447);
or U487 (N_487,In_1193,In_1745);
nand U488 (N_488,In_1864,In_176);
nand U489 (N_489,In_528,In_2208);
and U490 (N_490,In_299,In_1724);
nor U491 (N_491,In_739,In_2319);
and U492 (N_492,In_2080,In_1415);
or U493 (N_493,In_1290,In_656);
nor U494 (N_494,In_792,In_1625);
nor U495 (N_495,In_966,In_2133);
nor U496 (N_496,In_871,In_1227);
and U497 (N_497,In_2121,In_828);
and U498 (N_498,In_1812,In_1468);
or U499 (N_499,In_675,In_1889);
xor U500 (N_500,In_348,In_282);
xor U501 (N_501,In_1735,In_365);
or U502 (N_502,In_2316,In_1872);
or U503 (N_503,In_251,In_1664);
xnor U504 (N_504,In_1119,In_1547);
nor U505 (N_505,In_1449,In_1759);
nand U506 (N_506,In_237,In_2234);
nor U507 (N_507,In_1259,In_1158);
nor U508 (N_508,In_757,In_1801);
nor U509 (N_509,In_842,In_1634);
xor U510 (N_510,In_378,In_1038);
nand U511 (N_511,In_33,In_1552);
nand U512 (N_512,In_1196,In_321);
nor U513 (N_513,In_289,In_1890);
nand U514 (N_514,In_2176,In_351);
and U515 (N_515,In_1089,In_1623);
nand U516 (N_516,In_1215,In_763);
nor U517 (N_517,In_606,In_887);
nor U518 (N_518,In_2223,In_1914);
nand U519 (N_519,In_2305,In_2297);
nand U520 (N_520,In_1743,In_975);
or U521 (N_521,In_553,In_838);
and U522 (N_522,In_1894,In_1232);
or U523 (N_523,In_1339,In_891);
nor U524 (N_524,In_1010,In_967);
nand U525 (N_525,In_2096,In_1004);
xor U526 (N_526,In_2034,In_2246);
nor U527 (N_527,In_1139,In_2393);
and U528 (N_528,In_1527,In_153);
or U529 (N_529,In_1118,In_1684);
or U530 (N_530,In_122,In_1609);
and U531 (N_531,In_977,In_1851);
nand U532 (N_532,In_1127,In_95);
nand U533 (N_533,In_1140,In_815);
and U534 (N_534,In_2474,In_2431);
nor U535 (N_535,In_1422,In_2253);
nand U536 (N_536,In_621,In_1202);
nor U537 (N_537,In_1100,In_2370);
and U538 (N_538,In_1754,In_62);
nand U539 (N_539,In_515,In_1109);
nor U540 (N_540,In_761,In_2428);
xor U541 (N_541,In_1717,In_2180);
and U542 (N_542,In_1795,In_1800);
or U543 (N_543,In_670,In_837);
nor U544 (N_544,In_1816,In_1736);
nor U545 (N_545,In_901,In_835);
or U546 (N_546,In_1857,In_983);
nor U547 (N_547,In_310,In_1844);
or U548 (N_548,In_1356,In_540);
and U549 (N_549,In_2311,In_2074);
or U550 (N_550,In_442,In_1827);
nor U551 (N_551,In_1836,In_220);
and U552 (N_552,In_2205,In_2029);
nand U553 (N_553,In_42,In_330);
nand U554 (N_554,In_1312,In_986);
or U555 (N_555,In_40,In_829);
and U556 (N_556,In_2491,In_613);
and U557 (N_557,In_1151,In_1999);
nand U558 (N_558,In_2479,In_950);
and U559 (N_559,In_313,In_589);
nand U560 (N_560,In_1371,In_1794);
nor U561 (N_561,In_2395,In_1969);
and U562 (N_562,In_2236,In_992);
nand U563 (N_563,In_1466,In_1762);
xnor U564 (N_564,In_1884,In_2489);
or U565 (N_565,In_1130,In_1472);
or U566 (N_566,In_1053,In_2440);
nand U567 (N_567,In_244,In_505);
xnor U568 (N_568,In_889,In_1298);
and U569 (N_569,In_2041,In_126);
nand U570 (N_570,In_1594,In_513);
nand U571 (N_571,In_110,In_974);
nand U572 (N_572,In_1033,In_1364);
or U573 (N_573,In_1752,In_1854);
or U574 (N_574,In_2185,In_2168);
nand U575 (N_575,In_1005,In_1102);
nand U576 (N_576,In_642,In_298);
xor U577 (N_577,In_897,In_2366);
nor U578 (N_578,In_919,In_736);
or U579 (N_579,In_1317,In_1965);
nand U580 (N_580,In_2464,In_550);
xor U581 (N_581,In_760,In_2478);
nor U582 (N_582,In_1935,In_874);
and U583 (N_583,In_1016,In_1520);
and U584 (N_584,In_643,In_898);
nor U585 (N_585,In_159,In_1435);
nor U586 (N_586,In_1026,In_547);
nand U587 (N_587,In_1500,In_2348);
or U588 (N_588,In_1394,In_1262);
or U589 (N_589,In_1421,In_866);
nor U590 (N_590,In_916,In_444);
nor U591 (N_591,In_225,In_1747);
and U592 (N_592,In_381,In_2107);
nor U593 (N_593,In_47,In_795);
or U594 (N_594,In_1123,In_1439);
and U595 (N_595,In_1399,In_1895);
nand U596 (N_596,In_1170,In_1721);
nor U597 (N_597,In_1756,In_152);
or U598 (N_598,In_395,In_1845);
nand U599 (N_599,In_741,In_1832);
nor U600 (N_600,In_1751,In_2410);
nor U601 (N_601,In_76,In_664);
nand U602 (N_602,In_2429,In_1081);
nand U603 (N_603,In_1994,In_2182);
and U604 (N_604,In_1431,In_71);
nor U605 (N_605,In_1838,In_1322);
nor U606 (N_606,In_1823,In_1309);
and U607 (N_607,In_1507,In_923);
xor U608 (N_608,In_605,In_1488);
and U609 (N_609,In_1749,In_2083);
nand U610 (N_610,In_2239,In_296);
or U611 (N_611,In_2267,In_1995);
nand U612 (N_612,In_2122,In_1989);
and U613 (N_613,In_1651,In_2026);
or U614 (N_614,In_335,In_1911);
nor U615 (N_615,In_83,In_1964);
nor U616 (N_616,In_1071,In_894);
and U617 (N_617,In_1913,In_720);
nor U618 (N_618,In_481,In_2299);
nand U619 (N_619,In_512,In_1125);
or U620 (N_620,In_527,In_1842);
or U621 (N_621,In_301,In_1958);
nor U622 (N_622,In_1362,In_2488);
and U623 (N_623,In_502,In_454);
and U624 (N_624,In_538,In_409);
nand U625 (N_625,In_946,In_2495);
nor U626 (N_626,In_419,In_801);
nand U627 (N_627,In_1896,In_1160);
and U628 (N_628,In_338,In_85);
nand U629 (N_629,In_2254,In_2262);
nand U630 (N_630,In_12,In_1129);
or U631 (N_631,In_1986,In_947);
nand U632 (N_632,In_745,In_208);
nor U633 (N_633,In_2017,In_463);
xor U634 (N_634,In_2394,In_845);
or U635 (N_635,In_1474,In_91);
nor U636 (N_636,In_1035,In_2141);
nor U637 (N_637,In_1960,In_1190);
nand U638 (N_638,In_155,In_1242);
xnor U639 (N_639,In_428,In_1779);
or U640 (N_640,In_1434,In_1284);
or U641 (N_641,In_2298,In_1981);
xor U642 (N_642,In_1136,In_1383);
nor U643 (N_643,In_174,In_1283);
nor U644 (N_644,In_1618,In_431);
and U645 (N_645,In_1301,In_738);
or U646 (N_646,In_434,In_459);
or U647 (N_647,In_1727,In_2292);
nand U648 (N_648,In_2396,In_746);
nor U649 (N_649,In_20,In_2467);
nor U650 (N_650,In_1040,In_492);
and U651 (N_651,In_316,In_1834);
or U652 (N_652,In_1880,In_2258);
nor U653 (N_653,In_1649,In_2391);
and U654 (N_654,In_1849,In_1548);
nand U655 (N_655,In_2015,In_73);
or U656 (N_656,In_1173,In_1907);
xor U657 (N_657,In_1776,In_1511);
nand U658 (N_658,In_1230,In_1360);
and U659 (N_659,In_765,In_2213);
or U660 (N_660,In_1323,In_1084);
or U661 (N_661,In_647,In_339);
nand U662 (N_662,In_1764,In_1122);
and U663 (N_663,In_2250,In_2336);
xor U664 (N_664,In_1628,In_396);
nand U665 (N_665,In_2330,In_2092);
nor U666 (N_666,In_706,In_52);
and U667 (N_667,In_1581,In_457);
or U668 (N_668,In_1726,In_535);
or U669 (N_669,In_169,In_2285);
nor U670 (N_670,In_616,In_295);
nor U671 (N_671,In_1479,In_1606);
and U672 (N_672,In_1297,In_1728);
nor U673 (N_673,In_1338,In_315);
nor U674 (N_674,In_504,In_786);
nor U675 (N_675,In_1487,In_369);
xnor U676 (N_676,In_1659,In_2163);
nor U677 (N_677,In_566,In_2006);
or U678 (N_678,In_1111,In_267);
nand U679 (N_679,In_1925,In_1042);
or U680 (N_680,In_1034,In_2420);
or U681 (N_681,In_639,In_2244);
xor U682 (N_682,In_1596,In_1222);
nor U683 (N_683,In_235,In_2264);
nand U684 (N_684,In_494,In_1929);
nor U685 (N_685,In_991,In_1517);
xor U686 (N_686,In_2005,In_2408);
xnor U687 (N_687,In_680,In_1855);
nand U688 (N_688,In_204,In_2329);
nor U689 (N_689,In_1121,In_1104);
nor U690 (N_690,In_629,In_2162);
xnor U691 (N_691,In_2457,In_1510);
nand U692 (N_692,In_2064,In_1402);
and U693 (N_693,In_1384,In_1428);
nor U694 (N_694,In_2494,In_1117);
nor U695 (N_695,In_632,In_2111);
nand U696 (N_696,In_734,In_1382);
and U697 (N_697,In_996,In_753);
nor U698 (N_698,In_2369,In_1938);
and U699 (N_699,In_1147,In_1982);
or U700 (N_700,In_660,In_1616);
xor U701 (N_701,In_1157,In_2397);
or U702 (N_702,In_577,In_1021);
and U703 (N_703,In_374,In_1194);
or U704 (N_704,In_1266,In_1739);
or U705 (N_705,In_603,In_931);
xor U706 (N_706,In_1828,In_1475);
or U707 (N_707,In_1593,In_559);
nor U708 (N_708,In_1588,In_104);
and U709 (N_709,In_1619,In_1590);
or U710 (N_710,In_1450,In_662);
or U711 (N_711,In_2327,In_1706);
nand U712 (N_712,In_1216,In_683);
nor U713 (N_713,In_1876,In_203);
or U714 (N_714,In_1305,In_2416);
or U715 (N_715,In_2376,In_970);
nor U716 (N_716,In_869,In_2047);
nand U717 (N_717,In_336,In_1247);
nor U718 (N_718,In_488,In_2098);
nor U719 (N_719,In_868,In_290);
or U720 (N_720,In_2349,In_2178);
nand U721 (N_721,In_1586,In_2284);
nor U722 (N_722,In_21,In_1172);
and U723 (N_723,In_1519,In_1978);
and U724 (N_724,In_1405,In_1473);
and U725 (N_725,In_690,In_1336);
or U726 (N_726,In_909,In_693);
nand U727 (N_727,In_1796,In_582);
or U728 (N_728,In_2039,In_1977);
nand U729 (N_729,In_38,In_709);
nor U730 (N_730,In_819,In_2287);
nand U731 (N_731,In_1692,In_364);
or U732 (N_732,In_346,In_708);
xor U733 (N_733,In_1198,In_802);
nor U734 (N_734,In_1031,In_1306);
or U735 (N_735,In_811,In_1452);
nor U736 (N_736,In_688,In_964);
and U737 (N_737,In_1947,In_2104);
and U738 (N_738,In_1375,In_562);
nand U739 (N_739,In_406,In_836);
nand U740 (N_740,In_2219,In_520);
nor U741 (N_741,In_989,In_1060);
nor U742 (N_742,In_1627,In_415);
nand U743 (N_743,In_186,In_448);
xor U744 (N_744,In_2481,In_1710);
and U745 (N_745,In_1243,In_2102);
or U746 (N_746,In_397,In_1589);
nand U747 (N_747,In_1400,In_948);
or U748 (N_748,In_1062,In_484);
or U749 (N_749,In_273,In_518);
and U750 (N_750,In_2200,In_933);
nor U751 (N_751,In_2470,In_2273);
and U752 (N_752,In_255,In_281);
and U753 (N_753,In_376,In_998);
and U754 (N_754,In_1670,In_754);
nand U755 (N_755,In_921,In_1766);
nor U756 (N_756,In_1950,In_1376);
xor U757 (N_757,In_304,In_1826);
or U758 (N_758,In_920,In_1106);
and U759 (N_759,In_620,In_1813);
nor U760 (N_760,In_2030,In_343);
and U761 (N_761,In_1469,In_2194);
or U762 (N_762,In_124,In_401);
and U763 (N_763,In_189,In_2455);
or U764 (N_764,In_2375,In_286);
nor U765 (N_765,In_1091,In_1918);
nand U766 (N_766,In_2062,In_2436);
nand U767 (N_767,In_1056,In_1390);
or U768 (N_768,In_2344,In_1987);
nor U769 (N_769,In_1398,In_1809);
xor U770 (N_770,In_2212,In_2268);
xnor U771 (N_771,In_2190,In_814);
and U772 (N_772,In_1601,In_1653);
and U773 (N_773,In_1729,In_1436);
xnor U774 (N_774,In_1614,In_115);
nand U775 (N_775,In_1381,In_2434);
nand U776 (N_776,In_166,In_402);
nand U777 (N_777,In_2049,In_1401);
nor U778 (N_778,In_1482,In_67);
nor U779 (N_779,In_2320,In_350);
xnor U780 (N_780,In_1534,In_2484);
and U781 (N_781,In_1107,In_2089);
or U782 (N_782,In_833,In_256);
or U783 (N_783,In_1263,In_1285);
or U784 (N_784,In_1971,In_529);
nand U785 (N_785,In_1934,In_287);
and U786 (N_786,In_2166,In_438);
nor U787 (N_787,In_1904,In_560);
nor U788 (N_788,In_640,In_1244);
and U789 (N_789,In_1008,In_1516);
nand U790 (N_790,In_26,In_2226);
and U791 (N_791,In_2191,In_326);
nor U792 (N_792,In_2450,In_2132);
or U793 (N_793,In_1404,In_327);
and U794 (N_794,In_5,In_615);
xor U795 (N_795,In_150,In_187);
and U796 (N_796,In_687,In_704);
and U797 (N_797,In_1580,In_756);
and U798 (N_798,In_113,In_332);
xor U799 (N_799,In_707,In_1006);
nand U800 (N_800,In_1932,In_2101);
xnor U801 (N_801,In_384,In_758);
nand U802 (N_802,In_53,In_1447);
and U803 (N_803,In_972,In_1019);
nor U804 (N_804,In_762,In_2001);
and U805 (N_805,In_1272,In_1574);
or U806 (N_806,In_2345,In_323);
and U807 (N_807,In_2188,In_92);
and U808 (N_808,In_2334,In_564);
and U809 (N_809,In_1069,In_2425);
or U810 (N_810,In_2445,In_2317);
nand U811 (N_811,In_2310,In_116);
nor U812 (N_812,In_604,In_631);
or U813 (N_813,In_1738,In_1817);
or U814 (N_814,In_883,In_59);
nor U815 (N_815,In_1485,In_1457);
xnor U816 (N_816,In_587,In_1974);
xor U817 (N_817,In_712,In_377);
nor U818 (N_818,In_417,In_864);
and U819 (N_819,In_1654,In_750);
nand U820 (N_820,In_788,In_1493);
and U821 (N_821,In_1819,In_1289);
nor U822 (N_822,In_1953,In_506);
nand U823 (N_823,In_387,In_1017);
or U824 (N_824,In_143,In_1391);
nor U825 (N_825,In_379,In_2487);
and U826 (N_826,In_1785,In_957);
or U827 (N_827,In_2,In_617);
nor U828 (N_828,In_1214,In_1630);
nor U829 (N_829,In_987,In_2033);
nand U830 (N_830,In_1731,In_1453);
nor U831 (N_831,In_1483,In_925);
nor U832 (N_832,In_793,In_1624);
nand U833 (N_833,In_490,In_1278);
and U834 (N_834,In_1543,In_716);
or U835 (N_835,In_551,In_1686);
nor U836 (N_836,In_1271,In_132);
and U837 (N_837,In_239,In_44);
nand U838 (N_838,In_1879,In_1810);
and U839 (N_839,In_1555,In_1532);
or U840 (N_840,In_1617,In_2364);
and U841 (N_841,In_2312,In_1585);
xor U842 (N_842,In_36,In_1145);
nor U843 (N_843,In_146,In_2137);
or U844 (N_844,In_857,In_1553);
or U845 (N_845,In_1086,In_548);
nand U846 (N_846,In_1154,In_1199);
nand U847 (N_847,In_650,In_1440);
or U848 (N_848,In_600,In_2451);
nand U849 (N_849,In_2164,In_2257);
and U850 (N_850,In_580,In_1967);
or U851 (N_851,In_700,In_2490);
nor U852 (N_852,In_2454,In_1564);
and U853 (N_853,In_1187,In_388);
or U854 (N_854,In_1128,In_2227);
xnor U855 (N_855,In_263,In_1791);
nor U856 (N_856,In_873,In_1696);
xor U857 (N_857,In_1408,In_202);
or U858 (N_858,In_2483,In_1430);
and U859 (N_859,In_254,In_1648);
nand U860 (N_860,In_1417,In_1184);
or U861 (N_861,In_1380,In_576);
nor U862 (N_862,In_1233,In_1883);
and U863 (N_863,In_1282,In_1632);
and U864 (N_864,In_980,In_1088);
nand U865 (N_865,In_681,In_129);
nor U866 (N_866,In_1411,In_285);
and U867 (N_867,In_588,In_1513);
nor U868 (N_868,In_657,In_1287);
nor U869 (N_869,In_1204,In_813);
nor U870 (N_870,In_368,In_2100);
or U871 (N_871,In_884,In_2075);
and U872 (N_872,In_93,In_2248);
nand U873 (N_873,In_840,In_325);
nor U874 (N_874,In_48,In_1097);
or U875 (N_875,In_2153,In_1037);
nand U876 (N_876,In_252,In_420);
or U877 (N_877,In_1281,In_1024);
nand U878 (N_878,In_939,In_2177);
nor U879 (N_879,In_752,In_796);
nor U880 (N_880,In_1655,In_1542);
and U881 (N_881,In_497,In_405);
and U882 (N_882,In_158,In_1662);
nor U883 (N_883,In_170,In_1218);
nor U884 (N_884,In_78,In_2300);
or U885 (N_885,In_11,In_578);
nand U886 (N_886,In_2302,In_804);
or U887 (N_887,In_1224,In_1229);
nand U888 (N_888,In_191,In_653);
and U889 (N_889,In_1171,In_2492);
nand U890 (N_890,In_1843,In_1315);
nor U891 (N_891,In_521,In_373);
nor U892 (N_892,In_2105,In_2472);
nor U893 (N_893,In_2423,In_418);
nor U894 (N_894,In_2139,In_2038);
or U895 (N_895,In_1134,In_1462);
xnor U896 (N_896,In_955,In_119);
or U897 (N_897,In_1862,In_265);
or U898 (N_898,In_2406,In_1980);
and U899 (N_899,In_1970,In_1211);
and U900 (N_900,In_1092,In_1048);
nor U901 (N_901,In_2313,In_1094);
nand U902 (N_902,In_2368,In_1502);
and U903 (N_903,In_1131,In_755);
and U904 (N_904,In_661,In_2120);
nor U905 (N_905,In_701,In_2407);
and U906 (N_906,In_270,In_1642);
nor U907 (N_907,In_1900,In_543);
or U908 (N_908,In_1940,In_654);
or U909 (N_909,In_1409,In_1612);
and U910 (N_910,In_1976,In_1438);
and U911 (N_911,In_230,In_2326);
nand U912 (N_912,In_737,In_1248);
and U913 (N_913,In_274,In_278);
nor U914 (N_914,In_1217,In_1508);
nand U915 (N_915,In_2333,In_1352);
nand U916 (N_916,In_2449,In_1427);
nand U917 (N_917,In_188,In_575);
xnor U918 (N_918,In_1395,In_2077);
nor U919 (N_919,In_1221,In_1626);
and U920 (N_920,In_1509,In_2146);
and U921 (N_921,In_2278,In_1054);
nor U922 (N_922,In_201,In_2392);
or U923 (N_923,In_2281,In_2130);
xnor U924 (N_924,In_710,In_1484);
or U925 (N_925,In_665,In_1114);
and U926 (N_926,In_192,In_277);
nor U927 (N_927,In_1495,In_1783);
and U928 (N_928,In_1014,In_2156);
nand U929 (N_929,In_985,In_1001);
xnor U930 (N_930,In_2441,In_914);
and U931 (N_931,In_1815,In_248);
xnor U932 (N_932,In_2093,In_1853);
or U933 (N_933,In_199,In_1968);
xor U934 (N_934,In_2409,In_2465);
and U935 (N_935,In_1470,In_1180);
nor U936 (N_936,In_2097,In_100);
or U937 (N_937,In_2158,In_173);
nand U938 (N_938,In_1497,In_391);
or U939 (N_939,In_2086,In_855);
and U940 (N_940,In_2043,In_45);
nor U941 (N_941,In_359,In_1867);
and U942 (N_942,In_2361,In_1164);
nor U943 (N_943,In_1830,In_1841);
nor U944 (N_944,In_2321,In_1899);
or U945 (N_945,In_1615,In_2019);
or U946 (N_946,In_1207,In_585);
nand U947 (N_947,In_1786,In_1910);
or U948 (N_948,In_1620,In_1525);
xor U949 (N_949,In_1708,In_685);
nand U950 (N_950,In_1159,In_123);
nand U951 (N_951,In_2399,In_1412);
or U952 (N_952,In_1231,In_2128);
xor U953 (N_953,In_1389,In_261);
xnor U954 (N_954,In_1582,In_1949);
and U955 (N_955,In_808,In_2087);
nand U956 (N_956,In_1476,In_544);
or U957 (N_957,In_1886,In_1789);
or U958 (N_958,In_219,In_522);
or U959 (N_959,In_2027,In_1023);
nor U960 (N_960,In_1656,In_361);
nor U961 (N_961,In_1750,In_1530);
nor U962 (N_962,In_1432,In_554);
nand U963 (N_963,In_1825,In_1770);
xor U964 (N_964,In_233,In_994);
nand U965 (N_965,In_1445,In_651);
and U966 (N_966,In_853,In_1108);
nand U967 (N_967,In_30,In_1388);
nor U968 (N_968,In_1461,In_1865);
nand U969 (N_969,In_2424,In_74);
nor U970 (N_970,In_2037,In_1592);
or U971 (N_971,In_545,In_1637);
nor U972 (N_972,In_960,In_112);
nor U973 (N_973,In_441,In_1459);
or U974 (N_974,In_1250,In_23);
nor U975 (N_975,In_2274,In_944);
xor U976 (N_976,In_1544,In_730);
nor U977 (N_977,In_2466,In_789);
and U978 (N_978,In_1050,In_1861);
xnor U979 (N_979,In_1148,In_703);
and U980 (N_980,In_1032,In_1074);
nor U981 (N_981,In_1631,In_245);
nor U982 (N_982,In_2013,In_2129);
and U983 (N_983,In_1255,In_1288);
nand U984 (N_984,In_2400,In_288);
nand U985 (N_985,In_2456,In_1093);
or U986 (N_986,In_2218,In_164);
and U987 (N_987,In_878,In_769);
nand U988 (N_988,In_1013,In_1571);
nand U989 (N_989,In_1835,In_151);
nor U990 (N_990,In_2372,In_2140);
nand U991 (N_991,In_912,In_1098);
nand U992 (N_992,In_179,In_1583);
or U993 (N_993,In_181,In_1146);
or U994 (N_994,In_193,In_2272);
and U995 (N_995,In_196,In_1997);
or U996 (N_996,In_1863,In_1733);
and U997 (N_997,In_637,In_774);
or U998 (N_998,In_1512,In_1039);
nand U999 (N_999,In_2339,In_764);
nor U1000 (N_1000,In_232,In_1643);
nand U1001 (N_1001,In_1923,In_1348);
nor U1002 (N_1002,In_780,In_1933);
or U1003 (N_1003,In_88,In_56);
nand U1004 (N_1004,In_995,In_427);
or U1005 (N_1005,In_2024,In_1963);
xnor U1006 (N_1006,In_1573,In_810);
nand U1007 (N_1007,In_125,In_1939);
and U1008 (N_1008,In_2136,In_888);
xor U1009 (N_1009,In_1419,In_1859);
nand U1010 (N_1010,In_2079,In_430);
and U1011 (N_1011,In_29,In_1683);
nand U1012 (N_1012,In_1941,In_1072);
nor U1013 (N_1013,In_383,In_218);
nand U1014 (N_1014,In_2263,In_1811);
xor U1015 (N_1015,In_1658,In_117);
xor U1016 (N_1016,In_626,In_1799);
nand U1017 (N_1017,In_435,In_2012);
xnor U1018 (N_1018,In_1645,In_1051);
or U1019 (N_1019,In_165,In_768);
nor U1020 (N_1020,In_2241,In_1561);
and U1021 (N_1021,In_55,In_19);
nand U1022 (N_1022,In_1503,In_81);
and U1023 (N_1023,In_1418,In_1711);
xnor U1024 (N_1024,In_557,In_1539);
nand U1025 (N_1025,In_1885,In_466);
and U1026 (N_1026,In_2203,In_1406);
and U1027 (N_1027,In_1201,In_72);
or U1028 (N_1028,In_1758,In_1852);
xor U1029 (N_1029,In_32,In_2390);
nor U1030 (N_1030,In_1183,In_659);
nand U1031 (N_1031,In_610,In_1279);
and U1032 (N_1032,In_2152,In_1860);
nor U1033 (N_1033,In_135,In_386);
xnor U1034 (N_1034,In_771,In_2204);
xor U1035 (N_1035,In_881,In_830);
nand U1036 (N_1036,In_1792,In_318);
nor U1037 (N_1037,In_1294,In_107);
nand U1038 (N_1038,In_8,In_1273);
nand U1039 (N_1039,In_1806,In_1666);
or U1040 (N_1040,In_1293,In_1413);
and U1041 (N_1041,In_1365,In_185);
nand U1042 (N_1042,In_118,In_111);
nor U1043 (N_1043,In_825,In_1808);
nor U1044 (N_1044,In_50,In_2127);
and U1045 (N_1045,In_149,In_940);
and U1046 (N_1046,In_812,In_1345);
nand U1047 (N_1047,In_87,In_1536);
and U1048 (N_1048,In_594,In_108);
or U1049 (N_1049,In_697,In_784);
nand U1050 (N_1050,In_532,In_94);
and U1051 (N_1051,In_334,In_1866);
or U1052 (N_1052,In_1491,In_2011);
nand U1053 (N_1053,In_136,In_1478);
nor U1054 (N_1054,In_2118,In_890);
xnor U1055 (N_1055,In_500,In_31);
nand U1056 (N_1056,In_773,In_779);
or U1057 (N_1057,In_1423,In_2073);
and U1058 (N_1058,In_1009,In_416);
xnor U1059 (N_1059,In_847,In_1073);
and U1060 (N_1060,In_959,In_1377);
nor U1061 (N_1061,In_1142,In_1064);
or U1062 (N_1062,In_412,In_1526);
and U1063 (N_1063,In_1410,In_2134);
or U1064 (N_1064,In_2051,In_1712);
xor U1065 (N_1065,In_2293,In_581);
nand U1066 (N_1066,In_820,In_1464);
nand U1067 (N_1067,In_2338,In_591);
and U1068 (N_1068,In_2382,In_1768);
and U1069 (N_1069,In_1022,In_291);
nand U1070 (N_1070,In_1782,In_1358);
nor U1071 (N_1071,In_2332,In_272);
nand U1072 (N_1072,In_1887,In_2044);
xor U1073 (N_1073,In_1120,In_356);
and U1074 (N_1074,In_1049,In_1261);
nand U1075 (N_1075,In_1531,In_39);
and U1076 (N_1076,In_453,In_28);
nand U1077 (N_1077,In_1152,In_1674);
nor U1078 (N_1078,In_66,In_1673);
nor U1079 (N_1079,In_831,In_1694);
and U1080 (N_1080,In_222,In_80);
nand U1081 (N_1081,In_1295,In_2022);
or U1082 (N_1082,In_2010,In_1124);
xnor U1083 (N_1083,In_1535,In_1238);
nor U1084 (N_1084,In_485,In_1426);
nand U1085 (N_1085,In_2216,In_666);
nand U1086 (N_1086,In_1200,In_14);
nor U1087 (N_1087,In_1587,In_1657);
and U1088 (N_1088,In_1898,In_1897);
nand U1089 (N_1089,In_483,In_1078);
nand U1090 (N_1090,In_2036,In_537);
and U1091 (N_1091,In_456,In_1797);
or U1092 (N_1092,In_1985,In_344);
or U1093 (N_1093,In_1156,In_280);
xnor U1094 (N_1094,In_1029,In_1350);
and U1095 (N_1095,In_2245,In_990);
nand U1096 (N_1096,In_1334,In_1275);
and U1097 (N_1097,In_976,In_684);
or U1098 (N_1098,In_910,In_2103);
nand U1099 (N_1099,In_679,In_900);
or U1100 (N_1100,In_1369,In_1537);
nor U1101 (N_1101,In_2269,In_2143);
or U1102 (N_1102,In_228,In_1952);
nand U1103 (N_1103,In_1236,In_200);
nand U1104 (N_1104,In_598,In_2430);
and U1105 (N_1105,In_207,In_1067);
nor U1106 (N_1106,In_246,In_1132);
nor U1107 (N_1107,In_367,In_2050);
or U1108 (N_1108,In_1496,In_1990);
or U1109 (N_1109,In_748,In_147);
or U1110 (N_1110,In_865,In_2048);
or U1111 (N_1111,In_1007,In_862);
or U1112 (N_1112,In_1327,In_1873);
or U1113 (N_1113,In_1875,In_1477);
nor U1114 (N_1114,In_1912,In_1372);
xor U1115 (N_1115,In_732,In_733);
xnor U1116 (N_1116,In_2458,In_70);
and U1117 (N_1117,In_1249,In_495);
or U1118 (N_1118,In_822,In_353);
or U1119 (N_1119,In_1002,In_103);
nand U1120 (N_1120,In_275,In_231);
xnor U1121 (N_1121,In_2004,In_46);
or U1122 (N_1122,In_1429,In_1905);
xor U1123 (N_1123,In_1045,In_797);
and U1124 (N_1124,In_1174,In_586);
or U1125 (N_1125,In_2207,In_511);
nand U1126 (N_1126,In_982,In_90);
nor U1127 (N_1127,In_355,In_2398);
nor U1128 (N_1128,In_1055,In_556);
nor U1129 (N_1129,In_770,In_2065);
nand U1130 (N_1130,In_1916,In_2184);
nand U1131 (N_1131,In_141,In_2421);
or U1132 (N_1132,In_337,In_1252);
xor U1133 (N_1133,In_1280,In_212);
or U1134 (N_1134,In_468,In_2059);
or U1135 (N_1135,In_2008,In_1228);
nand U1136 (N_1136,In_1304,In_1003);
and U1137 (N_1137,In_717,In_1443);
or U1138 (N_1138,In_1988,In_507);
or U1139 (N_1139,In_322,In_1681);
nor U1140 (N_1140,In_2418,In_776);
nor U1141 (N_1141,In_1256,In_850);
nor U1142 (N_1142,In_389,In_407);
or U1143 (N_1143,In_1260,In_2189);
nand U1144 (N_1144,In_524,In_1699);
or U1145 (N_1145,In_27,In_1246);
nand U1146 (N_1146,In_455,In_1155);
and U1147 (N_1147,In_892,In_533);
nor U1148 (N_1148,In_1757,In_602);
and U1149 (N_1149,In_1353,In_2459);
nor U1150 (N_1150,In_2347,In_314);
nor U1151 (N_1151,In_519,In_498);
or U1152 (N_1152,In_2291,In_1359);
and U1153 (N_1153,In_358,In_247);
nand U1154 (N_1154,In_2070,In_1533);
nand U1155 (N_1155,In_349,In_329);
nand U1156 (N_1156,In_711,In_501);
or U1157 (N_1157,In_2088,In_744);
nand U1158 (N_1158,In_2160,In_168);
and U1159 (N_1159,In_918,In_880);
and U1160 (N_1160,In_584,In_999);
or U1161 (N_1161,In_913,In_2198);
nand U1162 (N_1162,In_2056,In_809);
nor U1163 (N_1163,In_973,In_133);
and U1164 (N_1164,In_1882,In_411);
and U1165 (N_1165,In_1877,In_65);
xor U1166 (N_1166,In_1501,In_1166);
nand U1167 (N_1167,In_1105,In_2023);
or U1168 (N_1168,In_723,In_404);
and U1169 (N_1169,In_1597,In_2147);
nand U1170 (N_1170,In_2231,In_1219);
or U1171 (N_1171,In_1821,In_1209);
nand U1172 (N_1172,In_1704,In_834);
nor U1173 (N_1173,In_1442,In_1570);
or U1174 (N_1174,In_447,In_2233);
or U1175 (N_1175,In_259,In_423);
or U1176 (N_1176,In_2230,In_1363);
nand U1177 (N_1177,In_82,In_628);
nand U1178 (N_1178,In_929,In_1341);
nor U1179 (N_1179,In_1387,In_2142);
nor U1180 (N_1180,In_1771,In_9);
or U1181 (N_1181,In_224,In_907);
or U1182 (N_1182,In_1798,In_806);
nand U1183 (N_1183,In_209,In_2071);
nand U1184 (N_1184,In_747,In_2443);
nand U1185 (N_1185,In_2215,In_1636);
nor U1186 (N_1186,In_172,In_63);
nand U1187 (N_1187,In_1137,In_2363);
xor U1188 (N_1188,In_2210,In_2371);
or U1189 (N_1189,In_1944,In_676);
nand U1190 (N_1190,In_1629,In_1112);
nor U1191 (N_1191,In_1961,In_536);
and U1192 (N_1192,In_1165,In_1975);
xnor U1193 (N_1193,In_243,In_2149);
nor U1194 (N_1194,In_2301,In_1741);
and U1195 (N_1195,In_1324,In_1663);
nand U1196 (N_1196,In_1942,In_714);
and U1197 (N_1197,In_635,In_2360);
nor U1198 (N_1198,In_1719,In_1378);
nor U1199 (N_1199,In_1357,In_134);
and U1200 (N_1200,In_903,In_1258);
nand U1201 (N_1201,In_303,In_1254);
nor U1202 (N_1202,In_160,In_1962);
nor U1203 (N_1203,In_1212,In_137);
and U1204 (N_1204,In_422,In_482);
nor U1205 (N_1205,In_599,In_694);
nand U1206 (N_1206,In_508,In_1959);
and U1207 (N_1207,In_1044,In_114);
and U1208 (N_1208,In_1433,In_1635);
nor U1209 (N_1209,In_691,In_938);
nor U1210 (N_1210,In_1090,In_2009);
nand U1211 (N_1211,In_1927,In_1556);
nor U1212 (N_1212,In_308,In_2099);
nor U1213 (N_1213,In_1558,In_1274);
and U1214 (N_1214,In_2199,In_503);
nor U1215 (N_1215,In_493,In_1992);
or U1216 (N_1216,In_1893,In_1489);
and U1217 (N_1217,In_1577,In_229);
and U1218 (N_1218,In_269,In_895);
nor U1219 (N_1219,In_293,In_1471);
nand U1220 (N_1220,In_1915,In_1087);
or U1221 (N_1221,In_340,In_394);
nor U1222 (N_1222,In_1268,In_2171);
and U1223 (N_1223,In_464,In_826);
or U1224 (N_1224,In_781,In_937);
xor U1225 (N_1225,In_439,In_649);
or U1226 (N_1226,In_467,In_2426);
nand U1227 (N_1227,In_614,In_563);
nor U1228 (N_1228,In_682,In_1833);
xor U1229 (N_1229,In_1767,In_446);
xor U1230 (N_1230,In_2414,In_843);
or U1231 (N_1231,In_96,In_471);
or U1232 (N_1232,In_2135,In_823);
nand U1233 (N_1233,In_1308,In_1780);
or U1234 (N_1234,In_2192,In_2221);
or U1235 (N_1235,In_722,In_440);
or U1236 (N_1236,In_2229,In_1946);
and U1237 (N_1237,In_1220,In_1015);
nand U1238 (N_1238,In_2238,In_1515);
nand U1239 (N_1239,In_1891,In_217);
or U1240 (N_1240,In_89,In_705);
or U1241 (N_1241,In_1059,In_728);
xnor U1242 (N_1242,In_2306,In_1820);
nor U1243 (N_1243,In_611,In_2154);
nor U1244 (N_1244,In_283,In_574);
and U1245 (N_1245,In_2452,In_785);
nand U1246 (N_1246,In_1150,In_848);
nor U1247 (N_1247,In_1319,In_2383);
and U1248 (N_1248,In_1701,In_380);
and U1249 (N_1249,In_1070,In_1113);
nand U1250 (N_1250,In_1657,In_2315);
nand U1251 (N_1251,In_981,In_878);
and U1252 (N_1252,In_2147,In_2018);
nor U1253 (N_1253,In_1184,In_678);
nand U1254 (N_1254,In_2086,In_1220);
nor U1255 (N_1255,In_2355,In_1128);
and U1256 (N_1256,In_221,In_2439);
xor U1257 (N_1257,In_1600,In_1538);
and U1258 (N_1258,In_2048,In_2044);
xor U1259 (N_1259,In_1640,In_1976);
nor U1260 (N_1260,In_97,In_515);
or U1261 (N_1261,In_164,In_2111);
and U1262 (N_1262,In_2457,In_2189);
nand U1263 (N_1263,In_1436,In_304);
nand U1264 (N_1264,In_105,In_41);
or U1265 (N_1265,In_1488,In_556);
nor U1266 (N_1266,In_1952,In_582);
or U1267 (N_1267,In_389,In_41);
nand U1268 (N_1268,In_1494,In_1351);
and U1269 (N_1269,In_1298,In_1442);
nor U1270 (N_1270,In_2442,In_2050);
or U1271 (N_1271,In_929,In_398);
nand U1272 (N_1272,In_614,In_1159);
and U1273 (N_1273,In_1754,In_1453);
nand U1274 (N_1274,In_2438,In_1034);
nor U1275 (N_1275,In_1511,In_1938);
nor U1276 (N_1276,In_2,In_1395);
or U1277 (N_1277,In_437,In_2439);
and U1278 (N_1278,In_2006,In_1584);
and U1279 (N_1279,In_438,In_2090);
or U1280 (N_1280,In_1207,In_1308);
nor U1281 (N_1281,In_297,In_461);
and U1282 (N_1282,In_392,In_2328);
nand U1283 (N_1283,In_1434,In_2471);
nand U1284 (N_1284,In_2310,In_1265);
or U1285 (N_1285,In_439,In_1696);
nor U1286 (N_1286,In_2398,In_754);
nand U1287 (N_1287,In_2019,In_11);
nor U1288 (N_1288,In_1860,In_36);
nor U1289 (N_1289,In_2438,In_58);
or U1290 (N_1290,In_1260,In_2031);
nor U1291 (N_1291,In_1048,In_292);
nor U1292 (N_1292,In_1367,In_1759);
nand U1293 (N_1293,In_314,In_43);
xor U1294 (N_1294,In_1393,In_2045);
nand U1295 (N_1295,In_1410,In_1221);
nor U1296 (N_1296,In_961,In_572);
and U1297 (N_1297,In_1153,In_326);
or U1298 (N_1298,In_911,In_2074);
and U1299 (N_1299,In_2196,In_562);
nand U1300 (N_1300,In_1777,In_189);
nor U1301 (N_1301,In_1927,In_1138);
nand U1302 (N_1302,In_2158,In_2008);
nor U1303 (N_1303,In_2004,In_1864);
nand U1304 (N_1304,In_443,In_932);
nand U1305 (N_1305,In_1506,In_993);
or U1306 (N_1306,In_213,In_1918);
and U1307 (N_1307,In_41,In_784);
nor U1308 (N_1308,In_107,In_1515);
or U1309 (N_1309,In_1713,In_1491);
or U1310 (N_1310,In_1314,In_2251);
nor U1311 (N_1311,In_2146,In_2185);
and U1312 (N_1312,In_804,In_731);
or U1313 (N_1313,In_2260,In_599);
and U1314 (N_1314,In_896,In_527);
nand U1315 (N_1315,In_2327,In_1610);
or U1316 (N_1316,In_1879,In_1372);
xor U1317 (N_1317,In_1089,In_813);
and U1318 (N_1318,In_1670,In_2214);
or U1319 (N_1319,In_2100,In_2101);
xnor U1320 (N_1320,In_102,In_177);
and U1321 (N_1321,In_638,In_754);
and U1322 (N_1322,In_1485,In_2124);
nor U1323 (N_1323,In_2419,In_1883);
xnor U1324 (N_1324,In_9,In_2272);
nor U1325 (N_1325,In_1851,In_1050);
and U1326 (N_1326,In_1433,In_1338);
or U1327 (N_1327,In_1999,In_1178);
xor U1328 (N_1328,In_1742,In_1567);
nand U1329 (N_1329,In_1836,In_1899);
nand U1330 (N_1330,In_1138,In_1669);
and U1331 (N_1331,In_55,In_2051);
nand U1332 (N_1332,In_811,In_1241);
nor U1333 (N_1333,In_1033,In_1934);
or U1334 (N_1334,In_1073,In_250);
nand U1335 (N_1335,In_1011,In_835);
xor U1336 (N_1336,In_1332,In_1231);
or U1337 (N_1337,In_139,In_2311);
and U1338 (N_1338,In_1075,In_1247);
xor U1339 (N_1339,In_1346,In_2393);
nor U1340 (N_1340,In_1639,In_1031);
or U1341 (N_1341,In_2013,In_1399);
or U1342 (N_1342,In_2152,In_1715);
and U1343 (N_1343,In_1703,In_693);
or U1344 (N_1344,In_1161,In_933);
and U1345 (N_1345,In_1977,In_1974);
and U1346 (N_1346,In_2181,In_1612);
nor U1347 (N_1347,In_1560,In_87);
or U1348 (N_1348,In_1601,In_602);
or U1349 (N_1349,In_1475,In_1127);
xor U1350 (N_1350,In_1385,In_2274);
or U1351 (N_1351,In_2299,In_1521);
or U1352 (N_1352,In_1,In_812);
xnor U1353 (N_1353,In_225,In_900);
nor U1354 (N_1354,In_1445,In_59);
nand U1355 (N_1355,In_2258,In_2438);
and U1356 (N_1356,In_1080,In_804);
and U1357 (N_1357,In_2312,In_412);
and U1358 (N_1358,In_889,In_1060);
and U1359 (N_1359,In_2205,In_1303);
nor U1360 (N_1360,In_2104,In_1870);
xnor U1361 (N_1361,In_2490,In_1937);
nand U1362 (N_1362,In_1641,In_2127);
and U1363 (N_1363,In_1337,In_1335);
or U1364 (N_1364,In_1265,In_61);
or U1365 (N_1365,In_2308,In_767);
nand U1366 (N_1366,In_1177,In_148);
or U1367 (N_1367,In_195,In_674);
and U1368 (N_1368,In_844,In_1291);
nand U1369 (N_1369,In_368,In_229);
nor U1370 (N_1370,In_1515,In_509);
xor U1371 (N_1371,In_2382,In_37);
or U1372 (N_1372,In_2233,In_2468);
nand U1373 (N_1373,In_1541,In_1666);
and U1374 (N_1374,In_1185,In_2135);
xnor U1375 (N_1375,In_1970,In_1123);
xnor U1376 (N_1376,In_734,In_1861);
xor U1377 (N_1377,In_1479,In_1831);
or U1378 (N_1378,In_533,In_1275);
nor U1379 (N_1379,In_571,In_465);
or U1380 (N_1380,In_1372,In_2439);
nand U1381 (N_1381,In_1052,In_1035);
nor U1382 (N_1382,In_1247,In_712);
xnor U1383 (N_1383,In_2443,In_755);
and U1384 (N_1384,In_559,In_1177);
xnor U1385 (N_1385,In_974,In_1546);
and U1386 (N_1386,In_1460,In_1526);
and U1387 (N_1387,In_1775,In_1817);
nor U1388 (N_1388,In_1533,In_126);
nor U1389 (N_1389,In_550,In_336);
nor U1390 (N_1390,In_1715,In_1520);
nor U1391 (N_1391,In_2191,In_2142);
or U1392 (N_1392,In_2187,In_2371);
nand U1393 (N_1393,In_1100,In_2029);
nor U1394 (N_1394,In_500,In_1037);
nor U1395 (N_1395,In_1911,In_2361);
nand U1396 (N_1396,In_2073,In_812);
nand U1397 (N_1397,In_260,In_1846);
nor U1398 (N_1398,In_184,In_764);
and U1399 (N_1399,In_1326,In_1568);
nor U1400 (N_1400,In_1839,In_789);
or U1401 (N_1401,In_21,In_426);
or U1402 (N_1402,In_1918,In_2011);
xnor U1403 (N_1403,In_363,In_322);
and U1404 (N_1404,In_503,In_1189);
nand U1405 (N_1405,In_1201,In_1480);
or U1406 (N_1406,In_1818,In_1076);
nand U1407 (N_1407,In_199,In_265);
nor U1408 (N_1408,In_365,In_1930);
or U1409 (N_1409,In_193,In_2119);
or U1410 (N_1410,In_1034,In_1930);
xnor U1411 (N_1411,In_1041,In_854);
or U1412 (N_1412,In_2335,In_2396);
nor U1413 (N_1413,In_1911,In_191);
xnor U1414 (N_1414,In_875,In_224);
or U1415 (N_1415,In_1627,In_1029);
and U1416 (N_1416,In_1233,In_1777);
nand U1417 (N_1417,In_568,In_2128);
nand U1418 (N_1418,In_300,In_1748);
xor U1419 (N_1419,In_242,In_1267);
or U1420 (N_1420,In_1416,In_1632);
nand U1421 (N_1421,In_808,In_83);
nor U1422 (N_1422,In_555,In_2475);
and U1423 (N_1423,In_414,In_515);
and U1424 (N_1424,In_1297,In_1702);
or U1425 (N_1425,In_871,In_818);
or U1426 (N_1426,In_777,In_1090);
nand U1427 (N_1427,In_315,In_624);
or U1428 (N_1428,In_1735,In_162);
and U1429 (N_1429,In_61,In_1227);
nor U1430 (N_1430,In_1437,In_50);
or U1431 (N_1431,In_1850,In_968);
and U1432 (N_1432,In_2052,In_1517);
nor U1433 (N_1433,In_1194,In_2315);
or U1434 (N_1434,In_2062,In_65);
or U1435 (N_1435,In_1872,In_1923);
nor U1436 (N_1436,In_1467,In_548);
and U1437 (N_1437,In_608,In_1408);
nand U1438 (N_1438,In_1065,In_1711);
nand U1439 (N_1439,In_1000,In_857);
or U1440 (N_1440,In_332,In_843);
and U1441 (N_1441,In_2412,In_1265);
or U1442 (N_1442,In_301,In_678);
nor U1443 (N_1443,In_984,In_877);
nor U1444 (N_1444,In_963,In_1819);
and U1445 (N_1445,In_633,In_1065);
nand U1446 (N_1446,In_1754,In_1034);
nand U1447 (N_1447,In_702,In_1834);
nand U1448 (N_1448,In_647,In_1975);
nor U1449 (N_1449,In_2280,In_393);
and U1450 (N_1450,In_928,In_227);
nor U1451 (N_1451,In_324,In_1551);
nor U1452 (N_1452,In_913,In_2280);
and U1453 (N_1453,In_761,In_4);
nor U1454 (N_1454,In_1020,In_1815);
nand U1455 (N_1455,In_910,In_826);
or U1456 (N_1456,In_432,In_309);
nand U1457 (N_1457,In_905,In_1929);
nand U1458 (N_1458,In_173,In_1597);
nor U1459 (N_1459,In_366,In_923);
nand U1460 (N_1460,In_674,In_1627);
nand U1461 (N_1461,In_189,In_1004);
nand U1462 (N_1462,In_1955,In_461);
nor U1463 (N_1463,In_1561,In_1224);
nor U1464 (N_1464,In_739,In_200);
nor U1465 (N_1465,In_1181,In_1738);
nand U1466 (N_1466,In_637,In_2125);
nand U1467 (N_1467,In_1153,In_1506);
or U1468 (N_1468,In_1771,In_1847);
or U1469 (N_1469,In_1743,In_1448);
xnor U1470 (N_1470,In_1711,In_1796);
or U1471 (N_1471,In_1677,In_284);
nand U1472 (N_1472,In_320,In_1645);
and U1473 (N_1473,In_1607,In_2164);
nand U1474 (N_1474,In_2075,In_1447);
or U1475 (N_1475,In_2115,In_1769);
or U1476 (N_1476,In_325,In_1154);
nor U1477 (N_1477,In_1849,In_1025);
and U1478 (N_1478,In_196,In_2098);
and U1479 (N_1479,In_2078,In_43);
nor U1480 (N_1480,In_889,In_679);
nand U1481 (N_1481,In_1137,In_170);
xor U1482 (N_1482,In_7,In_559);
or U1483 (N_1483,In_2133,In_119);
nand U1484 (N_1484,In_2350,In_2486);
or U1485 (N_1485,In_797,In_2427);
xor U1486 (N_1486,In_1272,In_2462);
and U1487 (N_1487,In_430,In_1920);
nor U1488 (N_1488,In_1452,In_2050);
nor U1489 (N_1489,In_44,In_367);
xnor U1490 (N_1490,In_2260,In_474);
nor U1491 (N_1491,In_721,In_1679);
nor U1492 (N_1492,In_2056,In_548);
nor U1493 (N_1493,In_2379,In_1473);
nand U1494 (N_1494,In_1746,In_2301);
or U1495 (N_1495,In_1398,In_2080);
nor U1496 (N_1496,In_1397,In_1684);
xor U1497 (N_1497,In_1466,In_1022);
nor U1498 (N_1498,In_978,In_905);
xnor U1499 (N_1499,In_358,In_1275);
and U1500 (N_1500,In_2404,In_2421);
or U1501 (N_1501,In_2169,In_1904);
and U1502 (N_1502,In_287,In_1127);
nor U1503 (N_1503,In_2071,In_286);
and U1504 (N_1504,In_95,In_1228);
nor U1505 (N_1505,In_1057,In_2131);
or U1506 (N_1506,In_712,In_2449);
nand U1507 (N_1507,In_1884,In_1006);
or U1508 (N_1508,In_1685,In_690);
nand U1509 (N_1509,In_1912,In_1732);
nor U1510 (N_1510,In_902,In_2381);
nor U1511 (N_1511,In_2491,In_473);
nand U1512 (N_1512,In_2362,In_1748);
nor U1513 (N_1513,In_1295,In_82);
nand U1514 (N_1514,In_522,In_2286);
nor U1515 (N_1515,In_1682,In_1495);
nand U1516 (N_1516,In_104,In_774);
or U1517 (N_1517,In_1656,In_1077);
nand U1518 (N_1518,In_192,In_645);
or U1519 (N_1519,In_2409,In_1829);
xnor U1520 (N_1520,In_1509,In_671);
or U1521 (N_1521,In_63,In_1708);
and U1522 (N_1522,In_1332,In_218);
nand U1523 (N_1523,In_678,In_1853);
or U1524 (N_1524,In_2413,In_1372);
nor U1525 (N_1525,In_1763,In_291);
xor U1526 (N_1526,In_463,In_190);
nor U1527 (N_1527,In_2157,In_1214);
or U1528 (N_1528,In_293,In_280);
and U1529 (N_1529,In_1185,In_569);
nor U1530 (N_1530,In_1502,In_318);
or U1531 (N_1531,In_1796,In_378);
nand U1532 (N_1532,In_1990,In_1217);
or U1533 (N_1533,In_1619,In_1188);
nand U1534 (N_1534,In_1629,In_1280);
and U1535 (N_1535,In_205,In_1790);
and U1536 (N_1536,In_1936,In_677);
xor U1537 (N_1537,In_2372,In_2309);
xnor U1538 (N_1538,In_1791,In_1529);
or U1539 (N_1539,In_1347,In_1825);
and U1540 (N_1540,In_1745,In_89);
nand U1541 (N_1541,In_1148,In_244);
nand U1542 (N_1542,In_84,In_1807);
and U1543 (N_1543,In_960,In_358);
nor U1544 (N_1544,In_1563,In_1435);
or U1545 (N_1545,In_733,In_735);
and U1546 (N_1546,In_2018,In_828);
xnor U1547 (N_1547,In_2436,In_1139);
nor U1548 (N_1548,In_1751,In_2425);
or U1549 (N_1549,In_1829,In_2399);
and U1550 (N_1550,In_940,In_1562);
nor U1551 (N_1551,In_173,In_787);
nand U1552 (N_1552,In_1216,In_528);
nor U1553 (N_1553,In_1003,In_424);
nand U1554 (N_1554,In_1272,In_2061);
nand U1555 (N_1555,In_2270,In_1092);
nand U1556 (N_1556,In_1676,In_1570);
and U1557 (N_1557,In_2407,In_2314);
nand U1558 (N_1558,In_2247,In_1184);
and U1559 (N_1559,In_1014,In_931);
and U1560 (N_1560,In_430,In_2083);
xnor U1561 (N_1561,In_38,In_732);
xnor U1562 (N_1562,In_661,In_1891);
and U1563 (N_1563,In_254,In_1815);
nand U1564 (N_1564,In_1826,In_2256);
nor U1565 (N_1565,In_1519,In_2118);
nor U1566 (N_1566,In_801,In_2248);
nand U1567 (N_1567,In_1195,In_106);
or U1568 (N_1568,In_1614,In_513);
nand U1569 (N_1569,In_219,In_1457);
or U1570 (N_1570,In_980,In_1430);
nand U1571 (N_1571,In_2293,In_1175);
nand U1572 (N_1572,In_514,In_1243);
xor U1573 (N_1573,In_373,In_1113);
nand U1574 (N_1574,In_1884,In_1389);
or U1575 (N_1575,In_2319,In_969);
nor U1576 (N_1576,In_2172,In_1000);
nor U1577 (N_1577,In_2339,In_102);
xnor U1578 (N_1578,In_492,In_1945);
and U1579 (N_1579,In_1549,In_1923);
xor U1580 (N_1580,In_1822,In_76);
and U1581 (N_1581,In_1566,In_784);
nor U1582 (N_1582,In_1888,In_1392);
or U1583 (N_1583,In_956,In_2022);
and U1584 (N_1584,In_2318,In_743);
nand U1585 (N_1585,In_2495,In_2147);
nand U1586 (N_1586,In_1203,In_1251);
nor U1587 (N_1587,In_952,In_2373);
nand U1588 (N_1588,In_692,In_537);
or U1589 (N_1589,In_2001,In_1919);
nand U1590 (N_1590,In_2444,In_2383);
or U1591 (N_1591,In_951,In_1523);
nor U1592 (N_1592,In_2336,In_1260);
nand U1593 (N_1593,In_989,In_1373);
nor U1594 (N_1594,In_120,In_138);
or U1595 (N_1595,In_2355,In_308);
nand U1596 (N_1596,In_1326,In_1834);
nand U1597 (N_1597,In_2040,In_622);
nand U1598 (N_1598,In_48,In_299);
nand U1599 (N_1599,In_1748,In_1229);
or U1600 (N_1600,In_142,In_1316);
xor U1601 (N_1601,In_532,In_1368);
xor U1602 (N_1602,In_416,In_103);
xnor U1603 (N_1603,In_1812,In_209);
nor U1604 (N_1604,In_1200,In_539);
and U1605 (N_1605,In_2132,In_1164);
nand U1606 (N_1606,In_662,In_1114);
and U1607 (N_1607,In_331,In_2266);
nand U1608 (N_1608,In_751,In_754);
or U1609 (N_1609,In_2252,In_252);
and U1610 (N_1610,In_1081,In_369);
and U1611 (N_1611,In_276,In_1639);
nor U1612 (N_1612,In_1870,In_2200);
nand U1613 (N_1613,In_846,In_2283);
nor U1614 (N_1614,In_1580,In_128);
or U1615 (N_1615,In_478,In_312);
and U1616 (N_1616,In_2181,In_1626);
or U1617 (N_1617,In_1796,In_1910);
nor U1618 (N_1618,In_46,In_266);
and U1619 (N_1619,In_1466,In_1575);
nor U1620 (N_1620,In_201,In_290);
nor U1621 (N_1621,In_934,In_1151);
nor U1622 (N_1622,In_1037,In_1061);
and U1623 (N_1623,In_532,In_636);
nand U1624 (N_1624,In_1310,In_2087);
or U1625 (N_1625,In_1647,In_1037);
and U1626 (N_1626,In_637,In_1466);
xnor U1627 (N_1627,In_1724,In_1992);
nand U1628 (N_1628,In_1653,In_1174);
and U1629 (N_1629,In_661,In_2191);
or U1630 (N_1630,In_2069,In_549);
or U1631 (N_1631,In_1716,In_2191);
nand U1632 (N_1632,In_409,In_1138);
nor U1633 (N_1633,In_969,In_662);
and U1634 (N_1634,In_196,In_2018);
nand U1635 (N_1635,In_258,In_892);
nor U1636 (N_1636,In_681,In_369);
nor U1637 (N_1637,In_1914,In_2236);
or U1638 (N_1638,In_1692,In_1350);
and U1639 (N_1639,In_940,In_2003);
nor U1640 (N_1640,In_2057,In_2453);
or U1641 (N_1641,In_524,In_890);
xor U1642 (N_1642,In_1201,In_1945);
xor U1643 (N_1643,In_1872,In_1846);
xor U1644 (N_1644,In_1152,In_1325);
and U1645 (N_1645,In_1598,In_483);
nor U1646 (N_1646,In_443,In_663);
nand U1647 (N_1647,In_1147,In_1122);
or U1648 (N_1648,In_374,In_324);
nor U1649 (N_1649,In_2016,In_1264);
nor U1650 (N_1650,In_1063,In_974);
nand U1651 (N_1651,In_128,In_2329);
nor U1652 (N_1652,In_660,In_422);
and U1653 (N_1653,In_1545,In_1632);
nor U1654 (N_1654,In_1245,In_353);
nand U1655 (N_1655,In_242,In_2209);
and U1656 (N_1656,In_1751,In_784);
and U1657 (N_1657,In_1939,In_1472);
nor U1658 (N_1658,In_422,In_2178);
and U1659 (N_1659,In_1511,In_352);
or U1660 (N_1660,In_1910,In_1886);
or U1661 (N_1661,In_767,In_1942);
or U1662 (N_1662,In_2223,In_1722);
or U1663 (N_1663,In_1328,In_1745);
xnor U1664 (N_1664,In_1440,In_32);
or U1665 (N_1665,In_2310,In_218);
nor U1666 (N_1666,In_323,In_1879);
and U1667 (N_1667,In_2161,In_1017);
and U1668 (N_1668,In_334,In_530);
or U1669 (N_1669,In_2288,In_2070);
nor U1670 (N_1670,In_65,In_1907);
or U1671 (N_1671,In_1435,In_2360);
and U1672 (N_1672,In_160,In_1913);
nand U1673 (N_1673,In_981,In_1795);
nand U1674 (N_1674,In_383,In_2289);
or U1675 (N_1675,In_1237,In_675);
nand U1676 (N_1676,In_2434,In_2447);
and U1677 (N_1677,In_408,In_1870);
nand U1678 (N_1678,In_144,In_1374);
nand U1679 (N_1679,In_245,In_845);
nor U1680 (N_1680,In_2134,In_180);
nor U1681 (N_1681,In_1942,In_2374);
and U1682 (N_1682,In_1190,In_1143);
and U1683 (N_1683,In_78,In_2025);
xnor U1684 (N_1684,In_2180,In_1277);
nor U1685 (N_1685,In_2012,In_16);
or U1686 (N_1686,In_576,In_1871);
nor U1687 (N_1687,In_1570,In_1297);
xor U1688 (N_1688,In_1049,In_1422);
or U1689 (N_1689,In_131,In_2452);
and U1690 (N_1690,In_513,In_1260);
or U1691 (N_1691,In_307,In_2406);
or U1692 (N_1692,In_801,In_1285);
and U1693 (N_1693,In_1926,In_1328);
and U1694 (N_1694,In_510,In_1717);
and U1695 (N_1695,In_44,In_1364);
or U1696 (N_1696,In_448,In_2251);
nor U1697 (N_1697,In_2193,In_2496);
and U1698 (N_1698,In_244,In_228);
or U1699 (N_1699,In_669,In_392);
nand U1700 (N_1700,In_811,In_104);
or U1701 (N_1701,In_1381,In_462);
xnor U1702 (N_1702,In_1034,In_465);
xnor U1703 (N_1703,In_1217,In_49);
nor U1704 (N_1704,In_1768,In_348);
nand U1705 (N_1705,In_1431,In_682);
nand U1706 (N_1706,In_519,In_1375);
and U1707 (N_1707,In_1960,In_1987);
or U1708 (N_1708,In_529,In_1388);
nand U1709 (N_1709,In_14,In_1710);
nand U1710 (N_1710,In_1583,In_514);
or U1711 (N_1711,In_2154,In_1244);
nor U1712 (N_1712,In_236,In_2469);
nand U1713 (N_1713,In_48,In_1331);
nor U1714 (N_1714,In_917,In_453);
xnor U1715 (N_1715,In_1281,In_2351);
nand U1716 (N_1716,In_18,In_2410);
and U1717 (N_1717,In_1856,In_905);
and U1718 (N_1718,In_2224,In_1987);
nand U1719 (N_1719,In_2105,In_1856);
nor U1720 (N_1720,In_750,In_2150);
or U1721 (N_1721,In_1197,In_1234);
or U1722 (N_1722,In_32,In_2495);
or U1723 (N_1723,In_244,In_1008);
and U1724 (N_1724,In_579,In_1371);
nand U1725 (N_1725,In_893,In_883);
nand U1726 (N_1726,In_2461,In_198);
nand U1727 (N_1727,In_256,In_538);
or U1728 (N_1728,In_460,In_2419);
nand U1729 (N_1729,In_229,In_332);
and U1730 (N_1730,In_2060,In_134);
nand U1731 (N_1731,In_2242,In_2193);
or U1732 (N_1732,In_1177,In_1285);
nand U1733 (N_1733,In_304,In_1148);
nor U1734 (N_1734,In_2440,In_1021);
nor U1735 (N_1735,In_498,In_2082);
nor U1736 (N_1736,In_2318,In_519);
nor U1737 (N_1737,In_2087,In_61);
or U1738 (N_1738,In_1813,In_1173);
or U1739 (N_1739,In_2001,In_912);
nand U1740 (N_1740,In_760,In_400);
or U1741 (N_1741,In_893,In_2427);
and U1742 (N_1742,In_2271,In_489);
nor U1743 (N_1743,In_1767,In_1256);
nand U1744 (N_1744,In_1850,In_1528);
or U1745 (N_1745,In_2364,In_572);
nand U1746 (N_1746,In_1224,In_617);
and U1747 (N_1747,In_1534,In_1960);
or U1748 (N_1748,In_279,In_660);
xnor U1749 (N_1749,In_1221,In_25);
or U1750 (N_1750,In_1229,In_322);
nand U1751 (N_1751,In_1336,In_1018);
or U1752 (N_1752,In_93,In_1860);
and U1753 (N_1753,In_1481,In_2292);
and U1754 (N_1754,In_834,In_1573);
and U1755 (N_1755,In_2443,In_2178);
and U1756 (N_1756,In_958,In_2302);
nand U1757 (N_1757,In_146,In_1222);
or U1758 (N_1758,In_285,In_841);
xor U1759 (N_1759,In_706,In_1927);
and U1760 (N_1760,In_551,In_882);
nand U1761 (N_1761,In_1973,In_825);
nand U1762 (N_1762,In_746,In_1974);
nor U1763 (N_1763,In_1608,In_1922);
nor U1764 (N_1764,In_1318,In_1312);
and U1765 (N_1765,In_826,In_288);
xnor U1766 (N_1766,In_1164,In_623);
or U1767 (N_1767,In_2246,In_2317);
and U1768 (N_1768,In_276,In_1056);
nor U1769 (N_1769,In_2022,In_464);
and U1770 (N_1770,In_36,In_1013);
and U1771 (N_1771,In_1804,In_297);
nand U1772 (N_1772,In_640,In_439);
nand U1773 (N_1773,In_2284,In_500);
nand U1774 (N_1774,In_870,In_1960);
xor U1775 (N_1775,In_1362,In_893);
nor U1776 (N_1776,In_269,In_1607);
nor U1777 (N_1777,In_1697,In_1432);
and U1778 (N_1778,In_503,In_2328);
nor U1779 (N_1779,In_1086,In_144);
or U1780 (N_1780,In_2037,In_1709);
and U1781 (N_1781,In_1986,In_2018);
or U1782 (N_1782,In_499,In_2236);
and U1783 (N_1783,In_1154,In_2381);
or U1784 (N_1784,In_159,In_1168);
and U1785 (N_1785,In_754,In_1368);
nand U1786 (N_1786,In_1919,In_225);
nand U1787 (N_1787,In_1861,In_1943);
nand U1788 (N_1788,In_819,In_183);
and U1789 (N_1789,In_207,In_1926);
and U1790 (N_1790,In_2176,In_710);
nor U1791 (N_1791,In_1999,In_2374);
nor U1792 (N_1792,In_374,In_1682);
and U1793 (N_1793,In_157,In_603);
or U1794 (N_1794,In_1805,In_1637);
xnor U1795 (N_1795,In_2020,In_653);
or U1796 (N_1796,In_1129,In_1128);
and U1797 (N_1797,In_1965,In_1275);
or U1798 (N_1798,In_1457,In_1648);
or U1799 (N_1799,In_715,In_1219);
and U1800 (N_1800,In_1260,In_425);
nor U1801 (N_1801,In_136,In_1958);
nand U1802 (N_1802,In_1755,In_2293);
or U1803 (N_1803,In_1887,In_742);
nand U1804 (N_1804,In_1568,In_886);
xor U1805 (N_1805,In_1788,In_1452);
nand U1806 (N_1806,In_1748,In_1823);
nor U1807 (N_1807,In_1902,In_1836);
xor U1808 (N_1808,In_1296,In_529);
or U1809 (N_1809,In_1502,In_1004);
nand U1810 (N_1810,In_296,In_1065);
nor U1811 (N_1811,In_1017,In_2251);
nand U1812 (N_1812,In_2466,In_1524);
and U1813 (N_1813,In_1213,In_604);
nand U1814 (N_1814,In_486,In_1194);
or U1815 (N_1815,In_744,In_851);
nor U1816 (N_1816,In_2283,In_2409);
nor U1817 (N_1817,In_2317,In_1585);
xor U1818 (N_1818,In_1013,In_495);
nand U1819 (N_1819,In_196,In_308);
nor U1820 (N_1820,In_784,In_1662);
nor U1821 (N_1821,In_814,In_2203);
nand U1822 (N_1822,In_1813,In_907);
and U1823 (N_1823,In_2444,In_1795);
and U1824 (N_1824,In_1349,In_2300);
nand U1825 (N_1825,In_529,In_927);
or U1826 (N_1826,In_2219,In_1038);
and U1827 (N_1827,In_688,In_1425);
and U1828 (N_1828,In_2217,In_961);
nor U1829 (N_1829,In_1328,In_2491);
or U1830 (N_1830,In_1150,In_2311);
or U1831 (N_1831,In_510,In_67);
nor U1832 (N_1832,In_1399,In_2225);
nor U1833 (N_1833,In_1426,In_354);
or U1834 (N_1834,In_1996,In_202);
nor U1835 (N_1835,In_2239,In_2141);
nor U1836 (N_1836,In_1209,In_1766);
or U1837 (N_1837,In_2402,In_168);
xnor U1838 (N_1838,In_1599,In_1977);
xor U1839 (N_1839,In_296,In_1979);
and U1840 (N_1840,In_930,In_525);
nor U1841 (N_1841,In_1135,In_161);
nor U1842 (N_1842,In_1545,In_2050);
nor U1843 (N_1843,In_303,In_1794);
nand U1844 (N_1844,In_925,In_293);
nand U1845 (N_1845,In_300,In_2191);
xor U1846 (N_1846,In_621,In_399);
or U1847 (N_1847,In_1339,In_284);
or U1848 (N_1848,In_937,In_1901);
or U1849 (N_1849,In_1971,In_1370);
nand U1850 (N_1850,In_1684,In_2095);
nand U1851 (N_1851,In_1460,In_729);
or U1852 (N_1852,In_1801,In_55);
or U1853 (N_1853,In_1582,In_1443);
nand U1854 (N_1854,In_1518,In_2070);
nand U1855 (N_1855,In_1112,In_1546);
and U1856 (N_1856,In_931,In_2449);
and U1857 (N_1857,In_647,In_2130);
and U1858 (N_1858,In_2065,In_2326);
and U1859 (N_1859,In_580,In_924);
nor U1860 (N_1860,In_2344,In_2295);
nor U1861 (N_1861,In_1130,In_712);
nand U1862 (N_1862,In_1977,In_2264);
nor U1863 (N_1863,In_1906,In_970);
nor U1864 (N_1864,In_2316,In_1986);
and U1865 (N_1865,In_365,In_1440);
or U1866 (N_1866,In_145,In_50);
nor U1867 (N_1867,In_1455,In_170);
nor U1868 (N_1868,In_1711,In_1987);
or U1869 (N_1869,In_276,In_2104);
xor U1870 (N_1870,In_1126,In_694);
or U1871 (N_1871,In_475,In_154);
nand U1872 (N_1872,In_1267,In_1068);
and U1873 (N_1873,In_651,In_31);
nor U1874 (N_1874,In_447,In_2356);
nand U1875 (N_1875,In_947,In_1644);
nand U1876 (N_1876,In_226,In_6);
and U1877 (N_1877,In_1917,In_1185);
nor U1878 (N_1878,In_22,In_952);
and U1879 (N_1879,In_582,In_437);
or U1880 (N_1880,In_527,In_474);
xnor U1881 (N_1881,In_1378,In_470);
nor U1882 (N_1882,In_1413,In_2469);
nand U1883 (N_1883,In_2288,In_2343);
and U1884 (N_1884,In_706,In_1671);
and U1885 (N_1885,In_666,In_278);
and U1886 (N_1886,In_1593,In_97);
or U1887 (N_1887,In_2370,In_318);
nor U1888 (N_1888,In_1936,In_2433);
nand U1889 (N_1889,In_324,In_550);
nand U1890 (N_1890,In_135,In_1394);
and U1891 (N_1891,In_655,In_237);
or U1892 (N_1892,In_1624,In_808);
xor U1893 (N_1893,In_374,In_471);
nor U1894 (N_1894,In_2436,In_137);
nor U1895 (N_1895,In_1025,In_1825);
or U1896 (N_1896,In_449,In_571);
or U1897 (N_1897,In_1862,In_2390);
nor U1898 (N_1898,In_235,In_2473);
or U1899 (N_1899,In_329,In_310);
and U1900 (N_1900,In_1246,In_1839);
or U1901 (N_1901,In_790,In_1095);
nor U1902 (N_1902,In_741,In_1667);
nand U1903 (N_1903,In_1165,In_756);
nand U1904 (N_1904,In_848,In_371);
and U1905 (N_1905,In_2233,In_279);
nor U1906 (N_1906,In_1270,In_1750);
or U1907 (N_1907,In_2032,In_830);
nand U1908 (N_1908,In_1917,In_439);
or U1909 (N_1909,In_776,In_467);
xor U1910 (N_1910,In_404,In_1124);
or U1911 (N_1911,In_2427,In_1590);
nor U1912 (N_1912,In_2455,In_2188);
and U1913 (N_1913,In_2185,In_1576);
and U1914 (N_1914,In_515,In_1799);
or U1915 (N_1915,In_1543,In_267);
nand U1916 (N_1916,In_1626,In_880);
or U1917 (N_1917,In_2312,In_52);
nor U1918 (N_1918,In_2028,In_648);
nor U1919 (N_1919,In_375,In_1870);
nand U1920 (N_1920,In_484,In_2015);
and U1921 (N_1921,In_1285,In_2472);
and U1922 (N_1922,In_129,In_115);
nor U1923 (N_1923,In_2167,In_444);
nor U1924 (N_1924,In_810,In_990);
and U1925 (N_1925,In_2409,In_1321);
xnor U1926 (N_1926,In_1587,In_2281);
or U1927 (N_1927,In_209,In_1661);
and U1928 (N_1928,In_1393,In_911);
nor U1929 (N_1929,In_1295,In_1521);
and U1930 (N_1930,In_551,In_420);
or U1931 (N_1931,In_1023,In_2336);
xor U1932 (N_1932,In_2114,In_1324);
and U1933 (N_1933,In_2195,In_1054);
nand U1934 (N_1934,In_2468,In_590);
and U1935 (N_1935,In_1974,In_140);
nor U1936 (N_1936,In_1977,In_1028);
nand U1937 (N_1937,In_1336,In_2066);
and U1938 (N_1938,In_1581,In_2380);
or U1939 (N_1939,In_1652,In_1282);
nor U1940 (N_1940,In_94,In_2430);
nor U1941 (N_1941,In_2499,In_2015);
or U1942 (N_1942,In_275,In_1249);
nor U1943 (N_1943,In_1142,In_2193);
nand U1944 (N_1944,In_1506,In_567);
nand U1945 (N_1945,In_1269,In_1017);
xor U1946 (N_1946,In_1293,In_1730);
or U1947 (N_1947,In_1259,In_1748);
or U1948 (N_1948,In_2412,In_42);
and U1949 (N_1949,In_1831,In_1274);
nand U1950 (N_1950,In_248,In_630);
nor U1951 (N_1951,In_1831,In_1236);
or U1952 (N_1952,In_778,In_1581);
nor U1953 (N_1953,In_1384,In_2389);
or U1954 (N_1954,In_2105,In_122);
or U1955 (N_1955,In_633,In_1173);
nand U1956 (N_1956,In_1954,In_1492);
nand U1957 (N_1957,In_948,In_694);
and U1958 (N_1958,In_1590,In_161);
and U1959 (N_1959,In_295,In_2225);
or U1960 (N_1960,In_1891,In_1190);
and U1961 (N_1961,In_2278,In_786);
or U1962 (N_1962,In_1625,In_1463);
nor U1963 (N_1963,In_525,In_1698);
or U1964 (N_1964,In_900,In_1118);
or U1965 (N_1965,In_1326,In_1936);
nand U1966 (N_1966,In_2486,In_966);
or U1967 (N_1967,In_1242,In_1433);
nand U1968 (N_1968,In_1561,In_487);
nor U1969 (N_1969,In_434,In_2404);
nand U1970 (N_1970,In_1107,In_1037);
xnor U1971 (N_1971,In_162,In_436);
nor U1972 (N_1972,In_2455,In_791);
and U1973 (N_1973,In_1566,In_1974);
and U1974 (N_1974,In_2030,In_553);
and U1975 (N_1975,In_773,In_1185);
nor U1976 (N_1976,In_2468,In_1412);
and U1977 (N_1977,In_1155,In_2085);
nand U1978 (N_1978,In_1748,In_1933);
xnor U1979 (N_1979,In_2040,In_98);
or U1980 (N_1980,In_1050,In_1224);
and U1981 (N_1981,In_738,In_780);
xor U1982 (N_1982,In_564,In_883);
and U1983 (N_1983,In_1351,In_339);
and U1984 (N_1984,In_2493,In_1865);
nand U1985 (N_1985,In_2163,In_1049);
and U1986 (N_1986,In_918,In_992);
or U1987 (N_1987,In_473,In_689);
xor U1988 (N_1988,In_2259,In_2425);
or U1989 (N_1989,In_2403,In_1141);
nor U1990 (N_1990,In_1779,In_849);
or U1991 (N_1991,In_1482,In_121);
or U1992 (N_1992,In_2140,In_373);
and U1993 (N_1993,In_2210,In_867);
xnor U1994 (N_1994,In_1908,In_1429);
nand U1995 (N_1995,In_1434,In_2261);
and U1996 (N_1996,In_2103,In_38);
and U1997 (N_1997,In_907,In_2325);
and U1998 (N_1998,In_4,In_1669);
xnor U1999 (N_1999,In_81,In_1365);
nor U2000 (N_2000,In_1839,In_1988);
nand U2001 (N_2001,In_252,In_232);
or U2002 (N_2002,In_847,In_544);
xor U2003 (N_2003,In_1349,In_1538);
or U2004 (N_2004,In_1429,In_138);
and U2005 (N_2005,In_1046,In_1871);
and U2006 (N_2006,In_2006,In_1101);
nor U2007 (N_2007,In_579,In_86);
or U2008 (N_2008,In_695,In_493);
nand U2009 (N_2009,In_239,In_2006);
xnor U2010 (N_2010,In_1429,In_544);
nor U2011 (N_2011,In_688,In_1900);
nand U2012 (N_2012,In_344,In_1638);
nand U2013 (N_2013,In_1528,In_1162);
and U2014 (N_2014,In_605,In_1804);
or U2015 (N_2015,In_2240,In_1715);
xnor U2016 (N_2016,In_493,In_327);
nor U2017 (N_2017,In_836,In_680);
or U2018 (N_2018,In_1431,In_277);
or U2019 (N_2019,In_2456,In_473);
nand U2020 (N_2020,In_661,In_796);
and U2021 (N_2021,In_1755,In_761);
nand U2022 (N_2022,In_736,In_845);
and U2023 (N_2023,In_950,In_1593);
or U2024 (N_2024,In_1845,In_961);
and U2025 (N_2025,In_149,In_1204);
nor U2026 (N_2026,In_429,In_2358);
nor U2027 (N_2027,In_2415,In_331);
nor U2028 (N_2028,In_2317,In_852);
or U2029 (N_2029,In_1114,In_2031);
xor U2030 (N_2030,In_1923,In_1067);
and U2031 (N_2031,In_180,In_1034);
xor U2032 (N_2032,In_1159,In_1515);
and U2033 (N_2033,In_1740,In_341);
and U2034 (N_2034,In_1568,In_415);
nor U2035 (N_2035,In_290,In_1004);
and U2036 (N_2036,In_1993,In_1410);
nor U2037 (N_2037,In_2087,In_1151);
and U2038 (N_2038,In_2025,In_816);
or U2039 (N_2039,In_423,In_1841);
or U2040 (N_2040,In_1234,In_2497);
nor U2041 (N_2041,In_783,In_166);
and U2042 (N_2042,In_2111,In_1802);
or U2043 (N_2043,In_1425,In_1723);
nor U2044 (N_2044,In_2297,In_1253);
and U2045 (N_2045,In_563,In_1233);
nor U2046 (N_2046,In_797,In_1945);
nor U2047 (N_2047,In_1088,In_269);
nor U2048 (N_2048,In_481,In_89);
nor U2049 (N_2049,In_1016,In_1554);
nor U2050 (N_2050,In_1003,In_33);
nor U2051 (N_2051,In_25,In_2346);
xor U2052 (N_2052,In_1473,In_640);
or U2053 (N_2053,In_653,In_2329);
or U2054 (N_2054,In_453,In_2433);
nor U2055 (N_2055,In_1805,In_2492);
or U2056 (N_2056,In_1464,In_1213);
nor U2057 (N_2057,In_1537,In_1895);
nand U2058 (N_2058,In_1477,In_1356);
and U2059 (N_2059,In_1476,In_2007);
nand U2060 (N_2060,In_740,In_111);
or U2061 (N_2061,In_2475,In_1194);
or U2062 (N_2062,In_144,In_273);
and U2063 (N_2063,In_1891,In_1411);
and U2064 (N_2064,In_730,In_2038);
nand U2065 (N_2065,In_262,In_1759);
nand U2066 (N_2066,In_2265,In_2426);
and U2067 (N_2067,In_2164,In_946);
or U2068 (N_2068,In_2404,In_1122);
xor U2069 (N_2069,In_425,In_2095);
and U2070 (N_2070,In_2033,In_2162);
nor U2071 (N_2071,In_1111,In_1488);
nand U2072 (N_2072,In_2110,In_2140);
nor U2073 (N_2073,In_2287,In_2311);
xnor U2074 (N_2074,In_1189,In_150);
or U2075 (N_2075,In_568,In_1661);
or U2076 (N_2076,In_536,In_1442);
xor U2077 (N_2077,In_62,In_2342);
xor U2078 (N_2078,In_606,In_230);
nand U2079 (N_2079,In_1460,In_669);
nand U2080 (N_2080,In_99,In_2338);
nor U2081 (N_2081,In_698,In_2065);
xor U2082 (N_2082,In_868,In_454);
xor U2083 (N_2083,In_1517,In_301);
or U2084 (N_2084,In_1920,In_1615);
or U2085 (N_2085,In_352,In_996);
nand U2086 (N_2086,In_1846,In_1152);
and U2087 (N_2087,In_907,In_1858);
nand U2088 (N_2088,In_2190,In_150);
nand U2089 (N_2089,In_1422,In_53);
or U2090 (N_2090,In_378,In_1857);
nor U2091 (N_2091,In_96,In_1703);
and U2092 (N_2092,In_1363,In_387);
and U2093 (N_2093,In_1894,In_1158);
or U2094 (N_2094,In_1544,In_932);
and U2095 (N_2095,In_1933,In_2186);
and U2096 (N_2096,In_25,In_946);
or U2097 (N_2097,In_53,In_858);
nand U2098 (N_2098,In_1223,In_1004);
nand U2099 (N_2099,In_2145,In_188);
and U2100 (N_2100,In_605,In_19);
xor U2101 (N_2101,In_982,In_2202);
or U2102 (N_2102,In_1404,In_27);
xnor U2103 (N_2103,In_1370,In_956);
xnor U2104 (N_2104,In_630,In_1029);
nand U2105 (N_2105,In_994,In_630);
and U2106 (N_2106,In_1301,In_1501);
and U2107 (N_2107,In_2131,In_2094);
nand U2108 (N_2108,In_2123,In_797);
nor U2109 (N_2109,In_1980,In_1727);
or U2110 (N_2110,In_2478,In_2149);
nand U2111 (N_2111,In_1551,In_762);
xnor U2112 (N_2112,In_39,In_2494);
nor U2113 (N_2113,In_1297,In_943);
nor U2114 (N_2114,In_2243,In_1391);
nor U2115 (N_2115,In_1560,In_1893);
nand U2116 (N_2116,In_2370,In_93);
and U2117 (N_2117,In_395,In_2174);
or U2118 (N_2118,In_2115,In_1094);
and U2119 (N_2119,In_1838,In_1627);
xor U2120 (N_2120,In_554,In_2165);
xor U2121 (N_2121,In_2194,In_649);
or U2122 (N_2122,In_2033,In_1277);
or U2123 (N_2123,In_1438,In_906);
nor U2124 (N_2124,In_977,In_1836);
nand U2125 (N_2125,In_1380,In_1118);
or U2126 (N_2126,In_992,In_43);
xor U2127 (N_2127,In_432,In_590);
nor U2128 (N_2128,In_2384,In_560);
xnor U2129 (N_2129,In_1835,In_258);
or U2130 (N_2130,In_174,In_809);
and U2131 (N_2131,In_1578,In_1013);
nand U2132 (N_2132,In_18,In_2486);
or U2133 (N_2133,In_1593,In_884);
xor U2134 (N_2134,In_499,In_1369);
and U2135 (N_2135,In_1043,In_1124);
nand U2136 (N_2136,In_307,In_201);
and U2137 (N_2137,In_881,In_3);
nand U2138 (N_2138,In_1114,In_732);
or U2139 (N_2139,In_1100,In_382);
nor U2140 (N_2140,In_253,In_13);
and U2141 (N_2141,In_1405,In_1410);
or U2142 (N_2142,In_1520,In_625);
xnor U2143 (N_2143,In_1643,In_161);
xnor U2144 (N_2144,In_1360,In_2063);
nand U2145 (N_2145,In_1056,In_850);
or U2146 (N_2146,In_1394,In_1432);
nor U2147 (N_2147,In_2019,In_1381);
and U2148 (N_2148,In_1547,In_2330);
and U2149 (N_2149,In_712,In_2305);
and U2150 (N_2150,In_2107,In_1791);
and U2151 (N_2151,In_476,In_2034);
and U2152 (N_2152,In_2040,In_623);
nor U2153 (N_2153,In_512,In_1268);
nor U2154 (N_2154,In_823,In_2494);
nand U2155 (N_2155,In_1685,In_1841);
nor U2156 (N_2156,In_470,In_565);
nor U2157 (N_2157,In_1672,In_728);
or U2158 (N_2158,In_2229,In_1045);
and U2159 (N_2159,In_635,In_1822);
nor U2160 (N_2160,In_1899,In_430);
or U2161 (N_2161,In_338,In_2396);
nand U2162 (N_2162,In_1502,In_779);
nor U2163 (N_2163,In_721,In_2102);
nand U2164 (N_2164,In_2393,In_1547);
nor U2165 (N_2165,In_787,In_1052);
xnor U2166 (N_2166,In_987,In_896);
nor U2167 (N_2167,In_1870,In_1924);
and U2168 (N_2168,In_1337,In_1140);
nand U2169 (N_2169,In_2465,In_170);
or U2170 (N_2170,In_2128,In_1971);
or U2171 (N_2171,In_1646,In_166);
nand U2172 (N_2172,In_1545,In_206);
nand U2173 (N_2173,In_1873,In_2192);
and U2174 (N_2174,In_1409,In_1027);
xor U2175 (N_2175,In_993,In_437);
nand U2176 (N_2176,In_912,In_101);
nor U2177 (N_2177,In_659,In_1916);
nand U2178 (N_2178,In_954,In_2316);
nor U2179 (N_2179,In_1309,In_231);
and U2180 (N_2180,In_1967,In_1106);
nor U2181 (N_2181,In_2479,In_1878);
or U2182 (N_2182,In_721,In_2491);
and U2183 (N_2183,In_61,In_1218);
or U2184 (N_2184,In_1227,In_798);
nand U2185 (N_2185,In_427,In_13);
or U2186 (N_2186,In_85,In_399);
or U2187 (N_2187,In_2291,In_879);
and U2188 (N_2188,In_42,In_289);
or U2189 (N_2189,In_2315,In_2328);
nor U2190 (N_2190,In_355,In_541);
nand U2191 (N_2191,In_2386,In_1560);
and U2192 (N_2192,In_919,In_2443);
xnor U2193 (N_2193,In_1234,In_2305);
or U2194 (N_2194,In_1075,In_2390);
nand U2195 (N_2195,In_1928,In_1625);
nand U2196 (N_2196,In_1151,In_2320);
or U2197 (N_2197,In_1911,In_1646);
or U2198 (N_2198,In_1572,In_1416);
xnor U2199 (N_2199,In_1585,In_2403);
nor U2200 (N_2200,In_2032,In_1859);
and U2201 (N_2201,In_1639,In_683);
nor U2202 (N_2202,In_70,In_1562);
nor U2203 (N_2203,In_22,In_1954);
nand U2204 (N_2204,In_355,In_1488);
or U2205 (N_2205,In_1486,In_1136);
nand U2206 (N_2206,In_687,In_1789);
or U2207 (N_2207,In_1064,In_2332);
nand U2208 (N_2208,In_1062,In_1967);
xnor U2209 (N_2209,In_1978,In_1853);
or U2210 (N_2210,In_2416,In_1018);
and U2211 (N_2211,In_1846,In_1017);
xnor U2212 (N_2212,In_2277,In_982);
nor U2213 (N_2213,In_1512,In_1032);
nor U2214 (N_2214,In_87,In_964);
and U2215 (N_2215,In_510,In_1388);
xor U2216 (N_2216,In_1324,In_1109);
nor U2217 (N_2217,In_1370,In_1933);
and U2218 (N_2218,In_299,In_1677);
and U2219 (N_2219,In_1974,In_788);
nand U2220 (N_2220,In_1277,In_1881);
xnor U2221 (N_2221,In_1572,In_2360);
or U2222 (N_2222,In_973,In_330);
and U2223 (N_2223,In_588,In_1996);
xnor U2224 (N_2224,In_1066,In_1451);
nor U2225 (N_2225,In_913,In_905);
or U2226 (N_2226,In_665,In_1204);
nand U2227 (N_2227,In_2270,In_2018);
and U2228 (N_2228,In_733,In_165);
nor U2229 (N_2229,In_1499,In_1149);
or U2230 (N_2230,In_993,In_2462);
nor U2231 (N_2231,In_1451,In_50);
nand U2232 (N_2232,In_2392,In_1299);
nor U2233 (N_2233,In_1149,In_2483);
nor U2234 (N_2234,In_492,In_887);
nand U2235 (N_2235,In_527,In_25);
xor U2236 (N_2236,In_1408,In_546);
nand U2237 (N_2237,In_541,In_2496);
xnor U2238 (N_2238,In_1584,In_2137);
nand U2239 (N_2239,In_1785,In_2490);
nor U2240 (N_2240,In_1532,In_2314);
nand U2241 (N_2241,In_1963,In_2319);
nand U2242 (N_2242,In_2216,In_2417);
or U2243 (N_2243,In_1745,In_127);
nor U2244 (N_2244,In_1879,In_2369);
xor U2245 (N_2245,In_1914,In_387);
and U2246 (N_2246,In_1098,In_742);
xnor U2247 (N_2247,In_326,In_903);
nand U2248 (N_2248,In_1363,In_999);
nor U2249 (N_2249,In_1572,In_2296);
xor U2250 (N_2250,In_1612,In_28);
xnor U2251 (N_2251,In_704,In_1614);
and U2252 (N_2252,In_199,In_1618);
xnor U2253 (N_2253,In_306,In_1681);
and U2254 (N_2254,In_2022,In_2464);
nor U2255 (N_2255,In_696,In_2057);
nand U2256 (N_2256,In_2406,In_1318);
xnor U2257 (N_2257,In_261,In_2092);
nor U2258 (N_2258,In_278,In_237);
nand U2259 (N_2259,In_793,In_1596);
and U2260 (N_2260,In_1685,In_2163);
and U2261 (N_2261,In_329,In_1799);
and U2262 (N_2262,In_1691,In_89);
or U2263 (N_2263,In_1798,In_1416);
nand U2264 (N_2264,In_2181,In_974);
nor U2265 (N_2265,In_1011,In_1272);
and U2266 (N_2266,In_2496,In_1329);
or U2267 (N_2267,In_2255,In_1520);
and U2268 (N_2268,In_2272,In_394);
nor U2269 (N_2269,In_1245,In_1372);
and U2270 (N_2270,In_128,In_2258);
nand U2271 (N_2271,In_2281,In_507);
or U2272 (N_2272,In_1882,In_2197);
and U2273 (N_2273,In_1153,In_781);
nor U2274 (N_2274,In_1080,In_2122);
nand U2275 (N_2275,In_912,In_525);
and U2276 (N_2276,In_1373,In_1285);
or U2277 (N_2277,In_1280,In_38);
or U2278 (N_2278,In_2270,In_2391);
nand U2279 (N_2279,In_2420,In_388);
nand U2280 (N_2280,In_473,In_865);
or U2281 (N_2281,In_9,In_905);
nor U2282 (N_2282,In_1974,In_1691);
and U2283 (N_2283,In_63,In_1490);
or U2284 (N_2284,In_255,In_1925);
nand U2285 (N_2285,In_1293,In_1572);
nand U2286 (N_2286,In_1465,In_2115);
nor U2287 (N_2287,In_1865,In_290);
xor U2288 (N_2288,In_1107,In_1954);
nand U2289 (N_2289,In_958,In_163);
and U2290 (N_2290,In_863,In_468);
and U2291 (N_2291,In_375,In_746);
nor U2292 (N_2292,In_2237,In_2408);
or U2293 (N_2293,In_906,In_990);
nor U2294 (N_2294,In_266,In_556);
nand U2295 (N_2295,In_162,In_1191);
nand U2296 (N_2296,In_1442,In_442);
xor U2297 (N_2297,In_2007,In_517);
nor U2298 (N_2298,In_132,In_437);
and U2299 (N_2299,In_839,In_1379);
nor U2300 (N_2300,In_2056,In_1869);
and U2301 (N_2301,In_981,In_954);
or U2302 (N_2302,In_981,In_220);
and U2303 (N_2303,In_2243,In_1639);
nand U2304 (N_2304,In_2423,In_1999);
nand U2305 (N_2305,In_1126,In_1281);
xor U2306 (N_2306,In_775,In_1138);
or U2307 (N_2307,In_2483,In_1739);
or U2308 (N_2308,In_367,In_2409);
or U2309 (N_2309,In_2242,In_480);
nor U2310 (N_2310,In_1083,In_1126);
or U2311 (N_2311,In_2373,In_101);
and U2312 (N_2312,In_934,In_651);
nand U2313 (N_2313,In_2230,In_1784);
and U2314 (N_2314,In_1046,In_2318);
nand U2315 (N_2315,In_2107,In_329);
nor U2316 (N_2316,In_1393,In_1286);
and U2317 (N_2317,In_2294,In_1200);
xor U2318 (N_2318,In_1185,In_1556);
or U2319 (N_2319,In_684,In_1316);
nand U2320 (N_2320,In_310,In_255);
and U2321 (N_2321,In_1254,In_2260);
nand U2322 (N_2322,In_2134,In_2152);
nand U2323 (N_2323,In_50,In_525);
nand U2324 (N_2324,In_952,In_2424);
nand U2325 (N_2325,In_255,In_28);
nand U2326 (N_2326,In_2417,In_1711);
xnor U2327 (N_2327,In_709,In_1762);
xnor U2328 (N_2328,In_1849,In_679);
and U2329 (N_2329,In_1335,In_2093);
xor U2330 (N_2330,In_2076,In_1934);
xnor U2331 (N_2331,In_2011,In_2112);
nand U2332 (N_2332,In_411,In_2498);
and U2333 (N_2333,In_1752,In_1406);
or U2334 (N_2334,In_285,In_224);
nor U2335 (N_2335,In_652,In_1427);
and U2336 (N_2336,In_887,In_1283);
nor U2337 (N_2337,In_1311,In_1945);
and U2338 (N_2338,In_2403,In_485);
and U2339 (N_2339,In_2412,In_2055);
nand U2340 (N_2340,In_157,In_1616);
nand U2341 (N_2341,In_1403,In_1731);
and U2342 (N_2342,In_1672,In_1807);
and U2343 (N_2343,In_1200,In_612);
or U2344 (N_2344,In_294,In_1819);
nor U2345 (N_2345,In_144,In_1769);
and U2346 (N_2346,In_723,In_1621);
or U2347 (N_2347,In_1495,In_2464);
nor U2348 (N_2348,In_1185,In_678);
xor U2349 (N_2349,In_1653,In_2178);
or U2350 (N_2350,In_2148,In_778);
or U2351 (N_2351,In_1849,In_620);
or U2352 (N_2352,In_269,In_2183);
nand U2353 (N_2353,In_565,In_2235);
or U2354 (N_2354,In_990,In_1045);
nand U2355 (N_2355,In_2287,In_1428);
and U2356 (N_2356,In_138,In_2060);
and U2357 (N_2357,In_1442,In_2262);
nand U2358 (N_2358,In_340,In_712);
nor U2359 (N_2359,In_2313,In_1434);
nand U2360 (N_2360,In_297,In_491);
or U2361 (N_2361,In_781,In_554);
and U2362 (N_2362,In_1106,In_2207);
and U2363 (N_2363,In_811,In_1527);
nor U2364 (N_2364,In_1084,In_251);
nor U2365 (N_2365,In_541,In_2233);
or U2366 (N_2366,In_2341,In_1107);
and U2367 (N_2367,In_361,In_1374);
and U2368 (N_2368,In_1865,In_1720);
and U2369 (N_2369,In_3,In_2213);
xor U2370 (N_2370,In_1293,In_298);
xor U2371 (N_2371,In_244,In_2282);
nor U2372 (N_2372,In_2312,In_169);
nand U2373 (N_2373,In_2074,In_140);
and U2374 (N_2374,In_1908,In_81);
nor U2375 (N_2375,In_504,In_2022);
nand U2376 (N_2376,In_202,In_1376);
nand U2377 (N_2377,In_553,In_230);
or U2378 (N_2378,In_1875,In_1827);
nand U2379 (N_2379,In_1170,In_1357);
nor U2380 (N_2380,In_2326,In_1291);
nand U2381 (N_2381,In_1830,In_2341);
or U2382 (N_2382,In_1804,In_365);
xnor U2383 (N_2383,In_772,In_827);
and U2384 (N_2384,In_856,In_1926);
and U2385 (N_2385,In_1963,In_1571);
nand U2386 (N_2386,In_277,In_792);
or U2387 (N_2387,In_237,In_2087);
and U2388 (N_2388,In_0,In_688);
and U2389 (N_2389,In_1941,In_1499);
nand U2390 (N_2390,In_1063,In_720);
and U2391 (N_2391,In_447,In_1765);
or U2392 (N_2392,In_105,In_1608);
nor U2393 (N_2393,In_2347,In_174);
nor U2394 (N_2394,In_2468,In_362);
nand U2395 (N_2395,In_637,In_928);
nor U2396 (N_2396,In_733,In_2073);
nand U2397 (N_2397,In_1923,In_1291);
xnor U2398 (N_2398,In_1011,In_2298);
nand U2399 (N_2399,In_2150,In_319);
and U2400 (N_2400,In_689,In_745);
and U2401 (N_2401,In_847,In_256);
and U2402 (N_2402,In_900,In_990);
or U2403 (N_2403,In_160,In_2083);
nand U2404 (N_2404,In_2276,In_905);
xnor U2405 (N_2405,In_1754,In_1806);
nand U2406 (N_2406,In_1891,In_1016);
nor U2407 (N_2407,In_1035,In_716);
or U2408 (N_2408,In_2023,In_1770);
and U2409 (N_2409,In_1604,In_2025);
and U2410 (N_2410,In_100,In_409);
xnor U2411 (N_2411,In_272,In_946);
or U2412 (N_2412,In_462,In_81);
nand U2413 (N_2413,In_1786,In_2422);
and U2414 (N_2414,In_1608,In_543);
nand U2415 (N_2415,In_964,In_2474);
nand U2416 (N_2416,In_72,In_2022);
nand U2417 (N_2417,In_2195,In_1619);
or U2418 (N_2418,In_1087,In_70);
nand U2419 (N_2419,In_1962,In_1151);
xnor U2420 (N_2420,In_982,In_1406);
nor U2421 (N_2421,In_1611,In_1606);
nor U2422 (N_2422,In_2438,In_609);
xor U2423 (N_2423,In_999,In_270);
nand U2424 (N_2424,In_1673,In_1850);
nand U2425 (N_2425,In_31,In_176);
nor U2426 (N_2426,In_2290,In_1269);
or U2427 (N_2427,In_2184,In_312);
or U2428 (N_2428,In_19,In_1608);
nand U2429 (N_2429,In_1194,In_2266);
or U2430 (N_2430,In_213,In_1518);
or U2431 (N_2431,In_1126,In_1688);
nor U2432 (N_2432,In_1625,In_234);
nor U2433 (N_2433,In_1028,In_887);
xor U2434 (N_2434,In_1807,In_1887);
nor U2435 (N_2435,In_57,In_1406);
nor U2436 (N_2436,In_1871,In_1584);
or U2437 (N_2437,In_2404,In_1922);
and U2438 (N_2438,In_1757,In_492);
or U2439 (N_2439,In_1764,In_934);
nor U2440 (N_2440,In_1483,In_1589);
or U2441 (N_2441,In_178,In_382);
nand U2442 (N_2442,In_1522,In_391);
or U2443 (N_2443,In_1191,In_916);
and U2444 (N_2444,In_703,In_1971);
or U2445 (N_2445,In_1336,In_1986);
and U2446 (N_2446,In_721,In_638);
nand U2447 (N_2447,In_1505,In_1226);
nand U2448 (N_2448,In_889,In_892);
nand U2449 (N_2449,In_1307,In_2034);
xor U2450 (N_2450,In_291,In_1131);
nor U2451 (N_2451,In_2382,In_1191);
nand U2452 (N_2452,In_1354,In_2239);
xor U2453 (N_2453,In_1269,In_2278);
nand U2454 (N_2454,In_1073,In_2031);
nand U2455 (N_2455,In_1952,In_1794);
nand U2456 (N_2456,In_1283,In_1388);
nand U2457 (N_2457,In_252,In_697);
nand U2458 (N_2458,In_2473,In_134);
or U2459 (N_2459,In_1947,In_867);
xor U2460 (N_2460,In_1165,In_1882);
nand U2461 (N_2461,In_1330,In_994);
nor U2462 (N_2462,In_1962,In_681);
xnor U2463 (N_2463,In_2456,In_1926);
or U2464 (N_2464,In_818,In_1274);
nor U2465 (N_2465,In_1481,In_625);
nor U2466 (N_2466,In_1582,In_327);
nor U2467 (N_2467,In_2277,In_28);
or U2468 (N_2468,In_1880,In_665);
nand U2469 (N_2469,In_1072,In_533);
and U2470 (N_2470,In_1701,In_1483);
and U2471 (N_2471,In_1477,In_545);
or U2472 (N_2472,In_1941,In_2474);
nand U2473 (N_2473,In_587,In_2303);
nor U2474 (N_2474,In_188,In_446);
or U2475 (N_2475,In_1100,In_2414);
nor U2476 (N_2476,In_331,In_2126);
and U2477 (N_2477,In_1245,In_736);
nor U2478 (N_2478,In_1034,In_1595);
and U2479 (N_2479,In_2228,In_865);
nor U2480 (N_2480,In_1759,In_1211);
xnor U2481 (N_2481,In_1166,In_194);
xor U2482 (N_2482,In_284,In_2097);
or U2483 (N_2483,In_101,In_1717);
nand U2484 (N_2484,In_2120,In_1484);
nand U2485 (N_2485,In_278,In_2330);
and U2486 (N_2486,In_2184,In_1046);
nand U2487 (N_2487,In_1877,In_2371);
nand U2488 (N_2488,In_1648,In_714);
nand U2489 (N_2489,In_1006,In_211);
nand U2490 (N_2490,In_1717,In_179);
nor U2491 (N_2491,In_2487,In_2477);
nand U2492 (N_2492,In_1180,In_1403);
nor U2493 (N_2493,In_2203,In_1760);
nor U2494 (N_2494,In_429,In_1106);
and U2495 (N_2495,In_468,In_482);
and U2496 (N_2496,In_1213,In_485);
and U2497 (N_2497,In_430,In_376);
or U2498 (N_2498,In_1478,In_534);
nand U2499 (N_2499,In_2380,In_1027);
or U2500 (N_2500,N_1903,N_10);
or U2501 (N_2501,N_353,N_2240);
nand U2502 (N_2502,N_1191,N_2497);
nor U2503 (N_2503,N_796,N_1257);
or U2504 (N_2504,N_452,N_280);
nor U2505 (N_2505,N_832,N_1069);
nand U2506 (N_2506,N_1455,N_422);
nand U2507 (N_2507,N_51,N_174);
or U2508 (N_2508,N_413,N_118);
xnor U2509 (N_2509,N_626,N_2144);
nor U2510 (N_2510,N_133,N_1316);
nand U2511 (N_2511,N_1101,N_2351);
nor U2512 (N_2512,N_766,N_2025);
nor U2513 (N_2513,N_1969,N_8);
nor U2514 (N_2514,N_697,N_1471);
and U2515 (N_2515,N_1196,N_131);
nand U2516 (N_2516,N_2337,N_238);
and U2517 (N_2517,N_2410,N_1902);
nor U2518 (N_2518,N_527,N_850);
or U2519 (N_2519,N_783,N_2285);
or U2520 (N_2520,N_641,N_758);
or U2521 (N_2521,N_704,N_1401);
nor U2522 (N_2522,N_1839,N_1834);
nand U2523 (N_2523,N_244,N_838);
or U2524 (N_2524,N_763,N_1350);
nor U2525 (N_2525,N_135,N_2278);
or U2526 (N_2526,N_1231,N_2349);
and U2527 (N_2527,N_1108,N_872);
and U2528 (N_2528,N_2159,N_1097);
nand U2529 (N_2529,N_1750,N_1352);
or U2530 (N_2530,N_1692,N_310);
and U2531 (N_2531,N_540,N_2065);
and U2532 (N_2532,N_1922,N_774);
or U2533 (N_2533,N_706,N_1580);
or U2534 (N_2534,N_1657,N_568);
and U2535 (N_2535,N_543,N_726);
nor U2536 (N_2536,N_762,N_1203);
nor U2537 (N_2537,N_2475,N_1914);
xnor U2538 (N_2538,N_2369,N_1768);
and U2539 (N_2539,N_996,N_2268);
nand U2540 (N_2540,N_752,N_659);
nor U2541 (N_2541,N_582,N_1075);
xor U2542 (N_2542,N_349,N_152);
or U2543 (N_2543,N_879,N_1875);
or U2544 (N_2544,N_1267,N_567);
and U2545 (N_2545,N_2283,N_1439);
nor U2546 (N_2546,N_75,N_38);
nand U2547 (N_2547,N_846,N_1539);
nand U2548 (N_2548,N_2361,N_732);
nand U2549 (N_2549,N_2463,N_246);
and U2550 (N_2550,N_1452,N_1911);
nand U2551 (N_2551,N_1727,N_6);
or U2552 (N_2552,N_1438,N_259);
nor U2553 (N_2553,N_2284,N_1232);
and U2554 (N_2554,N_1858,N_1984);
and U2555 (N_2555,N_2163,N_1093);
nor U2556 (N_2556,N_1558,N_2400);
nand U2557 (N_2557,N_2030,N_594);
nand U2558 (N_2558,N_2033,N_27);
nor U2559 (N_2559,N_1104,N_648);
or U2560 (N_2560,N_2418,N_2239);
or U2561 (N_2561,N_2368,N_285);
or U2562 (N_2562,N_1652,N_1449);
nand U2563 (N_2563,N_702,N_1913);
nand U2564 (N_2564,N_2242,N_1724);
or U2565 (N_2565,N_1906,N_1251);
nand U2566 (N_2566,N_278,N_834);
nand U2567 (N_2567,N_2376,N_1714);
xor U2568 (N_2568,N_1562,N_1013);
nor U2569 (N_2569,N_656,N_689);
xor U2570 (N_2570,N_283,N_2063);
nand U2571 (N_2571,N_1145,N_986);
and U2572 (N_2572,N_1769,N_818);
nand U2573 (N_2573,N_2175,N_2004);
nor U2574 (N_2574,N_785,N_1931);
and U2575 (N_2575,N_58,N_853);
nand U2576 (N_2576,N_458,N_2314);
nand U2577 (N_2577,N_1125,N_86);
nand U2578 (N_2578,N_635,N_630);
or U2579 (N_2579,N_705,N_1956);
xnor U2580 (N_2580,N_268,N_2407);
xor U2581 (N_2581,N_424,N_234);
and U2582 (N_2582,N_1985,N_2392);
or U2583 (N_2583,N_1498,N_2069);
or U2584 (N_2584,N_959,N_1691);
nor U2585 (N_2585,N_1163,N_2243);
nand U2586 (N_2586,N_1374,N_1067);
xor U2587 (N_2587,N_631,N_509);
nand U2588 (N_2588,N_915,N_296);
nor U2589 (N_2589,N_1332,N_888);
and U2590 (N_2590,N_661,N_1699);
xor U2591 (N_2591,N_492,N_1754);
or U2592 (N_2592,N_2014,N_276);
and U2593 (N_2593,N_2120,N_1259);
nand U2594 (N_2594,N_849,N_562);
and U2595 (N_2595,N_974,N_511);
or U2596 (N_2596,N_1362,N_96);
nor U2597 (N_2597,N_2010,N_2062);
nand U2598 (N_2598,N_1668,N_2327);
or U2599 (N_2599,N_1269,N_2340);
nor U2600 (N_2600,N_730,N_2020);
nand U2601 (N_2601,N_1441,N_266);
xnor U2602 (N_2602,N_1572,N_1779);
nor U2603 (N_2603,N_228,N_2436);
and U2604 (N_2604,N_1701,N_465);
or U2605 (N_2605,N_2439,N_1043);
and U2606 (N_2606,N_297,N_333);
or U2607 (N_2607,N_129,N_72);
nor U2608 (N_2608,N_1174,N_1762);
nor U2609 (N_2609,N_1688,N_1373);
nor U2610 (N_2610,N_2305,N_2289);
nor U2611 (N_2611,N_1360,N_1087);
or U2612 (N_2612,N_230,N_1740);
nor U2613 (N_2613,N_636,N_1835);
nand U2614 (N_2614,N_1866,N_1965);
nand U2615 (N_2615,N_1932,N_1935);
or U2616 (N_2616,N_668,N_1066);
and U2617 (N_2617,N_1490,N_1518);
or U2618 (N_2618,N_698,N_182);
or U2619 (N_2619,N_1184,N_2344);
or U2620 (N_2620,N_2185,N_2323);
nor U2621 (N_2621,N_1406,N_1817);
nand U2622 (N_2622,N_2149,N_2419);
and U2623 (N_2623,N_1068,N_1283);
xor U2624 (N_2624,N_1496,N_1475);
nand U2625 (N_2625,N_1781,N_1504);
nand U2626 (N_2626,N_575,N_799);
or U2627 (N_2627,N_859,N_1032);
nor U2628 (N_2628,N_1534,N_136);
nand U2629 (N_2629,N_105,N_755);
and U2630 (N_2630,N_78,N_100);
or U2631 (N_2631,N_1274,N_1346);
and U2632 (N_2632,N_2059,N_253);
or U2633 (N_2633,N_1594,N_643);
and U2634 (N_2634,N_886,N_1164);
and U2635 (N_2635,N_1318,N_213);
nor U2636 (N_2636,N_176,N_2496);
nand U2637 (N_2637,N_2139,N_1343);
nand U2638 (N_2638,N_1017,N_1268);
and U2639 (N_2639,N_316,N_1695);
xnor U2640 (N_2640,N_2230,N_655);
and U2641 (N_2641,N_2355,N_1213);
and U2642 (N_2642,N_1419,N_2405);
or U2643 (N_2643,N_1160,N_1683);
nor U2644 (N_2644,N_1905,N_1025);
or U2645 (N_2645,N_1151,N_1199);
or U2646 (N_2646,N_2271,N_952);
nor U2647 (N_2647,N_1107,N_657);
nand U2648 (N_2648,N_776,N_1860);
nor U2649 (N_2649,N_2117,N_325);
and U2650 (N_2650,N_1838,N_203);
nand U2651 (N_2651,N_1859,N_1773);
and U2652 (N_2652,N_497,N_1673);
and U2653 (N_2653,N_1077,N_178);
or U2654 (N_2654,N_2077,N_2479);
nand U2655 (N_2655,N_104,N_1509);
nand U2656 (N_2656,N_1542,N_1885);
xnor U2657 (N_2657,N_1661,N_361);
and U2658 (N_2658,N_2259,N_1605);
nand U2659 (N_2659,N_2430,N_2125);
or U2660 (N_2660,N_98,N_814);
or U2661 (N_2661,N_2330,N_1638);
and U2662 (N_2662,N_110,N_194);
or U2663 (N_2663,N_1720,N_1870);
nor U2664 (N_2664,N_1624,N_548);
and U2665 (N_2665,N_79,N_2084);
nor U2666 (N_2666,N_700,N_1925);
xnor U2667 (N_2667,N_2241,N_1225);
nor U2668 (N_2668,N_1705,N_475);
and U2669 (N_2669,N_352,N_1815);
nor U2670 (N_2670,N_1726,N_2052);
xor U2671 (N_2671,N_1868,N_116);
and U2672 (N_2672,N_1791,N_94);
nand U2673 (N_2673,N_795,N_1864);
and U2674 (N_2674,N_2255,N_1823);
nor U2675 (N_2675,N_1016,N_1396);
nand U2676 (N_2676,N_271,N_20);
or U2677 (N_2677,N_1055,N_1982);
nor U2678 (N_2678,N_2491,N_2245);
or U2679 (N_2679,N_1584,N_1526);
nor U2680 (N_2680,N_1963,N_1124);
nor U2681 (N_2681,N_2450,N_593);
or U2682 (N_2682,N_897,N_320);
nand U2683 (N_2683,N_434,N_843);
nand U2684 (N_2684,N_808,N_1926);
or U2685 (N_2685,N_993,N_1139);
nor U2686 (N_2686,N_1631,N_374);
or U2687 (N_2687,N_1763,N_2232);
nand U2688 (N_2688,N_1429,N_1214);
or U2689 (N_2689,N_1824,N_580);
and U2690 (N_2690,N_63,N_1685);
and U2691 (N_2691,N_2,N_2143);
nor U2692 (N_2692,N_1376,N_715);
and U2693 (N_2693,N_2096,N_2132);
or U2694 (N_2694,N_651,N_1286);
xor U2695 (N_2695,N_977,N_910);
nor U2696 (N_2696,N_512,N_2391);
nor U2697 (N_2697,N_2022,N_1976);
nor U2698 (N_2698,N_852,N_1774);
and U2699 (N_2699,N_1521,N_1143);
and U2700 (N_2700,N_156,N_911);
or U2701 (N_2701,N_2473,N_2116);
xnor U2702 (N_2702,N_945,N_2028);
xnor U2703 (N_2703,N_1715,N_2320);
nand U2704 (N_2704,N_844,N_321);
nand U2705 (N_2705,N_24,N_1233);
nand U2706 (N_2706,N_347,N_967);
nor U2707 (N_2707,N_699,N_644);
nand U2708 (N_2708,N_2181,N_2451);
and U2709 (N_2709,N_2445,N_1460);
nand U2710 (N_2710,N_1201,N_2017);
nand U2711 (N_2711,N_2070,N_1871);
nand U2712 (N_2712,N_1748,N_2016);
nand U2713 (N_2713,N_341,N_56);
nor U2714 (N_2714,N_282,N_1023);
or U2715 (N_2715,N_1883,N_418);
nand U2716 (N_2716,N_145,N_893);
nand U2717 (N_2717,N_561,N_1123);
nand U2718 (N_2718,N_451,N_816);
or U2719 (N_2719,N_827,N_981);
nor U2720 (N_2720,N_1152,N_2466);
or U2721 (N_2721,N_2201,N_1492);
xor U2722 (N_2722,N_2262,N_1601);
xor U2723 (N_2723,N_2055,N_528);
or U2724 (N_2724,N_1867,N_2060);
xnor U2725 (N_2725,N_128,N_842);
nand U2726 (N_2726,N_1195,N_652);
nor U2727 (N_2727,N_1249,N_215);
nand U2728 (N_2728,N_1315,N_1091);
and U2729 (N_2729,N_1940,N_1877);
nand U2730 (N_2730,N_836,N_427);
and U2731 (N_2731,N_117,N_982);
or U2732 (N_2732,N_70,N_1153);
or U2733 (N_2733,N_556,N_1044);
nor U2734 (N_2734,N_461,N_1995);
or U2735 (N_2735,N_1957,N_1005);
or U2736 (N_2736,N_1060,N_1807);
or U2737 (N_2737,N_873,N_1592);
xor U2738 (N_2738,N_759,N_1928);
and U2739 (N_2739,N_1863,N_778);
or U2740 (N_2740,N_680,N_906);
and U2741 (N_2741,N_809,N_1743);
nor U2742 (N_2742,N_1072,N_2111);
nand U2743 (N_2743,N_902,N_480);
nor U2744 (N_2744,N_2115,N_210);
nand U2745 (N_2745,N_1056,N_1372);
xnor U2746 (N_2746,N_1747,N_694);
or U2747 (N_2747,N_1949,N_976);
nand U2748 (N_2748,N_264,N_924);
and U2749 (N_2749,N_254,N_149);
nand U2750 (N_2750,N_304,N_415);
nand U2751 (N_2751,N_1325,N_696);
or U2752 (N_2752,N_1390,N_542);
nand U2753 (N_2753,N_1892,N_1166);
nor U2754 (N_2754,N_52,N_483);
nand U2755 (N_2755,N_903,N_436);
and U2756 (N_2756,N_2295,N_731);
nand U2757 (N_2757,N_2308,N_1464);
or U2758 (N_2758,N_1793,N_1497);
nor U2759 (N_2759,N_1818,N_1583);
and U2760 (N_2760,N_170,N_2408);
or U2761 (N_2761,N_1992,N_1543);
or U2762 (N_2762,N_1796,N_33);
and U2763 (N_2763,N_274,N_380);
xor U2764 (N_2764,N_1567,N_1974);
nand U2765 (N_2765,N_2127,N_912);
or U2766 (N_2766,N_1742,N_1856);
nor U2767 (N_2767,N_1917,N_729);
and U2768 (N_2768,N_1819,N_1207);
nor U2769 (N_2769,N_627,N_1188);
or U2770 (N_2770,N_1425,N_1208);
nand U2771 (N_2771,N_2129,N_1338);
nand U2772 (N_2772,N_219,N_309);
nand U2773 (N_2773,N_1644,N_2388);
nand U2774 (N_2774,N_15,N_1553);
and U2775 (N_2775,N_1626,N_2264);
xor U2776 (N_2776,N_591,N_32);
nand U2777 (N_2777,N_2247,N_1099);
xor U2778 (N_2778,N_598,N_856);
or U2779 (N_2779,N_1936,N_181);
nand U2780 (N_2780,N_1921,N_1181);
xor U2781 (N_2781,N_633,N_1451);
nor U2782 (N_2782,N_944,N_1478);
or U2783 (N_2783,N_2048,N_1457);
nand U2784 (N_2784,N_1435,N_1218);
nand U2785 (N_2785,N_691,N_1198);
and U2786 (N_2786,N_1062,N_933);
nor U2787 (N_2787,N_490,N_1482);
nor U2788 (N_2788,N_1299,N_1680);
or U2789 (N_2789,N_1535,N_13);
or U2790 (N_2790,N_1453,N_2480);
nor U2791 (N_2791,N_1573,N_1663);
nand U2792 (N_2792,N_1275,N_450);
and U2793 (N_2793,N_2180,N_95);
and U2794 (N_2794,N_407,N_1317);
nor U2795 (N_2795,N_21,N_2394);
nand U2796 (N_2796,N_572,N_2218);
nor U2797 (N_2797,N_1412,N_1432);
and U2798 (N_2798,N_2402,N_1570);
nor U2799 (N_2799,N_187,N_47);
nand U2800 (N_2800,N_81,N_2036);
nand U2801 (N_2801,N_1065,N_1280);
nor U2802 (N_2802,N_35,N_820);
and U2803 (N_2803,N_124,N_1488);
or U2804 (N_2804,N_2279,N_1404);
or U2805 (N_2805,N_375,N_1057);
nor U2806 (N_2806,N_2409,N_302);
and U2807 (N_2807,N_870,N_1019);
and U2808 (N_2808,N_1349,N_2076);
nand U2809 (N_2809,N_357,N_2382);
or U2810 (N_2810,N_517,N_1293);
or U2811 (N_2811,N_1313,N_183);
nand U2812 (N_2812,N_447,N_348);
or U2813 (N_2813,N_2399,N_898);
nand U2814 (N_2814,N_1845,N_2119);
or U2815 (N_2815,N_1434,N_854);
xor U2816 (N_2816,N_1331,N_90);
or U2817 (N_2817,N_2341,N_2336);
nor U2818 (N_2818,N_980,N_1851);
or U2819 (N_2819,N_2104,N_2137);
nand U2820 (N_2820,N_1713,N_1884);
or U2821 (N_2821,N_392,N_2114);
or U2822 (N_2822,N_67,N_467);
or U2823 (N_2823,N_2487,N_1557);
nor U2824 (N_2824,N_1386,N_1508);
nand U2825 (N_2825,N_241,N_2265);
nor U2826 (N_2826,N_1989,N_1115);
nor U2827 (N_2827,N_1121,N_577);
xnor U2828 (N_2828,N_399,N_2001);
and U2829 (N_2829,N_269,N_750);
nor U2830 (N_2830,N_299,N_714);
or U2831 (N_2831,N_864,N_331);
nand U2832 (N_2832,N_1827,N_1944);
xnor U2833 (N_2833,N_227,N_1576);
or U2834 (N_2834,N_2133,N_36);
and U2835 (N_2835,N_2296,N_148);
or U2836 (N_2836,N_1290,N_516);
or U2837 (N_2837,N_1565,N_165);
and U2838 (N_2838,N_45,N_2403);
and U2839 (N_2839,N_603,N_2126);
or U2840 (N_2840,N_491,N_1972);
nand U2841 (N_2841,N_588,N_494);
nor U2842 (N_2842,N_365,N_1398);
nand U2843 (N_2843,N_1327,N_1671);
nor U2844 (N_2844,N_1383,N_760);
or U2845 (N_2845,N_943,N_1209);
nand U2846 (N_2846,N_584,N_1772);
nor U2847 (N_2847,N_616,N_994);
xnor U2848 (N_2848,N_679,N_1878);
or U2849 (N_2849,N_144,N_560);
and U2850 (N_2850,N_2188,N_289);
and U2851 (N_2851,N_1907,N_2363);
nor U2852 (N_2852,N_770,N_597);
or U2853 (N_2853,N_293,N_1582);
nor U2854 (N_2854,N_1459,N_1569);
and U2855 (N_2855,N_1837,N_80);
and U2856 (N_2856,N_416,N_1920);
nand U2857 (N_2857,N_1264,N_558);
or U2858 (N_2858,N_2307,N_526);
nand U2859 (N_2859,N_1623,N_11);
and U2860 (N_2860,N_1030,N_586);
xor U2861 (N_2861,N_524,N_1975);
and U2862 (N_2862,N_1222,N_1697);
or U2863 (N_2863,N_2426,N_874);
xor U2864 (N_2864,N_1880,N_2142);
and U2865 (N_2865,N_1456,N_242);
and U2866 (N_2866,N_544,N_1971);
xnor U2867 (N_2867,N_666,N_438);
or U2868 (N_2868,N_85,N_123);
or U2869 (N_2869,N_1096,N_1910);
nand U2870 (N_2870,N_1347,N_501);
or U2871 (N_2871,N_1825,N_231);
and U2872 (N_2872,N_1090,N_2103);
or U2873 (N_2873,N_42,N_1051);
nor U2874 (N_2874,N_367,N_1061);
xnor U2875 (N_2875,N_1258,N_18);
or U2876 (N_2876,N_1081,N_688);
or U2877 (N_2877,N_1901,N_1194);
nand U2878 (N_2878,N_1128,N_1706);
nand U2879 (N_2879,N_1639,N_692);
nor U2880 (N_2880,N_1756,N_1967);
nand U2881 (N_2881,N_724,N_2280);
or U2882 (N_2882,N_394,N_99);
or U2883 (N_2883,N_281,N_2113);
or U2884 (N_2884,N_946,N_1950);
or U2885 (N_2885,N_1462,N_1105);
nor U2886 (N_2886,N_2097,N_1585);
and U2887 (N_2887,N_1606,N_1448);
nand U2888 (N_2888,N_151,N_2182);
nand U2889 (N_2889,N_518,N_34);
and U2890 (N_2890,N_1618,N_1024);
nand U2891 (N_2891,N_150,N_2358);
nand U2892 (N_2892,N_1197,N_1118);
or U2893 (N_2893,N_960,N_2226);
xor U2894 (N_2894,N_1794,N_48);
and U2895 (N_2895,N_1552,N_1006);
and U2896 (N_2896,N_1089,N_286);
and U2897 (N_2897,N_419,N_1158);
or U2898 (N_2898,N_1555,N_2150);
and U2899 (N_2899,N_935,N_1896);
nand U2900 (N_2900,N_1000,N_909);
nand U2901 (N_2901,N_1244,N_2002);
nor U2902 (N_2902,N_1245,N_198);
nor U2903 (N_2903,N_954,N_1337);
nor U2904 (N_2904,N_405,N_953);
or U2905 (N_2905,N_1586,N_617);
and U2906 (N_2906,N_948,N_1046);
or U2907 (N_2907,N_1517,N_1465);
and U2908 (N_2908,N_638,N_1150);
nand U2909 (N_2909,N_312,N_2298);
and U2910 (N_2910,N_313,N_2197);
or U2911 (N_2911,N_1034,N_740);
xor U2912 (N_2912,N_334,N_1765);
nor U2913 (N_2913,N_904,N_2091);
nor U2914 (N_2914,N_335,N_1830);
nor U2915 (N_2915,N_384,N_1531);
or U2916 (N_2916,N_793,N_892);
nand U2917 (N_2917,N_847,N_1294);
or U2918 (N_2918,N_69,N_2156);
and U2919 (N_2919,N_2172,N_1650);
nor U2920 (N_2920,N_2095,N_2217);
and U2921 (N_2921,N_1252,N_1784);
and U2922 (N_2922,N_1523,N_2442);
and U2923 (N_2923,N_439,N_409);
nand U2924 (N_2924,N_2406,N_2166);
or U2925 (N_2925,N_1368,N_1733);
nand U2926 (N_2926,N_239,N_576);
nor U2927 (N_2927,N_772,N_1799);
nand U2928 (N_2928,N_172,N_248);
nand U2929 (N_2929,N_662,N_673);
or U2930 (N_2930,N_485,N_1271);
nand U2931 (N_2931,N_1402,N_163);
nor U2932 (N_2932,N_670,N_410);
and U2933 (N_2933,N_790,N_1395);
or U2934 (N_2934,N_663,N_634);
and U2935 (N_2935,N_2207,N_2362);
nand U2936 (N_2936,N_1148,N_127);
nor U2937 (N_2937,N_1205,N_1083);
and U2938 (N_2938,N_1603,N_681);
nand U2939 (N_2939,N_2089,N_498);
nand U2940 (N_2940,N_2420,N_2455);
or U2941 (N_2941,N_1662,N_2370);
or U2942 (N_2942,N_830,N_1446);
or U2943 (N_2943,N_2404,N_962);
or U2944 (N_2944,N_495,N_2495);
or U2945 (N_2945,N_1106,N_777);
nand U2946 (N_2946,N_1723,N_5);
nor U2947 (N_2947,N_1361,N_1649);
nand U2948 (N_2948,N_1022,N_1127);
and U2949 (N_2949,N_1304,N_1282);
or U2950 (N_2950,N_860,N_398);
nand U2951 (N_2951,N_1547,N_1216);
nor U2952 (N_2952,N_520,N_1516);
or U2953 (N_2953,N_2009,N_493);
and U2954 (N_2954,N_768,N_1767);
nor U2955 (N_2955,N_791,N_894);
and U2956 (N_2956,N_2481,N_1417);
xor U2957 (N_2957,N_1173,N_2231);
or U2958 (N_2958,N_1560,N_1597);
nand U2959 (N_2959,N_457,N_1011);
xor U2960 (N_2960,N_103,N_1073);
nand U2961 (N_2961,N_93,N_1080);
nand U2962 (N_2962,N_1745,N_2347);
nor U2963 (N_2963,N_1937,N_1832);
nand U2964 (N_2964,N_2177,N_471);
nor U2965 (N_2965,N_1728,N_1862);
and U2966 (N_2966,N_159,N_1602);
and U2967 (N_2967,N_857,N_472);
nor U2968 (N_2968,N_921,N_2401);
and U2969 (N_2969,N_2270,N_1161);
nor U2970 (N_2970,N_2049,N_1082);
nand U2971 (N_2971,N_2053,N_1996);
and U2972 (N_2972,N_1130,N_2469);
xor U2973 (N_2973,N_1176,N_332);
nand U2974 (N_2974,N_1549,N_1436);
and U2975 (N_2975,N_314,N_2353);
nand U2976 (N_2976,N_2338,N_292);
or U2977 (N_2977,N_525,N_2190);
nor U2978 (N_2978,N_473,N_1039);
and U2979 (N_2979,N_1698,N_1502);
nor U2980 (N_2980,N_2332,N_2488);
or U2981 (N_2981,N_1297,N_1421);
xnor U2982 (N_2982,N_1223,N_1110);
nand U2983 (N_2983,N_1276,N_319);
or U2984 (N_2984,N_1169,N_2396);
or U2985 (N_2985,N_1033,N_1408);
nand U2986 (N_2986,N_939,N_449);
nor U2987 (N_2987,N_1758,N_2274);
or U2988 (N_2988,N_2007,N_1979);
nand U2989 (N_2989,N_1563,N_1643);
nand U2990 (N_2990,N_2251,N_1546);
and U2991 (N_2991,N_2220,N_2141);
xor U2992 (N_2992,N_1770,N_2173);
or U2993 (N_2993,N_1693,N_841);
nor U2994 (N_2994,N_2041,N_914);
or U2995 (N_2995,N_1647,N_1635);
or U2996 (N_2996,N_1718,N_723);
nand U2997 (N_2997,N_126,N_660);
nand U2998 (N_2998,N_1734,N_28);
nand U2999 (N_2999,N_1443,N_1566);
nor U3000 (N_3000,N_161,N_1933);
or U3001 (N_3001,N_806,N_1394);
nand U3002 (N_3002,N_2378,N_1849);
xor U3003 (N_3003,N_2395,N_1886);
and U3004 (N_3004,N_1064,N_1146);
nand U3005 (N_3005,N_456,N_1589);
nand U3006 (N_3006,N_2412,N_2275);
or U3007 (N_3007,N_311,N_383);
nand U3008 (N_3008,N_581,N_166);
or U3009 (N_3009,N_2191,N_503);
or U3010 (N_3010,N_2294,N_2068);
and U3011 (N_3011,N_29,N_2209);
nor U3012 (N_3012,N_265,N_664);
nor U3013 (N_3013,N_1311,N_1595);
nor U3014 (N_3014,N_1147,N_1367);
and U3015 (N_3015,N_1593,N_1241);
nand U3016 (N_3016,N_2301,N_2387);
nor U3017 (N_3017,N_1112,N_2422);
nand U3018 (N_3018,N_1889,N_1804);
or U3019 (N_3019,N_2319,N_650);
nand U3020 (N_3020,N_345,N_1183);
nand U3021 (N_3021,N_2386,N_68);
nand U3022 (N_3022,N_250,N_324);
nor U3023 (N_3023,N_725,N_2484);
and U3024 (N_3024,N_1029,N_557);
and U3025 (N_3025,N_1575,N_1263);
or U3026 (N_3026,N_354,N_973);
and U3027 (N_3027,N_1776,N_477);
and U3028 (N_3028,N_1461,N_1608);
xnor U3029 (N_3029,N_428,N_2474);
and U3030 (N_3030,N_955,N_788);
xor U3031 (N_3031,N_779,N_2054);
or U3032 (N_3032,N_2123,N_2263);
nor U3033 (N_3033,N_887,N_2081);
and U3034 (N_3034,N_111,N_2210);
and U3035 (N_3035,N_1345,N_1749);
xor U3036 (N_3036,N_2183,N_1165);
xnor U3037 (N_3037,N_364,N_113);
and U3038 (N_3038,N_1186,N_592);
or U3039 (N_3039,N_890,N_211);
or U3040 (N_3040,N_2074,N_209);
and U3041 (N_3041,N_235,N_1525);
nand U3042 (N_3042,N_824,N_889);
nor U3043 (N_3043,N_1812,N_837);
and U3044 (N_3044,N_1709,N_1981);
or U3045 (N_3045,N_1841,N_275);
xnor U3046 (N_3046,N_753,N_1287);
and U3047 (N_3047,N_866,N_2499);
nor U3048 (N_3048,N_2078,N_845);
and U3049 (N_3049,N_2287,N_1308);
or U3050 (N_3050,N_486,N_2266);
and U3051 (N_3051,N_2008,N_487);
or U3052 (N_3052,N_1681,N_1364);
and U3053 (N_3053,N_1738,N_1717);
or U3054 (N_3054,N_1993,N_787);
and U3055 (N_3055,N_2064,N_46);
and U3056 (N_3056,N_1433,N_2187);
and U3057 (N_3057,N_2393,N_743);
and U3058 (N_3058,N_37,N_1619);
or U3059 (N_3059,N_14,N_1848);
nand U3060 (N_3060,N_1675,N_2493);
nand U3061 (N_3061,N_1366,N_1193);
nand U3062 (N_3062,N_185,N_2027);
and U3063 (N_3063,N_2380,N_1038);
and U3064 (N_3064,N_1800,N_716);
xnor U3065 (N_3065,N_1527,N_559);
nor U3066 (N_3066,N_880,N_2267);
nand U3067 (N_3067,N_1865,N_1466);
and U3068 (N_3068,N_1797,N_192);
nand U3069 (N_3069,N_2024,N_1312);
or U3070 (N_3070,N_1753,N_2431);
and U3071 (N_3071,N_77,N_130);
and U3072 (N_3072,N_158,N_1633);
nand U3073 (N_3073,N_1915,N_757);
nand U3074 (N_3074,N_162,N_1810);
xor U3075 (N_3075,N_83,N_1512);
and U3076 (N_3076,N_377,N_462);
and U3077 (N_3077,N_571,N_2212);
and U3078 (N_3078,N_91,N_2213);
nand U3079 (N_3079,N_1536,N_858);
or U3080 (N_3080,N_878,N_622);
nor U3081 (N_3081,N_1686,N_2331);
nor U3082 (N_3082,N_1484,N_1872);
and U3083 (N_3083,N_2321,N_1840);
and U3084 (N_3084,N_2427,N_2176);
and U3085 (N_3085,N_539,N_530);
xor U3086 (N_3086,N_810,N_1256);
nor U3087 (N_3087,N_896,N_1806);
and U3088 (N_3088,N_1588,N_1945);
nand U3089 (N_3089,N_1265,N_771);
nor U3090 (N_3090,N_247,N_833);
nor U3091 (N_3091,N_1759,N_1604);
or U3092 (N_3092,N_1070,N_2444);
and U3093 (N_3093,N_1899,N_602);
nor U3094 (N_3094,N_1356,N_532);
xor U3095 (N_3095,N_1326,N_1777);
nand U3096 (N_3096,N_189,N_322);
nand U3097 (N_3097,N_519,N_84);
and U3098 (N_3098,N_400,N_2494);
or U3099 (N_3099,N_1574,N_2367);
or U3100 (N_3100,N_2244,N_306);
or U3101 (N_3101,N_1532,N_667);
nor U3102 (N_3102,N_579,N_961);
nand U3103 (N_3103,N_905,N_479);
xor U3104 (N_3104,N_1544,N_329);
or U3105 (N_3105,N_2277,N_950);
and U3106 (N_3106,N_1687,N_999);
and U3107 (N_3107,N_1564,N_1904);
nand U3108 (N_3108,N_645,N_741);
xor U3109 (N_3109,N_1157,N_1873);
xnor U3110 (N_3110,N_260,N_1440);
nor U3111 (N_3111,N_883,N_1339);
and U3112 (N_3112,N_1300,N_1538);
or U3113 (N_3113,N_366,N_184);
and U3114 (N_3114,N_1141,N_885);
and U3115 (N_3115,N_2434,N_263);
nor U3116 (N_3116,N_2051,N_678);
or U3117 (N_3117,N_1998,N_425);
or U3118 (N_3118,N_940,N_344);
or U3119 (N_3119,N_262,N_1385);
nor U3120 (N_3120,N_1923,N_443);
xor U3121 (N_3121,N_1004,N_867);
or U3122 (N_3122,N_2257,N_1215);
nand U3123 (N_3123,N_76,N_1015);
nand U3124 (N_3124,N_140,N_1637);
xor U3125 (N_3125,N_1778,N_932);
nor U3126 (N_3126,N_1177,N_1820);
nor U3127 (N_3127,N_60,N_1003);
nor U3128 (N_3128,N_742,N_1514);
or U3129 (N_3129,N_2297,N_1008);
or U3130 (N_3130,N_1939,N_1510);
nand U3131 (N_3131,N_1175,N_975);
xnor U3132 (N_3132,N_1846,N_1371);
nand U3133 (N_3133,N_1405,N_318);
nand U3134 (N_3134,N_1036,N_800);
xnor U3135 (N_3135,N_204,N_2348);
nor U3136 (N_3136,N_2071,N_1210);
and U3137 (N_3137,N_1511,N_1918);
or U3138 (N_3138,N_2223,N_330);
nor U3139 (N_3139,N_2417,N_1515);
nor U3140 (N_3140,N_1874,N_737);
and U3141 (N_3141,N_1254,N_1735);
nor U3142 (N_3142,N_2169,N_4);
nand U3143 (N_3143,N_1955,N_31);
or U3144 (N_3144,N_2160,N_2174);
xnor U3145 (N_3145,N_1370,N_2476);
and U3146 (N_3146,N_1612,N_1237);
or U3147 (N_3147,N_1375,N_221);
nand U3148 (N_3148,N_417,N_2248);
and U3149 (N_3149,N_1250,N_1301);
or U3150 (N_3150,N_695,N_22);
nand U3151 (N_3151,N_1577,N_1500);
nor U3152 (N_3152,N_1014,N_1634);
and U3153 (N_3153,N_825,N_2222);
xnor U3154 (N_3154,N_745,N_876);
nand U3155 (N_3155,N_2359,N_764);
or U3156 (N_3156,N_925,N_2398);
xnor U3157 (N_3157,N_533,N_1752);
nor U3158 (N_3158,N_851,N_1305);
nand U3159 (N_3159,N_301,N_391);
or U3160 (N_3160,N_2005,N_2334);
nor U3161 (N_3161,N_444,N_831);
and U3162 (N_3162,N_751,N_1958);
nor U3163 (N_3163,N_1217,N_1071);
nand U3164 (N_3164,N_376,N_2411);
xor U3165 (N_3165,N_89,N_2276);
and U3166 (N_3166,N_157,N_336);
nand U3167 (N_3167,N_1785,N_1854);
nand U3168 (N_3168,N_1621,N_2189);
nand U3169 (N_3169,N_2015,N_202);
nand U3170 (N_3170,N_108,N_64);
or U3171 (N_3171,N_2164,N_1672);
or U3172 (N_3172,N_686,N_1829);
nor U3173 (N_3173,N_1964,N_2238);
nor U3174 (N_3174,N_288,N_1192);
and U3175 (N_3175,N_1027,N_2118);
and U3176 (N_3176,N_71,N_569);
xnor U3177 (N_3177,N_214,N_1495);
and U3178 (N_3178,N_240,N_971);
or U3179 (N_3179,N_1021,N_521);
and U3180 (N_3180,N_2306,N_917);
nand U3181 (N_3181,N_684,N_1092);
or U3182 (N_3182,N_1037,N_2440);
or U3183 (N_3183,N_2153,N_1211);
or U3184 (N_3184,N_1481,N_2086);
nand U3185 (N_3185,N_442,N_583);
nand U3186 (N_3186,N_1983,N_606);
and U3187 (N_3187,N_1653,N_446);
nand U3188 (N_3188,N_1489,N_207);
nor U3189 (N_3189,N_2031,N_1990);
or U3190 (N_3190,N_464,N_789);
nand U3191 (N_3191,N_173,N_1407);
or U3192 (N_3192,N_2194,N_2202);
nand U3193 (N_3193,N_1086,N_2152);
and U3194 (N_3194,N_373,N_346);
or U3195 (N_3195,N_2157,N_2161);
nor U3196 (N_3196,N_1420,N_1437);
xor U3197 (N_3197,N_1227,N_1413);
and U3198 (N_3198,N_1929,N_685);
or U3199 (N_3199,N_1467,N_1235);
and U3200 (N_3200,N_2346,N_1960);
nor U3201 (N_3201,N_1103,N_972);
nor U3202 (N_3202,N_197,N_964);
or U3203 (N_3203,N_585,N_1212);
nor U3204 (N_3204,N_1522,N_1684);
nor U3205 (N_3205,N_609,N_1454);
or U3206 (N_3206,N_1384,N_1716);
nand U3207 (N_3207,N_2130,N_1284);
or U3208 (N_3208,N_727,N_1897);
nor U3209 (N_3209,N_1261,N_482);
nand U3210 (N_3210,N_682,N_1548);
nand U3211 (N_3211,N_773,N_747);
nor U3212 (N_3212,N_1790,N_1391);
and U3213 (N_3213,N_1135,N_2316);
nor U3214 (N_3214,N_1501,N_701);
nand U3215 (N_3215,N_1279,N_2354);
nor U3216 (N_3216,N_2342,N_1048);
and U3217 (N_3217,N_1012,N_2236);
nor U3218 (N_3218,N_2040,N_2447);
or U3219 (N_3219,N_1942,N_1098);
or U3220 (N_3220,N_2377,N_1140);
and U3221 (N_3221,N_199,N_1599);
nand U3222 (N_3222,N_908,N_1078);
and U3223 (N_3223,N_619,N_1667);
nand U3224 (N_3224,N_500,N_2170);
or U3225 (N_3225,N_1994,N_295);
nand U3226 (N_3226,N_1002,N_988);
xor U3227 (N_3227,N_489,N_2158);
nand U3228 (N_3228,N_2311,N_2075);
nand U3229 (N_3229,N_270,N_997);
and U3230 (N_3230,N_369,N_624);
and U3231 (N_3231,N_459,N_1334);
nor U3232 (N_3232,N_305,N_811);
nand U3233 (N_3233,N_2026,N_1415);
nand U3234 (N_3234,N_1260,N_1598);
or U3235 (N_3235,N_1941,N_1551);
nor U3236 (N_3236,N_1393,N_2204);
or U3237 (N_3237,N_1529,N_1132);
nand U3238 (N_3238,N_640,N_188);
or U3239 (N_3239,N_2258,N_900);
nand U3240 (N_3240,N_1220,N_1946);
nor U3241 (N_3241,N_2093,N_2140);
xnor U3242 (N_3242,N_171,N_1659);
nand U3243 (N_3243,N_1156,N_403);
nor U3244 (N_3244,N_1696,N_615);
xnor U3245 (N_3245,N_1458,N_2366);
nand U3246 (N_3246,N_1893,N_2198);
nand U3247 (N_3247,N_2151,N_823);
and U3248 (N_3248,N_1200,N_291);
or U3249 (N_3249,N_1676,N_1798);
xnor U3250 (N_3250,N_1040,N_404);
nand U3251 (N_3251,N_1519,N_2148);
or U3252 (N_3252,N_803,N_343);
xnor U3253 (N_3253,N_2448,N_1185);
or U3254 (N_3254,N_1234,N_41);
nor U3255 (N_3255,N_807,N_1679);
nor U3256 (N_3256,N_2237,N_862);
or U3257 (N_3257,N_1842,N_2468);
xor U3258 (N_3258,N_1411,N_114);
nor U3259 (N_3259,N_390,N_632);
and U3260 (N_3260,N_1224,N_901);
nand U3261 (N_3261,N_1221,N_106);
and U3262 (N_3262,N_1288,N_1813);
or U3263 (N_3263,N_1587,N_1354);
nor U3264 (N_3264,N_1614,N_2383);
or U3265 (N_3265,N_984,N_621);
nand U3266 (N_3266,N_1302,N_1900);
or U3267 (N_3267,N_393,N_738);
nand U3268 (N_3268,N_1049,N_2102);
and U3269 (N_3269,N_1528,N_1485);
and U3270 (N_3270,N_920,N_395);
or U3271 (N_3271,N_711,N_1041);
or U3272 (N_3272,N_49,N_2066);
nand U3273 (N_3273,N_1600,N_1816);
or U3274 (N_3274,N_780,N_552);
or U3275 (N_3275,N_2090,N_2292);
nand U3276 (N_3276,N_2219,N_179);
nor U3277 (N_3277,N_761,N_2326);
and U3278 (N_3278,N_1491,N_92);
nor U3279 (N_3279,N_2039,N_1470);
nand U3280 (N_3280,N_1403,N_819);
and U3281 (N_3281,N_1291,N_1187);
or U3282 (N_3282,N_2425,N_649);
and U3283 (N_3283,N_2357,N_821);
or U3284 (N_3284,N_12,N_2215);
nor U3285 (N_3285,N_735,N_1887);
xor U3286 (N_3286,N_1855,N_440);
and U3287 (N_3287,N_1890,N_1533);
nor U3288 (N_3288,N_736,N_139);
xnor U3289 (N_3289,N_1285,N_1381);
and U3290 (N_3290,N_1962,N_881);
or U3291 (N_3291,N_1330,N_899);
xor U3292 (N_3292,N_177,N_931);
or U3293 (N_3293,N_125,N_2112);
or U3294 (N_3294,N_1379,N_1028);
nor U3295 (N_3295,N_2472,N_25);
and U3296 (N_3296,N_2029,N_1323);
nor U3297 (N_3297,N_1007,N_968);
or U3298 (N_3298,N_1978,N_1788);
and U3299 (N_3299,N_2269,N_1973);
nor U3300 (N_3300,N_628,N_2414);
nor U3301 (N_3301,N_551,N_676);
nor U3302 (N_3302,N_1322,N_828);
nand U3303 (N_3303,N_53,N_1909);
nor U3304 (N_3304,N_1578,N_463);
or U3305 (N_3305,N_1811,N_1359);
nand U3306 (N_3306,N_2312,N_1392);
xnor U3307 (N_3307,N_499,N_217);
xnor U3308 (N_3308,N_351,N_2073);
nand U3309 (N_3309,N_252,N_1930);
or U3310 (N_3310,N_1243,N_798);
and U3311 (N_3311,N_2045,N_595);
nand U3312 (N_3312,N_1953,N_1808);
xnor U3313 (N_3313,N_1468,N_1182);
nor U3314 (N_3314,N_496,N_929);
and U3315 (N_3315,N_460,N_1079);
or U3316 (N_3316,N_1766,N_978);
and U3317 (N_3317,N_2124,N_2449);
and U3318 (N_3318,N_748,N_647);
nand U3319 (N_3319,N_236,N_2246);
or U3320 (N_3320,N_1190,N_488);
nand U3321 (N_3321,N_625,N_414);
or U3322 (N_3322,N_1710,N_2100);
and U3323 (N_3323,N_1414,N_372);
or U3324 (N_3324,N_120,N_522);
or U3325 (N_3325,N_2390,N_1047);
nor U3326 (N_3326,N_2486,N_1240);
xnor U3327 (N_3327,N_2205,N_1530);
and U3328 (N_3328,N_958,N_1159);
and U3329 (N_3329,N_1289,N_1646);
or U3330 (N_3330,N_2136,N_1018);
and U3331 (N_3331,N_1568,N_1178);
nand U3332 (N_3332,N_1700,N_2489);
or U3333 (N_3333,N_1111,N_815);
and U3334 (N_3334,N_712,N_429);
nand U3335 (N_3335,N_249,N_208);
nand U3336 (N_3336,N_826,N_2385);
nor U3337 (N_3337,N_2293,N_2035);
nand U3338 (N_3338,N_2131,N_2441);
and U3339 (N_3339,N_1719,N_784);
nor U3340 (N_3340,N_1266,N_1058);
or U3341 (N_3341,N_147,N_1052);
nand U3342 (N_3342,N_2044,N_2286);
nand U3343 (N_3343,N_1270,N_547);
nand U3344 (N_3344,N_437,N_1581);
nor U3345 (N_3345,N_153,N_2196);
nand U3346 (N_3346,N_1389,N_2192);
nor U3347 (N_3347,N_2290,N_1879);
or U3348 (N_3348,N_1137,N_2225);
or U3349 (N_3349,N_2252,N_1801);
or U3350 (N_3350,N_1537,N_1682);
or U3351 (N_3351,N_277,N_1296);
or U3352 (N_3352,N_2433,N_2083);
or U3353 (N_3353,N_154,N_1755);
and U3354 (N_3354,N_739,N_1377);
and U3355 (N_3355,N_218,N_2082);
nand U3356 (N_3356,N_122,N_1246);
and U3357 (N_3357,N_2038,N_1857);
or U3358 (N_3358,N_1607,N_812);
or U3359 (N_3359,N_7,N_2186);
nand U3360 (N_3360,N_1179,N_1622);
nor U3361 (N_3361,N_937,N_1363);
nor U3362 (N_3362,N_2421,N_1122);
and U3363 (N_3363,N_378,N_607);
and U3364 (N_3364,N_2461,N_66);
nor U3365 (N_3365,N_2155,N_1894);
nand U3366 (N_3366,N_1814,N_1655);
and U3367 (N_3367,N_19,N_2423);
and U3368 (N_3368,N_992,N_1479);
nor U3369 (N_3369,N_1641,N_1760);
xnor U3370 (N_3370,N_74,N_913);
or U3371 (N_3371,N_421,N_1730);
nor U3372 (N_3372,N_1154,N_1084);
or U3373 (N_3373,N_861,N_1961);
or U3374 (N_3374,N_2254,N_983);
or U3375 (N_3375,N_690,N_387);
nor U3376 (N_3376,N_261,N_502);
and U3377 (N_3377,N_26,N_484);
or U3378 (N_3378,N_1219,N_1853);
and U3379 (N_3379,N_402,N_566);
nor U3380 (N_3380,N_1020,N_1229);
or U3381 (N_3381,N_1737,N_23);
or U3382 (N_3382,N_1658,N_612);
nor U3383 (N_3383,N_2235,N_1783);
or U3384 (N_3384,N_1524,N_642);
nand U3385 (N_3385,N_869,N_1499);
nand U3386 (N_3386,N_2373,N_1255);
nor U3387 (N_3387,N_1694,N_523);
nand U3388 (N_3388,N_168,N_1826);
nor U3389 (N_3389,N_797,N_298);
nor U3390 (N_3390,N_1054,N_990);
or U3391 (N_3391,N_1142,N_435);
and U3392 (N_3392,N_963,N_339);
nand U3393 (N_3393,N_2381,N_1010);
or U3394 (N_3394,N_175,N_2477);
nand U3395 (N_3395,N_54,N_1977);
nor U3396 (N_3396,N_40,N_608);
or U3397 (N_3397,N_1919,N_610);
xnor U3398 (N_3398,N_863,N_848);
xor U3399 (N_3399,N_989,N_767);
nand U3400 (N_3400,N_538,N_2492);
or U3401 (N_3401,N_119,N_2446);
and U3402 (N_3402,N_1426,N_710);
or U3403 (N_3403,N_441,N_1924);
nand U3404 (N_3404,N_2072,N_1645);
and U3405 (N_3405,N_550,N_1171);
xor U3406 (N_3406,N_2490,N_1273);
xor U3407 (N_3407,N_1712,N_2154);
or U3408 (N_3408,N_233,N_2281);
or U3409 (N_3409,N_101,N_362);
or U3410 (N_3410,N_1615,N_2339);
nand U3411 (N_3411,N_164,N_1725);
and U3412 (N_3412,N_817,N_2043);
nor U3413 (N_3413,N_2467,N_781);
or U3414 (N_3414,N_1307,N_570);
nand U3415 (N_3415,N_97,N_1131);
or U3416 (N_3416,N_191,N_720);
nand U3417 (N_3417,N_1095,N_1450);
or U3418 (N_3418,N_601,N_360);
or U3419 (N_3419,N_1369,N_2184);
nand U3420 (N_3420,N_17,N_1134);
xor U3421 (N_3421,N_216,N_1418);
or U3422 (N_3422,N_59,N_1422);
and U3423 (N_3423,N_1954,N_474);
or U3424 (N_3424,N_9,N_326);
nand U3425 (N_3425,N_1247,N_563);
or U3426 (N_3426,N_1999,N_1353);
or U3427 (N_3427,N_956,N_541);
or U3428 (N_3428,N_82,N_1732);
and U3429 (N_3429,N_979,N_2092);
or U3430 (N_3430,N_1117,N_919);
nand U3431 (N_3431,N_251,N_2195);
xnor U3432 (N_3432,N_1991,N_2375);
and U3433 (N_3433,N_2260,N_1206);
nor U3434 (N_3434,N_2233,N_2454);
nand U3435 (N_3435,N_2356,N_2080);
nand U3436 (N_3436,N_1847,N_1520);
and U3437 (N_3437,N_2145,N_1789);
nor U3438 (N_3438,N_1678,N_756);
and U3439 (N_3439,N_432,N_687);
nor U3440 (N_3440,N_717,N_553);
and U3441 (N_3441,N_205,N_2415);
or U3442 (N_3442,N_2034,N_2099);
or U3443 (N_3443,N_1616,N_2211);
or U3444 (N_3444,N_87,N_273);
or U3445 (N_3445,N_531,N_1545);
nor U3446 (N_3446,N_2253,N_1463);
nand U3447 (N_3447,N_141,N_1226);
and U3448 (N_3448,N_1591,N_1959);
and U3449 (N_3449,N_2013,N_504);
or U3450 (N_3450,N_359,N_1951);
and U3451 (N_3451,N_2288,N_167);
or U3452 (N_3452,N_1628,N_966);
and U3453 (N_3453,N_1665,N_1952);
nor U3454 (N_3454,N_1590,N_1507);
nor U3455 (N_3455,N_350,N_1248);
nand U3456 (N_3456,N_142,N_708);
xor U3457 (N_3457,N_794,N_2094);
nand U3458 (N_3458,N_1483,N_137);
or U3459 (N_3459,N_1351,N_1129);
nand U3460 (N_3460,N_229,N_2037);
or U3461 (N_3461,N_1613,N_408);
nand U3462 (N_3462,N_1431,N_1596);
xor U3463 (N_3463,N_1670,N_43);
nand U3464 (N_3464,N_1888,N_840);
nand U3465 (N_3465,N_2478,N_895);
and U3466 (N_3466,N_1342,N_1042);
nand U3467 (N_3467,N_431,N_618);
or U3468 (N_3468,N_1739,N_2303);
nor U3469 (N_3469,N_327,N_1494);
nand U3470 (N_3470,N_877,N_2462);
nand U3471 (N_3471,N_802,N_2250);
xnor U3472 (N_3472,N_596,N_669);
nand U3473 (N_3473,N_554,N_1986);
nand U3474 (N_3474,N_132,N_1721);
and U3475 (N_3475,N_328,N_381);
and U3476 (N_3476,N_1782,N_1640);
or U3477 (N_3477,N_2032,N_1380);
nor U3478 (N_3478,N_2304,N_303);
or U3479 (N_3479,N_2109,N_2085);
and U3480 (N_3480,N_455,N_1775);
and U3481 (N_3481,N_2216,N_574);
nand U3482 (N_3482,N_1792,N_426);
xnor U3483 (N_3483,N_1895,N_671);
nand U3484 (N_3484,N_115,N_907);
or U3485 (N_3485,N_951,N_2413);
or U3486 (N_3486,N_871,N_3);
nand U3487 (N_3487,N_1648,N_775);
and U3488 (N_3488,N_2224,N_1660);
nor U3489 (N_3489,N_1833,N_1741);
nor U3490 (N_3490,N_1674,N_272);
xnor U3491 (N_3491,N_1189,N_430);
xor U3492 (N_3492,N_1828,N_1324);
xnor U3493 (N_3493,N_2128,N_2465);
and U3494 (N_3494,N_226,N_1348);
nor U3495 (N_3495,N_1298,N_549);
or U3496 (N_3496,N_1120,N_1802);
nand U3497 (N_3497,N_1113,N_1410);
and U3498 (N_3498,N_1382,N_1844);
or U3499 (N_3499,N_2134,N_1882);
nor U3500 (N_3500,N_1321,N_1045);
or U3501 (N_3501,N_2098,N_2272);
and U3502 (N_3502,N_1009,N_674);
and U3503 (N_3503,N_1968,N_1319);
nor U3504 (N_3504,N_1116,N_481);
or U3505 (N_3505,N_2122,N_2322);
xor U3506 (N_3506,N_1262,N_693);
nand U3507 (N_3507,N_55,N_1609);
nand U3508 (N_3508,N_2121,N_2325);
and U3509 (N_3509,N_613,N_506);
or U3510 (N_3510,N_1357,N_2057);
or U3511 (N_3511,N_2498,N_2459);
nand U3512 (N_3512,N_822,N_193);
and U3513 (N_3513,N_2079,N_2019);
and U3514 (N_3514,N_1541,N_505);
xnor U3515 (N_3515,N_65,N_2299);
and U3516 (N_3516,N_44,N_1746);
xor U3517 (N_3517,N_406,N_1780);
nand U3518 (N_3518,N_2464,N_604);
nand U3519 (N_3519,N_1704,N_1409);
nand U3520 (N_3520,N_1442,N_2067);
and U3521 (N_3521,N_1100,N_1306);
or U3522 (N_3522,N_1610,N_1074);
or U3523 (N_3523,N_2256,N_1387);
nand U3524 (N_3524,N_1611,N_1831);
nor U3525 (N_3525,N_1554,N_1632);
and U3526 (N_3526,N_1035,N_195);
and U3527 (N_3527,N_1,N_1423);
nor U3528 (N_3528,N_2352,N_1328);
nand U3529 (N_3529,N_1278,N_1329);
nand U3530 (N_3530,N_138,N_294);
xnor U3531 (N_3531,N_355,N_1314);
and U3532 (N_3532,N_1102,N_865);
nor U3533 (N_3533,N_1388,N_470);
xor U3534 (N_3534,N_411,N_317);
and U3535 (N_3535,N_1168,N_0);
nand U3536 (N_3536,N_1861,N_1876);
and U3537 (N_3537,N_2234,N_792);
and U3538 (N_3538,N_39,N_683);
and U3539 (N_3539,N_1447,N_212);
or U3540 (N_3540,N_2324,N_396);
or U3541 (N_3541,N_1505,N_629);
nand U3542 (N_3542,N_2228,N_1063);
xnor U3543 (N_3543,N_1242,N_2011);
and U3544 (N_3544,N_1666,N_1677);
nor U3545 (N_3545,N_1757,N_2333);
or U3546 (N_3546,N_363,N_267);
xor U3547 (N_3547,N_782,N_1295);
or U3548 (N_3548,N_2227,N_2350);
and U3549 (N_3549,N_1803,N_805);
and U3550 (N_3550,N_2379,N_2214);
and U3551 (N_3551,N_469,N_2171);
nor U3552 (N_3552,N_1493,N_589);
nor U3553 (N_3553,N_412,N_2389);
and U3554 (N_3554,N_358,N_578);
nor U3555 (N_3555,N_2006,N_1970);
nand U3556 (N_3556,N_1703,N_1333);
and U3557 (N_3557,N_1550,N_1506);
nand U3558 (N_3558,N_1355,N_2428);
nand U3559 (N_3559,N_2437,N_1341);
xor U3560 (N_3560,N_918,N_1731);
and U3561 (N_3561,N_287,N_1559);
xnor U3562 (N_3562,N_754,N_2300);
nor U3563 (N_3563,N_1948,N_916);
and U3564 (N_3564,N_2282,N_2087);
nand U3565 (N_3565,N_323,N_510);
nor U3566 (N_3566,N_513,N_941);
nand U3567 (N_3567,N_57,N_454);
and U3568 (N_3568,N_1076,N_719);
nor U3569 (N_3569,N_928,N_2345);
or U3570 (N_3570,N_338,N_1358);
or U3571 (N_3571,N_112,N_2061);
xor U3572 (N_3572,N_2047,N_2056);
or U3573 (N_3573,N_107,N_926);
and U3574 (N_3574,N_1656,N_1891);
or U3575 (N_3575,N_2371,N_423);
nor U3576 (N_3576,N_927,N_420);
nand U3577 (N_3577,N_2193,N_555);
or U3578 (N_3578,N_453,N_1053);
or U3579 (N_3579,N_1805,N_196);
and U3580 (N_3580,N_1822,N_605);
xnor U3581 (N_3581,N_200,N_707);
and U3582 (N_3582,N_839,N_1744);
or U3583 (N_3583,N_1310,N_1630);
and U3584 (N_3584,N_1540,N_721);
nand U3585 (N_3585,N_677,N_2482);
nand U3586 (N_3586,N_991,N_2424);
and U3587 (N_3587,N_1180,N_565);
and U3588 (N_3588,N_1277,N_2485);
or U3589 (N_3589,N_1202,N_1430);
and U3590 (N_3590,N_2146,N_599);
xnor U3591 (N_3591,N_2452,N_1934);
and U3592 (N_3592,N_1272,N_257);
nand U3593 (N_3593,N_186,N_2167);
and U3594 (N_3594,N_1987,N_2058);
and U3595 (N_3595,N_2435,N_385);
nand U3596 (N_3596,N_2273,N_614);
or U3597 (N_3597,N_2088,N_1094);
nor U3598 (N_3598,N_804,N_1050);
nand U3599 (N_3599,N_654,N_564);
nand U3600 (N_3600,N_1136,N_2168);
xor U3601 (N_3601,N_1320,N_882);
xnor U3602 (N_3602,N_936,N_342);
and U3603 (N_3603,N_1503,N_573);
or U3604 (N_3604,N_949,N_734);
or U3605 (N_3605,N_746,N_623);
and U3606 (N_3606,N_1399,N_529);
xor U3607 (N_3607,N_938,N_1230);
or U3608 (N_3608,N_2483,N_1445);
nor U3609 (N_3609,N_1155,N_2178);
nand U3610 (N_3610,N_829,N_891);
nor U3611 (N_3611,N_1427,N_356);
nor U3612 (N_3612,N_1786,N_1764);
nor U3613 (N_3613,N_337,N_2206);
nor U3614 (N_3614,N_1109,N_1292);
nand U3615 (N_3615,N_1133,N_1469);
nor U3616 (N_3616,N_2000,N_478);
or U3617 (N_3617,N_1444,N_942);
nand U3618 (N_3618,N_1988,N_190);
or U3619 (N_3619,N_672,N_109);
or U3620 (N_3620,N_611,N_1836);
and U3621 (N_3621,N_2343,N_62);
or U3622 (N_3622,N_749,N_1980);
nand U3623 (N_3623,N_545,N_2315);
or U3624 (N_3624,N_813,N_445);
nand U3625 (N_3625,N_590,N_160);
nand U3626 (N_3626,N_1172,N_1898);
nor U3627 (N_3627,N_50,N_1625);
nor U3628 (N_3628,N_2458,N_1654);
nand U3629 (N_3629,N_1162,N_884);
nand U3630 (N_3630,N_2162,N_507);
nand U3631 (N_3631,N_2012,N_587);
nand U3632 (N_3632,N_2108,N_134);
or U3633 (N_3633,N_1620,N_1114);
nor U3634 (N_3634,N_1309,N_1303);
and U3635 (N_3635,N_279,N_546);
or U3636 (N_3636,N_1365,N_1167);
xor U3637 (N_3637,N_703,N_514);
nor U3638 (N_3638,N_2309,N_379);
or U3639 (N_3639,N_2438,N_1947);
nor U3640 (N_3640,N_2372,N_2397);
or U3641 (N_3641,N_675,N_1850);
and U3642 (N_3642,N_370,N_1809);
or U3643 (N_3643,N_1722,N_1881);
nor U3644 (N_3644,N_2147,N_2328);
xor U3645 (N_3645,N_468,N_1821);
xor U3646 (N_3646,N_2313,N_987);
and U3647 (N_3647,N_224,N_2471);
and U3648 (N_3648,N_1238,N_2229);
nor U3649 (N_3649,N_315,N_923);
xnor U3650 (N_3650,N_1736,N_875);
or U3651 (N_3651,N_2138,N_1476);
and U3652 (N_3652,N_1927,N_1477);
nand U3653 (N_3653,N_2364,N_1729);
nor U3654 (N_3654,N_222,N_206);
nor U3655 (N_3655,N_1424,N_1843);
xnor U3656 (N_3656,N_61,N_256);
or U3657 (N_3657,N_1711,N_245);
nor U3658 (N_3658,N_2101,N_1253);
and U3659 (N_3659,N_1473,N_476);
or U3660 (N_3660,N_1708,N_653);
nand U3661 (N_3661,N_466,N_382);
and U3662 (N_3662,N_947,N_1997);
or U3663 (N_3663,N_2365,N_1627);
or U3664 (N_3664,N_2249,N_16);
or U3665 (N_3665,N_600,N_1239);
nor U3666 (N_3666,N_243,N_1378);
xnor U3667 (N_3667,N_646,N_2261);
and U3668 (N_3668,N_639,N_2317);
nand U3669 (N_3669,N_1617,N_620);
nand U3670 (N_3670,N_284,N_1031);
nor U3671 (N_3671,N_300,N_448);
xor U3672 (N_3672,N_1651,N_201);
or U3673 (N_3673,N_769,N_2335);
or U3674 (N_3674,N_386,N_985);
nor U3675 (N_3675,N_1751,N_2203);
and U3676 (N_3676,N_1335,N_1787);
nor U3677 (N_3677,N_1579,N_1795);
and U3678 (N_3678,N_2105,N_2460);
nand U3679 (N_3679,N_718,N_515);
nand U3680 (N_3680,N_223,N_2457);
and U3681 (N_3681,N_388,N_2107);
nand U3682 (N_3682,N_2208,N_1636);
nand U3683 (N_3683,N_709,N_2318);
or U3684 (N_3684,N_2021,N_2443);
nor U3685 (N_3685,N_1486,N_765);
xnor U3686 (N_3686,N_237,N_855);
or U3687 (N_3687,N_1869,N_2470);
nand U3688 (N_3688,N_786,N_2429);
and U3689 (N_3689,N_433,N_1771);
nand U3690 (N_3690,N_308,N_1336);
nand U3691 (N_3691,N_368,N_1761);
nor U3692 (N_3692,N_255,N_2018);
and U3693 (N_3693,N_2432,N_73);
and U3694 (N_3694,N_934,N_536);
or U3695 (N_3695,N_1344,N_143);
nor U3696 (N_3696,N_1702,N_1912);
nor U3697 (N_3697,N_534,N_930);
or U3698 (N_3698,N_995,N_1689);
nor U3699 (N_3699,N_1001,N_2329);
and U3700 (N_3700,N_637,N_1561);
nand U3701 (N_3701,N_1938,N_868);
and U3702 (N_3702,N_2199,N_801);
or U3703 (N_3703,N_1707,N_2106);
and U3704 (N_3704,N_1088,N_1397);
nor U3705 (N_3705,N_665,N_713);
nor U3706 (N_3706,N_2384,N_1204);
nand U3707 (N_3707,N_2135,N_922);
nor U3708 (N_3708,N_1138,N_537);
nor U3709 (N_3709,N_1400,N_535);
nand U3710 (N_3710,N_733,N_1026);
nor U3711 (N_3711,N_998,N_1170);
xnor U3712 (N_3712,N_1472,N_2416);
and U3713 (N_3713,N_401,N_722);
xnor U3714 (N_3714,N_102,N_1474);
nand U3715 (N_3715,N_2003,N_728);
and U3716 (N_3716,N_1119,N_2374);
nand U3717 (N_3717,N_155,N_970);
nor U3718 (N_3718,N_1281,N_1340);
nor U3719 (N_3719,N_658,N_2165);
nor U3720 (N_3720,N_1916,N_1085);
xor U3721 (N_3721,N_2046,N_1416);
and U3722 (N_3722,N_2310,N_1059);
or U3723 (N_3723,N_508,N_835);
xnor U3724 (N_3724,N_146,N_220);
nor U3725 (N_3725,N_371,N_965);
and U3726 (N_3726,N_1236,N_1690);
and U3727 (N_3727,N_88,N_2456);
nand U3728 (N_3728,N_2179,N_1126);
xor U3729 (N_3729,N_957,N_180);
and U3730 (N_3730,N_1629,N_225);
xor U3731 (N_3731,N_1943,N_30);
nand U3732 (N_3732,N_2302,N_2453);
nor U3733 (N_3733,N_1487,N_1669);
nand U3734 (N_3734,N_258,N_1571);
xnor U3735 (N_3735,N_1852,N_290);
or U3736 (N_3736,N_744,N_232);
or U3737 (N_3737,N_2200,N_169);
nor U3738 (N_3738,N_2221,N_1428);
xor U3739 (N_3739,N_1966,N_2291);
or U3740 (N_3740,N_121,N_389);
and U3741 (N_3741,N_1149,N_340);
nand U3742 (N_3742,N_1513,N_2360);
and U3743 (N_3743,N_2050,N_1556);
nand U3744 (N_3744,N_397,N_1480);
and U3745 (N_3745,N_1642,N_1664);
nand U3746 (N_3746,N_969,N_2110);
or U3747 (N_3747,N_2023,N_1908);
and U3748 (N_3748,N_2042,N_1144);
nor U3749 (N_3749,N_307,N_1228);
xnor U3750 (N_3750,N_1433,N_1176);
and U3751 (N_3751,N_1234,N_997);
or U3752 (N_3752,N_1462,N_2437);
and U3753 (N_3753,N_32,N_1837);
and U3754 (N_3754,N_2437,N_1619);
xnor U3755 (N_3755,N_1477,N_433);
and U3756 (N_3756,N_1622,N_2423);
nand U3757 (N_3757,N_2307,N_1909);
or U3758 (N_3758,N_370,N_2374);
and U3759 (N_3759,N_17,N_3);
or U3760 (N_3760,N_1267,N_1205);
and U3761 (N_3761,N_388,N_1073);
and U3762 (N_3762,N_2013,N_24);
nor U3763 (N_3763,N_1899,N_1386);
nand U3764 (N_3764,N_1105,N_1446);
or U3765 (N_3765,N_1576,N_1811);
nand U3766 (N_3766,N_562,N_2369);
or U3767 (N_3767,N_1012,N_681);
xnor U3768 (N_3768,N_962,N_789);
or U3769 (N_3769,N_10,N_2466);
or U3770 (N_3770,N_436,N_1030);
nand U3771 (N_3771,N_257,N_2041);
or U3772 (N_3772,N_66,N_275);
or U3773 (N_3773,N_2336,N_265);
and U3774 (N_3774,N_1150,N_32);
and U3775 (N_3775,N_1360,N_1275);
nor U3776 (N_3776,N_155,N_936);
and U3777 (N_3777,N_1945,N_1624);
nor U3778 (N_3778,N_2164,N_1439);
and U3779 (N_3779,N_1821,N_1972);
nor U3780 (N_3780,N_1914,N_327);
nor U3781 (N_3781,N_388,N_959);
nand U3782 (N_3782,N_1522,N_207);
nand U3783 (N_3783,N_1337,N_2410);
nor U3784 (N_3784,N_1723,N_1437);
xnor U3785 (N_3785,N_2447,N_958);
or U3786 (N_3786,N_860,N_2207);
nand U3787 (N_3787,N_2372,N_1652);
nand U3788 (N_3788,N_2360,N_952);
nor U3789 (N_3789,N_61,N_1169);
nand U3790 (N_3790,N_1104,N_1113);
nand U3791 (N_3791,N_2331,N_1675);
nand U3792 (N_3792,N_643,N_1824);
xnor U3793 (N_3793,N_714,N_182);
nor U3794 (N_3794,N_614,N_679);
or U3795 (N_3795,N_841,N_467);
and U3796 (N_3796,N_94,N_1694);
or U3797 (N_3797,N_2280,N_2328);
nor U3798 (N_3798,N_391,N_203);
or U3799 (N_3799,N_1142,N_688);
and U3800 (N_3800,N_528,N_2351);
nor U3801 (N_3801,N_1194,N_1621);
or U3802 (N_3802,N_2170,N_2416);
or U3803 (N_3803,N_2476,N_973);
nand U3804 (N_3804,N_1246,N_1548);
and U3805 (N_3805,N_795,N_408);
or U3806 (N_3806,N_693,N_833);
nand U3807 (N_3807,N_1200,N_1154);
and U3808 (N_3808,N_237,N_1936);
nand U3809 (N_3809,N_88,N_1202);
xor U3810 (N_3810,N_901,N_2014);
xnor U3811 (N_3811,N_262,N_335);
or U3812 (N_3812,N_374,N_2026);
nor U3813 (N_3813,N_1385,N_210);
and U3814 (N_3814,N_1244,N_1926);
or U3815 (N_3815,N_1860,N_2410);
nor U3816 (N_3816,N_1411,N_402);
and U3817 (N_3817,N_736,N_1768);
nand U3818 (N_3818,N_1165,N_279);
or U3819 (N_3819,N_2332,N_2303);
nand U3820 (N_3820,N_138,N_399);
nand U3821 (N_3821,N_1436,N_458);
and U3822 (N_3822,N_2309,N_771);
or U3823 (N_3823,N_677,N_229);
nor U3824 (N_3824,N_1170,N_1300);
or U3825 (N_3825,N_428,N_1076);
nor U3826 (N_3826,N_1229,N_591);
or U3827 (N_3827,N_191,N_1595);
or U3828 (N_3828,N_1164,N_928);
and U3829 (N_3829,N_2457,N_2);
nor U3830 (N_3830,N_80,N_517);
nor U3831 (N_3831,N_2384,N_1214);
or U3832 (N_3832,N_2022,N_1029);
and U3833 (N_3833,N_1539,N_201);
and U3834 (N_3834,N_235,N_611);
nor U3835 (N_3835,N_954,N_338);
nor U3836 (N_3836,N_2191,N_1865);
nand U3837 (N_3837,N_2185,N_1686);
xor U3838 (N_3838,N_801,N_2417);
and U3839 (N_3839,N_1580,N_1038);
and U3840 (N_3840,N_1876,N_1854);
or U3841 (N_3841,N_1525,N_1335);
and U3842 (N_3842,N_1708,N_1273);
or U3843 (N_3843,N_725,N_2146);
nand U3844 (N_3844,N_1603,N_458);
and U3845 (N_3845,N_1889,N_1839);
nor U3846 (N_3846,N_2491,N_1939);
xnor U3847 (N_3847,N_1280,N_780);
nor U3848 (N_3848,N_503,N_527);
or U3849 (N_3849,N_1581,N_436);
and U3850 (N_3850,N_115,N_1003);
nor U3851 (N_3851,N_843,N_847);
nor U3852 (N_3852,N_1605,N_1544);
nor U3853 (N_3853,N_1927,N_2295);
and U3854 (N_3854,N_910,N_1501);
nand U3855 (N_3855,N_137,N_1258);
nor U3856 (N_3856,N_2471,N_905);
or U3857 (N_3857,N_31,N_312);
and U3858 (N_3858,N_321,N_2212);
and U3859 (N_3859,N_786,N_1409);
and U3860 (N_3860,N_814,N_2022);
nor U3861 (N_3861,N_1082,N_1812);
nor U3862 (N_3862,N_739,N_1116);
xor U3863 (N_3863,N_1382,N_727);
xor U3864 (N_3864,N_2296,N_1475);
nor U3865 (N_3865,N_1358,N_1310);
nor U3866 (N_3866,N_1811,N_1790);
and U3867 (N_3867,N_560,N_1841);
and U3868 (N_3868,N_1954,N_1065);
xnor U3869 (N_3869,N_780,N_246);
nor U3870 (N_3870,N_2176,N_2300);
nand U3871 (N_3871,N_1052,N_581);
and U3872 (N_3872,N_658,N_1415);
or U3873 (N_3873,N_1937,N_1833);
and U3874 (N_3874,N_2220,N_1249);
nor U3875 (N_3875,N_489,N_497);
and U3876 (N_3876,N_167,N_249);
nor U3877 (N_3877,N_116,N_734);
nand U3878 (N_3878,N_1737,N_1067);
or U3879 (N_3879,N_1174,N_41);
or U3880 (N_3880,N_2257,N_1814);
nand U3881 (N_3881,N_147,N_554);
and U3882 (N_3882,N_2321,N_1868);
or U3883 (N_3883,N_856,N_2420);
xor U3884 (N_3884,N_1450,N_901);
or U3885 (N_3885,N_381,N_965);
or U3886 (N_3886,N_2074,N_2094);
or U3887 (N_3887,N_1227,N_1087);
nand U3888 (N_3888,N_1614,N_1425);
nor U3889 (N_3889,N_642,N_1810);
xor U3890 (N_3890,N_1621,N_29);
nor U3891 (N_3891,N_290,N_1497);
or U3892 (N_3892,N_657,N_2055);
and U3893 (N_3893,N_225,N_2299);
or U3894 (N_3894,N_2250,N_844);
nor U3895 (N_3895,N_2053,N_2186);
and U3896 (N_3896,N_1684,N_270);
and U3897 (N_3897,N_1799,N_1468);
or U3898 (N_3898,N_695,N_2453);
or U3899 (N_3899,N_1468,N_2398);
or U3900 (N_3900,N_1303,N_1104);
nor U3901 (N_3901,N_2247,N_283);
nand U3902 (N_3902,N_425,N_962);
nor U3903 (N_3903,N_1395,N_2123);
xnor U3904 (N_3904,N_2209,N_1143);
or U3905 (N_3905,N_757,N_1762);
nand U3906 (N_3906,N_2056,N_2093);
nor U3907 (N_3907,N_730,N_407);
nand U3908 (N_3908,N_1873,N_1022);
or U3909 (N_3909,N_560,N_699);
or U3910 (N_3910,N_430,N_628);
nand U3911 (N_3911,N_2425,N_345);
nand U3912 (N_3912,N_1320,N_1460);
and U3913 (N_3913,N_2276,N_1385);
or U3914 (N_3914,N_25,N_2070);
and U3915 (N_3915,N_2059,N_1742);
and U3916 (N_3916,N_1139,N_45);
nand U3917 (N_3917,N_1849,N_346);
or U3918 (N_3918,N_2328,N_175);
and U3919 (N_3919,N_899,N_518);
nor U3920 (N_3920,N_459,N_872);
nor U3921 (N_3921,N_1358,N_2325);
or U3922 (N_3922,N_1674,N_1755);
or U3923 (N_3923,N_1957,N_1946);
nor U3924 (N_3924,N_1968,N_1667);
and U3925 (N_3925,N_715,N_1467);
nor U3926 (N_3926,N_316,N_1748);
xor U3927 (N_3927,N_594,N_959);
and U3928 (N_3928,N_702,N_176);
nand U3929 (N_3929,N_761,N_1294);
xor U3930 (N_3930,N_108,N_2284);
nand U3931 (N_3931,N_918,N_530);
nor U3932 (N_3932,N_2461,N_2104);
nand U3933 (N_3933,N_1332,N_2420);
nand U3934 (N_3934,N_480,N_1272);
or U3935 (N_3935,N_2466,N_527);
nor U3936 (N_3936,N_981,N_1920);
nand U3937 (N_3937,N_1,N_1764);
or U3938 (N_3938,N_112,N_397);
nor U3939 (N_3939,N_770,N_744);
and U3940 (N_3940,N_1846,N_770);
nand U3941 (N_3941,N_469,N_2430);
nand U3942 (N_3942,N_2439,N_1786);
and U3943 (N_3943,N_2179,N_2332);
nor U3944 (N_3944,N_1601,N_1750);
or U3945 (N_3945,N_1923,N_574);
nand U3946 (N_3946,N_607,N_1802);
nand U3947 (N_3947,N_2362,N_657);
nor U3948 (N_3948,N_727,N_2466);
or U3949 (N_3949,N_1896,N_2010);
or U3950 (N_3950,N_309,N_1528);
nor U3951 (N_3951,N_2273,N_2235);
or U3952 (N_3952,N_1638,N_2);
and U3953 (N_3953,N_1041,N_207);
nand U3954 (N_3954,N_1414,N_746);
xnor U3955 (N_3955,N_1894,N_2241);
xor U3956 (N_3956,N_987,N_2292);
or U3957 (N_3957,N_342,N_1591);
nand U3958 (N_3958,N_529,N_1293);
nor U3959 (N_3959,N_398,N_1224);
or U3960 (N_3960,N_151,N_302);
and U3961 (N_3961,N_835,N_219);
and U3962 (N_3962,N_1383,N_1713);
and U3963 (N_3963,N_267,N_1956);
or U3964 (N_3964,N_1055,N_2443);
or U3965 (N_3965,N_483,N_974);
nand U3966 (N_3966,N_1722,N_74);
nand U3967 (N_3967,N_2420,N_1674);
and U3968 (N_3968,N_1028,N_1384);
and U3969 (N_3969,N_1653,N_1567);
and U3970 (N_3970,N_1779,N_700);
and U3971 (N_3971,N_582,N_50);
or U3972 (N_3972,N_1504,N_538);
nor U3973 (N_3973,N_2306,N_1394);
nand U3974 (N_3974,N_37,N_2025);
nor U3975 (N_3975,N_173,N_516);
nand U3976 (N_3976,N_2343,N_2105);
nor U3977 (N_3977,N_2266,N_2405);
nor U3978 (N_3978,N_1693,N_1975);
and U3979 (N_3979,N_622,N_819);
nor U3980 (N_3980,N_1705,N_1376);
nand U3981 (N_3981,N_1429,N_2013);
and U3982 (N_3982,N_281,N_487);
nor U3983 (N_3983,N_2205,N_1308);
nand U3984 (N_3984,N_1492,N_919);
nand U3985 (N_3985,N_2027,N_1033);
nand U3986 (N_3986,N_407,N_589);
nor U3987 (N_3987,N_2254,N_2279);
and U3988 (N_3988,N_380,N_1516);
xor U3989 (N_3989,N_2275,N_553);
nor U3990 (N_3990,N_480,N_2251);
nor U3991 (N_3991,N_100,N_1688);
xnor U3992 (N_3992,N_2327,N_1950);
xor U3993 (N_3993,N_1306,N_621);
nor U3994 (N_3994,N_2374,N_1163);
and U3995 (N_3995,N_1159,N_323);
nor U3996 (N_3996,N_454,N_600);
xor U3997 (N_3997,N_1457,N_1506);
and U3998 (N_3998,N_313,N_684);
xnor U3999 (N_3999,N_2337,N_2000);
nand U4000 (N_4000,N_1790,N_565);
xnor U4001 (N_4001,N_1972,N_638);
xor U4002 (N_4002,N_1195,N_814);
or U4003 (N_4003,N_405,N_1281);
nand U4004 (N_4004,N_1077,N_1706);
xor U4005 (N_4005,N_2367,N_435);
and U4006 (N_4006,N_558,N_1690);
nor U4007 (N_4007,N_2452,N_147);
nor U4008 (N_4008,N_2162,N_743);
or U4009 (N_4009,N_1071,N_2266);
and U4010 (N_4010,N_113,N_1827);
and U4011 (N_4011,N_1165,N_330);
nor U4012 (N_4012,N_2071,N_1585);
nand U4013 (N_4013,N_903,N_2122);
nor U4014 (N_4014,N_1646,N_1581);
or U4015 (N_4015,N_1326,N_627);
and U4016 (N_4016,N_1537,N_639);
or U4017 (N_4017,N_1852,N_1144);
or U4018 (N_4018,N_244,N_195);
nand U4019 (N_4019,N_1839,N_1522);
nand U4020 (N_4020,N_1100,N_1152);
nand U4021 (N_4021,N_282,N_444);
nand U4022 (N_4022,N_2199,N_803);
nand U4023 (N_4023,N_1032,N_244);
xor U4024 (N_4024,N_1983,N_1589);
nand U4025 (N_4025,N_1326,N_2133);
and U4026 (N_4026,N_832,N_2088);
xnor U4027 (N_4027,N_2305,N_2061);
nor U4028 (N_4028,N_1581,N_1380);
xnor U4029 (N_4029,N_2126,N_1866);
nand U4030 (N_4030,N_217,N_2027);
nor U4031 (N_4031,N_1107,N_2198);
xor U4032 (N_4032,N_366,N_1901);
nand U4033 (N_4033,N_2188,N_1369);
or U4034 (N_4034,N_2059,N_1138);
nand U4035 (N_4035,N_1424,N_1458);
or U4036 (N_4036,N_1401,N_973);
nand U4037 (N_4037,N_1022,N_2360);
nand U4038 (N_4038,N_195,N_932);
or U4039 (N_4039,N_1610,N_561);
nand U4040 (N_4040,N_1672,N_1749);
nor U4041 (N_4041,N_426,N_162);
nor U4042 (N_4042,N_2476,N_2128);
nor U4043 (N_4043,N_1255,N_1032);
xor U4044 (N_4044,N_861,N_1802);
nand U4045 (N_4045,N_2147,N_939);
and U4046 (N_4046,N_2152,N_1053);
or U4047 (N_4047,N_215,N_1182);
or U4048 (N_4048,N_1958,N_2255);
nand U4049 (N_4049,N_739,N_851);
xor U4050 (N_4050,N_1429,N_1560);
or U4051 (N_4051,N_809,N_1862);
and U4052 (N_4052,N_2499,N_1990);
or U4053 (N_4053,N_1064,N_300);
nand U4054 (N_4054,N_506,N_313);
or U4055 (N_4055,N_1961,N_73);
nand U4056 (N_4056,N_1877,N_1459);
and U4057 (N_4057,N_916,N_1377);
or U4058 (N_4058,N_1037,N_2426);
xor U4059 (N_4059,N_336,N_2357);
nand U4060 (N_4060,N_1010,N_578);
and U4061 (N_4061,N_1653,N_540);
nor U4062 (N_4062,N_931,N_1068);
nor U4063 (N_4063,N_1631,N_1278);
nor U4064 (N_4064,N_1854,N_1331);
or U4065 (N_4065,N_2482,N_1930);
or U4066 (N_4066,N_1416,N_800);
nand U4067 (N_4067,N_742,N_1813);
and U4068 (N_4068,N_104,N_875);
nand U4069 (N_4069,N_2479,N_2027);
and U4070 (N_4070,N_1026,N_2243);
nor U4071 (N_4071,N_655,N_1103);
and U4072 (N_4072,N_1620,N_395);
and U4073 (N_4073,N_335,N_1031);
or U4074 (N_4074,N_747,N_1949);
xor U4075 (N_4075,N_1777,N_37);
xor U4076 (N_4076,N_1820,N_178);
and U4077 (N_4077,N_77,N_2038);
xor U4078 (N_4078,N_900,N_522);
nor U4079 (N_4079,N_749,N_883);
and U4080 (N_4080,N_1399,N_581);
and U4081 (N_4081,N_1896,N_2169);
or U4082 (N_4082,N_106,N_2017);
and U4083 (N_4083,N_2041,N_1667);
nor U4084 (N_4084,N_813,N_2407);
nand U4085 (N_4085,N_260,N_23);
and U4086 (N_4086,N_2017,N_1628);
and U4087 (N_4087,N_170,N_2389);
or U4088 (N_4088,N_98,N_2339);
nor U4089 (N_4089,N_643,N_35);
and U4090 (N_4090,N_606,N_756);
and U4091 (N_4091,N_2235,N_299);
and U4092 (N_4092,N_1753,N_922);
nand U4093 (N_4093,N_1960,N_649);
nand U4094 (N_4094,N_1029,N_2046);
or U4095 (N_4095,N_2447,N_485);
or U4096 (N_4096,N_321,N_280);
nor U4097 (N_4097,N_1165,N_775);
nor U4098 (N_4098,N_1679,N_84);
or U4099 (N_4099,N_2172,N_1364);
or U4100 (N_4100,N_145,N_1141);
nand U4101 (N_4101,N_2170,N_598);
and U4102 (N_4102,N_1948,N_240);
or U4103 (N_4103,N_1305,N_410);
and U4104 (N_4104,N_582,N_990);
nor U4105 (N_4105,N_8,N_1911);
or U4106 (N_4106,N_1350,N_2327);
nor U4107 (N_4107,N_2076,N_1139);
nand U4108 (N_4108,N_13,N_960);
or U4109 (N_4109,N_1346,N_2204);
nand U4110 (N_4110,N_1744,N_8);
or U4111 (N_4111,N_1277,N_658);
xnor U4112 (N_4112,N_1891,N_403);
or U4113 (N_4113,N_29,N_1289);
and U4114 (N_4114,N_2053,N_358);
nand U4115 (N_4115,N_579,N_95);
nand U4116 (N_4116,N_909,N_1515);
xor U4117 (N_4117,N_301,N_589);
nor U4118 (N_4118,N_1823,N_735);
and U4119 (N_4119,N_2247,N_2435);
and U4120 (N_4120,N_382,N_318);
xnor U4121 (N_4121,N_1856,N_331);
and U4122 (N_4122,N_1287,N_562);
nor U4123 (N_4123,N_1352,N_700);
nand U4124 (N_4124,N_1901,N_1124);
and U4125 (N_4125,N_138,N_921);
and U4126 (N_4126,N_918,N_980);
xor U4127 (N_4127,N_2046,N_1245);
or U4128 (N_4128,N_1565,N_1983);
and U4129 (N_4129,N_961,N_991);
nand U4130 (N_4130,N_1513,N_1854);
or U4131 (N_4131,N_1380,N_300);
and U4132 (N_4132,N_608,N_538);
or U4133 (N_4133,N_1235,N_1205);
nor U4134 (N_4134,N_471,N_1019);
nor U4135 (N_4135,N_721,N_1744);
and U4136 (N_4136,N_1236,N_1577);
and U4137 (N_4137,N_1521,N_2089);
nor U4138 (N_4138,N_945,N_274);
and U4139 (N_4139,N_408,N_2011);
nand U4140 (N_4140,N_2139,N_1149);
and U4141 (N_4141,N_2460,N_1226);
or U4142 (N_4142,N_2488,N_857);
xor U4143 (N_4143,N_933,N_1730);
nor U4144 (N_4144,N_100,N_578);
nand U4145 (N_4145,N_1417,N_1685);
nand U4146 (N_4146,N_2035,N_1481);
or U4147 (N_4147,N_1935,N_572);
nand U4148 (N_4148,N_1236,N_1420);
xor U4149 (N_4149,N_476,N_2127);
or U4150 (N_4150,N_527,N_691);
xor U4151 (N_4151,N_942,N_983);
xnor U4152 (N_4152,N_358,N_2228);
and U4153 (N_4153,N_2218,N_1266);
or U4154 (N_4154,N_968,N_95);
or U4155 (N_4155,N_588,N_1494);
and U4156 (N_4156,N_7,N_1828);
or U4157 (N_4157,N_1264,N_1627);
or U4158 (N_4158,N_471,N_893);
nand U4159 (N_4159,N_35,N_1287);
nor U4160 (N_4160,N_503,N_1126);
xnor U4161 (N_4161,N_372,N_1273);
or U4162 (N_4162,N_2096,N_189);
xor U4163 (N_4163,N_1268,N_1919);
nand U4164 (N_4164,N_1777,N_706);
and U4165 (N_4165,N_1982,N_1310);
nand U4166 (N_4166,N_1273,N_769);
nand U4167 (N_4167,N_2304,N_2325);
nand U4168 (N_4168,N_1119,N_718);
and U4169 (N_4169,N_2437,N_422);
nor U4170 (N_4170,N_1480,N_1011);
nor U4171 (N_4171,N_523,N_911);
nor U4172 (N_4172,N_2319,N_1832);
and U4173 (N_4173,N_1252,N_177);
or U4174 (N_4174,N_1350,N_1948);
nand U4175 (N_4175,N_1140,N_1158);
nor U4176 (N_4176,N_397,N_1225);
or U4177 (N_4177,N_1860,N_1718);
xor U4178 (N_4178,N_1526,N_2254);
and U4179 (N_4179,N_1106,N_1744);
and U4180 (N_4180,N_602,N_1991);
nor U4181 (N_4181,N_787,N_1136);
and U4182 (N_4182,N_1717,N_1220);
or U4183 (N_4183,N_2246,N_1243);
or U4184 (N_4184,N_2483,N_148);
nand U4185 (N_4185,N_1118,N_541);
or U4186 (N_4186,N_1861,N_1264);
xor U4187 (N_4187,N_851,N_1981);
or U4188 (N_4188,N_1397,N_741);
nand U4189 (N_4189,N_939,N_2471);
xor U4190 (N_4190,N_2262,N_1076);
nand U4191 (N_4191,N_2451,N_955);
or U4192 (N_4192,N_1285,N_392);
and U4193 (N_4193,N_1056,N_1586);
or U4194 (N_4194,N_356,N_1857);
nand U4195 (N_4195,N_1521,N_137);
nor U4196 (N_4196,N_884,N_1654);
nor U4197 (N_4197,N_2391,N_567);
nor U4198 (N_4198,N_1697,N_1706);
or U4199 (N_4199,N_1903,N_1555);
nor U4200 (N_4200,N_95,N_1086);
nand U4201 (N_4201,N_1778,N_1121);
and U4202 (N_4202,N_1924,N_1658);
nand U4203 (N_4203,N_505,N_0);
and U4204 (N_4204,N_1310,N_23);
or U4205 (N_4205,N_162,N_1417);
or U4206 (N_4206,N_365,N_686);
or U4207 (N_4207,N_1142,N_2071);
nand U4208 (N_4208,N_175,N_404);
xor U4209 (N_4209,N_1148,N_357);
nor U4210 (N_4210,N_854,N_1661);
or U4211 (N_4211,N_252,N_1529);
nand U4212 (N_4212,N_1901,N_1631);
nor U4213 (N_4213,N_49,N_1944);
and U4214 (N_4214,N_1894,N_2452);
nand U4215 (N_4215,N_835,N_726);
nand U4216 (N_4216,N_761,N_2142);
nor U4217 (N_4217,N_1184,N_1560);
or U4218 (N_4218,N_591,N_2246);
xnor U4219 (N_4219,N_473,N_1103);
nor U4220 (N_4220,N_859,N_727);
and U4221 (N_4221,N_2479,N_1468);
nand U4222 (N_4222,N_1935,N_2312);
nor U4223 (N_4223,N_1634,N_1782);
nor U4224 (N_4224,N_622,N_2020);
or U4225 (N_4225,N_922,N_1122);
xnor U4226 (N_4226,N_390,N_699);
and U4227 (N_4227,N_2357,N_1951);
nand U4228 (N_4228,N_450,N_1070);
or U4229 (N_4229,N_38,N_928);
nor U4230 (N_4230,N_1852,N_1524);
nor U4231 (N_4231,N_1735,N_1583);
nand U4232 (N_4232,N_941,N_1713);
and U4233 (N_4233,N_342,N_874);
nor U4234 (N_4234,N_2437,N_1658);
nand U4235 (N_4235,N_2163,N_2094);
nand U4236 (N_4236,N_2412,N_578);
nor U4237 (N_4237,N_741,N_1295);
nor U4238 (N_4238,N_1820,N_2040);
xnor U4239 (N_4239,N_2450,N_122);
or U4240 (N_4240,N_1123,N_788);
and U4241 (N_4241,N_35,N_1398);
nand U4242 (N_4242,N_2404,N_1406);
or U4243 (N_4243,N_328,N_2320);
or U4244 (N_4244,N_378,N_1781);
and U4245 (N_4245,N_1827,N_1705);
or U4246 (N_4246,N_1490,N_812);
xnor U4247 (N_4247,N_651,N_1183);
nand U4248 (N_4248,N_1522,N_2308);
nand U4249 (N_4249,N_599,N_1320);
nor U4250 (N_4250,N_469,N_166);
and U4251 (N_4251,N_2008,N_82);
xor U4252 (N_4252,N_2387,N_1133);
nor U4253 (N_4253,N_989,N_2486);
xnor U4254 (N_4254,N_2009,N_912);
nand U4255 (N_4255,N_1623,N_742);
or U4256 (N_4256,N_982,N_1460);
xnor U4257 (N_4257,N_2091,N_1649);
and U4258 (N_4258,N_780,N_1291);
xor U4259 (N_4259,N_2106,N_1576);
nand U4260 (N_4260,N_568,N_742);
or U4261 (N_4261,N_2483,N_2279);
or U4262 (N_4262,N_1708,N_1154);
and U4263 (N_4263,N_599,N_1035);
nand U4264 (N_4264,N_2110,N_1074);
and U4265 (N_4265,N_1885,N_2203);
or U4266 (N_4266,N_60,N_1436);
xnor U4267 (N_4267,N_521,N_1393);
and U4268 (N_4268,N_1847,N_750);
or U4269 (N_4269,N_1876,N_62);
nor U4270 (N_4270,N_1109,N_2378);
or U4271 (N_4271,N_1726,N_1241);
nor U4272 (N_4272,N_1210,N_1481);
xnor U4273 (N_4273,N_62,N_668);
nor U4274 (N_4274,N_1116,N_1414);
and U4275 (N_4275,N_2492,N_1456);
nand U4276 (N_4276,N_2333,N_1983);
xor U4277 (N_4277,N_976,N_2041);
and U4278 (N_4278,N_266,N_217);
xor U4279 (N_4279,N_408,N_333);
nor U4280 (N_4280,N_1083,N_2494);
or U4281 (N_4281,N_2177,N_2292);
or U4282 (N_4282,N_2247,N_305);
and U4283 (N_4283,N_215,N_1286);
xor U4284 (N_4284,N_438,N_949);
and U4285 (N_4285,N_1543,N_1309);
nand U4286 (N_4286,N_1477,N_2164);
xnor U4287 (N_4287,N_635,N_1024);
nand U4288 (N_4288,N_344,N_292);
nand U4289 (N_4289,N_989,N_637);
or U4290 (N_4290,N_819,N_1167);
nand U4291 (N_4291,N_526,N_1324);
and U4292 (N_4292,N_270,N_573);
nor U4293 (N_4293,N_1671,N_2008);
and U4294 (N_4294,N_1196,N_435);
nor U4295 (N_4295,N_2104,N_2127);
and U4296 (N_4296,N_978,N_1124);
nor U4297 (N_4297,N_125,N_821);
nand U4298 (N_4298,N_1847,N_142);
and U4299 (N_4299,N_259,N_1637);
nor U4300 (N_4300,N_894,N_1070);
nand U4301 (N_4301,N_1440,N_73);
or U4302 (N_4302,N_413,N_1089);
and U4303 (N_4303,N_944,N_1883);
or U4304 (N_4304,N_1685,N_1318);
and U4305 (N_4305,N_2244,N_1149);
nand U4306 (N_4306,N_2088,N_998);
xnor U4307 (N_4307,N_467,N_2102);
or U4308 (N_4308,N_136,N_1873);
or U4309 (N_4309,N_2234,N_13);
nor U4310 (N_4310,N_128,N_735);
nor U4311 (N_4311,N_2438,N_2032);
nor U4312 (N_4312,N_814,N_1598);
and U4313 (N_4313,N_1012,N_151);
or U4314 (N_4314,N_1159,N_2377);
nor U4315 (N_4315,N_2278,N_1328);
nand U4316 (N_4316,N_1957,N_914);
and U4317 (N_4317,N_1328,N_944);
nand U4318 (N_4318,N_1268,N_922);
and U4319 (N_4319,N_2023,N_2411);
nor U4320 (N_4320,N_2188,N_911);
nand U4321 (N_4321,N_1506,N_62);
nand U4322 (N_4322,N_1849,N_1935);
and U4323 (N_4323,N_1499,N_1272);
and U4324 (N_4324,N_506,N_2285);
or U4325 (N_4325,N_1596,N_1334);
or U4326 (N_4326,N_1906,N_290);
nor U4327 (N_4327,N_87,N_446);
and U4328 (N_4328,N_103,N_1787);
nor U4329 (N_4329,N_2476,N_1322);
or U4330 (N_4330,N_2257,N_369);
nor U4331 (N_4331,N_1003,N_1646);
xnor U4332 (N_4332,N_313,N_2386);
or U4333 (N_4333,N_1900,N_1571);
nand U4334 (N_4334,N_1144,N_2197);
nand U4335 (N_4335,N_981,N_1345);
nor U4336 (N_4336,N_2013,N_1973);
nand U4337 (N_4337,N_138,N_2142);
nor U4338 (N_4338,N_940,N_1532);
nor U4339 (N_4339,N_2434,N_611);
and U4340 (N_4340,N_2403,N_884);
or U4341 (N_4341,N_1706,N_564);
or U4342 (N_4342,N_2385,N_846);
nor U4343 (N_4343,N_1891,N_1122);
nor U4344 (N_4344,N_717,N_2093);
xnor U4345 (N_4345,N_999,N_1765);
or U4346 (N_4346,N_869,N_701);
nand U4347 (N_4347,N_1425,N_292);
or U4348 (N_4348,N_2016,N_255);
nor U4349 (N_4349,N_2465,N_2075);
and U4350 (N_4350,N_1922,N_301);
nand U4351 (N_4351,N_768,N_1507);
nand U4352 (N_4352,N_416,N_1318);
nand U4353 (N_4353,N_2128,N_244);
or U4354 (N_4354,N_963,N_1245);
nor U4355 (N_4355,N_721,N_1199);
nand U4356 (N_4356,N_1180,N_2465);
or U4357 (N_4357,N_1955,N_1754);
nor U4358 (N_4358,N_347,N_352);
or U4359 (N_4359,N_462,N_30);
and U4360 (N_4360,N_407,N_2408);
or U4361 (N_4361,N_135,N_1588);
nor U4362 (N_4362,N_774,N_2222);
or U4363 (N_4363,N_1524,N_550);
xor U4364 (N_4364,N_1774,N_498);
and U4365 (N_4365,N_2477,N_16);
xor U4366 (N_4366,N_277,N_2295);
or U4367 (N_4367,N_1461,N_1681);
or U4368 (N_4368,N_1066,N_2198);
or U4369 (N_4369,N_957,N_318);
nor U4370 (N_4370,N_2176,N_490);
and U4371 (N_4371,N_2070,N_186);
nand U4372 (N_4372,N_1550,N_563);
nor U4373 (N_4373,N_1009,N_1365);
and U4374 (N_4374,N_824,N_1813);
xnor U4375 (N_4375,N_1665,N_109);
nand U4376 (N_4376,N_1207,N_593);
or U4377 (N_4377,N_1473,N_2170);
nand U4378 (N_4378,N_1019,N_2416);
nand U4379 (N_4379,N_202,N_673);
xor U4380 (N_4380,N_2230,N_2275);
nor U4381 (N_4381,N_855,N_1499);
nor U4382 (N_4382,N_171,N_2447);
nand U4383 (N_4383,N_1768,N_1413);
nor U4384 (N_4384,N_1245,N_2240);
and U4385 (N_4385,N_1966,N_1639);
or U4386 (N_4386,N_735,N_1549);
nor U4387 (N_4387,N_946,N_2056);
xor U4388 (N_4388,N_677,N_942);
nand U4389 (N_4389,N_1759,N_1559);
nor U4390 (N_4390,N_1681,N_2436);
or U4391 (N_4391,N_1126,N_853);
and U4392 (N_4392,N_1695,N_1408);
nor U4393 (N_4393,N_741,N_2122);
or U4394 (N_4394,N_2046,N_697);
and U4395 (N_4395,N_1110,N_1174);
or U4396 (N_4396,N_274,N_1859);
nor U4397 (N_4397,N_1039,N_1891);
nor U4398 (N_4398,N_1881,N_1228);
nand U4399 (N_4399,N_1655,N_2254);
nand U4400 (N_4400,N_1188,N_2222);
nor U4401 (N_4401,N_563,N_853);
nand U4402 (N_4402,N_572,N_1175);
and U4403 (N_4403,N_1449,N_2212);
nor U4404 (N_4404,N_2274,N_1479);
or U4405 (N_4405,N_1350,N_205);
nor U4406 (N_4406,N_2159,N_1687);
xnor U4407 (N_4407,N_647,N_173);
and U4408 (N_4408,N_1994,N_1688);
nand U4409 (N_4409,N_2262,N_2134);
xor U4410 (N_4410,N_1946,N_895);
or U4411 (N_4411,N_1421,N_1781);
or U4412 (N_4412,N_1563,N_985);
nand U4413 (N_4413,N_971,N_2459);
nor U4414 (N_4414,N_38,N_199);
nand U4415 (N_4415,N_1561,N_51);
and U4416 (N_4416,N_273,N_1206);
and U4417 (N_4417,N_521,N_1169);
and U4418 (N_4418,N_1802,N_2276);
nor U4419 (N_4419,N_1947,N_1571);
nand U4420 (N_4420,N_303,N_1918);
nand U4421 (N_4421,N_2325,N_1699);
or U4422 (N_4422,N_500,N_974);
or U4423 (N_4423,N_2048,N_1152);
nand U4424 (N_4424,N_1211,N_1561);
nand U4425 (N_4425,N_722,N_2226);
or U4426 (N_4426,N_2095,N_1981);
or U4427 (N_4427,N_2445,N_920);
or U4428 (N_4428,N_1415,N_2490);
and U4429 (N_4429,N_103,N_1162);
or U4430 (N_4430,N_151,N_2132);
nor U4431 (N_4431,N_242,N_1236);
or U4432 (N_4432,N_314,N_2138);
or U4433 (N_4433,N_2074,N_1478);
nand U4434 (N_4434,N_535,N_1417);
nand U4435 (N_4435,N_1901,N_2037);
nor U4436 (N_4436,N_1338,N_315);
nor U4437 (N_4437,N_2192,N_1262);
nand U4438 (N_4438,N_692,N_1672);
xnor U4439 (N_4439,N_1442,N_1778);
nand U4440 (N_4440,N_1906,N_483);
or U4441 (N_4441,N_1018,N_1724);
nor U4442 (N_4442,N_2413,N_885);
and U4443 (N_4443,N_1861,N_1963);
and U4444 (N_4444,N_1526,N_2167);
nand U4445 (N_4445,N_1515,N_1732);
xnor U4446 (N_4446,N_1025,N_2194);
or U4447 (N_4447,N_1030,N_1593);
or U4448 (N_4448,N_2344,N_1824);
nand U4449 (N_4449,N_2306,N_38);
and U4450 (N_4450,N_1551,N_1858);
and U4451 (N_4451,N_144,N_507);
nor U4452 (N_4452,N_34,N_1368);
nand U4453 (N_4453,N_522,N_977);
nand U4454 (N_4454,N_1476,N_2444);
nor U4455 (N_4455,N_926,N_758);
nand U4456 (N_4456,N_1229,N_227);
or U4457 (N_4457,N_179,N_715);
nand U4458 (N_4458,N_2208,N_670);
or U4459 (N_4459,N_973,N_1030);
or U4460 (N_4460,N_627,N_2237);
or U4461 (N_4461,N_2043,N_398);
or U4462 (N_4462,N_187,N_2297);
nor U4463 (N_4463,N_1504,N_467);
or U4464 (N_4464,N_1800,N_2180);
or U4465 (N_4465,N_1437,N_1620);
xor U4466 (N_4466,N_1609,N_2444);
nand U4467 (N_4467,N_995,N_2059);
xor U4468 (N_4468,N_546,N_768);
and U4469 (N_4469,N_56,N_1544);
nor U4470 (N_4470,N_1191,N_1004);
nand U4471 (N_4471,N_1726,N_2223);
or U4472 (N_4472,N_1988,N_940);
nand U4473 (N_4473,N_1427,N_133);
and U4474 (N_4474,N_17,N_2444);
and U4475 (N_4475,N_1708,N_972);
and U4476 (N_4476,N_2278,N_880);
and U4477 (N_4477,N_1572,N_1122);
or U4478 (N_4478,N_65,N_354);
nand U4479 (N_4479,N_33,N_1544);
nand U4480 (N_4480,N_716,N_681);
xor U4481 (N_4481,N_116,N_2263);
and U4482 (N_4482,N_797,N_903);
nor U4483 (N_4483,N_1403,N_1529);
or U4484 (N_4484,N_580,N_1921);
or U4485 (N_4485,N_1642,N_1238);
nor U4486 (N_4486,N_186,N_808);
or U4487 (N_4487,N_924,N_2390);
and U4488 (N_4488,N_2150,N_2109);
xor U4489 (N_4489,N_1231,N_1627);
and U4490 (N_4490,N_379,N_941);
nor U4491 (N_4491,N_599,N_116);
nand U4492 (N_4492,N_2493,N_2257);
nor U4493 (N_4493,N_1125,N_1190);
nor U4494 (N_4494,N_71,N_541);
or U4495 (N_4495,N_2457,N_2459);
or U4496 (N_4496,N_558,N_636);
xor U4497 (N_4497,N_1714,N_626);
or U4498 (N_4498,N_1051,N_157);
and U4499 (N_4499,N_2413,N_2265);
nand U4500 (N_4500,N_2263,N_752);
and U4501 (N_4501,N_881,N_2471);
or U4502 (N_4502,N_1493,N_245);
and U4503 (N_4503,N_1334,N_2429);
and U4504 (N_4504,N_1766,N_105);
and U4505 (N_4505,N_1067,N_2187);
or U4506 (N_4506,N_941,N_1785);
or U4507 (N_4507,N_801,N_57);
or U4508 (N_4508,N_2221,N_1177);
nand U4509 (N_4509,N_2129,N_1317);
or U4510 (N_4510,N_2136,N_2130);
nor U4511 (N_4511,N_911,N_2290);
and U4512 (N_4512,N_2337,N_2418);
and U4513 (N_4513,N_293,N_957);
nand U4514 (N_4514,N_708,N_1269);
nand U4515 (N_4515,N_263,N_33);
nor U4516 (N_4516,N_166,N_153);
nor U4517 (N_4517,N_104,N_1086);
nand U4518 (N_4518,N_1020,N_2086);
xor U4519 (N_4519,N_619,N_1084);
and U4520 (N_4520,N_1237,N_498);
nand U4521 (N_4521,N_289,N_185);
and U4522 (N_4522,N_122,N_1130);
nor U4523 (N_4523,N_1119,N_1554);
nor U4524 (N_4524,N_142,N_839);
and U4525 (N_4525,N_1931,N_1422);
or U4526 (N_4526,N_718,N_238);
xor U4527 (N_4527,N_1132,N_1586);
or U4528 (N_4528,N_1936,N_2225);
or U4529 (N_4529,N_575,N_2150);
nand U4530 (N_4530,N_660,N_414);
nor U4531 (N_4531,N_1038,N_1429);
nor U4532 (N_4532,N_450,N_1821);
nand U4533 (N_4533,N_1351,N_431);
and U4534 (N_4534,N_171,N_2061);
nand U4535 (N_4535,N_589,N_366);
nor U4536 (N_4536,N_1247,N_1964);
or U4537 (N_4537,N_890,N_922);
nor U4538 (N_4538,N_2069,N_333);
or U4539 (N_4539,N_1965,N_2229);
nand U4540 (N_4540,N_1729,N_410);
nand U4541 (N_4541,N_2311,N_748);
nor U4542 (N_4542,N_1104,N_1225);
or U4543 (N_4543,N_2478,N_885);
and U4544 (N_4544,N_577,N_1297);
or U4545 (N_4545,N_2350,N_2051);
nand U4546 (N_4546,N_27,N_307);
and U4547 (N_4547,N_190,N_2410);
or U4548 (N_4548,N_2011,N_1799);
or U4549 (N_4549,N_926,N_1359);
or U4550 (N_4550,N_287,N_100);
nor U4551 (N_4551,N_175,N_1682);
and U4552 (N_4552,N_814,N_577);
and U4553 (N_4553,N_1558,N_2265);
or U4554 (N_4554,N_324,N_1546);
and U4555 (N_4555,N_1443,N_733);
and U4556 (N_4556,N_1086,N_1200);
nand U4557 (N_4557,N_94,N_370);
xnor U4558 (N_4558,N_1616,N_1183);
nand U4559 (N_4559,N_2169,N_649);
and U4560 (N_4560,N_1058,N_311);
nand U4561 (N_4561,N_480,N_1786);
nor U4562 (N_4562,N_938,N_365);
nand U4563 (N_4563,N_720,N_2306);
or U4564 (N_4564,N_897,N_2299);
nand U4565 (N_4565,N_1848,N_2197);
and U4566 (N_4566,N_1423,N_2437);
nand U4567 (N_4567,N_466,N_1288);
xor U4568 (N_4568,N_2430,N_1894);
nand U4569 (N_4569,N_1019,N_1611);
nor U4570 (N_4570,N_1334,N_1559);
or U4571 (N_4571,N_1057,N_1066);
nor U4572 (N_4572,N_1914,N_1491);
or U4573 (N_4573,N_1844,N_1174);
nor U4574 (N_4574,N_486,N_1367);
xor U4575 (N_4575,N_1282,N_1212);
nor U4576 (N_4576,N_563,N_2368);
and U4577 (N_4577,N_1520,N_1125);
and U4578 (N_4578,N_1497,N_2067);
nor U4579 (N_4579,N_134,N_1934);
and U4580 (N_4580,N_232,N_1305);
nand U4581 (N_4581,N_1618,N_356);
and U4582 (N_4582,N_1504,N_1155);
or U4583 (N_4583,N_1642,N_561);
and U4584 (N_4584,N_196,N_2364);
nand U4585 (N_4585,N_1840,N_782);
nand U4586 (N_4586,N_2055,N_875);
nand U4587 (N_4587,N_1928,N_207);
and U4588 (N_4588,N_718,N_490);
nor U4589 (N_4589,N_454,N_2334);
nor U4590 (N_4590,N_2120,N_1374);
nand U4591 (N_4591,N_1661,N_2258);
or U4592 (N_4592,N_1206,N_211);
or U4593 (N_4593,N_8,N_2384);
nor U4594 (N_4594,N_1996,N_401);
nor U4595 (N_4595,N_1556,N_1386);
and U4596 (N_4596,N_1018,N_762);
nor U4597 (N_4597,N_1959,N_295);
xor U4598 (N_4598,N_595,N_1849);
nor U4599 (N_4599,N_2178,N_2277);
nor U4600 (N_4600,N_923,N_1182);
nor U4601 (N_4601,N_933,N_51);
nand U4602 (N_4602,N_2012,N_1616);
and U4603 (N_4603,N_2468,N_2245);
or U4604 (N_4604,N_292,N_2095);
or U4605 (N_4605,N_41,N_1492);
or U4606 (N_4606,N_1070,N_71);
or U4607 (N_4607,N_2009,N_2270);
or U4608 (N_4608,N_2358,N_689);
and U4609 (N_4609,N_421,N_165);
or U4610 (N_4610,N_1800,N_423);
or U4611 (N_4611,N_1415,N_1554);
nor U4612 (N_4612,N_267,N_407);
and U4613 (N_4613,N_2155,N_2403);
nor U4614 (N_4614,N_1114,N_261);
xnor U4615 (N_4615,N_2078,N_2337);
or U4616 (N_4616,N_191,N_2374);
nor U4617 (N_4617,N_443,N_1298);
or U4618 (N_4618,N_1311,N_444);
or U4619 (N_4619,N_1952,N_1404);
and U4620 (N_4620,N_757,N_2312);
and U4621 (N_4621,N_285,N_1285);
nand U4622 (N_4622,N_1351,N_904);
nor U4623 (N_4623,N_2374,N_2477);
xnor U4624 (N_4624,N_929,N_1517);
or U4625 (N_4625,N_2184,N_1992);
or U4626 (N_4626,N_1653,N_1272);
nor U4627 (N_4627,N_285,N_2289);
or U4628 (N_4628,N_435,N_1019);
and U4629 (N_4629,N_116,N_702);
nor U4630 (N_4630,N_1875,N_1723);
nand U4631 (N_4631,N_2341,N_1321);
nor U4632 (N_4632,N_88,N_1664);
or U4633 (N_4633,N_981,N_487);
nor U4634 (N_4634,N_2114,N_719);
or U4635 (N_4635,N_1455,N_1581);
and U4636 (N_4636,N_2430,N_2118);
or U4637 (N_4637,N_1957,N_918);
nor U4638 (N_4638,N_2005,N_904);
or U4639 (N_4639,N_403,N_1901);
or U4640 (N_4640,N_1526,N_2178);
nor U4641 (N_4641,N_167,N_131);
and U4642 (N_4642,N_1927,N_558);
nand U4643 (N_4643,N_2094,N_687);
or U4644 (N_4644,N_2017,N_1701);
and U4645 (N_4645,N_2275,N_2262);
nor U4646 (N_4646,N_1125,N_1986);
or U4647 (N_4647,N_1699,N_2427);
nand U4648 (N_4648,N_779,N_726);
and U4649 (N_4649,N_147,N_2024);
or U4650 (N_4650,N_68,N_2376);
nor U4651 (N_4651,N_1124,N_1591);
and U4652 (N_4652,N_256,N_677);
nor U4653 (N_4653,N_2085,N_997);
nand U4654 (N_4654,N_446,N_2466);
xor U4655 (N_4655,N_1092,N_200);
and U4656 (N_4656,N_1751,N_2274);
and U4657 (N_4657,N_933,N_1482);
and U4658 (N_4658,N_740,N_890);
nor U4659 (N_4659,N_2218,N_2032);
or U4660 (N_4660,N_1369,N_569);
nand U4661 (N_4661,N_970,N_2383);
and U4662 (N_4662,N_286,N_298);
nand U4663 (N_4663,N_1837,N_1361);
xor U4664 (N_4664,N_2176,N_1722);
and U4665 (N_4665,N_436,N_2225);
nand U4666 (N_4666,N_1920,N_2181);
and U4667 (N_4667,N_1651,N_1636);
nand U4668 (N_4668,N_1042,N_1483);
or U4669 (N_4669,N_369,N_2455);
nand U4670 (N_4670,N_589,N_1654);
nor U4671 (N_4671,N_16,N_180);
or U4672 (N_4672,N_1771,N_2022);
nand U4673 (N_4673,N_1394,N_1823);
nor U4674 (N_4674,N_1844,N_349);
xor U4675 (N_4675,N_579,N_1041);
and U4676 (N_4676,N_1823,N_885);
nor U4677 (N_4677,N_184,N_1128);
xor U4678 (N_4678,N_1089,N_1905);
nor U4679 (N_4679,N_174,N_1096);
nand U4680 (N_4680,N_589,N_2248);
nand U4681 (N_4681,N_1389,N_990);
xor U4682 (N_4682,N_260,N_259);
nor U4683 (N_4683,N_1029,N_1921);
nor U4684 (N_4684,N_769,N_1459);
nand U4685 (N_4685,N_1755,N_772);
or U4686 (N_4686,N_2077,N_129);
or U4687 (N_4687,N_218,N_2234);
nor U4688 (N_4688,N_148,N_1661);
nand U4689 (N_4689,N_896,N_1106);
and U4690 (N_4690,N_621,N_696);
and U4691 (N_4691,N_2476,N_512);
and U4692 (N_4692,N_2163,N_1563);
nor U4693 (N_4693,N_2241,N_490);
or U4694 (N_4694,N_51,N_80);
and U4695 (N_4695,N_659,N_1565);
nand U4696 (N_4696,N_1363,N_2036);
and U4697 (N_4697,N_179,N_303);
nor U4698 (N_4698,N_683,N_2409);
and U4699 (N_4699,N_1051,N_1650);
nand U4700 (N_4700,N_759,N_2237);
or U4701 (N_4701,N_872,N_1286);
and U4702 (N_4702,N_818,N_1878);
or U4703 (N_4703,N_500,N_200);
nand U4704 (N_4704,N_2400,N_1865);
xnor U4705 (N_4705,N_568,N_1126);
nand U4706 (N_4706,N_84,N_1476);
and U4707 (N_4707,N_2481,N_1205);
and U4708 (N_4708,N_2180,N_1014);
xor U4709 (N_4709,N_1863,N_2225);
nand U4710 (N_4710,N_239,N_2233);
and U4711 (N_4711,N_2021,N_1733);
nand U4712 (N_4712,N_569,N_1529);
and U4713 (N_4713,N_1682,N_59);
nor U4714 (N_4714,N_761,N_623);
or U4715 (N_4715,N_1091,N_1705);
nor U4716 (N_4716,N_1447,N_2109);
nor U4717 (N_4717,N_300,N_1704);
or U4718 (N_4718,N_899,N_416);
xnor U4719 (N_4719,N_840,N_880);
and U4720 (N_4720,N_1593,N_531);
nor U4721 (N_4721,N_1236,N_962);
nor U4722 (N_4722,N_46,N_2485);
and U4723 (N_4723,N_426,N_2069);
and U4724 (N_4724,N_1302,N_1052);
and U4725 (N_4725,N_1693,N_2234);
xnor U4726 (N_4726,N_2209,N_1522);
nor U4727 (N_4727,N_667,N_1950);
nand U4728 (N_4728,N_493,N_1332);
or U4729 (N_4729,N_1189,N_1591);
nor U4730 (N_4730,N_220,N_1822);
nand U4731 (N_4731,N_1091,N_1071);
nor U4732 (N_4732,N_197,N_1202);
nor U4733 (N_4733,N_190,N_1400);
or U4734 (N_4734,N_2230,N_1019);
or U4735 (N_4735,N_1731,N_1126);
or U4736 (N_4736,N_555,N_423);
nor U4737 (N_4737,N_814,N_2493);
or U4738 (N_4738,N_761,N_2254);
nor U4739 (N_4739,N_1287,N_599);
or U4740 (N_4740,N_2452,N_814);
nand U4741 (N_4741,N_1434,N_1949);
xnor U4742 (N_4742,N_708,N_2015);
nor U4743 (N_4743,N_1457,N_557);
nand U4744 (N_4744,N_1693,N_1594);
or U4745 (N_4745,N_1168,N_722);
nor U4746 (N_4746,N_584,N_245);
nor U4747 (N_4747,N_497,N_1453);
nand U4748 (N_4748,N_1003,N_1799);
or U4749 (N_4749,N_1491,N_2216);
or U4750 (N_4750,N_1895,N_2284);
or U4751 (N_4751,N_293,N_1192);
and U4752 (N_4752,N_2148,N_723);
nand U4753 (N_4753,N_925,N_1392);
or U4754 (N_4754,N_1965,N_2445);
and U4755 (N_4755,N_260,N_57);
nor U4756 (N_4756,N_2295,N_2275);
or U4757 (N_4757,N_2421,N_1640);
and U4758 (N_4758,N_46,N_461);
xor U4759 (N_4759,N_1421,N_1595);
or U4760 (N_4760,N_1537,N_2244);
or U4761 (N_4761,N_97,N_1054);
nor U4762 (N_4762,N_524,N_1581);
or U4763 (N_4763,N_1744,N_1442);
nor U4764 (N_4764,N_964,N_543);
nand U4765 (N_4765,N_2179,N_263);
nor U4766 (N_4766,N_1860,N_2076);
xor U4767 (N_4767,N_1555,N_72);
nand U4768 (N_4768,N_1259,N_99);
or U4769 (N_4769,N_1294,N_217);
nand U4770 (N_4770,N_1395,N_1137);
nand U4771 (N_4771,N_1071,N_1673);
or U4772 (N_4772,N_2265,N_1286);
and U4773 (N_4773,N_326,N_1226);
nor U4774 (N_4774,N_585,N_774);
xnor U4775 (N_4775,N_660,N_75);
and U4776 (N_4776,N_1390,N_12);
nand U4777 (N_4777,N_1345,N_980);
and U4778 (N_4778,N_3,N_1073);
or U4779 (N_4779,N_35,N_1470);
and U4780 (N_4780,N_1563,N_1407);
or U4781 (N_4781,N_972,N_1298);
nor U4782 (N_4782,N_438,N_1534);
nand U4783 (N_4783,N_1264,N_870);
and U4784 (N_4784,N_1091,N_610);
or U4785 (N_4785,N_26,N_330);
nand U4786 (N_4786,N_2366,N_208);
nand U4787 (N_4787,N_2121,N_2243);
nand U4788 (N_4788,N_1616,N_895);
or U4789 (N_4789,N_1307,N_236);
and U4790 (N_4790,N_505,N_1419);
and U4791 (N_4791,N_453,N_1546);
and U4792 (N_4792,N_1789,N_2350);
nand U4793 (N_4793,N_263,N_3);
xnor U4794 (N_4794,N_1098,N_1874);
or U4795 (N_4795,N_153,N_602);
nand U4796 (N_4796,N_219,N_287);
and U4797 (N_4797,N_2127,N_1431);
nand U4798 (N_4798,N_1722,N_161);
or U4799 (N_4799,N_1497,N_988);
xor U4800 (N_4800,N_337,N_2384);
nand U4801 (N_4801,N_822,N_1753);
or U4802 (N_4802,N_996,N_866);
and U4803 (N_4803,N_1941,N_631);
or U4804 (N_4804,N_222,N_1279);
nand U4805 (N_4805,N_2071,N_1709);
or U4806 (N_4806,N_2407,N_1726);
nand U4807 (N_4807,N_505,N_565);
nor U4808 (N_4808,N_433,N_784);
and U4809 (N_4809,N_465,N_73);
nand U4810 (N_4810,N_2225,N_726);
nand U4811 (N_4811,N_2270,N_701);
or U4812 (N_4812,N_829,N_1171);
nor U4813 (N_4813,N_1642,N_1824);
nor U4814 (N_4814,N_2373,N_439);
or U4815 (N_4815,N_1205,N_927);
and U4816 (N_4816,N_31,N_556);
nor U4817 (N_4817,N_2452,N_1909);
nor U4818 (N_4818,N_2351,N_1571);
nand U4819 (N_4819,N_2438,N_561);
nand U4820 (N_4820,N_872,N_285);
or U4821 (N_4821,N_1771,N_2213);
nor U4822 (N_4822,N_1035,N_320);
and U4823 (N_4823,N_1918,N_30);
and U4824 (N_4824,N_1005,N_1680);
or U4825 (N_4825,N_969,N_1454);
or U4826 (N_4826,N_1251,N_1349);
nand U4827 (N_4827,N_1132,N_272);
nor U4828 (N_4828,N_1593,N_911);
nor U4829 (N_4829,N_679,N_942);
nor U4830 (N_4830,N_828,N_1649);
and U4831 (N_4831,N_2440,N_1924);
or U4832 (N_4832,N_472,N_574);
nand U4833 (N_4833,N_1500,N_1040);
nand U4834 (N_4834,N_779,N_2000);
or U4835 (N_4835,N_1677,N_1377);
or U4836 (N_4836,N_521,N_1071);
nor U4837 (N_4837,N_213,N_283);
nand U4838 (N_4838,N_961,N_1235);
nor U4839 (N_4839,N_1011,N_1609);
nand U4840 (N_4840,N_1192,N_2351);
nand U4841 (N_4841,N_692,N_307);
or U4842 (N_4842,N_2350,N_2423);
nor U4843 (N_4843,N_1099,N_1089);
nor U4844 (N_4844,N_1522,N_2371);
and U4845 (N_4845,N_2407,N_1814);
and U4846 (N_4846,N_595,N_1748);
nand U4847 (N_4847,N_1059,N_1214);
and U4848 (N_4848,N_992,N_1590);
xor U4849 (N_4849,N_745,N_1277);
or U4850 (N_4850,N_2357,N_1145);
or U4851 (N_4851,N_1934,N_997);
and U4852 (N_4852,N_900,N_1222);
and U4853 (N_4853,N_1557,N_1072);
nor U4854 (N_4854,N_2239,N_827);
nand U4855 (N_4855,N_2340,N_1044);
and U4856 (N_4856,N_700,N_1420);
nor U4857 (N_4857,N_1060,N_7);
nor U4858 (N_4858,N_2277,N_1286);
and U4859 (N_4859,N_160,N_1658);
nor U4860 (N_4860,N_219,N_587);
and U4861 (N_4861,N_911,N_2180);
and U4862 (N_4862,N_1243,N_1111);
or U4863 (N_4863,N_476,N_507);
and U4864 (N_4864,N_2237,N_53);
nand U4865 (N_4865,N_2018,N_53);
nand U4866 (N_4866,N_1365,N_2295);
or U4867 (N_4867,N_1367,N_1650);
nor U4868 (N_4868,N_2007,N_1187);
nand U4869 (N_4869,N_718,N_1569);
nor U4870 (N_4870,N_1212,N_983);
or U4871 (N_4871,N_1603,N_212);
or U4872 (N_4872,N_777,N_1795);
nand U4873 (N_4873,N_479,N_2377);
xnor U4874 (N_4874,N_204,N_2495);
nor U4875 (N_4875,N_170,N_2346);
nor U4876 (N_4876,N_1145,N_489);
nand U4877 (N_4877,N_1400,N_1595);
or U4878 (N_4878,N_1029,N_1584);
or U4879 (N_4879,N_350,N_2080);
xor U4880 (N_4880,N_1082,N_675);
and U4881 (N_4881,N_743,N_78);
nor U4882 (N_4882,N_533,N_1686);
nor U4883 (N_4883,N_2437,N_499);
or U4884 (N_4884,N_2342,N_1895);
xor U4885 (N_4885,N_223,N_1170);
xnor U4886 (N_4886,N_405,N_1065);
or U4887 (N_4887,N_1042,N_1994);
xor U4888 (N_4888,N_343,N_1703);
nor U4889 (N_4889,N_2469,N_1731);
and U4890 (N_4890,N_1867,N_1726);
nor U4891 (N_4891,N_121,N_1017);
nor U4892 (N_4892,N_2068,N_285);
nor U4893 (N_4893,N_701,N_1638);
xor U4894 (N_4894,N_1159,N_2285);
or U4895 (N_4895,N_1608,N_2284);
nand U4896 (N_4896,N_417,N_2337);
nand U4897 (N_4897,N_2423,N_454);
nor U4898 (N_4898,N_540,N_125);
nand U4899 (N_4899,N_231,N_697);
xnor U4900 (N_4900,N_645,N_1202);
nor U4901 (N_4901,N_2092,N_856);
nand U4902 (N_4902,N_749,N_2072);
nor U4903 (N_4903,N_2178,N_1966);
nand U4904 (N_4904,N_473,N_2293);
nor U4905 (N_4905,N_521,N_730);
and U4906 (N_4906,N_1151,N_78);
nand U4907 (N_4907,N_1642,N_1311);
or U4908 (N_4908,N_2403,N_2273);
or U4909 (N_4909,N_2,N_438);
nor U4910 (N_4910,N_162,N_2219);
nand U4911 (N_4911,N_1052,N_877);
nand U4912 (N_4912,N_152,N_362);
nand U4913 (N_4913,N_1801,N_744);
nor U4914 (N_4914,N_123,N_2407);
nor U4915 (N_4915,N_1858,N_2481);
xnor U4916 (N_4916,N_509,N_2466);
nand U4917 (N_4917,N_460,N_1524);
nand U4918 (N_4918,N_127,N_1249);
or U4919 (N_4919,N_1650,N_102);
and U4920 (N_4920,N_2242,N_1445);
and U4921 (N_4921,N_1566,N_2195);
nand U4922 (N_4922,N_1902,N_2153);
or U4923 (N_4923,N_2010,N_381);
nor U4924 (N_4924,N_273,N_708);
or U4925 (N_4925,N_2492,N_1331);
xnor U4926 (N_4926,N_1123,N_866);
and U4927 (N_4927,N_1968,N_1916);
and U4928 (N_4928,N_1073,N_1437);
or U4929 (N_4929,N_307,N_275);
nand U4930 (N_4930,N_969,N_1885);
nand U4931 (N_4931,N_331,N_412);
nor U4932 (N_4932,N_1108,N_1473);
and U4933 (N_4933,N_1538,N_237);
nor U4934 (N_4934,N_2230,N_2439);
or U4935 (N_4935,N_1752,N_23);
and U4936 (N_4936,N_575,N_663);
and U4937 (N_4937,N_63,N_2335);
xnor U4938 (N_4938,N_2321,N_1632);
and U4939 (N_4939,N_1438,N_982);
xnor U4940 (N_4940,N_973,N_2066);
and U4941 (N_4941,N_1057,N_761);
and U4942 (N_4942,N_2040,N_664);
or U4943 (N_4943,N_1240,N_2084);
nand U4944 (N_4944,N_2061,N_1767);
or U4945 (N_4945,N_184,N_867);
xor U4946 (N_4946,N_233,N_1061);
nand U4947 (N_4947,N_1515,N_1003);
nor U4948 (N_4948,N_289,N_543);
nor U4949 (N_4949,N_173,N_2477);
nor U4950 (N_4950,N_1778,N_2284);
or U4951 (N_4951,N_288,N_307);
nand U4952 (N_4952,N_2158,N_670);
or U4953 (N_4953,N_1548,N_600);
nand U4954 (N_4954,N_1533,N_2229);
or U4955 (N_4955,N_1858,N_1950);
or U4956 (N_4956,N_1350,N_2373);
xor U4957 (N_4957,N_2015,N_1701);
nand U4958 (N_4958,N_881,N_1938);
nand U4959 (N_4959,N_1519,N_2141);
or U4960 (N_4960,N_2408,N_1317);
nor U4961 (N_4961,N_2015,N_1508);
nand U4962 (N_4962,N_2317,N_1704);
or U4963 (N_4963,N_1954,N_697);
xor U4964 (N_4964,N_1080,N_444);
and U4965 (N_4965,N_2086,N_1855);
nor U4966 (N_4966,N_1464,N_1936);
or U4967 (N_4967,N_503,N_2158);
and U4968 (N_4968,N_1346,N_648);
nand U4969 (N_4969,N_1570,N_708);
and U4970 (N_4970,N_207,N_1329);
or U4971 (N_4971,N_1409,N_881);
nor U4972 (N_4972,N_2188,N_2110);
or U4973 (N_4973,N_1906,N_1662);
or U4974 (N_4974,N_391,N_2461);
nand U4975 (N_4975,N_463,N_1438);
and U4976 (N_4976,N_2182,N_115);
nor U4977 (N_4977,N_352,N_947);
and U4978 (N_4978,N_1122,N_1318);
or U4979 (N_4979,N_2230,N_67);
or U4980 (N_4980,N_1756,N_352);
nor U4981 (N_4981,N_66,N_1445);
nor U4982 (N_4982,N_221,N_1983);
or U4983 (N_4983,N_634,N_1858);
and U4984 (N_4984,N_2238,N_1356);
or U4985 (N_4985,N_1842,N_446);
and U4986 (N_4986,N_831,N_975);
nand U4987 (N_4987,N_1204,N_1541);
and U4988 (N_4988,N_626,N_318);
xor U4989 (N_4989,N_1107,N_176);
nor U4990 (N_4990,N_1635,N_2075);
nand U4991 (N_4991,N_2128,N_2051);
xnor U4992 (N_4992,N_1751,N_140);
and U4993 (N_4993,N_1322,N_1233);
and U4994 (N_4994,N_214,N_1297);
or U4995 (N_4995,N_437,N_1843);
or U4996 (N_4996,N_1480,N_1460);
or U4997 (N_4997,N_1600,N_357);
nor U4998 (N_4998,N_60,N_1794);
and U4999 (N_4999,N_1604,N_1036);
xnor U5000 (N_5000,N_3788,N_4008);
and U5001 (N_5001,N_2733,N_3344);
nand U5002 (N_5002,N_3781,N_2533);
and U5003 (N_5003,N_3698,N_4808);
nor U5004 (N_5004,N_3951,N_3246);
nor U5005 (N_5005,N_4246,N_3553);
nand U5006 (N_5006,N_4159,N_3879);
or U5007 (N_5007,N_4579,N_3319);
nor U5008 (N_5008,N_4940,N_3403);
nor U5009 (N_5009,N_4670,N_4158);
and U5010 (N_5010,N_4882,N_2896);
nor U5011 (N_5011,N_3852,N_3619);
nand U5012 (N_5012,N_3596,N_3439);
xor U5013 (N_5013,N_2655,N_3661);
nand U5014 (N_5014,N_4618,N_4464);
and U5015 (N_5015,N_4713,N_4910);
and U5016 (N_5016,N_2900,N_4253);
nor U5017 (N_5017,N_2717,N_3093);
xnor U5018 (N_5018,N_4161,N_3881);
or U5019 (N_5019,N_2992,N_2786);
nor U5020 (N_5020,N_3701,N_3212);
nand U5021 (N_5021,N_3767,N_3373);
or U5022 (N_5022,N_4728,N_4594);
nand U5023 (N_5023,N_3548,N_2707);
nand U5024 (N_5024,N_2701,N_2735);
nor U5025 (N_5025,N_4827,N_3886);
and U5026 (N_5026,N_2930,N_3032);
nand U5027 (N_5027,N_4771,N_2544);
nor U5028 (N_5028,N_2874,N_2702);
nand U5029 (N_5029,N_3709,N_2609);
and U5030 (N_5030,N_3053,N_4915);
and U5031 (N_5031,N_3140,N_4991);
nand U5032 (N_5032,N_2644,N_3685);
nand U5033 (N_5033,N_4147,N_4197);
nand U5034 (N_5034,N_4118,N_2798);
or U5035 (N_5035,N_2954,N_3324);
or U5036 (N_5036,N_2864,N_4558);
nand U5037 (N_5037,N_4261,N_2673);
and U5038 (N_5038,N_3106,N_2570);
or U5039 (N_5039,N_3449,N_2723);
and U5040 (N_5040,N_3916,N_3102);
and U5041 (N_5041,N_3637,N_3014);
or U5042 (N_5042,N_3476,N_4078);
nor U5043 (N_5043,N_2618,N_2805);
and U5044 (N_5044,N_2780,N_3578);
or U5045 (N_5045,N_4825,N_4793);
or U5046 (N_5046,N_3110,N_4073);
and U5047 (N_5047,N_3227,N_3390);
nand U5048 (N_5048,N_3871,N_3037);
or U5049 (N_5049,N_3622,N_3535);
and U5050 (N_5050,N_2984,N_4730);
and U5051 (N_5051,N_4964,N_4623);
xnor U5052 (N_5052,N_2546,N_4205);
nor U5053 (N_5053,N_3529,N_4887);
and U5054 (N_5054,N_3338,N_3672);
and U5055 (N_5055,N_4692,N_4050);
or U5056 (N_5056,N_2695,N_4584);
nand U5057 (N_5057,N_4251,N_4903);
nor U5058 (N_5058,N_3104,N_4489);
nand U5059 (N_5059,N_3311,N_3552);
and U5060 (N_5060,N_2776,N_2699);
nand U5061 (N_5061,N_2950,N_3854);
nand U5062 (N_5062,N_4537,N_3010);
and U5063 (N_5063,N_3209,N_3714);
xnor U5064 (N_5064,N_4933,N_4060);
or U5065 (N_5065,N_2710,N_2636);
nand U5066 (N_5066,N_3623,N_2678);
and U5067 (N_5067,N_2576,N_3550);
nor U5068 (N_5068,N_2648,N_3090);
xor U5069 (N_5069,N_4637,N_4459);
or U5070 (N_5070,N_4313,N_4001);
nand U5071 (N_5071,N_3254,N_3676);
nand U5072 (N_5072,N_4708,N_3420);
xor U5073 (N_5073,N_4206,N_3967);
or U5074 (N_5074,N_4444,N_3187);
nor U5075 (N_5075,N_2854,N_3423);
and U5076 (N_5076,N_3411,N_3241);
nor U5077 (N_5077,N_3895,N_4066);
nor U5078 (N_5078,N_4653,N_3494);
or U5079 (N_5079,N_4519,N_4006);
nor U5080 (N_5080,N_2846,N_3720);
and U5081 (N_5081,N_4768,N_2907);
nor U5082 (N_5082,N_3351,N_4611);
or U5083 (N_5083,N_3989,N_2745);
nand U5084 (N_5084,N_2899,N_3841);
or U5085 (N_5085,N_4819,N_4898);
nand U5086 (N_5086,N_2602,N_4457);
xor U5087 (N_5087,N_3480,N_3786);
or U5088 (N_5088,N_2993,N_4113);
or U5089 (N_5089,N_2961,N_4757);
nor U5090 (N_5090,N_3772,N_4862);
nand U5091 (N_5091,N_3092,N_3581);
nand U5092 (N_5092,N_4559,N_3129);
nand U5093 (N_5093,N_4121,N_2782);
or U5094 (N_5094,N_2860,N_3611);
or U5095 (N_5095,N_3865,N_4296);
xnor U5096 (N_5096,N_3127,N_4650);
nand U5097 (N_5097,N_3911,N_3229);
and U5098 (N_5098,N_3280,N_2525);
and U5099 (N_5099,N_3418,N_3337);
and U5100 (N_5100,N_3148,N_2698);
nand U5101 (N_5101,N_2785,N_3600);
or U5102 (N_5102,N_2720,N_2687);
nor U5103 (N_5103,N_4271,N_4076);
or U5104 (N_5104,N_4082,N_3632);
nand U5105 (N_5105,N_4520,N_2944);
or U5106 (N_5106,N_3931,N_2939);
and U5107 (N_5107,N_2728,N_3851);
and U5108 (N_5108,N_4247,N_4353);
nor U5109 (N_5109,N_4326,N_4487);
nor U5110 (N_5110,N_3308,N_2621);
nor U5111 (N_5111,N_3584,N_3188);
or U5112 (N_5112,N_4681,N_2787);
nor U5113 (N_5113,N_3215,N_4171);
and U5114 (N_5114,N_3897,N_4644);
nand U5115 (N_5115,N_3486,N_3519);
nor U5116 (N_5116,N_3583,N_3828);
nor U5117 (N_5117,N_2884,N_4508);
and U5118 (N_5118,N_4621,N_3673);
xnor U5119 (N_5119,N_3873,N_4877);
nor U5120 (N_5120,N_3953,N_2691);
or U5121 (N_5121,N_4983,N_3204);
nand U5122 (N_5122,N_4456,N_4088);
nor U5123 (N_5123,N_3235,N_3960);
and U5124 (N_5124,N_3779,N_2591);
nor U5125 (N_5125,N_2784,N_3791);
nand U5126 (N_5126,N_2643,N_4996);
nor U5127 (N_5127,N_4542,N_4229);
or U5128 (N_5128,N_3674,N_3913);
nor U5129 (N_5129,N_3904,N_4327);
or U5130 (N_5130,N_4291,N_2604);
or U5131 (N_5131,N_4678,N_4303);
or U5132 (N_5132,N_4902,N_2561);
or U5133 (N_5133,N_4695,N_2937);
nand U5134 (N_5134,N_4166,N_3936);
or U5135 (N_5135,N_3538,N_2966);
xor U5136 (N_5136,N_3225,N_2799);
and U5137 (N_5137,N_3207,N_4477);
and U5138 (N_5138,N_3432,N_3360);
xnor U5139 (N_5139,N_4010,N_2836);
nor U5140 (N_5140,N_3840,N_4866);
nand U5141 (N_5141,N_4475,N_2975);
or U5142 (N_5142,N_3075,N_3620);
or U5143 (N_5143,N_4484,N_4410);
and U5144 (N_5144,N_4179,N_4574);
nor U5145 (N_5145,N_4259,N_3665);
nand U5146 (N_5146,N_4414,N_3797);
or U5147 (N_5147,N_2955,N_3256);
or U5148 (N_5148,N_3971,N_2886);
nand U5149 (N_5149,N_4553,N_2504);
and U5150 (N_5150,N_4657,N_3986);
xor U5151 (N_5151,N_3065,N_4037);
or U5152 (N_5152,N_4919,N_3787);
nand U5153 (N_5153,N_4596,N_4361);
and U5154 (N_5154,N_3316,N_4545);
or U5155 (N_5155,N_4378,N_4912);
or U5156 (N_5156,N_4510,N_4944);
xnor U5157 (N_5157,N_4130,N_4927);
and U5158 (N_5158,N_3570,N_3071);
or U5159 (N_5159,N_3066,N_3638);
and U5160 (N_5160,N_4565,N_3966);
and U5161 (N_5161,N_3700,N_4196);
or U5162 (N_5162,N_4977,N_4907);
nand U5163 (N_5163,N_3660,N_3226);
nor U5164 (N_5164,N_2759,N_3430);
xnor U5165 (N_5165,N_3183,N_3702);
and U5166 (N_5166,N_4764,N_4632);
or U5167 (N_5167,N_4425,N_3518);
nand U5168 (N_5168,N_2771,N_4112);
nor U5169 (N_5169,N_3194,N_2573);
nor U5170 (N_5170,N_2942,N_3557);
or U5171 (N_5171,N_4045,N_4195);
or U5172 (N_5172,N_2818,N_3663);
or U5173 (N_5173,N_4330,N_4573);
and U5174 (N_5174,N_4672,N_3682);
or U5175 (N_5175,N_4065,N_2817);
nor U5176 (N_5176,N_4294,N_4548);
nor U5177 (N_5177,N_4200,N_2658);
nor U5178 (N_5178,N_3626,N_4265);
or U5179 (N_5179,N_3166,N_3330);
or U5180 (N_5180,N_2920,N_4923);
or U5181 (N_5181,N_4472,N_3461);
nand U5182 (N_5182,N_2861,N_4356);
nand U5183 (N_5183,N_4879,N_4116);
nand U5184 (N_5184,N_4350,N_4298);
and U5185 (N_5185,N_3908,N_4125);
nand U5186 (N_5186,N_4406,N_4640);
nand U5187 (N_5187,N_3694,N_3243);
xnor U5188 (N_5188,N_4231,N_4607);
or U5189 (N_5189,N_4354,N_4040);
or U5190 (N_5190,N_3442,N_3425);
and U5191 (N_5191,N_2888,N_3516);
xnor U5192 (N_5192,N_3048,N_3363);
nor U5193 (N_5193,N_3558,N_3485);
xor U5194 (N_5194,N_2902,N_2885);
or U5195 (N_5195,N_4756,N_2528);
nor U5196 (N_5196,N_3107,N_2571);
nor U5197 (N_5197,N_4582,N_4871);
nor U5198 (N_5198,N_4384,N_2791);
nor U5199 (N_5199,N_4697,N_3124);
and U5200 (N_5200,N_3902,N_4945);
nand U5201 (N_5201,N_3408,N_4921);
nor U5202 (N_5202,N_2822,N_4067);
and U5203 (N_5203,N_4509,N_4020);
and U5204 (N_5204,N_4900,N_4114);
xnor U5205 (N_5205,N_3298,N_3864);
nor U5206 (N_5206,N_4424,N_4168);
or U5207 (N_5207,N_4086,N_4693);
nor U5208 (N_5208,N_2671,N_2632);
and U5209 (N_5209,N_3070,N_2606);
nand U5210 (N_5210,N_4990,N_3927);
nor U5211 (N_5211,N_3659,N_2685);
nand U5212 (N_5212,N_3136,N_4306);
or U5213 (N_5213,N_2789,N_3909);
or U5214 (N_5214,N_2923,N_4057);
nor U5215 (N_5215,N_2697,N_4227);
nor U5216 (N_5216,N_3024,N_2826);
nand U5217 (N_5217,N_3524,N_4207);
or U5218 (N_5218,N_3677,N_4436);
nor U5219 (N_5219,N_4393,N_4034);
nand U5220 (N_5220,N_2670,N_2819);
or U5221 (N_5221,N_4101,N_3991);
nor U5222 (N_5222,N_2514,N_3891);
and U5223 (N_5223,N_3507,N_2672);
nand U5224 (N_5224,N_3151,N_3364);
nand U5225 (N_5225,N_4613,N_3798);
nand U5226 (N_5226,N_3887,N_4257);
nor U5227 (N_5227,N_3283,N_4776);
xnor U5228 (N_5228,N_4396,N_4975);
and U5229 (N_5229,N_4843,N_3356);
nor U5230 (N_5230,N_4790,N_4884);
nand U5231 (N_5231,N_3567,N_4173);
and U5232 (N_5232,N_4646,N_2929);
nor U5233 (N_5233,N_3970,N_2773);
and U5234 (N_5234,N_2897,N_2712);
nand U5235 (N_5235,N_3457,N_4598);
and U5236 (N_5236,N_3859,N_4019);
nor U5237 (N_5237,N_2622,N_4575);
and U5238 (N_5238,N_3341,N_3009);
nor U5239 (N_5239,N_3441,N_4624);
and U5240 (N_5240,N_2970,N_3291);
or U5241 (N_5241,N_3296,N_3635);
and U5242 (N_5242,N_4238,N_3631);
nor U5243 (N_5243,N_3842,N_3762);
xor U5244 (N_5244,N_4138,N_4465);
nor U5245 (N_5245,N_3975,N_2904);
xnor U5246 (N_5246,N_3693,N_2778);
nor U5247 (N_5247,N_3132,N_2536);
and U5248 (N_5248,N_3336,N_4781);
or U5249 (N_5249,N_4743,N_2869);
or U5250 (N_5250,N_2565,N_2501);
or U5251 (N_5251,N_4920,N_3613);
nand U5252 (N_5252,N_3310,N_4749);
nor U5253 (N_5253,N_3618,N_4324);
nand U5254 (N_5254,N_4844,N_4534);
nor U5255 (N_5255,N_3979,N_2535);
or U5256 (N_5256,N_2914,N_2530);
nand U5257 (N_5257,N_2972,N_4667);
or U5258 (N_5258,N_4276,N_4911);
nor U5259 (N_5259,N_3750,N_2509);
or U5260 (N_5260,N_4452,N_4184);
nor U5261 (N_5261,N_4469,N_3816);
nor U5262 (N_5262,N_4704,N_3625);
and U5263 (N_5263,N_4616,N_2765);
and U5264 (N_5264,N_3656,N_3086);
nor U5265 (N_5265,N_3705,N_4219);
nand U5266 (N_5266,N_3521,N_4141);
nand U5267 (N_5267,N_3747,N_4023);
and U5268 (N_5268,N_2520,N_3387);
nand U5269 (N_5269,N_2585,N_3329);
and U5270 (N_5270,N_3860,N_4543);
or U5271 (N_5271,N_2906,N_4333);
or U5272 (N_5272,N_3028,N_4146);
nand U5273 (N_5273,N_3534,N_2666);
and U5274 (N_5274,N_4003,N_3681);
and U5275 (N_5275,N_3393,N_3769);
nand U5276 (N_5276,N_3091,N_3250);
xnor U5277 (N_5277,N_3046,N_3097);
or U5278 (N_5278,N_3251,N_4727);
and U5279 (N_5279,N_4740,N_2743);
and U5280 (N_5280,N_2856,N_3717);
xor U5281 (N_5281,N_3907,N_3906);
nor U5282 (N_5282,N_4712,N_4571);
nand U5283 (N_5283,N_4810,N_3383);
nand U5284 (N_5284,N_3811,N_4674);
and U5285 (N_5285,N_4342,N_3560);
nand U5286 (N_5286,N_4395,N_3574);
nand U5287 (N_5287,N_4343,N_2951);
nand U5288 (N_5288,N_4698,N_3733);
nor U5289 (N_5289,N_3263,N_4531);
nand U5290 (N_5290,N_2729,N_3527);
or U5291 (N_5291,N_4736,N_3332);
nor U5292 (N_5292,N_2746,N_4556);
nor U5293 (N_5293,N_2957,N_3643);
nor U5294 (N_5294,N_2919,N_4011);
nand U5295 (N_5295,N_2596,N_4665);
or U5296 (N_5296,N_2724,N_4015);
xor U5297 (N_5297,N_3051,N_4400);
and U5298 (N_5298,N_4815,N_2564);
nor U5299 (N_5299,N_4677,N_2676);
nor U5300 (N_5300,N_4555,N_4172);
nor U5301 (N_5301,N_3794,N_2508);
and U5302 (N_5302,N_3147,N_2619);
or U5303 (N_5303,N_4965,N_2597);
xnor U5304 (N_5304,N_3844,N_4385);
nand U5305 (N_5305,N_2736,N_4336);
or U5306 (N_5306,N_4572,N_2763);
or U5307 (N_5307,N_3784,N_3857);
and U5308 (N_5308,N_4560,N_2711);
nand U5309 (N_5309,N_3780,N_2892);
or U5310 (N_5310,N_2660,N_4522);
nor U5311 (N_5311,N_3477,N_2522);
or U5312 (N_5312,N_3386,N_3131);
nor U5313 (N_5313,N_2667,N_4694);
and U5314 (N_5314,N_4714,N_2580);
nor U5315 (N_5315,N_4612,N_3861);
or U5316 (N_5316,N_3939,N_3868);
xor U5317 (N_5317,N_3023,N_4331);
and U5318 (N_5318,N_4024,N_3369);
or U5319 (N_5319,N_3743,N_3876);
xnor U5320 (N_5320,N_2777,N_4164);
nand U5321 (N_5321,N_2754,N_3427);
and U5322 (N_5322,N_4929,N_4413);
nor U5323 (N_5323,N_3604,N_4144);
nand U5324 (N_5324,N_4804,N_4512);
and U5325 (N_5325,N_4634,N_2713);
nand U5326 (N_5326,N_4422,N_4075);
xor U5327 (N_5327,N_3142,N_2503);
nor U5328 (N_5328,N_3862,N_3029);
nor U5329 (N_5329,N_2583,N_3785);
nor U5330 (N_5330,N_4734,N_3407);
nor U5331 (N_5331,N_4250,N_2753);
nand U5332 (N_5332,N_2719,N_4586);
or U5333 (N_5333,N_4935,N_2615);
nor U5334 (N_5334,N_3735,N_3082);
nand U5335 (N_5335,N_4583,N_3912);
nand U5336 (N_5336,N_4187,N_4357);
or U5337 (N_5337,N_3502,N_3154);
xor U5338 (N_5338,N_4193,N_2824);
xor U5339 (N_5339,N_4833,N_3465);
nand U5340 (N_5340,N_3260,N_4329);
nor U5341 (N_5341,N_3447,N_3122);
and U5342 (N_5342,N_2908,N_3079);
or U5343 (N_5343,N_2761,N_4111);
and U5344 (N_5344,N_4286,N_3575);
and U5345 (N_5345,N_3850,N_3822);
and U5346 (N_5346,N_3398,N_2934);
nor U5347 (N_5347,N_2837,N_4865);
and U5348 (N_5348,N_2624,N_2965);
or U5349 (N_5349,N_4236,N_3168);
or U5350 (N_5350,N_3684,N_4163);
nor U5351 (N_5351,N_2545,N_3703);
or U5352 (N_5352,N_4769,N_3888);
nor U5353 (N_5353,N_3832,N_4706);
nor U5354 (N_5354,N_2633,N_3541);
or U5355 (N_5355,N_3985,N_4850);
nand U5356 (N_5356,N_4098,N_3954);
or U5357 (N_5357,N_3493,N_4334);
and U5358 (N_5358,N_3957,N_4131);
and U5359 (N_5359,N_3526,N_3824);
nand U5360 (N_5360,N_4948,N_3820);
nand U5361 (N_5361,N_4540,N_4212);
nand U5362 (N_5362,N_3139,N_4174);
xor U5363 (N_5363,N_4471,N_3466);
or U5364 (N_5364,N_2738,N_2989);
and U5365 (N_5365,N_3252,N_3505);
nor U5366 (N_5366,N_3357,N_3930);
or U5367 (N_5367,N_2627,N_4069);
and U5368 (N_5368,N_3670,N_2981);
xor U5369 (N_5369,N_4022,N_4847);
nand U5370 (N_5370,N_3597,N_3812);
or U5371 (N_5371,N_3917,N_4982);
nor U5372 (N_5372,N_4619,N_3491);
nand U5373 (N_5373,N_3504,N_4861);
or U5374 (N_5374,N_4533,N_4602);
and U5375 (N_5375,N_3293,N_4304);
and U5376 (N_5376,N_3737,N_3867);
or U5377 (N_5377,N_2502,N_4763);
and U5378 (N_5378,N_4938,N_3544);
nand U5379 (N_5379,N_4435,N_4660);
nand U5380 (N_5380,N_2556,N_3899);
and U5381 (N_5381,N_4590,N_3577);
nand U5382 (N_5382,N_3531,N_4784);
nor U5383 (N_5383,N_3016,N_4245);
or U5384 (N_5384,N_4679,N_2605);
xor U5385 (N_5385,N_2858,N_3355);
xnor U5386 (N_5386,N_4450,N_3872);
xnor U5387 (N_5387,N_2629,N_4416);
or U5388 (N_5388,N_4243,N_4242);
nand U5389 (N_5389,N_4483,N_3839);
nand U5390 (N_5390,N_2531,N_3445);
or U5391 (N_5391,N_3005,N_4638);
or U5392 (N_5392,N_3932,N_4526);
or U5393 (N_5393,N_4789,N_3394);
or U5394 (N_5394,N_2646,N_3175);
xnor U5395 (N_5395,N_3008,N_3572);
and U5396 (N_5396,N_3173,N_4668);
nor U5397 (N_5397,N_4755,N_4169);
and U5398 (N_5398,N_3094,N_4221);
nand U5399 (N_5399,N_3453,N_2529);
and U5400 (N_5400,N_4322,N_3602);
and U5401 (N_5401,N_4760,N_4440);
xor U5402 (N_5402,N_4405,N_3468);
nor U5403 (N_5403,N_4893,N_4585);
nand U5404 (N_5404,N_2757,N_4924);
nor U5405 (N_5405,N_3883,N_3025);
and U5406 (N_5406,N_2749,N_3655);
nor U5407 (N_5407,N_4104,N_3484);
nor U5408 (N_5408,N_2642,N_4610);
and U5409 (N_5409,N_2625,N_4490);
nand U5410 (N_5410,N_3367,N_4423);
and U5411 (N_5411,N_4094,N_2767);
nor U5412 (N_5412,N_4345,N_3216);
xor U5413 (N_5413,N_2750,N_4237);
nand U5414 (N_5414,N_2808,N_3039);
and U5415 (N_5415,N_4828,N_3013);
xnor U5416 (N_5416,N_4204,N_3300);
nand U5417 (N_5417,N_4316,N_3181);
and U5418 (N_5418,N_4642,N_4787);
xor U5419 (N_5419,N_4899,N_4255);
nor U5420 (N_5420,N_4143,N_4030);
nand U5421 (N_5421,N_3495,N_2659);
nor U5422 (N_5422,N_4747,N_4569);
xor U5423 (N_5423,N_4711,N_2991);
or U5424 (N_5424,N_2579,N_4930);
nand U5425 (N_5425,N_3179,N_3734);
and U5426 (N_5426,N_3419,N_4680);
and U5427 (N_5427,N_3948,N_3706);
and U5428 (N_5428,N_2927,N_3133);
or U5429 (N_5429,N_4960,N_4052);
or U5430 (N_5430,N_3918,N_4922);
nor U5431 (N_5431,N_4805,N_4439);
xor U5432 (N_5432,N_3691,N_4408);
xor U5433 (N_5433,N_3205,N_3189);
and U5434 (N_5434,N_4382,N_3903);
nor U5435 (N_5435,N_4185,N_3633);
or U5436 (N_5436,N_3406,N_3267);
or U5437 (N_5437,N_3138,N_4675);
and U5438 (N_5438,N_2600,N_3829);
nor U5439 (N_5439,N_4407,N_2800);
or U5440 (N_5440,N_4687,N_2898);
and U5441 (N_5441,N_3358,N_3582);
nor U5442 (N_5442,N_3346,N_4177);
or U5443 (N_5443,N_3368,N_4103);
or U5444 (N_5444,N_2994,N_3451);
or U5445 (N_5445,N_4403,N_2704);
and U5446 (N_5446,N_4148,N_2973);
and U5447 (N_5447,N_2862,N_4417);
or U5448 (N_5448,N_4901,N_2731);
xnor U5449 (N_5449,N_2500,N_2842);
nand U5450 (N_5450,N_3745,N_4344);
or U5451 (N_5451,N_3487,N_4394);
or U5452 (N_5452,N_2523,N_4419);
and U5453 (N_5453,N_4310,N_3514);
or U5454 (N_5454,N_4441,N_3072);
or U5455 (N_5455,N_2703,N_2859);
or U5456 (N_5456,N_4036,N_4552);
nand U5457 (N_5457,N_4005,N_3874);
nand U5458 (N_5458,N_3371,N_3392);
nand U5459 (N_5459,N_2969,N_2540);
and U5460 (N_5460,N_2557,N_3472);
nand U5461 (N_5461,N_2882,N_2558);
and U5462 (N_5462,N_3253,N_4364);
nor U5463 (N_5463,N_4525,N_3551);
and U5464 (N_5464,N_3404,N_2893);
and U5465 (N_5465,N_2512,N_4803);
nor U5466 (N_5466,N_4617,N_4791);
or U5467 (N_5467,N_4709,N_4830);
and U5468 (N_5468,N_4188,N_4376);
and U5469 (N_5469,N_3580,N_4254);
or U5470 (N_5470,N_3501,N_2868);
nor U5471 (N_5471,N_3185,N_2527);
and U5472 (N_5472,N_3087,N_3223);
nor U5473 (N_5473,N_3322,N_3033);
or U5474 (N_5474,N_4550,N_4216);
and U5475 (N_5475,N_3349,N_3776);
nor U5476 (N_5476,N_2823,N_4399);
nand U5477 (N_5477,N_4102,N_3509);
and U5478 (N_5478,N_3807,N_4014);
and U5479 (N_5479,N_4949,N_3146);
nor U5480 (N_5480,N_3808,N_3438);
and U5481 (N_5481,N_3340,N_3981);
nor U5482 (N_5482,N_2963,N_3914);
or U5483 (N_5483,N_3778,N_2567);
or U5484 (N_5484,N_2948,N_4274);
nor U5485 (N_5485,N_2510,N_4707);
or U5486 (N_5486,N_4941,N_3257);
xor U5487 (N_5487,N_3601,N_4026);
nand U5488 (N_5488,N_3576,N_4135);
nor U5489 (N_5489,N_3058,N_2883);
or U5490 (N_5490,N_4986,N_4044);
xor U5491 (N_5491,N_4659,N_2537);
xnor U5492 (N_5492,N_3821,N_3218);
xnor U5493 (N_5493,N_3117,N_4081);
nand U5494 (N_5494,N_3803,N_4054);
and U5495 (N_5495,N_2737,N_4429);
or U5496 (N_5496,N_3297,N_4943);
xnor U5497 (N_5497,N_2524,N_4988);
or U5498 (N_5498,N_4953,N_2569);
nor U5499 (N_5499,N_2613,N_4122);
and U5500 (N_5500,N_3000,N_3827);
and U5501 (N_5501,N_4028,N_3289);
and U5502 (N_5502,N_4663,N_4873);
nor U5503 (N_5503,N_3753,N_2631);
nor U5504 (N_5504,N_3513,N_3915);
nor U5505 (N_5505,N_4473,N_2905);
or U5506 (N_5506,N_4870,N_2584);
or U5507 (N_5507,N_4032,N_2518);
xnor U5508 (N_5508,N_2867,N_3946);
or U5509 (N_5509,N_3019,N_4217);
nor U5510 (N_5510,N_4127,N_4980);
and U5511 (N_5511,N_3458,N_3269);
and U5512 (N_5512,N_4317,N_3727);
nor U5513 (N_5513,N_3239,N_4120);
or U5514 (N_5514,N_2964,N_4753);
or U5515 (N_5515,N_2925,N_4346);
and U5516 (N_5516,N_3830,N_4775);
nand U5517 (N_5517,N_3116,N_2766);
xor U5518 (N_5518,N_3961,N_4639);
nand U5519 (N_5519,N_4314,N_3983);
nand U5520 (N_5520,N_3758,N_4448);
or U5521 (N_5521,N_3802,N_2811);
nor U5522 (N_5522,N_3563,N_3943);
or U5523 (N_5523,N_3999,N_3098);
and U5524 (N_5524,N_3742,N_3648);
or U5525 (N_5525,N_4107,N_4090);
or U5526 (N_5526,N_3435,N_4315);
nand U5527 (N_5527,N_4951,N_4318);
nor U5528 (N_5528,N_4320,N_2865);
nor U5529 (N_5529,N_4485,N_3566);
xnor U5530 (N_5530,N_3621,N_3467);
or U5531 (N_5531,N_4530,N_4047);
nor U5532 (N_5532,N_4124,N_2903);
or U5533 (N_5533,N_4852,N_4658);
or U5534 (N_5534,N_3591,N_3678);
or U5535 (N_5535,N_4332,N_4411);
or U5536 (N_5536,N_3856,N_3063);
nand U5537 (N_5537,N_3994,N_4249);
or U5538 (N_5538,N_4954,N_2852);
or U5539 (N_5539,N_3057,N_3374);
nor U5540 (N_5540,N_3230,N_4189);
nand U5541 (N_5541,N_3177,N_3771);
or U5542 (N_5542,N_4311,N_2668);
and U5543 (N_5543,N_3021,N_3801);
nor U5544 (N_5544,N_4557,N_4701);
and U5545 (N_5545,N_3074,N_2692);
or U5546 (N_5546,N_3174,N_4956);
nand U5547 (N_5547,N_4853,N_2542);
and U5548 (N_5548,N_4561,N_3492);
or U5549 (N_5549,N_4772,N_3628);
and U5550 (N_5550,N_4162,N_4963);
or U5551 (N_5551,N_2839,N_2889);
nand U5552 (N_5552,N_3882,N_3402);
nor U5553 (N_5553,N_2995,N_3379);
or U5554 (N_5554,N_3636,N_4750);
nor U5555 (N_5555,N_3593,N_2551);
or U5556 (N_5556,N_2742,N_4063);
and U5557 (N_5557,N_4738,N_4645);
nand U5558 (N_5558,N_4795,N_2592);
nor U5559 (N_5559,N_3089,N_3905);
and U5560 (N_5560,N_4241,N_4266);
nor U5561 (N_5561,N_2947,N_3149);
or U5562 (N_5562,N_4942,N_3757);
and U5563 (N_5563,N_3049,N_4751);
nand U5564 (N_5564,N_4494,N_3059);
nand U5565 (N_5565,N_4035,N_3232);
nand U5566 (N_5566,N_4767,N_3426);
nor U5567 (N_5567,N_3217,N_3067);
and U5568 (N_5568,N_3615,N_3878);
nand U5569 (N_5569,N_4012,N_3272);
or U5570 (N_5570,N_3306,N_4739);
xor U5571 (N_5571,N_3546,N_4213);
or U5572 (N_5572,N_4401,N_4592);
and U5573 (N_5573,N_3270,N_4972);
nand U5574 (N_5574,N_4779,N_2873);
or U5575 (N_5575,N_4588,N_4816);
or U5576 (N_5576,N_2933,N_2755);
and U5577 (N_5577,N_2727,N_4302);
nor U5578 (N_5578,N_3547,N_2875);
or U5579 (N_5579,N_4372,N_2628);
xnor U5580 (N_5580,N_4774,N_4608);
nor U5581 (N_5581,N_3099,N_4077);
nand U5582 (N_5582,N_4863,N_3559);
xor U5583 (N_5583,N_2938,N_3069);
nand U5584 (N_5584,N_4683,N_3268);
nand U5585 (N_5585,N_3157,N_2657);
nand U5586 (N_5586,N_4794,N_2513);
nand U5587 (N_5587,N_2519,N_3723);
nand U5588 (N_5588,N_3923,N_3167);
nand U5589 (N_5589,N_3653,N_2696);
nor U5590 (N_5590,N_3599,N_2578);
and U5591 (N_5591,N_3305,N_3760);
nand U5592 (N_5592,N_4281,N_3366);
or U5593 (N_5593,N_3325,N_3412);
nand U5594 (N_5594,N_3228,N_3616);
nor U5595 (N_5595,N_2801,N_4813);
nand U5596 (N_5596,N_3503,N_2857);
and U5597 (N_5597,N_3764,N_3896);
nand U5598 (N_5598,N_3834,N_3343);
and U5599 (N_5599,N_2814,N_4041);
nand U5600 (N_5600,N_3130,N_3429);
nor U5601 (N_5601,N_3853,N_3444);
nor U5602 (N_5602,N_4115,N_4589);
nand U5603 (N_5603,N_2638,N_3141);
or U5604 (N_5604,N_2971,N_4062);
nor U5605 (N_5605,N_3848,N_3384);
or U5606 (N_5606,N_4149,N_3805);
nand U5607 (N_5607,N_3708,N_4046);
nand U5608 (N_5608,N_4380,N_2559);
nand U5609 (N_5609,N_3378,N_3481);
nand U5610 (N_5610,N_3721,N_4925);
nand U5611 (N_5611,N_4128,N_3288);
and U5612 (N_5612,N_4547,N_3799);
nor U5613 (N_5613,N_2610,N_4631);
nor U5614 (N_5614,N_3299,N_4818);
nor U5615 (N_5615,N_4962,N_4239);
or U5616 (N_5616,N_3261,N_3922);
or U5617 (N_5617,N_4199,N_4742);
or U5618 (N_5618,N_2976,N_3399);
nor U5619 (N_5619,N_2953,N_4984);
nand U5620 (N_5620,N_4055,N_3328);
nand U5621 (N_5621,N_3645,N_3273);
and U5622 (N_5622,N_3199,N_4995);
or U5623 (N_5623,N_3644,N_3161);
and U5624 (N_5624,N_2507,N_4615);
or U5625 (N_5625,N_4209,N_4386);
xnor U5626 (N_5626,N_3434,N_3084);
nand U5627 (N_5627,N_4931,N_3800);
and U5628 (N_5628,N_4913,N_2788);
nor U5629 (N_5629,N_2774,N_4273);
nor U5630 (N_5630,N_3083,N_3522);
nand U5631 (N_5631,N_3125,N_3696);
and U5632 (N_5632,N_2781,N_4068);
or U5633 (N_5633,N_4338,N_2996);
xor U5634 (N_5634,N_2881,N_3007);
or U5635 (N_5635,N_4095,N_3947);
xor U5636 (N_5636,N_4967,N_4491);
nand U5637 (N_5637,N_3755,N_3456);
nor U5638 (N_5638,N_3055,N_4745);
or U5639 (N_5639,N_3763,N_4300);
or U5640 (N_5640,N_4689,N_2877);
xnor U5641 (N_5641,N_3353,N_3980);
and U5642 (N_5642,N_4297,N_4591);
or U5643 (N_5643,N_3112,N_3790);
and U5644 (N_5644,N_3135,N_3639);
nand U5645 (N_5645,N_3898,N_4716);
or U5646 (N_5646,N_3282,N_4083);
nand U5647 (N_5647,N_4834,N_3624);
nor U5648 (N_5648,N_3100,N_3352);
nand U5649 (N_5649,N_4224,N_2949);
nor U5650 (N_5650,N_4845,N_3666);
nand U5651 (N_5651,N_3222,N_2768);
or U5652 (N_5652,N_4812,N_3164);
nand U5653 (N_5653,N_4262,N_4890);
and U5654 (N_5654,N_4946,N_3258);
and U5655 (N_5655,N_3095,N_3077);
nand U5656 (N_5656,N_3679,N_2566);
and U5657 (N_5657,N_4222,N_3265);
nor U5658 (N_5658,N_4564,N_3080);
or U5659 (N_5659,N_3396,N_3950);
nor U5660 (N_5660,N_4754,N_3191);
nand U5661 (N_5661,N_3713,N_3793);
xnor U5662 (N_5662,N_4109,N_2677);
nor U5663 (N_5663,N_4897,N_3606);
xnor U5664 (N_5664,N_4252,N_4373);
nor U5665 (N_5665,N_3400,N_3050);
nand U5666 (N_5666,N_4748,N_3517);
and U5667 (N_5667,N_3115,N_4947);
or U5668 (N_5668,N_2516,N_3262);
or U5669 (N_5669,N_4495,N_4976);
or U5670 (N_5670,N_4497,N_2714);
or U5671 (N_5671,N_4328,N_2752);
or U5672 (N_5672,N_3313,N_3375);
nor U5673 (N_5673,N_4389,N_4688);
or U5674 (N_5674,N_3925,N_4662);
nand U5675 (N_5675,N_2616,N_4321);
or U5676 (N_5676,N_4883,N_3026);
or U5677 (N_5677,N_3823,N_3770);
xor U5678 (N_5678,N_4595,N_3347);
nand U5679 (N_5679,N_3835,N_4482);
and U5680 (N_5680,N_4817,N_3556);
xnor U5681 (N_5681,N_3473,N_2816);
nor U5682 (N_5682,N_2834,N_4208);
nand U5683 (N_5683,N_3197,N_3497);
or U5684 (N_5684,N_2640,N_4374);
nor U5685 (N_5685,N_2708,N_3076);
or U5686 (N_5686,N_3963,N_3469);
and U5687 (N_5687,N_4987,N_3119);
and U5688 (N_5688,N_3726,N_3782);
and U5689 (N_5689,N_3038,N_4841);
xnor U5690 (N_5690,N_3031,N_3278);
nand U5691 (N_5691,N_4966,N_3945);
nand U5692 (N_5692,N_4106,N_3652);
nand U5693 (N_5693,N_3796,N_4438);
or U5694 (N_5694,N_2682,N_3213);
xnor U5695 (N_5695,N_3610,N_3833);
or U5696 (N_5696,N_4622,N_3751);
nand U5697 (N_5697,N_3894,N_2730);
and U5698 (N_5698,N_2828,N_2563);
nand U5699 (N_5699,N_4896,N_4136);
and U5700 (N_5700,N_4493,N_3942);
xor U5701 (N_5701,N_2845,N_3955);
nor U5702 (N_5702,N_2855,N_4282);
nor U5703 (N_5703,N_4521,N_2807);
nor U5704 (N_5704,N_3537,N_4358);
or U5705 (N_5705,N_4479,N_4268);
xnor U5706 (N_5706,N_3738,N_3573);
nand U5707 (N_5707,N_3244,N_2764);
or U5708 (N_5708,N_2612,N_3342);
and U5709 (N_5709,N_2555,N_4539);
or U5710 (N_5710,N_3416,N_2718);
or U5711 (N_5711,N_3200,N_4165);
xnor U5712 (N_5712,N_4758,N_2779);
xnor U5713 (N_5713,N_4156,N_2539);
and U5714 (N_5714,N_4501,N_3047);
or U5715 (N_5715,N_4492,N_3792);
and U5716 (N_5716,N_3397,N_3499);
xnor U5717 (N_5717,N_2651,N_4682);
nor U5718 (N_5718,N_3650,N_4614);
nor U5719 (N_5719,N_3765,N_3933);
and U5720 (N_5720,N_2686,N_3036);
and U5721 (N_5721,N_3587,N_2878);
xnor U5722 (N_5722,N_3964,N_3692);
nor U5723 (N_5723,N_2910,N_4234);
xnor U5724 (N_5724,N_2999,N_4025);
and U5725 (N_5725,N_4874,N_3858);
or U5726 (N_5726,N_3795,N_4009);
or U5727 (N_5727,N_4703,N_4280);
nand U5728 (N_5728,N_3523,N_4004);
nand U5729 (N_5729,N_4064,N_3178);
nor U5730 (N_5730,N_4800,N_4061);
and U5731 (N_5731,N_4604,N_4186);
and U5732 (N_5732,N_4837,N_4746);
nor U5733 (N_5733,N_4323,N_2803);
and U5734 (N_5734,N_3783,N_3471);
and U5735 (N_5735,N_3018,N_2663);
and U5736 (N_5736,N_3773,N_2841);
nor U5737 (N_5737,N_4341,N_4524);
and U5738 (N_5738,N_3536,N_3221);
nor U5739 (N_5739,N_4039,N_4969);
xnor U5740 (N_5740,N_2594,N_2598);
or U5741 (N_5741,N_3237,N_3042);
nor U5742 (N_5742,N_4474,N_3843);
nand U5743 (N_5743,N_4299,N_3277);
or U5744 (N_5744,N_4443,N_2921);
and U5745 (N_5745,N_3990,N_3292);
and U5746 (N_5746,N_4860,N_3992);
nand U5747 (N_5747,N_3884,N_3249);
or U5748 (N_5748,N_4059,N_4397);
nor U5749 (N_5749,N_2588,N_3462);
nand U5750 (N_5750,N_2772,N_4655);
or U5751 (N_5751,N_3220,N_4686);
and U5752 (N_5752,N_2634,N_4309);
and U5753 (N_5753,N_4627,N_4783);
or U5754 (N_5754,N_4857,N_3686);
and U5755 (N_5755,N_4402,N_3595);
nand U5756 (N_5756,N_2716,N_3974);
or U5757 (N_5757,N_3711,N_4858);
or U5758 (N_5758,N_2827,N_4699);
nor U5759 (N_5759,N_4952,N_4263);
xor U5760 (N_5760,N_4481,N_3203);
nor U5761 (N_5761,N_3506,N_4351);
xnor U5762 (N_5762,N_2932,N_3609);
nor U5763 (N_5763,N_4587,N_3826);
or U5764 (N_5764,N_3062,N_4463);
or U5765 (N_5765,N_4752,N_4048);
and U5766 (N_5766,N_4726,N_3303);
nor U5767 (N_5767,N_3170,N_3478);
and U5768 (N_5768,N_3376,N_3836);
or U5769 (N_5769,N_4412,N_4718);
or U5770 (N_5770,N_4528,N_3640);
or U5771 (N_5771,N_3440,N_3761);
and U5772 (N_5772,N_2922,N_2532);
nor U5773 (N_5773,N_4287,N_4272);
xnor U5774 (N_5774,N_4721,N_3437);
nand U5775 (N_5775,N_4599,N_4581);
nand U5776 (N_5776,N_2608,N_3061);
nor U5777 (N_5777,N_4451,N_4134);
nor U5778 (N_5778,N_3120,N_4427);
nor U5779 (N_5779,N_3688,N_4108);
and U5780 (N_5780,N_2806,N_4319);
and U5781 (N_5781,N_3561,N_3159);
nand U5782 (N_5782,N_3339,N_2960);
xor U5783 (N_5783,N_4782,N_4541);
or U5784 (N_5784,N_4225,N_3323);
or U5785 (N_5785,N_4498,N_3171);
and U5786 (N_5786,N_2760,N_4021);
or U5787 (N_5787,N_3984,N_2879);
nand U5788 (N_5788,N_3831,N_3555);
nand U5789 (N_5789,N_3929,N_3040);
and U5790 (N_5790,N_4446,N_2586);
and U5791 (N_5791,N_3482,N_4366);
nand U5792 (N_5792,N_3489,N_3012);
and U5793 (N_5793,N_3539,N_4089);
xor U5794 (N_5794,N_4458,N_4453);
nand U5795 (N_5795,N_4349,N_3627);
and U5796 (N_5796,N_2998,N_3034);
nor U5797 (N_5797,N_4183,N_2952);
or U5798 (N_5798,N_4381,N_3877);
nor U5799 (N_5799,N_3331,N_2652);
or U5800 (N_5800,N_3345,N_4580);
and U5801 (N_5801,N_4864,N_2812);
nor U5802 (N_5802,N_3307,N_3710);
nor U5803 (N_5803,N_3658,N_4160);
xor U5804 (N_5804,N_3545,N_3003);
nand U5805 (N_5805,N_4178,N_2967);
and U5806 (N_5806,N_4228,N_2684);
nor U5807 (N_5807,N_4151,N_4460);
or U5808 (N_5808,N_3103,N_3295);
nand U5809 (N_5809,N_2795,N_3956);
or U5810 (N_5810,N_2574,N_4839);
or U5811 (N_5811,N_4702,N_3184);
nor U5812 (N_5812,N_3276,N_2700);
nor U5813 (N_5813,N_3333,N_2829);
nor U5814 (N_5814,N_3454,N_3410);
and U5815 (N_5815,N_3450,N_3976);
xor U5816 (N_5816,N_4532,N_3890);
or U5817 (N_5817,N_4985,N_4359);
nor U5818 (N_5818,N_4806,N_3287);
nand U5819 (N_5819,N_2851,N_2940);
nor U5820 (N_5820,N_3549,N_3749);
or U5821 (N_5821,N_4308,N_4880);
and U5822 (N_5822,N_4486,N_4868);
and U5823 (N_5823,N_4720,N_2581);
nor U5824 (N_5824,N_3326,N_2726);
or U5825 (N_5825,N_4829,N_4240);
nand U5826 (N_5826,N_4507,N_3689);
nor U5827 (N_5827,N_4516,N_3114);
nor U5828 (N_5828,N_4878,N_3362);
and U5829 (N_5829,N_2866,N_3377);
and U5830 (N_5830,N_3145,N_3759);
nand U5831 (N_5831,N_3101,N_4367);
nor U5832 (N_5832,N_3134,N_4700);
nand U5833 (N_5833,N_4370,N_3417);
nor U5834 (N_5834,N_4499,N_4855);
nand U5835 (N_5835,N_3421,N_4277);
nor U5836 (N_5836,N_3290,N_4649);
nor U5837 (N_5837,N_3152,N_3671);
and U5838 (N_5838,N_2543,N_4535);
or U5839 (N_5839,N_2962,N_4684);
or U5840 (N_5840,N_3096,N_3388);
nand U5841 (N_5841,N_3715,N_3234);
nor U5842 (N_5842,N_2918,N_3683);
nand U5843 (N_5843,N_2732,N_4462);
or U5844 (N_5844,N_2912,N_3015);
nor U5845 (N_5845,N_3605,N_3662);
nor U5846 (N_5846,N_2541,N_3027);
nand U5847 (N_5847,N_3334,N_3206);
nand U5848 (N_5848,N_2769,N_2935);
and U5849 (N_5849,N_2611,N_4968);
and U5850 (N_5850,N_3697,N_4223);
nand U5851 (N_5851,N_4233,N_4371);
or U5852 (N_5852,N_3603,N_2987);
and U5853 (N_5853,N_2637,N_3748);
and U5854 (N_5854,N_2810,N_4696);
xnor U5855 (N_5855,N_2630,N_4428);
or U5856 (N_5856,N_3752,N_2815);
and U5857 (N_5857,N_4759,N_2880);
xor U5858 (N_5858,N_3428,N_4831);
or U5859 (N_5859,N_2830,N_3813);
nand U5860 (N_5860,N_3525,N_4056);
nor U5861 (N_5861,N_3348,N_3810);
or U5862 (N_5862,N_4335,N_4470);
or U5863 (N_5863,N_2748,N_2974);
nor U5864 (N_5864,N_4958,N_4365);
xnor U5865 (N_5865,N_4383,N_2977);
nor U5866 (N_5866,N_4049,N_4822);
or U5867 (N_5867,N_4279,N_4363);
or U5868 (N_5868,N_2762,N_4091);
nand U5869 (N_5869,N_3910,N_3372);
or U5870 (N_5870,N_3919,N_3825);
nor U5871 (N_5871,N_4626,N_3612);
and U5872 (N_5872,N_4916,N_4989);
xnor U5873 (N_5873,N_2715,N_3474);
nor U5874 (N_5874,N_3542,N_2891);
or U5875 (N_5875,N_3460,N_3712);
nand U5876 (N_5876,N_4180,N_4889);
nand U5877 (N_5877,N_2538,N_3255);
nand U5878 (N_5878,N_4167,N_4362);
nor U5879 (N_5879,N_2988,N_4766);
xor U5880 (N_5880,N_3937,N_4220);
nor U5881 (N_5881,N_4226,N_2783);
xor U5882 (N_5882,N_4797,N_4620);
and U5883 (N_5883,N_4100,N_4904);
or U5884 (N_5884,N_2946,N_4881);
and U5885 (N_5885,N_3654,N_3817);
and U5886 (N_5886,N_4339,N_3286);
xnor U5887 (N_5887,N_4869,N_3448);
and U5888 (N_5888,N_4071,N_2870);
nand U5889 (N_5889,N_3113,N_3245);
nor U5890 (N_5890,N_4554,N_4671);
nor U5891 (N_5891,N_2876,N_4278);
nand U5892 (N_5892,N_3530,N_3370);
and U5893 (N_5893,N_2980,N_3866);
nand U5894 (N_5894,N_3317,N_4430);
or U5895 (N_5895,N_3695,N_4885);
nor U5896 (N_5896,N_3996,N_3554);
nand U5897 (N_5897,N_2688,N_3498);
nand U5898 (N_5898,N_3608,N_3818);
or U5899 (N_5899,N_3202,N_3318);
or U5900 (N_5900,N_4544,N_2694);
or U5901 (N_5901,N_4605,N_2850);
nand U5902 (N_5902,N_3350,N_2917);
nor U5903 (N_5903,N_4093,N_4211);
or U5904 (N_5904,N_4230,N_4867);
or U5905 (N_5905,N_2553,N_4284);
nand U5906 (N_5906,N_3464,N_4959);
nor U5907 (N_5907,N_4398,N_3592);
nor U5908 (N_5908,N_2639,N_4936);
nand U5909 (N_5909,N_4762,N_2813);
and U5910 (N_5910,N_4119,N_2751);
xnor U5911 (N_5911,N_4051,N_3043);
nor U5912 (N_5912,N_2835,N_3236);
or U5913 (N_5913,N_4737,N_3172);
xnor U5914 (N_5914,N_4191,N_2958);
nand U5915 (N_5915,N_2844,N_4515);
xnor U5916 (N_5916,N_4404,N_3880);
xor U5917 (N_5917,N_3294,N_3335);
nor U5918 (N_5918,N_4842,N_3634);
nor U5919 (N_5919,N_2894,N_4145);
nor U5920 (N_5920,N_4717,N_4523);
nand U5921 (N_5921,N_4609,N_3588);
xor U5922 (N_5922,N_4043,N_2548);
and U5923 (N_5923,N_4647,N_2607);
or U5924 (N_5924,N_3846,N_2679);
nor U5925 (N_5925,N_3809,N_4377);
and U5926 (N_5926,N_2956,N_4053);
or U5927 (N_5927,N_4437,N_4097);
nor U5928 (N_5928,N_3081,N_3248);
nand U5929 (N_5929,N_4017,N_2593);
nor U5930 (N_5930,N_3214,N_3607);
and U5931 (N_5931,N_3391,N_4391);
nand U5932 (N_5932,N_4181,N_3938);
or U5933 (N_5933,N_3657,N_4765);
nand U5934 (N_5934,N_3921,N_3496);
or U5935 (N_5935,N_3651,N_3617);
xnor U5936 (N_5936,N_2849,N_2654);
nand U5937 (N_5937,N_3837,N_4434);
or U5938 (N_5938,N_3052,N_2911);
or U5939 (N_5939,N_3470,N_2582);
nand U5940 (N_5940,N_4013,N_3892);
and U5941 (N_5941,N_2554,N_2821);
xor U5942 (N_5942,N_4392,N_3321);
nor U5943 (N_5943,N_4468,N_2599);
nand U5944 (N_5944,N_4455,N_3732);
or U5945 (N_5945,N_3728,N_3586);
and U5946 (N_5946,N_3924,N_4648);
nor U5947 (N_5947,N_3078,N_2505);
and U5948 (N_5948,N_4293,N_4002);
or U5949 (N_5949,N_4182,N_4505);
nor U5950 (N_5950,N_3314,N_3118);
nor U5951 (N_5951,N_2978,N_3274);
nand U5952 (N_5952,N_4788,N_3182);
xnor U5953 (N_5953,N_3598,N_4214);
nor U5954 (N_5954,N_4999,N_3137);
and U5955 (N_5955,N_3126,N_4937);
xnor U5956 (N_5956,N_3565,N_3382);
nand U5957 (N_5957,N_4476,N_3885);
nand U5958 (N_5958,N_3312,N_4210);
or U5959 (N_5959,N_3804,N_3044);
nand U5960 (N_5960,N_4133,N_4856);
and U5961 (N_5961,N_2669,N_4809);
nor U5962 (N_5962,N_3144,N_3889);
and U5963 (N_5963,N_4955,N_3160);
nand U5964 (N_5964,N_4379,N_3845);
or U5965 (N_5965,N_3285,N_4529);
nor U5966 (N_5966,N_3777,N_3952);
xnor U5967 (N_5967,N_3301,N_3901);
nand U5968 (N_5968,N_4513,N_2792);
and U5969 (N_5969,N_4641,N_2809);
xnor U5970 (N_5970,N_3528,N_3729);
and U5971 (N_5971,N_2936,N_3155);
or U5972 (N_5972,N_4849,N_4387);
xor U5973 (N_5973,N_3564,N_4551);
and U5974 (N_5974,N_3405,N_2706);
xor U5975 (N_5975,N_3928,N_3668);
xor U5976 (N_5976,N_4305,N_4137);
xor U5977 (N_5977,N_3754,N_4722);
nor U5978 (N_5978,N_4673,N_4801);
and U5979 (N_5979,N_4578,N_4415);
nor U5980 (N_5980,N_3855,N_4312);
or U5981 (N_5981,N_3192,N_4724);
or U5982 (N_5982,N_3035,N_3520);
nor U5983 (N_5983,N_4518,N_3479);
and U5984 (N_5984,N_4950,N_4527);
or U5985 (N_5985,N_4732,N_4432);
and U5986 (N_5986,N_2568,N_4823);
or U5987 (N_5987,N_3266,N_3242);
and U5988 (N_5988,N_3121,N_4731);
nor U5989 (N_5989,N_2709,N_3510);
nor U5990 (N_5990,N_2871,N_4854);
nor U5991 (N_5991,N_4337,N_4288);
nor U5992 (N_5992,N_4503,N_4974);
nand U5993 (N_5993,N_2744,N_4886);
and U5994 (N_5994,N_2661,N_3045);
nand U5995 (N_5995,N_4478,N_4175);
nor U5996 (N_5996,N_4725,N_4292);
or U5997 (N_5997,N_3463,N_3483);
nor U5998 (N_5998,N_2680,N_4875);
or U5999 (N_5999,N_2725,N_3354);
or U6000 (N_6000,N_3998,N_3073);
xor U6001 (N_6001,N_3969,N_4347);
or U6002 (N_6002,N_4629,N_3365);
nor U6003 (N_6003,N_3958,N_2990);
nor U6004 (N_6004,N_3193,N_3279);
nand U6005 (N_6005,N_4202,N_3022);
or U6006 (N_6006,N_4562,N_3169);
or U6007 (N_6007,N_3736,N_3540);
and U6008 (N_6008,N_3893,N_3436);
or U6009 (N_6009,N_3186,N_3224);
nor U6010 (N_6010,N_2681,N_4129);
nor U6011 (N_6011,N_2617,N_4390);
xor U6012 (N_6012,N_4832,N_3198);
and U6013 (N_6013,N_2575,N_3869);
and U6014 (N_6014,N_2982,N_4979);
and U6015 (N_6015,N_3109,N_4538);
and U6016 (N_6016,N_4256,N_3240);
nand U6017 (N_6017,N_4203,N_3571);
nor U6018 (N_6018,N_3201,N_4894);
nor U6019 (N_6019,N_4016,N_2552);
or U6020 (N_6020,N_3163,N_4110);
nor U6021 (N_6021,N_4480,N_3543);
or U6022 (N_6022,N_2683,N_4723);
nand U6023 (N_6023,N_2577,N_2603);
nor U6024 (N_6024,N_2645,N_4710);
nand U6025 (N_6025,N_4836,N_4905);
or U6026 (N_6026,N_2739,N_2740);
nand U6027 (N_6027,N_4536,N_3690);
and U6028 (N_6028,N_4628,N_2915);
nand U6029 (N_6029,N_3875,N_4514);
and U6030 (N_6030,N_3972,N_4994);
xnor U6031 (N_6031,N_2589,N_4656);
nand U6032 (N_6032,N_3041,N_4729);
nand U6033 (N_6033,N_4997,N_2928);
or U6034 (N_6034,N_2562,N_2831);
or U6035 (N_6035,N_2985,N_4635);
xor U6036 (N_6036,N_4664,N_4447);
xor U6037 (N_6037,N_3940,N_3649);
nand U6038 (N_6038,N_3271,N_4418);
nor U6039 (N_6039,N_3719,N_2941);
nor U6040 (N_6040,N_4283,N_2656);
nor U6041 (N_6041,N_2665,N_3162);
or U6042 (N_6042,N_4235,N_4741);
nor U6043 (N_6043,N_4301,N_2515);
or U6044 (N_6044,N_3962,N_4908);
nand U6045 (N_6045,N_3259,N_2926);
or U6046 (N_6046,N_4690,N_4973);
xnor U6047 (N_6047,N_2931,N_4153);
nand U6048 (N_6048,N_4570,N_4601);
and U6049 (N_6049,N_4517,N_4192);
or U6050 (N_6050,N_2797,N_3128);
or U6051 (N_6051,N_3211,N_3006);
nor U6052 (N_6052,N_2820,N_2901);
nor U6053 (N_6053,N_3315,N_4773);
nor U6054 (N_6054,N_4449,N_2997);
and U6055 (N_6055,N_4070,N_2550);
xnor U6056 (N_6056,N_3594,N_3190);
nand U6057 (N_6057,N_2833,N_2526);
xor U6058 (N_6058,N_2770,N_3870);
nor U6059 (N_6059,N_4431,N_2983);
nor U6060 (N_6060,N_3231,N_3395);
and U6061 (N_6061,N_3020,N_2517);
nand U6062 (N_6062,N_3060,N_3459);
xor U6063 (N_6063,N_4891,N_3730);
and U6064 (N_6064,N_4577,N_4851);
nand U6065 (N_6065,N_2968,N_4080);
or U6066 (N_6066,N_2986,N_4079);
xnor U6067 (N_6067,N_2560,N_4348);
nand U6068 (N_6068,N_2887,N_4633);
nand U6069 (N_6069,N_4792,N_3309);
and U6070 (N_6070,N_3532,N_3105);
or U6071 (N_6071,N_3424,N_4123);
and U6072 (N_6072,N_3304,N_2924);
and U6073 (N_6073,N_4285,N_4676);
nand U6074 (N_6074,N_4576,N_4295);
nor U6075 (N_6075,N_3987,N_2848);
or U6076 (N_6076,N_3165,N_3327);
nand U6077 (N_6077,N_3741,N_3085);
and U6078 (N_6078,N_4194,N_4691);
and U6079 (N_6079,N_4152,N_3926);
or U6080 (N_6080,N_3508,N_3589);
or U6081 (N_6081,N_2653,N_4496);
nor U6082 (N_6082,N_4215,N_4651);
nor U6083 (N_6083,N_4625,N_4467);
and U6084 (N_6084,N_3446,N_4661);
nand U6085 (N_6085,N_2675,N_3806);
or U6086 (N_6086,N_3590,N_3443);
or U6087 (N_6087,N_3646,N_3030);
or U6088 (N_6088,N_4705,N_4506);
or U6089 (N_6089,N_2840,N_4033);
nor U6090 (N_6090,N_4031,N_3675);
and U6091 (N_6091,N_3068,N_3562);
xnor U6092 (N_6092,N_4072,N_4566);
and U6093 (N_6093,N_3475,N_4914);
and U6094 (N_6094,N_3359,N_2916);
nor U6095 (N_6095,N_2793,N_4170);
and U6096 (N_6096,N_3156,N_4872);
nand U6097 (N_6097,N_3284,N_2572);
and U6098 (N_6098,N_3988,N_2959);
xnor U6099 (N_6099,N_3774,N_4770);
xor U6100 (N_6100,N_4669,N_4846);
nor U6101 (N_6101,N_2721,N_3054);
nand U6102 (N_6102,N_2853,N_4970);
nand U6103 (N_6103,N_3756,N_4368);
nor U6104 (N_6104,N_3585,N_4360);
nand U6105 (N_6105,N_3233,N_3944);
nor U6106 (N_6106,N_4340,N_4811);
or U6107 (N_6107,N_3195,N_4777);
nor U6108 (N_6108,N_2635,N_3011);
or U6109 (N_6109,N_3150,N_4892);
or U6110 (N_6110,N_3707,N_3642);
nand U6111 (N_6111,N_3579,N_4735);
or U6112 (N_6112,N_4821,N_4928);
nor U6113 (N_6113,N_4085,N_3431);
or U6114 (N_6114,N_2943,N_2549);
nor U6115 (N_6115,N_4971,N_2872);
nand U6116 (N_6116,N_3740,N_3997);
or U6117 (N_6117,N_2547,N_4150);
or U6118 (N_6118,N_3977,N_4018);
and U6119 (N_6119,N_2979,N_4190);
nor U6120 (N_6120,N_2664,N_4918);
and U6121 (N_6121,N_3180,N_4007);
and U6122 (N_6122,N_3143,N_3724);
and U6123 (N_6123,N_3819,N_4140);
or U6124 (N_6124,N_4932,N_2705);
and U6125 (N_6125,N_3385,N_3002);
and U6126 (N_6126,N_4654,N_4369);
nand U6127 (N_6127,N_3718,N_2756);
nand U6128 (N_6128,N_4926,N_4375);
or U6129 (N_6129,N_2747,N_3433);
and U6130 (N_6130,N_4895,N_2945);
or U6131 (N_6131,N_2838,N_4838);
and U6132 (N_6132,N_4961,N_3959);
and U6133 (N_6133,N_2595,N_4859);
nand U6134 (N_6134,N_3900,N_4643);
xor U6135 (N_6135,N_2662,N_3361);
or U6136 (N_6136,N_4176,N_2626);
nand U6137 (N_6137,N_3847,N_3455);
or U6138 (N_6138,N_3935,N_3088);
or U6139 (N_6139,N_4715,N_3641);
nor U6140 (N_6140,N_3302,N_4096);
and U6141 (N_6141,N_4270,N_4275);
nand U6142 (N_6142,N_4814,N_4157);
and U6143 (N_6143,N_4388,N_2843);
nand U6144 (N_6144,N_2804,N_3687);
or U6145 (N_6145,N_2722,N_3123);
nand U6146 (N_6146,N_2825,N_4906);
and U6147 (N_6147,N_2590,N_4038);
or U6148 (N_6148,N_4198,N_3775);
or U6149 (N_6149,N_2913,N_3630);
or U6150 (N_6150,N_4939,N_4600);
and U6151 (N_6151,N_4289,N_4888);
or U6152 (N_6152,N_2511,N_2758);
nand U6153 (N_6153,N_2796,N_4909);
nor U6154 (N_6154,N_4421,N_3629);
or U6155 (N_6155,N_4126,N_2689);
nor U6156 (N_6156,N_2741,N_4630);
and U6157 (N_6157,N_3978,N_3934);
nand U6158 (N_6158,N_3515,N_3973);
or U6159 (N_6159,N_3389,N_2832);
nor U6160 (N_6160,N_3568,N_3422);
nor U6161 (N_6161,N_2623,N_4504);
nor U6162 (N_6162,N_3949,N_3111);
nor U6163 (N_6163,N_3153,N_4232);
and U6164 (N_6164,N_2534,N_3680);
nor U6165 (N_6165,N_2521,N_3647);
nor U6166 (N_6166,N_3413,N_4511);
xnor U6167 (N_6167,N_2649,N_3664);
nor U6168 (N_6168,N_2693,N_3512);
or U6169 (N_6169,N_2863,N_4502);
nor U6170 (N_6170,N_4835,N_4244);
xnor U6171 (N_6171,N_3838,N_4454);
or U6172 (N_6172,N_3725,N_4848);
nor U6173 (N_6173,N_2690,N_3208);
xnor U6174 (N_6174,N_3158,N_4084);
or U6175 (N_6175,N_3699,N_3409);
or U6176 (N_6176,N_2734,N_4981);
or U6177 (N_6177,N_3768,N_4258);
and U6178 (N_6178,N_4099,N_3414);
or U6179 (N_6179,N_3744,N_2647);
nor U6180 (N_6180,N_3275,N_4652);
and U6181 (N_6181,N_3320,N_2847);
nor U6182 (N_6182,N_2587,N_3511);
nand U6183 (N_6183,N_2650,N_3210);
nand U6184 (N_6184,N_4719,N_4087);
nand U6185 (N_6185,N_3415,N_3380);
and U6186 (N_6186,N_4409,N_3017);
or U6187 (N_6187,N_4799,N_4820);
or U6188 (N_6188,N_4042,N_3849);
xor U6189 (N_6189,N_3815,N_4058);
or U6190 (N_6190,N_4092,N_2620);
xor U6191 (N_6191,N_2895,N_4603);
nor U6192 (N_6192,N_3533,N_2601);
nor U6193 (N_6193,N_3982,N_4917);
or U6194 (N_6194,N_3614,N_4786);
or U6195 (N_6195,N_4105,N_4978);
nand U6196 (N_6196,N_3196,N_4957);
nand U6197 (N_6197,N_2909,N_4029);
or U6198 (N_6198,N_4445,N_3789);
and U6199 (N_6199,N_4248,N_4798);
or U6200 (N_6200,N_3004,N_2614);
nor U6201 (N_6201,N_4155,N_4132);
or U6202 (N_6202,N_3064,N_4563);
or U6203 (N_6203,N_2802,N_3281);
nand U6204 (N_6204,N_3739,N_3968);
xor U6205 (N_6205,N_4290,N_4264);
nand U6206 (N_6206,N_4267,N_4606);
or U6207 (N_6207,N_3993,N_3731);
nand U6208 (N_6208,N_3452,N_4593);
xnor U6209 (N_6209,N_4154,N_4461);
and U6210 (N_6210,N_3247,N_4568);
nand U6211 (N_6211,N_3056,N_3669);
nor U6212 (N_6212,N_2641,N_3108);
nand U6213 (N_6213,N_4307,N_3264);
or U6214 (N_6214,N_3490,N_4840);
or U6215 (N_6215,N_2794,N_4027);
nor U6216 (N_6216,N_2506,N_4488);
nand U6217 (N_6217,N_3401,N_4824);
or U6218 (N_6218,N_3569,N_4780);
nand U6219 (N_6219,N_4442,N_4796);
nand U6220 (N_6220,N_4802,N_3746);
and U6221 (N_6221,N_4744,N_3965);
nand U6222 (N_6222,N_3176,N_4934);
nand U6223 (N_6223,N_4466,N_4355);
and U6224 (N_6224,N_3001,N_4546);
or U6225 (N_6225,N_4636,N_4218);
xnor U6226 (N_6226,N_4807,N_4074);
and U6227 (N_6227,N_3381,N_4117);
or U6228 (N_6228,N_4785,N_3704);
nand U6229 (N_6229,N_4733,N_4420);
or U6230 (N_6230,N_4000,N_3920);
or U6231 (N_6231,N_4597,N_2775);
nor U6232 (N_6232,N_4666,N_3941);
or U6233 (N_6233,N_3488,N_4260);
or U6234 (N_6234,N_4352,N_2890);
nand U6235 (N_6235,N_3814,N_3667);
nor U6236 (N_6236,N_4201,N_3500);
nor U6237 (N_6237,N_4269,N_4992);
nor U6238 (N_6238,N_2790,N_2674);
xor U6239 (N_6239,N_4826,N_4500);
and U6240 (N_6240,N_4426,N_4761);
and U6241 (N_6241,N_3722,N_3766);
xnor U6242 (N_6242,N_3995,N_3219);
or U6243 (N_6243,N_3863,N_4685);
or U6244 (N_6244,N_4993,N_4998);
nand U6245 (N_6245,N_4876,N_4567);
or U6246 (N_6246,N_4325,N_4549);
or U6247 (N_6247,N_4139,N_4778);
nor U6248 (N_6248,N_3238,N_4433);
and U6249 (N_6249,N_3716,N_4142);
or U6250 (N_6250,N_4014,N_2733);
nand U6251 (N_6251,N_4911,N_4080);
nor U6252 (N_6252,N_2813,N_4002);
nor U6253 (N_6253,N_4768,N_3979);
nand U6254 (N_6254,N_3962,N_3065);
nor U6255 (N_6255,N_4177,N_4483);
nor U6256 (N_6256,N_4437,N_4138);
or U6257 (N_6257,N_2677,N_3395);
nor U6258 (N_6258,N_4628,N_3245);
or U6259 (N_6259,N_3961,N_4728);
xnor U6260 (N_6260,N_4489,N_4584);
xnor U6261 (N_6261,N_3793,N_3008);
or U6262 (N_6262,N_4467,N_3795);
xor U6263 (N_6263,N_3080,N_3949);
and U6264 (N_6264,N_4256,N_3607);
xor U6265 (N_6265,N_4581,N_2678);
nor U6266 (N_6266,N_4367,N_4765);
or U6267 (N_6267,N_4420,N_3119);
nand U6268 (N_6268,N_3197,N_3499);
and U6269 (N_6269,N_4724,N_2597);
and U6270 (N_6270,N_2891,N_4476);
or U6271 (N_6271,N_3935,N_2906);
nand U6272 (N_6272,N_3120,N_3823);
nand U6273 (N_6273,N_4652,N_2802);
or U6274 (N_6274,N_2511,N_3893);
nor U6275 (N_6275,N_4287,N_3048);
xor U6276 (N_6276,N_3690,N_3947);
nand U6277 (N_6277,N_3513,N_4977);
and U6278 (N_6278,N_4358,N_2990);
nor U6279 (N_6279,N_3894,N_3241);
and U6280 (N_6280,N_3767,N_4629);
nand U6281 (N_6281,N_4397,N_3986);
or U6282 (N_6282,N_4695,N_3985);
xnor U6283 (N_6283,N_3322,N_4986);
xor U6284 (N_6284,N_3851,N_2709);
nand U6285 (N_6285,N_4983,N_4014);
nand U6286 (N_6286,N_3411,N_3513);
xor U6287 (N_6287,N_4910,N_3382);
nor U6288 (N_6288,N_3103,N_2792);
or U6289 (N_6289,N_4720,N_3550);
or U6290 (N_6290,N_4482,N_3400);
nand U6291 (N_6291,N_4324,N_3561);
xor U6292 (N_6292,N_3511,N_4328);
and U6293 (N_6293,N_4576,N_3946);
nand U6294 (N_6294,N_3076,N_2798);
and U6295 (N_6295,N_2888,N_4603);
nor U6296 (N_6296,N_2660,N_4440);
and U6297 (N_6297,N_3110,N_4954);
xor U6298 (N_6298,N_4585,N_4101);
or U6299 (N_6299,N_2827,N_4369);
xor U6300 (N_6300,N_2997,N_3560);
nor U6301 (N_6301,N_3207,N_4982);
nor U6302 (N_6302,N_4368,N_2915);
or U6303 (N_6303,N_3183,N_3560);
and U6304 (N_6304,N_4001,N_4718);
or U6305 (N_6305,N_4234,N_3105);
or U6306 (N_6306,N_3233,N_3828);
or U6307 (N_6307,N_3879,N_4423);
or U6308 (N_6308,N_3512,N_3329);
or U6309 (N_6309,N_4467,N_2888);
xor U6310 (N_6310,N_4822,N_3258);
nand U6311 (N_6311,N_3809,N_4128);
nand U6312 (N_6312,N_4101,N_2788);
nor U6313 (N_6313,N_4257,N_4127);
xor U6314 (N_6314,N_4819,N_3242);
nand U6315 (N_6315,N_4107,N_4204);
xor U6316 (N_6316,N_3223,N_2676);
nor U6317 (N_6317,N_3893,N_4904);
and U6318 (N_6318,N_3787,N_3904);
xor U6319 (N_6319,N_4793,N_4520);
nor U6320 (N_6320,N_4404,N_3219);
or U6321 (N_6321,N_4545,N_3697);
and U6322 (N_6322,N_4373,N_4723);
and U6323 (N_6323,N_2733,N_2704);
or U6324 (N_6324,N_4310,N_3839);
or U6325 (N_6325,N_3628,N_2649);
or U6326 (N_6326,N_4252,N_2779);
xnor U6327 (N_6327,N_4359,N_4081);
nor U6328 (N_6328,N_4781,N_3962);
or U6329 (N_6329,N_3852,N_3833);
xor U6330 (N_6330,N_3100,N_3599);
or U6331 (N_6331,N_3261,N_2614);
nor U6332 (N_6332,N_2600,N_4326);
or U6333 (N_6333,N_4741,N_4276);
xnor U6334 (N_6334,N_2893,N_2674);
nand U6335 (N_6335,N_4142,N_4895);
nand U6336 (N_6336,N_4864,N_3012);
nor U6337 (N_6337,N_3699,N_3617);
nand U6338 (N_6338,N_3733,N_4427);
and U6339 (N_6339,N_4215,N_4816);
nor U6340 (N_6340,N_4404,N_3064);
nand U6341 (N_6341,N_3548,N_4767);
nor U6342 (N_6342,N_4820,N_3634);
and U6343 (N_6343,N_2762,N_2710);
or U6344 (N_6344,N_4573,N_3096);
nand U6345 (N_6345,N_2876,N_2825);
nor U6346 (N_6346,N_4038,N_3468);
and U6347 (N_6347,N_3102,N_4647);
nand U6348 (N_6348,N_3026,N_2790);
or U6349 (N_6349,N_4861,N_4320);
nor U6350 (N_6350,N_3083,N_3100);
nor U6351 (N_6351,N_3841,N_4368);
nand U6352 (N_6352,N_3067,N_3111);
xor U6353 (N_6353,N_3050,N_2537);
nor U6354 (N_6354,N_4048,N_3714);
and U6355 (N_6355,N_4084,N_3773);
and U6356 (N_6356,N_3776,N_3245);
nor U6357 (N_6357,N_2976,N_4924);
xnor U6358 (N_6358,N_4021,N_3812);
xnor U6359 (N_6359,N_2764,N_2964);
nand U6360 (N_6360,N_4788,N_3017);
or U6361 (N_6361,N_2691,N_4892);
nor U6362 (N_6362,N_2705,N_4592);
nand U6363 (N_6363,N_4523,N_3028);
nor U6364 (N_6364,N_4984,N_2734);
and U6365 (N_6365,N_3010,N_4748);
nand U6366 (N_6366,N_4200,N_3344);
xor U6367 (N_6367,N_3945,N_2630);
or U6368 (N_6368,N_3720,N_3143);
nand U6369 (N_6369,N_4873,N_4343);
and U6370 (N_6370,N_3264,N_2536);
or U6371 (N_6371,N_3861,N_3139);
nand U6372 (N_6372,N_3140,N_3603);
or U6373 (N_6373,N_4922,N_3176);
nand U6374 (N_6374,N_3586,N_3310);
or U6375 (N_6375,N_4008,N_4570);
nor U6376 (N_6376,N_3377,N_4671);
and U6377 (N_6377,N_3700,N_3544);
nor U6378 (N_6378,N_3595,N_4329);
or U6379 (N_6379,N_2577,N_2745);
or U6380 (N_6380,N_4624,N_3207);
and U6381 (N_6381,N_4576,N_4941);
nor U6382 (N_6382,N_4253,N_2807);
xor U6383 (N_6383,N_2637,N_3197);
nand U6384 (N_6384,N_4648,N_3746);
or U6385 (N_6385,N_3290,N_2606);
or U6386 (N_6386,N_4293,N_4744);
and U6387 (N_6387,N_4833,N_2574);
and U6388 (N_6388,N_4740,N_3190);
xnor U6389 (N_6389,N_3328,N_3214);
and U6390 (N_6390,N_4138,N_3260);
nand U6391 (N_6391,N_3365,N_2828);
nand U6392 (N_6392,N_4023,N_3216);
nor U6393 (N_6393,N_4581,N_4791);
nor U6394 (N_6394,N_4981,N_4754);
and U6395 (N_6395,N_2532,N_2624);
nand U6396 (N_6396,N_3146,N_4189);
or U6397 (N_6397,N_4104,N_2678);
nor U6398 (N_6398,N_3187,N_3436);
xnor U6399 (N_6399,N_4261,N_3292);
and U6400 (N_6400,N_3277,N_3432);
nor U6401 (N_6401,N_4163,N_4288);
nor U6402 (N_6402,N_3746,N_3093);
and U6403 (N_6403,N_3958,N_4184);
or U6404 (N_6404,N_3184,N_4294);
nor U6405 (N_6405,N_3117,N_3290);
or U6406 (N_6406,N_4944,N_3367);
or U6407 (N_6407,N_4887,N_3321);
nand U6408 (N_6408,N_3782,N_2986);
nor U6409 (N_6409,N_2974,N_3608);
and U6410 (N_6410,N_3613,N_4130);
nor U6411 (N_6411,N_3869,N_4683);
and U6412 (N_6412,N_4354,N_3456);
nor U6413 (N_6413,N_4499,N_4702);
or U6414 (N_6414,N_3104,N_4042);
or U6415 (N_6415,N_3874,N_3750);
nand U6416 (N_6416,N_3155,N_2555);
or U6417 (N_6417,N_2662,N_4927);
or U6418 (N_6418,N_4921,N_4390);
or U6419 (N_6419,N_3241,N_4094);
nand U6420 (N_6420,N_2592,N_4021);
nor U6421 (N_6421,N_3032,N_3523);
nand U6422 (N_6422,N_2871,N_4766);
xnor U6423 (N_6423,N_4340,N_3369);
xnor U6424 (N_6424,N_3036,N_3054);
nor U6425 (N_6425,N_3281,N_3252);
or U6426 (N_6426,N_3470,N_4603);
or U6427 (N_6427,N_3936,N_3400);
and U6428 (N_6428,N_4049,N_3128);
or U6429 (N_6429,N_3950,N_2799);
or U6430 (N_6430,N_4675,N_3029);
nand U6431 (N_6431,N_3921,N_4558);
or U6432 (N_6432,N_4458,N_4604);
nor U6433 (N_6433,N_4025,N_4863);
and U6434 (N_6434,N_4407,N_3602);
nor U6435 (N_6435,N_2586,N_3295);
nor U6436 (N_6436,N_4698,N_2863);
nor U6437 (N_6437,N_2531,N_4156);
or U6438 (N_6438,N_4389,N_4885);
nor U6439 (N_6439,N_3331,N_4352);
nor U6440 (N_6440,N_4574,N_3175);
and U6441 (N_6441,N_3335,N_2657);
or U6442 (N_6442,N_4397,N_3680);
and U6443 (N_6443,N_4929,N_4834);
or U6444 (N_6444,N_3209,N_4841);
and U6445 (N_6445,N_2630,N_3611);
nor U6446 (N_6446,N_2995,N_3403);
nand U6447 (N_6447,N_2894,N_4228);
xnor U6448 (N_6448,N_4962,N_2693);
or U6449 (N_6449,N_4139,N_3803);
or U6450 (N_6450,N_4082,N_4162);
or U6451 (N_6451,N_3855,N_4032);
xor U6452 (N_6452,N_2929,N_2630);
nand U6453 (N_6453,N_2814,N_4714);
nand U6454 (N_6454,N_3481,N_2861);
nand U6455 (N_6455,N_3252,N_3438);
nand U6456 (N_6456,N_4096,N_3847);
nand U6457 (N_6457,N_3167,N_4607);
and U6458 (N_6458,N_4833,N_3921);
or U6459 (N_6459,N_3687,N_2639);
nand U6460 (N_6460,N_3434,N_4407);
nand U6461 (N_6461,N_3522,N_3548);
and U6462 (N_6462,N_3080,N_3853);
and U6463 (N_6463,N_4799,N_4222);
and U6464 (N_6464,N_4630,N_3757);
xnor U6465 (N_6465,N_3447,N_2913);
nand U6466 (N_6466,N_3031,N_2801);
and U6467 (N_6467,N_3278,N_4220);
or U6468 (N_6468,N_3488,N_4693);
or U6469 (N_6469,N_2869,N_3086);
and U6470 (N_6470,N_4327,N_3822);
nor U6471 (N_6471,N_3232,N_3621);
or U6472 (N_6472,N_2732,N_3266);
and U6473 (N_6473,N_3305,N_4851);
xor U6474 (N_6474,N_3948,N_3303);
and U6475 (N_6475,N_3952,N_4328);
nand U6476 (N_6476,N_2931,N_4622);
or U6477 (N_6477,N_3336,N_2580);
nor U6478 (N_6478,N_3592,N_4972);
nor U6479 (N_6479,N_3215,N_3018);
xnor U6480 (N_6480,N_4886,N_3164);
or U6481 (N_6481,N_4317,N_3466);
nor U6482 (N_6482,N_4780,N_3777);
nor U6483 (N_6483,N_4503,N_4961);
and U6484 (N_6484,N_3165,N_4987);
nand U6485 (N_6485,N_4943,N_4759);
and U6486 (N_6486,N_3984,N_4416);
nand U6487 (N_6487,N_4386,N_4455);
nor U6488 (N_6488,N_4168,N_3971);
and U6489 (N_6489,N_3524,N_2866);
or U6490 (N_6490,N_3249,N_4716);
and U6491 (N_6491,N_2524,N_4962);
xnor U6492 (N_6492,N_4687,N_3102);
nand U6493 (N_6493,N_4035,N_3865);
and U6494 (N_6494,N_4952,N_4298);
or U6495 (N_6495,N_3789,N_3270);
and U6496 (N_6496,N_2711,N_3735);
nand U6497 (N_6497,N_4569,N_4916);
nor U6498 (N_6498,N_3905,N_4010);
or U6499 (N_6499,N_3801,N_3626);
or U6500 (N_6500,N_3562,N_4464);
or U6501 (N_6501,N_2830,N_3667);
nor U6502 (N_6502,N_4676,N_3750);
and U6503 (N_6503,N_3712,N_3487);
nand U6504 (N_6504,N_3577,N_4474);
nor U6505 (N_6505,N_3872,N_3881);
or U6506 (N_6506,N_3530,N_3889);
nor U6507 (N_6507,N_4394,N_2708);
or U6508 (N_6508,N_3123,N_3199);
xnor U6509 (N_6509,N_3325,N_2711);
nor U6510 (N_6510,N_4517,N_3065);
or U6511 (N_6511,N_4098,N_3420);
nor U6512 (N_6512,N_4159,N_2925);
or U6513 (N_6513,N_4660,N_3700);
or U6514 (N_6514,N_4363,N_4464);
nor U6515 (N_6515,N_2623,N_4903);
xnor U6516 (N_6516,N_2769,N_3506);
xnor U6517 (N_6517,N_3426,N_4540);
nand U6518 (N_6518,N_2631,N_4521);
nor U6519 (N_6519,N_3230,N_3437);
nand U6520 (N_6520,N_4275,N_2715);
and U6521 (N_6521,N_2529,N_2742);
xnor U6522 (N_6522,N_3172,N_4570);
nor U6523 (N_6523,N_4194,N_3671);
nand U6524 (N_6524,N_4266,N_2638);
nor U6525 (N_6525,N_3373,N_3335);
nand U6526 (N_6526,N_4600,N_2634);
nand U6527 (N_6527,N_4101,N_3161);
and U6528 (N_6528,N_4371,N_4494);
and U6529 (N_6529,N_3631,N_3003);
nand U6530 (N_6530,N_2748,N_2681);
and U6531 (N_6531,N_3196,N_4129);
xor U6532 (N_6532,N_2754,N_3683);
nor U6533 (N_6533,N_2786,N_3803);
and U6534 (N_6534,N_4644,N_2885);
and U6535 (N_6535,N_3609,N_4108);
and U6536 (N_6536,N_3248,N_3188);
nor U6537 (N_6537,N_3346,N_2989);
or U6538 (N_6538,N_3614,N_4959);
nand U6539 (N_6539,N_2639,N_4532);
nand U6540 (N_6540,N_3660,N_3665);
xor U6541 (N_6541,N_4889,N_3752);
xnor U6542 (N_6542,N_4144,N_2895);
nand U6543 (N_6543,N_3444,N_2665);
nor U6544 (N_6544,N_4096,N_3672);
nand U6545 (N_6545,N_4166,N_4135);
nor U6546 (N_6546,N_3391,N_3943);
xnor U6547 (N_6547,N_4370,N_3687);
nand U6548 (N_6548,N_4212,N_3381);
and U6549 (N_6549,N_3449,N_3169);
or U6550 (N_6550,N_3811,N_3813);
or U6551 (N_6551,N_4930,N_3784);
and U6552 (N_6552,N_2935,N_4588);
nor U6553 (N_6553,N_3409,N_4343);
and U6554 (N_6554,N_3977,N_2519);
and U6555 (N_6555,N_4882,N_4670);
or U6556 (N_6556,N_4466,N_4484);
nand U6557 (N_6557,N_3905,N_4184);
or U6558 (N_6558,N_4306,N_4497);
nand U6559 (N_6559,N_2593,N_3323);
xor U6560 (N_6560,N_4487,N_3366);
and U6561 (N_6561,N_2801,N_4087);
nand U6562 (N_6562,N_3754,N_4738);
or U6563 (N_6563,N_2934,N_2731);
and U6564 (N_6564,N_4333,N_3939);
nand U6565 (N_6565,N_4131,N_2592);
nand U6566 (N_6566,N_4565,N_2568);
or U6567 (N_6567,N_3166,N_4349);
nor U6568 (N_6568,N_4129,N_4793);
nand U6569 (N_6569,N_4010,N_2845);
nor U6570 (N_6570,N_4072,N_4248);
xnor U6571 (N_6571,N_2878,N_4536);
nor U6572 (N_6572,N_2802,N_4302);
or U6573 (N_6573,N_3958,N_3631);
and U6574 (N_6574,N_4287,N_2912);
or U6575 (N_6575,N_3505,N_3157);
and U6576 (N_6576,N_3795,N_3895);
xnor U6577 (N_6577,N_4101,N_4132);
nand U6578 (N_6578,N_4598,N_3924);
and U6579 (N_6579,N_4120,N_3542);
or U6580 (N_6580,N_4753,N_3950);
nor U6581 (N_6581,N_4914,N_3801);
and U6582 (N_6582,N_4836,N_3797);
nand U6583 (N_6583,N_2772,N_3223);
nor U6584 (N_6584,N_2828,N_3846);
nand U6585 (N_6585,N_3884,N_3058);
xor U6586 (N_6586,N_3673,N_4165);
or U6587 (N_6587,N_3275,N_3956);
xnor U6588 (N_6588,N_2661,N_4511);
or U6589 (N_6589,N_2756,N_4614);
or U6590 (N_6590,N_3248,N_3317);
nand U6591 (N_6591,N_2515,N_2729);
nor U6592 (N_6592,N_3252,N_3121);
or U6593 (N_6593,N_2945,N_3572);
or U6594 (N_6594,N_4396,N_3364);
and U6595 (N_6595,N_4322,N_3109);
or U6596 (N_6596,N_3133,N_2773);
or U6597 (N_6597,N_4964,N_3472);
nor U6598 (N_6598,N_4253,N_4309);
and U6599 (N_6599,N_3336,N_3346);
nand U6600 (N_6600,N_3619,N_3080);
nand U6601 (N_6601,N_3386,N_2757);
and U6602 (N_6602,N_3255,N_4716);
or U6603 (N_6603,N_3098,N_2722);
nor U6604 (N_6604,N_4913,N_2831);
nand U6605 (N_6605,N_3921,N_3732);
or U6606 (N_6606,N_2834,N_3288);
and U6607 (N_6607,N_4297,N_3632);
and U6608 (N_6608,N_2721,N_4066);
and U6609 (N_6609,N_4379,N_3004);
or U6610 (N_6610,N_3619,N_4961);
nand U6611 (N_6611,N_3417,N_3018);
nand U6612 (N_6612,N_4292,N_4377);
or U6613 (N_6613,N_4382,N_2987);
nor U6614 (N_6614,N_2569,N_3571);
or U6615 (N_6615,N_3832,N_3143);
and U6616 (N_6616,N_4908,N_3751);
or U6617 (N_6617,N_4890,N_4635);
xor U6618 (N_6618,N_4555,N_4275);
and U6619 (N_6619,N_4709,N_3862);
nor U6620 (N_6620,N_4801,N_2843);
or U6621 (N_6621,N_4910,N_4630);
nand U6622 (N_6622,N_2529,N_4391);
nand U6623 (N_6623,N_4964,N_3405);
and U6624 (N_6624,N_3974,N_4589);
or U6625 (N_6625,N_3480,N_2681);
nor U6626 (N_6626,N_3699,N_4827);
nand U6627 (N_6627,N_4213,N_4409);
nand U6628 (N_6628,N_3168,N_3529);
and U6629 (N_6629,N_4121,N_4576);
xor U6630 (N_6630,N_3890,N_4040);
nand U6631 (N_6631,N_2843,N_3463);
nor U6632 (N_6632,N_4173,N_4336);
or U6633 (N_6633,N_4674,N_3035);
or U6634 (N_6634,N_3704,N_4984);
or U6635 (N_6635,N_3205,N_4010);
nand U6636 (N_6636,N_4894,N_2787);
and U6637 (N_6637,N_3764,N_3342);
and U6638 (N_6638,N_3980,N_2548);
nor U6639 (N_6639,N_4576,N_4041);
and U6640 (N_6640,N_3588,N_4460);
and U6641 (N_6641,N_2554,N_3075);
nand U6642 (N_6642,N_4187,N_4387);
nand U6643 (N_6643,N_4382,N_3558);
nand U6644 (N_6644,N_3067,N_4959);
nand U6645 (N_6645,N_4301,N_3405);
nor U6646 (N_6646,N_4379,N_4789);
and U6647 (N_6647,N_4534,N_4000);
nand U6648 (N_6648,N_4155,N_3862);
xnor U6649 (N_6649,N_4127,N_3268);
nand U6650 (N_6650,N_2818,N_3767);
nor U6651 (N_6651,N_4168,N_3583);
and U6652 (N_6652,N_3335,N_4942);
nand U6653 (N_6653,N_3584,N_3838);
nor U6654 (N_6654,N_4492,N_4654);
nand U6655 (N_6655,N_3546,N_2575);
nor U6656 (N_6656,N_4574,N_4386);
and U6657 (N_6657,N_3798,N_3687);
and U6658 (N_6658,N_3091,N_4721);
or U6659 (N_6659,N_3157,N_4984);
and U6660 (N_6660,N_2774,N_3648);
nor U6661 (N_6661,N_2590,N_3008);
or U6662 (N_6662,N_3257,N_4116);
or U6663 (N_6663,N_4240,N_3406);
nor U6664 (N_6664,N_4089,N_3198);
nand U6665 (N_6665,N_4304,N_4141);
xor U6666 (N_6666,N_4351,N_4935);
nand U6667 (N_6667,N_4552,N_2753);
and U6668 (N_6668,N_2979,N_3313);
xnor U6669 (N_6669,N_3756,N_3207);
and U6670 (N_6670,N_4776,N_2724);
nand U6671 (N_6671,N_2973,N_2733);
nand U6672 (N_6672,N_4582,N_3332);
nor U6673 (N_6673,N_4865,N_4508);
nor U6674 (N_6674,N_3954,N_3808);
and U6675 (N_6675,N_2583,N_3655);
or U6676 (N_6676,N_3684,N_4767);
and U6677 (N_6677,N_2758,N_3028);
nor U6678 (N_6678,N_4832,N_4464);
nand U6679 (N_6679,N_2582,N_4806);
nand U6680 (N_6680,N_2797,N_2757);
and U6681 (N_6681,N_3447,N_3380);
nor U6682 (N_6682,N_3404,N_2535);
or U6683 (N_6683,N_4140,N_3146);
and U6684 (N_6684,N_2557,N_3813);
and U6685 (N_6685,N_3703,N_4168);
nand U6686 (N_6686,N_4419,N_4442);
or U6687 (N_6687,N_3060,N_4777);
and U6688 (N_6688,N_4186,N_2823);
nand U6689 (N_6689,N_2780,N_3472);
and U6690 (N_6690,N_4526,N_4390);
or U6691 (N_6691,N_4639,N_3067);
nor U6692 (N_6692,N_4501,N_2985);
xor U6693 (N_6693,N_3740,N_2755);
nor U6694 (N_6694,N_4018,N_3331);
nor U6695 (N_6695,N_3357,N_3374);
and U6696 (N_6696,N_3068,N_4463);
and U6697 (N_6697,N_4477,N_3586);
xnor U6698 (N_6698,N_3851,N_3863);
and U6699 (N_6699,N_3104,N_4750);
nor U6700 (N_6700,N_3086,N_2868);
nand U6701 (N_6701,N_4654,N_3335);
xnor U6702 (N_6702,N_3094,N_3970);
and U6703 (N_6703,N_4400,N_4908);
nand U6704 (N_6704,N_4744,N_4406);
nor U6705 (N_6705,N_3080,N_3656);
and U6706 (N_6706,N_3930,N_3273);
nor U6707 (N_6707,N_3542,N_4143);
or U6708 (N_6708,N_2701,N_3006);
and U6709 (N_6709,N_4757,N_2969);
and U6710 (N_6710,N_3872,N_3526);
or U6711 (N_6711,N_4339,N_2636);
xnor U6712 (N_6712,N_2632,N_4991);
nand U6713 (N_6713,N_4195,N_4936);
nor U6714 (N_6714,N_3682,N_4122);
nor U6715 (N_6715,N_3189,N_3683);
or U6716 (N_6716,N_4372,N_2886);
nand U6717 (N_6717,N_4231,N_2863);
nor U6718 (N_6718,N_3842,N_3497);
and U6719 (N_6719,N_3733,N_2727);
nand U6720 (N_6720,N_3381,N_2517);
nor U6721 (N_6721,N_3967,N_4792);
and U6722 (N_6722,N_3720,N_4286);
or U6723 (N_6723,N_4653,N_4337);
nand U6724 (N_6724,N_4010,N_3375);
or U6725 (N_6725,N_3018,N_2668);
nor U6726 (N_6726,N_4002,N_3021);
nor U6727 (N_6727,N_4581,N_2738);
or U6728 (N_6728,N_2741,N_4837);
nand U6729 (N_6729,N_2847,N_4390);
and U6730 (N_6730,N_3679,N_4945);
nor U6731 (N_6731,N_3292,N_3774);
nor U6732 (N_6732,N_4219,N_2627);
nor U6733 (N_6733,N_3018,N_2608);
or U6734 (N_6734,N_4494,N_3938);
or U6735 (N_6735,N_3412,N_4063);
or U6736 (N_6736,N_4625,N_3216);
nand U6737 (N_6737,N_4014,N_4664);
nand U6738 (N_6738,N_4604,N_4449);
and U6739 (N_6739,N_4895,N_3677);
nand U6740 (N_6740,N_4242,N_2763);
or U6741 (N_6741,N_2895,N_4536);
nand U6742 (N_6742,N_3982,N_4034);
nand U6743 (N_6743,N_4344,N_2592);
and U6744 (N_6744,N_3195,N_4574);
nand U6745 (N_6745,N_2680,N_2729);
and U6746 (N_6746,N_3137,N_3919);
and U6747 (N_6747,N_3530,N_4456);
or U6748 (N_6748,N_3546,N_2505);
xnor U6749 (N_6749,N_4342,N_3064);
or U6750 (N_6750,N_3324,N_2565);
or U6751 (N_6751,N_3176,N_3632);
or U6752 (N_6752,N_2914,N_3640);
nand U6753 (N_6753,N_3171,N_2671);
and U6754 (N_6754,N_3437,N_3855);
or U6755 (N_6755,N_2564,N_4477);
nor U6756 (N_6756,N_3505,N_4494);
or U6757 (N_6757,N_3031,N_4100);
and U6758 (N_6758,N_2563,N_2871);
and U6759 (N_6759,N_3205,N_3127);
nor U6760 (N_6760,N_4015,N_4731);
nor U6761 (N_6761,N_2650,N_2880);
nand U6762 (N_6762,N_3582,N_3076);
nand U6763 (N_6763,N_3184,N_3625);
nand U6764 (N_6764,N_4066,N_4945);
nand U6765 (N_6765,N_2951,N_4306);
or U6766 (N_6766,N_4595,N_4690);
xor U6767 (N_6767,N_2632,N_2965);
and U6768 (N_6768,N_4621,N_4801);
or U6769 (N_6769,N_3537,N_4766);
nand U6770 (N_6770,N_4511,N_3772);
and U6771 (N_6771,N_3210,N_3572);
and U6772 (N_6772,N_4124,N_2934);
or U6773 (N_6773,N_4650,N_4107);
nor U6774 (N_6774,N_3517,N_4110);
xnor U6775 (N_6775,N_3287,N_3465);
and U6776 (N_6776,N_4705,N_2908);
nor U6777 (N_6777,N_4940,N_2950);
nor U6778 (N_6778,N_2624,N_3595);
and U6779 (N_6779,N_3070,N_3544);
nand U6780 (N_6780,N_3119,N_4838);
nand U6781 (N_6781,N_4135,N_3736);
nor U6782 (N_6782,N_4912,N_4688);
nor U6783 (N_6783,N_4274,N_3676);
xor U6784 (N_6784,N_3998,N_4743);
nand U6785 (N_6785,N_2987,N_2680);
or U6786 (N_6786,N_4612,N_2834);
nor U6787 (N_6787,N_3308,N_4980);
nor U6788 (N_6788,N_4468,N_3753);
nor U6789 (N_6789,N_2964,N_3350);
nand U6790 (N_6790,N_2966,N_4633);
and U6791 (N_6791,N_3888,N_4453);
or U6792 (N_6792,N_2784,N_3389);
nand U6793 (N_6793,N_2565,N_4321);
and U6794 (N_6794,N_4961,N_2503);
or U6795 (N_6795,N_3725,N_3254);
xor U6796 (N_6796,N_3861,N_4171);
or U6797 (N_6797,N_4236,N_3178);
and U6798 (N_6798,N_3336,N_2621);
nand U6799 (N_6799,N_2678,N_4301);
nand U6800 (N_6800,N_2739,N_3319);
and U6801 (N_6801,N_4932,N_3869);
and U6802 (N_6802,N_3291,N_2591);
or U6803 (N_6803,N_3565,N_4275);
or U6804 (N_6804,N_3569,N_3730);
or U6805 (N_6805,N_3252,N_3495);
xor U6806 (N_6806,N_4749,N_4470);
nor U6807 (N_6807,N_4664,N_4807);
and U6808 (N_6808,N_3225,N_3849);
nand U6809 (N_6809,N_4672,N_3458);
nor U6810 (N_6810,N_4147,N_4551);
nor U6811 (N_6811,N_4503,N_4360);
xnor U6812 (N_6812,N_3259,N_4831);
nand U6813 (N_6813,N_3613,N_3411);
nor U6814 (N_6814,N_4285,N_3216);
nor U6815 (N_6815,N_3366,N_4462);
nand U6816 (N_6816,N_3467,N_3277);
nand U6817 (N_6817,N_3995,N_4546);
nand U6818 (N_6818,N_3469,N_4684);
xor U6819 (N_6819,N_2894,N_4474);
and U6820 (N_6820,N_4152,N_3870);
or U6821 (N_6821,N_3860,N_4771);
xnor U6822 (N_6822,N_2501,N_4719);
nor U6823 (N_6823,N_2649,N_3926);
or U6824 (N_6824,N_3898,N_3399);
nor U6825 (N_6825,N_2918,N_4992);
xnor U6826 (N_6826,N_4672,N_4919);
or U6827 (N_6827,N_3497,N_3667);
nand U6828 (N_6828,N_3554,N_3342);
nand U6829 (N_6829,N_3844,N_3562);
or U6830 (N_6830,N_2640,N_3266);
nor U6831 (N_6831,N_3878,N_2762);
and U6832 (N_6832,N_3621,N_3529);
nand U6833 (N_6833,N_3532,N_4012);
or U6834 (N_6834,N_4745,N_4495);
xnor U6835 (N_6835,N_4971,N_3681);
or U6836 (N_6836,N_2872,N_4037);
and U6837 (N_6837,N_3277,N_4916);
and U6838 (N_6838,N_3767,N_4192);
nor U6839 (N_6839,N_3386,N_4655);
nand U6840 (N_6840,N_4081,N_4048);
and U6841 (N_6841,N_4194,N_3337);
xnor U6842 (N_6842,N_3017,N_2660);
or U6843 (N_6843,N_3138,N_4176);
nor U6844 (N_6844,N_3926,N_3500);
or U6845 (N_6845,N_3071,N_3095);
nand U6846 (N_6846,N_3993,N_2741);
and U6847 (N_6847,N_3673,N_4383);
nor U6848 (N_6848,N_4583,N_4697);
and U6849 (N_6849,N_4863,N_3532);
nor U6850 (N_6850,N_4279,N_4660);
nand U6851 (N_6851,N_2810,N_2984);
nor U6852 (N_6852,N_4170,N_3870);
nand U6853 (N_6853,N_4979,N_4511);
nor U6854 (N_6854,N_3152,N_3405);
and U6855 (N_6855,N_3463,N_2751);
nor U6856 (N_6856,N_2511,N_2870);
and U6857 (N_6857,N_2691,N_3919);
nor U6858 (N_6858,N_4235,N_4290);
or U6859 (N_6859,N_3438,N_3178);
or U6860 (N_6860,N_2661,N_3994);
nand U6861 (N_6861,N_3276,N_4511);
nand U6862 (N_6862,N_3586,N_4859);
and U6863 (N_6863,N_3156,N_2864);
nor U6864 (N_6864,N_2539,N_4452);
nand U6865 (N_6865,N_4752,N_2614);
nor U6866 (N_6866,N_4934,N_3791);
or U6867 (N_6867,N_4117,N_3384);
and U6868 (N_6868,N_3874,N_3067);
or U6869 (N_6869,N_3593,N_4767);
nor U6870 (N_6870,N_2671,N_2604);
xor U6871 (N_6871,N_2537,N_4656);
nand U6872 (N_6872,N_2608,N_4407);
nor U6873 (N_6873,N_4528,N_3236);
nand U6874 (N_6874,N_4680,N_3560);
nand U6875 (N_6875,N_4908,N_3981);
or U6876 (N_6876,N_3476,N_3840);
and U6877 (N_6877,N_3718,N_4024);
or U6878 (N_6878,N_4361,N_4924);
or U6879 (N_6879,N_2614,N_4384);
or U6880 (N_6880,N_3457,N_4270);
or U6881 (N_6881,N_2545,N_4486);
and U6882 (N_6882,N_3539,N_2745);
nand U6883 (N_6883,N_3058,N_3597);
xor U6884 (N_6884,N_4566,N_4739);
and U6885 (N_6885,N_4125,N_3411);
xor U6886 (N_6886,N_3788,N_4214);
xor U6887 (N_6887,N_3955,N_2964);
or U6888 (N_6888,N_3996,N_4670);
nand U6889 (N_6889,N_2559,N_4473);
and U6890 (N_6890,N_4660,N_4017);
nor U6891 (N_6891,N_3375,N_4034);
and U6892 (N_6892,N_2987,N_2603);
nor U6893 (N_6893,N_4115,N_4658);
nand U6894 (N_6894,N_2513,N_2580);
or U6895 (N_6895,N_4406,N_3654);
nand U6896 (N_6896,N_4214,N_4942);
or U6897 (N_6897,N_3398,N_3550);
nand U6898 (N_6898,N_4973,N_2717);
xnor U6899 (N_6899,N_4481,N_4018);
nor U6900 (N_6900,N_3190,N_3152);
and U6901 (N_6901,N_4392,N_3521);
nand U6902 (N_6902,N_3545,N_3299);
and U6903 (N_6903,N_3750,N_4128);
and U6904 (N_6904,N_4494,N_3087);
and U6905 (N_6905,N_3675,N_3305);
and U6906 (N_6906,N_4277,N_4302);
or U6907 (N_6907,N_4469,N_3321);
and U6908 (N_6908,N_3640,N_4969);
nor U6909 (N_6909,N_4015,N_2974);
or U6910 (N_6910,N_3452,N_4333);
or U6911 (N_6911,N_3983,N_2916);
xnor U6912 (N_6912,N_4102,N_2928);
nor U6913 (N_6913,N_4629,N_4588);
nand U6914 (N_6914,N_4949,N_4551);
or U6915 (N_6915,N_4660,N_3611);
xnor U6916 (N_6916,N_3905,N_2971);
or U6917 (N_6917,N_3312,N_2984);
nand U6918 (N_6918,N_4724,N_4398);
nor U6919 (N_6919,N_2560,N_4158);
or U6920 (N_6920,N_4340,N_3798);
xor U6921 (N_6921,N_3957,N_4089);
xnor U6922 (N_6922,N_3073,N_3333);
nand U6923 (N_6923,N_4821,N_3740);
nand U6924 (N_6924,N_2903,N_2764);
nand U6925 (N_6925,N_2825,N_3242);
nor U6926 (N_6926,N_3501,N_2597);
nor U6927 (N_6927,N_4159,N_4151);
nor U6928 (N_6928,N_3509,N_2702);
nand U6929 (N_6929,N_4531,N_4132);
nand U6930 (N_6930,N_4637,N_4887);
or U6931 (N_6931,N_4350,N_2736);
nor U6932 (N_6932,N_2505,N_4446);
nand U6933 (N_6933,N_4055,N_3103);
and U6934 (N_6934,N_4617,N_2769);
nand U6935 (N_6935,N_3828,N_4611);
nand U6936 (N_6936,N_3753,N_3001);
nor U6937 (N_6937,N_4739,N_4353);
nor U6938 (N_6938,N_3607,N_3635);
and U6939 (N_6939,N_2572,N_3762);
or U6940 (N_6940,N_4075,N_2631);
nor U6941 (N_6941,N_4516,N_2556);
nor U6942 (N_6942,N_2895,N_3629);
nand U6943 (N_6943,N_3047,N_4065);
nand U6944 (N_6944,N_4685,N_3534);
nand U6945 (N_6945,N_4344,N_3641);
nand U6946 (N_6946,N_4717,N_4314);
and U6947 (N_6947,N_2805,N_2847);
or U6948 (N_6948,N_4656,N_4733);
nor U6949 (N_6949,N_4926,N_2648);
xor U6950 (N_6950,N_2973,N_3726);
nor U6951 (N_6951,N_2515,N_4355);
nor U6952 (N_6952,N_3109,N_3368);
nand U6953 (N_6953,N_3438,N_4989);
xor U6954 (N_6954,N_2655,N_3391);
xnor U6955 (N_6955,N_4205,N_4530);
nor U6956 (N_6956,N_2726,N_2932);
nand U6957 (N_6957,N_3083,N_4264);
nor U6958 (N_6958,N_3905,N_4174);
nor U6959 (N_6959,N_2573,N_2795);
or U6960 (N_6960,N_4002,N_4145);
or U6961 (N_6961,N_2698,N_4542);
nand U6962 (N_6962,N_3391,N_4591);
or U6963 (N_6963,N_4902,N_3450);
or U6964 (N_6964,N_3343,N_4638);
nor U6965 (N_6965,N_3894,N_3387);
or U6966 (N_6966,N_2500,N_4312);
and U6967 (N_6967,N_3734,N_3175);
or U6968 (N_6968,N_3811,N_2635);
and U6969 (N_6969,N_4330,N_3212);
nand U6970 (N_6970,N_4542,N_2559);
nor U6971 (N_6971,N_3584,N_3494);
nand U6972 (N_6972,N_4477,N_4363);
nor U6973 (N_6973,N_2877,N_2630);
or U6974 (N_6974,N_3902,N_4971);
and U6975 (N_6975,N_3870,N_3438);
xor U6976 (N_6976,N_3335,N_2941);
or U6977 (N_6977,N_4230,N_4065);
nor U6978 (N_6978,N_3386,N_3435);
or U6979 (N_6979,N_2682,N_4885);
nor U6980 (N_6980,N_4209,N_4823);
or U6981 (N_6981,N_4165,N_3517);
nor U6982 (N_6982,N_4695,N_4924);
nor U6983 (N_6983,N_4169,N_2933);
and U6984 (N_6984,N_4633,N_4916);
or U6985 (N_6985,N_4988,N_4982);
nor U6986 (N_6986,N_4973,N_3322);
nor U6987 (N_6987,N_3179,N_3131);
xnor U6988 (N_6988,N_2797,N_4354);
nand U6989 (N_6989,N_2893,N_3200);
or U6990 (N_6990,N_3301,N_3140);
nand U6991 (N_6991,N_2790,N_4772);
and U6992 (N_6992,N_3506,N_4565);
nor U6993 (N_6993,N_3148,N_3026);
nor U6994 (N_6994,N_2922,N_4689);
or U6995 (N_6995,N_4301,N_3835);
or U6996 (N_6996,N_3379,N_2935);
nand U6997 (N_6997,N_2731,N_4925);
and U6998 (N_6998,N_3084,N_4987);
or U6999 (N_6999,N_2798,N_2587);
nor U7000 (N_7000,N_4034,N_4824);
nand U7001 (N_7001,N_3238,N_4554);
nand U7002 (N_7002,N_3540,N_3438);
nand U7003 (N_7003,N_4876,N_3255);
or U7004 (N_7004,N_2873,N_4349);
nand U7005 (N_7005,N_2934,N_2813);
and U7006 (N_7006,N_4410,N_3002);
nor U7007 (N_7007,N_3269,N_2787);
xor U7008 (N_7008,N_2687,N_4144);
nor U7009 (N_7009,N_3784,N_3325);
nand U7010 (N_7010,N_3533,N_2675);
or U7011 (N_7011,N_3880,N_3868);
nand U7012 (N_7012,N_4089,N_3809);
and U7013 (N_7013,N_3946,N_2621);
nand U7014 (N_7014,N_2637,N_4876);
or U7015 (N_7015,N_4629,N_3887);
nor U7016 (N_7016,N_4380,N_4878);
nor U7017 (N_7017,N_2758,N_2707);
and U7018 (N_7018,N_4230,N_4702);
or U7019 (N_7019,N_3375,N_4686);
xor U7020 (N_7020,N_3963,N_4837);
and U7021 (N_7021,N_3083,N_4422);
nand U7022 (N_7022,N_3325,N_2800);
or U7023 (N_7023,N_3268,N_4635);
and U7024 (N_7024,N_4398,N_3083);
and U7025 (N_7025,N_4542,N_2915);
nand U7026 (N_7026,N_3030,N_4729);
or U7027 (N_7027,N_3189,N_3229);
nand U7028 (N_7028,N_3472,N_3083);
and U7029 (N_7029,N_3145,N_4655);
nor U7030 (N_7030,N_2517,N_2601);
xnor U7031 (N_7031,N_2901,N_3145);
nand U7032 (N_7032,N_4003,N_3526);
and U7033 (N_7033,N_4581,N_2860);
nand U7034 (N_7034,N_4620,N_4991);
xnor U7035 (N_7035,N_3280,N_4721);
nand U7036 (N_7036,N_3442,N_4290);
and U7037 (N_7037,N_4980,N_3430);
nor U7038 (N_7038,N_3984,N_2628);
nor U7039 (N_7039,N_3945,N_2929);
nor U7040 (N_7040,N_2632,N_4874);
xor U7041 (N_7041,N_3534,N_2583);
nor U7042 (N_7042,N_2735,N_2690);
and U7043 (N_7043,N_4254,N_2884);
or U7044 (N_7044,N_3264,N_3458);
or U7045 (N_7045,N_3123,N_4359);
nor U7046 (N_7046,N_2716,N_3269);
and U7047 (N_7047,N_3788,N_3224);
nor U7048 (N_7048,N_3726,N_3126);
or U7049 (N_7049,N_4944,N_2670);
or U7050 (N_7050,N_2999,N_2844);
nor U7051 (N_7051,N_4628,N_2878);
nor U7052 (N_7052,N_3480,N_3888);
nor U7053 (N_7053,N_4248,N_3934);
and U7054 (N_7054,N_4666,N_2995);
nand U7055 (N_7055,N_4195,N_4616);
nand U7056 (N_7056,N_3840,N_2715);
xnor U7057 (N_7057,N_2605,N_3340);
and U7058 (N_7058,N_2610,N_4972);
nand U7059 (N_7059,N_4452,N_3065);
xnor U7060 (N_7060,N_4723,N_3632);
xnor U7061 (N_7061,N_2502,N_2797);
nor U7062 (N_7062,N_2876,N_4066);
nor U7063 (N_7063,N_2864,N_4417);
or U7064 (N_7064,N_4216,N_4619);
or U7065 (N_7065,N_4854,N_2867);
nor U7066 (N_7066,N_3408,N_2930);
or U7067 (N_7067,N_2642,N_4690);
nand U7068 (N_7068,N_4489,N_4586);
nand U7069 (N_7069,N_4310,N_2507);
nor U7070 (N_7070,N_3481,N_4688);
or U7071 (N_7071,N_3755,N_4346);
xnor U7072 (N_7072,N_3822,N_2589);
nand U7073 (N_7073,N_2753,N_3494);
nor U7074 (N_7074,N_4201,N_3561);
or U7075 (N_7075,N_4715,N_4047);
nor U7076 (N_7076,N_4340,N_4794);
or U7077 (N_7077,N_4485,N_4550);
xor U7078 (N_7078,N_3793,N_4122);
or U7079 (N_7079,N_3483,N_2887);
nor U7080 (N_7080,N_3554,N_2566);
or U7081 (N_7081,N_3682,N_4077);
xor U7082 (N_7082,N_2994,N_4634);
or U7083 (N_7083,N_4587,N_4068);
nor U7084 (N_7084,N_4259,N_3304);
nand U7085 (N_7085,N_2692,N_4972);
nor U7086 (N_7086,N_2966,N_3606);
nand U7087 (N_7087,N_3042,N_2508);
and U7088 (N_7088,N_4617,N_3127);
or U7089 (N_7089,N_3467,N_3444);
and U7090 (N_7090,N_2927,N_2800);
and U7091 (N_7091,N_2694,N_4746);
nand U7092 (N_7092,N_3118,N_4719);
or U7093 (N_7093,N_3170,N_3699);
and U7094 (N_7094,N_2505,N_3439);
nand U7095 (N_7095,N_2898,N_2918);
and U7096 (N_7096,N_4084,N_3387);
xor U7097 (N_7097,N_4719,N_4731);
nor U7098 (N_7098,N_3899,N_2791);
or U7099 (N_7099,N_4941,N_2738);
and U7100 (N_7100,N_2903,N_3288);
xnor U7101 (N_7101,N_3704,N_2654);
nor U7102 (N_7102,N_3210,N_3152);
nand U7103 (N_7103,N_3748,N_3859);
xnor U7104 (N_7104,N_4848,N_2782);
and U7105 (N_7105,N_4413,N_4948);
and U7106 (N_7106,N_2671,N_3513);
nor U7107 (N_7107,N_2711,N_4023);
xor U7108 (N_7108,N_2932,N_3246);
nor U7109 (N_7109,N_2700,N_2977);
or U7110 (N_7110,N_2589,N_4423);
xor U7111 (N_7111,N_3633,N_4440);
or U7112 (N_7112,N_4419,N_3569);
and U7113 (N_7113,N_4075,N_4471);
nand U7114 (N_7114,N_3555,N_4633);
nor U7115 (N_7115,N_3339,N_3094);
or U7116 (N_7116,N_3365,N_4395);
nand U7117 (N_7117,N_3340,N_3582);
and U7118 (N_7118,N_4850,N_4878);
or U7119 (N_7119,N_4358,N_2611);
nor U7120 (N_7120,N_3848,N_4144);
or U7121 (N_7121,N_4719,N_4960);
nor U7122 (N_7122,N_2897,N_3650);
xnor U7123 (N_7123,N_3412,N_4543);
xor U7124 (N_7124,N_2954,N_3336);
and U7125 (N_7125,N_3089,N_3116);
nor U7126 (N_7126,N_2855,N_4784);
nor U7127 (N_7127,N_3133,N_3564);
and U7128 (N_7128,N_2796,N_2827);
or U7129 (N_7129,N_3838,N_2606);
and U7130 (N_7130,N_2852,N_4348);
xor U7131 (N_7131,N_4769,N_3175);
and U7132 (N_7132,N_2965,N_4654);
or U7133 (N_7133,N_2939,N_3936);
nor U7134 (N_7134,N_4676,N_2618);
and U7135 (N_7135,N_2628,N_3598);
and U7136 (N_7136,N_2963,N_4815);
or U7137 (N_7137,N_4500,N_2567);
nand U7138 (N_7138,N_3933,N_3605);
nand U7139 (N_7139,N_2557,N_2657);
or U7140 (N_7140,N_3019,N_2838);
and U7141 (N_7141,N_3771,N_4187);
or U7142 (N_7142,N_4243,N_2794);
and U7143 (N_7143,N_3322,N_2617);
nand U7144 (N_7144,N_4635,N_4054);
or U7145 (N_7145,N_3921,N_4865);
and U7146 (N_7146,N_2558,N_4020);
or U7147 (N_7147,N_3113,N_4932);
nor U7148 (N_7148,N_3436,N_2813);
and U7149 (N_7149,N_2892,N_4433);
and U7150 (N_7150,N_4603,N_3061);
and U7151 (N_7151,N_3478,N_3862);
nand U7152 (N_7152,N_2598,N_4793);
nand U7153 (N_7153,N_3432,N_4723);
nor U7154 (N_7154,N_3555,N_3911);
nand U7155 (N_7155,N_2627,N_4790);
nand U7156 (N_7156,N_3843,N_3440);
and U7157 (N_7157,N_3356,N_3003);
or U7158 (N_7158,N_2507,N_3576);
nand U7159 (N_7159,N_3764,N_3111);
nor U7160 (N_7160,N_4041,N_3269);
and U7161 (N_7161,N_3470,N_2604);
nor U7162 (N_7162,N_4242,N_3851);
and U7163 (N_7163,N_3730,N_2673);
and U7164 (N_7164,N_4848,N_2841);
and U7165 (N_7165,N_3774,N_4977);
xnor U7166 (N_7166,N_4188,N_4020);
or U7167 (N_7167,N_4986,N_2875);
nor U7168 (N_7168,N_3481,N_4466);
or U7169 (N_7169,N_4011,N_4135);
or U7170 (N_7170,N_3034,N_2869);
nor U7171 (N_7171,N_3214,N_2596);
nand U7172 (N_7172,N_3856,N_2616);
xnor U7173 (N_7173,N_4930,N_3878);
nor U7174 (N_7174,N_4066,N_2858);
nand U7175 (N_7175,N_4216,N_2787);
xnor U7176 (N_7176,N_2885,N_3281);
nor U7177 (N_7177,N_4667,N_3458);
or U7178 (N_7178,N_2806,N_3108);
nand U7179 (N_7179,N_3680,N_4909);
nor U7180 (N_7180,N_4551,N_4902);
and U7181 (N_7181,N_2858,N_3168);
xor U7182 (N_7182,N_3896,N_4079);
or U7183 (N_7183,N_3763,N_3868);
and U7184 (N_7184,N_3332,N_3239);
and U7185 (N_7185,N_4104,N_4731);
or U7186 (N_7186,N_2548,N_2716);
nand U7187 (N_7187,N_3496,N_2652);
and U7188 (N_7188,N_2857,N_3874);
or U7189 (N_7189,N_4766,N_2714);
and U7190 (N_7190,N_3467,N_3255);
nand U7191 (N_7191,N_3208,N_3614);
nor U7192 (N_7192,N_3925,N_2732);
nand U7193 (N_7193,N_2886,N_2895);
or U7194 (N_7194,N_2779,N_3360);
nor U7195 (N_7195,N_3694,N_3205);
or U7196 (N_7196,N_2610,N_3920);
nor U7197 (N_7197,N_3283,N_3773);
xnor U7198 (N_7198,N_4696,N_4703);
or U7199 (N_7199,N_4605,N_4830);
nor U7200 (N_7200,N_4442,N_2827);
nor U7201 (N_7201,N_3228,N_3547);
nand U7202 (N_7202,N_4841,N_2812);
nand U7203 (N_7203,N_4025,N_4126);
nor U7204 (N_7204,N_4613,N_3694);
nor U7205 (N_7205,N_2878,N_3537);
nand U7206 (N_7206,N_2572,N_3370);
nor U7207 (N_7207,N_3258,N_4909);
and U7208 (N_7208,N_3701,N_4909);
nor U7209 (N_7209,N_3707,N_3906);
nand U7210 (N_7210,N_4941,N_4181);
or U7211 (N_7211,N_4827,N_4754);
nand U7212 (N_7212,N_3360,N_4887);
and U7213 (N_7213,N_4262,N_4040);
and U7214 (N_7214,N_4592,N_3045);
and U7215 (N_7215,N_3336,N_2814);
and U7216 (N_7216,N_4045,N_4508);
nand U7217 (N_7217,N_4224,N_3422);
nor U7218 (N_7218,N_2991,N_3498);
or U7219 (N_7219,N_3771,N_4924);
nand U7220 (N_7220,N_2882,N_4625);
or U7221 (N_7221,N_3204,N_4490);
or U7222 (N_7222,N_3955,N_3967);
and U7223 (N_7223,N_4439,N_3990);
nand U7224 (N_7224,N_3635,N_3439);
or U7225 (N_7225,N_4468,N_2585);
xnor U7226 (N_7226,N_4270,N_4328);
nand U7227 (N_7227,N_4818,N_4998);
nand U7228 (N_7228,N_3751,N_3092);
or U7229 (N_7229,N_3406,N_4451);
and U7230 (N_7230,N_3580,N_4854);
nor U7231 (N_7231,N_3183,N_4721);
nand U7232 (N_7232,N_4503,N_4707);
or U7233 (N_7233,N_4538,N_3427);
nor U7234 (N_7234,N_3844,N_3040);
or U7235 (N_7235,N_3649,N_2902);
and U7236 (N_7236,N_3601,N_4710);
nand U7237 (N_7237,N_4318,N_4891);
or U7238 (N_7238,N_4748,N_3996);
or U7239 (N_7239,N_2505,N_2729);
or U7240 (N_7240,N_2986,N_3483);
xnor U7241 (N_7241,N_3664,N_2580);
nand U7242 (N_7242,N_4692,N_3762);
xor U7243 (N_7243,N_3326,N_3412);
nand U7244 (N_7244,N_2642,N_2540);
nand U7245 (N_7245,N_4714,N_4445);
nand U7246 (N_7246,N_3920,N_3511);
or U7247 (N_7247,N_3012,N_3911);
and U7248 (N_7248,N_2984,N_4498);
or U7249 (N_7249,N_2945,N_2803);
nand U7250 (N_7250,N_3959,N_2942);
xor U7251 (N_7251,N_2508,N_3338);
or U7252 (N_7252,N_3656,N_3575);
nor U7253 (N_7253,N_2985,N_3364);
nand U7254 (N_7254,N_2901,N_3119);
and U7255 (N_7255,N_3848,N_2807);
nor U7256 (N_7256,N_2732,N_3880);
nor U7257 (N_7257,N_4295,N_2679);
and U7258 (N_7258,N_4372,N_4062);
nand U7259 (N_7259,N_4695,N_2813);
and U7260 (N_7260,N_3620,N_4615);
and U7261 (N_7261,N_2514,N_3985);
and U7262 (N_7262,N_3107,N_4043);
xnor U7263 (N_7263,N_4155,N_3806);
nand U7264 (N_7264,N_4840,N_3115);
and U7265 (N_7265,N_3157,N_4190);
and U7266 (N_7266,N_3373,N_3599);
and U7267 (N_7267,N_2834,N_4399);
and U7268 (N_7268,N_2724,N_4540);
and U7269 (N_7269,N_4233,N_2729);
xor U7270 (N_7270,N_4894,N_2634);
nor U7271 (N_7271,N_3455,N_2619);
xor U7272 (N_7272,N_4717,N_4661);
or U7273 (N_7273,N_4385,N_3959);
or U7274 (N_7274,N_4013,N_2788);
xnor U7275 (N_7275,N_4940,N_4427);
nor U7276 (N_7276,N_2898,N_4954);
xnor U7277 (N_7277,N_3330,N_4499);
nor U7278 (N_7278,N_3405,N_3746);
nand U7279 (N_7279,N_3005,N_4951);
and U7280 (N_7280,N_3967,N_2864);
nor U7281 (N_7281,N_4108,N_4600);
nand U7282 (N_7282,N_3737,N_3359);
and U7283 (N_7283,N_3920,N_2624);
and U7284 (N_7284,N_3831,N_3199);
and U7285 (N_7285,N_3405,N_3195);
nand U7286 (N_7286,N_4938,N_3812);
nor U7287 (N_7287,N_4482,N_4794);
and U7288 (N_7288,N_4502,N_4200);
nand U7289 (N_7289,N_4984,N_4824);
xor U7290 (N_7290,N_4870,N_2818);
nand U7291 (N_7291,N_3678,N_3163);
and U7292 (N_7292,N_4325,N_2959);
or U7293 (N_7293,N_3779,N_2942);
nand U7294 (N_7294,N_3235,N_3520);
or U7295 (N_7295,N_3345,N_3998);
nor U7296 (N_7296,N_3617,N_4514);
or U7297 (N_7297,N_3500,N_2707);
nand U7298 (N_7298,N_3385,N_4648);
nor U7299 (N_7299,N_3387,N_4523);
nand U7300 (N_7300,N_3738,N_3564);
xor U7301 (N_7301,N_2990,N_4723);
xnor U7302 (N_7302,N_3333,N_4900);
nand U7303 (N_7303,N_4164,N_3033);
xor U7304 (N_7304,N_4397,N_2805);
nor U7305 (N_7305,N_2507,N_4487);
nor U7306 (N_7306,N_3888,N_3885);
and U7307 (N_7307,N_2700,N_4109);
nor U7308 (N_7308,N_3849,N_2937);
nor U7309 (N_7309,N_4869,N_4708);
and U7310 (N_7310,N_3700,N_4046);
nor U7311 (N_7311,N_3950,N_3801);
xor U7312 (N_7312,N_4765,N_4750);
and U7313 (N_7313,N_4123,N_3193);
nor U7314 (N_7314,N_3464,N_4966);
and U7315 (N_7315,N_4603,N_3920);
xor U7316 (N_7316,N_4273,N_4062);
and U7317 (N_7317,N_3977,N_2627);
or U7318 (N_7318,N_4243,N_3841);
and U7319 (N_7319,N_3596,N_4819);
nor U7320 (N_7320,N_4304,N_4723);
or U7321 (N_7321,N_4589,N_2578);
nor U7322 (N_7322,N_3763,N_2627);
nor U7323 (N_7323,N_4497,N_4294);
nand U7324 (N_7324,N_4784,N_2651);
and U7325 (N_7325,N_3268,N_4670);
and U7326 (N_7326,N_2888,N_4679);
or U7327 (N_7327,N_4221,N_3214);
xnor U7328 (N_7328,N_2654,N_4192);
nand U7329 (N_7329,N_3754,N_4391);
and U7330 (N_7330,N_4162,N_4712);
nor U7331 (N_7331,N_4882,N_2798);
or U7332 (N_7332,N_3599,N_4739);
nand U7333 (N_7333,N_4426,N_4162);
nand U7334 (N_7334,N_4043,N_4547);
xnor U7335 (N_7335,N_2693,N_2712);
nor U7336 (N_7336,N_3351,N_3669);
or U7337 (N_7337,N_4032,N_4265);
and U7338 (N_7338,N_3918,N_4336);
nand U7339 (N_7339,N_4154,N_3012);
nor U7340 (N_7340,N_2533,N_4300);
xnor U7341 (N_7341,N_2790,N_4744);
or U7342 (N_7342,N_2843,N_2694);
xnor U7343 (N_7343,N_2817,N_4221);
or U7344 (N_7344,N_4143,N_4209);
or U7345 (N_7345,N_4768,N_2974);
nor U7346 (N_7346,N_2952,N_3276);
or U7347 (N_7347,N_4290,N_3094);
or U7348 (N_7348,N_4188,N_3040);
or U7349 (N_7349,N_3946,N_2615);
nor U7350 (N_7350,N_4412,N_4160);
or U7351 (N_7351,N_4787,N_4579);
nor U7352 (N_7352,N_4990,N_3365);
nor U7353 (N_7353,N_3355,N_4959);
nor U7354 (N_7354,N_3745,N_3456);
nor U7355 (N_7355,N_3248,N_2534);
and U7356 (N_7356,N_3888,N_4891);
nand U7357 (N_7357,N_3266,N_4204);
nand U7358 (N_7358,N_2851,N_2747);
or U7359 (N_7359,N_4404,N_3955);
xnor U7360 (N_7360,N_4563,N_3218);
nor U7361 (N_7361,N_4296,N_2733);
nand U7362 (N_7362,N_4150,N_4925);
nor U7363 (N_7363,N_3464,N_3152);
and U7364 (N_7364,N_3395,N_3590);
nor U7365 (N_7365,N_2686,N_4938);
and U7366 (N_7366,N_3215,N_4208);
and U7367 (N_7367,N_2623,N_2633);
nand U7368 (N_7368,N_4777,N_3473);
nand U7369 (N_7369,N_4666,N_4531);
nand U7370 (N_7370,N_4786,N_4864);
and U7371 (N_7371,N_2992,N_4101);
xor U7372 (N_7372,N_3282,N_3224);
and U7373 (N_7373,N_4430,N_3960);
nor U7374 (N_7374,N_4000,N_3960);
and U7375 (N_7375,N_3954,N_2952);
nor U7376 (N_7376,N_3500,N_4226);
and U7377 (N_7377,N_4996,N_2535);
nand U7378 (N_7378,N_3792,N_2830);
nor U7379 (N_7379,N_3337,N_3308);
xor U7380 (N_7380,N_4451,N_2638);
nor U7381 (N_7381,N_4730,N_4942);
and U7382 (N_7382,N_2776,N_4040);
and U7383 (N_7383,N_2801,N_4229);
nor U7384 (N_7384,N_4866,N_4391);
or U7385 (N_7385,N_3978,N_3803);
nor U7386 (N_7386,N_3144,N_3243);
and U7387 (N_7387,N_4812,N_4476);
and U7388 (N_7388,N_3558,N_2591);
nor U7389 (N_7389,N_3569,N_4941);
nand U7390 (N_7390,N_4691,N_4186);
nand U7391 (N_7391,N_4941,N_3183);
nor U7392 (N_7392,N_3339,N_3354);
and U7393 (N_7393,N_4382,N_4252);
or U7394 (N_7394,N_3881,N_2681);
nor U7395 (N_7395,N_3037,N_2970);
nor U7396 (N_7396,N_3965,N_4115);
xor U7397 (N_7397,N_3437,N_3678);
nor U7398 (N_7398,N_3597,N_2962);
xor U7399 (N_7399,N_3219,N_3852);
or U7400 (N_7400,N_4655,N_3531);
and U7401 (N_7401,N_2745,N_3151);
nand U7402 (N_7402,N_4278,N_4838);
and U7403 (N_7403,N_3675,N_3969);
or U7404 (N_7404,N_4809,N_3408);
nand U7405 (N_7405,N_2956,N_2517);
nand U7406 (N_7406,N_3828,N_2950);
nor U7407 (N_7407,N_4353,N_3082);
and U7408 (N_7408,N_3479,N_4101);
or U7409 (N_7409,N_3628,N_2954);
or U7410 (N_7410,N_3783,N_3817);
or U7411 (N_7411,N_4449,N_3151);
or U7412 (N_7412,N_2807,N_4677);
nor U7413 (N_7413,N_2638,N_4101);
nand U7414 (N_7414,N_2546,N_3225);
or U7415 (N_7415,N_4009,N_3473);
nor U7416 (N_7416,N_3137,N_4707);
and U7417 (N_7417,N_4231,N_2787);
and U7418 (N_7418,N_3834,N_4119);
and U7419 (N_7419,N_3182,N_2864);
and U7420 (N_7420,N_4579,N_3856);
nand U7421 (N_7421,N_3086,N_3995);
and U7422 (N_7422,N_4021,N_3977);
or U7423 (N_7423,N_4028,N_4695);
and U7424 (N_7424,N_4187,N_4712);
nor U7425 (N_7425,N_4842,N_4753);
nor U7426 (N_7426,N_3101,N_2696);
nor U7427 (N_7427,N_2805,N_4344);
nor U7428 (N_7428,N_3203,N_3085);
and U7429 (N_7429,N_3100,N_2872);
and U7430 (N_7430,N_4502,N_3097);
nand U7431 (N_7431,N_3938,N_3437);
nor U7432 (N_7432,N_3686,N_3190);
or U7433 (N_7433,N_2881,N_4020);
xor U7434 (N_7434,N_3628,N_3314);
nand U7435 (N_7435,N_4204,N_4128);
xnor U7436 (N_7436,N_4250,N_4520);
nor U7437 (N_7437,N_4500,N_3041);
xnor U7438 (N_7438,N_3330,N_4253);
nand U7439 (N_7439,N_3429,N_4484);
and U7440 (N_7440,N_2860,N_2649);
or U7441 (N_7441,N_3447,N_3666);
and U7442 (N_7442,N_4766,N_2539);
nor U7443 (N_7443,N_3316,N_4259);
xor U7444 (N_7444,N_2618,N_2982);
nor U7445 (N_7445,N_2728,N_4857);
nor U7446 (N_7446,N_3212,N_3089);
xor U7447 (N_7447,N_4832,N_3489);
nor U7448 (N_7448,N_3973,N_2763);
nor U7449 (N_7449,N_4128,N_2548);
and U7450 (N_7450,N_4524,N_3438);
and U7451 (N_7451,N_3162,N_3546);
nor U7452 (N_7452,N_4446,N_3753);
nand U7453 (N_7453,N_3027,N_4551);
nor U7454 (N_7454,N_3321,N_4674);
or U7455 (N_7455,N_4083,N_4329);
and U7456 (N_7456,N_3665,N_3910);
nor U7457 (N_7457,N_3599,N_3833);
and U7458 (N_7458,N_3386,N_4628);
nor U7459 (N_7459,N_2621,N_4250);
nor U7460 (N_7460,N_2540,N_4277);
nor U7461 (N_7461,N_4382,N_4105);
or U7462 (N_7462,N_3512,N_3136);
or U7463 (N_7463,N_4667,N_4970);
and U7464 (N_7464,N_4979,N_2957);
nand U7465 (N_7465,N_2738,N_2923);
xor U7466 (N_7466,N_2528,N_3707);
nand U7467 (N_7467,N_4816,N_4539);
or U7468 (N_7468,N_3184,N_2609);
and U7469 (N_7469,N_3237,N_3036);
and U7470 (N_7470,N_2811,N_3600);
nor U7471 (N_7471,N_4002,N_3739);
xor U7472 (N_7472,N_3390,N_3940);
nor U7473 (N_7473,N_4605,N_3065);
xnor U7474 (N_7474,N_2994,N_3601);
nor U7475 (N_7475,N_2917,N_3197);
and U7476 (N_7476,N_4590,N_2961);
or U7477 (N_7477,N_4929,N_3779);
xor U7478 (N_7478,N_4979,N_4135);
nand U7479 (N_7479,N_4049,N_3002);
nor U7480 (N_7480,N_2680,N_4175);
and U7481 (N_7481,N_2643,N_4313);
or U7482 (N_7482,N_4441,N_2570);
xnor U7483 (N_7483,N_3241,N_3347);
or U7484 (N_7484,N_3993,N_3142);
nand U7485 (N_7485,N_2953,N_3418);
or U7486 (N_7486,N_3117,N_4576);
and U7487 (N_7487,N_4756,N_2547);
nand U7488 (N_7488,N_4185,N_4033);
or U7489 (N_7489,N_3437,N_3446);
or U7490 (N_7490,N_2741,N_2945);
and U7491 (N_7491,N_2927,N_4675);
or U7492 (N_7492,N_4171,N_2864);
or U7493 (N_7493,N_3170,N_2981);
nand U7494 (N_7494,N_3377,N_4734);
or U7495 (N_7495,N_4974,N_4920);
nor U7496 (N_7496,N_3599,N_2839);
nor U7497 (N_7497,N_2954,N_2565);
xnor U7498 (N_7498,N_2984,N_3691);
and U7499 (N_7499,N_3970,N_4450);
and U7500 (N_7500,N_6260,N_6938);
nand U7501 (N_7501,N_5097,N_5203);
and U7502 (N_7502,N_5341,N_5169);
or U7503 (N_7503,N_7471,N_5268);
or U7504 (N_7504,N_7314,N_5763);
or U7505 (N_7505,N_6604,N_7028);
xnor U7506 (N_7506,N_6226,N_5312);
nand U7507 (N_7507,N_5325,N_6431);
and U7508 (N_7508,N_6791,N_6977);
nand U7509 (N_7509,N_5824,N_5062);
or U7510 (N_7510,N_5012,N_7371);
and U7511 (N_7511,N_5231,N_6259);
nor U7512 (N_7512,N_6637,N_5354);
nand U7513 (N_7513,N_5099,N_7243);
xnor U7514 (N_7514,N_5044,N_6150);
and U7515 (N_7515,N_5077,N_6053);
xnor U7516 (N_7516,N_5800,N_7275);
or U7517 (N_7517,N_7043,N_7153);
nand U7518 (N_7518,N_6082,N_5749);
nand U7519 (N_7519,N_5886,N_6099);
or U7520 (N_7520,N_6972,N_6366);
and U7521 (N_7521,N_6342,N_6327);
and U7522 (N_7522,N_7173,N_5756);
nand U7523 (N_7523,N_6732,N_5738);
or U7524 (N_7524,N_6687,N_6591);
and U7525 (N_7525,N_6577,N_5730);
nor U7526 (N_7526,N_5794,N_5467);
nand U7527 (N_7527,N_5092,N_5436);
nand U7528 (N_7528,N_5880,N_6896);
xnor U7529 (N_7529,N_7041,N_5226);
nor U7530 (N_7530,N_5858,N_6971);
and U7531 (N_7531,N_6098,N_5120);
or U7532 (N_7532,N_6521,N_7181);
nand U7533 (N_7533,N_7320,N_5248);
and U7534 (N_7534,N_5121,N_5629);
and U7535 (N_7535,N_7435,N_7364);
and U7536 (N_7536,N_7042,N_5750);
or U7537 (N_7537,N_5619,N_6237);
nor U7538 (N_7538,N_6111,N_5257);
nand U7539 (N_7539,N_6831,N_5442);
nor U7540 (N_7540,N_6446,N_5844);
and U7541 (N_7541,N_5389,N_6454);
nor U7542 (N_7542,N_5335,N_6176);
nand U7543 (N_7543,N_6912,N_6549);
or U7544 (N_7544,N_5412,N_6235);
nor U7545 (N_7545,N_5684,N_5328);
nor U7546 (N_7546,N_5019,N_5520);
nand U7547 (N_7547,N_6215,N_5899);
xnor U7548 (N_7548,N_6566,N_5586);
nor U7549 (N_7549,N_6136,N_5941);
nand U7550 (N_7550,N_6069,N_6090);
nand U7551 (N_7551,N_6390,N_7218);
nand U7552 (N_7552,N_6878,N_6149);
and U7553 (N_7553,N_7140,N_5770);
or U7554 (N_7554,N_5283,N_6655);
and U7555 (N_7555,N_6444,N_6122);
nand U7556 (N_7556,N_5584,N_7497);
nand U7557 (N_7557,N_6120,N_5994);
nor U7558 (N_7558,N_7118,N_7369);
and U7559 (N_7559,N_6401,N_5218);
nor U7560 (N_7560,N_6983,N_5713);
or U7561 (N_7561,N_6561,N_5219);
nor U7562 (N_7562,N_5543,N_6834);
or U7563 (N_7563,N_6658,N_5262);
nand U7564 (N_7564,N_5188,N_5965);
and U7565 (N_7565,N_6633,N_6994);
nor U7566 (N_7566,N_6715,N_6282);
nor U7567 (N_7567,N_6460,N_5392);
nor U7568 (N_7568,N_6776,N_5876);
or U7569 (N_7569,N_6712,N_7341);
or U7570 (N_7570,N_5228,N_6389);
nor U7571 (N_7571,N_6100,N_5346);
nand U7572 (N_7572,N_5212,N_6334);
nor U7573 (N_7573,N_5802,N_6175);
nor U7574 (N_7574,N_5846,N_7160);
nand U7575 (N_7575,N_5680,N_6234);
xnor U7576 (N_7576,N_6246,N_5276);
or U7577 (N_7577,N_5109,N_7293);
nor U7578 (N_7578,N_6699,N_5870);
or U7579 (N_7579,N_5871,N_5816);
xnor U7580 (N_7580,N_5801,N_7002);
nor U7581 (N_7581,N_5477,N_6611);
nand U7582 (N_7582,N_7003,N_5060);
nand U7583 (N_7583,N_6719,N_6425);
nor U7584 (N_7584,N_7139,N_6110);
nand U7585 (N_7585,N_6770,N_6932);
xor U7586 (N_7586,N_6574,N_7068);
and U7587 (N_7587,N_5417,N_6157);
nor U7588 (N_7588,N_6199,N_5175);
and U7589 (N_7589,N_5926,N_6899);
nand U7590 (N_7590,N_5494,N_6908);
nand U7591 (N_7591,N_5665,N_6598);
nand U7592 (N_7592,N_5768,N_5727);
nor U7593 (N_7593,N_5697,N_5920);
nand U7594 (N_7594,N_6336,N_6459);
nor U7595 (N_7595,N_6347,N_6991);
and U7596 (N_7596,N_7361,N_6421);
and U7597 (N_7597,N_5183,N_5516);
nor U7598 (N_7598,N_7337,N_5910);
or U7599 (N_7599,N_5551,N_5464);
nor U7600 (N_7600,N_5894,N_5326);
and U7601 (N_7601,N_5435,N_6513);
nand U7602 (N_7602,N_7481,N_6754);
nand U7603 (N_7603,N_5017,N_5433);
nor U7604 (N_7604,N_6393,N_5990);
and U7605 (N_7605,N_5925,N_5302);
or U7606 (N_7606,N_7020,N_6382);
nand U7607 (N_7607,N_5461,N_5029);
nor U7608 (N_7608,N_5042,N_7257);
and U7609 (N_7609,N_6553,N_5180);
xnor U7610 (N_7610,N_5654,N_5174);
or U7611 (N_7611,N_5995,N_5122);
nand U7612 (N_7612,N_5480,N_6021);
nand U7613 (N_7613,N_6974,N_7036);
or U7614 (N_7614,N_5891,N_6548);
nand U7615 (N_7615,N_7116,N_6490);
nand U7616 (N_7616,N_6755,N_6473);
nand U7617 (N_7617,N_6484,N_5033);
nand U7618 (N_7618,N_6000,N_7027);
and U7619 (N_7619,N_6312,N_7047);
nor U7620 (N_7620,N_5934,N_5372);
or U7621 (N_7621,N_5245,N_7237);
nor U7622 (N_7622,N_5274,N_5428);
or U7623 (N_7623,N_7133,N_7071);
nor U7624 (N_7624,N_6154,N_5306);
nor U7625 (N_7625,N_6787,N_5708);
or U7626 (N_7626,N_6092,N_6284);
or U7627 (N_7627,N_5655,N_6358);
or U7628 (N_7628,N_5152,N_5553);
xor U7629 (N_7629,N_6057,N_5488);
nor U7630 (N_7630,N_6860,N_6560);
nor U7631 (N_7631,N_6159,N_6047);
or U7632 (N_7632,N_5695,N_5625);
xnor U7633 (N_7633,N_5474,N_7468);
nor U7634 (N_7634,N_6918,N_5585);
and U7635 (N_7635,N_6089,N_5015);
nand U7636 (N_7636,N_6507,N_7374);
nand U7637 (N_7637,N_7455,N_6919);
and U7638 (N_7638,N_7394,N_5783);
and U7639 (N_7639,N_7034,N_6813);
nor U7640 (N_7640,N_6769,N_6863);
nor U7641 (N_7641,N_6703,N_5361);
and U7642 (N_7642,N_7021,N_6868);
nand U7643 (N_7643,N_5492,N_5338);
nand U7644 (N_7644,N_7297,N_6893);
nand U7645 (N_7645,N_6224,N_5451);
nor U7646 (N_7646,N_5378,N_7015);
nand U7647 (N_7647,N_6391,N_6188);
and U7648 (N_7648,N_7215,N_6816);
nor U7649 (N_7649,N_5052,N_6422);
or U7650 (N_7650,N_6432,N_5754);
or U7651 (N_7651,N_6048,N_5736);
and U7652 (N_7652,N_5342,N_5829);
and U7653 (N_7653,N_6094,N_6172);
and U7654 (N_7654,N_5281,N_5278);
and U7655 (N_7655,N_6556,N_6563);
or U7656 (N_7656,N_5963,N_5444);
nand U7657 (N_7657,N_6790,N_6420);
and U7658 (N_7658,N_7113,N_6360);
xor U7659 (N_7659,N_6998,N_6876);
or U7660 (N_7660,N_5500,N_6608);
nor U7661 (N_7661,N_5637,N_6151);
nor U7662 (N_7662,N_7454,N_5315);
or U7663 (N_7663,N_6626,N_5298);
nand U7664 (N_7664,N_6130,N_7208);
nor U7665 (N_7665,N_5303,N_7357);
xnor U7666 (N_7666,N_6323,N_5172);
or U7667 (N_7667,N_5096,N_7379);
nor U7668 (N_7668,N_7209,N_5836);
nor U7669 (N_7669,N_5462,N_5513);
and U7670 (N_7670,N_5463,N_6129);
nand U7671 (N_7671,N_5550,N_6445);
nand U7672 (N_7672,N_7233,N_7194);
and U7673 (N_7673,N_5159,N_5571);
nand U7674 (N_7674,N_5205,N_6929);
nand U7675 (N_7675,N_5470,N_6798);
or U7676 (N_7676,N_5536,N_5771);
nand U7677 (N_7677,N_6913,N_5983);
or U7678 (N_7678,N_5631,N_7039);
or U7679 (N_7679,N_5230,N_5577);
or U7680 (N_7680,N_6081,N_6286);
xor U7681 (N_7681,N_6522,N_7235);
and U7682 (N_7682,N_6709,N_5757);
nand U7683 (N_7683,N_5630,N_6239);
nor U7684 (N_7684,N_5943,N_5616);
or U7685 (N_7685,N_6836,N_6250);
xor U7686 (N_7686,N_5072,N_5093);
nand U7687 (N_7687,N_6737,N_7044);
or U7688 (N_7688,N_7007,N_6964);
and U7689 (N_7689,N_5251,N_5959);
and U7690 (N_7690,N_7001,N_5234);
or U7691 (N_7691,N_6984,N_6631);
nor U7692 (N_7692,N_6486,N_5530);
nand U7693 (N_7693,N_5517,N_5569);
nor U7694 (N_7694,N_6030,N_7158);
nor U7695 (N_7695,N_6435,N_5991);
or U7696 (N_7696,N_6480,N_6669);
and U7697 (N_7697,N_5032,N_7350);
xnor U7698 (N_7698,N_5945,N_7360);
nand U7699 (N_7699,N_6008,N_7413);
or U7700 (N_7700,N_6299,N_7114);
nand U7701 (N_7701,N_6781,N_5216);
and U7702 (N_7702,N_5425,N_6520);
nor U7703 (N_7703,N_6346,N_6031);
nand U7704 (N_7704,N_7256,N_6039);
and U7705 (N_7705,N_7095,N_5366);
nand U7706 (N_7706,N_6487,N_6541);
nor U7707 (N_7707,N_6070,N_7366);
nor U7708 (N_7708,N_6332,N_6620);
or U7709 (N_7709,N_7420,N_6305);
nor U7710 (N_7710,N_6468,N_6397);
and U7711 (N_7711,N_5731,N_7059);
and U7712 (N_7712,N_6281,N_5656);
nor U7713 (N_7713,N_7060,N_6704);
nand U7714 (N_7714,N_7424,N_6132);
or U7715 (N_7715,N_5336,N_7087);
and U7716 (N_7716,N_6850,N_6204);
or U7717 (N_7717,N_5322,N_5168);
nand U7718 (N_7718,N_6488,N_6195);
or U7719 (N_7719,N_5021,N_5901);
and U7720 (N_7720,N_6551,N_6858);
nand U7721 (N_7721,N_6121,N_7473);
nand U7722 (N_7722,N_5080,N_7339);
or U7723 (N_7723,N_6362,N_6605);
nand U7724 (N_7724,N_6174,N_6838);
and U7725 (N_7725,N_7202,N_7014);
xor U7726 (N_7726,N_6536,N_6666);
and U7727 (N_7727,N_7382,N_6124);
xnor U7728 (N_7728,N_7469,N_7197);
nand U7729 (N_7729,N_5084,N_6399);
xor U7730 (N_7730,N_7229,N_5562);
or U7731 (N_7731,N_5013,N_5030);
or U7732 (N_7732,N_5971,N_6276);
and U7733 (N_7733,N_6163,N_6768);
nand U7734 (N_7734,N_7412,N_6368);
nor U7735 (N_7735,N_6474,N_5086);
or U7736 (N_7736,N_7093,N_6529);
and U7737 (N_7737,N_5604,N_5842);
and U7738 (N_7738,N_6001,N_6270);
nand U7739 (N_7739,N_6245,N_6871);
xnor U7740 (N_7740,N_5137,N_5862);
and U7741 (N_7741,N_6958,N_5307);
or U7742 (N_7742,N_5568,N_5985);
nor U7743 (N_7743,N_5284,N_7164);
xor U7744 (N_7744,N_5566,N_7092);
nor U7745 (N_7745,N_6872,N_6212);
and U7746 (N_7746,N_5744,N_5046);
and U7747 (N_7747,N_6557,N_7057);
or U7748 (N_7748,N_7037,N_5064);
nand U7749 (N_7749,N_7077,N_5496);
or U7750 (N_7750,N_5753,N_7423);
nand U7751 (N_7751,N_5495,N_7405);
xnor U7752 (N_7752,N_5944,N_7462);
nand U7753 (N_7753,N_6503,N_5673);
and U7754 (N_7754,N_7288,N_5652);
and U7755 (N_7755,N_5523,N_7415);
or U7756 (N_7756,N_6202,N_5459);
nand U7757 (N_7757,N_5831,N_5045);
nand U7758 (N_7758,N_5647,N_5238);
or U7759 (N_7759,N_6580,N_5194);
nand U7760 (N_7760,N_5337,N_5821);
or U7761 (N_7761,N_5117,N_6131);
nor U7762 (N_7762,N_6895,N_5385);
and U7763 (N_7763,N_6624,N_6192);
and U7764 (N_7764,N_5690,N_5332);
or U7765 (N_7765,N_5683,N_5712);
xnor U7766 (N_7766,N_6293,N_6359);
or U7767 (N_7767,N_7000,N_6277);
nor U7768 (N_7768,N_6238,N_5192);
or U7769 (N_7769,N_7207,N_5161);
nand U7770 (N_7770,N_5643,N_5005);
xor U7771 (N_7771,N_5634,N_7389);
or U7772 (N_7772,N_5349,N_6470);
nor U7773 (N_7773,N_5884,N_5449);
and U7774 (N_7774,N_6583,N_7403);
and U7775 (N_7775,N_7024,N_5733);
and U7776 (N_7776,N_6355,N_7079);
and U7777 (N_7777,N_6430,N_6706);
nand U7778 (N_7778,N_5674,N_7226);
and U7779 (N_7779,N_5726,N_5171);
nand U7780 (N_7780,N_5747,N_6603);
nor U7781 (N_7781,N_6379,N_6980);
and U7782 (N_7782,N_5393,N_7308);
and U7783 (N_7783,N_5331,N_5196);
or U7784 (N_7784,N_5138,N_6833);
or U7785 (N_7785,N_7120,N_5297);
and U7786 (N_7786,N_6266,N_5431);
and U7787 (N_7787,N_7284,N_7063);
or U7788 (N_7788,N_5798,N_6927);
nor U7789 (N_7789,N_5782,N_6668);
xnor U7790 (N_7790,N_7427,N_6573);
xor U7791 (N_7791,N_7102,N_6437);
and U7792 (N_7792,N_6640,N_5575);
nand U7793 (N_7793,N_7285,N_6128);
or U7794 (N_7794,N_5486,N_6112);
xnor U7795 (N_7795,N_6800,N_7245);
and U7796 (N_7796,N_6537,N_7483);
nand U7797 (N_7797,N_6588,N_5678);
nor U7798 (N_7798,N_5107,N_5922);
and U7799 (N_7799,N_7182,N_6644);
and U7800 (N_7800,N_7219,N_7480);
nand U7801 (N_7801,N_6823,N_7432);
or U7802 (N_7802,N_5221,N_6153);
nor U7803 (N_7803,N_5693,N_7484);
xor U7804 (N_7804,N_6877,N_5839);
nand U7805 (N_7805,N_5528,N_7330);
nand U7806 (N_7806,N_5270,N_6595);
and U7807 (N_7807,N_5947,N_5102);
nand U7808 (N_7808,N_6279,N_5125);
nor U7809 (N_7809,N_5993,N_7175);
nor U7810 (N_7810,N_5623,N_7258);
nor U7811 (N_7811,N_5848,N_5371);
or U7812 (N_7812,N_5058,N_6967);
nand U7813 (N_7813,N_5984,N_6632);
nor U7814 (N_7814,N_7367,N_6410);
nand U7815 (N_7815,N_5182,N_6020);
nand U7816 (N_7816,N_6254,N_7107);
nand U7817 (N_7817,N_6278,N_6308);
nor U7818 (N_7818,N_7310,N_6680);
and U7819 (N_7819,N_5565,N_6394);
nand U7820 (N_7820,N_5157,N_6329);
nand U7821 (N_7821,N_5904,N_5454);
and U7822 (N_7822,N_7298,N_6141);
or U7823 (N_7823,N_5620,N_6073);
nor U7824 (N_7824,N_7378,N_5438);
and U7825 (N_7825,N_6331,N_6819);
and U7826 (N_7826,N_6406,N_6027);
xnor U7827 (N_7827,N_6814,N_5432);
or U7828 (N_7828,N_6223,N_6744);
or U7829 (N_7829,N_7381,N_5511);
and U7830 (N_7830,N_5469,N_5557);
nor U7831 (N_7831,N_6171,N_6975);
nor U7832 (N_7832,N_6702,N_6742);
nand U7833 (N_7833,N_6880,N_5386);
nand U7834 (N_7834,N_5003,N_5612);
and U7835 (N_7835,N_5900,N_6063);
and U7836 (N_7836,N_5919,N_6181);
nand U7837 (N_7837,N_7008,N_5721);
or U7838 (N_7838,N_6014,N_5069);
or U7839 (N_7839,N_7248,N_6185);
or U7840 (N_7840,N_5139,N_6652);
or U7841 (N_7841,N_5826,N_5924);
xnor U7842 (N_7842,N_6255,N_6959);
nor U7843 (N_7843,N_6808,N_5942);
and U7844 (N_7844,N_5751,N_6736);
nor U7845 (N_7845,N_6690,N_5987);
or U7846 (N_7846,N_5938,N_7477);
and U7847 (N_7847,N_6085,N_7206);
or U7848 (N_7848,N_5008,N_5746);
and U7849 (N_7849,N_5561,N_5388);
xnor U7850 (N_7850,N_5186,N_6585);
nor U7851 (N_7851,N_6679,N_7163);
xor U7852 (N_7852,N_5074,N_5155);
or U7853 (N_7853,N_7242,N_5752);
and U7854 (N_7854,N_5741,N_6989);
nand U7855 (N_7855,N_5930,N_6267);
and U7856 (N_7856,N_5447,N_5698);
nand U7857 (N_7857,N_6726,N_7395);
and U7858 (N_7858,N_6933,N_7377);
and U7859 (N_7859,N_6518,N_5936);
and U7860 (N_7860,N_5970,N_7200);
nor U7861 (N_7861,N_5755,N_6214);
or U7862 (N_7862,N_6888,N_6201);
or U7863 (N_7863,N_6493,N_7017);
xnor U7864 (N_7864,N_5398,N_5319);
nor U7865 (N_7865,N_5351,N_6367);
nor U7866 (N_7866,N_7333,N_5081);
and U7867 (N_7867,N_7273,N_5272);
nor U7868 (N_7868,N_5394,N_6718);
or U7869 (N_7869,N_7165,N_5031);
nor U7870 (N_7870,N_6567,N_6155);
or U7871 (N_7871,N_6562,N_6012);
or U7872 (N_7872,N_6458,N_7434);
and U7873 (N_7873,N_6618,N_5692);
or U7874 (N_7874,N_7383,N_5650);
nand U7875 (N_7875,N_6965,N_5540);
nand U7876 (N_7876,N_6761,N_5705);
or U7877 (N_7877,N_6407,N_6166);
or U7878 (N_7878,N_7190,N_7272);
nor U7879 (N_7879,N_5148,N_7023);
nand U7880 (N_7880,N_6685,N_5440);
nand U7881 (N_7881,N_6182,N_6852);
or U7882 (N_7882,N_5113,N_6427);
and U7883 (N_7883,N_5701,N_5601);
and U7884 (N_7884,N_5864,N_6928);
nand U7885 (N_7885,N_5885,N_5147);
nor U7886 (N_7886,N_5506,N_6630);
nand U7887 (N_7887,N_6987,N_5723);
xor U7888 (N_7888,N_7254,N_5198);
nand U7889 (N_7889,N_7217,N_5381);
nor U7890 (N_7890,N_5819,N_5524);
nand U7891 (N_7891,N_6638,N_6211);
or U7892 (N_7892,N_5016,N_5413);
nand U7893 (N_7893,N_6449,N_5580);
nor U7894 (N_7894,N_7072,N_7408);
and U7895 (N_7895,N_5256,N_6935);
nor U7896 (N_7896,N_5908,N_5410);
and U7897 (N_7897,N_5989,N_5696);
and U7898 (N_7898,N_6263,N_6409);
or U7899 (N_7899,N_7046,N_5881);
and U7900 (N_7900,N_7121,N_7051);
nand U7901 (N_7901,N_6050,N_6827);
and U7902 (N_7902,N_5593,N_5711);
nand U7903 (N_7903,N_5764,N_6647);
or U7904 (N_7904,N_7445,N_6601);
nand U7905 (N_7905,N_7451,N_6721);
and U7906 (N_7906,N_7104,N_7195);
or U7907 (N_7907,N_5600,N_6649);
and U7908 (N_7908,N_5905,N_6165);
xor U7909 (N_7909,N_5460,N_6290);
and U7910 (N_7910,N_7425,N_5290);
nand U7911 (N_7911,N_6496,N_6784);
or U7912 (N_7912,N_6506,N_6043);
or U7913 (N_7913,N_7355,N_7204);
or U7914 (N_7914,N_5423,N_6572);
xnor U7915 (N_7915,N_6351,N_7253);
or U7916 (N_7916,N_5402,N_6997);
nand U7917 (N_7917,N_7391,N_5572);
xor U7918 (N_7918,N_5422,N_7436);
or U7919 (N_7919,N_6956,N_5377);
nor U7920 (N_7920,N_7183,N_6797);
nor U7921 (N_7921,N_5067,N_5057);
nor U7922 (N_7922,N_5691,N_5788);
nand U7923 (N_7923,N_6571,N_6426);
nor U7924 (N_7924,N_6302,N_5966);
xnor U7925 (N_7925,N_5745,N_7280);
and U7926 (N_7926,N_5807,N_5988);
or U7927 (N_7927,N_5050,N_7187);
and U7928 (N_7928,N_6416,N_7111);
nand U7929 (N_7929,N_5646,N_7363);
and U7930 (N_7930,N_7301,N_6249);
or U7931 (N_7931,N_5728,N_7441);
and U7932 (N_7932,N_7287,N_5531);
or U7933 (N_7933,N_6711,N_5158);
or U7934 (N_7934,N_5441,N_7141);
and U7935 (N_7935,N_5363,N_6142);
nor U7936 (N_7936,N_6418,N_6477);
nor U7937 (N_7937,N_6384,N_7212);
nand U7938 (N_7938,N_7167,N_6526);
nor U7939 (N_7939,N_6064,N_6225);
and U7940 (N_7940,N_5641,N_5118);
nand U7941 (N_7941,N_6764,N_5823);
or U7942 (N_7942,N_5666,N_5808);
xor U7943 (N_7943,N_5254,N_5855);
nor U7944 (N_7944,N_7213,N_7127);
nor U7945 (N_7945,N_5888,N_6862);
xor U7946 (N_7946,N_6095,N_6482);
xor U7947 (N_7947,N_5838,N_5668);
nand U7948 (N_7948,N_6613,N_6102);
nand U7949 (N_7949,N_5418,N_6137);
and U7950 (N_7950,N_7365,N_6147);
nor U7951 (N_7951,N_5209,N_5964);
nand U7952 (N_7952,N_5865,N_6514);
or U7953 (N_7953,N_6535,N_6954);
nand U7954 (N_7954,N_6162,N_5275);
xor U7955 (N_7955,N_6478,N_5797);
nor U7956 (N_7956,N_7075,N_5103);
nor U7957 (N_7957,N_7013,N_6544);
nand U7958 (N_7958,N_6909,N_7388);
or U7959 (N_7959,N_6330,N_6208);
nor U7960 (N_7960,N_6320,N_7085);
nor U7961 (N_7961,N_6545,N_7495);
nand U7962 (N_7962,N_7407,N_6476);
or U7963 (N_7963,N_7159,N_6735);
nor U7964 (N_7964,N_7033,N_5887);
or U7965 (N_7965,N_6222,N_5301);
and U7966 (N_7966,N_7313,N_5707);
nand U7967 (N_7967,N_6058,N_6350);
nand U7968 (N_7968,N_5061,N_5709);
and U7969 (N_7969,N_7125,N_6939);
or U7970 (N_7970,N_6156,N_5853);
and U7971 (N_7971,N_5260,N_7440);
nor U7972 (N_7972,N_7205,N_5804);
and U7973 (N_7973,N_5352,N_7069);
nor U7974 (N_7974,N_5515,N_6206);
and U7975 (N_7975,N_6855,N_7180);
and U7976 (N_7976,N_7155,N_6848);
and U7977 (N_7977,N_6055,N_6584);
nor U7978 (N_7978,N_5603,N_5043);
xnor U7979 (N_7979,N_6947,N_5403);
and U7980 (N_7980,N_7119,N_6576);
nand U7981 (N_7981,N_5973,N_5617);
and U7982 (N_7982,N_6766,N_6772);
xor U7983 (N_7983,N_5505,N_5976);
nand U7984 (N_7984,N_6803,N_6375);
nand U7985 (N_7985,N_6906,N_6722);
nor U7986 (N_7986,N_6148,N_6291);
or U7987 (N_7987,N_7409,N_6361);
or U7988 (N_7988,N_7249,N_7225);
and U7989 (N_7989,N_5979,N_7305);
nand U7990 (N_7990,N_6625,N_6849);
nor U7991 (N_7991,N_5591,N_6752);
nor U7992 (N_7992,N_6785,N_5376);
nand U7993 (N_7993,N_6412,N_7324);
nor U7994 (N_7994,N_7074,N_5784);
xnor U7995 (N_7995,N_5390,N_6904);
and U7996 (N_7996,N_6372,N_6970);
or U7997 (N_7997,N_5574,N_6428);
or U7998 (N_7998,N_6118,N_5588);
or U7999 (N_7999,N_5261,N_6845);
nor U8000 (N_8000,N_5089,N_6882);
nor U8001 (N_8001,N_6728,N_6317);
xor U8002 (N_8002,N_5368,N_6309);
xnor U8003 (N_8003,N_7344,N_7128);
nand U8004 (N_8004,N_7099,N_6804);
or U8005 (N_8005,N_6341,N_6106);
and U8006 (N_8006,N_6499,N_7384);
nor U8007 (N_8007,N_6258,N_5189);
nand U8008 (N_8008,N_5578,N_6140);
and U8009 (N_8009,N_6794,N_7134);
xnor U8010 (N_8010,N_6930,N_6472);
nor U8011 (N_8011,N_7376,N_5841);
and U8012 (N_8012,N_7005,N_7117);
nand U8013 (N_8013,N_6925,N_6657);
nand U8014 (N_8014,N_6104,N_6515);
or U8015 (N_8015,N_6024,N_7016);
nand U8016 (N_8016,N_7472,N_6639);
nor U8017 (N_8017,N_5615,N_6753);
and U8018 (N_8018,N_6292,N_6433);
and U8019 (N_8019,N_7169,N_5645);
or U8020 (N_8020,N_7453,N_6310);
nor U8021 (N_8021,N_6240,N_6992);
and U8022 (N_8022,N_5642,N_6883);
and U8023 (N_8023,N_5380,N_6253);
or U8024 (N_8024,N_5404,N_6558);
nor U8025 (N_8025,N_7385,N_5953);
and U8026 (N_8026,N_5471,N_6619);
xnor U8027 (N_8027,N_5890,N_5676);
nor U8028 (N_8028,N_5407,N_5236);
or U8029 (N_8029,N_5840,N_5405);
xor U8030 (N_8030,N_6530,N_6673);
nand U8031 (N_8031,N_7426,N_6108);
or U8032 (N_8032,N_6288,N_7038);
nand U8033 (N_8033,N_6979,N_6842);
nor U8034 (N_8034,N_5179,N_5482);
nand U8035 (N_8035,N_6607,N_5535);
nand U8036 (N_8036,N_7231,N_5142);
nand U8037 (N_8037,N_6228,N_5555);
nand U8038 (N_8038,N_7354,N_6133);
and U8039 (N_8039,N_6554,N_5859);
and U8040 (N_8040,N_6453,N_6579);
nor U8041 (N_8041,N_5197,N_6217);
xnor U8042 (N_8042,N_6773,N_7326);
or U8043 (N_8043,N_7422,N_6636);
nand U8044 (N_8044,N_6189,N_5025);
nand U8045 (N_8045,N_5559,N_7315);
nand U8046 (N_8046,N_5508,N_7397);
or U8047 (N_8047,N_6191,N_5285);
and U8048 (N_8048,N_7349,N_5448);
and U8049 (N_8049,N_6623,N_7496);
nand U8050 (N_8050,N_7211,N_5348);
nand U8051 (N_8051,N_7278,N_5825);
and U8052 (N_8052,N_6581,N_6378);
xnor U8053 (N_8053,N_6948,N_7252);
nand U8054 (N_8054,N_6550,N_5658);
xnor U8055 (N_8055,N_5490,N_6101);
nand U8056 (N_8056,N_5126,N_6910);
and U8057 (N_8057,N_7457,N_6186);
nor U8058 (N_8058,N_5857,N_7410);
or U8059 (N_8059,N_6243,N_5329);
and U8060 (N_8060,N_5076,N_7261);
or U8061 (N_8061,N_5453,N_5609);
and U8062 (N_8062,N_6807,N_5957);
or U8063 (N_8063,N_7241,N_6143);
and U8064 (N_8064,N_6645,N_6916);
or U8065 (N_8065,N_5048,N_5367);
and U8066 (N_8066,N_6606,N_6661);
nand U8067 (N_8067,N_5040,N_5362);
xnor U8068 (N_8068,N_6667,N_5539);
nand U8069 (N_8069,N_5415,N_5101);
and U8070 (N_8070,N_6738,N_6303);
nor U8071 (N_8071,N_5686,N_6628);
and U8072 (N_8072,N_5774,N_5547);
nand U8073 (N_8073,N_6621,N_5724);
or U8074 (N_8074,N_6127,N_6009);
xor U8075 (N_8075,N_6894,N_5408);
or U8076 (N_8076,N_6516,N_7049);
xor U8077 (N_8077,N_6086,N_6796);
nand U8078 (N_8078,N_6065,N_5160);
nand U8079 (N_8079,N_6083,N_6252);
nand U8080 (N_8080,N_6392,N_6693);
and U8081 (N_8081,N_5271,N_5455);
nand U8082 (N_8082,N_5960,N_5140);
nor U8083 (N_8083,N_6835,N_5071);
nor U8084 (N_8084,N_5079,N_6067);
xnor U8085 (N_8085,N_5739,N_6400);
and U8086 (N_8086,N_6914,N_5977);
nor U8087 (N_8087,N_5735,N_5187);
nor U8088 (N_8088,N_6398,N_6602);
or U8089 (N_8089,N_5982,N_5563);
or U8090 (N_8090,N_6475,N_5507);
and U8091 (N_8091,N_5475,N_6565);
nor U8092 (N_8092,N_5956,N_5769);
nor U8093 (N_8093,N_6751,N_5560);
nor U8094 (N_8094,N_6296,N_6966);
or U8095 (N_8095,N_5805,N_5590);
or U8096 (N_8096,N_6700,N_5426);
and U8097 (N_8097,N_5716,N_5622);
or U8098 (N_8098,N_7157,N_5677);
nand U8099 (N_8099,N_5070,N_6646);
or U8100 (N_8100,N_5780,N_5124);
nor U8101 (N_8101,N_6135,N_6046);
xnor U8102 (N_8102,N_7295,N_5384);
or U8103 (N_8103,N_7129,N_6178);
and U8104 (N_8104,N_5420,N_6114);
and U8105 (N_8105,N_6168,N_5310);
and U8106 (N_8106,N_5128,N_5318);
nor U8107 (N_8107,N_6694,N_7149);
and U8108 (N_8108,N_6547,N_5883);
nand U8109 (N_8109,N_5054,N_6374);
nor U8110 (N_8110,N_6404,N_6869);
and U8111 (N_8111,N_6450,N_6733);
nor U8112 (N_8112,N_5776,N_6256);
nor U8113 (N_8113,N_5063,N_6622);
or U8114 (N_8114,N_6665,N_6231);
nor U8115 (N_8115,N_7234,N_6789);
xor U8116 (N_8116,N_5785,N_6117);
and U8117 (N_8117,N_5485,N_6600);
or U8118 (N_8118,N_5204,N_7123);
and U8119 (N_8119,N_5534,N_7239);
nand U8120 (N_8120,N_5849,N_6826);
and U8121 (N_8121,N_7147,N_6750);
nor U8122 (N_8122,N_5667,N_5594);
nand U8123 (N_8123,N_5258,N_6257);
nand U8124 (N_8124,N_6011,N_7054);
xnor U8125 (N_8125,N_6386,N_7067);
xor U8126 (N_8126,N_5662,N_6886);
nand U8127 (N_8127,N_6993,N_5589);
or U8128 (N_8128,N_5409,N_5512);
nor U8129 (N_8129,N_7091,N_6139);
or U8130 (N_8130,N_5813,N_6898);
or U8131 (N_8131,N_7475,N_5323);
nor U8132 (N_8132,N_5759,N_6423);
nor U8133 (N_8133,N_6040,N_6889);
nor U8134 (N_8134,N_5468,N_5703);
or U8135 (N_8135,N_6701,N_6678);
xor U8136 (N_8136,N_5974,N_5567);
nand U8137 (N_8137,N_6955,N_5526);
xor U8138 (N_8138,N_5670,N_6280);
and U8139 (N_8139,N_6248,N_6677);
nor U8140 (N_8140,N_7490,N_5867);
nor U8141 (N_8141,N_6846,N_6822);
nor U8142 (N_8142,N_5694,N_5786);
nand U8143 (N_8143,N_7094,N_6152);
and U8144 (N_8144,N_7061,N_6339);
or U8145 (N_8145,N_5651,N_7429);
xnor U8146 (N_8146,N_7487,N_7387);
nand U8147 (N_8147,N_5817,N_7431);
or U8148 (N_8148,N_6395,N_7018);
xnor U8149 (N_8149,N_6749,N_6648);
and U8150 (N_8150,N_6697,N_7345);
or U8151 (N_8151,N_6837,N_6532);
or U8152 (N_8152,N_5240,N_7090);
and U8153 (N_8153,N_5777,N_6328);
nand U8154 (N_8154,N_6173,N_6995);
nor U8155 (N_8155,N_6061,N_6616);
nand U8156 (N_8156,N_6643,N_6370);
nor U8157 (N_8157,N_5660,N_5664);
nand U8158 (N_8158,N_6448,N_5522);
nor U8159 (N_8159,N_5932,N_5743);
or U8160 (N_8160,N_5207,N_6654);
nand U8161 (N_8161,N_7004,N_7031);
or U8162 (N_8162,N_5682,N_5835);
or U8163 (N_8163,N_6546,N_5151);
nand U8164 (N_8164,N_5949,N_6313);
or U8165 (N_8165,N_5065,N_5457);
and U8166 (N_8166,N_7089,N_5847);
and U8167 (N_8167,N_6840,N_6663);
nor U8168 (N_8168,N_5969,N_5837);
or U8169 (N_8169,N_6821,N_7312);
xor U8170 (N_8170,N_6874,N_6466);
and U8171 (N_8171,N_6216,N_5320);
and U8172 (N_8172,N_5596,N_5129);
nand U8173 (N_8173,N_6905,N_7185);
and U8174 (N_8174,N_6442,N_5446);
and U8175 (N_8175,N_5347,N_6036);
and U8176 (N_8176,N_5626,N_6716);
or U8177 (N_8177,N_6403,N_5259);
xnor U8178 (N_8178,N_7456,N_6025);
and U8179 (N_8179,N_5353,N_5399);
nor U8180 (N_8180,N_7221,N_7176);
nor U8181 (N_8181,N_6824,N_7268);
or U8182 (N_8182,N_6922,N_5163);
and U8183 (N_8183,N_5178,N_7414);
nor U8184 (N_8184,N_6818,N_6641);
or U8185 (N_8185,N_6538,N_7131);
nor U8186 (N_8186,N_5424,N_7066);
nand U8187 (N_8187,N_7292,N_6731);
nand U8188 (N_8188,N_6865,N_5244);
and U8189 (N_8189,N_6324,N_6345);
xnor U8190 (N_8190,N_5950,N_5465);
or U8191 (N_8191,N_7009,N_6978);
and U8192 (N_8192,N_7098,N_7096);
and U8193 (N_8193,N_7416,N_7110);
nor U8194 (N_8194,N_7136,N_6946);
xor U8195 (N_8195,N_7486,N_7448);
nor U8196 (N_8196,N_6109,N_6285);
and U8197 (N_8197,N_7115,N_6926);
nor U8198 (N_8198,N_5324,N_5355);
or U8199 (N_8199,N_5153,N_6113);
and U8200 (N_8200,N_6505,N_7331);
xnor U8201 (N_8201,N_5227,N_6745);
xor U8202 (N_8202,N_5689,N_5915);
or U8203 (N_8203,N_5912,N_5790);
xor U8204 (N_8204,N_5277,N_6032);
and U8205 (N_8205,N_6066,N_6782);
or U8206 (N_8206,N_6962,N_6635);
and U8207 (N_8207,N_6167,N_5809);
or U8208 (N_8208,N_6512,N_5980);
and U8209 (N_8209,N_5525,N_6501);
xnor U8210 (N_8210,N_6004,N_6672);
nand U8211 (N_8211,N_7442,N_7491);
nor U8212 (N_8212,N_6792,N_7452);
or U8213 (N_8213,N_6158,N_5317);
and U8214 (N_8214,N_6596,N_5878);
nor U8215 (N_8215,N_6028,N_5653);
and U8216 (N_8216,N_6170,N_6943);
nand U8217 (N_8217,N_7222,N_5502);
and U8218 (N_8218,N_6734,N_6016);
and U8219 (N_8219,N_5114,N_7168);
or U8220 (N_8220,N_7336,N_5445);
nor U8221 (N_8221,N_5748,N_6533);
nand U8222 (N_8222,N_5439,N_7319);
or U8223 (N_8223,N_5037,N_6023);
nand U8224 (N_8224,N_5098,N_7150);
or U8225 (N_8225,N_6125,N_5100);
nor U8226 (N_8226,N_6126,N_5533);
or U8227 (N_8227,N_6767,N_6957);
or U8228 (N_8228,N_6464,N_5856);
or U8229 (N_8229,N_6268,N_6042);
xor U8230 (N_8230,N_5373,N_5552);
nand U8231 (N_8231,N_6951,N_6969);
nor U8232 (N_8232,N_7179,N_5434);
and U8233 (N_8233,N_6924,N_5215);
and U8234 (N_8234,N_6740,N_5799);
nand U8235 (N_8235,N_5679,N_6037);
nand U8236 (N_8236,N_6720,N_5233);
xor U8237 (N_8237,N_5264,N_6319);
or U8238 (N_8238,N_6034,N_6315);
nand U8239 (N_8239,N_5532,N_7230);
nor U8240 (N_8240,N_7461,N_6318);
or U8241 (N_8241,N_7177,N_7465);
or U8242 (N_8242,N_6615,N_5199);
or U8243 (N_8243,N_5917,N_5370);
and U8244 (N_8244,N_6662,N_5927);
nand U8245 (N_8245,N_5487,N_6218);
nand U8246 (N_8246,N_6417,N_5929);
and U8247 (N_8247,N_6381,N_5165);
xor U8248 (N_8248,N_6756,N_5872);
or U8249 (N_8249,N_7406,N_6578);
nor U8250 (N_8250,N_6138,N_6200);
nand U8251 (N_8251,N_5288,N_5211);
or U8252 (N_8252,N_6900,N_5229);
nand U8253 (N_8253,N_5632,N_6080);
nor U8254 (N_8254,N_6710,N_6463);
and U8255 (N_8255,N_6614,N_6589);
xnor U8256 (N_8256,N_6002,N_7126);
and U8257 (N_8257,N_5430,N_6451);
and U8258 (N_8258,N_6262,N_6504);
or U8259 (N_8259,N_6941,N_7323);
nor U8260 (N_8260,N_6760,N_5006);
nor U8261 (N_8261,N_6273,N_7400);
or U8262 (N_8262,N_7100,N_6999);
nand U8263 (N_8263,N_5149,N_7251);
nand U8264 (N_8264,N_5243,N_5828);
or U8265 (N_8265,N_7282,N_7450);
or U8266 (N_8266,N_5663,N_5661);
nand U8267 (N_8267,N_5028,N_6942);
and U8268 (N_8268,N_6479,N_5011);
and U8269 (N_8269,N_7277,N_5822);
or U8270 (N_8270,N_6543,N_5111);
nand U8271 (N_8271,N_6795,N_5395);
or U8272 (N_8272,N_5239,N_5510);
and U8273 (N_8273,N_5918,N_6847);
or U8274 (N_8274,N_7380,N_5599);
or U8275 (N_8275,N_6832,N_5339);
and U8276 (N_8276,N_7232,N_6413);
and U8277 (N_8277,N_5350,N_7340);
nand U8278 (N_8278,N_6380,N_5644);
nor U8279 (N_8279,N_5897,N_7105);
or U8280 (N_8280,N_5742,N_7335);
nand U8281 (N_8281,N_6233,N_6870);
xor U8282 (N_8282,N_6272,N_6077);
nand U8283 (N_8283,N_7170,N_6660);
nand U8284 (N_8284,N_5007,N_7386);
and U8285 (N_8285,N_6686,N_6659);
or U8286 (N_8286,N_5191,N_5518);
nor U8287 (N_8287,N_5954,N_6038);
nor U8288 (N_8288,N_7303,N_7011);
or U8289 (N_8289,N_7271,N_5892);
nor U8290 (N_8290,N_7025,N_5869);
nand U8291 (N_8291,N_6976,N_7191);
and U8292 (N_8292,N_6612,N_6229);
nand U8293 (N_8293,N_5289,N_6707);
nand U8294 (N_8294,N_6953,N_5700);
and U8295 (N_8295,N_5791,N_5962);
nand U8296 (N_8296,N_5613,N_7198);
or U8297 (N_8297,N_7053,N_6227);
nand U8298 (N_8298,N_7390,N_7489);
or U8299 (N_8299,N_5955,N_5489);
or U8300 (N_8300,N_6019,N_7396);
nand U8301 (N_8301,N_6078,N_6076);
and U8302 (N_8302,N_5544,N_6307);
and U8303 (N_8303,N_5146,N_5879);
and U8304 (N_8304,N_5898,N_5483);
or U8305 (N_8305,N_5843,N_6003);
or U8306 (N_8306,N_7130,N_6817);
or U8307 (N_8307,N_6344,N_7056);
and U8308 (N_8308,N_5514,N_6568);
nor U8309 (N_8309,N_6590,N_5053);
nor U8310 (N_8310,N_5833,N_7493);
or U8311 (N_8311,N_6371,N_7368);
nand U8312 (N_8312,N_5997,N_5732);
and U8313 (N_8313,N_6569,N_5570);
nand U8314 (N_8314,N_5141,N_5018);
or U8315 (N_8315,N_5049,N_7088);
nand U8316 (N_8316,N_5308,N_7145);
nand U8317 (N_8317,N_5906,N_7498);
nor U8318 (N_8318,N_6364,N_6483);
and U8319 (N_8319,N_6439,N_6387);
nor U8320 (N_8320,N_5996,N_5911);
or U8321 (N_8321,N_5232,N_5291);
or U8322 (N_8322,N_7138,N_5581);
and U8323 (N_8323,N_7154,N_7266);
and U8324 (N_8324,N_5704,N_6917);
or U8325 (N_8325,N_5173,N_5611);
nor U8326 (N_8326,N_5875,N_5456);
or U8327 (N_8327,N_6314,N_6748);
and U8328 (N_8328,N_7283,N_5548);
and U8329 (N_8329,N_6041,N_6920);
nand U8330 (N_8330,N_6029,N_7076);
xnor U8331 (N_8331,N_5145,N_5247);
nor U8332 (N_8332,N_7398,N_5340);
xnor U8333 (N_8333,N_6103,N_5830);
and U8334 (N_8334,N_7291,N_5066);
and U8335 (N_8335,N_5214,N_5313);
or U8336 (N_8336,N_6134,N_7358);
and U8337 (N_8337,N_5250,N_6696);
nor U8338 (N_8338,N_6071,N_6123);
nand U8339 (N_8339,N_5091,N_5687);
nor U8340 (N_8340,N_7463,N_7332);
or U8341 (N_8341,N_6297,N_5521);
xor U8342 (N_8342,N_5280,N_5937);
and U8343 (N_8343,N_5316,N_7467);
or U8344 (N_8344,N_6656,N_6322);
or U8345 (N_8345,N_7351,N_5176);
or U8346 (N_8346,N_6294,N_6915);
or U8347 (N_8347,N_5729,N_5767);
or U8348 (N_8348,N_7137,N_5414);
nand U8349 (N_8349,N_6447,N_6179);
nor U8350 (N_8350,N_5916,N_5978);
nor U8351 (N_8351,N_5217,N_5010);
and U8352 (N_8352,N_6241,N_5095);
xnor U8353 (N_8353,N_6146,N_6436);
nand U8354 (N_8354,N_5541,N_7055);
and U8355 (N_8355,N_7108,N_7352);
xor U8356 (N_8356,N_6921,N_5734);
or U8357 (N_8357,N_7488,N_5133);
nor U8358 (N_8358,N_5714,N_7375);
nor U8359 (N_8359,N_7322,N_5452);
and U8360 (N_8360,N_5587,N_6617);
nand U8361 (N_8361,N_5860,N_6806);
and U8362 (N_8362,N_6841,N_6708);
nand U8363 (N_8363,N_6861,N_6843);
nor U8364 (N_8364,N_5014,N_7240);
xnor U8365 (N_8365,N_6045,N_6084);
or U8366 (N_8366,N_6783,N_6940);
xor U8367 (N_8367,N_6670,N_6952);
or U8368 (N_8368,N_6306,N_5608);
nor U8369 (N_8369,N_6741,N_7327);
xor U8370 (N_8370,N_6119,N_6799);
or U8371 (N_8371,N_7262,N_5811);
nor U8372 (N_8372,N_6242,N_5024);
or U8373 (N_8373,N_5778,N_6509);
or U8374 (N_8374,N_5400,N_6511);
nand U8375 (N_8375,N_6552,N_7460);
or U8376 (N_8376,N_6853,N_5252);
or U8377 (N_8377,N_7263,N_7144);
xnor U8378 (N_8378,N_5803,N_6060);
nor U8379 (N_8379,N_6338,N_6866);
nand U8380 (N_8380,N_6356,N_5967);
nor U8381 (N_8381,N_5190,N_6717);
and U8382 (N_8382,N_6337,N_6471);
xor U8383 (N_8383,N_6879,N_5419);
and U8384 (N_8384,N_7458,N_5968);
and U8385 (N_8385,N_5246,N_7019);
or U8386 (N_8386,N_5762,N_5542);
and U8387 (N_8387,N_6295,N_5210);
nor U8388 (N_8388,N_5773,N_5688);
or U8389 (N_8389,N_5699,N_5725);
xor U8390 (N_8390,N_5815,N_5443);
nor U8391 (N_8391,N_5206,N_5498);
nor U8392 (N_8392,N_6854,N_7404);
or U8393 (N_8393,N_6177,N_6586);
and U8394 (N_8394,N_6988,N_5476);
and U8395 (N_8395,N_6867,N_5056);
and U8396 (N_8396,N_6438,N_7276);
and U8397 (N_8397,N_5266,N_6534);
or U8398 (N_8398,N_7178,N_7080);
xor U8399 (N_8399,N_5618,N_5851);
nand U8400 (N_8400,N_6609,N_5556);
or U8401 (N_8401,N_6494,N_6013);
and U8402 (N_8402,N_5923,N_7210);
nand U8403 (N_8403,N_7238,N_6705);
nand U8404 (N_8404,N_7362,N_6990);
xnor U8405 (N_8405,N_7318,N_6363);
or U8406 (N_8406,N_5041,N_5614);
or U8407 (N_8407,N_6097,N_7296);
nor U8408 (N_8408,N_6684,N_5391);
or U8409 (N_8409,N_5863,N_6582);
nor U8410 (N_8410,N_5235,N_5576);
nor U8411 (N_8411,N_6691,N_6497);
and U8412 (N_8412,N_6365,N_5200);
nand U8413 (N_8413,N_7299,N_5546);
and U8414 (N_8414,N_6311,N_5304);
and U8415 (N_8415,N_7012,N_7439);
nor U8416 (N_8416,N_6209,N_5116);
nand U8417 (N_8417,N_6096,N_5951);
or U8418 (N_8418,N_7470,N_7459);
nand U8419 (N_8419,N_5610,N_5633);
xor U8420 (N_8420,N_7267,N_7216);
and U8421 (N_8421,N_7269,N_6072);
or U8422 (N_8422,N_6049,N_7040);
and U8423 (N_8423,N_6244,N_6221);
nand U8424 (N_8424,N_6357,N_6443);
nor U8425 (N_8425,N_5717,N_5009);
and U8426 (N_8426,N_7192,N_5224);
and U8427 (N_8427,N_5579,N_5027);
xor U8428 (N_8428,N_6369,N_6205);
nor U8429 (N_8429,N_7048,N_7485);
nor U8430 (N_8430,N_6903,N_7449);
nand U8431 (N_8431,N_6519,N_5669);
or U8432 (N_8432,N_7433,N_5627);
nand U8433 (N_8433,N_6196,N_7476);
xnor U8434 (N_8434,N_6396,N_5406);
nor U8435 (N_8435,N_6105,N_6779);
xnor U8436 (N_8436,N_5999,N_7199);
nor U8437 (N_8437,N_5628,N_7402);
xnor U8438 (N_8438,N_7304,N_5573);
nor U8439 (N_8439,N_5827,N_5493);
and U8440 (N_8440,N_7010,N_6683);
nor U8441 (N_8441,N_6996,N_6115);
xnor U8442 (N_8442,N_5772,N_5143);
and U8443 (N_8443,N_6193,N_5672);
nand U8444 (N_8444,N_5681,N_7172);
nor U8445 (N_8445,N_7166,N_5877);
or U8446 (N_8446,N_5657,N_6017);
nor U8447 (N_8447,N_6289,N_6385);
nand U8448 (N_8448,N_6007,N_6033);
nand U8449 (N_8449,N_7083,N_6269);
xnor U8450 (N_8450,N_5365,N_5648);
and U8451 (N_8451,N_5948,N_6161);
nor U8452 (N_8452,N_6981,N_7132);
nand U8453 (N_8453,N_7184,N_7328);
and U8454 (N_8454,N_6651,N_6074);
or U8455 (N_8455,N_6283,N_5020);
nand U8456 (N_8456,N_5595,N_6839);
nor U8457 (N_8457,N_6844,N_5255);
and U8458 (N_8458,N_5334,N_5921);
nor U8459 (N_8459,N_5237,N_5914);
and U8460 (N_8460,N_5383,N_6326);
nor U8461 (N_8461,N_6570,N_7466);
nand U8462 (N_8462,N_5852,N_7045);
xnor U8463 (N_8463,N_6671,N_5715);
or U8464 (N_8464,N_7464,N_5110);
or U8465 (N_8465,N_5002,N_5273);
nand U8466 (N_8466,N_6730,N_5000);
nor U8467 (N_8467,N_7329,N_7035);
or U8468 (N_8468,N_6873,N_6945);
xor U8469 (N_8469,N_5127,N_6739);
nand U8470 (N_8470,N_6907,N_6219);
nand U8471 (N_8471,N_6775,N_6316);
and U8472 (N_8472,N_7255,N_5537);
nor U8473 (N_8473,N_5893,N_7347);
nand U8474 (N_8474,N_6759,N_7188);
nand U8475 (N_8475,N_7279,N_6901);
nand U8476 (N_8476,N_6184,N_5082);
nor U8477 (N_8477,N_6725,N_6236);
or U8478 (N_8478,N_5499,N_7342);
or U8479 (N_8479,N_6461,N_5760);
and U8480 (N_8480,N_6884,N_6207);
and U8481 (N_8481,N_5806,N_5850);
or U8482 (N_8482,N_5638,N_5087);
xnor U8483 (N_8483,N_7084,N_6825);
and U8484 (N_8484,N_7274,N_6887);
nand U8485 (N_8485,N_5106,N_5509);
or U8486 (N_8486,N_5090,N_7492);
and U8487 (N_8487,N_7348,N_7307);
nor U8488 (N_8488,N_5134,N_6674);
and U8489 (N_8489,N_6376,N_5026);
nor U8490 (N_8490,N_7446,N_5222);
and U8491 (N_8491,N_7152,N_5538);
xnor U8492 (N_8492,N_5166,N_7161);
nor U8493 (N_8493,N_6681,N_7325);
and U8494 (N_8494,N_6747,N_6771);
nor U8495 (N_8495,N_5416,N_5105);
nor U8496 (N_8496,N_7289,N_5882);
xnor U8497 (N_8497,N_5360,N_5343);
nand U8498 (N_8498,N_6809,N_7482);
and U8499 (N_8499,N_5267,N_5299);
xor U8500 (N_8500,N_6650,N_6440);
or U8501 (N_8501,N_6688,N_5793);
xnor U8502 (N_8502,N_5820,N_6714);
nor U8503 (N_8503,N_6251,N_7214);
or U8504 (N_8504,N_5379,N_5775);
or U8505 (N_8505,N_6689,N_6664);
nor U8506 (N_8506,N_7058,N_5201);
nand U8507 (N_8507,N_6352,N_7135);
nand U8508 (N_8508,N_5558,N_5022);
xnor U8509 (N_8509,N_5549,N_5112);
nand U8510 (N_8510,N_6287,N_6525);
nand U8511 (N_8511,N_5583,N_5810);
xor U8512 (N_8512,N_5059,N_6187);
nand U8513 (N_8513,N_5779,N_7444);
and U8514 (N_8514,N_7443,N_6634);
and U8515 (N_8515,N_7103,N_6087);
nor U8516 (N_8516,N_7109,N_6890);
and U8517 (N_8517,N_6786,N_6743);
and U8518 (N_8518,N_5181,N_5935);
or U8519 (N_8519,N_6197,N_6692);
and U8520 (N_8520,N_5387,N_5931);
nor U8521 (N_8521,N_5998,N_5001);
nand U8522 (N_8522,N_6829,N_5889);
nand U8523 (N_8523,N_6923,N_5792);
nor U8524 (N_8524,N_6455,N_5868);
xnor U8525 (N_8525,N_6564,N_5940);
nand U8526 (N_8526,N_6815,N_6931);
xnor U8527 (N_8527,N_6949,N_6793);
nand U8528 (N_8528,N_6321,N_5369);
xnor U8529 (N_8529,N_6675,N_7421);
and U8530 (N_8530,N_5854,N_6763);
or U8531 (N_8531,N_6729,N_7417);
nor U8532 (N_8532,N_6820,N_5903);
and U8533 (N_8533,N_5004,N_7078);
nand U8534 (N_8534,N_5279,N_5253);
and U8535 (N_8535,N_5294,N_6891);
nor U8536 (N_8536,N_7321,N_7437);
and U8537 (N_8537,N_6502,N_6510);
nand U8538 (N_8538,N_5812,N_7143);
or U8539 (N_8539,N_5873,N_6183);
xor U8540 (N_8540,N_7265,N_5458);
or U8541 (N_8541,N_5396,N_5737);
and U8542 (N_8542,N_5427,N_7438);
and U8543 (N_8543,N_5135,N_6758);
or U8544 (N_8544,N_7499,N_6968);
or U8545 (N_8545,N_5554,N_6642);
or U8546 (N_8546,N_5374,N_5223);
and U8547 (N_8547,N_6944,N_6180);
nand U8548 (N_8548,N_5429,N_5036);
and U8549 (N_8549,N_6062,N_5592);
or U8550 (N_8550,N_7065,N_6335);
nor U8551 (N_8551,N_5972,N_5722);
and U8552 (N_8552,N_5675,N_5702);
nor U8553 (N_8553,N_6746,N_5119);
and U8554 (N_8554,N_6203,N_6429);
and U8555 (N_8555,N_5055,N_6051);
or U8556 (N_8556,N_7250,N_6059);
or U8557 (N_8557,N_6088,N_5115);
nand U8558 (N_8558,N_5981,N_5286);
xnor U8559 (N_8559,N_7029,N_6653);
nor U8560 (N_8560,N_6145,N_5123);
or U8561 (N_8561,N_7334,N_5333);
nor U8562 (N_8562,N_5184,N_6304);
nand U8563 (N_8563,N_5845,N_5602);
nor U8564 (N_8564,N_7064,N_5639);
or U8565 (N_8565,N_5478,N_6780);
nand U8566 (N_8566,N_7193,N_7196);
or U8567 (N_8567,N_6353,N_5330);
or U8568 (N_8568,N_6348,N_5607);
or U8569 (N_8569,N_6462,N_5621);
nand U8570 (N_8570,N_6052,N_6777);
and U8571 (N_8571,N_5185,N_6343);
or U8572 (N_8572,N_7162,N_6851);
nand U8573 (N_8573,N_6934,N_6811);
xnor U8574 (N_8574,N_5582,N_5718);
or U8575 (N_8575,N_6801,N_5720);
nor U8576 (N_8576,N_5104,N_7338);
or U8577 (N_8577,N_7478,N_6093);
and U8578 (N_8578,N_7174,N_6539);
nand U8579 (N_8579,N_7399,N_7264);
nand U8580 (N_8580,N_5958,N_6723);
nor U8581 (N_8581,N_6441,N_7070);
nand U8582 (N_8582,N_5939,N_5564);
or U8583 (N_8583,N_6575,N_5640);
or U8584 (N_8584,N_7106,N_7246);
nor U8585 (N_8585,N_7224,N_6079);
or U8586 (N_8586,N_5896,N_6986);
and U8587 (N_8587,N_6724,N_6213);
or U8588 (N_8588,N_6164,N_6340);
nor U8589 (N_8589,N_5758,N_5309);
nand U8590 (N_8590,N_6434,N_5130);
nor U8591 (N_8591,N_5671,N_5144);
nor U8592 (N_8592,N_7343,N_5986);
xnor U8593 (N_8593,N_5242,N_5287);
nor U8594 (N_8594,N_5766,N_5088);
and U8595 (N_8595,N_6275,N_5397);
and U8596 (N_8596,N_6875,N_6405);
nand U8597 (N_8597,N_5636,N_5193);
xnor U8598 (N_8598,N_5597,N_7030);
nor U8599 (N_8599,N_7032,N_7247);
nand U8600 (N_8600,N_5902,N_5832);
nor U8601 (N_8601,N_5472,N_6300);
or U8602 (N_8602,N_7201,N_5933);
or U8603 (N_8603,N_5635,N_6107);
nor U8604 (N_8604,N_7223,N_7062);
or U8605 (N_8605,N_6812,N_7203);
or U8606 (N_8606,N_6402,N_6411);
nor U8607 (N_8607,N_7189,N_5295);
nor U8608 (N_8608,N_5545,N_7294);
nor U8609 (N_8609,N_6542,N_7474);
and U8610 (N_8610,N_5382,N_5263);
nand U8611 (N_8611,N_6523,N_6424);
nor U8612 (N_8612,N_6936,N_6713);
or U8613 (N_8613,N_5094,N_5605);
or U8614 (N_8614,N_5411,N_6015);
or U8615 (N_8615,N_5761,N_6116);
nor U8616 (N_8616,N_6830,N_6274);
nand U8617 (N_8617,N_7447,N_7086);
and U8618 (N_8618,N_5131,N_7370);
and U8619 (N_8619,N_5529,N_5907);
and U8620 (N_8620,N_6271,N_7171);
and U8621 (N_8621,N_6419,N_5085);
nor U8622 (N_8622,N_6190,N_6698);
nand U8623 (N_8623,N_6857,N_5083);
nor U8624 (N_8624,N_6982,N_5344);
nand U8625 (N_8625,N_5437,N_6491);
and U8626 (N_8626,N_5292,N_7430);
nand U8627 (N_8627,N_7418,N_5156);
or U8628 (N_8628,N_5038,N_6727);
nor U8629 (N_8629,N_5249,N_6349);
xor U8630 (N_8630,N_5154,N_5034);
nand U8631 (N_8631,N_7244,N_5132);
nor U8632 (N_8632,N_5473,N_6856);
nand U8633 (N_8633,N_5606,N_6500);
nor U8634 (N_8634,N_5519,N_5164);
nand U8635 (N_8635,N_7082,N_7392);
nand U8636 (N_8636,N_7006,N_6006);
nand U8637 (N_8637,N_6527,N_6973);
or U8638 (N_8638,N_5162,N_5866);
nor U8639 (N_8639,N_6963,N_6555);
and U8640 (N_8640,N_5035,N_7373);
nor U8641 (N_8641,N_7220,N_6005);
or U8642 (N_8642,N_6091,N_5527);
and U8643 (N_8643,N_5765,N_6498);
nor U8644 (N_8644,N_6026,N_6897);
nor U8645 (N_8645,N_7270,N_6881);
nor U8646 (N_8646,N_5311,N_6528);
and U8647 (N_8647,N_6068,N_7306);
nand U8648 (N_8648,N_5598,N_6610);
nand U8649 (N_8649,N_6298,N_5364);
xnor U8650 (N_8650,N_7281,N_5296);
nor U8651 (N_8651,N_6950,N_7372);
xnor U8652 (N_8652,N_5649,N_5504);
or U8653 (N_8653,N_7359,N_6765);
nor U8654 (N_8654,N_6592,N_5269);
nor U8655 (N_8655,N_6373,N_6230);
nand U8656 (N_8656,N_6517,N_7081);
or U8657 (N_8657,N_5874,N_7026);
nor U8658 (N_8658,N_6778,N_6265);
and U8659 (N_8659,N_6325,N_5710);
nor U8660 (N_8660,N_5108,N_5282);
nor U8661 (N_8661,N_7356,N_5167);
or U8662 (N_8662,N_6902,N_5195);
nand U8663 (N_8663,N_6018,N_6264);
nand U8664 (N_8664,N_6682,N_7290);
nor U8665 (N_8665,N_6960,N_5624);
or U8666 (N_8666,N_6210,N_6599);
and U8667 (N_8667,N_7101,N_6022);
or U8668 (N_8668,N_7302,N_7148);
nand U8669 (N_8669,N_6465,N_6354);
or U8670 (N_8670,N_5136,N_7052);
nor U8671 (N_8671,N_5913,N_6757);
nor U8672 (N_8672,N_7151,N_5208);
or U8673 (N_8673,N_5789,N_5491);
nor U8674 (N_8674,N_6593,N_6864);
and U8675 (N_8675,N_5450,N_7073);
or U8676 (N_8676,N_7353,N_5909);
nor U8677 (N_8677,N_6054,N_5241);
nor U8678 (N_8678,N_6597,N_5047);
nor U8679 (N_8679,N_5356,N_7186);
or U8680 (N_8680,N_6383,N_6144);
nor U8681 (N_8681,N_5787,N_7227);
nand U8682 (N_8682,N_6961,N_7122);
xor U8683 (N_8683,N_5068,N_6587);
nor U8684 (N_8684,N_6388,N_6774);
xnor U8685 (N_8685,N_6676,N_6415);
nor U8686 (N_8686,N_5075,N_5305);
nor U8687 (N_8687,N_5659,N_5073);
nor U8688 (N_8688,N_5314,N_6075);
or U8689 (N_8689,N_6892,N_5814);
or U8690 (N_8690,N_5795,N_5357);
and U8691 (N_8691,N_7346,N_7124);
xor U8692 (N_8692,N_6594,N_6885);
nor U8693 (N_8693,N_5359,N_5401);
nor U8694 (N_8694,N_7300,N_5992);
nor U8695 (N_8695,N_7316,N_7097);
and U8696 (N_8696,N_6056,N_5321);
or U8697 (N_8697,N_5327,N_6627);
or U8698 (N_8698,N_6044,N_6492);
xnor U8699 (N_8699,N_6810,N_7494);
nor U8700 (N_8700,N_6481,N_7050);
xnor U8701 (N_8701,N_7401,N_5740);
nor U8702 (N_8702,N_6414,N_5265);
and U8703 (N_8703,N_5501,N_6010);
nand U8704 (N_8704,N_6802,N_6301);
or U8705 (N_8705,N_6859,N_6194);
and U8706 (N_8706,N_7260,N_6452);
and U8707 (N_8707,N_7259,N_5685);
nor U8708 (N_8708,N_5497,N_6629);
nand U8709 (N_8709,N_6508,N_5781);
nand U8710 (N_8710,N_5023,N_5928);
nand U8711 (N_8711,N_7228,N_5293);
nor U8712 (N_8712,N_5952,N_7146);
and U8713 (N_8713,N_6828,N_7022);
and U8714 (N_8714,N_7309,N_6457);
nor U8715 (N_8715,N_6485,N_5818);
or U8716 (N_8716,N_5961,N_6985);
nand U8717 (N_8717,N_7311,N_5834);
nor U8718 (N_8718,N_6220,N_5375);
nor U8719 (N_8719,N_5051,N_5225);
nor U8720 (N_8720,N_7286,N_5039);
nor U8721 (N_8721,N_6762,N_7479);
xnor U8722 (N_8722,N_5895,N_6377);
or U8723 (N_8723,N_5479,N_5078);
nor U8724 (N_8724,N_5220,N_5300);
and U8725 (N_8725,N_6232,N_6467);
nand U8726 (N_8726,N_5706,N_5719);
or U8727 (N_8727,N_6524,N_6937);
nor U8728 (N_8728,N_5213,N_6531);
or U8729 (N_8729,N_7393,N_7317);
nor U8730 (N_8730,N_6035,N_5861);
nor U8731 (N_8731,N_7419,N_6408);
nand U8732 (N_8732,N_6169,N_7411);
and U8733 (N_8733,N_5202,N_6805);
nand U8734 (N_8734,N_6160,N_5503);
nand U8735 (N_8735,N_6695,N_5484);
or U8736 (N_8736,N_7142,N_6261);
and U8737 (N_8737,N_5481,N_6489);
nor U8738 (N_8738,N_6198,N_6495);
and U8739 (N_8739,N_5946,N_7236);
nor U8740 (N_8740,N_5170,N_6540);
nand U8741 (N_8741,N_5796,N_5421);
nor U8742 (N_8742,N_6469,N_6247);
xor U8743 (N_8743,N_5150,N_6911);
and U8744 (N_8744,N_6456,N_7112);
nor U8745 (N_8745,N_6788,N_7428);
and U8746 (N_8746,N_5358,N_6559);
and U8747 (N_8747,N_5177,N_5975);
nand U8748 (N_8748,N_6333,N_5466);
and U8749 (N_8749,N_7156,N_5345);
nand U8750 (N_8750,N_7282,N_5765);
nand U8751 (N_8751,N_5850,N_6536);
and U8752 (N_8752,N_7125,N_5607);
and U8753 (N_8753,N_5878,N_6937);
nor U8754 (N_8754,N_6773,N_5488);
or U8755 (N_8755,N_6516,N_5495);
and U8756 (N_8756,N_5023,N_7442);
and U8757 (N_8757,N_7077,N_6595);
nor U8758 (N_8758,N_7391,N_7435);
nor U8759 (N_8759,N_7088,N_7466);
nand U8760 (N_8760,N_6506,N_5258);
or U8761 (N_8761,N_5711,N_5044);
xnor U8762 (N_8762,N_7303,N_5393);
and U8763 (N_8763,N_7402,N_5255);
nand U8764 (N_8764,N_5261,N_5522);
and U8765 (N_8765,N_5705,N_6395);
nand U8766 (N_8766,N_6254,N_7364);
nor U8767 (N_8767,N_7067,N_6554);
xnor U8768 (N_8768,N_6645,N_5550);
nor U8769 (N_8769,N_7474,N_5743);
xnor U8770 (N_8770,N_5335,N_5003);
nand U8771 (N_8771,N_7198,N_6222);
or U8772 (N_8772,N_6013,N_5693);
xor U8773 (N_8773,N_6136,N_5302);
nor U8774 (N_8774,N_6743,N_5134);
nand U8775 (N_8775,N_6470,N_5125);
nand U8776 (N_8776,N_6810,N_5092);
or U8777 (N_8777,N_6460,N_6070);
or U8778 (N_8778,N_5643,N_6925);
xor U8779 (N_8779,N_5278,N_6327);
nand U8780 (N_8780,N_5243,N_7443);
nor U8781 (N_8781,N_6628,N_7020);
nand U8782 (N_8782,N_5415,N_5466);
nor U8783 (N_8783,N_6717,N_7368);
nand U8784 (N_8784,N_5821,N_6407);
nand U8785 (N_8785,N_6768,N_5582);
nand U8786 (N_8786,N_6244,N_7090);
nand U8787 (N_8787,N_6501,N_6454);
or U8788 (N_8788,N_7394,N_5264);
nor U8789 (N_8789,N_5195,N_7334);
and U8790 (N_8790,N_5671,N_7428);
nand U8791 (N_8791,N_6511,N_6148);
nand U8792 (N_8792,N_6958,N_5011);
and U8793 (N_8793,N_6482,N_5650);
and U8794 (N_8794,N_7101,N_6949);
nand U8795 (N_8795,N_6748,N_5844);
nand U8796 (N_8796,N_5614,N_6115);
xor U8797 (N_8797,N_6029,N_5853);
nand U8798 (N_8798,N_6303,N_5487);
nor U8799 (N_8799,N_5297,N_7443);
nand U8800 (N_8800,N_7180,N_5541);
and U8801 (N_8801,N_7317,N_7407);
nand U8802 (N_8802,N_6170,N_7148);
or U8803 (N_8803,N_6649,N_6129);
or U8804 (N_8804,N_6349,N_6653);
or U8805 (N_8805,N_7455,N_5146);
nand U8806 (N_8806,N_6563,N_6087);
xnor U8807 (N_8807,N_6334,N_7308);
nor U8808 (N_8808,N_7189,N_6098);
nand U8809 (N_8809,N_5885,N_5447);
nor U8810 (N_8810,N_7009,N_6178);
or U8811 (N_8811,N_6990,N_5311);
xnor U8812 (N_8812,N_6618,N_7027);
xor U8813 (N_8813,N_6385,N_6016);
and U8814 (N_8814,N_6884,N_5118);
and U8815 (N_8815,N_6740,N_7337);
nor U8816 (N_8816,N_6655,N_5960);
and U8817 (N_8817,N_7329,N_7363);
nand U8818 (N_8818,N_5274,N_5559);
nor U8819 (N_8819,N_7419,N_6072);
or U8820 (N_8820,N_5939,N_7171);
nand U8821 (N_8821,N_5461,N_6523);
or U8822 (N_8822,N_5151,N_6607);
nand U8823 (N_8823,N_7097,N_6757);
nand U8824 (N_8824,N_6972,N_7390);
nor U8825 (N_8825,N_5618,N_5546);
nor U8826 (N_8826,N_6050,N_7284);
nor U8827 (N_8827,N_7253,N_5193);
nor U8828 (N_8828,N_5188,N_7441);
or U8829 (N_8829,N_5403,N_5835);
nor U8830 (N_8830,N_6660,N_7192);
or U8831 (N_8831,N_5699,N_6579);
nor U8832 (N_8832,N_6114,N_6452);
nor U8833 (N_8833,N_6012,N_5648);
and U8834 (N_8834,N_6850,N_5506);
nand U8835 (N_8835,N_6952,N_6984);
or U8836 (N_8836,N_7057,N_5897);
or U8837 (N_8837,N_6025,N_5597);
or U8838 (N_8838,N_6648,N_5617);
nand U8839 (N_8839,N_5225,N_7276);
nor U8840 (N_8840,N_5428,N_5632);
nand U8841 (N_8841,N_5221,N_5491);
and U8842 (N_8842,N_6062,N_6366);
nand U8843 (N_8843,N_5033,N_7219);
or U8844 (N_8844,N_7212,N_6927);
and U8845 (N_8845,N_7190,N_5543);
or U8846 (N_8846,N_5785,N_5236);
nor U8847 (N_8847,N_5997,N_5570);
xnor U8848 (N_8848,N_6370,N_5939);
nor U8849 (N_8849,N_5221,N_6963);
nor U8850 (N_8850,N_5881,N_5107);
xor U8851 (N_8851,N_5936,N_7032);
or U8852 (N_8852,N_5705,N_7454);
nand U8853 (N_8853,N_5249,N_5100);
or U8854 (N_8854,N_5262,N_6310);
or U8855 (N_8855,N_5874,N_7405);
and U8856 (N_8856,N_7437,N_6160);
nand U8857 (N_8857,N_7344,N_6377);
and U8858 (N_8858,N_6910,N_5411);
nor U8859 (N_8859,N_6857,N_6259);
or U8860 (N_8860,N_5928,N_6592);
and U8861 (N_8861,N_6429,N_5538);
and U8862 (N_8862,N_6680,N_7072);
nand U8863 (N_8863,N_7158,N_6854);
and U8864 (N_8864,N_6516,N_5556);
and U8865 (N_8865,N_7455,N_5790);
nand U8866 (N_8866,N_5819,N_5556);
and U8867 (N_8867,N_6402,N_5016);
nor U8868 (N_8868,N_6999,N_6829);
or U8869 (N_8869,N_6225,N_7252);
xor U8870 (N_8870,N_6009,N_7102);
or U8871 (N_8871,N_5389,N_7052);
or U8872 (N_8872,N_5356,N_6862);
nand U8873 (N_8873,N_6221,N_6078);
nor U8874 (N_8874,N_6507,N_5871);
nand U8875 (N_8875,N_6683,N_5834);
xnor U8876 (N_8876,N_5686,N_7407);
nor U8877 (N_8877,N_6985,N_6701);
or U8878 (N_8878,N_7350,N_6285);
or U8879 (N_8879,N_6478,N_6121);
and U8880 (N_8880,N_6057,N_5073);
or U8881 (N_8881,N_7341,N_5880);
nor U8882 (N_8882,N_6978,N_6264);
nand U8883 (N_8883,N_7460,N_7200);
nor U8884 (N_8884,N_7176,N_5693);
nand U8885 (N_8885,N_6828,N_7085);
nor U8886 (N_8886,N_6786,N_7006);
and U8887 (N_8887,N_6569,N_6880);
nor U8888 (N_8888,N_5943,N_6145);
or U8889 (N_8889,N_7152,N_7288);
nor U8890 (N_8890,N_6860,N_6309);
nand U8891 (N_8891,N_6367,N_7268);
nand U8892 (N_8892,N_6085,N_5800);
and U8893 (N_8893,N_5688,N_6586);
nor U8894 (N_8894,N_5007,N_5414);
nand U8895 (N_8895,N_6794,N_7083);
nor U8896 (N_8896,N_5144,N_5757);
nor U8897 (N_8897,N_5660,N_5021);
nor U8898 (N_8898,N_5670,N_6827);
nand U8899 (N_8899,N_6249,N_5543);
xor U8900 (N_8900,N_7096,N_6806);
nor U8901 (N_8901,N_6867,N_5470);
xnor U8902 (N_8902,N_6321,N_5276);
nand U8903 (N_8903,N_7457,N_5764);
and U8904 (N_8904,N_5504,N_7492);
or U8905 (N_8905,N_6533,N_6895);
nand U8906 (N_8906,N_5634,N_6811);
nor U8907 (N_8907,N_6290,N_5218);
nand U8908 (N_8908,N_5423,N_5424);
nor U8909 (N_8909,N_5965,N_7094);
and U8910 (N_8910,N_6951,N_6435);
or U8911 (N_8911,N_6133,N_7453);
and U8912 (N_8912,N_5148,N_7044);
and U8913 (N_8913,N_5812,N_6483);
nand U8914 (N_8914,N_5269,N_5877);
nand U8915 (N_8915,N_6180,N_6594);
nor U8916 (N_8916,N_6722,N_6021);
nand U8917 (N_8917,N_6235,N_5836);
xor U8918 (N_8918,N_5857,N_5836);
nor U8919 (N_8919,N_6544,N_7096);
and U8920 (N_8920,N_5497,N_6368);
and U8921 (N_8921,N_5958,N_6537);
nor U8922 (N_8922,N_5841,N_6082);
nand U8923 (N_8923,N_5093,N_7013);
or U8924 (N_8924,N_5083,N_7145);
and U8925 (N_8925,N_5123,N_5280);
nor U8926 (N_8926,N_6658,N_7324);
or U8927 (N_8927,N_5738,N_7351);
nand U8928 (N_8928,N_5035,N_5060);
or U8929 (N_8929,N_6503,N_5395);
or U8930 (N_8930,N_6657,N_5533);
nor U8931 (N_8931,N_6464,N_5434);
or U8932 (N_8932,N_5639,N_7370);
or U8933 (N_8933,N_7278,N_6624);
or U8934 (N_8934,N_7493,N_5152);
and U8935 (N_8935,N_5452,N_5743);
nand U8936 (N_8936,N_6518,N_6749);
xnor U8937 (N_8937,N_7198,N_5428);
nor U8938 (N_8938,N_5828,N_5211);
and U8939 (N_8939,N_5050,N_6028);
xor U8940 (N_8940,N_5748,N_5430);
and U8941 (N_8941,N_6265,N_7385);
nor U8942 (N_8942,N_5716,N_7442);
and U8943 (N_8943,N_6912,N_6248);
or U8944 (N_8944,N_6221,N_6442);
and U8945 (N_8945,N_5798,N_5634);
or U8946 (N_8946,N_6844,N_7264);
and U8947 (N_8947,N_7237,N_6496);
nand U8948 (N_8948,N_6601,N_5807);
or U8949 (N_8949,N_6602,N_5924);
and U8950 (N_8950,N_5001,N_7249);
nand U8951 (N_8951,N_6020,N_6607);
nor U8952 (N_8952,N_5207,N_5077);
and U8953 (N_8953,N_6690,N_5500);
or U8954 (N_8954,N_6305,N_6397);
nand U8955 (N_8955,N_5122,N_5459);
nor U8956 (N_8956,N_6246,N_6545);
nand U8957 (N_8957,N_7330,N_6141);
nor U8958 (N_8958,N_6661,N_7077);
nor U8959 (N_8959,N_5142,N_6699);
xor U8960 (N_8960,N_5692,N_6863);
nor U8961 (N_8961,N_6204,N_7486);
and U8962 (N_8962,N_6736,N_7473);
and U8963 (N_8963,N_6971,N_5059);
nor U8964 (N_8964,N_5714,N_6951);
nand U8965 (N_8965,N_6320,N_7460);
nand U8966 (N_8966,N_6014,N_6375);
and U8967 (N_8967,N_5509,N_6587);
nand U8968 (N_8968,N_5846,N_6331);
and U8969 (N_8969,N_5990,N_6482);
nor U8970 (N_8970,N_7355,N_7146);
or U8971 (N_8971,N_5087,N_6937);
nor U8972 (N_8972,N_6450,N_6333);
xor U8973 (N_8973,N_5835,N_5008);
and U8974 (N_8974,N_7499,N_6498);
or U8975 (N_8975,N_6282,N_6097);
nor U8976 (N_8976,N_6276,N_5105);
xnor U8977 (N_8977,N_7317,N_6729);
nand U8978 (N_8978,N_7075,N_7165);
nand U8979 (N_8979,N_7013,N_7039);
nor U8980 (N_8980,N_6784,N_5464);
or U8981 (N_8981,N_7334,N_6954);
and U8982 (N_8982,N_6592,N_5248);
nor U8983 (N_8983,N_6106,N_5924);
and U8984 (N_8984,N_5057,N_7461);
or U8985 (N_8985,N_5302,N_5827);
and U8986 (N_8986,N_6129,N_5569);
or U8987 (N_8987,N_7423,N_5096);
xor U8988 (N_8988,N_6635,N_5849);
xnor U8989 (N_8989,N_7389,N_5860);
nor U8990 (N_8990,N_6255,N_6102);
or U8991 (N_8991,N_7097,N_5953);
and U8992 (N_8992,N_5954,N_6280);
nand U8993 (N_8993,N_5548,N_6944);
nand U8994 (N_8994,N_5675,N_5923);
and U8995 (N_8995,N_5998,N_6132);
or U8996 (N_8996,N_6153,N_5087);
nor U8997 (N_8997,N_6189,N_5683);
and U8998 (N_8998,N_6044,N_6602);
and U8999 (N_8999,N_5466,N_6385);
or U9000 (N_9000,N_5339,N_5623);
and U9001 (N_9001,N_6045,N_5304);
or U9002 (N_9002,N_6171,N_5478);
or U9003 (N_9003,N_5646,N_5883);
or U9004 (N_9004,N_6267,N_5447);
or U9005 (N_9005,N_6297,N_5747);
nor U9006 (N_9006,N_6592,N_6376);
nor U9007 (N_9007,N_5589,N_7262);
nand U9008 (N_9008,N_6854,N_5949);
nand U9009 (N_9009,N_6557,N_7342);
nor U9010 (N_9010,N_5170,N_5423);
nand U9011 (N_9011,N_5779,N_5318);
nor U9012 (N_9012,N_5786,N_5686);
xor U9013 (N_9013,N_6575,N_5688);
and U9014 (N_9014,N_5684,N_5911);
nand U9015 (N_9015,N_6584,N_5430);
or U9016 (N_9016,N_7016,N_7351);
nor U9017 (N_9017,N_6965,N_7492);
or U9018 (N_9018,N_6975,N_7091);
or U9019 (N_9019,N_7402,N_7025);
and U9020 (N_9020,N_6802,N_6590);
xor U9021 (N_9021,N_6197,N_6797);
and U9022 (N_9022,N_6279,N_6340);
and U9023 (N_9023,N_7202,N_5730);
nand U9024 (N_9024,N_5088,N_5029);
or U9025 (N_9025,N_5208,N_5713);
nand U9026 (N_9026,N_6154,N_5075);
or U9027 (N_9027,N_7103,N_6538);
and U9028 (N_9028,N_6355,N_5416);
or U9029 (N_9029,N_5791,N_6804);
nor U9030 (N_9030,N_6950,N_5663);
nand U9031 (N_9031,N_5013,N_5859);
nand U9032 (N_9032,N_6961,N_6852);
nor U9033 (N_9033,N_6096,N_5989);
and U9034 (N_9034,N_6563,N_7239);
and U9035 (N_9035,N_6778,N_6185);
xor U9036 (N_9036,N_7354,N_6969);
nand U9037 (N_9037,N_6954,N_5199);
or U9038 (N_9038,N_6146,N_7329);
or U9039 (N_9039,N_7096,N_6225);
nor U9040 (N_9040,N_5891,N_6570);
nand U9041 (N_9041,N_7284,N_7184);
or U9042 (N_9042,N_5382,N_6795);
xor U9043 (N_9043,N_5880,N_6504);
and U9044 (N_9044,N_5321,N_6161);
and U9045 (N_9045,N_7327,N_6759);
and U9046 (N_9046,N_5468,N_5272);
or U9047 (N_9047,N_6120,N_5770);
nor U9048 (N_9048,N_6817,N_7324);
xor U9049 (N_9049,N_5066,N_6595);
nand U9050 (N_9050,N_5630,N_5205);
nor U9051 (N_9051,N_5783,N_6479);
xor U9052 (N_9052,N_5493,N_7267);
nand U9053 (N_9053,N_6671,N_5736);
and U9054 (N_9054,N_5563,N_5150);
nand U9055 (N_9055,N_5938,N_5720);
nand U9056 (N_9056,N_7406,N_6853);
or U9057 (N_9057,N_6330,N_5969);
or U9058 (N_9058,N_5097,N_6491);
nor U9059 (N_9059,N_6783,N_7325);
nand U9060 (N_9060,N_5538,N_5555);
nand U9061 (N_9061,N_6629,N_6257);
nor U9062 (N_9062,N_7135,N_5623);
and U9063 (N_9063,N_6504,N_5906);
and U9064 (N_9064,N_6230,N_7373);
and U9065 (N_9065,N_6072,N_7085);
and U9066 (N_9066,N_7406,N_5636);
or U9067 (N_9067,N_7429,N_5406);
xnor U9068 (N_9068,N_5470,N_5320);
or U9069 (N_9069,N_6874,N_7385);
and U9070 (N_9070,N_7226,N_6906);
or U9071 (N_9071,N_7422,N_5621);
and U9072 (N_9072,N_6576,N_6935);
nand U9073 (N_9073,N_6194,N_6799);
or U9074 (N_9074,N_7037,N_6575);
nand U9075 (N_9075,N_5013,N_6529);
nand U9076 (N_9076,N_6152,N_7488);
nor U9077 (N_9077,N_5497,N_5590);
nand U9078 (N_9078,N_7433,N_6442);
or U9079 (N_9079,N_6212,N_5788);
xor U9080 (N_9080,N_6063,N_6940);
nand U9081 (N_9081,N_5572,N_6759);
or U9082 (N_9082,N_5644,N_6631);
or U9083 (N_9083,N_5975,N_7413);
xnor U9084 (N_9084,N_5704,N_6469);
xor U9085 (N_9085,N_6951,N_5592);
or U9086 (N_9086,N_7357,N_6246);
and U9087 (N_9087,N_6169,N_7132);
nor U9088 (N_9088,N_5200,N_7364);
nand U9089 (N_9089,N_6118,N_6653);
or U9090 (N_9090,N_6030,N_5866);
nor U9091 (N_9091,N_7060,N_7364);
nor U9092 (N_9092,N_5422,N_6382);
and U9093 (N_9093,N_6971,N_6993);
or U9094 (N_9094,N_6111,N_6121);
nor U9095 (N_9095,N_6789,N_7341);
nor U9096 (N_9096,N_7245,N_7101);
nand U9097 (N_9097,N_5304,N_6890);
nor U9098 (N_9098,N_6515,N_6118);
and U9099 (N_9099,N_7099,N_5853);
nor U9100 (N_9100,N_5356,N_7305);
or U9101 (N_9101,N_7430,N_6969);
nor U9102 (N_9102,N_5607,N_7388);
nor U9103 (N_9103,N_5587,N_5093);
and U9104 (N_9104,N_7276,N_6791);
nor U9105 (N_9105,N_7197,N_7334);
xor U9106 (N_9106,N_7379,N_5655);
nor U9107 (N_9107,N_6015,N_5650);
nor U9108 (N_9108,N_7329,N_5489);
nor U9109 (N_9109,N_7058,N_6355);
or U9110 (N_9110,N_5241,N_7367);
xnor U9111 (N_9111,N_5806,N_7221);
or U9112 (N_9112,N_7023,N_6627);
or U9113 (N_9113,N_5509,N_5006);
or U9114 (N_9114,N_6658,N_7321);
nand U9115 (N_9115,N_7034,N_5873);
or U9116 (N_9116,N_7184,N_6239);
and U9117 (N_9117,N_6191,N_6329);
nor U9118 (N_9118,N_5951,N_5316);
and U9119 (N_9119,N_5886,N_5616);
or U9120 (N_9120,N_5137,N_7241);
or U9121 (N_9121,N_5619,N_5863);
or U9122 (N_9122,N_7284,N_5566);
nor U9123 (N_9123,N_5607,N_6901);
nand U9124 (N_9124,N_7483,N_6534);
nor U9125 (N_9125,N_5647,N_7310);
xnor U9126 (N_9126,N_7229,N_6824);
nand U9127 (N_9127,N_5346,N_6923);
and U9128 (N_9128,N_5683,N_5432);
or U9129 (N_9129,N_5741,N_6576);
xor U9130 (N_9130,N_6438,N_5349);
xor U9131 (N_9131,N_6296,N_7192);
or U9132 (N_9132,N_5083,N_5318);
nor U9133 (N_9133,N_5654,N_7479);
and U9134 (N_9134,N_6324,N_5698);
nand U9135 (N_9135,N_6186,N_6910);
nand U9136 (N_9136,N_5490,N_6963);
or U9137 (N_9137,N_5745,N_6195);
and U9138 (N_9138,N_6157,N_6407);
nor U9139 (N_9139,N_7318,N_7012);
nand U9140 (N_9140,N_5329,N_6094);
and U9141 (N_9141,N_5746,N_5547);
nand U9142 (N_9142,N_6135,N_6418);
or U9143 (N_9143,N_5396,N_5699);
or U9144 (N_9144,N_6294,N_6213);
nand U9145 (N_9145,N_7241,N_6316);
or U9146 (N_9146,N_7294,N_6998);
nand U9147 (N_9147,N_5838,N_7079);
nand U9148 (N_9148,N_7101,N_7094);
and U9149 (N_9149,N_5847,N_7314);
or U9150 (N_9150,N_5473,N_6154);
xnor U9151 (N_9151,N_6236,N_6895);
nor U9152 (N_9152,N_7320,N_5033);
or U9153 (N_9153,N_6140,N_7302);
nor U9154 (N_9154,N_6252,N_6690);
and U9155 (N_9155,N_6392,N_5340);
nor U9156 (N_9156,N_5080,N_5470);
or U9157 (N_9157,N_6915,N_5122);
or U9158 (N_9158,N_6114,N_6970);
nand U9159 (N_9159,N_5062,N_5781);
and U9160 (N_9160,N_6035,N_7096);
nor U9161 (N_9161,N_5803,N_5997);
nor U9162 (N_9162,N_6778,N_6423);
nor U9163 (N_9163,N_6311,N_5136);
or U9164 (N_9164,N_6032,N_6952);
and U9165 (N_9165,N_6068,N_7218);
nand U9166 (N_9166,N_5616,N_5084);
nand U9167 (N_9167,N_6156,N_7286);
nor U9168 (N_9168,N_6072,N_5477);
or U9169 (N_9169,N_5833,N_7313);
nand U9170 (N_9170,N_6248,N_6089);
nand U9171 (N_9171,N_7234,N_7261);
or U9172 (N_9172,N_6741,N_5183);
nor U9173 (N_9173,N_5097,N_6705);
nor U9174 (N_9174,N_7141,N_5386);
or U9175 (N_9175,N_6941,N_6488);
or U9176 (N_9176,N_6118,N_6419);
nand U9177 (N_9177,N_7211,N_6686);
nor U9178 (N_9178,N_7059,N_6117);
nor U9179 (N_9179,N_5557,N_5820);
nor U9180 (N_9180,N_5935,N_6530);
or U9181 (N_9181,N_5156,N_5229);
or U9182 (N_9182,N_5325,N_6402);
or U9183 (N_9183,N_7134,N_6920);
xor U9184 (N_9184,N_6842,N_5396);
or U9185 (N_9185,N_6240,N_5978);
or U9186 (N_9186,N_7368,N_7097);
nor U9187 (N_9187,N_7072,N_5790);
or U9188 (N_9188,N_5477,N_6463);
nand U9189 (N_9189,N_7447,N_5009);
nor U9190 (N_9190,N_6063,N_6943);
and U9191 (N_9191,N_5787,N_7126);
nand U9192 (N_9192,N_6670,N_5534);
nand U9193 (N_9193,N_5689,N_7062);
and U9194 (N_9194,N_5109,N_6944);
or U9195 (N_9195,N_6845,N_5571);
nand U9196 (N_9196,N_5550,N_6072);
and U9197 (N_9197,N_7434,N_5688);
nand U9198 (N_9198,N_5861,N_5361);
nand U9199 (N_9199,N_5639,N_5967);
nor U9200 (N_9200,N_5524,N_6379);
nor U9201 (N_9201,N_6595,N_7201);
and U9202 (N_9202,N_5520,N_5256);
and U9203 (N_9203,N_5544,N_6902);
nor U9204 (N_9204,N_6715,N_5522);
and U9205 (N_9205,N_6005,N_6341);
or U9206 (N_9206,N_6083,N_5111);
and U9207 (N_9207,N_6208,N_5294);
or U9208 (N_9208,N_6496,N_6323);
and U9209 (N_9209,N_6651,N_7206);
or U9210 (N_9210,N_7088,N_7398);
nand U9211 (N_9211,N_6984,N_6765);
nor U9212 (N_9212,N_6803,N_5360);
nor U9213 (N_9213,N_7210,N_5757);
or U9214 (N_9214,N_7075,N_6365);
or U9215 (N_9215,N_5990,N_7333);
and U9216 (N_9216,N_5699,N_5062);
nor U9217 (N_9217,N_7498,N_6731);
xor U9218 (N_9218,N_7167,N_5922);
nand U9219 (N_9219,N_6609,N_7317);
nand U9220 (N_9220,N_6974,N_5194);
nand U9221 (N_9221,N_6051,N_6950);
and U9222 (N_9222,N_6838,N_5955);
nand U9223 (N_9223,N_7359,N_6145);
nor U9224 (N_9224,N_5177,N_5384);
nand U9225 (N_9225,N_7321,N_5784);
nand U9226 (N_9226,N_6768,N_6536);
and U9227 (N_9227,N_6412,N_7029);
nor U9228 (N_9228,N_6246,N_6253);
or U9229 (N_9229,N_5569,N_6903);
or U9230 (N_9230,N_5079,N_5309);
nor U9231 (N_9231,N_5856,N_6870);
nor U9232 (N_9232,N_7045,N_6516);
nor U9233 (N_9233,N_7411,N_5634);
xnor U9234 (N_9234,N_5177,N_7485);
nand U9235 (N_9235,N_5483,N_7475);
nand U9236 (N_9236,N_5088,N_6280);
and U9237 (N_9237,N_6039,N_6988);
and U9238 (N_9238,N_6235,N_6263);
or U9239 (N_9239,N_7469,N_7367);
or U9240 (N_9240,N_5182,N_7438);
or U9241 (N_9241,N_5453,N_5251);
or U9242 (N_9242,N_5978,N_6611);
or U9243 (N_9243,N_6152,N_5352);
or U9244 (N_9244,N_6570,N_5108);
nor U9245 (N_9245,N_6805,N_5657);
nand U9246 (N_9246,N_6725,N_5987);
nand U9247 (N_9247,N_5737,N_6683);
xnor U9248 (N_9248,N_6502,N_6055);
nor U9249 (N_9249,N_6789,N_7301);
and U9250 (N_9250,N_6224,N_5463);
or U9251 (N_9251,N_6106,N_6296);
or U9252 (N_9252,N_6303,N_6736);
and U9253 (N_9253,N_5786,N_7459);
or U9254 (N_9254,N_5705,N_6160);
xor U9255 (N_9255,N_6683,N_5342);
nand U9256 (N_9256,N_7257,N_5349);
or U9257 (N_9257,N_5719,N_6442);
nor U9258 (N_9258,N_5854,N_6419);
and U9259 (N_9259,N_6968,N_5538);
nand U9260 (N_9260,N_5813,N_5391);
and U9261 (N_9261,N_7390,N_7176);
xnor U9262 (N_9262,N_7140,N_6333);
nor U9263 (N_9263,N_6594,N_7367);
nand U9264 (N_9264,N_7473,N_7210);
nand U9265 (N_9265,N_5823,N_6017);
xor U9266 (N_9266,N_6171,N_6359);
nand U9267 (N_9267,N_5730,N_7454);
xor U9268 (N_9268,N_6434,N_7071);
and U9269 (N_9269,N_6342,N_6938);
nand U9270 (N_9270,N_7154,N_6858);
and U9271 (N_9271,N_5925,N_5344);
nand U9272 (N_9272,N_7201,N_6038);
and U9273 (N_9273,N_6727,N_5650);
xnor U9274 (N_9274,N_6298,N_6153);
nor U9275 (N_9275,N_7414,N_6319);
xnor U9276 (N_9276,N_7215,N_7403);
nor U9277 (N_9277,N_7250,N_5046);
and U9278 (N_9278,N_6558,N_6576);
or U9279 (N_9279,N_6203,N_6431);
xnor U9280 (N_9280,N_5317,N_7307);
or U9281 (N_9281,N_6912,N_7366);
nand U9282 (N_9282,N_7354,N_6971);
and U9283 (N_9283,N_7213,N_5941);
nor U9284 (N_9284,N_5966,N_5713);
and U9285 (N_9285,N_5756,N_5775);
and U9286 (N_9286,N_6410,N_7226);
or U9287 (N_9287,N_7258,N_5450);
and U9288 (N_9288,N_7458,N_5235);
and U9289 (N_9289,N_6089,N_7347);
or U9290 (N_9290,N_5149,N_7360);
and U9291 (N_9291,N_7179,N_7459);
and U9292 (N_9292,N_7305,N_5408);
nor U9293 (N_9293,N_6727,N_5642);
nor U9294 (N_9294,N_6967,N_7186);
nor U9295 (N_9295,N_7400,N_7213);
nor U9296 (N_9296,N_6409,N_6736);
xnor U9297 (N_9297,N_6677,N_7197);
nand U9298 (N_9298,N_5526,N_7390);
or U9299 (N_9299,N_6687,N_7162);
xor U9300 (N_9300,N_6639,N_5979);
and U9301 (N_9301,N_5626,N_5796);
xnor U9302 (N_9302,N_6622,N_7167);
and U9303 (N_9303,N_7358,N_6562);
nand U9304 (N_9304,N_7100,N_7419);
nand U9305 (N_9305,N_6670,N_5917);
and U9306 (N_9306,N_6222,N_6288);
nor U9307 (N_9307,N_6070,N_6349);
and U9308 (N_9308,N_5811,N_7456);
xnor U9309 (N_9309,N_7466,N_7194);
xnor U9310 (N_9310,N_5192,N_5928);
nor U9311 (N_9311,N_5886,N_7123);
and U9312 (N_9312,N_5698,N_5686);
nor U9313 (N_9313,N_7317,N_6112);
nand U9314 (N_9314,N_7171,N_6517);
xnor U9315 (N_9315,N_6046,N_6178);
nor U9316 (N_9316,N_7366,N_5172);
nor U9317 (N_9317,N_5028,N_6567);
and U9318 (N_9318,N_6256,N_6988);
nand U9319 (N_9319,N_6873,N_5685);
or U9320 (N_9320,N_6222,N_5433);
or U9321 (N_9321,N_5526,N_5696);
nand U9322 (N_9322,N_5528,N_5705);
nand U9323 (N_9323,N_5155,N_6763);
or U9324 (N_9324,N_5906,N_6591);
nand U9325 (N_9325,N_7253,N_6378);
and U9326 (N_9326,N_5105,N_5290);
nor U9327 (N_9327,N_7259,N_5791);
nor U9328 (N_9328,N_5087,N_6555);
and U9329 (N_9329,N_7214,N_6419);
or U9330 (N_9330,N_5104,N_5308);
and U9331 (N_9331,N_7357,N_5614);
or U9332 (N_9332,N_5834,N_6616);
or U9333 (N_9333,N_5660,N_6110);
or U9334 (N_9334,N_6994,N_5407);
or U9335 (N_9335,N_5074,N_7357);
and U9336 (N_9336,N_5283,N_6783);
and U9337 (N_9337,N_6963,N_5762);
xor U9338 (N_9338,N_5608,N_5708);
or U9339 (N_9339,N_5047,N_5401);
or U9340 (N_9340,N_5651,N_5775);
nand U9341 (N_9341,N_6812,N_5144);
nor U9342 (N_9342,N_5450,N_7119);
nor U9343 (N_9343,N_5671,N_6881);
nor U9344 (N_9344,N_6401,N_6129);
xnor U9345 (N_9345,N_6192,N_5304);
and U9346 (N_9346,N_6049,N_7018);
xor U9347 (N_9347,N_7416,N_5038);
or U9348 (N_9348,N_5184,N_5309);
nor U9349 (N_9349,N_5154,N_7084);
nand U9350 (N_9350,N_6755,N_6394);
nor U9351 (N_9351,N_6984,N_6940);
nor U9352 (N_9352,N_5811,N_6016);
xor U9353 (N_9353,N_6138,N_6302);
nand U9354 (N_9354,N_6540,N_5788);
and U9355 (N_9355,N_6726,N_5241);
or U9356 (N_9356,N_6418,N_6946);
or U9357 (N_9357,N_7211,N_6546);
nor U9358 (N_9358,N_6378,N_5561);
nand U9359 (N_9359,N_6647,N_5883);
or U9360 (N_9360,N_5462,N_5143);
nand U9361 (N_9361,N_6750,N_5292);
nor U9362 (N_9362,N_5410,N_6711);
nor U9363 (N_9363,N_5290,N_5240);
and U9364 (N_9364,N_5135,N_5429);
nor U9365 (N_9365,N_6983,N_5102);
nor U9366 (N_9366,N_6843,N_5623);
and U9367 (N_9367,N_7298,N_5426);
or U9368 (N_9368,N_5972,N_6158);
xnor U9369 (N_9369,N_7073,N_7286);
xnor U9370 (N_9370,N_5114,N_7414);
xor U9371 (N_9371,N_6178,N_5540);
nor U9372 (N_9372,N_5954,N_6528);
xor U9373 (N_9373,N_6586,N_5864);
nand U9374 (N_9374,N_6214,N_6445);
or U9375 (N_9375,N_5850,N_6633);
or U9376 (N_9376,N_5510,N_6753);
nor U9377 (N_9377,N_7205,N_5950);
nand U9378 (N_9378,N_5606,N_6011);
or U9379 (N_9379,N_5933,N_6673);
nor U9380 (N_9380,N_6489,N_6787);
nand U9381 (N_9381,N_7011,N_5594);
nor U9382 (N_9382,N_7114,N_5547);
or U9383 (N_9383,N_6593,N_5522);
and U9384 (N_9384,N_5643,N_6040);
nor U9385 (N_9385,N_6379,N_5243);
nor U9386 (N_9386,N_7119,N_5297);
nor U9387 (N_9387,N_6287,N_5544);
and U9388 (N_9388,N_6381,N_7314);
nor U9389 (N_9389,N_5866,N_5905);
and U9390 (N_9390,N_6864,N_5409);
and U9391 (N_9391,N_5970,N_6113);
nand U9392 (N_9392,N_6393,N_5480);
and U9393 (N_9393,N_6188,N_5288);
nand U9394 (N_9394,N_6746,N_6072);
xnor U9395 (N_9395,N_5912,N_5823);
or U9396 (N_9396,N_5988,N_7374);
nor U9397 (N_9397,N_5007,N_6080);
nor U9398 (N_9398,N_6299,N_6784);
nand U9399 (N_9399,N_5864,N_6929);
xor U9400 (N_9400,N_7219,N_6624);
nor U9401 (N_9401,N_6562,N_6829);
or U9402 (N_9402,N_6893,N_5965);
nand U9403 (N_9403,N_5021,N_7036);
nand U9404 (N_9404,N_5615,N_7085);
and U9405 (N_9405,N_5532,N_6088);
and U9406 (N_9406,N_6253,N_6107);
and U9407 (N_9407,N_5587,N_5454);
or U9408 (N_9408,N_5623,N_6530);
nor U9409 (N_9409,N_5462,N_6853);
nor U9410 (N_9410,N_6290,N_7117);
nand U9411 (N_9411,N_5614,N_6064);
and U9412 (N_9412,N_5839,N_7305);
or U9413 (N_9413,N_6533,N_5280);
nor U9414 (N_9414,N_5136,N_6397);
nand U9415 (N_9415,N_6612,N_6382);
nand U9416 (N_9416,N_5919,N_6352);
and U9417 (N_9417,N_5138,N_6878);
nor U9418 (N_9418,N_6329,N_5554);
nor U9419 (N_9419,N_5275,N_5098);
or U9420 (N_9420,N_7268,N_7275);
or U9421 (N_9421,N_6393,N_5305);
or U9422 (N_9422,N_5492,N_7393);
nor U9423 (N_9423,N_7392,N_5834);
nand U9424 (N_9424,N_7366,N_5089);
xor U9425 (N_9425,N_6674,N_6704);
xnor U9426 (N_9426,N_6474,N_5865);
nor U9427 (N_9427,N_6119,N_6247);
nor U9428 (N_9428,N_7390,N_6237);
nor U9429 (N_9429,N_5361,N_7194);
nor U9430 (N_9430,N_5978,N_6762);
or U9431 (N_9431,N_5251,N_6980);
or U9432 (N_9432,N_6089,N_6027);
or U9433 (N_9433,N_6293,N_5549);
or U9434 (N_9434,N_6791,N_5909);
xnor U9435 (N_9435,N_6468,N_6551);
nor U9436 (N_9436,N_5779,N_7199);
xnor U9437 (N_9437,N_7408,N_6926);
nor U9438 (N_9438,N_6949,N_5704);
xnor U9439 (N_9439,N_6936,N_6779);
xnor U9440 (N_9440,N_7266,N_5368);
and U9441 (N_9441,N_6778,N_5867);
and U9442 (N_9442,N_5712,N_6554);
xnor U9443 (N_9443,N_6026,N_5545);
xor U9444 (N_9444,N_6573,N_7453);
or U9445 (N_9445,N_7497,N_7331);
or U9446 (N_9446,N_5609,N_6244);
or U9447 (N_9447,N_7360,N_7235);
nand U9448 (N_9448,N_6853,N_5697);
and U9449 (N_9449,N_5607,N_6997);
or U9450 (N_9450,N_5429,N_5022);
or U9451 (N_9451,N_7059,N_6617);
nand U9452 (N_9452,N_5276,N_6524);
nor U9453 (N_9453,N_6223,N_7334);
nor U9454 (N_9454,N_6383,N_5200);
xnor U9455 (N_9455,N_7222,N_5262);
nor U9456 (N_9456,N_5179,N_5779);
nand U9457 (N_9457,N_6576,N_5430);
and U9458 (N_9458,N_5090,N_5593);
nor U9459 (N_9459,N_5492,N_5555);
or U9460 (N_9460,N_7331,N_6580);
nand U9461 (N_9461,N_6389,N_5523);
nand U9462 (N_9462,N_6371,N_6157);
or U9463 (N_9463,N_6294,N_6755);
or U9464 (N_9464,N_6236,N_6342);
xnor U9465 (N_9465,N_6828,N_5345);
or U9466 (N_9466,N_6697,N_7462);
or U9467 (N_9467,N_7084,N_6290);
or U9468 (N_9468,N_7284,N_5733);
nand U9469 (N_9469,N_7289,N_6191);
and U9470 (N_9470,N_6519,N_6945);
or U9471 (N_9471,N_6142,N_5813);
nor U9472 (N_9472,N_7248,N_7114);
and U9473 (N_9473,N_6130,N_6529);
and U9474 (N_9474,N_6592,N_7280);
nand U9475 (N_9475,N_7477,N_6427);
or U9476 (N_9476,N_5918,N_6009);
xor U9477 (N_9477,N_6946,N_6419);
nand U9478 (N_9478,N_5877,N_6769);
nand U9479 (N_9479,N_6614,N_6254);
or U9480 (N_9480,N_6082,N_6882);
or U9481 (N_9481,N_7311,N_5185);
and U9482 (N_9482,N_6412,N_6267);
or U9483 (N_9483,N_5437,N_6900);
and U9484 (N_9484,N_5187,N_6013);
nand U9485 (N_9485,N_6187,N_5150);
nor U9486 (N_9486,N_5657,N_6196);
and U9487 (N_9487,N_5184,N_6845);
and U9488 (N_9488,N_7415,N_6746);
nand U9489 (N_9489,N_5757,N_6263);
nor U9490 (N_9490,N_6594,N_7495);
xnor U9491 (N_9491,N_7252,N_5101);
nand U9492 (N_9492,N_6802,N_6547);
nor U9493 (N_9493,N_5327,N_5475);
nand U9494 (N_9494,N_7235,N_5975);
or U9495 (N_9495,N_6836,N_6867);
or U9496 (N_9496,N_7016,N_6787);
and U9497 (N_9497,N_5170,N_5715);
or U9498 (N_9498,N_5975,N_6754);
or U9499 (N_9499,N_7122,N_5985);
nand U9500 (N_9500,N_5138,N_6058);
nand U9501 (N_9501,N_7380,N_5936);
or U9502 (N_9502,N_7441,N_5568);
nor U9503 (N_9503,N_5518,N_6699);
nand U9504 (N_9504,N_7044,N_5505);
and U9505 (N_9505,N_5403,N_5964);
xnor U9506 (N_9506,N_5757,N_5026);
and U9507 (N_9507,N_6667,N_6143);
or U9508 (N_9508,N_7034,N_5909);
and U9509 (N_9509,N_7471,N_6460);
nor U9510 (N_9510,N_5847,N_7244);
or U9511 (N_9511,N_7421,N_5406);
nor U9512 (N_9512,N_5889,N_7434);
nand U9513 (N_9513,N_5825,N_7390);
or U9514 (N_9514,N_7065,N_5490);
nand U9515 (N_9515,N_6657,N_7016);
and U9516 (N_9516,N_6191,N_7493);
or U9517 (N_9517,N_5175,N_5286);
or U9518 (N_9518,N_5550,N_5813);
nor U9519 (N_9519,N_5394,N_5416);
and U9520 (N_9520,N_6711,N_6996);
nand U9521 (N_9521,N_5935,N_6863);
and U9522 (N_9522,N_5813,N_5417);
nor U9523 (N_9523,N_6001,N_5463);
and U9524 (N_9524,N_5109,N_5501);
and U9525 (N_9525,N_6595,N_5929);
nor U9526 (N_9526,N_6953,N_5991);
nand U9527 (N_9527,N_5300,N_5562);
nor U9528 (N_9528,N_5715,N_6132);
nand U9529 (N_9529,N_5050,N_6487);
nor U9530 (N_9530,N_6105,N_5969);
and U9531 (N_9531,N_5857,N_5197);
or U9532 (N_9532,N_6686,N_5783);
or U9533 (N_9533,N_6402,N_5145);
nor U9534 (N_9534,N_6314,N_6227);
nand U9535 (N_9535,N_5784,N_5701);
nand U9536 (N_9536,N_7126,N_7144);
nor U9537 (N_9537,N_6360,N_5935);
or U9538 (N_9538,N_6323,N_6012);
nor U9539 (N_9539,N_6140,N_6875);
nor U9540 (N_9540,N_6414,N_7293);
or U9541 (N_9541,N_5619,N_5145);
xor U9542 (N_9542,N_6849,N_5942);
or U9543 (N_9543,N_5078,N_5149);
xnor U9544 (N_9544,N_5243,N_6174);
and U9545 (N_9545,N_6237,N_6671);
nor U9546 (N_9546,N_6694,N_6769);
or U9547 (N_9547,N_5148,N_6845);
and U9548 (N_9548,N_6535,N_7064);
xnor U9549 (N_9549,N_5390,N_5795);
or U9550 (N_9550,N_6153,N_7211);
and U9551 (N_9551,N_7154,N_5178);
nor U9552 (N_9552,N_5061,N_5923);
and U9553 (N_9553,N_6304,N_6894);
nor U9554 (N_9554,N_6202,N_5107);
nor U9555 (N_9555,N_6191,N_6093);
and U9556 (N_9556,N_5799,N_7445);
nand U9557 (N_9557,N_5539,N_6760);
nor U9558 (N_9558,N_7403,N_6386);
nor U9559 (N_9559,N_6092,N_7473);
or U9560 (N_9560,N_7454,N_6046);
and U9561 (N_9561,N_5209,N_5673);
nand U9562 (N_9562,N_6812,N_6747);
and U9563 (N_9563,N_6078,N_5531);
and U9564 (N_9564,N_6251,N_5502);
nor U9565 (N_9565,N_6302,N_6961);
and U9566 (N_9566,N_7337,N_6785);
or U9567 (N_9567,N_6687,N_5275);
or U9568 (N_9568,N_5710,N_6360);
or U9569 (N_9569,N_6668,N_7447);
or U9570 (N_9570,N_5301,N_7330);
nand U9571 (N_9571,N_5804,N_6596);
and U9572 (N_9572,N_6678,N_5568);
or U9573 (N_9573,N_5538,N_5492);
and U9574 (N_9574,N_6358,N_5681);
or U9575 (N_9575,N_5498,N_7190);
nor U9576 (N_9576,N_7250,N_7126);
nand U9577 (N_9577,N_5926,N_5852);
nand U9578 (N_9578,N_5356,N_7074);
and U9579 (N_9579,N_7287,N_6945);
and U9580 (N_9580,N_7184,N_6556);
and U9581 (N_9581,N_5969,N_6472);
or U9582 (N_9582,N_7278,N_6219);
and U9583 (N_9583,N_6731,N_6939);
nand U9584 (N_9584,N_5364,N_5736);
and U9585 (N_9585,N_6701,N_7035);
nor U9586 (N_9586,N_7432,N_5946);
nor U9587 (N_9587,N_6679,N_6696);
nand U9588 (N_9588,N_6096,N_5773);
or U9589 (N_9589,N_7147,N_5852);
or U9590 (N_9590,N_7360,N_5304);
xnor U9591 (N_9591,N_6533,N_5140);
nand U9592 (N_9592,N_6724,N_5505);
xnor U9593 (N_9593,N_5730,N_6072);
and U9594 (N_9594,N_5461,N_6953);
nand U9595 (N_9595,N_7017,N_5661);
or U9596 (N_9596,N_7062,N_7270);
and U9597 (N_9597,N_7135,N_6600);
and U9598 (N_9598,N_5403,N_7341);
nor U9599 (N_9599,N_5596,N_5449);
nand U9600 (N_9600,N_5812,N_5507);
or U9601 (N_9601,N_7425,N_5389);
xor U9602 (N_9602,N_5481,N_6879);
nor U9603 (N_9603,N_7401,N_5983);
nor U9604 (N_9604,N_7207,N_5043);
nand U9605 (N_9605,N_5598,N_6700);
nand U9606 (N_9606,N_5896,N_6584);
or U9607 (N_9607,N_6280,N_6008);
nand U9608 (N_9608,N_5641,N_7366);
or U9609 (N_9609,N_6051,N_6968);
and U9610 (N_9610,N_6611,N_7000);
nand U9611 (N_9611,N_7268,N_6994);
or U9612 (N_9612,N_6538,N_5182);
nand U9613 (N_9613,N_5537,N_6481);
nor U9614 (N_9614,N_7470,N_5403);
and U9615 (N_9615,N_6367,N_6443);
or U9616 (N_9616,N_6889,N_7038);
or U9617 (N_9617,N_5997,N_5386);
nand U9618 (N_9618,N_5016,N_6696);
and U9619 (N_9619,N_5825,N_6337);
nor U9620 (N_9620,N_5477,N_6811);
and U9621 (N_9621,N_5653,N_6851);
nand U9622 (N_9622,N_7355,N_6558);
and U9623 (N_9623,N_5093,N_7407);
nand U9624 (N_9624,N_7307,N_5789);
and U9625 (N_9625,N_6446,N_6348);
or U9626 (N_9626,N_6436,N_5158);
and U9627 (N_9627,N_6884,N_6379);
and U9628 (N_9628,N_5254,N_7466);
or U9629 (N_9629,N_5483,N_5378);
or U9630 (N_9630,N_7051,N_7266);
and U9631 (N_9631,N_6048,N_7029);
nand U9632 (N_9632,N_7229,N_5966);
xnor U9633 (N_9633,N_6045,N_5226);
nor U9634 (N_9634,N_6208,N_5120);
xnor U9635 (N_9635,N_6510,N_6231);
nand U9636 (N_9636,N_5353,N_5601);
nor U9637 (N_9637,N_5059,N_7348);
nand U9638 (N_9638,N_6352,N_6304);
nor U9639 (N_9639,N_5827,N_7473);
nand U9640 (N_9640,N_5960,N_7342);
and U9641 (N_9641,N_5641,N_6279);
or U9642 (N_9642,N_7129,N_5232);
or U9643 (N_9643,N_5228,N_5525);
and U9644 (N_9644,N_7135,N_6285);
or U9645 (N_9645,N_7387,N_5223);
nand U9646 (N_9646,N_6741,N_5748);
nor U9647 (N_9647,N_6610,N_5597);
nor U9648 (N_9648,N_7122,N_6435);
or U9649 (N_9649,N_6406,N_7147);
and U9650 (N_9650,N_5074,N_6239);
nor U9651 (N_9651,N_7059,N_6050);
nor U9652 (N_9652,N_5045,N_5136);
and U9653 (N_9653,N_7329,N_5152);
or U9654 (N_9654,N_7093,N_5967);
nand U9655 (N_9655,N_6965,N_6686);
and U9656 (N_9656,N_6925,N_6553);
and U9657 (N_9657,N_6650,N_5114);
or U9658 (N_9658,N_5747,N_5081);
nor U9659 (N_9659,N_6228,N_7223);
nand U9660 (N_9660,N_6559,N_7462);
and U9661 (N_9661,N_6358,N_5977);
and U9662 (N_9662,N_6160,N_7483);
nand U9663 (N_9663,N_6737,N_5629);
and U9664 (N_9664,N_5578,N_5661);
nand U9665 (N_9665,N_6481,N_5220);
nor U9666 (N_9666,N_5288,N_6471);
nor U9667 (N_9667,N_6996,N_5657);
nor U9668 (N_9668,N_5320,N_7020);
xnor U9669 (N_9669,N_7138,N_6513);
xor U9670 (N_9670,N_5342,N_5297);
xnor U9671 (N_9671,N_5687,N_5435);
or U9672 (N_9672,N_5027,N_5789);
or U9673 (N_9673,N_5694,N_5112);
or U9674 (N_9674,N_6544,N_5585);
nor U9675 (N_9675,N_7373,N_5125);
xnor U9676 (N_9676,N_5395,N_5937);
or U9677 (N_9677,N_5051,N_7237);
or U9678 (N_9678,N_5161,N_7117);
or U9679 (N_9679,N_6270,N_7321);
or U9680 (N_9680,N_5335,N_7161);
nor U9681 (N_9681,N_6511,N_5195);
or U9682 (N_9682,N_6206,N_5974);
or U9683 (N_9683,N_6875,N_6944);
xor U9684 (N_9684,N_5743,N_6176);
xor U9685 (N_9685,N_6219,N_6798);
nand U9686 (N_9686,N_5344,N_6959);
and U9687 (N_9687,N_7242,N_6335);
nor U9688 (N_9688,N_5178,N_6872);
or U9689 (N_9689,N_6754,N_7157);
nor U9690 (N_9690,N_6042,N_7436);
or U9691 (N_9691,N_6509,N_5777);
and U9692 (N_9692,N_5356,N_5186);
nand U9693 (N_9693,N_5715,N_5257);
xor U9694 (N_9694,N_6965,N_7289);
nand U9695 (N_9695,N_6540,N_6250);
and U9696 (N_9696,N_6930,N_6846);
and U9697 (N_9697,N_5469,N_5750);
and U9698 (N_9698,N_6037,N_6695);
or U9699 (N_9699,N_6354,N_5915);
nor U9700 (N_9700,N_6371,N_6901);
nand U9701 (N_9701,N_5863,N_6072);
xnor U9702 (N_9702,N_7302,N_6539);
nand U9703 (N_9703,N_6839,N_7396);
nor U9704 (N_9704,N_6437,N_7151);
and U9705 (N_9705,N_5466,N_5455);
xnor U9706 (N_9706,N_6173,N_5071);
nand U9707 (N_9707,N_6318,N_5453);
xnor U9708 (N_9708,N_5839,N_7035);
or U9709 (N_9709,N_6365,N_6180);
nor U9710 (N_9710,N_7069,N_6085);
nor U9711 (N_9711,N_5851,N_6192);
or U9712 (N_9712,N_5417,N_7068);
nand U9713 (N_9713,N_6356,N_5395);
and U9714 (N_9714,N_6291,N_5834);
or U9715 (N_9715,N_6100,N_5618);
nor U9716 (N_9716,N_6843,N_6279);
nor U9717 (N_9717,N_6525,N_7344);
or U9718 (N_9718,N_5679,N_7178);
and U9719 (N_9719,N_5415,N_6765);
nand U9720 (N_9720,N_7371,N_6607);
nand U9721 (N_9721,N_6500,N_6084);
nand U9722 (N_9722,N_5550,N_5664);
or U9723 (N_9723,N_5921,N_5979);
and U9724 (N_9724,N_7045,N_6136);
nor U9725 (N_9725,N_7448,N_5800);
nor U9726 (N_9726,N_7474,N_5085);
and U9727 (N_9727,N_7483,N_6253);
and U9728 (N_9728,N_6539,N_6807);
nor U9729 (N_9729,N_6489,N_5041);
or U9730 (N_9730,N_6340,N_5389);
or U9731 (N_9731,N_5173,N_7346);
nor U9732 (N_9732,N_6198,N_5254);
xnor U9733 (N_9733,N_6852,N_5813);
nor U9734 (N_9734,N_5414,N_5881);
nor U9735 (N_9735,N_7480,N_6335);
nor U9736 (N_9736,N_7033,N_6390);
xor U9737 (N_9737,N_5257,N_5205);
nand U9738 (N_9738,N_5207,N_6762);
nor U9739 (N_9739,N_7278,N_5445);
nand U9740 (N_9740,N_6844,N_6297);
nand U9741 (N_9741,N_7105,N_6310);
nand U9742 (N_9742,N_6930,N_6985);
and U9743 (N_9743,N_6315,N_6325);
nand U9744 (N_9744,N_5991,N_7303);
or U9745 (N_9745,N_6750,N_5311);
nor U9746 (N_9746,N_6136,N_6670);
nand U9747 (N_9747,N_7171,N_6209);
or U9748 (N_9748,N_5054,N_5705);
or U9749 (N_9749,N_6860,N_5900);
xor U9750 (N_9750,N_5566,N_5247);
nor U9751 (N_9751,N_5674,N_5388);
and U9752 (N_9752,N_5581,N_5574);
nor U9753 (N_9753,N_5751,N_6354);
nor U9754 (N_9754,N_5634,N_6412);
and U9755 (N_9755,N_5042,N_6433);
or U9756 (N_9756,N_5112,N_6852);
xnor U9757 (N_9757,N_6699,N_7203);
or U9758 (N_9758,N_7185,N_5670);
nor U9759 (N_9759,N_6401,N_7064);
nor U9760 (N_9760,N_7065,N_6267);
and U9761 (N_9761,N_5952,N_6309);
and U9762 (N_9762,N_5736,N_6731);
and U9763 (N_9763,N_6506,N_7082);
nand U9764 (N_9764,N_5914,N_5429);
or U9765 (N_9765,N_6196,N_6048);
and U9766 (N_9766,N_5371,N_5307);
xor U9767 (N_9767,N_5700,N_6697);
xnor U9768 (N_9768,N_6504,N_6110);
nor U9769 (N_9769,N_7302,N_5038);
and U9770 (N_9770,N_6200,N_7371);
or U9771 (N_9771,N_5095,N_6787);
nand U9772 (N_9772,N_7203,N_5075);
nand U9773 (N_9773,N_7259,N_6689);
or U9774 (N_9774,N_7426,N_5707);
nor U9775 (N_9775,N_5379,N_6024);
nor U9776 (N_9776,N_6989,N_6722);
or U9777 (N_9777,N_5609,N_5055);
nand U9778 (N_9778,N_6744,N_7069);
nand U9779 (N_9779,N_6602,N_7241);
and U9780 (N_9780,N_6815,N_5885);
and U9781 (N_9781,N_5377,N_6467);
or U9782 (N_9782,N_6541,N_5849);
and U9783 (N_9783,N_7193,N_5538);
nand U9784 (N_9784,N_7160,N_7162);
nor U9785 (N_9785,N_7184,N_5159);
xnor U9786 (N_9786,N_7367,N_5931);
xnor U9787 (N_9787,N_5626,N_5422);
or U9788 (N_9788,N_6207,N_6968);
and U9789 (N_9789,N_5161,N_5654);
nor U9790 (N_9790,N_5804,N_5592);
nor U9791 (N_9791,N_5899,N_6464);
or U9792 (N_9792,N_6243,N_5532);
or U9793 (N_9793,N_7031,N_7203);
nand U9794 (N_9794,N_5297,N_6174);
nor U9795 (N_9795,N_5558,N_5462);
nor U9796 (N_9796,N_6437,N_5092);
and U9797 (N_9797,N_6632,N_5667);
and U9798 (N_9798,N_7149,N_6850);
nand U9799 (N_9799,N_7039,N_7165);
nand U9800 (N_9800,N_6637,N_5155);
or U9801 (N_9801,N_5032,N_5915);
or U9802 (N_9802,N_7437,N_7479);
and U9803 (N_9803,N_5163,N_7395);
nor U9804 (N_9804,N_6677,N_5179);
nor U9805 (N_9805,N_6414,N_5729);
and U9806 (N_9806,N_7372,N_7346);
nand U9807 (N_9807,N_7033,N_5022);
nand U9808 (N_9808,N_7270,N_6230);
xnor U9809 (N_9809,N_5686,N_5684);
xnor U9810 (N_9810,N_7123,N_5233);
and U9811 (N_9811,N_5580,N_7373);
or U9812 (N_9812,N_5697,N_5366);
nor U9813 (N_9813,N_7082,N_6436);
nand U9814 (N_9814,N_5230,N_7268);
nor U9815 (N_9815,N_7419,N_6993);
or U9816 (N_9816,N_6846,N_7319);
nor U9817 (N_9817,N_6531,N_6878);
nor U9818 (N_9818,N_7152,N_6274);
nand U9819 (N_9819,N_6054,N_6098);
nor U9820 (N_9820,N_5559,N_5697);
or U9821 (N_9821,N_7399,N_6195);
nand U9822 (N_9822,N_6832,N_6863);
xnor U9823 (N_9823,N_6426,N_5780);
nor U9824 (N_9824,N_6918,N_5460);
or U9825 (N_9825,N_5892,N_5750);
nor U9826 (N_9826,N_5798,N_5129);
or U9827 (N_9827,N_7317,N_7073);
or U9828 (N_9828,N_7352,N_5912);
or U9829 (N_9829,N_6965,N_7397);
and U9830 (N_9830,N_6888,N_6283);
nor U9831 (N_9831,N_6709,N_5761);
nor U9832 (N_9832,N_5147,N_5802);
xor U9833 (N_9833,N_5307,N_5612);
xor U9834 (N_9834,N_5830,N_6551);
xnor U9835 (N_9835,N_6187,N_5359);
or U9836 (N_9836,N_5213,N_5453);
nor U9837 (N_9837,N_6033,N_6681);
and U9838 (N_9838,N_7005,N_5816);
and U9839 (N_9839,N_6287,N_5817);
nor U9840 (N_9840,N_5954,N_5097);
or U9841 (N_9841,N_5265,N_7367);
or U9842 (N_9842,N_5812,N_6154);
xor U9843 (N_9843,N_7058,N_6732);
nor U9844 (N_9844,N_6210,N_5947);
and U9845 (N_9845,N_5273,N_7396);
nor U9846 (N_9846,N_6092,N_6243);
and U9847 (N_9847,N_6060,N_5832);
nor U9848 (N_9848,N_5639,N_5886);
nor U9849 (N_9849,N_6334,N_6841);
or U9850 (N_9850,N_7117,N_5575);
or U9851 (N_9851,N_7082,N_5107);
nor U9852 (N_9852,N_7222,N_5715);
nor U9853 (N_9853,N_5291,N_5877);
and U9854 (N_9854,N_5258,N_5903);
or U9855 (N_9855,N_7189,N_5469);
nand U9856 (N_9856,N_5937,N_5831);
nor U9857 (N_9857,N_7179,N_6816);
nor U9858 (N_9858,N_6372,N_7110);
and U9859 (N_9859,N_7431,N_6324);
or U9860 (N_9860,N_6876,N_6165);
xnor U9861 (N_9861,N_6485,N_5723);
or U9862 (N_9862,N_5824,N_5938);
nor U9863 (N_9863,N_5866,N_5518);
nand U9864 (N_9864,N_5112,N_7357);
nor U9865 (N_9865,N_6608,N_7404);
nor U9866 (N_9866,N_6484,N_5799);
nand U9867 (N_9867,N_7025,N_6531);
nor U9868 (N_9868,N_7001,N_5184);
nor U9869 (N_9869,N_5217,N_6922);
and U9870 (N_9870,N_5281,N_6814);
or U9871 (N_9871,N_6280,N_6613);
or U9872 (N_9872,N_5352,N_5110);
nor U9873 (N_9873,N_7418,N_7021);
or U9874 (N_9874,N_5009,N_5718);
nand U9875 (N_9875,N_7062,N_6331);
nor U9876 (N_9876,N_5645,N_6301);
nor U9877 (N_9877,N_7329,N_5933);
nor U9878 (N_9878,N_6916,N_7124);
nor U9879 (N_9879,N_5343,N_7336);
nor U9880 (N_9880,N_6749,N_6586);
xor U9881 (N_9881,N_5849,N_7069);
and U9882 (N_9882,N_5001,N_5728);
or U9883 (N_9883,N_5552,N_6425);
nor U9884 (N_9884,N_5680,N_5479);
nor U9885 (N_9885,N_6557,N_5487);
and U9886 (N_9886,N_5584,N_7033);
xnor U9887 (N_9887,N_5242,N_6538);
xnor U9888 (N_9888,N_6672,N_7396);
nor U9889 (N_9889,N_7047,N_6599);
and U9890 (N_9890,N_7444,N_6793);
and U9891 (N_9891,N_6894,N_6617);
nor U9892 (N_9892,N_6105,N_6795);
nand U9893 (N_9893,N_7203,N_5803);
or U9894 (N_9894,N_6286,N_6978);
or U9895 (N_9895,N_6200,N_5699);
nand U9896 (N_9896,N_5630,N_5350);
or U9897 (N_9897,N_6458,N_6683);
or U9898 (N_9898,N_5489,N_7355);
or U9899 (N_9899,N_6374,N_5657);
and U9900 (N_9900,N_7423,N_7268);
xnor U9901 (N_9901,N_5626,N_5909);
nand U9902 (N_9902,N_5130,N_6181);
and U9903 (N_9903,N_5260,N_7084);
and U9904 (N_9904,N_5373,N_6692);
nand U9905 (N_9905,N_5952,N_5138);
or U9906 (N_9906,N_5478,N_5695);
nor U9907 (N_9907,N_6017,N_5356);
nor U9908 (N_9908,N_5556,N_5180);
xnor U9909 (N_9909,N_5400,N_5443);
or U9910 (N_9910,N_5321,N_5244);
nor U9911 (N_9911,N_6044,N_7110);
xnor U9912 (N_9912,N_6838,N_6061);
or U9913 (N_9913,N_6498,N_6398);
nand U9914 (N_9914,N_5622,N_6144);
and U9915 (N_9915,N_5782,N_5037);
nand U9916 (N_9916,N_6021,N_6531);
and U9917 (N_9917,N_6988,N_6931);
and U9918 (N_9918,N_5125,N_6681);
xor U9919 (N_9919,N_5222,N_7114);
nor U9920 (N_9920,N_7313,N_7273);
and U9921 (N_9921,N_5831,N_5255);
and U9922 (N_9922,N_6477,N_6257);
nor U9923 (N_9923,N_6685,N_5113);
and U9924 (N_9924,N_7189,N_6786);
nor U9925 (N_9925,N_6258,N_6526);
nand U9926 (N_9926,N_5325,N_5115);
and U9927 (N_9927,N_5074,N_5442);
nor U9928 (N_9928,N_5949,N_6370);
nand U9929 (N_9929,N_7215,N_5987);
nand U9930 (N_9930,N_7053,N_5621);
or U9931 (N_9931,N_6618,N_5884);
nor U9932 (N_9932,N_5139,N_6506);
and U9933 (N_9933,N_5268,N_7126);
or U9934 (N_9934,N_6589,N_5377);
and U9935 (N_9935,N_6153,N_6293);
and U9936 (N_9936,N_6684,N_7092);
nor U9937 (N_9937,N_5829,N_7062);
nor U9938 (N_9938,N_5493,N_6095);
or U9939 (N_9939,N_6706,N_5787);
xor U9940 (N_9940,N_5947,N_6656);
nor U9941 (N_9941,N_5475,N_6281);
and U9942 (N_9942,N_5571,N_7028);
or U9943 (N_9943,N_6861,N_6456);
or U9944 (N_9944,N_7438,N_6458);
nor U9945 (N_9945,N_5032,N_6655);
nor U9946 (N_9946,N_5236,N_5501);
nand U9947 (N_9947,N_6861,N_5531);
nor U9948 (N_9948,N_5988,N_5193);
or U9949 (N_9949,N_6180,N_5364);
or U9950 (N_9950,N_7404,N_6538);
or U9951 (N_9951,N_6201,N_6542);
nor U9952 (N_9952,N_7168,N_7284);
nand U9953 (N_9953,N_5819,N_5166);
or U9954 (N_9954,N_5969,N_7193);
nor U9955 (N_9955,N_6582,N_6474);
nand U9956 (N_9956,N_5092,N_6605);
nor U9957 (N_9957,N_5071,N_7290);
nor U9958 (N_9958,N_5879,N_5995);
or U9959 (N_9959,N_5361,N_6567);
nand U9960 (N_9960,N_5076,N_6595);
or U9961 (N_9961,N_7407,N_6870);
and U9962 (N_9962,N_6173,N_6004);
and U9963 (N_9963,N_6255,N_7322);
and U9964 (N_9964,N_7362,N_6830);
or U9965 (N_9965,N_5545,N_6364);
and U9966 (N_9966,N_6703,N_5968);
nor U9967 (N_9967,N_5528,N_6247);
or U9968 (N_9968,N_6540,N_6677);
nand U9969 (N_9969,N_6975,N_5764);
nand U9970 (N_9970,N_5392,N_6453);
or U9971 (N_9971,N_6026,N_5221);
xnor U9972 (N_9972,N_5748,N_6895);
nand U9973 (N_9973,N_6223,N_6290);
or U9974 (N_9974,N_7345,N_5224);
or U9975 (N_9975,N_7494,N_6193);
or U9976 (N_9976,N_5406,N_6053);
nand U9977 (N_9977,N_6796,N_5819);
xnor U9978 (N_9978,N_5200,N_6350);
nor U9979 (N_9979,N_6043,N_6834);
nand U9980 (N_9980,N_6022,N_6790);
nor U9981 (N_9981,N_6073,N_5981);
xor U9982 (N_9982,N_5408,N_5755);
nor U9983 (N_9983,N_5234,N_6459);
or U9984 (N_9984,N_7018,N_6580);
nor U9985 (N_9985,N_6471,N_6449);
nand U9986 (N_9986,N_5445,N_5331);
xnor U9987 (N_9987,N_6311,N_6226);
xnor U9988 (N_9988,N_5389,N_6631);
and U9989 (N_9989,N_6655,N_5314);
nor U9990 (N_9990,N_5137,N_6562);
or U9991 (N_9991,N_6488,N_5987);
and U9992 (N_9992,N_7046,N_6479);
nand U9993 (N_9993,N_6168,N_6065);
nand U9994 (N_9994,N_5371,N_6835);
xnor U9995 (N_9995,N_6522,N_5758);
and U9996 (N_9996,N_6003,N_5097);
nand U9997 (N_9997,N_6456,N_6158);
nand U9998 (N_9998,N_6046,N_7211);
xnor U9999 (N_9999,N_5705,N_6492);
or U10000 (N_10000,N_7946,N_9438);
or U10001 (N_10001,N_9108,N_9532);
nand U10002 (N_10002,N_9258,N_8373);
and U10003 (N_10003,N_9703,N_9304);
nor U10004 (N_10004,N_8986,N_7882);
and U10005 (N_10005,N_7582,N_9422);
or U10006 (N_10006,N_8261,N_9209);
nand U10007 (N_10007,N_8442,N_9733);
or U10008 (N_10008,N_9364,N_7999);
and U10009 (N_10009,N_9833,N_9693);
nor U10010 (N_10010,N_7903,N_7804);
nor U10011 (N_10011,N_8733,N_9016);
and U10012 (N_10012,N_9037,N_9701);
xor U10013 (N_10013,N_8761,N_8651);
or U10014 (N_10014,N_8289,N_9850);
or U10015 (N_10015,N_8087,N_7566);
nand U10016 (N_10016,N_7696,N_8911);
nor U10017 (N_10017,N_9759,N_8328);
or U10018 (N_10018,N_9130,N_8740);
xnor U10019 (N_10019,N_8735,N_7931);
nand U10020 (N_10020,N_9869,N_9349);
or U10021 (N_10021,N_8010,N_8209);
xnor U10022 (N_10022,N_8746,N_7857);
and U10023 (N_10023,N_9932,N_8538);
or U10024 (N_10024,N_7586,N_9107);
or U10025 (N_10025,N_8562,N_9671);
or U10026 (N_10026,N_9250,N_7686);
and U10027 (N_10027,N_7834,N_8815);
and U10028 (N_10028,N_7912,N_8426);
or U10029 (N_10029,N_9231,N_9921);
or U10030 (N_10030,N_9604,N_9573);
or U10031 (N_10031,N_8549,N_7744);
nand U10032 (N_10032,N_7928,N_8490);
nor U10033 (N_10033,N_9112,N_9399);
nor U10034 (N_10034,N_9688,N_8688);
and U10035 (N_10035,N_7802,N_9819);
nor U10036 (N_10036,N_8276,N_8903);
xor U10037 (N_10037,N_9172,N_9760);
xor U10038 (N_10038,N_8309,N_8904);
xor U10039 (N_10039,N_7665,N_9907);
nor U10040 (N_10040,N_9502,N_7898);
nor U10041 (N_10041,N_9060,N_7574);
and U10042 (N_10042,N_9911,N_8559);
nand U10043 (N_10043,N_8491,N_9451);
xnor U10044 (N_10044,N_8874,N_9981);
or U10045 (N_10045,N_9647,N_9941);
or U10046 (N_10046,N_9135,N_8131);
nand U10047 (N_10047,N_8629,N_8274);
and U10048 (N_10048,N_7752,N_9221);
or U10049 (N_10049,N_7572,N_9335);
nand U10050 (N_10050,N_7821,N_7695);
and U10051 (N_10051,N_9627,N_8308);
nor U10052 (N_10052,N_9073,N_7532);
or U10053 (N_10053,N_9961,N_7934);
xnor U10054 (N_10054,N_9249,N_7758);
nand U10055 (N_10055,N_8482,N_7925);
nand U10056 (N_10056,N_9722,N_7693);
and U10057 (N_10057,N_7539,N_8083);
and U10058 (N_10058,N_8163,N_8546);
nand U10059 (N_10059,N_7808,N_9238);
or U10060 (N_10060,N_9425,N_8727);
nor U10061 (N_10061,N_9928,N_9577);
or U10062 (N_10062,N_9998,N_8254);
or U10063 (N_10063,N_8719,N_9867);
nand U10064 (N_10064,N_7593,N_8056);
and U10065 (N_10065,N_7690,N_9835);
or U10066 (N_10066,N_8435,N_8027);
and U10067 (N_10067,N_9610,N_9939);
nand U10068 (N_10068,N_8392,N_8013);
and U10069 (N_10069,N_8714,N_9456);
xor U10070 (N_10070,N_8601,N_9235);
and U10071 (N_10071,N_7987,N_8658);
and U10072 (N_10072,N_9333,N_7552);
and U10073 (N_10073,N_9536,N_8967);
or U10074 (N_10074,N_9718,N_9484);
xnor U10075 (N_10075,N_8657,N_8793);
xnor U10076 (N_10076,N_8600,N_9372);
xor U10077 (N_10077,N_8989,N_9297);
nand U10078 (N_10078,N_8397,N_8560);
nand U10079 (N_10079,N_9291,N_8246);
and U10080 (N_10080,N_9470,N_8036);
and U10081 (N_10081,N_8631,N_8234);
and U10082 (N_10082,N_8304,N_8186);
and U10083 (N_10083,N_7543,N_7516);
nor U10084 (N_10084,N_9368,N_9567);
and U10085 (N_10085,N_9500,N_7520);
nand U10086 (N_10086,N_8220,N_8148);
and U10087 (N_10087,N_8350,N_9924);
nor U10088 (N_10088,N_9408,N_8647);
and U10089 (N_10089,N_9972,N_7775);
or U10090 (N_10090,N_9487,N_8138);
nor U10091 (N_10091,N_8336,N_8934);
or U10092 (N_10092,N_8583,N_9239);
nand U10093 (N_10093,N_9452,N_9247);
xor U10094 (N_10094,N_8883,N_9793);
nand U10095 (N_10095,N_8360,N_9667);
and U10096 (N_10096,N_9363,N_9350);
nand U10097 (N_10097,N_8505,N_8499);
nor U10098 (N_10098,N_9863,N_8528);
nand U10099 (N_10099,N_7880,N_8994);
and U10100 (N_10100,N_7745,N_7932);
nor U10101 (N_10101,N_8949,N_7832);
and U10102 (N_10102,N_7678,N_8099);
nand U10103 (N_10103,N_8877,N_8170);
or U10104 (N_10104,N_7778,N_9906);
and U10105 (N_10105,N_8586,N_9785);
and U10106 (N_10106,N_9728,N_7637);
or U10107 (N_10107,N_8094,N_8756);
nand U10108 (N_10108,N_8625,N_9462);
or U10109 (N_10109,N_9008,N_8645);
and U10110 (N_10110,N_8782,N_7746);
or U10111 (N_10111,N_8997,N_9529);
xor U10112 (N_10112,N_9582,N_9136);
and U10113 (N_10113,N_8451,N_8481);
xor U10114 (N_10114,N_8928,N_9988);
nand U10115 (N_10115,N_7776,N_7883);
nor U10116 (N_10116,N_9881,N_9549);
nand U10117 (N_10117,N_8324,N_7813);
nand U10118 (N_10118,N_7535,N_7551);
or U10119 (N_10119,N_9358,N_9384);
and U10120 (N_10120,N_9809,N_8823);
or U10121 (N_10121,N_8085,N_8759);
xor U10122 (N_10122,N_9465,N_8183);
nor U10123 (N_10123,N_8074,N_9200);
and U10124 (N_10124,N_8193,N_8568);
nand U10125 (N_10125,N_9361,N_7651);
nor U10126 (N_10126,N_7647,N_8409);
nand U10127 (N_10127,N_9413,N_8743);
nand U10128 (N_10128,N_9146,N_8580);
and U10129 (N_10129,N_9613,N_8582);
nor U10130 (N_10130,N_7526,N_9575);
and U10131 (N_10131,N_8101,N_7640);
or U10132 (N_10132,N_9806,N_8908);
nor U10133 (N_10133,N_9829,N_8256);
nand U10134 (N_10134,N_7954,N_8547);
nand U10135 (N_10135,N_9755,N_8766);
and U10136 (N_10136,N_8984,N_9486);
nand U10137 (N_10137,N_7591,N_7700);
or U10138 (N_10138,N_8914,N_8872);
xnor U10139 (N_10139,N_9475,N_9959);
or U10140 (N_10140,N_7867,N_9746);
xor U10141 (N_10141,N_9898,N_9531);
nand U10142 (N_10142,N_9587,N_7772);
and U10143 (N_10143,N_8891,N_7740);
and U10144 (N_10144,N_7994,N_7565);
nor U10145 (N_10145,N_8362,N_7998);
or U10146 (N_10146,N_8369,N_7580);
or U10147 (N_10147,N_9915,N_8152);
or U10148 (N_10148,N_9689,N_8952);
and U10149 (N_10149,N_9257,N_7988);
nand U10150 (N_10150,N_7975,N_9884);
and U10151 (N_10151,N_9786,N_8382);
and U10152 (N_10152,N_8253,N_8439);
xor U10153 (N_10153,N_8455,N_9749);
and U10154 (N_10154,N_7504,N_9449);
nor U10155 (N_10155,N_8709,N_8410);
or U10156 (N_10156,N_7915,N_8454);
nand U10157 (N_10157,N_7781,N_9878);
and U10158 (N_10158,N_9712,N_8948);
xor U10159 (N_10159,N_9679,N_8805);
nand U10160 (N_10160,N_7791,N_9044);
nor U10161 (N_10161,N_9735,N_9986);
or U10162 (N_10162,N_8749,N_7818);
or U10163 (N_10163,N_8955,N_9454);
xnor U10164 (N_10164,N_7762,N_9427);
or U10165 (N_10165,N_9153,N_8178);
nor U10166 (N_10166,N_7542,N_7664);
nand U10167 (N_10167,N_9930,N_9094);
nor U10168 (N_10168,N_9894,N_7659);
or U10169 (N_10169,N_7506,N_8998);
xnor U10170 (N_10170,N_8831,N_8752);
nor U10171 (N_10171,N_8205,N_7942);
nand U10172 (N_10172,N_9958,N_9453);
or U10173 (N_10173,N_9841,N_9284);
nor U10174 (N_10174,N_9710,N_9559);
nor U10175 (N_10175,N_8999,N_9338);
nor U10176 (N_10176,N_8970,N_7757);
and U10177 (N_10177,N_9705,N_9217);
and U10178 (N_10178,N_8540,N_8912);
nand U10179 (N_10179,N_9858,N_7841);
nor U10180 (N_10180,N_7798,N_8195);
nor U10181 (N_10181,N_8694,N_8469);
nand U10182 (N_10182,N_8222,N_8809);
or U10183 (N_10183,N_8945,N_8450);
or U10184 (N_10184,N_8850,N_7560);
or U10185 (N_10185,N_9123,N_8281);
and U10186 (N_10186,N_7793,N_8407);
xnor U10187 (N_10187,N_8069,N_8251);
nor U10188 (N_10188,N_7812,N_8058);
nand U10189 (N_10189,N_9652,N_7519);
nor U10190 (N_10190,N_8247,N_9090);
nor U10191 (N_10191,N_7581,N_8555);
nor U10192 (N_10192,N_7761,N_7767);
or U10193 (N_10193,N_9659,N_8242);
nand U10194 (N_10194,N_8834,N_9052);
or U10195 (N_10195,N_9187,N_8897);
and U10196 (N_10196,N_8574,N_9723);
xor U10197 (N_10197,N_7536,N_9158);
nor U10198 (N_10198,N_7939,N_8239);
and U10199 (N_10199,N_9311,N_9109);
nor U10200 (N_10200,N_7789,N_7773);
and U10201 (N_10201,N_9691,N_9264);
nand U10202 (N_10202,N_8849,N_9043);
nand U10203 (N_10203,N_9820,N_7685);
nand U10204 (N_10204,N_9715,N_8497);
or U10205 (N_10205,N_7610,N_7531);
nor U10206 (N_10206,N_7787,N_8682);
nand U10207 (N_10207,N_9070,N_7937);
xnor U10208 (N_10208,N_8621,N_8861);
nor U10209 (N_10209,N_8594,N_9560);
and U10210 (N_10210,N_8475,N_9104);
nand U10211 (N_10211,N_9514,N_7839);
xor U10212 (N_10212,N_9828,N_9357);
or U10213 (N_10213,N_8366,N_7684);
nand U10214 (N_10214,N_9325,N_8436);
and U10215 (N_10215,N_9448,N_9195);
nor U10216 (N_10216,N_9547,N_8327);
nand U10217 (N_10217,N_8526,N_8859);
nor U10218 (N_10218,N_8930,N_8660);
or U10219 (N_10219,N_8656,N_9240);
nand U10220 (N_10220,N_9161,N_8768);
or U10221 (N_10221,N_9039,N_8609);
or U10222 (N_10222,N_9354,N_9155);
nor U10223 (N_10223,N_8020,N_9134);
or U10224 (N_10224,N_9129,N_8618);
nor U10225 (N_10225,N_7710,N_7889);
nor U10226 (N_10226,N_9446,N_7753);
nand U10227 (N_10227,N_8964,N_9836);
nand U10228 (N_10228,N_8187,N_8889);
nor U10229 (N_10229,N_7972,N_8430);
nor U10230 (N_10230,N_7719,N_9504);
and U10231 (N_10231,N_7800,N_7615);
or U10232 (N_10232,N_7731,N_9555);
or U10233 (N_10233,N_7784,N_7725);
nor U10234 (N_10234,N_7720,N_7661);
or U10235 (N_10235,N_9694,N_8567);
nand U10236 (N_10236,N_7973,N_9381);
or U10237 (N_10237,N_9685,N_9199);
xnor U10238 (N_10238,N_8884,N_7632);
nor U10239 (N_10239,N_8675,N_9101);
or U10240 (N_10240,N_9375,N_8478);
nand U10241 (N_10241,N_7514,N_9886);
nand U10242 (N_10242,N_8194,N_9089);
or U10243 (N_10243,N_9795,N_7783);
and U10244 (N_10244,N_7518,N_8344);
nor U10245 (N_10245,N_7865,N_8981);
nand U10246 (N_10246,N_8700,N_9498);
and U10247 (N_10247,N_9117,N_9439);
nor U10248 (N_10248,N_8520,N_7698);
nand U10249 (N_10249,N_8100,N_7616);
or U10250 (N_10250,N_8090,N_8638);
and U10251 (N_10251,N_7517,N_8312);
and U10252 (N_10252,N_8725,N_9927);
nand U10253 (N_10253,N_9063,N_8875);
or U10254 (N_10254,N_8093,N_8046);
nor U10255 (N_10255,N_8742,N_7823);
nor U10256 (N_10256,N_7782,N_8781);
and U10257 (N_10257,N_7962,N_8622);
and U10258 (N_10258,N_9663,N_9233);
or U10259 (N_10259,N_8288,N_9579);
and U10260 (N_10260,N_8716,N_9434);
and U10261 (N_10261,N_9821,N_8798);
nand U10262 (N_10262,N_8221,N_9692);
and U10263 (N_10263,N_9492,N_8367);
nand U10264 (N_10264,N_7851,N_8991);
nor U10265 (N_10265,N_8257,N_9113);
or U10266 (N_10266,N_7741,N_9651);
and U10267 (N_10267,N_9519,N_8443);
nand U10268 (N_10268,N_8018,N_8134);
or U10269 (N_10269,N_9208,N_8424);
and U10270 (N_10270,N_9513,N_8208);
nor U10271 (N_10271,N_8236,N_9708);
or U10272 (N_10272,N_9156,N_8917);
nand U10273 (N_10273,N_8990,N_8077);
nand U10274 (N_10274,N_7828,N_9218);
xor U10275 (N_10275,N_7952,N_9159);
nand U10276 (N_10276,N_9441,N_7612);
and U10277 (N_10277,N_9846,N_8370);
and U10278 (N_10278,N_7985,N_8286);
or U10279 (N_10279,N_7525,N_9175);
and U10280 (N_10280,N_9936,N_9406);
or U10281 (N_10281,N_7922,N_9457);
nand U10282 (N_10282,N_9526,N_8411);
or U10283 (N_10283,N_9080,N_7672);
nand U10284 (N_10284,N_8472,N_9933);
and U10285 (N_10285,N_8920,N_9724);
and U10286 (N_10286,N_7623,N_7620);
nor U10287 (N_10287,N_8376,N_8206);
or U10288 (N_10288,N_7614,N_8347);
and U10289 (N_10289,N_8713,N_9009);
nor U10290 (N_10290,N_9267,N_9962);
or U10291 (N_10291,N_7528,N_9459);
or U10292 (N_10292,N_9750,N_8154);
or U10293 (N_10293,N_7707,N_8707);
and U10294 (N_10294,N_7763,N_8937);
nor U10295 (N_10295,N_7881,N_8202);
nor U10296 (N_10296,N_9277,N_8953);
nand U10297 (N_10297,N_9509,N_9100);
nor U10298 (N_10298,N_7562,N_9802);
nor U10299 (N_10299,N_8364,N_8825);
or U10300 (N_10300,N_8591,N_8237);
nand U10301 (N_10301,N_7971,N_8294);
xnor U10302 (N_10302,N_8425,N_8837);
nand U10303 (N_10303,N_8541,N_9160);
and U10304 (N_10304,N_9864,N_7554);
nand U10305 (N_10305,N_9803,N_7508);
nor U10306 (N_10306,N_8975,N_9322);
nor U10307 (N_10307,N_9995,N_8285);
nor U10308 (N_10308,N_8806,N_8144);
or U10309 (N_10309,N_7642,N_7897);
and U10310 (N_10310,N_7792,N_7852);
nand U10311 (N_10311,N_7564,N_9516);
xnor U10312 (N_10312,N_9030,N_9676);
and U10313 (N_10313,N_9312,N_8507);
nand U10314 (N_10314,N_9120,N_9271);
nor U10315 (N_10315,N_9093,N_8462);
nand U10316 (N_10316,N_9203,N_8744);
xnor U10317 (N_10317,N_8189,N_8685);
or U10318 (N_10318,N_8810,N_8676);
nand U10319 (N_10319,N_9789,N_8244);
and U10320 (N_10320,N_9507,N_8264);
or U10321 (N_10321,N_9654,N_8649);
or U10322 (N_10322,N_8722,N_8856);
and U10323 (N_10323,N_9642,N_9868);
and U10324 (N_10324,N_8732,N_8597);
xnor U10325 (N_10325,N_9949,N_9814);
nand U10326 (N_10326,N_9404,N_9281);
or U10327 (N_10327,N_8946,N_8433);
nand U10328 (N_10328,N_8203,N_8042);
nand U10329 (N_10329,N_9403,N_8331);
xor U10330 (N_10330,N_8755,N_8581);
nand U10331 (N_10331,N_7904,N_8282);
and U10332 (N_10332,N_9031,N_8318);
nor U10333 (N_10333,N_9272,N_8476);
or U10334 (N_10334,N_8092,N_9489);
or U10335 (N_10335,N_7935,N_8035);
nand U10336 (N_10336,N_8182,N_9818);
or U10337 (N_10337,N_8137,N_7955);
xnor U10338 (N_10338,N_8471,N_9853);
nor U10339 (N_10339,N_7588,N_7618);
and U10340 (N_10340,N_8391,N_9817);
nand U10341 (N_10341,N_9079,N_7630);
or U10342 (N_10342,N_9309,N_9002);
nor U10343 (N_10343,N_9816,N_9234);
or U10344 (N_10344,N_8672,N_8215);
or U10345 (N_10345,N_8412,N_8474);
xnor U10346 (N_10346,N_8200,N_9256);
or U10347 (N_10347,N_8233,N_9882);
and U10348 (N_10348,N_9164,N_9618);
and U10349 (N_10349,N_8386,N_9762);
or U10350 (N_10350,N_7596,N_7980);
or U10351 (N_10351,N_9274,N_9334);
nand U10352 (N_10352,N_8579,N_9677);
nor U10353 (N_10353,N_9469,N_8315);
nand U10354 (N_10354,N_9352,N_9464);
or U10355 (N_10355,N_7811,N_9860);
and U10356 (N_10356,N_9143,N_9213);
nor U10357 (N_10357,N_8057,N_7894);
nand U10358 (N_10358,N_7599,N_9024);
xor U10359 (N_10359,N_9388,N_9788);
xnor U10360 (N_10360,N_8537,N_9808);
and U10361 (N_10361,N_9308,N_7703);
nand U10362 (N_10362,N_9974,N_8155);
or U10363 (N_10363,N_9952,N_8860);
xor U10364 (N_10364,N_8635,N_8669);
or U10365 (N_10365,N_9483,N_8053);
nand U10366 (N_10366,N_8852,N_9241);
or U10367 (N_10367,N_9386,N_8223);
nor U10368 (N_10368,N_7578,N_8295);
xnor U10369 (N_10369,N_9222,N_9026);
or U10370 (N_10370,N_8045,N_9268);
and U10371 (N_10371,N_9313,N_9518);
nand U10372 (N_10372,N_9626,N_8403);
nand U10373 (N_10373,N_8695,N_8033);
or U10374 (N_10374,N_9077,N_7673);
or U10375 (N_10375,N_9300,N_7675);
or U10376 (N_10376,N_8941,N_8062);
and U10377 (N_10377,N_7859,N_7683);
nand U10378 (N_10378,N_8011,N_9690);
nor U10379 (N_10379,N_8570,N_9811);
nand U10380 (N_10380,N_9551,N_7501);
nor U10381 (N_10381,N_8627,N_9251);
and U10382 (N_10382,N_9299,N_9485);
nor U10383 (N_10383,N_9632,N_8771);
nor U10384 (N_10384,N_8265,N_7826);
and U10385 (N_10385,N_7936,N_8380);
or U10386 (N_10386,N_7995,N_8484);
and U10387 (N_10387,N_9049,N_8530);
and U10388 (N_10388,N_8477,N_9302);
and U10389 (N_10389,N_9584,N_9510);
and U10390 (N_10390,N_8630,N_8835);
nand U10391 (N_10391,N_8923,N_9893);
nor U10392 (N_10392,N_9048,N_8379);
and U10393 (N_10393,N_8689,N_8381);
and U10394 (N_10394,N_8136,N_7723);
or U10395 (N_10395,N_9503,N_7510);
nand U10396 (N_10396,N_7633,N_9373);
nor U10397 (N_10397,N_8351,N_8836);
nand U10398 (N_10398,N_7991,N_9657);
or U10399 (N_10399,N_8414,N_9145);
nand U10400 (N_10400,N_9463,N_9356);
or U10401 (N_10401,N_9047,N_8792);
xnor U10402 (N_10402,N_8738,N_7641);
or U10403 (N_10403,N_7885,N_8841);
nand U10404 (N_10404,N_7626,N_8263);
nand U10405 (N_10405,N_8071,N_8204);
nand U10406 (N_10406,N_8933,N_8047);
or U10407 (N_10407,N_9607,N_9188);
nand U10408 (N_10408,N_8429,N_8159);
and U10409 (N_10409,N_9612,N_9431);
nand U10410 (N_10410,N_8905,N_9353);
or U10411 (N_10411,N_9371,N_8198);
nor U10412 (N_10412,N_8993,N_8824);
nor U10413 (N_10413,N_7921,N_8420);
and U10414 (N_10414,N_8015,N_9597);
or U10415 (N_10415,N_9849,N_8663);
nand U10416 (N_10416,N_8019,N_9367);
nand U10417 (N_10417,N_9336,N_8321);
xor U10418 (N_10418,N_9269,N_8977);
and U10419 (N_10419,N_7639,N_8338);
nand U10420 (N_10420,N_7919,N_8465);
xnor U10421 (N_10421,N_8863,N_8219);
nand U10422 (N_10422,N_9768,N_7544);
nand U10423 (N_10423,N_8985,N_8697);
or U10424 (N_10424,N_9989,N_9606);
nor U10425 (N_10425,N_9056,N_8396);
or U10426 (N_10426,N_8365,N_8633);
and U10427 (N_10427,N_7644,N_7742);
nor U10428 (N_10428,N_9067,N_9407);
and U10429 (N_10429,N_8646,N_7905);
and U10430 (N_10430,N_8565,N_8156);
and U10431 (N_10431,N_8119,N_9620);
xor U10432 (N_10432,N_8736,N_9339);
or U10433 (N_10433,N_7704,N_7896);
or U10434 (N_10434,N_8624,N_8238);
nand U10435 (N_10435,N_8421,N_8241);
xor U10436 (N_10436,N_7602,N_8302);
and U10437 (N_10437,N_9540,N_9224);
or U10438 (N_10438,N_8003,N_9097);
xnor U10439 (N_10439,N_8385,N_8662);
nor U10440 (N_10440,N_9292,N_7901);
and U10441 (N_10441,N_7691,N_8395);
nor U10442 (N_10442,N_9205,N_7879);
and U10443 (N_10443,N_8717,N_8516);
or U10444 (N_10444,N_9912,N_8383);
or U10445 (N_10445,N_8607,N_8388);
nand U10446 (N_10446,N_9098,N_8778);
and U10447 (N_10447,N_7561,N_9976);
nor U10448 (N_10448,N_8361,N_8073);
nor U10449 (N_10449,N_9609,N_8199);
xnor U10450 (N_10450,N_8728,N_7825);
nor U10451 (N_10451,N_8269,N_9660);
xnor U10452 (N_10452,N_8005,N_8864);
nor U10453 (N_10453,N_7847,N_9523);
nand U10454 (N_10454,N_9698,N_9596);
nand U10455 (N_10455,N_8402,N_8561);
xor U10456 (N_10456,N_7521,N_8001);
nor U10457 (N_10457,N_9730,N_9535);
nor U10458 (N_10458,N_9937,N_9103);
and U10459 (N_10459,N_9824,N_9005);
nor U10460 (N_10460,N_7829,N_8218);
or U10461 (N_10461,N_8514,N_7712);
xor U10462 (N_10462,N_8374,N_8287);
nor U10463 (N_10463,N_9279,N_9887);
or U10464 (N_10464,N_9641,N_9925);
nand U10465 (N_10465,N_8457,N_8612);
nor U10466 (N_10466,N_7820,N_8616);
xnor U10467 (N_10467,N_9854,N_8483);
nand U10468 (N_10468,N_7957,N_8593);
and U10469 (N_10469,N_8311,N_8319);
or U10470 (N_10470,N_9740,N_9889);
or U10471 (N_10471,N_8335,N_9374);
nand U10472 (N_10472,N_9359,N_8317);
or U10473 (N_10473,N_8487,N_9592);
nand U10474 (N_10474,N_8250,N_9702);
or U10475 (N_10475,N_9148,N_7785);
and U10476 (N_10476,N_9650,N_8988);
nand U10477 (N_10477,N_9711,N_9955);
or U10478 (N_10478,N_9751,N_8963);
nand U10479 (N_10479,N_8940,N_9400);
and U10480 (N_10480,N_7981,N_7537);
nand U10481 (N_10481,N_9013,N_9466);
xor U10482 (N_10482,N_9416,N_8765);
nor U10483 (N_10483,N_7965,N_9001);
nand U10484 (N_10484,N_7576,N_8384);
nand U10485 (N_10485,N_7682,N_9387);
nand U10486 (N_10486,N_9266,N_9042);
nor U10487 (N_10487,N_8339,N_9402);
nor U10488 (N_10488,N_8117,N_8006);
or U10489 (N_10489,N_8811,N_8639);
and U10490 (N_10490,N_7730,N_9140);
nand U10491 (N_10491,N_9614,N_8827);
nand U10492 (N_10492,N_8348,N_8297);
and U10493 (N_10493,N_7674,N_9035);
nand U10494 (N_10494,N_8213,N_9390);
or U10495 (N_10495,N_9902,N_7702);
nor U10496 (N_10496,N_9774,N_8853);
nor U10497 (N_10497,N_7838,N_8915);
or U10498 (N_10498,N_8983,N_9993);
nor U10499 (N_10499,N_8463,N_7966);
nor U10500 (N_10500,N_9658,N_8800);
nand U10501 (N_10501,N_8158,N_8779);
or U10502 (N_10502,N_9246,N_8479);
xor U10503 (N_10503,N_8394,N_8126);
xnor U10504 (N_10504,N_7734,N_8783);
or U10505 (N_10505,N_7967,N_9377);
or U10506 (N_10506,N_8773,N_9591);
nand U10507 (N_10507,N_8648,N_9191);
nor U10508 (N_10508,N_9877,N_8508);
nor U10509 (N_10509,N_9283,N_9355);
or U10510 (N_10510,N_8552,N_9787);
nor U10511 (N_10511,N_8762,N_8803);
nand U10512 (N_10512,N_8091,N_8924);
xnor U10513 (N_10513,N_9538,N_8842);
and U10514 (N_10514,N_8532,N_8626);
nor U10515 (N_10515,N_9741,N_7628);
nand U10516 (N_10516,N_9649,N_8828);
nor U10517 (N_10517,N_8720,N_7527);
nor U10518 (N_10518,N_8865,N_7646);
or U10519 (N_10519,N_9069,N_9149);
or U10520 (N_10520,N_7856,N_7715);
nor U10521 (N_10521,N_7729,N_7652);
or U10522 (N_10522,N_9275,N_8775);
nor U10523 (N_10523,N_9180,N_8017);
nand U10524 (N_10524,N_8192,N_8323);
nor U10525 (N_10525,N_9141,N_8470);
nand U10526 (N_10526,N_8217,N_9997);
and U10527 (N_10527,N_8343,N_9920);
or U10528 (N_10528,N_7587,N_9985);
nand U10529 (N_10529,N_8228,N_9611);
and U10530 (N_10530,N_7713,N_7884);
or U10531 (N_10531,N_9978,N_7502);
nor U10532 (N_10532,N_8518,N_9916);
and U10533 (N_10533,N_8168,N_9321);
xnor U10534 (N_10534,N_9289,N_9904);
xnor U10535 (N_10535,N_8708,N_8909);
or U10536 (N_10536,N_7636,N_8652);
xor U10537 (N_10537,N_9015,N_9253);
xor U10538 (N_10538,N_7805,N_9706);
nand U10539 (N_10539,N_8067,N_9074);
nor U10540 (N_10540,N_9054,N_8341);
or U10541 (N_10541,N_7846,N_7941);
xor U10542 (N_10542,N_8854,N_7609);
nand U10543 (N_10543,N_8147,N_9038);
and U10544 (N_10544,N_9960,N_8900);
or U10545 (N_10545,N_9447,N_9252);
and U10546 (N_10546,N_9186,N_8588);
xor U10547 (N_10547,N_7709,N_8065);
nor U10548 (N_10548,N_8231,N_8081);
or U10549 (N_10549,N_7540,N_9935);
and U10550 (N_10550,N_7803,N_8543);
nand U10551 (N_10551,N_8566,N_8851);
nor U10552 (N_10552,N_9624,N_8862);
or U10553 (N_10553,N_9414,N_8650);
nand U10554 (N_10554,N_8172,N_9947);
and U10555 (N_10555,N_9595,N_7875);
and U10556 (N_10556,N_9940,N_7648);
and U10557 (N_10557,N_8971,N_9494);
nand U10558 (N_10558,N_7613,N_8034);
xnor U10559 (N_10559,N_9797,N_9201);
and U10560 (N_10560,N_8509,N_9348);
or U10561 (N_10561,N_7887,N_7786);
xnor U10562 (N_10562,N_9131,N_8730);
xor U10563 (N_10563,N_8692,N_7906);
or U10564 (N_10564,N_8245,N_9497);
nor U10565 (N_10565,N_9528,N_8180);
xor U10566 (N_10566,N_9530,N_9326);
or U10567 (N_10567,N_9633,N_7604);
and U10568 (N_10568,N_9273,N_8699);
nor U10569 (N_10569,N_8529,N_9617);
nand U10570 (N_10570,N_9493,N_7862);
nor U10571 (N_10571,N_8060,N_8807);
nor U10572 (N_10572,N_8125,N_9426);
xnor U10573 (N_10573,N_8356,N_9794);
nand U10574 (N_10574,N_7908,N_9581);
nor U10575 (N_10575,N_9979,N_7933);
nand U10576 (N_10576,N_8527,N_8968);
or U10577 (N_10577,N_8899,N_9669);
and U10578 (N_10578,N_9126,N_8417);
nand U10579 (N_10579,N_9545,N_7692);
and U10580 (N_10580,N_9765,N_9083);
nand U10581 (N_10581,N_8059,N_9351);
and U10582 (N_10582,N_8129,N_8642);
or U10583 (N_10583,N_9185,N_9496);
and U10584 (N_10584,N_9092,N_8534);
xnor U10585 (N_10585,N_9472,N_7816);
nor U10586 (N_10586,N_7627,N_9481);
xnor U10587 (N_10587,N_9294,N_8459);
nand U10588 (N_10588,N_9539,N_9522);
nand U10589 (N_10589,N_8110,N_7770);
nand U10590 (N_10590,N_7953,N_7667);
and U10591 (N_10591,N_8307,N_7631);
nand U10592 (N_10592,N_8785,N_9491);
nor U10593 (N_10593,N_7924,N_8095);
and U10594 (N_10594,N_9286,N_9444);
nand U10595 (N_10595,N_7559,N_9842);
nor U10596 (N_10596,N_9973,N_9687);
or U10597 (N_10597,N_8240,N_9410);
nor U10598 (N_10598,N_9619,N_7976);
nand U10599 (N_10599,N_7914,N_9244);
or U10600 (N_10600,N_8096,N_7754);
or U10601 (N_10601,N_9964,N_7993);
nor U10602 (N_10602,N_8346,N_7721);
nand U10603 (N_10603,N_9945,N_9556);
nand U10604 (N_10604,N_7681,N_7766);
nor U10605 (N_10605,N_9332,N_9807);
or U10606 (N_10606,N_9380,N_8636);
nand U10607 (N_10607,N_7550,N_8961);
nor U10608 (N_10608,N_9629,N_8830);
nand U10609 (N_10609,N_9554,N_7666);
or U10610 (N_10610,N_9023,N_9319);
and U10611 (N_10611,N_9541,N_7997);
nor U10612 (N_10612,N_9848,N_7663);
nand U10613 (N_10613,N_8079,N_9914);
nand U10614 (N_10614,N_8604,N_7680);
nand U10615 (N_10615,N_9996,N_8721);
nand U10616 (N_10616,N_7662,N_9918);
nor U10617 (N_10617,N_8995,N_8037);
or U10618 (N_10618,N_8748,N_8216);
or U10619 (N_10619,N_9415,N_9082);
nor U10620 (N_10620,N_7749,N_8817);
or U10621 (N_10621,N_7671,N_8935);
or U10622 (N_10622,N_8705,N_9151);
and U10623 (N_10623,N_7579,N_9550);
nor U10624 (N_10624,N_8372,N_8916);
nor U10625 (N_10625,N_9673,N_8075);
or U10626 (N_10626,N_8826,N_8965);
and U10627 (N_10627,N_9285,N_8249);
nand U10628 (N_10628,N_9713,N_9563);
or U10629 (N_10629,N_7687,N_7843);
or U10630 (N_10630,N_8846,N_7807);
or U10631 (N_10631,N_9739,N_9784);
nor U10632 (N_10632,N_8486,N_8655);
or U10633 (N_10633,N_8028,N_8548);
and U10634 (N_10634,N_8641,N_8122);
or U10635 (N_10635,N_7619,N_7617);
or U10636 (N_10636,N_9132,N_8608);
nand U10637 (N_10637,N_8829,N_8270);
nand U10638 (N_10638,N_8796,N_9330);
and U10639 (N_10639,N_9505,N_7739);
nor U10640 (N_10640,N_7590,N_8214);
and U10641 (N_10641,N_9719,N_9953);
nor U10642 (N_10642,N_9324,N_7585);
nor U10643 (N_10643,N_8363,N_9303);
or U10644 (N_10644,N_9139,N_8894);
nand U10645 (N_10645,N_9471,N_9754);
nand U10646 (N_10646,N_9640,N_9232);
xor U10647 (N_10647,N_8277,N_8504);
and U10648 (N_10648,N_9091,N_8524);
and U10649 (N_10649,N_8922,N_9678);
nand U10650 (N_10650,N_9382,N_9150);
xor U10651 (N_10651,N_8545,N_8039);
nand U10652 (N_10652,N_8051,N_7606);
or U10653 (N_10653,N_9675,N_8804);
and U10654 (N_10654,N_8974,N_9517);
xor U10655 (N_10655,N_8165,N_9118);
xnor U10656 (N_10656,N_9033,N_9176);
nor U10657 (N_10657,N_8767,N_8954);
xor U10658 (N_10658,N_9874,N_8167);
and U10659 (N_10659,N_9561,N_8333);
nand U10660 (N_10660,N_8306,N_9019);
nand U10661 (N_10661,N_8787,N_7892);
nand U10662 (N_10662,N_8764,N_9245);
or U10663 (N_10663,N_9910,N_8229);
nand U10664 (N_10664,N_8305,N_9194);
and U10665 (N_10665,N_8467,N_9420);
xor U10666 (N_10666,N_8089,N_8603);
nor U10667 (N_10667,N_9394,N_8501);
xnor U10668 (N_10668,N_9022,N_9166);
and U10669 (N_10669,N_7601,N_8741);
and U10670 (N_10670,N_9460,N_8919);
and U10671 (N_10671,N_7780,N_8670);
nand U10672 (N_10672,N_7589,N_8135);
nand U10673 (N_10673,N_9778,N_8906);
and U10674 (N_10674,N_8976,N_7716);
and U10675 (N_10675,N_7797,N_7759);
and U10676 (N_10676,N_9021,N_9791);
and U10677 (N_10677,N_7529,N_8248);
nand U10678 (N_10678,N_8683,N_9656);
or U10679 (N_10679,N_9036,N_9331);
and U10680 (N_10680,N_7992,N_8659);
nor U10681 (N_10681,N_8123,N_8525);
xnor U10682 (N_10682,N_7556,N_7533);
or U10683 (N_10683,N_8445,N_7607);
nor U10684 (N_10684,N_9411,N_9111);
and U10685 (N_10685,N_9346,N_8038);
and U10686 (N_10686,N_8704,N_8173);
nand U10687 (N_10687,N_9296,N_8855);
and U10688 (N_10688,N_8892,N_7523);
and U10689 (N_10689,N_9125,N_8886);
or U10690 (N_10690,N_9211,N_9508);
and U10691 (N_10691,N_9365,N_9704);
or U10692 (N_10692,N_8686,N_8437);
and U10693 (N_10693,N_8927,N_8243);
nor U10694 (N_10694,N_7907,N_8441);
xnor U10695 (N_10695,N_9775,N_8066);
nor U10696 (N_10696,N_7982,N_9401);
and U10697 (N_10697,N_8878,N_9553);
or U10698 (N_10698,N_7795,N_9576);
and U10699 (N_10699,N_9792,N_9899);
nand U10700 (N_10700,N_9051,N_9202);
nand U10701 (N_10701,N_9716,N_9182);
and U10702 (N_10702,N_7831,N_7960);
nor U10703 (N_10703,N_8666,N_9752);
and U10704 (N_10704,N_8072,N_8519);
nor U10705 (N_10705,N_9225,N_9003);
nor U10706 (N_10706,N_8495,N_9119);
and U10707 (N_10707,N_9598,N_8784);
nand U10708 (N_10708,N_8177,N_8428);
or U10709 (N_10709,N_9564,N_8857);
nand U10710 (N_10710,N_7923,N_9480);
or U10711 (N_10711,N_9636,N_9572);
or U10712 (N_10712,N_9905,N_7886);
and U10713 (N_10713,N_8016,N_8197);
xnor U10714 (N_10714,N_8161,N_8150);
or U10715 (N_10715,N_7577,N_7751);
xor U10716 (N_10716,N_8706,N_9665);
and U10717 (N_10717,N_9737,N_8644);
nor U10718 (N_10718,N_7801,N_8398);
nor U10719 (N_10719,N_8115,N_7679);
xor U10720 (N_10720,N_8105,N_8873);
or U10721 (N_10721,N_8111,N_9050);
nand U10722 (N_10722,N_7768,N_8054);
or U10723 (N_10723,N_8821,N_8196);
and U10724 (N_10724,N_9944,N_8230);
nand U10725 (N_10725,N_8556,N_8040);
and U10726 (N_10726,N_7555,N_7891);
or U10727 (N_10727,N_8596,N_7819);
or U10728 (N_10728,N_7711,N_9743);
or U10729 (N_10729,N_8614,N_9398);
or U10730 (N_10730,N_9590,N_9557);
or U10731 (N_10731,N_7645,N_8097);
and U10732 (N_10732,N_7929,N_7872);
nor U10733 (N_10733,N_8572,N_8406);
and U10734 (N_10734,N_8521,N_8368);
xor U10735 (N_10735,N_9138,N_8461);
and U10736 (N_10736,N_8992,N_7547);
or U10737 (N_10737,N_8456,N_8480);
and U10738 (N_10738,N_9228,N_8751);
or U10739 (N_10739,N_8640,N_9975);
xnor U10740 (N_10740,N_8352,N_8359);
or U10741 (N_10741,N_8535,N_9804);
nor U10742 (N_10742,N_8127,N_9174);
nand U10743 (N_10743,N_9943,N_8757);
and U10744 (N_10744,N_8665,N_9866);
and U10745 (N_10745,N_8296,N_8316);
nor U10746 (N_10746,N_8109,N_7511);
and U10747 (N_10747,N_9423,N_8925);
nand U10748 (N_10748,N_9800,N_9801);
or U10749 (N_10749,N_9027,N_7515);
and U10750 (N_10750,N_9062,N_8086);
or U10751 (N_10751,N_9128,N_8334);
or U10752 (N_10752,N_8799,N_8814);
and U10753 (N_10753,N_9890,N_7625);
or U10754 (N_10754,N_7822,N_8102);
nor U10755 (N_10755,N_8958,N_9495);
xor U10756 (N_10756,N_9879,N_9223);
nand U10757 (N_10757,N_8332,N_7689);
or U10758 (N_10758,N_8325,N_8754);
nand U10759 (N_10759,N_9834,N_7854);
nand U10760 (N_10760,N_9602,N_8292);
nor U10761 (N_10761,N_9436,N_9435);
nand U10762 (N_10762,N_9011,N_7600);
or U10763 (N_10763,N_9709,N_9230);
or U10764 (N_10764,N_8266,N_8598);
or U10765 (N_10765,N_8996,N_9370);
and U10766 (N_10766,N_8179,N_9458);
nor U10767 (N_10767,N_9546,N_8226);
nor U10768 (N_10768,N_9455,N_9193);
or U10769 (N_10769,N_9383,N_8512);
xor U10770 (N_10770,N_9421,N_8790);
nor U10771 (N_10771,N_8871,N_9695);
nor U10772 (N_10772,N_9085,N_9883);
and U10773 (N_10773,N_9717,N_9210);
and U10774 (N_10774,N_8980,N_9830);
nand U10775 (N_10775,N_8653,N_9583);
or U10776 (N_10776,N_7916,N_8982);
nand U10777 (N_10777,N_8024,N_8354);
and U10778 (N_10778,N_9206,N_8936);
nor U10779 (N_10779,N_7598,N_9639);
xnor U10780 (N_10780,N_8592,N_8291);
and U10781 (N_10781,N_8585,N_8731);
and U10782 (N_10782,N_8816,N_8921);
nor U10783 (N_10783,N_9968,N_8224);
nor U10784 (N_10784,N_8910,N_9327);
nand U10785 (N_10785,N_9574,N_8513);
and U10786 (N_10786,N_9171,N_9666);
or U10787 (N_10787,N_8446,N_7624);
nor U10788 (N_10788,N_9442,N_8468);
nor U10789 (N_10789,N_8723,N_7974);
nand U10790 (N_10790,N_8531,N_9773);
and U10791 (N_10791,N_7990,N_8500);
and U10792 (N_10792,N_8702,N_9337);
nand U10793 (N_10793,N_7809,N_9142);
nand U10794 (N_10794,N_9599,N_7964);
or U10795 (N_10795,N_7567,N_9908);
nand U10796 (N_10796,N_9810,N_9731);
and U10797 (N_10797,N_7824,N_8275);
xor U10798 (N_10798,N_8671,N_9862);
nand U10799 (N_10799,N_7557,N_9732);
xnor U10800 (N_10800,N_9197,N_9075);
nor U10801 (N_10801,N_7817,N_9183);
or U10802 (N_10802,N_8503,N_7958);
or U10803 (N_10803,N_8674,N_8943);
or U10804 (N_10804,N_8210,N_9734);
or U10805 (N_10805,N_9896,N_9488);
and U10806 (N_10806,N_9181,N_9419);
or U10807 (N_10807,N_8690,N_9055);
or U10808 (N_10808,N_7977,N_9263);
nor U10809 (N_10809,N_7864,N_9570);
or U10810 (N_10810,N_8893,N_7876);
nand U10811 (N_10811,N_8843,N_9084);
nand U10812 (N_10812,N_8108,N_8419);
and U10813 (N_10813,N_7638,N_8511);
or U10814 (N_10814,N_7658,N_8776);
or U10815 (N_10815,N_9293,N_9000);
nand U10816 (N_10816,N_9991,N_7747);
or U10817 (N_10817,N_9154,N_9931);
nor U10818 (N_10818,N_9796,N_7878);
or U10819 (N_10819,N_9861,N_7845);
nand U10820 (N_10820,N_8617,N_9344);
and U10821 (N_10821,N_8498,N_7959);
nand U10822 (N_10822,N_8340,N_8064);
nor U10823 (N_10823,N_9888,N_8342);
xor U10824 (N_10824,N_7979,N_7902);
xnor U10825 (N_10825,N_7595,N_8303);
nor U10826 (N_10826,N_8082,N_7649);
and U10827 (N_10827,N_8235,N_8262);
nor U10828 (N_10828,N_9053,N_7956);
or U10829 (N_10829,N_9812,N_9468);
and U10830 (N_10830,N_9032,N_9086);
nand U10831 (N_10831,N_9544,N_7737);
nand U10832 (N_10832,N_7705,N_8438);
nand U10833 (N_10833,N_9781,N_9102);
and U10834 (N_10834,N_9025,N_8268);
and U10835 (N_10835,N_7806,N_8602);
and U10836 (N_10836,N_8820,N_8164);
and U10837 (N_10837,N_9018,N_7755);
and U10838 (N_10838,N_7718,N_7500);
or U10839 (N_10839,N_7608,N_7706);
nand U10840 (N_10840,N_8794,N_8128);
nor U10841 (N_10841,N_7910,N_9198);
nand U10842 (N_10842,N_8718,N_9680);
nand U10843 (N_10843,N_9990,N_7603);
nand U10844 (N_10844,N_9064,N_9615);
nor U10845 (N_10845,N_8901,N_8496);
xnor U10846 (N_10846,N_9347,N_7858);
or U10847 (N_10847,N_9162,N_9674);
xor U10848 (N_10848,N_9376,N_8962);
nor U10849 (N_10849,N_7629,N_8632);
xor U10850 (N_10850,N_8619,N_7724);
nor U10851 (N_10851,N_8278,N_8049);
and U10852 (N_10852,N_8310,N_8280);
and U10853 (N_10853,N_8026,N_9323);
nand U10854 (N_10854,N_7656,N_9396);
or U10855 (N_10855,N_9621,N_8290);
or U10856 (N_10856,N_8691,N_7563);
nand U10857 (N_10857,N_7694,N_8870);
or U10858 (N_10858,N_9066,N_9727);
nand U10859 (N_10859,N_9443,N_7909);
and U10860 (N_10860,N_9880,N_9721);
nor U10861 (N_10861,N_9059,N_9605);
or U10862 (N_10862,N_8885,N_8371);
xor U10863 (N_10863,N_8404,N_7558);
and U10864 (N_10864,N_8114,N_8201);
nor U10865 (N_10865,N_8139,N_9987);
and U10866 (N_10866,N_9635,N_9317);
and U10867 (N_10867,N_7842,N_9984);
nand U10868 (N_10868,N_8611,N_9412);
or U10869 (N_10869,N_7871,N_9923);
nand U10870 (N_10870,N_7969,N_9477);
or U10871 (N_10871,N_7653,N_8458);
xor U10872 (N_10872,N_9777,N_7777);
or U10873 (N_10873,N_9010,N_8405);
or U10874 (N_10874,N_8032,N_9068);
nor U10875 (N_10875,N_8162,N_7996);
and U10876 (N_10876,N_7835,N_9585);
nand U10877 (N_10877,N_9971,N_8595);
or U10878 (N_10878,N_9764,N_8227);
and U10879 (N_10879,N_8780,N_8668);
and U10880 (N_10880,N_8797,N_7788);
nor U10881 (N_10881,N_8149,N_8427);
nor U10882 (N_10882,N_9490,N_7986);
and U10883 (N_10883,N_9061,N_8088);
nand U10884 (N_10884,N_7968,N_9865);
and U10885 (N_10885,N_8637,N_9087);
xor U10886 (N_10886,N_8701,N_7927);
or U10887 (N_10887,N_7949,N_9643);
nor U10888 (N_10888,N_9512,N_8729);
nand U10889 (N_10889,N_9919,N_9088);
nor U10890 (N_10890,N_8605,N_9078);
xor U10891 (N_10891,N_8349,N_7699);
nor U10892 (N_10892,N_8031,N_7668);
nor U10893 (N_10893,N_9844,N_7874);
nor U10894 (N_10894,N_8973,N_8413);
nor U10895 (N_10895,N_8577,N_7810);
nor U10896 (N_10896,N_8926,N_9648);
or U10897 (N_10897,N_9580,N_8734);
or U10898 (N_10898,N_9196,N_8599);
nand U10899 (N_10899,N_7553,N_8522);
nand U10900 (N_10900,N_8401,N_9783);
or U10901 (N_10901,N_9725,N_9859);
and U10902 (N_10902,N_8536,N_8418);
nand U10903 (N_10903,N_9870,N_8118);
and U10904 (N_10904,N_9533,N_8422);
and U10905 (N_10905,N_8050,N_8022);
or U10906 (N_10906,N_9770,N_9994);
xor U10907 (N_10907,N_8314,N_9963);
nand U10908 (N_10908,N_8055,N_8387);
nand U10909 (N_10909,N_9895,N_8190);
nand U10910 (N_10910,N_9236,N_9305);
and U10911 (N_10911,N_9366,N_9173);
and U10912 (N_10912,N_8184,N_8408);
or U10913 (N_10913,N_8063,N_7570);
nand U10914 (N_10914,N_8932,N_8822);
nor U10915 (N_10915,N_8684,N_9855);
and U10916 (N_10916,N_8061,N_9065);
nor U10917 (N_10917,N_8399,N_9753);
nor U10918 (N_10918,N_8876,N_7541);
or U10919 (N_10919,N_9769,N_8869);
nor U10920 (N_10920,N_9780,N_8791);
nand U10921 (N_10921,N_7660,N_7509);
and U10922 (N_10922,N_7657,N_9316);
nand U10923 (N_10923,N_7918,N_9170);
nor U10924 (N_10924,N_9057,N_8750);
and U10925 (N_10925,N_9782,N_9204);
or U10926 (N_10926,N_7584,N_9771);
nor U10927 (N_10927,N_9805,N_8473);
and U10928 (N_10928,N_8786,N_9314);
nand U10929 (N_10929,N_9184,N_8448);
or U10930 (N_10930,N_9748,N_7534);
or U10931 (N_10931,N_7947,N_9168);
and U10932 (N_10932,N_8259,N_7849);
nand U10933 (N_10933,N_8007,N_9114);
or U10934 (N_10934,N_8553,N_8378);
nor U10935 (N_10935,N_8726,N_9588);
nand U10936 (N_10936,N_8389,N_8978);
nand U10937 (N_10937,N_8188,N_9871);
nor U10938 (N_10938,N_9558,N_8551);
nand U10939 (N_10939,N_7978,N_8564);
nor U10940 (N_10940,N_9847,N_8416);
and U10941 (N_10941,N_8939,N_8320);
and U10942 (N_10942,N_7895,N_8358);
xor U10943 (N_10943,N_7853,N_9261);
nor U10944 (N_10944,N_9440,N_8533);
and U10945 (N_10945,N_8845,N_7844);
nor U10946 (N_10946,N_8715,N_7799);
xor U10947 (N_10947,N_8818,N_8643);
nor U10948 (N_10948,N_8023,N_7848);
nand U10949 (N_10949,N_8710,N_8542);
nand U10950 (N_10950,N_8048,N_7961);
xor U10951 (N_10951,N_9901,N_7938);
and U10952 (N_10952,N_7688,N_9226);
xnor U10953 (N_10953,N_9761,N_8758);
nor U10954 (N_10954,N_8232,N_9395);
xor U10955 (N_10955,N_8769,N_9726);
nor U10956 (N_10956,N_7732,N_9369);
nor U10957 (N_10957,N_7855,N_9948);
or U10958 (N_10958,N_9707,N_9012);
and U10959 (N_10959,N_9568,N_8142);
nor U10960 (N_10960,N_9342,N_7873);
and U10961 (N_10961,N_9478,N_8944);
nor U10962 (N_10962,N_8107,N_8014);
or U10963 (N_10963,N_8449,N_8175);
nor U10964 (N_10964,N_9220,N_9099);
and U10965 (N_10965,N_7654,N_8739);
and U10966 (N_10966,N_8867,N_9840);
and U10967 (N_10967,N_9857,N_9799);
nor U10968 (N_10968,N_7575,N_9608);
or U10969 (N_10969,N_9825,N_7983);
and U10970 (N_10970,N_7697,N_7948);
nor U10971 (N_10971,N_8145,N_8931);
and U10972 (N_10972,N_9437,N_8434);
nand U10973 (N_10973,N_8301,N_9520);
nor U10974 (N_10974,N_9875,N_9124);
nor U10975 (N_10975,N_9813,N_8116);
nand U10976 (N_10976,N_9071,N_9270);
nor U10977 (N_10977,N_9637,N_8987);
or U10978 (N_10978,N_9681,N_9900);
nor U10979 (N_10979,N_8176,N_9329);
nand U10980 (N_10980,N_7790,N_8098);
and U10981 (N_10981,N_8896,N_9742);
xnor U10982 (N_10982,N_8661,N_9307);
xor U10983 (N_10983,N_9105,N_9262);
nor U10984 (N_10984,N_9430,N_9646);
and U10985 (N_10985,N_8185,N_7538);
and U10986 (N_10986,N_9219,N_8299);
and U10987 (N_10987,N_9525,N_7774);
or U10988 (N_10988,N_7861,N_8613);
nand U10989 (N_10989,N_8103,N_9007);
nor U10990 (N_10990,N_8423,N_7677);
nor U10991 (N_10991,N_9653,N_9938);
nor U10992 (N_10992,N_8008,N_8606);
and U10993 (N_10993,N_7951,N_7913);
nand U10994 (N_10994,N_9137,N_9165);
nor U10995 (N_10995,N_7568,N_9965);
nand U10996 (N_10996,N_9826,N_9664);
or U10997 (N_10997,N_9757,N_7837);
nand U10998 (N_10998,N_8678,N_8724);
nor U10999 (N_10999,N_8124,N_9006);
and U11000 (N_11000,N_9683,N_8907);
and U11001 (N_11001,N_8554,N_9116);
or U11002 (N_11002,N_9046,N_8106);
xnor U11003 (N_11003,N_9552,N_8569);
or U11004 (N_11004,N_9360,N_9772);
nand U11005 (N_11005,N_9970,N_8887);
nand U11006 (N_11006,N_7866,N_8913);
nand U11007 (N_11007,N_7771,N_7701);
and U11008 (N_11008,N_8942,N_9798);
xor U11009 (N_11009,N_9756,N_8012);
and U11010 (N_11010,N_7670,N_9569);
nand U11011 (N_11011,N_9216,N_8840);
and U11012 (N_11012,N_9474,N_8400);
or U11013 (N_11013,N_8972,N_8753);
or U11014 (N_11014,N_7611,N_8252);
or U11015 (N_11015,N_8112,N_8329);
or U11016 (N_11016,N_9897,N_9720);
nor U11017 (N_11017,N_7530,N_7714);
nand U11018 (N_11018,N_9121,N_7597);
and U11019 (N_11019,N_9243,N_8025);
nor U11020 (N_11020,N_9179,N_9362);
or U11021 (N_11021,N_8120,N_7635);
and U11022 (N_11022,N_9543,N_8151);
and U11023 (N_11023,N_9290,N_8584);
nand U11024 (N_11024,N_8390,N_9482);
and U11025 (N_11025,N_8571,N_7863);
xor U11026 (N_11026,N_8898,N_8272);
nand U11027 (N_11027,N_8355,N_9954);
nor U11028 (N_11028,N_8677,N_9696);
or U11029 (N_11029,N_9515,N_9571);
nor U11030 (N_11030,N_9004,N_7870);
nand U11031 (N_11031,N_7869,N_9926);
nor U11032 (N_11032,N_9638,N_8868);
nor U11033 (N_11033,N_9622,N_7943);
or U11034 (N_11034,N_7764,N_7836);
nand U11035 (N_11035,N_8882,N_7513);
nand U11036 (N_11036,N_8000,N_9418);
nand U11037 (N_11037,N_9144,N_9594);
or U11038 (N_11038,N_8431,N_9276);
and U11039 (N_11039,N_8696,N_9506);
and U11040 (N_11040,N_7708,N_9320);
nor U11041 (N_11041,N_9391,N_7622);
nand U11042 (N_11042,N_8517,N_9287);
nand U11043 (N_11043,N_7583,N_7840);
xor U11044 (N_11044,N_7899,N_8357);
nor U11045 (N_11045,N_9432,N_9815);
nor U11046 (N_11046,N_9946,N_8460);
xor U11047 (N_11047,N_7893,N_8777);
and U11048 (N_11048,N_8488,N_8772);
nor U11049 (N_11049,N_9461,N_9429);
and U11050 (N_11050,N_9189,N_9831);
nand U11051 (N_11051,N_9790,N_9450);
or U11052 (N_11052,N_8258,N_8880);
and U11053 (N_11053,N_9122,N_7621);
nor U11054 (N_11054,N_9524,N_9668);
nor U11055 (N_11055,N_9913,N_8833);
or U11056 (N_11056,N_8712,N_7794);
xnor U11057 (N_11057,N_9956,N_9178);
nand U11058 (N_11058,N_9845,N_7888);
nand U11059 (N_11059,N_7569,N_9542);
or U11060 (N_11060,N_8628,N_9115);
nand U11061 (N_11061,N_9328,N_7522);
nand U11062 (N_11062,N_9127,N_8703);
or U11063 (N_11063,N_9045,N_8747);
nand U11064 (N_11064,N_8789,N_7850);
and U11065 (N_11065,N_7650,N_9700);
and U11066 (N_11066,N_8464,N_9565);
and U11067 (N_11067,N_9630,N_7827);
nor U11068 (N_11068,N_7926,N_8132);
or U11069 (N_11069,N_9345,N_9254);
and U11070 (N_11070,N_8169,N_8030);
or U11071 (N_11071,N_8271,N_8654);
or U11072 (N_11072,N_8890,N_9917);
xor U11073 (N_11073,N_9822,N_7727);
nand U11074 (N_11074,N_8615,N_9343);
xor U11075 (N_11075,N_8550,N_8002);
nor U11076 (N_11076,N_9738,N_9631);
and U11077 (N_11077,N_9229,N_8440);
or U11078 (N_11078,N_7738,N_8634);
and U11079 (N_11079,N_8966,N_9872);
and U11080 (N_11080,N_8104,N_7728);
or U11081 (N_11081,N_9950,N_8956);
nor U11082 (N_11082,N_9909,N_9295);
nor U11083 (N_11083,N_8664,N_9389);
nand U11084 (N_11084,N_9237,N_8377);
nand U11085 (N_11085,N_9385,N_9315);
or U11086 (N_11086,N_8174,N_8191);
nor U11087 (N_11087,N_9521,N_9744);
nand U11088 (N_11088,N_8557,N_8832);
or U11089 (N_11089,N_8313,N_9603);
nor U11090 (N_11090,N_8029,N_9977);
nor U11091 (N_11091,N_8808,N_9586);
nor U11092 (N_11092,N_7592,N_7722);
and U11093 (N_11093,N_8004,N_9467);
nand U11094 (N_11094,N_9957,N_8763);
or U11095 (N_11095,N_8760,N_8415);
xor U11096 (N_11096,N_9409,N_7507);
or U11097 (N_11097,N_9623,N_8068);
nor U11098 (N_11098,N_8506,N_7877);
and U11099 (N_11099,N_8711,N_7634);
xor U11100 (N_11100,N_8801,N_8959);
xor U11101 (N_11101,N_9686,N_9424);
xor U11102 (N_11102,N_8084,N_8673);
or U11103 (N_11103,N_8515,N_9951);
or U11104 (N_11104,N_9655,N_8745);
and U11105 (N_11105,N_7963,N_7548);
or U11106 (N_11106,N_8141,N_8432);
and U11107 (N_11107,N_9672,N_8812);
nor U11108 (N_11108,N_9499,N_8578);
xnor U11109 (N_11109,N_9392,N_8623);
or U11110 (N_11110,N_9662,N_9473);
nand U11111 (N_11111,N_8510,N_7643);
and U11112 (N_11112,N_9980,N_9259);
xor U11113 (N_11113,N_9157,N_9999);
and U11114 (N_11114,N_8895,N_9682);
nor U11115 (N_11115,N_8298,N_9167);
nand U11116 (N_11116,N_7830,N_8819);
nand U11117 (N_11117,N_9227,N_9190);
nand U11118 (N_11118,N_8225,N_9017);
or U11119 (N_11119,N_9670,N_8866);
or U11120 (N_11120,N_9766,N_7733);
or U11121 (N_11121,N_8575,N_8353);
or U11122 (N_11122,N_9340,N_9779);
nand U11123 (N_11123,N_8044,N_8502);
and U11124 (N_11124,N_9697,N_9282);
nor U11125 (N_11125,N_9058,N_8680);
xnor U11126 (N_11126,N_9527,N_8293);
nor U11127 (N_11127,N_9729,N_8452);
and U11128 (N_11128,N_8888,N_8485);
or U11129 (N_11129,N_8938,N_9593);
nor U11130 (N_11130,N_8679,N_7760);
and U11131 (N_11131,N_9280,N_8610);
nand U11132 (N_11132,N_8802,N_9578);
xor U11133 (N_11133,N_8687,N_7930);
xor U11134 (N_11134,N_8858,N_8492);
or U11135 (N_11135,N_7573,N_8879);
nor U11136 (N_11136,N_9736,N_7524);
and U11137 (N_11137,N_8951,N_8041);
and U11138 (N_11138,N_7743,N_7796);
nor U11139 (N_11139,N_7756,N_7546);
or U11140 (N_11140,N_9758,N_9966);
and U11141 (N_11141,N_9843,N_7989);
and U11142 (N_11142,N_8140,N_9537);
and U11143 (N_11143,N_9856,N_9876);
or U11144 (N_11144,N_7769,N_9763);
or U11145 (N_11145,N_8693,N_8146);
or U11146 (N_11146,N_9417,N_8160);
nor U11147 (N_11147,N_8052,N_7735);
or U11148 (N_11148,N_9767,N_7717);
and U11149 (N_11149,N_9072,N_9922);
nor U11150 (N_11150,N_8080,N_7860);
or U11151 (N_11151,N_9566,N_7815);
nor U11152 (N_11152,N_9776,N_8076);
and U11153 (N_11153,N_9479,N_9445);
nand U11154 (N_11154,N_9747,N_8283);
nor U11155 (N_11155,N_9215,N_7950);
or U11156 (N_11156,N_8255,N_9827);
and U11157 (N_11157,N_8043,N_8260);
nand U11158 (N_11158,N_8589,N_9601);
nor U11159 (N_11159,N_9177,N_7890);
nor U11160 (N_11160,N_8576,N_9823);
or U11161 (N_11161,N_8143,N_9378);
nor U11162 (N_11162,N_8375,N_9892);
and U11163 (N_11163,N_9306,N_8957);
or U11164 (N_11164,N_9838,N_9278);
xnor U11165 (N_11165,N_8447,N_9832);
xnor U11166 (N_11166,N_9152,N_9942);
nand U11167 (N_11167,N_9885,N_9645);
xnor U11168 (N_11168,N_8947,N_7900);
nor U11169 (N_11169,N_9163,N_9837);
xnor U11170 (N_11170,N_8326,N_7944);
nor U11171 (N_11171,N_8207,N_8563);
and U11172 (N_11172,N_8838,N_9029);
or U11173 (N_11173,N_9076,N_9625);
or U11174 (N_11174,N_8279,N_8345);
or U11175 (N_11175,N_8681,N_9983);
nor U11176 (N_11176,N_8918,N_8121);
or U11177 (N_11177,N_7669,N_8070);
and U11178 (N_11178,N_9310,N_9851);
and U11179 (N_11179,N_8590,N_8539);
nor U11180 (N_11180,N_8133,N_8494);
and U11181 (N_11181,N_7545,N_7571);
nor U11182 (N_11182,N_8847,N_9301);
xor U11183 (N_11183,N_8181,N_9110);
nor U11184 (N_11184,N_9248,N_7945);
and U11185 (N_11185,N_8113,N_9982);
nand U11186 (N_11186,N_8667,N_9298);
and U11187 (N_11187,N_9969,N_9433);
and U11188 (N_11188,N_9397,N_8902);
xnor U11189 (N_11189,N_9661,N_7920);
nand U11190 (N_11190,N_8171,N_8929);
or U11191 (N_11191,N_7503,N_9634);
nand U11192 (N_11192,N_9839,N_8620);
nand U11193 (N_11193,N_8267,N_7940);
nor U11194 (N_11194,N_9242,N_9873);
or U11195 (N_11195,N_9040,N_7736);
nor U11196 (N_11196,N_8813,N_9106);
and U11197 (N_11197,N_9288,N_8393);
nand U11198 (N_11198,N_7655,N_9501);
or U11199 (N_11199,N_7765,N_8489);
nor U11200 (N_11200,N_8788,N_9014);
xor U11201 (N_11201,N_8284,N_7911);
or U11202 (N_11202,N_9147,N_9745);
and U11203 (N_11203,N_8573,N_9476);
xor U11204 (N_11204,N_9699,N_8544);
or U11205 (N_11205,N_7512,N_9260);
nor U11206 (N_11206,N_9212,N_8960);
xnor U11207 (N_11207,N_8770,N_9891);
nand U11208 (N_11208,N_9600,N_9929);
or U11209 (N_11209,N_8587,N_8078);
nor U11210 (N_11210,N_8969,N_8698);
xnor U11211 (N_11211,N_9020,N_9379);
and U11212 (N_11212,N_8153,N_9562);
and U11213 (N_11213,N_9684,N_8848);
and U11214 (N_11214,N_9034,N_8844);
or U11215 (N_11215,N_9133,N_7726);
nand U11216 (N_11216,N_9041,N_8322);
or U11217 (N_11217,N_8021,N_8330);
nor U11218 (N_11218,N_7779,N_7917);
and U11219 (N_11219,N_9628,N_8273);
nor U11220 (N_11220,N_8558,N_9644);
and U11221 (N_11221,N_9405,N_8337);
xnor U11222 (N_11222,N_8493,N_9169);
xor U11223 (N_11223,N_9318,N_8166);
nand U11224 (N_11224,N_8009,N_9214);
xor U11225 (N_11225,N_9028,N_8523);
nand U11226 (N_11226,N_8444,N_9428);
nand U11227 (N_11227,N_9589,N_9265);
or U11228 (N_11228,N_9207,N_8466);
nand U11229 (N_11229,N_7868,N_8212);
nand U11230 (N_11230,N_7549,N_7984);
nand U11231 (N_11231,N_8130,N_8157);
nor U11232 (N_11232,N_9192,N_8453);
xor U11233 (N_11233,N_9081,N_7605);
nand U11234 (N_11234,N_7505,N_8881);
nand U11235 (N_11235,N_7814,N_7833);
xor U11236 (N_11236,N_9616,N_7970);
nor U11237 (N_11237,N_9511,N_8774);
and U11238 (N_11238,N_9096,N_8211);
nand U11239 (N_11239,N_9992,N_7748);
nor U11240 (N_11240,N_9095,N_8300);
xnor U11241 (N_11241,N_9967,N_7594);
or U11242 (N_11242,N_8979,N_7750);
nand U11243 (N_11243,N_9341,N_9903);
nand U11244 (N_11244,N_9255,N_9714);
and U11245 (N_11245,N_8950,N_7676);
nand U11246 (N_11246,N_9852,N_8737);
and U11247 (N_11247,N_9393,N_8839);
or U11248 (N_11248,N_9534,N_9548);
or U11249 (N_11249,N_8795,N_9934);
and U11250 (N_11250,N_9044,N_7876);
and U11251 (N_11251,N_8489,N_9619);
or U11252 (N_11252,N_9076,N_8780);
nor U11253 (N_11253,N_8113,N_9738);
nor U11254 (N_11254,N_9943,N_9493);
and U11255 (N_11255,N_9685,N_9810);
xnor U11256 (N_11256,N_7649,N_9413);
nor U11257 (N_11257,N_9874,N_9785);
nor U11258 (N_11258,N_8157,N_8766);
nor U11259 (N_11259,N_9971,N_8982);
and U11260 (N_11260,N_9513,N_9386);
or U11261 (N_11261,N_9479,N_9021);
and U11262 (N_11262,N_8829,N_9963);
or U11263 (N_11263,N_9303,N_8314);
or U11264 (N_11264,N_7779,N_9360);
and U11265 (N_11265,N_8788,N_9645);
and U11266 (N_11266,N_9700,N_9940);
and U11267 (N_11267,N_8094,N_7734);
nor U11268 (N_11268,N_9247,N_8977);
and U11269 (N_11269,N_9236,N_7830);
xor U11270 (N_11270,N_7978,N_7553);
xnor U11271 (N_11271,N_7941,N_7634);
xor U11272 (N_11272,N_9166,N_8037);
and U11273 (N_11273,N_9028,N_8862);
nor U11274 (N_11274,N_8985,N_9128);
or U11275 (N_11275,N_9948,N_9134);
and U11276 (N_11276,N_9122,N_8682);
or U11277 (N_11277,N_7606,N_8669);
or U11278 (N_11278,N_9628,N_8679);
nand U11279 (N_11279,N_8150,N_7969);
nand U11280 (N_11280,N_7662,N_9256);
xnor U11281 (N_11281,N_7816,N_7516);
and U11282 (N_11282,N_8040,N_7515);
and U11283 (N_11283,N_8386,N_9538);
nor U11284 (N_11284,N_8607,N_9557);
or U11285 (N_11285,N_8253,N_7525);
nand U11286 (N_11286,N_9012,N_8392);
or U11287 (N_11287,N_9423,N_9273);
and U11288 (N_11288,N_7862,N_8450);
xor U11289 (N_11289,N_7665,N_7513);
nand U11290 (N_11290,N_9374,N_8745);
or U11291 (N_11291,N_8571,N_9468);
nand U11292 (N_11292,N_8982,N_8574);
and U11293 (N_11293,N_8509,N_9119);
xnor U11294 (N_11294,N_8607,N_9360);
xor U11295 (N_11295,N_7618,N_7945);
and U11296 (N_11296,N_9991,N_8560);
or U11297 (N_11297,N_7997,N_9856);
or U11298 (N_11298,N_9186,N_7888);
nand U11299 (N_11299,N_8136,N_7939);
xnor U11300 (N_11300,N_9402,N_9234);
or U11301 (N_11301,N_8334,N_9482);
nand U11302 (N_11302,N_9512,N_8072);
nand U11303 (N_11303,N_8226,N_8734);
and U11304 (N_11304,N_7792,N_8292);
nand U11305 (N_11305,N_9619,N_9218);
and U11306 (N_11306,N_7571,N_9550);
nand U11307 (N_11307,N_9185,N_8427);
nand U11308 (N_11308,N_9758,N_7609);
xnor U11309 (N_11309,N_7873,N_9596);
nor U11310 (N_11310,N_8662,N_8552);
nand U11311 (N_11311,N_8516,N_9979);
and U11312 (N_11312,N_8101,N_7994);
or U11313 (N_11313,N_9262,N_9195);
xnor U11314 (N_11314,N_7790,N_8880);
and U11315 (N_11315,N_8958,N_9691);
or U11316 (N_11316,N_8972,N_9707);
nand U11317 (N_11317,N_9930,N_9445);
nor U11318 (N_11318,N_9547,N_8822);
nand U11319 (N_11319,N_8400,N_9893);
or U11320 (N_11320,N_7782,N_9763);
nand U11321 (N_11321,N_8399,N_7704);
nand U11322 (N_11322,N_7843,N_7768);
or U11323 (N_11323,N_9196,N_8014);
nor U11324 (N_11324,N_8097,N_9769);
xor U11325 (N_11325,N_9070,N_9900);
and U11326 (N_11326,N_8662,N_8425);
xor U11327 (N_11327,N_8223,N_7659);
or U11328 (N_11328,N_9667,N_7962);
or U11329 (N_11329,N_8238,N_9753);
and U11330 (N_11330,N_7968,N_8140);
or U11331 (N_11331,N_9367,N_8344);
nand U11332 (N_11332,N_7534,N_8767);
xnor U11333 (N_11333,N_9127,N_7786);
nor U11334 (N_11334,N_8402,N_7942);
and U11335 (N_11335,N_8141,N_8888);
xor U11336 (N_11336,N_8484,N_8302);
nand U11337 (N_11337,N_8153,N_9579);
or U11338 (N_11338,N_7783,N_9859);
or U11339 (N_11339,N_9113,N_9160);
and U11340 (N_11340,N_7985,N_9441);
nand U11341 (N_11341,N_8958,N_8157);
nand U11342 (N_11342,N_7618,N_9673);
nor U11343 (N_11343,N_7814,N_8311);
nand U11344 (N_11344,N_8741,N_9876);
or U11345 (N_11345,N_9685,N_8881);
nand U11346 (N_11346,N_9396,N_8012);
or U11347 (N_11347,N_9635,N_8510);
or U11348 (N_11348,N_9296,N_9236);
and U11349 (N_11349,N_8747,N_8659);
or U11350 (N_11350,N_9730,N_8083);
and U11351 (N_11351,N_9991,N_9256);
xor U11352 (N_11352,N_9014,N_8564);
nand U11353 (N_11353,N_8857,N_7967);
nand U11354 (N_11354,N_9014,N_7624);
or U11355 (N_11355,N_8009,N_8970);
nand U11356 (N_11356,N_7771,N_8095);
nand U11357 (N_11357,N_7607,N_8707);
and U11358 (N_11358,N_9593,N_8072);
nand U11359 (N_11359,N_8286,N_9252);
nand U11360 (N_11360,N_9269,N_8649);
nand U11361 (N_11361,N_8841,N_9792);
nand U11362 (N_11362,N_9794,N_7790);
or U11363 (N_11363,N_8457,N_8446);
and U11364 (N_11364,N_9904,N_9853);
and U11365 (N_11365,N_7655,N_7747);
and U11366 (N_11366,N_9482,N_9832);
or U11367 (N_11367,N_9349,N_9558);
nand U11368 (N_11368,N_9178,N_7911);
nand U11369 (N_11369,N_9763,N_9828);
nor U11370 (N_11370,N_8260,N_9022);
nand U11371 (N_11371,N_8505,N_8685);
nor U11372 (N_11372,N_8634,N_8639);
and U11373 (N_11373,N_8944,N_8965);
and U11374 (N_11374,N_9472,N_8167);
or U11375 (N_11375,N_9541,N_8190);
or U11376 (N_11376,N_9424,N_8019);
and U11377 (N_11377,N_8909,N_9452);
and U11378 (N_11378,N_8739,N_9683);
nor U11379 (N_11379,N_8159,N_8459);
and U11380 (N_11380,N_7588,N_9800);
and U11381 (N_11381,N_7698,N_8485);
and U11382 (N_11382,N_9301,N_9599);
or U11383 (N_11383,N_9749,N_8625);
and U11384 (N_11384,N_8290,N_7583);
nand U11385 (N_11385,N_8248,N_8808);
or U11386 (N_11386,N_8819,N_8190);
and U11387 (N_11387,N_7620,N_7673);
and U11388 (N_11388,N_7660,N_7539);
nand U11389 (N_11389,N_9838,N_9202);
nand U11390 (N_11390,N_9389,N_9850);
nor U11391 (N_11391,N_9350,N_8924);
and U11392 (N_11392,N_9261,N_8808);
and U11393 (N_11393,N_8095,N_8569);
or U11394 (N_11394,N_8318,N_7555);
xor U11395 (N_11395,N_8415,N_9159);
xor U11396 (N_11396,N_9896,N_7626);
nand U11397 (N_11397,N_7954,N_8326);
nor U11398 (N_11398,N_9624,N_9127);
nor U11399 (N_11399,N_9760,N_9230);
nand U11400 (N_11400,N_9521,N_9967);
or U11401 (N_11401,N_9600,N_8565);
and U11402 (N_11402,N_8694,N_7975);
nor U11403 (N_11403,N_8401,N_7707);
or U11404 (N_11404,N_8760,N_8109);
nand U11405 (N_11405,N_9145,N_8405);
and U11406 (N_11406,N_8984,N_8229);
xor U11407 (N_11407,N_8112,N_9001);
nor U11408 (N_11408,N_8915,N_8326);
and U11409 (N_11409,N_7537,N_9879);
and U11410 (N_11410,N_9223,N_8914);
or U11411 (N_11411,N_8800,N_8614);
or U11412 (N_11412,N_7536,N_8566);
or U11413 (N_11413,N_8582,N_9186);
nor U11414 (N_11414,N_8821,N_9065);
nand U11415 (N_11415,N_7611,N_8544);
nand U11416 (N_11416,N_8229,N_9353);
and U11417 (N_11417,N_8210,N_8076);
nor U11418 (N_11418,N_8276,N_9508);
nor U11419 (N_11419,N_9981,N_7842);
nor U11420 (N_11420,N_7835,N_8971);
and U11421 (N_11421,N_9619,N_9591);
and U11422 (N_11422,N_9069,N_9915);
and U11423 (N_11423,N_8378,N_9298);
nand U11424 (N_11424,N_9732,N_8372);
and U11425 (N_11425,N_9504,N_9246);
and U11426 (N_11426,N_8566,N_9751);
and U11427 (N_11427,N_7642,N_8159);
nor U11428 (N_11428,N_9412,N_7584);
nand U11429 (N_11429,N_7608,N_8710);
or U11430 (N_11430,N_9313,N_9401);
nor U11431 (N_11431,N_8972,N_7765);
and U11432 (N_11432,N_7756,N_9083);
nor U11433 (N_11433,N_7672,N_9023);
nor U11434 (N_11434,N_8275,N_9007);
or U11435 (N_11435,N_7638,N_7880);
xor U11436 (N_11436,N_8665,N_8743);
nand U11437 (N_11437,N_8367,N_8777);
nor U11438 (N_11438,N_9145,N_7616);
or U11439 (N_11439,N_8037,N_9546);
or U11440 (N_11440,N_8213,N_7506);
nor U11441 (N_11441,N_9959,N_8267);
and U11442 (N_11442,N_8776,N_7714);
and U11443 (N_11443,N_9609,N_7538);
nand U11444 (N_11444,N_7976,N_9898);
nand U11445 (N_11445,N_8431,N_9775);
nor U11446 (N_11446,N_8271,N_8930);
nand U11447 (N_11447,N_9402,N_8781);
and U11448 (N_11448,N_7554,N_8826);
and U11449 (N_11449,N_8294,N_7828);
xor U11450 (N_11450,N_7999,N_9647);
and U11451 (N_11451,N_7814,N_9697);
nor U11452 (N_11452,N_7560,N_8725);
nor U11453 (N_11453,N_7514,N_8556);
xnor U11454 (N_11454,N_9570,N_9983);
and U11455 (N_11455,N_8522,N_7568);
or U11456 (N_11456,N_8096,N_8912);
nor U11457 (N_11457,N_7749,N_9250);
nor U11458 (N_11458,N_7551,N_8674);
and U11459 (N_11459,N_8307,N_8243);
nor U11460 (N_11460,N_8968,N_9678);
nor U11461 (N_11461,N_9523,N_9736);
or U11462 (N_11462,N_9909,N_8363);
nand U11463 (N_11463,N_8404,N_8119);
nor U11464 (N_11464,N_9715,N_8219);
and U11465 (N_11465,N_7561,N_9551);
or U11466 (N_11466,N_7986,N_9669);
and U11467 (N_11467,N_8421,N_7862);
nor U11468 (N_11468,N_9067,N_9128);
and U11469 (N_11469,N_8835,N_7868);
or U11470 (N_11470,N_8571,N_9186);
nor U11471 (N_11471,N_9625,N_8963);
xor U11472 (N_11472,N_7997,N_9359);
nor U11473 (N_11473,N_9433,N_9706);
nand U11474 (N_11474,N_8932,N_8836);
and U11475 (N_11475,N_9488,N_7552);
nor U11476 (N_11476,N_7517,N_9162);
and U11477 (N_11477,N_9951,N_7822);
and U11478 (N_11478,N_9244,N_8678);
or U11479 (N_11479,N_8748,N_8413);
xnor U11480 (N_11480,N_8897,N_7659);
and U11481 (N_11481,N_9471,N_9455);
nand U11482 (N_11482,N_9063,N_7983);
nand U11483 (N_11483,N_9833,N_9432);
xor U11484 (N_11484,N_8443,N_9190);
and U11485 (N_11485,N_9195,N_9805);
or U11486 (N_11486,N_9029,N_8778);
nor U11487 (N_11487,N_8767,N_8265);
xnor U11488 (N_11488,N_7927,N_9492);
nand U11489 (N_11489,N_8971,N_9716);
and U11490 (N_11490,N_8482,N_9254);
or U11491 (N_11491,N_7563,N_8398);
xor U11492 (N_11492,N_9571,N_8501);
nand U11493 (N_11493,N_9859,N_7861);
nor U11494 (N_11494,N_9498,N_7988);
xor U11495 (N_11495,N_7700,N_8305);
or U11496 (N_11496,N_8414,N_8285);
and U11497 (N_11497,N_8524,N_7973);
or U11498 (N_11498,N_8435,N_9356);
nor U11499 (N_11499,N_9531,N_7830);
and U11500 (N_11500,N_8333,N_8560);
or U11501 (N_11501,N_8226,N_9031);
or U11502 (N_11502,N_8538,N_8062);
nor U11503 (N_11503,N_9776,N_9291);
or U11504 (N_11504,N_9764,N_8166);
or U11505 (N_11505,N_9863,N_8422);
and U11506 (N_11506,N_7844,N_8907);
and U11507 (N_11507,N_9486,N_9926);
nand U11508 (N_11508,N_8240,N_9533);
and U11509 (N_11509,N_8571,N_7638);
nand U11510 (N_11510,N_9977,N_8708);
nand U11511 (N_11511,N_8773,N_9752);
nor U11512 (N_11512,N_8256,N_8060);
nor U11513 (N_11513,N_9592,N_7637);
and U11514 (N_11514,N_8060,N_9603);
nor U11515 (N_11515,N_9123,N_7613);
nor U11516 (N_11516,N_9417,N_8625);
nand U11517 (N_11517,N_9993,N_7530);
nand U11518 (N_11518,N_8376,N_7679);
nand U11519 (N_11519,N_7561,N_8501);
or U11520 (N_11520,N_9798,N_9988);
and U11521 (N_11521,N_8984,N_9889);
nand U11522 (N_11522,N_8444,N_7653);
or U11523 (N_11523,N_9273,N_8710);
nand U11524 (N_11524,N_9958,N_8581);
and U11525 (N_11525,N_8941,N_7970);
and U11526 (N_11526,N_8888,N_8459);
and U11527 (N_11527,N_9592,N_9116);
xnor U11528 (N_11528,N_9341,N_9794);
or U11529 (N_11529,N_8826,N_8204);
xor U11530 (N_11530,N_9170,N_9187);
and U11531 (N_11531,N_8453,N_9845);
nand U11532 (N_11532,N_7634,N_9620);
nor U11533 (N_11533,N_7774,N_7512);
nand U11534 (N_11534,N_8186,N_7644);
or U11535 (N_11535,N_9494,N_9363);
nand U11536 (N_11536,N_8815,N_8219);
xnor U11537 (N_11537,N_8580,N_8959);
nor U11538 (N_11538,N_7632,N_9439);
xor U11539 (N_11539,N_8650,N_9657);
nor U11540 (N_11540,N_9296,N_9298);
and U11541 (N_11541,N_9624,N_9722);
nor U11542 (N_11542,N_9915,N_9838);
or U11543 (N_11543,N_8805,N_9557);
nand U11544 (N_11544,N_9746,N_8779);
xor U11545 (N_11545,N_8327,N_9953);
nand U11546 (N_11546,N_9167,N_8229);
or U11547 (N_11547,N_9734,N_9693);
and U11548 (N_11548,N_9025,N_9654);
nand U11549 (N_11549,N_9754,N_8371);
and U11550 (N_11550,N_9144,N_9451);
nand U11551 (N_11551,N_8742,N_9962);
nand U11552 (N_11552,N_8243,N_7927);
and U11553 (N_11553,N_9188,N_7717);
or U11554 (N_11554,N_9149,N_8492);
or U11555 (N_11555,N_9059,N_9774);
nor U11556 (N_11556,N_9515,N_7631);
and U11557 (N_11557,N_9036,N_9397);
and U11558 (N_11558,N_7923,N_8654);
or U11559 (N_11559,N_7940,N_8788);
nand U11560 (N_11560,N_9036,N_7576);
or U11561 (N_11561,N_8424,N_8011);
or U11562 (N_11562,N_8475,N_9728);
or U11563 (N_11563,N_9305,N_8910);
and U11564 (N_11564,N_9862,N_8915);
or U11565 (N_11565,N_8708,N_9997);
nand U11566 (N_11566,N_7667,N_9279);
and U11567 (N_11567,N_9464,N_9157);
nand U11568 (N_11568,N_7674,N_7514);
nand U11569 (N_11569,N_9668,N_9196);
nor U11570 (N_11570,N_8825,N_8031);
xor U11571 (N_11571,N_9301,N_8316);
and U11572 (N_11572,N_8807,N_9102);
nor U11573 (N_11573,N_9830,N_7985);
nor U11574 (N_11574,N_9537,N_9897);
nor U11575 (N_11575,N_9727,N_7890);
and U11576 (N_11576,N_9700,N_9779);
nand U11577 (N_11577,N_9166,N_8323);
or U11578 (N_11578,N_7530,N_9320);
nand U11579 (N_11579,N_9551,N_8960);
nor U11580 (N_11580,N_9240,N_8354);
or U11581 (N_11581,N_8061,N_8141);
and U11582 (N_11582,N_9258,N_7977);
nor U11583 (N_11583,N_7994,N_7755);
nand U11584 (N_11584,N_8056,N_8280);
nor U11585 (N_11585,N_7746,N_9348);
and U11586 (N_11586,N_9490,N_9872);
nand U11587 (N_11587,N_8588,N_8247);
xor U11588 (N_11588,N_9663,N_8979);
and U11589 (N_11589,N_9827,N_9691);
nand U11590 (N_11590,N_9340,N_9073);
nor U11591 (N_11591,N_8591,N_7777);
nand U11592 (N_11592,N_9361,N_8164);
nand U11593 (N_11593,N_9494,N_9313);
or U11594 (N_11594,N_8779,N_8080);
nand U11595 (N_11595,N_9850,N_7861);
and U11596 (N_11596,N_9452,N_9707);
and U11597 (N_11597,N_9571,N_8449);
or U11598 (N_11598,N_7883,N_7567);
xnor U11599 (N_11599,N_8153,N_9587);
nand U11600 (N_11600,N_9059,N_8232);
nor U11601 (N_11601,N_9263,N_9135);
nor U11602 (N_11602,N_9517,N_8657);
nor U11603 (N_11603,N_8342,N_8231);
or U11604 (N_11604,N_9028,N_8722);
nor U11605 (N_11605,N_7867,N_7897);
nor U11606 (N_11606,N_8781,N_7935);
and U11607 (N_11607,N_9413,N_8316);
nor U11608 (N_11608,N_9860,N_9510);
and U11609 (N_11609,N_9246,N_9043);
and U11610 (N_11610,N_9584,N_8221);
xnor U11611 (N_11611,N_7853,N_7896);
or U11612 (N_11612,N_7954,N_7829);
or U11613 (N_11613,N_9929,N_8875);
nand U11614 (N_11614,N_7544,N_8583);
nand U11615 (N_11615,N_9245,N_7823);
and U11616 (N_11616,N_9397,N_9326);
or U11617 (N_11617,N_9532,N_8509);
and U11618 (N_11618,N_9356,N_8941);
nor U11619 (N_11619,N_8901,N_9124);
and U11620 (N_11620,N_8028,N_9025);
and U11621 (N_11621,N_9051,N_7872);
nor U11622 (N_11622,N_7549,N_7816);
nor U11623 (N_11623,N_7891,N_8706);
nor U11624 (N_11624,N_7919,N_8385);
nor U11625 (N_11625,N_8407,N_9773);
or U11626 (N_11626,N_9775,N_8740);
and U11627 (N_11627,N_8507,N_8156);
or U11628 (N_11628,N_9549,N_7816);
or U11629 (N_11629,N_8228,N_7955);
or U11630 (N_11630,N_8248,N_7550);
nor U11631 (N_11631,N_9113,N_9304);
nor U11632 (N_11632,N_7860,N_9866);
or U11633 (N_11633,N_8598,N_9709);
xnor U11634 (N_11634,N_8631,N_7676);
and U11635 (N_11635,N_8393,N_9355);
and U11636 (N_11636,N_8698,N_9349);
and U11637 (N_11637,N_8059,N_8721);
or U11638 (N_11638,N_9467,N_9972);
or U11639 (N_11639,N_9302,N_7937);
and U11640 (N_11640,N_8391,N_7674);
nor U11641 (N_11641,N_8451,N_8980);
and U11642 (N_11642,N_9480,N_9197);
and U11643 (N_11643,N_7770,N_9259);
nand U11644 (N_11644,N_8237,N_8403);
or U11645 (N_11645,N_8729,N_7551);
or U11646 (N_11646,N_9640,N_8799);
or U11647 (N_11647,N_7587,N_7964);
and U11648 (N_11648,N_9827,N_9009);
xor U11649 (N_11649,N_9497,N_7620);
nor U11650 (N_11650,N_8820,N_8910);
and U11651 (N_11651,N_9239,N_8931);
nand U11652 (N_11652,N_9967,N_8423);
and U11653 (N_11653,N_7608,N_7994);
or U11654 (N_11654,N_8849,N_7624);
nor U11655 (N_11655,N_9567,N_9578);
nand U11656 (N_11656,N_9154,N_8473);
nand U11657 (N_11657,N_9825,N_8315);
or U11658 (N_11658,N_8131,N_8196);
nand U11659 (N_11659,N_8190,N_9894);
nand U11660 (N_11660,N_9455,N_8722);
nor U11661 (N_11661,N_7878,N_8410);
nand U11662 (N_11662,N_8840,N_8699);
nor U11663 (N_11663,N_9812,N_8960);
nor U11664 (N_11664,N_8244,N_8931);
or U11665 (N_11665,N_7823,N_9512);
and U11666 (N_11666,N_8529,N_9321);
or U11667 (N_11667,N_8229,N_9563);
nand U11668 (N_11668,N_9300,N_8407);
nor U11669 (N_11669,N_9791,N_8057);
nor U11670 (N_11670,N_8535,N_9195);
nand U11671 (N_11671,N_8792,N_7980);
and U11672 (N_11672,N_9952,N_8583);
and U11673 (N_11673,N_8931,N_9794);
or U11674 (N_11674,N_9559,N_8452);
nor U11675 (N_11675,N_7907,N_9168);
xor U11676 (N_11676,N_8869,N_7719);
or U11677 (N_11677,N_9644,N_9890);
and U11678 (N_11678,N_9284,N_8129);
and U11679 (N_11679,N_8560,N_8677);
and U11680 (N_11680,N_9385,N_8487);
and U11681 (N_11681,N_9507,N_8432);
and U11682 (N_11682,N_8476,N_9068);
or U11683 (N_11683,N_9005,N_7894);
nand U11684 (N_11684,N_9854,N_8101);
and U11685 (N_11685,N_9260,N_9807);
and U11686 (N_11686,N_8098,N_9476);
and U11687 (N_11687,N_7501,N_9627);
and U11688 (N_11688,N_8020,N_7881);
or U11689 (N_11689,N_7795,N_9984);
or U11690 (N_11690,N_8949,N_9535);
nand U11691 (N_11691,N_9171,N_7603);
and U11692 (N_11692,N_8237,N_9957);
xor U11693 (N_11693,N_8780,N_7528);
and U11694 (N_11694,N_9380,N_9922);
nor U11695 (N_11695,N_8801,N_9739);
nand U11696 (N_11696,N_8909,N_7643);
nand U11697 (N_11697,N_9813,N_9375);
nand U11698 (N_11698,N_8480,N_7648);
nor U11699 (N_11699,N_7559,N_9017);
and U11700 (N_11700,N_8771,N_8352);
nor U11701 (N_11701,N_7702,N_8390);
nand U11702 (N_11702,N_9002,N_8074);
and U11703 (N_11703,N_8631,N_9266);
and U11704 (N_11704,N_7865,N_9112);
nor U11705 (N_11705,N_8515,N_8362);
and U11706 (N_11706,N_9566,N_8464);
and U11707 (N_11707,N_9620,N_7525);
or U11708 (N_11708,N_8635,N_9101);
xnor U11709 (N_11709,N_9312,N_9061);
nor U11710 (N_11710,N_9755,N_7596);
and U11711 (N_11711,N_7660,N_8287);
or U11712 (N_11712,N_7868,N_7923);
nand U11713 (N_11713,N_8227,N_9715);
or U11714 (N_11714,N_8451,N_7509);
and U11715 (N_11715,N_8551,N_8599);
nor U11716 (N_11716,N_9335,N_9920);
nand U11717 (N_11717,N_9226,N_8784);
nor U11718 (N_11718,N_9150,N_9570);
nand U11719 (N_11719,N_8490,N_8079);
or U11720 (N_11720,N_8376,N_8857);
or U11721 (N_11721,N_7982,N_9982);
or U11722 (N_11722,N_7807,N_7842);
nand U11723 (N_11723,N_8065,N_9658);
or U11724 (N_11724,N_7925,N_7959);
and U11725 (N_11725,N_9771,N_9130);
nor U11726 (N_11726,N_9257,N_7511);
nand U11727 (N_11727,N_9467,N_9005);
nand U11728 (N_11728,N_8661,N_9964);
and U11729 (N_11729,N_8688,N_8566);
or U11730 (N_11730,N_8000,N_8077);
nor U11731 (N_11731,N_9470,N_8207);
or U11732 (N_11732,N_7836,N_9428);
nor U11733 (N_11733,N_9481,N_8022);
nand U11734 (N_11734,N_9951,N_9600);
and U11735 (N_11735,N_8379,N_8879);
nor U11736 (N_11736,N_9471,N_9265);
nor U11737 (N_11737,N_8664,N_9302);
nor U11738 (N_11738,N_7902,N_7813);
nor U11739 (N_11739,N_8796,N_9434);
or U11740 (N_11740,N_8784,N_8516);
and U11741 (N_11741,N_8452,N_8015);
or U11742 (N_11742,N_9429,N_8202);
and U11743 (N_11743,N_7855,N_8445);
nand U11744 (N_11744,N_9235,N_9857);
and U11745 (N_11745,N_9114,N_7959);
nand U11746 (N_11746,N_7557,N_9814);
or U11747 (N_11747,N_9745,N_7510);
nor U11748 (N_11748,N_9711,N_9143);
xnor U11749 (N_11749,N_9965,N_7817);
nor U11750 (N_11750,N_8669,N_7966);
and U11751 (N_11751,N_9653,N_8734);
and U11752 (N_11752,N_8052,N_9392);
nor U11753 (N_11753,N_9224,N_7973);
and U11754 (N_11754,N_9196,N_9002);
and U11755 (N_11755,N_9198,N_7724);
xor U11756 (N_11756,N_8899,N_9915);
and U11757 (N_11757,N_8118,N_8720);
nor U11758 (N_11758,N_9043,N_8847);
nor U11759 (N_11759,N_8913,N_7997);
nand U11760 (N_11760,N_8612,N_9309);
nor U11761 (N_11761,N_7820,N_7675);
or U11762 (N_11762,N_8688,N_8847);
and U11763 (N_11763,N_8373,N_8360);
nand U11764 (N_11764,N_7852,N_9217);
or U11765 (N_11765,N_9828,N_7518);
nor U11766 (N_11766,N_7968,N_9226);
or U11767 (N_11767,N_9751,N_8771);
and U11768 (N_11768,N_9339,N_8722);
or U11769 (N_11769,N_8242,N_9390);
and U11770 (N_11770,N_8918,N_7891);
nor U11771 (N_11771,N_8877,N_8728);
and U11772 (N_11772,N_9593,N_7668);
nor U11773 (N_11773,N_9730,N_8419);
and U11774 (N_11774,N_9108,N_9972);
or U11775 (N_11775,N_8573,N_8669);
and U11776 (N_11776,N_9420,N_7741);
nor U11777 (N_11777,N_8959,N_8788);
and U11778 (N_11778,N_7936,N_9293);
and U11779 (N_11779,N_7832,N_7836);
xor U11780 (N_11780,N_8717,N_8648);
nand U11781 (N_11781,N_8976,N_9532);
or U11782 (N_11782,N_8154,N_8562);
or U11783 (N_11783,N_9607,N_9151);
nand U11784 (N_11784,N_8841,N_9011);
and U11785 (N_11785,N_8655,N_8194);
or U11786 (N_11786,N_9175,N_8187);
and U11787 (N_11787,N_9939,N_8452);
and U11788 (N_11788,N_8755,N_9998);
and U11789 (N_11789,N_8141,N_8518);
nor U11790 (N_11790,N_9990,N_8615);
xor U11791 (N_11791,N_8255,N_8639);
or U11792 (N_11792,N_7699,N_9183);
nand U11793 (N_11793,N_9836,N_8742);
or U11794 (N_11794,N_7670,N_8378);
and U11795 (N_11795,N_8992,N_8936);
and U11796 (N_11796,N_8615,N_9717);
nor U11797 (N_11797,N_8666,N_7739);
and U11798 (N_11798,N_9435,N_8030);
nor U11799 (N_11799,N_9592,N_8132);
and U11800 (N_11800,N_9044,N_8790);
or U11801 (N_11801,N_9864,N_8180);
or U11802 (N_11802,N_8413,N_9406);
nor U11803 (N_11803,N_9466,N_7702);
and U11804 (N_11804,N_7690,N_8333);
xnor U11805 (N_11805,N_8433,N_9719);
nor U11806 (N_11806,N_9942,N_8294);
and U11807 (N_11807,N_7549,N_7901);
xor U11808 (N_11808,N_9057,N_7503);
or U11809 (N_11809,N_9310,N_8285);
and U11810 (N_11810,N_9532,N_8256);
nand U11811 (N_11811,N_9308,N_7996);
or U11812 (N_11812,N_8886,N_9226);
nor U11813 (N_11813,N_9175,N_7678);
or U11814 (N_11814,N_8474,N_8282);
nand U11815 (N_11815,N_7516,N_7720);
or U11816 (N_11816,N_9866,N_7859);
nand U11817 (N_11817,N_8694,N_7705);
xor U11818 (N_11818,N_9858,N_7537);
nor U11819 (N_11819,N_9552,N_8441);
and U11820 (N_11820,N_9540,N_9463);
nand U11821 (N_11821,N_7963,N_8479);
xor U11822 (N_11822,N_8086,N_8914);
nand U11823 (N_11823,N_8146,N_9592);
nor U11824 (N_11824,N_9432,N_7747);
nor U11825 (N_11825,N_8910,N_9026);
and U11826 (N_11826,N_9929,N_9281);
xnor U11827 (N_11827,N_7906,N_9319);
nor U11828 (N_11828,N_8261,N_9019);
and U11829 (N_11829,N_7708,N_7881);
or U11830 (N_11830,N_7723,N_8361);
xor U11831 (N_11831,N_7851,N_8197);
and U11832 (N_11832,N_7867,N_7688);
and U11833 (N_11833,N_7801,N_9937);
nor U11834 (N_11834,N_9299,N_8645);
or U11835 (N_11835,N_9791,N_7913);
nand U11836 (N_11836,N_8172,N_9999);
or U11837 (N_11837,N_9748,N_7941);
nor U11838 (N_11838,N_9039,N_7536);
nand U11839 (N_11839,N_8242,N_8523);
nor U11840 (N_11840,N_7947,N_7810);
nand U11841 (N_11841,N_8254,N_7613);
xor U11842 (N_11842,N_8838,N_9967);
nand U11843 (N_11843,N_7543,N_8708);
nor U11844 (N_11844,N_7727,N_8577);
or U11845 (N_11845,N_8366,N_8426);
and U11846 (N_11846,N_7998,N_9539);
and U11847 (N_11847,N_9063,N_8386);
or U11848 (N_11848,N_9473,N_9797);
or U11849 (N_11849,N_9704,N_8215);
nand U11850 (N_11850,N_9471,N_9886);
and U11851 (N_11851,N_9517,N_9148);
and U11852 (N_11852,N_9624,N_8436);
nand U11853 (N_11853,N_8579,N_8451);
nand U11854 (N_11854,N_7943,N_8553);
xnor U11855 (N_11855,N_8538,N_9543);
nor U11856 (N_11856,N_7680,N_8531);
nand U11857 (N_11857,N_7740,N_8011);
xor U11858 (N_11858,N_9831,N_8481);
and U11859 (N_11859,N_9695,N_7688);
and U11860 (N_11860,N_8782,N_8965);
or U11861 (N_11861,N_9702,N_9758);
or U11862 (N_11862,N_7941,N_7841);
and U11863 (N_11863,N_9949,N_9324);
nor U11864 (N_11864,N_9703,N_8916);
and U11865 (N_11865,N_8979,N_9781);
nand U11866 (N_11866,N_7629,N_9811);
nand U11867 (N_11867,N_9234,N_8850);
and U11868 (N_11868,N_9331,N_9756);
xnor U11869 (N_11869,N_7738,N_8704);
or U11870 (N_11870,N_8919,N_8890);
nor U11871 (N_11871,N_9961,N_8363);
and U11872 (N_11872,N_7534,N_8432);
xnor U11873 (N_11873,N_8497,N_7953);
xor U11874 (N_11874,N_8769,N_8378);
nor U11875 (N_11875,N_9378,N_9521);
nand U11876 (N_11876,N_8146,N_8785);
nor U11877 (N_11877,N_8878,N_8752);
nand U11878 (N_11878,N_9856,N_8466);
or U11879 (N_11879,N_8782,N_9763);
or U11880 (N_11880,N_9695,N_7544);
nand U11881 (N_11881,N_9635,N_8990);
nor U11882 (N_11882,N_9009,N_7700);
xor U11883 (N_11883,N_9601,N_8729);
xor U11884 (N_11884,N_8644,N_8567);
nor U11885 (N_11885,N_8685,N_9982);
or U11886 (N_11886,N_8174,N_9156);
nand U11887 (N_11887,N_8237,N_9642);
nor U11888 (N_11888,N_7865,N_9340);
nor U11889 (N_11889,N_8084,N_8407);
and U11890 (N_11890,N_8141,N_8221);
or U11891 (N_11891,N_8984,N_8347);
and U11892 (N_11892,N_9220,N_9961);
and U11893 (N_11893,N_8224,N_9502);
and U11894 (N_11894,N_8534,N_9222);
and U11895 (N_11895,N_8373,N_9345);
and U11896 (N_11896,N_7767,N_8148);
and U11897 (N_11897,N_8433,N_9132);
nand U11898 (N_11898,N_8809,N_7674);
nor U11899 (N_11899,N_8309,N_8996);
and U11900 (N_11900,N_9366,N_9304);
nand U11901 (N_11901,N_8705,N_7654);
or U11902 (N_11902,N_9544,N_8358);
nor U11903 (N_11903,N_9525,N_9821);
and U11904 (N_11904,N_9414,N_7988);
and U11905 (N_11905,N_8709,N_9085);
nor U11906 (N_11906,N_9632,N_8435);
nand U11907 (N_11907,N_9621,N_9708);
and U11908 (N_11908,N_8447,N_9435);
nor U11909 (N_11909,N_9667,N_8651);
and U11910 (N_11910,N_9755,N_7994);
xor U11911 (N_11911,N_9936,N_7554);
or U11912 (N_11912,N_9610,N_7586);
nand U11913 (N_11913,N_9194,N_9467);
and U11914 (N_11914,N_8922,N_8871);
nand U11915 (N_11915,N_9705,N_7764);
and U11916 (N_11916,N_7918,N_9740);
or U11917 (N_11917,N_9597,N_8654);
nor U11918 (N_11918,N_9373,N_9360);
or U11919 (N_11919,N_7634,N_7512);
and U11920 (N_11920,N_9999,N_9255);
nand U11921 (N_11921,N_7627,N_9251);
nand U11922 (N_11922,N_8920,N_8662);
nand U11923 (N_11923,N_9304,N_9066);
and U11924 (N_11924,N_9078,N_9383);
nor U11925 (N_11925,N_8470,N_8950);
nor U11926 (N_11926,N_9752,N_8786);
nor U11927 (N_11927,N_9595,N_8517);
and U11928 (N_11928,N_9438,N_8777);
nor U11929 (N_11929,N_9828,N_8456);
and U11930 (N_11930,N_8075,N_8444);
xnor U11931 (N_11931,N_7716,N_7637);
xor U11932 (N_11932,N_9887,N_7579);
or U11933 (N_11933,N_8167,N_7504);
nor U11934 (N_11934,N_8806,N_8071);
and U11935 (N_11935,N_8661,N_9429);
and U11936 (N_11936,N_9396,N_7520);
or U11937 (N_11937,N_9296,N_7918);
or U11938 (N_11938,N_9629,N_7715);
nor U11939 (N_11939,N_9774,N_8651);
and U11940 (N_11940,N_9146,N_9355);
xor U11941 (N_11941,N_8968,N_9621);
nand U11942 (N_11942,N_9895,N_9589);
nand U11943 (N_11943,N_9097,N_7551);
xnor U11944 (N_11944,N_7560,N_8853);
or U11945 (N_11945,N_9146,N_9606);
nor U11946 (N_11946,N_7532,N_9600);
and U11947 (N_11947,N_9840,N_9548);
xnor U11948 (N_11948,N_8389,N_7925);
and U11949 (N_11949,N_8988,N_8762);
nor U11950 (N_11950,N_8840,N_9450);
nor U11951 (N_11951,N_9965,N_7538);
nand U11952 (N_11952,N_7604,N_7683);
or U11953 (N_11953,N_7716,N_8570);
or U11954 (N_11954,N_9938,N_9990);
nor U11955 (N_11955,N_9145,N_8712);
nand U11956 (N_11956,N_7679,N_9302);
nand U11957 (N_11957,N_9395,N_8474);
xor U11958 (N_11958,N_8282,N_9555);
or U11959 (N_11959,N_8881,N_7669);
nor U11960 (N_11960,N_7936,N_9950);
or U11961 (N_11961,N_8381,N_9683);
nand U11962 (N_11962,N_7805,N_8983);
nand U11963 (N_11963,N_9139,N_9301);
nand U11964 (N_11964,N_8029,N_7934);
nand U11965 (N_11965,N_8610,N_8101);
xnor U11966 (N_11966,N_8944,N_8312);
nor U11967 (N_11967,N_9012,N_7767);
or U11968 (N_11968,N_8184,N_8567);
nor U11969 (N_11969,N_9898,N_9511);
and U11970 (N_11970,N_9361,N_9629);
or U11971 (N_11971,N_9992,N_9781);
nor U11972 (N_11972,N_9658,N_9422);
or U11973 (N_11973,N_9803,N_7651);
nor U11974 (N_11974,N_7594,N_8157);
nor U11975 (N_11975,N_7591,N_7631);
nor U11976 (N_11976,N_7677,N_7807);
and U11977 (N_11977,N_9420,N_7796);
nand U11978 (N_11978,N_8221,N_8085);
nand U11979 (N_11979,N_9236,N_9293);
and U11980 (N_11980,N_9990,N_9304);
xnor U11981 (N_11981,N_8823,N_8653);
xor U11982 (N_11982,N_7682,N_9010);
xor U11983 (N_11983,N_8960,N_9743);
or U11984 (N_11984,N_8870,N_7769);
or U11985 (N_11985,N_8487,N_8029);
or U11986 (N_11986,N_7883,N_8885);
nor U11987 (N_11987,N_8418,N_9037);
and U11988 (N_11988,N_9515,N_8902);
or U11989 (N_11989,N_8690,N_9128);
nor U11990 (N_11990,N_8396,N_7514);
or U11991 (N_11991,N_8683,N_8641);
xnor U11992 (N_11992,N_8451,N_9501);
xnor U11993 (N_11993,N_8200,N_8959);
xnor U11994 (N_11994,N_8406,N_7764);
or U11995 (N_11995,N_7712,N_8496);
nand U11996 (N_11996,N_8085,N_8669);
xnor U11997 (N_11997,N_9851,N_9060);
and U11998 (N_11998,N_7582,N_8917);
xnor U11999 (N_11999,N_8223,N_9336);
nand U12000 (N_12000,N_7539,N_9515);
or U12001 (N_12001,N_9770,N_9750);
or U12002 (N_12002,N_8205,N_9724);
nand U12003 (N_12003,N_8072,N_8489);
nor U12004 (N_12004,N_8745,N_8643);
nand U12005 (N_12005,N_9245,N_9683);
or U12006 (N_12006,N_8066,N_9834);
nand U12007 (N_12007,N_9694,N_8006);
or U12008 (N_12008,N_8055,N_9153);
or U12009 (N_12009,N_9360,N_9064);
nor U12010 (N_12010,N_7632,N_7665);
nand U12011 (N_12011,N_8711,N_8657);
nand U12012 (N_12012,N_8284,N_7724);
nand U12013 (N_12013,N_8565,N_8465);
and U12014 (N_12014,N_8534,N_8620);
and U12015 (N_12015,N_7750,N_7707);
and U12016 (N_12016,N_9413,N_8620);
and U12017 (N_12017,N_9984,N_8399);
or U12018 (N_12018,N_7574,N_9639);
or U12019 (N_12019,N_9244,N_8306);
nor U12020 (N_12020,N_9960,N_8651);
and U12021 (N_12021,N_8465,N_8817);
nor U12022 (N_12022,N_8769,N_8609);
nand U12023 (N_12023,N_8550,N_8207);
or U12024 (N_12024,N_9316,N_8163);
and U12025 (N_12025,N_9877,N_8336);
and U12026 (N_12026,N_7589,N_8284);
nor U12027 (N_12027,N_7977,N_8579);
nand U12028 (N_12028,N_8943,N_9713);
nor U12029 (N_12029,N_7606,N_7597);
nand U12030 (N_12030,N_9013,N_8285);
nor U12031 (N_12031,N_7866,N_8916);
xnor U12032 (N_12032,N_9945,N_9673);
and U12033 (N_12033,N_8828,N_8636);
and U12034 (N_12034,N_7834,N_8043);
or U12035 (N_12035,N_7713,N_9530);
nand U12036 (N_12036,N_7786,N_9440);
nand U12037 (N_12037,N_9744,N_8665);
nor U12038 (N_12038,N_8870,N_9797);
nor U12039 (N_12039,N_7998,N_8176);
nand U12040 (N_12040,N_9954,N_9856);
nor U12041 (N_12041,N_7560,N_7840);
xor U12042 (N_12042,N_8983,N_9560);
nor U12043 (N_12043,N_9634,N_7609);
nand U12044 (N_12044,N_8870,N_8546);
nand U12045 (N_12045,N_7797,N_8145);
or U12046 (N_12046,N_9735,N_8743);
and U12047 (N_12047,N_8177,N_8971);
or U12048 (N_12048,N_7726,N_9097);
nand U12049 (N_12049,N_7943,N_8885);
nand U12050 (N_12050,N_7584,N_9258);
nand U12051 (N_12051,N_7564,N_9290);
nand U12052 (N_12052,N_9044,N_8472);
and U12053 (N_12053,N_9524,N_9017);
nor U12054 (N_12054,N_9215,N_8399);
xnor U12055 (N_12055,N_9686,N_8931);
nand U12056 (N_12056,N_7842,N_8933);
nand U12057 (N_12057,N_9183,N_8698);
or U12058 (N_12058,N_9290,N_8078);
and U12059 (N_12059,N_8098,N_9064);
and U12060 (N_12060,N_9457,N_9911);
nor U12061 (N_12061,N_9154,N_8639);
or U12062 (N_12062,N_7629,N_7758);
or U12063 (N_12063,N_9905,N_7586);
or U12064 (N_12064,N_9745,N_7627);
xnor U12065 (N_12065,N_7914,N_8749);
nand U12066 (N_12066,N_8038,N_8238);
nor U12067 (N_12067,N_9300,N_7724);
and U12068 (N_12068,N_9503,N_8028);
nand U12069 (N_12069,N_9865,N_8950);
nor U12070 (N_12070,N_9773,N_8611);
nor U12071 (N_12071,N_8245,N_8222);
and U12072 (N_12072,N_7500,N_8596);
and U12073 (N_12073,N_7941,N_8914);
xnor U12074 (N_12074,N_8689,N_9929);
xnor U12075 (N_12075,N_9720,N_8017);
nand U12076 (N_12076,N_9846,N_7775);
xnor U12077 (N_12077,N_8687,N_8558);
or U12078 (N_12078,N_8580,N_9101);
nor U12079 (N_12079,N_8739,N_8897);
or U12080 (N_12080,N_9110,N_9665);
and U12081 (N_12081,N_7974,N_7879);
and U12082 (N_12082,N_8685,N_7564);
nor U12083 (N_12083,N_8451,N_9171);
and U12084 (N_12084,N_8161,N_7751);
nand U12085 (N_12085,N_8605,N_9324);
or U12086 (N_12086,N_9426,N_9439);
and U12087 (N_12087,N_8106,N_9562);
and U12088 (N_12088,N_8968,N_7943);
and U12089 (N_12089,N_9604,N_9905);
nor U12090 (N_12090,N_8528,N_8950);
or U12091 (N_12091,N_9321,N_9183);
or U12092 (N_12092,N_8138,N_9805);
or U12093 (N_12093,N_8105,N_7904);
nand U12094 (N_12094,N_9832,N_8511);
nor U12095 (N_12095,N_8666,N_9156);
nand U12096 (N_12096,N_9226,N_8781);
or U12097 (N_12097,N_8519,N_8533);
nand U12098 (N_12098,N_9320,N_9481);
nand U12099 (N_12099,N_9709,N_8435);
or U12100 (N_12100,N_8397,N_9556);
or U12101 (N_12101,N_8212,N_8552);
xnor U12102 (N_12102,N_9417,N_9672);
nor U12103 (N_12103,N_8879,N_8200);
xnor U12104 (N_12104,N_8610,N_9303);
nor U12105 (N_12105,N_9075,N_9521);
xnor U12106 (N_12106,N_7792,N_7517);
nor U12107 (N_12107,N_9284,N_7544);
or U12108 (N_12108,N_8790,N_7741);
xor U12109 (N_12109,N_8796,N_7772);
nor U12110 (N_12110,N_8790,N_7502);
or U12111 (N_12111,N_9422,N_7629);
xor U12112 (N_12112,N_8243,N_7506);
nand U12113 (N_12113,N_9011,N_7791);
nor U12114 (N_12114,N_9608,N_7681);
nor U12115 (N_12115,N_7957,N_8346);
nand U12116 (N_12116,N_9213,N_8059);
or U12117 (N_12117,N_9642,N_9109);
nand U12118 (N_12118,N_9121,N_9015);
xor U12119 (N_12119,N_7526,N_9589);
and U12120 (N_12120,N_9043,N_9046);
and U12121 (N_12121,N_7513,N_8925);
or U12122 (N_12122,N_8393,N_9432);
and U12123 (N_12123,N_8191,N_9188);
xor U12124 (N_12124,N_9789,N_9908);
nor U12125 (N_12125,N_9528,N_8293);
and U12126 (N_12126,N_8029,N_8771);
nor U12127 (N_12127,N_9475,N_8607);
nor U12128 (N_12128,N_8070,N_9469);
xor U12129 (N_12129,N_9748,N_7635);
nand U12130 (N_12130,N_9050,N_7603);
xnor U12131 (N_12131,N_9470,N_9154);
nand U12132 (N_12132,N_9000,N_9403);
nand U12133 (N_12133,N_7562,N_9442);
or U12134 (N_12134,N_9214,N_9920);
nand U12135 (N_12135,N_8835,N_9172);
and U12136 (N_12136,N_9294,N_9847);
nor U12137 (N_12137,N_8357,N_8258);
or U12138 (N_12138,N_8456,N_7549);
nor U12139 (N_12139,N_8489,N_7856);
nand U12140 (N_12140,N_8595,N_7540);
nand U12141 (N_12141,N_7550,N_9591);
nor U12142 (N_12142,N_8530,N_8483);
xnor U12143 (N_12143,N_9183,N_7581);
nor U12144 (N_12144,N_8897,N_8502);
or U12145 (N_12145,N_9429,N_8453);
xnor U12146 (N_12146,N_9935,N_8105);
nor U12147 (N_12147,N_7562,N_8310);
nor U12148 (N_12148,N_7961,N_8852);
or U12149 (N_12149,N_9626,N_8444);
and U12150 (N_12150,N_8390,N_9412);
and U12151 (N_12151,N_9134,N_9263);
and U12152 (N_12152,N_7797,N_8872);
and U12153 (N_12153,N_7911,N_9179);
or U12154 (N_12154,N_7701,N_9902);
nor U12155 (N_12155,N_8351,N_8152);
nor U12156 (N_12156,N_8179,N_8862);
nor U12157 (N_12157,N_9615,N_8047);
nand U12158 (N_12158,N_9466,N_7816);
nor U12159 (N_12159,N_9755,N_8087);
nor U12160 (N_12160,N_8626,N_9411);
or U12161 (N_12161,N_9722,N_8549);
xnor U12162 (N_12162,N_8226,N_8750);
xor U12163 (N_12163,N_9925,N_7575);
or U12164 (N_12164,N_9011,N_9291);
or U12165 (N_12165,N_7511,N_8368);
xnor U12166 (N_12166,N_8771,N_9366);
xnor U12167 (N_12167,N_8066,N_9090);
or U12168 (N_12168,N_9873,N_9664);
nor U12169 (N_12169,N_7886,N_8093);
nor U12170 (N_12170,N_9820,N_9802);
nor U12171 (N_12171,N_8821,N_8447);
nand U12172 (N_12172,N_9216,N_9692);
and U12173 (N_12173,N_9298,N_9047);
nand U12174 (N_12174,N_9027,N_8198);
xor U12175 (N_12175,N_9125,N_9158);
xor U12176 (N_12176,N_9868,N_9296);
xor U12177 (N_12177,N_7602,N_9908);
and U12178 (N_12178,N_9836,N_8866);
and U12179 (N_12179,N_7951,N_8578);
nand U12180 (N_12180,N_8893,N_8967);
nor U12181 (N_12181,N_8448,N_7757);
nand U12182 (N_12182,N_7650,N_9668);
or U12183 (N_12183,N_7916,N_9465);
nand U12184 (N_12184,N_7997,N_9783);
nor U12185 (N_12185,N_8737,N_8167);
or U12186 (N_12186,N_9211,N_8144);
or U12187 (N_12187,N_7641,N_7942);
nor U12188 (N_12188,N_7552,N_8236);
or U12189 (N_12189,N_9955,N_7792);
nor U12190 (N_12190,N_8995,N_9906);
nor U12191 (N_12191,N_7658,N_8419);
or U12192 (N_12192,N_9575,N_9846);
nand U12193 (N_12193,N_8401,N_9996);
nand U12194 (N_12194,N_7558,N_7921);
nand U12195 (N_12195,N_8429,N_8675);
nand U12196 (N_12196,N_7793,N_9663);
nor U12197 (N_12197,N_8658,N_9733);
or U12198 (N_12198,N_8144,N_8601);
and U12199 (N_12199,N_8511,N_8160);
or U12200 (N_12200,N_8688,N_8854);
xnor U12201 (N_12201,N_7582,N_8730);
and U12202 (N_12202,N_8757,N_9685);
or U12203 (N_12203,N_9341,N_8354);
nor U12204 (N_12204,N_7724,N_9651);
or U12205 (N_12205,N_8479,N_9010);
nor U12206 (N_12206,N_9875,N_9583);
or U12207 (N_12207,N_9612,N_8599);
or U12208 (N_12208,N_8829,N_8531);
nor U12209 (N_12209,N_8557,N_9576);
nor U12210 (N_12210,N_9343,N_9133);
nand U12211 (N_12211,N_8787,N_9507);
nor U12212 (N_12212,N_9024,N_8928);
nand U12213 (N_12213,N_8449,N_9049);
or U12214 (N_12214,N_9561,N_9355);
nand U12215 (N_12215,N_9653,N_8540);
nand U12216 (N_12216,N_7513,N_7996);
xor U12217 (N_12217,N_8621,N_8136);
or U12218 (N_12218,N_9758,N_8967);
nand U12219 (N_12219,N_8149,N_8707);
and U12220 (N_12220,N_9466,N_9331);
nand U12221 (N_12221,N_9421,N_9165);
and U12222 (N_12222,N_7683,N_8016);
nor U12223 (N_12223,N_8171,N_9540);
nor U12224 (N_12224,N_9580,N_7542);
nand U12225 (N_12225,N_8367,N_9376);
nand U12226 (N_12226,N_9703,N_8291);
nor U12227 (N_12227,N_7612,N_9619);
or U12228 (N_12228,N_9123,N_9589);
or U12229 (N_12229,N_7819,N_9015);
xor U12230 (N_12230,N_7610,N_7852);
xnor U12231 (N_12231,N_8851,N_8633);
xor U12232 (N_12232,N_7503,N_8286);
xor U12233 (N_12233,N_9474,N_9519);
nand U12234 (N_12234,N_8691,N_9809);
nor U12235 (N_12235,N_8858,N_9443);
or U12236 (N_12236,N_9537,N_9268);
and U12237 (N_12237,N_9635,N_8308);
xnor U12238 (N_12238,N_8110,N_9369);
nor U12239 (N_12239,N_7832,N_9605);
nand U12240 (N_12240,N_8038,N_9588);
and U12241 (N_12241,N_9698,N_7780);
nor U12242 (N_12242,N_9250,N_9539);
xnor U12243 (N_12243,N_7871,N_8476);
nand U12244 (N_12244,N_9247,N_8286);
nor U12245 (N_12245,N_9044,N_9070);
and U12246 (N_12246,N_9416,N_8211);
nor U12247 (N_12247,N_8753,N_9863);
and U12248 (N_12248,N_9384,N_8348);
nor U12249 (N_12249,N_7525,N_7891);
nand U12250 (N_12250,N_8425,N_9613);
and U12251 (N_12251,N_9634,N_8004);
or U12252 (N_12252,N_7651,N_9522);
nand U12253 (N_12253,N_9678,N_7564);
and U12254 (N_12254,N_8980,N_9709);
or U12255 (N_12255,N_9115,N_9634);
xnor U12256 (N_12256,N_8361,N_9346);
and U12257 (N_12257,N_8223,N_8492);
and U12258 (N_12258,N_8694,N_8641);
and U12259 (N_12259,N_7569,N_9831);
or U12260 (N_12260,N_8648,N_8331);
and U12261 (N_12261,N_9798,N_8744);
nor U12262 (N_12262,N_9548,N_9317);
and U12263 (N_12263,N_9687,N_7753);
or U12264 (N_12264,N_9157,N_8267);
or U12265 (N_12265,N_9437,N_9306);
or U12266 (N_12266,N_8653,N_7978);
nand U12267 (N_12267,N_9419,N_9088);
xor U12268 (N_12268,N_9526,N_9403);
nor U12269 (N_12269,N_8019,N_9407);
xnor U12270 (N_12270,N_8331,N_8635);
and U12271 (N_12271,N_9548,N_8688);
or U12272 (N_12272,N_7913,N_9293);
and U12273 (N_12273,N_7615,N_7509);
and U12274 (N_12274,N_7516,N_9480);
and U12275 (N_12275,N_9173,N_9375);
and U12276 (N_12276,N_8865,N_8638);
nor U12277 (N_12277,N_9763,N_8847);
and U12278 (N_12278,N_8610,N_8880);
or U12279 (N_12279,N_8953,N_9929);
nor U12280 (N_12280,N_7832,N_8987);
or U12281 (N_12281,N_9124,N_9007);
or U12282 (N_12282,N_9758,N_8771);
or U12283 (N_12283,N_8872,N_8156);
or U12284 (N_12284,N_8446,N_9827);
nand U12285 (N_12285,N_9876,N_8688);
and U12286 (N_12286,N_8455,N_7826);
or U12287 (N_12287,N_9277,N_8022);
or U12288 (N_12288,N_7580,N_8511);
nand U12289 (N_12289,N_7729,N_8500);
xor U12290 (N_12290,N_9185,N_9465);
and U12291 (N_12291,N_8039,N_7904);
and U12292 (N_12292,N_9584,N_9879);
or U12293 (N_12293,N_9814,N_9749);
and U12294 (N_12294,N_7744,N_8208);
xnor U12295 (N_12295,N_7748,N_8861);
nand U12296 (N_12296,N_8962,N_9044);
xor U12297 (N_12297,N_9755,N_9649);
xor U12298 (N_12298,N_9139,N_7605);
or U12299 (N_12299,N_9285,N_7630);
and U12300 (N_12300,N_7653,N_9905);
nand U12301 (N_12301,N_8752,N_9369);
and U12302 (N_12302,N_9708,N_9805);
and U12303 (N_12303,N_8920,N_8534);
or U12304 (N_12304,N_7906,N_9720);
or U12305 (N_12305,N_7905,N_9540);
nor U12306 (N_12306,N_8729,N_7970);
nand U12307 (N_12307,N_8110,N_9554);
or U12308 (N_12308,N_9085,N_9300);
and U12309 (N_12309,N_8045,N_9287);
nand U12310 (N_12310,N_7754,N_9914);
or U12311 (N_12311,N_9015,N_9043);
nand U12312 (N_12312,N_9464,N_8875);
xor U12313 (N_12313,N_9140,N_8580);
nor U12314 (N_12314,N_8407,N_9087);
xnor U12315 (N_12315,N_9548,N_7991);
nor U12316 (N_12316,N_9659,N_8604);
or U12317 (N_12317,N_9948,N_9770);
or U12318 (N_12318,N_7539,N_9397);
nor U12319 (N_12319,N_7748,N_8834);
nor U12320 (N_12320,N_9296,N_9314);
and U12321 (N_12321,N_9539,N_9809);
xnor U12322 (N_12322,N_8234,N_8166);
nor U12323 (N_12323,N_8110,N_8858);
and U12324 (N_12324,N_9099,N_9614);
nand U12325 (N_12325,N_8886,N_8114);
xnor U12326 (N_12326,N_7963,N_8130);
or U12327 (N_12327,N_9149,N_8674);
nand U12328 (N_12328,N_9449,N_9838);
nand U12329 (N_12329,N_9339,N_8519);
nor U12330 (N_12330,N_9619,N_8505);
nand U12331 (N_12331,N_9104,N_9979);
and U12332 (N_12332,N_8679,N_9290);
nand U12333 (N_12333,N_8372,N_8039);
nor U12334 (N_12334,N_8412,N_7874);
nand U12335 (N_12335,N_8053,N_9908);
nor U12336 (N_12336,N_9939,N_9920);
nand U12337 (N_12337,N_8096,N_8862);
or U12338 (N_12338,N_8263,N_8750);
and U12339 (N_12339,N_8876,N_8250);
and U12340 (N_12340,N_8465,N_8154);
and U12341 (N_12341,N_8196,N_9839);
or U12342 (N_12342,N_9210,N_9348);
nor U12343 (N_12343,N_8535,N_9767);
nor U12344 (N_12344,N_8876,N_7596);
nand U12345 (N_12345,N_8494,N_7795);
or U12346 (N_12346,N_9045,N_8985);
and U12347 (N_12347,N_9016,N_8140);
nor U12348 (N_12348,N_9711,N_9372);
nand U12349 (N_12349,N_9549,N_9931);
nor U12350 (N_12350,N_9483,N_8215);
and U12351 (N_12351,N_8289,N_7917);
nand U12352 (N_12352,N_9617,N_9810);
or U12353 (N_12353,N_7871,N_8514);
and U12354 (N_12354,N_9584,N_9790);
and U12355 (N_12355,N_8195,N_9055);
or U12356 (N_12356,N_7933,N_9303);
and U12357 (N_12357,N_8885,N_8031);
and U12358 (N_12358,N_9175,N_9331);
and U12359 (N_12359,N_7990,N_7635);
nand U12360 (N_12360,N_9926,N_8276);
or U12361 (N_12361,N_7864,N_9784);
and U12362 (N_12362,N_9590,N_8667);
nor U12363 (N_12363,N_9483,N_8935);
nor U12364 (N_12364,N_8005,N_9835);
or U12365 (N_12365,N_8487,N_9517);
nand U12366 (N_12366,N_9607,N_9592);
nand U12367 (N_12367,N_7747,N_8917);
nand U12368 (N_12368,N_8227,N_8087);
nand U12369 (N_12369,N_8622,N_8965);
nor U12370 (N_12370,N_9142,N_7576);
and U12371 (N_12371,N_8095,N_8876);
and U12372 (N_12372,N_9299,N_9918);
or U12373 (N_12373,N_9540,N_7613);
nor U12374 (N_12374,N_8948,N_8691);
nor U12375 (N_12375,N_9878,N_8576);
nor U12376 (N_12376,N_7834,N_9385);
nand U12377 (N_12377,N_8314,N_8481);
and U12378 (N_12378,N_8219,N_7549);
nand U12379 (N_12379,N_8154,N_8188);
nand U12380 (N_12380,N_8631,N_9980);
or U12381 (N_12381,N_7603,N_7743);
nand U12382 (N_12382,N_8605,N_9870);
nand U12383 (N_12383,N_9782,N_8855);
nand U12384 (N_12384,N_8038,N_8919);
nand U12385 (N_12385,N_7694,N_9174);
and U12386 (N_12386,N_9603,N_9111);
nand U12387 (N_12387,N_7761,N_8238);
and U12388 (N_12388,N_9628,N_8200);
or U12389 (N_12389,N_8319,N_9556);
and U12390 (N_12390,N_9543,N_9753);
xnor U12391 (N_12391,N_8710,N_8480);
or U12392 (N_12392,N_8848,N_8067);
nor U12393 (N_12393,N_9701,N_9007);
nor U12394 (N_12394,N_7836,N_8957);
and U12395 (N_12395,N_8176,N_8525);
or U12396 (N_12396,N_9051,N_8907);
and U12397 (N_12397,N_9203,N_8695);
nor U12398 (N_12398,N_8783,N_8787);
nand U12399 (N_12399,N_9043,N_8806);
and U12400 (N_12400,N_9689,N_8414);
nand U12401 (N_12401,N_7924,N_9422);
and U12402 (N_12402,N_7551,N_8970);
and U12403 (N_12403,N_9112,N_7505);
and U12404 (N_12404,N_9554,N_7959);
nand U12405 (N_12405,N_9610,N_8796);
or U12406 (N_12406,N_7949,N_8567);
or U12407 (N_12407,N_8258,N_9822);
nand U12408 (N_12408,N_8866,N_8265);
or U12409 (N_12409,N_8279,N_9575);
xnor U12410 (N_12410,N_8756,N_7505);
nor U12411 (N_12411,N_9829,N_7953);
xnor U12412 (N_12412,N_9870,N_9041);
or U12413 (N_12413,N_8514,N_9316);
nor U12414 (N_12414,N_8947,N_8870);
nand U12415 (N_12415,N_7696,N_9904);
nor U12416 (N_12416,N_8834,N_9295);
nor U12417 (N_12417,N_8686,N_9553);
nor U12418 (N_12418,N_8030,N_7810);
and U12419 (N_12419,N_8498,N_8169);
nand U12420 (N_12420,N_7709,N_8318);
or U12421 (N_12421,N_8249,N_7719);
xnor U12422 (N_12422,N_8920,N_8539);
nor U12423 (N_12423,N_8784,N_9504);
and U12424 (N_12424,N_8982,N_9005);
nor U12425 (N_12425,N_8843,N_8493);
or U12426 (N_12426,N_8174,N_7977);
and U12427 (N_12427,N_9881,N_9293);
nor U12428 (N_12428,N_9164,N_9913);
or U12429 (N_12429,N_7872,N_9617);
nand U12430 (N_12430,N_9713,N_8270);
or U12431 (N_12431,N_9660,N_9804);
or U12432 (N_12432,N_9477,N_7912);
nand U12433 (N_12433,N_9767,N_8554);
and U12434 (N_12434,N_9011,N_9196);
nand U12435 (N_12435,N_7748,N_7647);
or U12436 (N_12436,N_7993,N_9118);
xor U12437 (N_12437,N_9571,N_9601);
nor U12438 (N_12438,N_7888,N_9711);
nor U12439 (N_12439,N_7761,N_8873);
or U12440 (N_12440,N_7809,N_8110);
or U12441 (N_12441,N_7624,N_8824);
nand U12442 (N_12442,N_7945,N_8634);
nand U12443 (N_12443,N_9867,N_8816);
or U12444 (N_12444,N_9340,N_8140);
xor U12445 (N_12445,N_9530,N_9989);
or U12446 (N_12446,N_9646,N_7682);
and U12447 (N_12447,N_8104,N_7765);
nand U12448 (N_12448,N_8089,N_9228);
or U12449 (N_12449,N_7524,N_8114);
nor U12450 (N_12450,N_8704,N_8915);
nand U12451 (N_12451,N_9488,N_8186);
nor U12452 (N_12452,N_9478,N_8443);
or U12453 (N_12453,N_9062,N_8319);
nor U12454 (N_12454,N_9225,N_7792);
and U12455 (N_12455,N_8686,N_8819);
nand U12456 (N_12456,N_9604,N_8099);
and U12457 (N_12457,N_9449,N_8738);
and U12458 (N_12458,N_7921,N_7976);
or U12459 (N_12459,N_8566,N_9494);
nand U12460 (N_12460,N_9379,N_8579);
and U12461 (N_12461,N_8804,N_7953);
nand U12462 (N_12462,N_9929,N_9090);
nor U12463 (N_12463,N_8452,N_7946);
or U12464 (N_12464,N_9470,N_9852);
nand U12465 (N_12465,N_9414,N_8812);
nand U12466 (N_12466,N_9892,N_9256);
or U12467 (N_12467,N_8857,N_9034);
or U12468 (N_12468,N_8547,N_9334);
nand U12469 (N_12469,N_9269,N_8115);
nor U12470 (N_12470,N_7718,N_7807);
and U12471 (N_12471,N_9457,N_8888);
and U12472 (N_12472,N_9223,N_7745);
nand U12473 (N_12473,N_9377,N_8328);
xnor U12474 (N_12474,N_9994,N_9062);
or U12475 (N_12475,N_7730,N_9707);
nor U12476 (N_12476,N_8194,N_8363);
nor U12477 (N_12477,N_8828,N_9659);
nand U12478 (N_12478,N_7830,N_9562);
or U12479 (N_12479,N_9130,N_7695);
nand U12480 (N_12480,N_9745,N_8180);
nor U12481 (N_12481,N_8055,N_8729);
xnor U12482 (N_12482,N_7903,N_9641);
or U12483 (N_12483,N_9244,N_9789);
or U12484 (N_12484,N_8678,N_9285);
and U12485 (N_12485,N_9096,N_7970);
nand U12486 (N_12486,N_9196,N_7751);
nand U12487 (N_12487,N_8310,N_8189);
xor U12488 (N_12488,N_9972,N_7840);
and U12489 (N_12489,N_9637,N_9140);
nor U12490 (N_12490,N_9420,N_9533);
nand U12491 (N_12491,N_7811,N_7944);
nor U12492 (N_12492,N_7972,N_9834);
nand U12493 (N_12493,N_8070,N_8169);
and U12494 (N_12494,N_8188,N_8521);
or U12495 (N_12495,N_9046,N_9128);
xnor U12496 (N_12496,N_7668,N_8469);
nand U12497 (N_12497,N_7520,N_9198);
and U12498 (N_12498,N_8364,N_8860);
and U12499 (N_12499,N_8179,N_7643);
and U12500 (N_12500,N_11989,N_10853);
nand U12501 (N_12501,N_10357,N_11058);
or U12502 (N_12502,N_12420,N_11637);
or U12503 (N_12503,N_10280,N_10966);
and U12504 (N_12504,N_10737,N_12066);
nor U12505 (N_12505,N_12361,N_10332);
or U12506 (N_12506,N_11268,N_10151);
xor U12507 (N_12507,N_12118,N_12431);
nand U12508 (N_12508,N_10697,N_10906);
nor U12509 (N_12509,N_12327,N_12235);
and U12510 (N_12510,N_11606,N_11972);
nand U12511 (N_12511,N_11082,N_10176);
nand U12512 (N_12512,N_11091,N_10169);
or U12513 (N_12513,N_10682,N_10041);
nand U12514 (N_12514,N_10857,N_11676);
nand U12515 (N_12515,N_10081,N_10931);
nor U12516 (N_12516,N_12297,N_10091);
nor U12517 (N_12517,N_11025,N_11877);
nor U12518 (N_12518,N_10377,N_11469);
nand U12519 (N_12519,N_10586,N_11516);
nor U12520 (N_12520,N_10662,N_11296);
or U12521 (N_12521,N_12243,N_11643);
nand U12522 (N_12522,N_11067,N_10406);
and U12523 (N_12523,N_11856,N_12165);
nand U12524 (N_12524,N_11874,N_12425);
xnor U12525 (N_12525,N_12147,N_11880);
or U12526 (N_12526,N_10202,N_12496);
nand U12527 (N_12527,N_11159,N_10884);
and U12528 (N_12528,N_10367,N_10088);
nor U12529 (N_12529,N_11299,N_10923);
nor U12530 (N_12530,N_10944,N_11841);
nor U12531 (N_12531,N_11817,N_11656);
nor U12532 (N_12532,N_11133,N_11172);
and U12533 (N_12533,N_10901,N_11384);
nand U12534 (N_12534,N_11364,N_11899);
and U12535 (N_12535,N_10532,N_11881);
xor U12536 (N_12536,N_10218,N_12416);
nor U12537 (N_12537,N_10313,N_11706);
or U12538 (N_12538,N_10842,N_12368);
or U12539 (N_12539,N_11087,N_10032);
nand U12540 (N_12540,N_11106,N_11331);
or U12541 (N_12541,N_10397,N_10368);
nor U12542 (N_12542,N_11430,N_10914);
or U12543 (N_12543,N_12444,N_10413);
xor U12544 (N_12544,N_12291,N_10083);
or U12545 (N_12545,N_10993,N_10732);
or U12546 (N_12546,N_11807,N_10131);
nor U12547 (N_12547,N_11935,N_11465);
xor U12548 (N_12548,N_11089,N_11586);
xnor U12549 (N_12549,N_10744,N_10150);
nand U12550 (N_12550,N_10433,N_11502);
nand U12551 (N_12551,N_11815,N_11065);
nor U12552 (N_12552,N_11314,N_11996);
nor U12553 (N_12553,N_11302,N_10781);
nand U12554 (N_12554,N_10025,N_11205);
and U12555 (N_12555,N_11851,N_10861);
nand U12556 (N_12556,N_11327,N_11351);
xor U12557 (N_12557,N_11278,N_11190);
nand U12558 (N_12558,N_11990,N_10859);
or U12559 (N_12559,N_11372,N_10269);
xnor U12560 (N_12560,N_11128,N_10801);
nor U12561 (N_12561,N_10386,N_11948);
xnor U12562 (N_12562,N_10001,N_11201);
nand U12563 (N_12563,N_12175,N_12299);
or U12564 (N_12564,N_10704,N_11934);
nand U12565 (N_12565,N_11052,N_11869);
or U12566 (N_12566,N_11657,N_10190);
nand U12567 (N_12567,N_11322,N_11170);
and U12568 (N_12568,N_12041,N_10359);
nand U12569 (N_12569,N_11311,N_10265);
or U12570 (N_12570,N_11005,N_11902);
xnor U12571 (N_12571,N_10608,N_11235);
nand U12572 (N_12572,N_10547,N_12447);
nand U12573 (N_12573,N_11876,N_11720);
nand U12574 (N_12574,N_12206,N_10317);
nor U12575 (N_12575,N_10450,N_10974);
nand U12576 (N_12576,N_10896,N_10680);
or U12577 (N_12577,N_10266,N_12240);
xnor U12578 (N_12578,N_10749,N_10309);
and U12579 (N_12579,N_11439,N_10205);
or U12580 (N_12580,N_11511,N_11672);
nand U12581 (N_12581,N_10883,N_12126);
nand U12582 (N_12582,N_11432,N_12064);
nor U12583 (N_12583,N_11885,N_11111);
xor U12584 (N_12584,N_12346,N_10183);
nor U12585 (N_12585,N_12472,N_11028);
or U12586 (N_12586,N_11486,N_11472);
or U12587 (N_12587,N_10271,N_11580);
or U12588 (N_12588,N_10063,N_11335);
nand U12589 (N_12589,N_12079,N_11233);
nand U12590 (N_12590,N_12424,N_11552);
and U12591 (N_12591,N_11821,N_10870);
xnor U12592 (N_12592,N_10015,N_12104);
nor U12593 (N_12593,N_11218,N_12109);
and U12594 (N_12594,N_11797,N_12320);
or U12595 (N_12595,N_10724,N_10513);
and U12596 (N_12596,N_12469,N_12199);
and U12597 (N_12597,N_12323,N_12253);
or U12598 (N_12598,N_10132,N_11558);
nor U12599 (N_12599,N_10037,N_11733);
and U12600 (N_12600,N_12061,N_10741);
nand U12601 (N_12601,N_12497,N_12358);
nor U12602 (N_12602,N_10172,N_10438);
nand U12603 (N_12603,N_12234,N_10486);
nor U12604 (N_12604,N_11875,N_10130);
xnor U12605 (N_12605,N_10773,N_11269);
nand U12606 (N_12606,N_10338,N_10283);
or U12607 (N_12607,N_11452,N_10666);
nor U12608 (N_12608,N_11811,N_12399);
xor U12609 (N_12609,N_12308,N_11464);
and U12610 (N_12610,N_12107,N_11313);
and U12611 (N_12611,N_12459,N_11217);
xnor U12612 (N_12612,N_10849,N_11346);
nand U12613 (N_12613,N_12316,N_11491);
xor U12614 (N_12614,N_11015,N_12488);
nor U12615 (N_12615,N_11588,N_11993);
nor U12616 (N_12616,N_10412,N_12266);
nand U12617 (N_12617,N_11461,N_12355);
xnor U12618 (N_12618,N_11768,N_11496);
nor U12619 (N_12619,N_10559,N_11199);
nand U12620 (N_12620,N_10108,N_10659);
or U12621 (N_12621,N_12169,N_11510);
nor U12622 (N_12622,N_11569,N_11009);
and U12623 (N_12623,N_10067,N_11288);
and U12624 (N_12624,N_12189,N_10587);
nor U12625 (N_12625,N_10573,N_10620);
and U12626 (N_12626,N_12385,N_10237);
nand U12627 (N_12627,N_11281,N_11828);
and U12628 (N_12628,N_10527,N_10447);
nor U12629 (N_12629,N_10153,N_10622);
nand U12630 (N_12630,N_10679,N_11363);
nor U12631 (N_12631,N_10575,N_10181);
nor U12632 (N_12632,N_11029,N_10435);
or U12633 (N_12633,N_12010,N_10648);
nor U12634 (N_12634,N_11203,N_10495);
nand U12635 (N_12635,N_11919,N_10717);
nand U12636 (N_12636,N_11515,N_12337);
and U12637 (N_12637,N_12057,N_10196);
nor U12638 (N_12638,N_10654,N_12367);
nand U12639 (N_12639,N_12384,N_11225);
or U12640 (N_12640,N_12335,N_11227);
nor U12641 (N_12641,N_10248,N_11774);
nor U12642 (N_12642,N_10674,N_10752);
and U12643 (N_12643,N_10696,N_12436);
and U12644 (N_12644,N_11147,N_10427);
xnor U12645 (N_12645,N_11859,N_11303);
or U12646 (N_12646,N_10734,N_10841);
nand U12647 (N_12647,N_12054,N_12260);
and U12648 (N_12648,N_10018,N_10369);
nand U12649 (N_12649,N_11531,N_11783);
nor U12650 (N_12650,N_12003,N_10467);
and U12651 (N_12651,N_11011,N_12482);
nor U12652 (N_12652,N_11426,N_11553);
nor U12653 (N_12653,N_10492,N_11534);
and U12654 (N_12654,N_12491,N_12035);
nand U12655 (N_12655,N_12303,N_12124);
xnor U12656 (N_12656,N_11727,N_11631);
and U12657 (N_12657,N_11548,N_12056);
or U12658 (N_12658,N_12078,N_10158);
nand U12659 (N_12659,N_10574,N_10556);
xor U12660 (N_12660,N_11286,N_11295);
nand U12661 (N_12661,N_10557,N_10077);
or U12662 (N_12662,N_10410,N_11107);
nor U12663 (N_12663,N_12471,N_10156);
nor U12664 (N_12664,N_12418,N_10723);
or U12665 (N_12665,N_11766,N_10405);
and U12666 (N_12666,N_11812,N_12004);
or U12667 (N_12667,N_10913,N_12142);
nand U12668 (N_12668,N_12307,N_11800);
and U12669 (N_12669,N_10321,N_10824);
or U12670 (N_12670,N_11057,N_10881);
nand U12671 (N_12671,N_10889,N_12429);
xor U12672 (N_12672,N_12073,N_11060);
or U12673 (N_12673,N_12071,N_10634);
nand U12674 (N_12674,N_10805,N_12152);
or U12675 (N_12675,N_10470,N_10258);
and U12676 (N_12676,N_11238,N_10508);
or U12677 (N_12677,N_10845,N_10710);
and U12678 (N_12678,N_11010,N_11930);
nor U12679 (N_12679,N_10910,N_10291);
nand U12680 (N_12680,N_10817,N_11032);
or U12681 (N_12681,N_10670,N_11559);
xnor U12682 (N_12682,N_11158,N_10459);
or U12683 (N_12683,N_11273,N_11002);
and U12684 (N_12684,N_11256,N_12298);
and U12685 (N_12685,N_11370,N_12406);
nor U12686 (N_12686,N_10808,N_10693);
or U12687 (N_12687,N_11577,N_11751);
and U12688 (N_12688,N_11801,N_10558);
and U12689 (N_12689,N_12435,N_11382);
xor U12690 (N_12690,N_11261,N_10758);
and U12691 (N_12691,N_12033,N_10024);
nor U12692 (N_12692,N_10136,N_10102);
nand U12693 (N_12693,N_11879,N_10942);
nand U12694 (N_12694,N_11603,N_10929);
nand U12695 (N_12695,N_11762,N_12250);
and U12696 (N_12696,N_12373,N_10355);
nor U12697 (N_12697,N_12221,N_10580);
or U12698 (N_12698,N_10312,N_10086);
and U12699 (N_12699,N_10457,N_10612);
nand U12700 (N_12700,N_12392,N_10822);
nor U12701 (N_12701,N_10113,N_10366);
nand U12702 (N_12702,N_11663,N_11118);
nor U12703 (N_12703,N_10154,N_10166);
nor U12704 (N_12704,N_11674,N_10968);
and U12705 (N_12705,N_11664,N_10227);
or U12706 (N_12706,N_10058,N_11914);
and U12707 (N_12707,N_10485,N_11964);
and U12708 (N_12708,N_11143,N_11232);
and U12709 (N_12709,N_12315,N_10745);
or U12710 (N_12710,N_12467,N_11799);
or U12711 (N_12711,N_11419,N_12014);
and U12712 (N_12712,N_10493,N_10468);
and U12713 (N_12713,N_11734,N_12100);
nand U12714 (N_12714,N_11488,N_10123);
nor U12715 (N_12715,N_11916,N_10542);
nand U12716 (N_12716,N_12473,N_11520);
nor U12717 (N_12717,N_11629,N_12359);
and U12718 (N_12718,N_10767,N_11323);
nor U12719 (N_12719,N_10033,N_12087);
nor U12720 (N_12720,N_10323,N_11283);
xnor U12721 (N_12721,N_12188,N_10727);
xor U12722 (N_12722,N_11195,N_10263);
and U12723 (N_12723,N_10792,N_11215);
nand U12724 (N_12724,N_11245,N_12131);
or U12725 (N_12725,N_11350,N_11478);
and U12726 (N_12726,N_10617,N_10992);
or U12727 (N_12727,N_11064,N_12149);
or U12728 (N_12728,N_12486,N_10152);
nor U12729 (N_12729,N_11229,N_10221);
or U12730 (N_12730,N_10610,N_10898);
nor U12731 (N_12731,N_10217,N_10628);
or U12732 (N_12732,N_10353,N_11100);
xor U12733 (N_12733,N_12099,N_12351);
and U12734 (N_12734,N_10199,N_11844);
nand U12735 (N_12735,N_11099,N_12452);
nand U12736 (N_12736,N_12246,N_10403);
and U12737 (N_12737,N_12249,N_10192);
and U12738 (N_12738,N_11981,N_12463);
nor U12739 (N_12739,N_11682,N_11980);
nor U12740 (N_12740,N_10897,N_12415);
nor U12741 (N_12741,N_10769,N_12094);
and U12742 (N_12742,N_10633,N_10442);
nand U12743 (N_12743,N_10489,N_11700);
and U12744 (N_12744,N_11458,N_11627);
nor U12745 (N_12745,N_11825,N_10615);
and U12746 (N_12746,N_11389,N_10932);
and U12747 (N_12747,N_11449,N_11022);
nand U12748 (N_12748,N_11598,N_10938);
or U12749 (N_12749,N_11354,N_11713);
and U12750 (N_12750,N_10160,N_11416);
nand U12751 (N_12751,N_12423,N_12024);
and U12752 (N_12752,N_10415,N_11001);
or U12753 (N_12753,N_10950,N_11396);
nand U12754 (N_12754,N_10969,N_10996);
and U12755 (N_12755,N_11081,N_10719);
or U12756 (N_12756,N_10478,N_10943);
nand U12757 (N_12757,N_10834,N_10742);
or U12758 (N_12758,N_12440,N_10625);
nor U12759 (N_12759,N_11780,N_11388);
nand U12760 (N_12760,N_12052,N_12151);
nor U12761 (N_12761,N_11505,N_10385);
or U12762 (N_12762,N_10224,N_10706);
or U12763 (N_12763,N_10678,N_10303);
nor U12764 (N_12764,N_10296,N_10106);
nand U12765 (N_12765,N_10677,N_11581);
nand U12766 (N_12766,N_12322,N_12158);
nor U12767 (N_12767,N_10319,N_10751);
nor U12768 (N_12768,N_11892,N_10148);
or U12769 (N_12769,N_11884,N_12215);
xor U12770 (N_12770,N_10311,N_12095);
and U12771 (N_12771,N_10909,N_11526);
xnor U12772 (N_12772,N_11633,N_11114);
nand U12773 (N_12773,N_11392,N_10429);
xor U12774 (N_12774,N_12251,N_10827);
nand U12775 (N_12775,N_12047,N_10970);
nand U12776 (N_12776,N_10236,N_10243);
nand U12777 (N_12777,N_11110,N_11873);
nand U12778 (N_12778,N_11787,N_11379);
xor U12779 (N_12779,N_10596,N_10920);
nor U12780 (N_12780,N_10491,N_10935);
nor U12781 (N_12781,N_11101,N_11518);
or U12782 (N_12782,N_10066,N_10515);
xor U12783 (N_12783,N_11315,N_10206);
and U12784 (N_12784,N_10093,N_12461);
and U12785 (N_12785,N_12101,N_11312);
and U12786 (N_12786,N_10268,N_11513);
nand U12787 (N_12787,N_11810,N_10120);
or U12788 (N_12788,N_12049,N_10940);
nand U12789 (N_12789,N_12313,N_12224);
and U12790 (N_12790,N_11166,N_10304);
nand U12791 (N_12791,N_10541,N_12374);
xor U12792 (N_12792,N_12258,N_11152);
nand U12793 (N_12793,N_11375,N_11122);
nand U12794 (N_12794,N_11231,N_10637);
xnor U12795 (N_12795,N_10585,N_10843);
nor U12796 (N_12796,N_11670,N_11503);
or U12797 (N_12797,N_11560,N_11198);
or U12798 (N_12798,N_11541,N_11482);
and U12799 (N_12799,N_11297,N_10064);
xor U12800 (N_12800,N_10655,N_11043);
nand U12801 (N_12801,N_12160,N_11251);
or U12802 (N_12802,N_12289,N_10975);
nand U12803 (N_12803,N_11417,N_12086);
xor U12804 (N_12804,N_11320,N_11454);
nand U12805 (N_12805,N_10245,N_12362);
nand U12806 (N_12806,N_10535,N_10246);
nand U12807 (N_12807,N_11747,N_11954);
and U12808 (N_12808,N_12190,N_12178);
xor U12809 (N_12809,N_10971,N_10840);
nand U12810 (N_12810,N_11903,N_11535);
nand U12811 (N_12811,N_10770,N_11249);
or U12812 (N_12812,N_10418,N_10978);
or U12813 (N_12813,N_12377,N_12139);
xor U12814 (N_12814,N_12204,N_12364);
or U12815 (N_12815,N_12287,N_12120);
nor U12816 (N_12816,N_10480,N_12470);
nor U12817 (N_12817,N_10097,N_12348);
or U12818 (N_12818,N_11255,N_11895);
and U12819 (N_12819,N_12405,N_10301);
nand U12820 (N_12820,N_10600,N_10383);
xor U12821 (N_12821,N_10220,N_12051);
or U12822 (N_12822,N_11489,N_10354);
nor U12823 (N_12823,N_10345,N_11070);
or U12824 (N_12824,N_10168,N_10287);
or U12825 (N_12825,N_10004,N_12237);
nand U12826 (N_12826,N_10384,N_11784);
nor U12827 (N_12827,N_12172,N_11196);
and U12828 (N_12828,N_11786,N_12219);
xor U12829 (N_12829,N_10563,N_11007);
nor U12830 (N_12830,N_10420,N_11049);
nor U12831 (N_12831,N_10340,N_10533);
and U12832 (N_12832,N_10228,N_12218);
or U12833 (N_12833,N_12474,N_10238);
nand U12834 (N_12834,N_10143,N_11130);
nor U12835 (N_12835,N_11492,N_10635);
or U12836 (N_12836,N_11102,N_11938);
or U12837 (N_12837,N_12422,N_12026);
and U12838 (N_12838,N_10663,N_12343);
and U12839 (N_12839,N_11069,N_11969);
or U12840 (N_12840,N_12228,N_10979);
nand U12841 (N_12841,N_11076,N_11846);
nand U12842 (N_12842,N_11153,N_10488);
nand U12843 (N_12843,N_11694,N_11487);
nor U12844 (N_12844,N_11123,N_11855);
or U12845 (N_12845,N_11186,N_10255);
nand U12846 (N_12846,N_12257,N_12354);
nand U12847 (N_12847,N_12011,N_11715);
nor U12848 (N_12848,N_10646,N_10144);
and U12849 (N_12849,N_11355,N_10708);
nand U12850 (N_12850,N_10084,N_11023);
nor U12851 (N_12851,N_11726,N_10440);
or U12852 (N_12852,N_10203,N_11500);
nand U12853 (N_12853,N_11391,N_12338);
nor U12854 (N_12854,N_11613,N_12113);
and U12855 (N_12855,N_10096,N_10484);
or U12856 (N_12856,N_11748,N_11723);
or U12857 (N_12857,N_10525,N_11517);
nand U12858 (N_12858,N_10242,N_10430);
or U12859 (N_12859,N_10452,N_11642);
nand U12860 (N_12860,N_11839,N_11804);
and U12861 (N_12861,N_10788,N_11362);
nand U12862 (N_12862,N_10416,N_10510);
nand U12863 (N_12863,N_12283,N_12388);
nand U12864 (N_12864,N_10284,N_10964);
nand U12865 (N_12865,N_10721,N_11330);
and U12866 (N_12866,N_12311,N_10239);
and U12867 (N_12867,N_12458,N_10134);
and U12868 (N_12868,N_11253,N_10581);
and U12869 (N_12869,N_10611,N_12164);
and U12870 (N_12870,N_12127,N_10838);
nor U12871 (N_12871,N_11909,N_11294);
or U12872 (N_12872,N_10045,N_10330);
nor U12873 (N_12873,N_11094,N_11448);
xor U12874 (N_12874,N_10856,N_11175);
nand U12875 (N_12875,N_10748,N_11451);
nor U12876 (N_12876,N_11952,N_11926);
nand U12877 (N_12877,N_10034,N_11574);
or U12878 (N_12878,N_11737,N_11178);
nor U12879 (N_12879,N_10370,N_11533);
xor U12880 (N_12880,N_11809,N_10735);
and U12881 (N_12881,N_10014,N_10137);
nand U12882 (N_12882,N_10867,N_10234);
or U12883 (N_12883,N_11347,N_10656);
nor U12884 (N_12884,N_11671,N_12083);
nor U12885 (N_12885,N_11477,N_10240);
and U12886 (N_12886,N_10772,N_10851);
and U12887 (N_12887,N_11866,N_12209);
nor U12888 (N_12888,N_11805,N_12382);
and U12889 (N_12889,N_10048,N_10591);
and U12890 (N_12890,N_11474,N_11490);
and U12891 (N_12891,N_10963,N_11886);
or U12892 (N_12892,N_11863,N_10082);
nand U12893 (N_12893,N_12349,N_12143);
nand U12894 (N_12894,N_11565,N_11582);
or U12895 (N_12895,N_11522,N_12363);
xnor U12896 (N_12896,N_12075,N_10194);
and U12897 (N_12897,N_12088,N_12376);
or U12898 (N_12898,N_12050,N_11068);
xnor U12899 (N_12899,N_11549,N_11008);
nand U12900 (N_12900,N_10872,N_12441);
and U12901 (N_12901,N_11039,N_12412);
xor U12902 (N_12902,N_12252,N_10177);
nor U12903 (N_12903,N_10946,N_10251);
xor U12904 (N_12904,N_11872,N_10423);
or U12905 (N_12905,N_10927,N_10750);
nand U12906 (N_12906,N_10564,N_11894);
or U12907 (N_12907,N_11424,N_10703);
nand U12908 (N_12908,N_11536,N_12340);
xnor U12909 (N_12909,N_10302,N_11026);
and U12910 (N_12910,N_11662,N_11006);
nor U12911 (N_12911,N_10138,N_12210);
xnor U12912 (N_12912,N_11135,N_11438);
and U12913 (N_12913,N_10279,N_10878);
nor U12914 (N_12914,N_11483,N_10035);
or U12915 (N_12915,N_12329,N_11126);
xor U12916 (N_12916,N_11705,N_12437);
or U12917 (N_12917,N_11842,N_10813);
xor U12918 (N_12918,N_12053,N_11612);
nor U12919 (N_12919,N_10707,N_10020);
or U12920 (N_12920,N_12034,N_12305);
and U12921 (N_12921,N_12080,N_10277);
and U12922 (N_12922,N_10374,N_10879);
or U12923 (N_12923,N_10393,N_11113);
or U12924 (N_12924,N_11083,N_11401);
and U12925 (N_12925,N_12007,N_11695);
or U12926 (N_12926,N_12451,N_10560);
and U12927 (N_12927,N_11193,N_10695);
xnor U12928 (N_12928,N_10375,N_10607);
nor U12929 (N_12929,N_10888,N_11016);
and U12930 (N_12930,N_10661,N_12048);
nand U12931 (N_12931,N_12492,N_11259);
nand U12932 (N_12932,N_11777,N_12356);
xnor U12933 (N_12933,N_10826,N_12063);
and U12934 (N_12934,N_10554,N_11305);
nand U12935 (N_12935,N_11437,N_11162);
or U12936 (N_12936,N_10590,N_11494);
nor U12937 (N_12937,N_11962,N_10522);
nand U12938 (N_12938,N_10264,N_10804);
and U12939 (N_12939,N_12085,N_12301);
and U12940 (N_12940,N_11585,N_12110);
nor U12941 (N_12941,N_11736,N_11444);
nand U12942 (N_12942,N_12325,N_10733);
nand U12943 (N_12943,N_11779,N_11325);
nand U12944 (N_12944,N_11827,N_11306);
nand U12945 (N_12945,N_11361,N_10046);
nand U12946 (N_12946,N_10521,N_11802);
nor U12947 (N_12947,N_11931,N_11223);
nor U12948 (N_12948,N_11624,N_11862);
nand U12949 (N_12949,N_11738,N_12205);
and U12950 (N_12950,N_11149,N_10825);
or U12951 (N_12951,N_11040,N_11376);
xor U12952 (N_12952,N_10672,N_12417);
nor U12953 (N_12953,N_11790,N_10163);
or U12954 (N_12954,N_11408,N_10503);
nand U12955 (N_12955,N_12197,N_12000);
nor U12956 (N_12956,N_10967,N_11374);
xor U12957 (N_12957,N_11803,N_11189);
nand U12958 (N_12958,N_11240,N_11403);
nand U12959 (N_12959,N_12031,N_12128);
and U12960 (N_12960,N_10730,N_11760);
nor U12961 (N_12961,N_10523,N_10076);
nor U12962 (N_12962,N_11258,N_11630);
nand U12963 (N_12963,N_11224,N_12401);
and U12964 (N_12964,N_11021,N_10908);
nor U12965 (N_12965,N_10601,N_12130);
xnor U12966 (N_12966,N_12220,N_11648);
or U12967 (N_12967,N_12187,N_11079);
xor U12968 (N_12968,N_11719,N_10829);
and U12969 (N_12969,N_10331,N_10299);
or U12970 (N_12970,N_12438,N_10161);
or U12971 (N_12971,N_10776,N_11334);
xor U12972 (N_12972,N_11634,N_11666);
and U12973 (N_12973,N_12453,N_12006);
nand U12974 (N_12974,N_10828,N_10140);
nor U12975 (N_12975,N_11252,N_11826);
and U12976 (N_12976,N_11117,N_11945);
or U12977 (N_12977,N_10977,N_10987);
nor U12978 (N_12978,N_12292,N_11213);
or U12979 (N_12979,N_11431,N_11460);
and U12980 (N_12980,N_11929,N_11528);
nand U12981 (N_12981,N_12465,N_10915);
xor U12982 (N_12982,N_10683,N_12350);
or U12983 (N_12983,N_11858,N_11922);
nor U12984 (N_12984,N_12016,N_10589);
and U12985 (N_12985,N_11242,N_10185);
nor U12986 (N_12986,N_11184,N_10428);
and U12987 (N_12987,N_10774,N_10193);
or U12988 (N_12988,N_12233,N_10945);
and U12989 (N_12989,N_11659,N_11537);
and U12990 (N_12990,N_10497,N_11708);
nand U12991 (N_12991,N_12168,N_10286);
nand U12992 (N_12992,N_10261,N_10069);
and U12993 (N_12993,N_12186,N_11453);
nand U12994 (N_12994,N_10373,N_12179);
and U12995 (N_12995,N_11729,N_10959);
nor U12996 (N_12996,N_11078,N_10209);
and U12997 (N_12997,N_11932,N_11254);
and U12998 (N_12998,N_11973,N_10653);
nor U12999 (N_12999,N_12009,N_10226);
or U13000 (N_13000,N_11605,N_11684);
and U13001 (N_13001,N_12093,N_11608);
nor U13002 (N_13002,N_11157,N_10074);
nor U13003 (N_13003,N_10387,N_11567);
and U13004 (N_13004,N_12030,N_12201);
or U13005 (N_13005,N_10962,N_12036);
or U13006 (N_13006,N_11310,N_11829);
or U13007 (N_13007,N_11385,N_10784);
or U13008 (N_13008,N_12409,N_11206);
nand U13009 (N_13009,N_10809,N_11466);
and U13010 (N_13010,N_10262,N_10762);
nand U13011 (N_13011,N_10725,N_10200);
xor U13012 (N_13012,N_12060,N_11204);
and U13013 (N_13013,N_10419,N_10458);
or U13014 (N_13014,N_11626,N_12309);
nand U13015 (N_13015,N_10544,N_10019);
or U13016 (N_13016,N_10043,N_11968);
or U13017 (N_13017,N_10934,N_10999);
or U13018 (N_13018,N_10215,N_11088);
nor U13019 (N_13019,N_10641,N_10009);
xor U13020 (N_13020,N_11542,N_12331);
nor U13021 (N_13021,N_10517,N_11045);
nor U13022 (N_13022,N_11234,N_10986);
or U13023 (N_13023,N_11712,N_11883);
nor U13024 (N_13024,N_11187,N_12236);
nor U13025 (N_13025,N_11757,N_11673);
and U13026 (N_13026,N_10787,N_10957);
nor U13027 (N_13027,N_10951,N_11092);
nor U13028 (N_13028,N_11589,N_11300);
nand U13029 (N_13029,N_10765,N_11731);
nor U13030 (N_13030,N_11985,N_11562);
nand U13031 (N_13031,N_11228,N_11947);
and U13032 (N_13032,N_11806,N_12259);
and U13033 (N_13033,N_10244,N_10214);
nand U13034 (N_13034,N_10441,N_11308);
or U13035 (N_13035,N_12432,N_10731);
nand U13036 (N_13036,N_12194,N_11813);
nor U13037 (N_13037,N_11262,N_10551);
nor U13038 (N_13038,N_11405,N_12111);
and U13039 (N_13039,N_10536,N_11167);
xor U13040 (N_13040,N_10911,N_10546);
xor U13041 (N_13041,N_10068,N_12394);
nand U13042 (N_13042,N_12499,N_11640);
and U13043 (N_13043,N_11814,N_12145);
nand U13044 (N_13044,N_10939,N_10380);
or U13045 (N_13045,N_10668,N_12150);
nor U13046 (N_13046,N_10080,N_11446);
nor U13047 (N_13047,N_11638,N_10461);
xor U13048 (N_13048,N_10095,N_11940);
xnor U13049 (N_13049,N_11014,N_12494);
and U13050 (N_13050,N_11440,N_11871);
nor U13051 (N_13051,N_11688,N_12138);
and U13052 (N_13052,N_10119,N_10389);
and U13053 (N_13053,N_12267,N_11572);
or U13054 (N_13054,N_11776,N_11910);
nor U13055 (N_13055,N_10783,N_10689);
and U13056 (N_13056,N_11739,N_12454);
nand U13057 (N_13057,N_10799,N_10116);
and U13058 (N_13058,N_11868,N_11377);
nor U13059 (N_13059,N_11820,N_11365);
and U13060 (N_13060,N_11888,N_10223);
and U13061 (N_13061,N_11546,N_10071);
nand U13062 (N_13062,N_10746,N_11597);
xor U13063 (N_13063,N_11501,N_11073);
xnor U13064 (N_13064,N_12062,N_10230);
and U13065 (N_13065,N_10577,N_10047);
or U13066 (N_13066,N_10676,N_12097);
nor U13067 (N_13067,N_10390,N_12319);
nor U13068 (N_13068,N_10588,N_11329);
xor U13069 (N_13069,N_11366,N_11030);
nand U13070 (N_13070,N_10073,N_10167);
nand U13071 (N_13071,N_11746,N_11764);
and U13072 (N_13072,N_11595,N_12277);
and U13073 (N_13073,N_10211,N_11378);
nand U13074 (N_13074,N_10424,N_10627);
nor U13075 (N_13075,N_11020,N_10421);
nor U13076 (N_13076,N_10320,N_11428);
nor U13077 (N_13077,N_11556,N_10973);
and U13078 (N_13078,N_11650,N_10629);
nor U13079 (N_13079,N_11808,N_10334);
nor U13080 (N_13080,N_12293,N_10222);
xnor U13081 (N_13081,N_10961,N_10814);
nor U13082 (N_13082,N_10763,N_11349);
nor U13083 (N_13083,N_10007,N_12103);
and U13084 (N_13084,N_11665,N_11290);
nand U13085 (N_13085,N_12183,N_10552);
nor U13086 (N_13086,N_11848,N_10649);
nand U13087 (N_13087,N_12391,N_10907);
xnor U13088 (N_13088,N_12200,N_10107);
xor U13089 (N_13089,N_11753,N_11066);
nor U13090 (N_13090,N_10482,N_10318);
nor U13091 (N_13091,N_11840,N_10686);
nor U13092 (N_13092,N_10276,N_10779);
and U13093 (N_13093,N_10567,N_11845);
nand U13094 (N_13094,N_11115,N_11925);
or U13095 (N_13095,N_10378,N_11696);
nor U13096 (N_13096,N_10038,N_11024);
or U13097 (N_13097,N_12371,N_10534);
nand U13098 (N_13098,N_11398,N_10605);
or U13099 (N_13099,N_12493,N_10391);
or U13100 (N_13100,N_11169,N_11918);
nor U13101 (N_13101,N_11358,N_11950);
nand U13102 (N_13102,N_12232,N_10854);
and U13103 (N_13103,N_10791,N_11660);
nor U13104 (N_13104,N_11248,N_10868);
nand U13105 (N_13105,N_12328,N_10728);
or U13106 (N_13106,N_11765,N_10050);
and U13107 (N_13107,N_11609,N_10902);
and U13108 (N_13108,N_11093,N_12370);
and U13109 (N_13109,N_11975,N_10810);
and U13110 (N_13110,N_11367,N_11514);
nor U13111 (N_13111,N_10476,N_10688);
nand U13112 (N_13112,N_10145,N_10411);
and U13113 (N_13113,N_12137,N_12229);
nand U13114 (N_13114,N_10984,N_11749);
and U13115 (N_13115,N_12450,N_12156);
xnor U13116 (N_13116,N_10778,N_12106);
xor U13117 (N_13117,N_10989,N_10692);
xor U13118 (N_13118,N_12428,N_10718);
or U13119 (N_13119,N_11509,N_10316);
nand U13120 (N_13120,N_10658,N_10343);
xnor U13121 (N_13121,N_11080,N_12092);
nor U13122 (N_13122,N_10855,N_11755);
nand U13123 (N_13123,N_10926,N_12114);
nand U13124 (N_13124,N_10593,N_12390);
or U13125 (N_13125,N_10178,N_12067);
and U13126 (N_13126,N_11455,N_11923);
nor U13127 (N_13127,N_10475,N_11678);
or U13128 (N_13128,N_12261,N_12002);
nand U13129 (N_13129,N_10499,N_10363);
xnor U13130 (N_13130,N_12369,N_10062);
or U13131 (N_13131,N_11138,N_11908);
and U13132 (N_13132,N_10213,N_11831);
nand U13133 (N_13133,N_11617,N_11984);
and U13134 (N_13134,N_11475,N_10858);
xnor U13135 (N_13135,N_12202,N_12173);
and U13136 (N_13136,N_12193,N_11140);
and U13137 (N_13137,N_12005,N_10850);
nor U13138 (N_13138,N_11041,N_11004);
nand U13139 (N_13139,N_12198,N_11900);
xor U13140 (N_13140,N_11145,N_10139);
xnor U13141 (N_13141,N_10379,N_11623);
xnor U13142 (N_13142,N_10117,N_11200);
nand U13143 (N_13143,N_11917,N_11220);
nand U13144 (N_13144,N_12468,N_10466);
and U13145 (N_13145,N_11270,N_12115);
or U13146 (N_13146,N_11271,N_10545);
and U13147 (N_13147,N_11304,N_11338);
nor U13148 (N_13148,N_12091,N_12353);
and U13149 (N_13149,N_11527,N_10681);
or U13150 (N_13150,N_12400,N_11027);
or U13151 (N_13151,N_10454,N_12207);
nand U13152 (N_13152,N_11698,N_10432);
or U13153 (N_13153,N_10988,N_11380);
and U13154 (N_13154,N_10754,N_11961);
nor U13155 (N_13155,N_12330,N_11732);
or U13156 (N_13156,N_10191,N_12366);
nand U13157 (N_13157,N_10578,N_11274);
or U13158 (N_13158,N_10669,N_10165);
and U13159 (N_13159,N_11921,N_10761);
nor U13160 (N_13160,N_10162,N_11773);
or U13161 (N_13161,N_11796,N_11097);
xnor U13162 (N_13162,N_12105,N_10282);
nand U13163 (N_13163,N_11661,N_11999);
nor U13164 (N_13164,N_12116,N_11710);
or U13165 (N_13165,N_11139,N_11263);
nor U13166 (N_13166,N_10636,N_12333);
nand U13167 (N_13167,N_11512,N_10631);
nor U13168 (N_13168,N_12077,N_10174);
nor U13169 (N_13169,N_11901,N_11924);
and U13170 (N_13170,N_12407,N_11530);
nor U13171 (N_13171,N_10362,N_11788);
nor U13172 (N_13172,N_11373,N_12332);
nand U13173 (N_13173,N_11155,N_11415);
or U13174 (N_13174,N_11284,N_10016);
or U13175 (N_13175,N_10260,N_11775);
or U13176 (N_13176,N_11793,N_11276);
and U13177 (N_13177,N_10930,N_10832);
or U13178 (N_13178,N_10250,N_10711);
xnor U13179 (N_13179,N_10060,N_12129);
nor U13180 (N_13180,N_10109,N_10396);
nor U13181 (N_13181,N_10408,N_11681);
or U13182 (N_13182,N_11761,N_10955);
or U13183 (N_13183,N_11905,N_12008);
nand U13184 (N_13184,N_12108,N_11730);
nand U13185 (N_13185,N_11600,N_10281);
nand U13186 (N_13186,N_10960,N_10401);
nand U13187 (N_13187,N_10027,N_10232);
and U13188 (N_13188,N_11125,N_12378);
and U13189 (N_13189,N_12271,N_11960);
nand U13190 (N_13190,N_12483,N_11709);
xnor U13191 (N_13191,N_12191,N_12387);
nor U13192 (N_13192,N_10831,N_10464);
nand U13193 (N_13193,N_11823,N_12217);
and U13194 (N_13194,N_12360,N_12180);
nand U13195 (N_13195,N_11979,N_11571);
nand U13196 (N_13196,N_11949,N_11570);
or U13197 (N_13197,N_12028,N_11576);
xnor U13198 (N_13198,N_11898,N_10188);
and U13199 (N_13199,N_11946,N_12445);
and U13200 (N_13200,N_10180,N_12427);
or U13201 (N_13201,N_10954,N_12042);
nand U13202 (N_13202,N_10905,N_12490);
nand U13203 (N_13203,N_10715,N_10372);
or U13204 (N_13204,N_10182,N_11053);
nor U13205 (N_13205,N_10571,N_10549);
nor U13206 (N_13206,N_10882,N_12081);
and U13207 (N_13207,N_10186,N_12302);
and U13208 (N_13208,N_10023,N_10864);
and U13209 (N_13209,N_10490,N_12241);
nor U13210 (N_13210,N_11942,N_10341);
xor U13211 (N_13211,N_10462,N_10446);
or U13212 (N_13212,N_12433,N_10700);
nor U13213 (N_13213,N_10453,N_10876);
and U13214 (N_13214,N_11395,N_10124);
and U13215 (N_13215,N_11018,N_11789);
and U13216 (N_13216,N_10111,N_12282);
and U13217 (N_13217,N_10500,N_10146);
or U13218 (N_13218,N_10099,N_10983);
nor U13219 (N_13219,N_11485,N_10075);
xnor U13220 (N_13220,N_11402,N_12112);
nand U13221 (N_13221,N_10051,N_11752);
nand U13222 (N_13222,N_12037,N_10899);
and U13223 (N_13223,N_11033,N_11785);
nand U13224 (N_13224,N_12426,N_11596);
or U13225 (N_13225,N_11371,N_10506);
nor U13226 (N_13226,N_12027,N_10101);
and U13227 (N_13227,N_10691,N_10065);
or U13228 (N_13228,N_11309,N_11740);
nand U13229 (N_13229,N_10057,N_11368);
nand U13230 (N_13230,N_11702,N_11561);
xnor U13231 (N_13231,N_11843,N_11291);
nor U13232 (N_13232,N_12134,N_11413);
or U13233 (N_13233,N_11104,N_10125);
or U13234 (N_13234,N_11770,N_11653);
and U13235 (N_13235,N_10847,N_12023);
nand U13236 (N_13236,N_11012,N_12466);
and U13237 (N_13237,N_11471,N_11939);
or U13238 (N_13238,N_11414,N_10392);
nand U13239 (N_13239,N_11156,N_10039);
or U13240 (N_13240,N_11061,N_11019);
or U13241 (N_13241,N_11202,N_11163);
nand U13242 (N_13242,N_12029,N_11105);
nand U13243 (N_13243,N_10642,N_10122);
nand U13244 (N_13244,N_10460,N_11754);
nand U13245 (N_13245,N_12022,N_10823);
nor U13246 (N_13246,N_11992,N_12397);
and U13247 (N_13247,N_10671,N_11602);
and U13248 (N_13248,N_12345,N_11359);
nand U13249 (N_13249,N_11280,N_11644);
nor U13250 (N_13250,N_10616,N_10965);
nand U13251 (N_13251,N_11344,N_11707);
nand U13252 (N_13252,N_10141,N_11085);
xnor U13253 (N_13253,N_10640,N_11792);
and U13254 (N_13254,N_11680,N_11063);
and U13255 (N_13255,N_10249,N_11154);
and U13256 (N_13256,N_12020,N_12379);
and U13257 (N_13257,N_12347,N_11957);
or U13258 (N_13258,N_10474,N_11607);
or U13259 (N_13259,N_10289,N_11741);
nand U13260 (N_13260,N_11264,N_11499);
nor U13261 (N_13261,N_10815,N_11669);
and U13262 (N_13262,N_10570,N_11328);
and U13263 (N_13263,N_11332,N_11459);
and U13264 (N_13264,N_11614,N_11540);
nand U13265 (N_13265,N_10647,N_10483);
nand U13266 (N_13266,N_10597,N_10818);
and U13267 (N_13267,N_10339,N_12017);
xnor U13268 (N_13268,N_10916,N_10465);
or U13269 (N_13269,N_10714,N_12403);
or U13270 (N_13270,N_11293,N_11610);
or U13271 (N_13271,N_10630,N_10118);
nor U13272 (N_13272,N_11691,N_10651);
and U13273 (N_13273,N_10326,N_11357);
nand U13274 (N_13274,N_10990,N_11445);
and U13275 (N_13275,N_11246,N_10598);
and U13276 (N_13276,N_11599,N_10110);
nand U13277 (N_13277,N_10644,N_10953);
or U13278 (N_13278,N_10272,N_11121);
and U13279 (N_13279,N_11208,N_11319);
nand U13280 (N_13280,N_11622,N_11852);
or U13281 (N_13281,N_12306,N_10133);
xnor U13282 (N_13282,N_12495,N_10836);
and U13283 (N_13283,N_10364,N_11551);
xor U13284 (N_13284,N_12174,N_10294);
and U13285 (N_13285,N_11641,N_10548);
nor U13286 (N_13286,N_11239,N_10325);
and U13287 (N_13287,N_12032,N_10098);
nand U13288 (N_13288,N_11250,N_11318);
nand U13289 (N_13289,N_10445,N_10404);
nor U13290 (N_13290,N_11017,N_12072);
and U13291 (N_13291,N_12276,N_11655);
or U13292 (N_13292,N_11194,N_11497);
or U13293 (N_13293,N_10078,N_11216);
nand U13294 (N_13294,N_11759,N_11955);
or U13295 (N_13295,N_12247,N_12341);
and U13296 (N_13296,N_10195,N_10871);
nand U13297 (N_13297,N_12170,N_10090);
or U13298 (N_13298,N_11473,N_10837);
nand U13299 (N_13299,N_10409,N_10582);
nand U13300 (N_13300,N_11457,N_10233);
and U13301 (N_13301,N_12439,N_12226);
or U13302 (N_13302,N_11352,N_10673);
nand U13303 (N_13303,N_11575,N_10736);
nand U13304 (N_13304,N_11177,N_11978);
nor U13305 (N_13305,N_11824,N_10348);
nor U13306 (N_13306,N_11971,N_10885);
and U13307 (N_13307,N_12195,N_12146);
nor U13308 (N_13308,N_10306,N_12336);
xor U13309 (N_13309,N_10241,N_10275);
nor U13310 (N_13310,N_10094,N_10830);
and U13311 (N_13311,N_10198,N_11508);
and U13312 (N_13312,N_10716,N_11095);
xnor U13313 (N_13313,N_11882,N_10835);
nand U13314 (N_13314,N_11654,N_10894);
nor U13315 (N_13315,N_11904,N_11834);
nand U13316 (N_13316,N_12402,N_10793);
xor U13317 (N_13317,N_12290,N_11188);
or U13318 (N_13318,N_12352,N_10775);
or U13319 (N_13319,N_11356,N_10701);
and U13320 (N_13320,N_12295,N_10594);
and U13321 (N_13321,N_12380,N_12211);
nor U13322 (N_13322,N_10526,N_11277);
xnor U13323 (N_13323,N_10664,N_12074);
or U13324 (N_13324,N_12270,N_12181);
and U13325 (N_13325,N_11243,N_11119);
nand U13326 (N_13326,N_10444,N_10726);
or U13327 (N_13327,N_11647,N_11420);
nor U13328 (N_13328,N_11480,N_11721);
nor U13329 (N_13329,N_11544,N_12058);
and U13330 (N_13330,N_12019,N_10003);
and U13331 (N_13331,N_10512,N_11179);
xor U13332 (N_13332,N_12121,N_12279);
xnor U13333 (N_13333,N_10494,N_11456);
or U13334 (N_13334,N_12192,N_12312);
nor U13335 (N_13335,N_11447,N_11890);
and U13336 (N_13336,N_10524,N_10479);
nor U13337 (N_13337,N_11937,N_10797);
nor U13338 (N_13338,N_10956,N_10371);
nor U13339 (N_13339,N_10786,N_10487);
nand U13340 (N_13340,N_11129,N_12479);
nand U13341 (N_13341,N_12133,N_11781);
and U13342 (N_13342,N_11479,N_11763);
xor U13343 (N_13343,N_10295,N_11718);
and U13344 (N_13344,N_12317,N_11878);
nor U13345 (N_13345,N_12065,N_11435);
and U13346 (N_13346,N_10833,N_11219);
and U13347 (N_13347,N_10860,N_11481);
and U13348 (N_13348,N_10862,N_11711);
nand U13349 (N_13349,N_11970,N_11976);
or U13350 (N_13350,N_12489,N_12155);
or U13351 (N_13351,N_11977,N_11745);
nand U13352 (N_13352,N_11742,N_10425);
nor U13353 (N_13353,N_10811,N_11525);
and U13354 (N_13354,N_11404,N_12296);
nand U13355 (N_13355,N_10297,N_11038);
or U13356 (N_13356,N_10212,N_11381);
nand U13357 (N_13357,N_10157,N_10040);
or U13358 (N_13358,N_11912,N_10807);
and U13359 (N_13359,N_11722,N_11689);
nand U13360 (N_13360,N_11151,N_11835);
nand U13361 (N_13361,N_10055,N_11072);
and U13362 (N_13362,N_10231,N_10365);
nor U13363 (N_13363,N_11226,N_11645);
nand U13364 (N_13364,N_11791,N_11098);
nor U13365 (N_13365,N_12119,N_11550);
xor U13366 (N_13366,N_11047,N_11176);
nand U13367 (N_13367,N_12314,N_11307);
nor U13368 (N_13368,N_10972,N_10336);
nand U13369 (N_13369,N_11084,N_10298);
nor U13370 (N_13370,N_11998,N_10991);
nor U13371 (N_13371,N_11409,N_11275);
and U13372 (N_13372,N_11836,N_11604);
or U13373 (N_13373,N_10031,N_11538);
nand U13374 (N_13374,N_11036,N_10257);
xnor U13375 (N_13375,N_10006,N_10170);
or U13376 (N_13376,N_11191,N_11222);
or U13377 (N_13377,N_11498,N_10358);
nand U13378 (N_13378,N_12446,N_10755);
or U13379 (N_13379,N_10344,N_12015);
or U13380 (N_13380,N_10981,N_11441);
or U13381 (N_13381,N_10537,N_10267);
nor U13382 (N_13382,N_11573,N_12184);
or U13383 (N_13383,N_11555,N_11867);
nor U13384 (N_13384,N_10756,N_10740);
nor U13385 (N_13385,N_10768,N_11928);
or U13386 (N_13386,N_11615,N_10518);
nor U13387 (N_13387,N_12256,N_12284);
nor U13388 (N_13388,N_10274,N_12254);
and U13389 (N_13389,N_11686,N_10619);
nand U13390 (N_13390,N_10684,N_10948);
nand U13391 (N_13391,N_10005,N_10505);
nand U13392 (N_13392,N_11724,N_11336);
and U13393 (N_13393,N_11077,N_11383);
or U13394 (N_13394,N_12045,N_10865);
and U13395 (N_13395,N_10904,N_11519);
nand U13396 (N_13396,N_11758,N_12082);
nand U13397 (N_13397,N_10509,N_12222);
and U13398 (N_13398,N_12043,N_11247);
nor U13399 (N_13399,N_11584,N_11701);
or U13400 (N_13400,N_10550,N_11593);
nor U13401 (N_13401,N_10869,N_11651);
or U13402 (N_13402,N_12144,N_11340);
and U13403 (N_13403,N_10437,N_11137);
nand U13404 (N_13404,N_10399,N_10771);
or U13405 (N_13405,N_12098,N_10877);
or U13406 (N_13406,N_10980,N_12484);
and U13407 (N_13407,N_11554,N_11854);
nand U13408 (N_13408,N_11628,N_10947);
nor U13409 (N_13409,N_10922,N_12089);
and U13410 (N_13410,N_10443,N_10639);
and U13411 (N_13411,N_11966,N_11816);
and U13412 (N_13412,N_12478,N_11427);
nor U13413 (N_13413,N_10103,N_12395);
and U13414 (N_13414,N_10451,N_11463);
or U13415 (N_13415,N_10753,N_11988);
and U13416 (N_13416,N_11911,N_10463);
or U13417 (N_13417,N_11590,N_11075);
nand U13418 (N_13418,N_10456,N_12040);
or U13419 (N_13419,N_10936,N_11051);
nand U13420 (N_13420,N_12038,N_10766);
xnor U13421 (N_13421,N_10952,N_11830);
and U13422 (N_13422,N_10667,N_10402);
nand U13423 (N_13423,N_12456,N_11387);
and U13424 (N_13424,N_11442,N_12230);
nand U13425 (N_13425,N_11059,N_12269);
nand U13426 (N_13426,N_10632,N_10599);
nand U13427 (N_13427,N_10012,N_10398);
nor U13428 (N_13428,N_11173,N_10614);
xor U13429 (N_13429,N_11865,N_10407);
nor U13430 (N_13430,N_10764,N_10056);
or U13431 (N_13431,N_11406,N_10802);
nor U13432 (N_13432,N_11578,N_10481);
or U13433 (N_13433,N_10328,N_11316);
or U13434 (N_13434,N_12117,N_10713);
or U13435 (N_13435,N_12326,N_12386);
nor U13436 (N_13436,N_12039,N_11639);
and U13437 (N_13437,N_11963,N_11282);
nor U13438 (N_13438,N_12227,N_11794);
nand U13439 (N_13439,N_11849,N_10757);
xnor U13440 (N_13440,N_11422,N_10652);
or U13441 (N_13441,N_12096,N_12213);
nand U13442 (N_13442,N_12272,N_12464);
and U13443 (N_13443,N_10665,N_11959);
or U13444 (N_13444,N_12268,N_11772);
or U13445 (N_13445,N_11687,N_10197);
nor U13446 (N_13446,N_10722,N_11345);
or U13447 (N_13447,N_12344,N_10886);
nand U13448 (N_13448,N_11257,N_10937);
nand U13449 (N_13449,N_10675,N_12167);
or U13450 (N_13450,N_10529,N_10606);
or U13451 (N_13451,N_11165,N_11625);
nand U13452 (N_13452,N_12214,N_12408);
and U13453 (N_13453,N_12148,N_11756);
or U13454 (N_13454,N_11983,N_11735);
nor U13455 (N_13455,N_10052,N_10207);
nor U13456 (N_13456,N_11450,N_10121);
or U13457 (N_13457,N_10042,N_10112);
or U13458 (N_13458,N_11348,N_10994);
nand U13459 (N_13459,N_11048,N_11974);
and U13460 (N_13460,N_11601,N_11668);
nor U13461 (N_13461,N_10660,N_12125);
or U13462 (N_13462,N_10584,N_10013);
and U13463 (N_13463,N_11164,N_10893);
nand U13464 (N_13464,N_11692,N_10844);
or U13465 (N_13465,N_12487,N_11180);
nor U13466 (N_13466,N_10645,N_11353);
or U13467 (N_13467,N_11860,N_10114);
nand U13468 (N_13468,N_11127,N_11292);
and U13469 (N_13469,N_11621,N_12448);
nor U13470 (N_13470,N_11425,N_11850);
nand U13471 (N_13471,N_12090,N_10738);
nor U13472 (N_13472,N_11272,N_10875);
xor U13473 (N_13473,N_10092,N_11493);
nor U13474 (N_13474,N_12102,N_10469);
or U13475 (N_13475,N_11853,N_11108);
nand U13476 (N_13476,N_12383,N_10887);
nand U13477 (N_13477,N_10928,N_12264);
and U13478 (N_13478,N_11951,N_12273);
or U13479 (N_13479,N_11716,N_10555);
nand U13480 (N_13480,N_10059,N_11214);
or U13481 (N_13481,N_10816,N_11539);
and U13482 (N_13482,N_10903,N_12421);
or U13483 (N_13483,N_10699,N_11725);
nand U13484 (N_13484,N_11462,N_10142);
and U13485 (N_13485,N_11658,N_10958);
and U13486 (N_13486,N_10252,N_10812);
or U13487 (N_13487,N_10798,N_11046);
xnor U13488 (N_13488,N_10204,N_10002);
nor U13489 (N_13489,N_10327,N_12475);
nand U13490 (N_13490,N_11397,N_10519);
nand U13491 (N_13491,N_10022,N_12159);
nor U13492 (N_13492,N_10511,N_11611);
and U13493 (N_13493,N_11236,N_10709);
nand U13494 (N_13494,N_10997,N_11798);
nor U13495 (N_13495,N_11649,N_11326);
nor U13496 (N_13496,N_11394,N_10866);
and U13497 (N_13497,N_10253,N_12203);
nor U13498 (N_13498,N_10643,N_10173);
nand U13499 (N_13499,N_10270,N_10976);
or U13500 (N_13500,N_10070,N_11897);
nand U13501 (N_13501,N_11171,N_10543);
nor U13502 (N_13502,N_10105,N_10189);
or U13503 (N_13503,N_10449,N_11837);
and U13504 (N_13504,N_10624,N_10011);
or U13505 (N_13505,N_11504,N_12245);
nand U13506 (N_13506,N_10561,N_12321);
xor U13507 (N_13507,N_10164,N_11632);
nor U13508 (N_13508,N_10531,N_10949);
xnor U13509 (N_13509,N_10029,N_11861);
and U13510 (N_13510,N_11887,N_10147);
nand U13511 (N_13511,N_11543,N_12171);
nand U13512 (N_13512,N_11568,N_11564);
nor U13513 (N_13513,N_10026,N_12166);
nand U13514 (N_13514,N_11547,N_10592);
nand U13515 (N_13515,N_10623,N_10259);
nand U13516 (N_13516,N_10874,N_12122);
nand U13517 (N_13517,N_10455,N_10852);
or U13518 (N_13518,N_10933,N_11390);
xor U13519 (N_13519,N_11423,N_11265);
nand U13520 (N_13520,N_10626,N_11646);
or U13521 (N_13521,N_10800,N_11210);
nor U13522 (N_13522,N_10054,N_12123);
nand U13523 (N_13523,N_11044,N_10595);
or U13524 (N_13524,N_11421,N_10720);
and U13525 (N_13525,N_11339,N_10179);
and U13526 (N_13526,N_12381,N_11819);
nand U13527 (N_13527,N_10300,N_10690);
nor U13528 (N_13528,N_10087,N_10982);
nor U13529 (N_13529,N_11965,N_10382);
nor U13530 (N_13530,N_12430,N_11035);
nor U13531 (N_13531,N_11197,N_10135);
nand U13532 (N_13532,N_11341,N_11260);
or U13533 (N_13533,N_10126,N_10216);
nand U13534 (N_13534,N_10347,N_12288);
or U13535 (N_13535,N_10613,N_11591);
nand U13536 (N_13536,N_10702,N_10028);
xnor U13537 (N_13537,N_12177,N_11109);
and U13538 (N_13538,N_11467,N_11468);
nor U13539 (N_13539,N_11652,N_10895);
and U13540 (N_13540,N_11042,N_11704);
or U13541 (N_13541,N_11620,N_10159);
nor U13542 (N_13542,N_10210,N_12480);
or U13543 (N_13543,N_11000,N_12375);
or U13544 (N_13544,N_10290,N_11750);
and U13545 (N_13545,N_11237,N_10568);
and U13546 (N_13546,N_10657,N_10924);
nand U13547 (N_13547,N_11889,N_11523);
and U13548 (N_13548,N_12141,N_11131);
or U13549 (N_13549,N_12342,N_11470);
or U13550 (N_13550,N_10917,N_10171);
nor U13551 (N_13551,N_12339,N_12462);
and U13552 (N_13552,N_11545,N_11412);
or U13553 (N_13553,N_10566,N_11838);
xor U13554 (N_13554,N_12157,N_10030);
xnor U13555 (N_13555,N_12196,N_10569);
or U13556 (N_13556,N_11301,N_10603);
nor U13557 (N_13557,N_11289,N_10376);
nand U13558 (N_13558,N_11717,N_12069);
and U13559 (N_13559,N_11062,N_11847);
or U13560 (N_13560,N_10848,N_10925);
and U13561 (N_13561,N_10439,N_11267);
nand U13562 (N_13562,N_10583,N_10307);
or U13563 (N_13563,N_11386,N_12013);
and U13564 (N_13564,N_11324,N_10395);
and U13565 (N_13565,N_11160,N_10698);
or U13566 (N_13566,N_12318,N_10900);
nand U13567 (N_13567,N_11714,N_11212);
xor U13568 (N_13568,N_11096,N_10400);
or U13569 (N_13569,N_11279,N_12239);
or U13570 (N_13570,N_10414,N_12162);
nand U13571 (N_13571,N_12046,N_11594);
and U13572 (N_13572,N_12485,N_11943);
nand U13573 (N_13573,N_10072,N_12182);
or U13574 (N_13574,N_11181,N_10729);
or U13575 (N_13575,N_10333,N_10229);
nand U13576 (N_13576,N_11436,N_12334);
and U13577 (N_13577,N_10743,N_11697);
and U13578 (N_13578,N_11144,N_12357);
nor U13579 (N_13579,N_11141,N_11495);
and U13580 (N_13580,N_10846,N_12242);
xor U13581 (N_13581,N_12025,N_12413);
and U13582 (N_13582,N_12262,N_10350);
nand U13583 (N_13583,N_10789,N_12255);
and U13584 (N_13584,N_10225,N_10609);
and U13585 (N_13585,N_10017,N_11778);
or U13586 (N_13586,N_11864,N_11994);
or U13587 (N_13587,N_10540,N_11557);
nor U13588 (N_13588,N_10351,N_10739);
nand U13589 (N_13589,N_12476,N_11592);
and U13590 (N_13590,N_11266,N_11566);
or U13591 (N_13591,N_10941,N_10760);
nor U13592 (N_13592,N_11579,N_11587);
nand U13593 (N_13593,N_10010,N_10863);
and U13594 (N_13594,N_12154,N_11211);
and U13595 (N_13595,N_11679,N_12059);
or U13596 (N_13596,N_12212,N_10329);
and U13597 (N_13597,N_12443,N_12410);
or U13598 (N_13598,N_10349,N_11893);
nor U13599 (N_13599,N_11833,N_10394);
and U13600 (N_13600,N_11667,N_11037);
nor U13601 (N_13601,N_10507,N_10293);
nor U13602 (N_13602,N_12498,N_10806);
nand U13603 (N_13603,N_11675,N_10254);
nor U13604 (N_13604,N_11185,N_11635);
or U13605 (N_13605,N_10360,N_10422);
nor U13606 (N_13606,N_12281,N_10381);
or U13607 (N_13607,N_10516,N_11429);
or U13608 (N_13608,N_12275,N_11771);
and U13609 (N_13609,N_11991,N_11743);
nand U13610 (N_13610,N_11116,N_12238);
nor U13611 (N_13611,N_10998,N_10361);
nand U13612 (N_13612,N_10530,N_11953);
and U13613 (N_13613,N_12404,N_11031);
or U13614 (N_13614,N_11244,N_10638);
nor U13615 (N_13615,N_11507,N_10308);
nand U13616 (N_13616,N_10155,N_11936);
or U13617 (N_13617,N_10880,N_12055);
or U13618 (N_13618,N_11476,N_11563);
or U13619 (N_13619,N_10921,N_11360);
nand U13620 (N_13620,N_10079,N_10426);
or U13621 (N_13621,N_12455,N_12389);
or U13622 (N_13622,N_11209,N_11174);
or U13623 (N_13623,N_10129,N_11677);
nand U13624 (N_13624,N_12434,N_11685);
and U13625 (N_13625,N_11054,N_11618);
nand U13626 (N_13626,N_11896,N_11411);
xor U13627 (N_13627,N_11086,N_10705);
or U13628 (N_13628,N_11132,N_11124);
nand U13629 (N_13629,N_11521,N_11134);
nor U13630 (N_13630,N_11443,N_11337);
nor U13631 (N_13631,N_11907,N_10650);
and U13632 (N_13632,N_10247,N_10528);
nand U13633 (N_13633,N_11241,N_11927);
or U13634 (N_13634,N_11693,N_11183);
nand U13635 (N_13635,N_11941,N_11056);
nand U13636 (N_13636,N_10201,N_12414);
and U13637 (N_13637,N_10819,N_11317);
nor U13638 (N_13638,N_10278,N_11987);
nand U13639 (N_13639,N_10892,N_10175);
nand U13640 (N_13640,N_12185,N_10000);
nor U13641 (N_13641,N_12457,N_12176);
nand U13642 (N_13642,N_10115,N_11857);
nand U13643 (N_13643,N_11529,N_11410);
xnor U13644 (N_13644,N_10712,N_11532);
and U13645 (N_13645,N_11230,N_11583);
and U13646 (N_13646,N_11146,N_11055);
or U13647 (N_13647,N_11683,N_10621);
nor U13648 (N_13648,N_10256,N_10448);
and U13649 (N_13649,N_10985,N_10685);
or U13650 (N_13650,N_12263,N_12365);
and U13651 (N_13651,N_10008,N_10049);
nand U13652 (N_13652,N_10044,N_10061);
and U13653 (N_13653,N_11920,N_12274);
nor U13654 (N_13654,N_11221,N_11182);
and U13655 (N_13655,N_10342,N_12140);
and U13656 (N_13656,N_12076,N_11997);
nor U13657 (N_13657,N_11619,N_11207);
xor U13658 (N_13658,N_12161,N_12278);
nand U13659 (N_13659,N_12225,N_10127);
nand U13660 (N_13660,N_10796,N_12460);
or U13661 (N_13661,N_11744,N_11013);
nand U13662 (N_13662,N_11168,N_11136);
and U13663 (N_13663,N_11285,N_10820);
nand U13664 (N_13664,N_12001,N_11074);
or U13665 (N_13665,N_11399,N_10777);
nand U13666 (N_13666,N_10995,N_11090);
nor U13667 (N_13667,N_10288,N_11071);
or U13668 (N_13668,N_10021,N_10572);
or U13669 (N_13669,N_12153,N_12477);
nor U13670 (N_13670,N_10790,N_11103);
nor U13671 (N_13671,N_11407,N_11120);
and U13672 (N_13672,N_12018,N_11524);
or U13673 (N_13673,N_11956,N_12304);
and U13674 (N_13674,N_11321,N_12310);
nand U13675 (N_13675,N_11161,N_12084);
or U13676 (N_13676,N_10759,N_11148);
nor U13677 (N_13677,N_10839,N_11967);
or U13678 (N_13678,N_10919,N_10314);
nand U13679 (N_13679,N_12208,N_11369);
nand U13680 (N_13680,N_11034,N_11418);
nand U13681 (N_13681,N_10472,N_12419);
nand U13682 (N_13682,N_11484,N_11690);
nor U13683 (N_13683,N_11703,N_10305);
or U13684 (N_13684,N_12248,N_10565);
nor U13685 (N_13685,N_11832,N_12481);
xnor U13686 (N_13686,N_11142,N_11986);
nand U13687 (N_13687,N_10520,N_11870);
nand U13688 (N_13688,N_12044,N_10337);
and U13689 (N_13689,N_11287,N_10471);
and U13690 (N_13690,N_11616,N_12244);
nand U13691 (N_13691,N_12442,N_10496);
xnor U13692 (N_13692,N_11333,N_10498);
or U13693 (N_13693,N_11400,N_11958);
or U13694 (N_13694,N_10602,N_10436);
nor U13695 (N_13695,N_10891,N_10803);
nor U13696 (N_13696,N_11767,N_10504);
nand U13697 (N_13697,N_10795,N_11891);
and U13698 (N_13698,N_10208,N_10315);
or U13699 (N_13699,N_10310,N_10912);
nor U13700 (N_13700,N_10576,N_10324);
or U13701 (N_13701,N_11506,N_10356);
nor U13702 (N_13702,N_10473,N_12324);
and U13703 (N_13703,N_10149,N_12285);
nand U13704 (N_13704,N_10694,N_12411);
or U13705 (N_13705,N_12231,N_11782);
nand U13706 (N_13706,N_10085,N_11822);
xnor U13707 (N_13707,N_10089,N_10285);
nand U13708 (N_13708,N_10747,N_10539);
nand U13709 (N_13709,N_12132,N_10100);
nand U13710 (N_13710,N_10782,N_12449);
and U13711 (N_13711,N_10434,N_12163);
or U13712 (N_13712,N_11995,N_12012);
nand U13713 (N_13713,N_10918,N_12135);
nor U13714 (N_13714,N_11915,N_10273);
nor U13715 (N_13715,N_10562,N_11699);
or U13716 (N_13716,N_10184,N_11795);
and U13717 (N_13717,N_11050,N_11112);
and U13718 (N_13718,N_12070,N_10292);
nand U13719 (N_13719,N_10618,N_11913);
xnor U13720 (N_13720,N_12286,N_10346);
or U13721 (N_13721,N_10553,N_11393);
or U13722 (N_13722,N_10128,N_12396);
xnor U13723 (N_13723,N_10579,N_10890);
or U13724 (N_13724,N_10335,N_12398);
and U13725 (N_13725,N_12223,N_12300);
or U13726 (N_13726,N_10502,N_11944);
or U13727 (N_13727,N_10187,N_10687);
nor U13728 (N_13728,N_10501,N_10417);
or U13729 (N_13729,N_12068,N_10104);
and U13730 (N_13730,N_11342,N_11192);
or U13731 (N_13731,N_12393,N_10785);
xnor U13732 (N_13732,N_10873,N_10514);
nand U13733 (N_13733,N_10053,N_12294);
and U13734 (N_13734,N_11728,N_11150);
or U13735 (N_13735,N_10604,N_10219);
nor U13736 (N_13736,N_11982,N_10322);
xor U13737 (N_13737,N_10431,N_11298);
or U13738 (N_13738,N_11433,N_11343);
or U13739 (N_13739,N_11769,N_12216);
and U13740 (N_13740,N_10780,N_10821);
or U13741 (N_13741,N_10388,N_12021);
and U13742 (N_13742,N_11906,N_11003);
and U13743 (N_13743,N_11636,N_10794);
or U13744 (N_13744,N_11933,N_10036);
or U13745 (N_13745,N_10352,N_12280);
or U13746 (N_13746,N_10538,N_10235);
and U13747 (N_13747,N_10477,N_12372);
or U13748 (N_13748,N_12136,N_11434);
and U13749 (N_13749,N_12265,N_11818);
nor U13750 (N_13750,N_11567,N_12110);
or U13751 (N_13751,N_11873,N_12284);
and U13752 (N_13752,N_11947,N_12404);
xnor U13753 (N_13753,N_10886,N_11815);
or U13754 (N_13754,N_11918,N_12082);
nor U13755 (N_13755,N_10998,N_10262);
nand U13756 (N_13756,N_12095,N_11336);
and U13757 (N_13757,N_11981,N_11788);
nor U13758 (N_13758,N_11058,N_11675);
nor U13759 (N_13759,N_10623,N_11896);
nor U13760 (N_13760,N_11253,N_10391);
and U13761 (N_13761,N_11514,N_11642);
nor U13762 (N_13762,N_12111,N_10343);
and U13763 (N_13763,N_11840,N_11816);
nand U13764 (N_13764,N_10348,N_11634);
nor U13765 (N_13765,N_12052,N_12259);
nand U13766 (N_13766,N_11727,N_10688);
and U13767 (N_13767,N_12296,N_10195);
nor U13768 (N_13768,N_10119,N_11627);
nand U13769 (N_13769,N_10344,N_12212);
and U13770 (N_13770,N_12052,N_11155);
or U13771 (N_13771,N_11933,N_11279);
or U13772 (N_13772,N_11777,N_12113);
and U13773 (N_13773,N_11052,N_11138);
or U13774 (N_13774,N_12324,N_11462);
or U13775 (N_13775,N_11182,N_10597);
and U13776 (N_13776,N_10330,N_10535);
nand U13777 (N_13777,N_11632,N_11450);
or U13778 (N_13778,N_11454,N_10529);
or U13779 (N_13779,N_11229,N_10723);
or U13780 (N_13780,N_10017,N_10451);
or U13781 (N_13781,N_10031,N_10821);
and U13782 (N_13782,N_11999,N_11430);
nand U13783 (N_13783,N_11802,N_11352);
and U13784 (N_13784,N_10835,N_10165);
or U13785 (N_13785,N_12027,N_10884);
or U13786 (N_13786,N_11981,N_11403);
and U13787 (N_13787,N_10328,N_10060);
nor U13788 (N_13788,N_11558,N_11017);
and U13789 (N_13789,N_11468,N_12346);
or U13790 (N_13790,N_11152,N_12290);
and U13791 (N_13791,N_12186,N_11660);
xnor U13792 (N_13792,N_10720,N_11078);
nand U13793 (N_13793,N_11485,N_10929);
nor U13794 (N_13794,N_10863,N_10673);
nand U13795 (N_13795,N_10299,N_12198);
or U13796 (N_13796,N_10683,N_10747);
and U13797 (N_13797,N_12067,N_12306);
xnor U13798 (N_13798,N_11111,N_10725);
nor U13799 (N_13799,N_11026,N_12127);
nand U13800 (N_13800,N_11611,N_11368);
nand U13801 (N_13801,N_10832,N_10139);
or U13802 (N_13802,N_11097,N_10962);
or U13803 (N_13803,N_11790,N_10456);
xor U13804 (N_13804,N_11157,N_11642);
xnor U13805 (N_13805,N_11649,N_12317);
or U13806 (N_13806,N_10754,N_12357);
and U13807 (N_13807,N_12026,N_10528);
or U13808 (N_13808,N_12015,N_11593);
xnor U13809 (N_13809,N_12302,N_11233);
and U13810 (N_13810,N_11672,N_10379);
and U13811 (N_13811,N_10824,N_10790);
nand U13812 (N_13812,N_10680,N_11423);
nor U13813 (N_13813,N_12006,N_11413);
or U13814 (N_13814,N_12485,N_11246);
nor U13815 (N_13815,N_10404,N_10300);
nor U13816 (N_13816,N_11062,N_10062);
nand U13817 (N_13817,N_10885,N_10937);
nor U13818 (N_13818,N_11975,N_10377);
or U13819 (N_13819,N_10844,N_10001);
or U13820 (N_13820,N_10542,N_11732);
nor U13821 (N_13821,N_12022,N_12233);
xnor U13822 (N_13822,N_12358,N_11365);
xor U13823 (N_13823,N_11718,N_11984);
nor U13824 (N_13824,N_11850,N_11433);
or U13825 (N_13825,N_10443,N_11312);
or U13826 (N_13826,N_10353,N_10605);
xor U13827 (N_13827,N_11229,N_11986);
xor U13828 (N_13828,N_11164,N_11200);
and U13829 (N_13829,N_11816,N_10839);
or U13830 (N_13830,N_12465,N_10791);
nor U13831 (N_13831,N_12467,N_11713);
or U13832 (N_13832,N_11306,N_10996);
nand U13833 (N_13833,N_11970,N_11704);
and U13834 (N_13834,N_12345,N_11480);
and U13835 (N_13835,N_10446,N_12098);
or U13836 (N_13836,N_12266,N_12341);
nand U13837 (N_13837,N_11832,N_12355);
and U13838 (N_13838,N_10673,N_10075);
nand U13839 (N_13839,N_12348,N_12235);
nand U13840 (N_13840,N_10495,N_12405);
xnor U13841 (N_13841,N_11388,N_10659);
and U13842 (N_13842,N_12115,N_11216);
nor U13843 (N_13843,N_10060,N_11361);
nor U13844 (N_13844,N_10039,N_10789);
nor U13845 (N_13845,N_11443,N_10146);
nor U13846 (N_13846,N_10192,N_10587);
nand U13847 (N_13847,N_11723,N_11657);
nor U13848 (N_13848,N_10404,N_12346);
nor U13849 (N_13849,N_11387,N_11153);
nor U13850 (N_13850,N_11015,N_10244);
nor U13851 (N_13851,N_11570,N_11187);
nor U13852 (N_13852,N_10948,N_10670);
or U13853 (N_13853,N_10425,N_12078);
nor U13854 (N_13854,N_11532,N_12217);
or U13855 (N_13855,N_11670,N_12149);
or U13856 (N_13856,N_11783,N_10129);
and U13857 (N_13857,N_10907,N_10846);
and U13858 (N_13858,N_10440,N_11871);
and U13859 (N_13859,N_10808,N_12075);
nand U13860 (N_13860,N_10396,N_11546);
and U13861 (N_13861,N_11043,N_12181);
nand U13862 (N_13862,N_11893,N_10924);
and U13863 (N_13863,N_11717,N_10891);
and U13864 (N_13864,N_10532,N_10677);
xnor U13865 (N_13865,N_10902,N_12396);
nand U13866 (N_13866,N_11448,N_10977);
or U13867 (N_13867,N_12104,N_10293);
nor U13868 (N_13868,N_11631,N_11936);
nor U13869 (N_13869,N_11547,N_11715);
or U13870 (N_13870,N_10226,N_12153);
nand U13871 (N_13871,N_10110,N_12313);
and U13872 (N_13872,N_10306,N_11586);
nor U13873 (N_13873,N_11300,N_11982);
xnor U13874 (N_13874,N_11266,N_12431);
and U13875 (N_13875,N_11612,N_11546);
nor U13876 (N_13876,N_10511,N_10564);
xnor U13877 (N_13877,N_11828,N_11186);
nor U13878 (N_13878,N_12439,N_10091);
nor U13879 (N_13879,N_11352,N_11628);
and U13880 (N_13880,N_12188,N_11307);
and U13881 (N_13881,N_11161,N_10615);
xnor U13882 (N_13882,N_11489,N_11443);
nor U13883 (N_13883,N_11430,N_12227);
nand U13884 (N_13884,N_12350,N_10544);
xor U13885 (N_13885,N_12280,N_11673);
nor U13886 (N_13886,N_12352,N_10451);
nor U13887 (N_13887,N_12214,N_10526);
nor U13888 (N_13888,N_11388,N_10677);
nor U13889 (N_13889,N_12206,N_11441);
nor U13890 (N_13890,N_11155,N_12350);
nor U13891 (N_13891,N_11299,N_11801);
nand U13892 (N_13892,N_11252,N_11371);
nor U13893 (N_13893,N_11915,N_12154);
nand U13894 (N_13894,N_11273,N_11186);
and U13895 (N_13895,N_11909,N_12346);
xor U13896 (N_13896,N_12042,N_10475);
xor U13897 (N_13897,N_10518,N_10375);
nand U13898 (N_13898,N_12485,N_11579);
and U13899 (N_13899,N_11163,N_11849);
nor U13900 (N_13900,N_10760,N_11085);
or U13901 (N_13901,N_10213,N_11451);
nand U13902 (N_13902,N_11131,N_11697);
nor U13903 (N_13903,N_12393,N_12057);
and U13904 (N_13904,N_10936,N_10511);
nand U13905 (N_13905,N_12243,N_12422);
nand U13906 (N_13906,N_10525,N_10617);
nand U13907 (N_13907,N_10624,N_12004);
and U13908 (N_13908,N_10071,N_10950);
nand U13909 (N_13909,N_10642,N_11845);
nand U13910 (N_13910,N_10481,N_11607);
or U13911 (N_13911,N_10558,N_11077);
nand U13912 (N_13912,N_12020,N_12072);
nand U13913 (N_13913,N_11347,N_10167);
nand U13914 (N_13914,N_10587,N_11010);
nor U13915 (N_13915,N_11644,N_10333);
and U13916 (N_13916,N_10808,N_10535);
and U13917 (N_13917,N_10254,N_10065);
nand U13918 (N_13918,N_10126,N_10598);
or U13919 (N_13919,N_12185,N_11083);
nand U13920 (N_13920,N_12346,N_11961);
nor U13921 (N_13921,N_11516,N_10343);
and U13922 (N_13922,N_11895,N_10025);
xnor U13923 (N_13923,N_11054,N_10378);
and U13924 (N_13924,N_12325,N_10595);
or U13925 (N_13925,N_10543,N_10626);
or U13926 (N_13926,N_12180,N_12231);
or U13927 (N_13927,N_10253,N_10358);
nor U13928 (N_13928,N_12176,N_11031);
or U13929 (N_13929,N_12256,N_12303);
or U13930 (N_13930,N_11485,N_10483);
nor U13931 (N_13931,N_10076,N_11282);
nand U13932 (N_13932,N_12304,N_11018);
nand U13933 (N_13933,N_10679,N_10045);
nor U13934 (N_13934,N_10773,N_11052);
and U13935 (N_13935,N_10884,N_11448);
and U13936 (N_13936,N_10015,N_10274);
or U13937 (N_13937,N_10718,N_10855);
nand U13938 (N_13938,N_12068,N_10283);
nor U13939 (N_13939,N_11722,N_12206);
and U13940 (N_13940,N_10165,N_10620);
and U13941 (N_13941,N_10192,N_10099);
or U13942 (N_13942,N_12168,N_11104);
or U13943 (N_13943,N_11414,N_11694);
and U13944 (N_13944,N_10228,N_10984);
and U13945 (N_13945,N_10737,N_10314);
nor U13946 (N_13946,N_10636,N_11627);
nor U13947 (N_13947,N_12172,N_11874);
nor U13948 (N_13948,N_10642,N_11549);
and U13949 (N_13949,N_10578,N_11880);
or U13950 (N_13950,N_10486,N_10681);
nand U13951 (N_13951,N_10089,N_11939);
nand U13952 (N_13952,N_10046,N_11268);
nand U13953 (N_13953,N_11454,N_12493);
nand U13954 (N_13954,N_10309,N_12468);
nor U13955 (N_13955,N_11925,N_10995);
or U13956 (N_13956,N_12083,N_10890);
and U13957 (N_13957,N_11320,N_10323);
nand U13958 (N_13958,N_11669,N_10268);
or U13959 (N_13959,N_10219,N_10560);
and U13960 (N_13960,N_11041,N_11323);
or U13961 (N_13961,N_12379,N_10997);
nor U13962 (N_13962,N_10637,N_12115);
nand U13963 (N_13963,N_10900,N_11817);
nor U13964 (N_13964,N_10323,N_10269);
nand U13965 (N_13965,N_10780,N_10379);
nand U13966 (N_13966,N_11744,N_11090);
nor U13967 (N_13967,N_11475,N_11550);
and U13968 (N_13968,N_10495,N_11685);
nand U13969 (N_13969,N_12441,N_11237);
xor U13970 (N_13970,N_11552,N_11806);
nor U13971 (N_13971,N_10024,N_10769);
or U13972 (N_13972,N_11842,N_10081);
nand U13973 (N_13973,N_12140,N_12341);
and U13974 (N_13974,N_10402,N_12273);
nor U13975 (N_13975,N_10224,N_10300);
and U13976 (N_13976,N_12488,N_12101);
and U13977 (N_13977,N_12273,N_11162);
nor U13978 (N_13978,N_11249,N_10513);
nand U13979 (N_13979,N_11081,N_10019);
nand U13980 (N_13980,N_10986,N_10036);
xnor U13981 (N_13981,N_10962,N_10025);
nand U13982 (N_13982,N_11277,N_12192);
nand U13983 (N_13983,N_10783,N_10014);
or U13984 (N_13984,N_11394,N_10507);
nand U13985 (N_13985,N_10588,N_10070);
nand U13986 (N_13986,N_12400,N_10142);
xor U13987 (N_13987,N_11844,N_12253);
nor U13988 (N_13988,N_11545,N_11863);
nand U13989 (N_13989,N_10684,N_10857);
nor U13990 (N_13990,N_12226,N_10893);
or U13991 (N_13991,N_11407,N_10654);
nor U13992 (N_13992,N_10835,N_10095);
or U13993 (N_13993,N_10980,N_12137);
and U13994 (N_13994,N_11435,N_11763);
and U13995 (N_13995,N_11067,N_11561);
nand U13996 (N_13996,N_11090,N_11660);
xnor U13997 (N_13997,N_10509,N_11468);
nand U13998 (N_13998,N_10824,N_10604);
or U13999 (N_13999,N_12023,N_10935);
nor U14000 (N_14000,N_10226,N_11139);
and U14001 (N_14001,N_11703,N_11773);
xor U14002 (N_14002,N_11890,N_10574);
nor U14003 (N_14003,N_10189,N_11907);
or U14004 (N_14004,N_11163,N_10595);
nor U14005 (N_14005,N_10221,N_10003);
nand U14006 (N_14006,N_10682,N_12031);
nor U14007 (N_14007,N_12142,N_12016);
xnor U14008 (N_14008,N_12491,N_11317);
and U14009 (N_14009,N_10575,N_10892);
xnor U14010 (N_14010,N_10923,N_10510);
or U14011 (N_14011,N_10375,N_10114);
xor U14012 (N_14012,N_11062,N_10695);
and U14013 (N_14013,N_12243,N_11067);
nand U14014 (N_14014,N_11792,N_10113);
nor U14015 (N_14015,N_12439,N_12168);
nor U14016 (N_14016,N_11522,N_10420);
and U14017 (N_14017,N_11654,N_10385);
xnor U14018 (N_14018,N_11930,N_10581);
and U14019 (N_14019,N_10251,N_10174);
nand U14020 (N_14020,N_11890,N_11388);
and U14021 (N_14021,N_12270,N_11849);
nand U14022 (N_14022,N_11436,N_12479);
xor U14023 (N_14023,N_10904,N_10680);
or U14024 (N_14024,N_11345,N_10935);
or U14025 (N_14025,N_11139,N_11764);
and U14026 (N_14026,N_10258,N_10488);
nor U14027 (N_14027,N_12457,N_10469);
or U14028 (N_14028,N_11132,N_10218);
nor U14029 (N_14029,N_11687,N_12385);
nand U14030 (N_14030,N_10856,N_11948);
or U14031 (N_14031,N_12095,N_10938);
xnor U14032 (N_14032,N_11879,N_12058);
and U14033 (N_14033,N_11463,N_10385);
and U14034 (N_14034,N_11714,N_12266);
and U14035 (N_14035,N_12004,N_11514);
nor U14036 (N_14036,N_10249,N_10444);
nor U14037 (N_14037,N_10997,N_10420);
and U14038 (N_14038,N_11000,N_11099);
nand U14039 (N_14039,N_10971,N_12268);
and U14040 (N_14040,N_11712,N_11604);
or U14041 (N_14041,N_11115,N_11890);
and U14042 (N_14042,N_11105,N_12141);
nor U14043 (N_14043,N_11549,N_10858);
nor U14044 (N_14044,N_10390,N_11961);
or U14045 (N_14045,N_10154,N_10632);
and U14046 (N_14046,N_12402,N_11520);
nand U14047 (N_14047,N_11537,N_10214);
nor U14048 (N_14048,N_11200,N_12484);
nor U14049 (N_14049,N_10301,N_10409);
xor U14050 (N_14050,N_11677,N_10849);
or U14051 (N_14051,N_10312,N_10167);
or U14052 (N_14052,N_10114,N_12265);
and U14053 (N_14053,N_11621,N_12266);
xor U14054 (N_14054,N_10248,N_10218);
nand U14055 (N_14055,N_12281,N_11416);
nor U14056 (N_14056,N_10449,N_12419);
and U14057 (N_14057,N_10137,N_11223);
or U14058 (N_14058,N_10436,N_10028);
nand U14059 (N_14059,N_11742,N_11263);
or U14060 (N_14060,N_10018,N_10612);
nand U14061 (N_14061,N_10188,N_10696);
nor U14062 (N_14062,N_10801,N_10687);
and U14063 (N_14063,N_12379,N_11888);
and U14064 (N_14064,N_11304,N_12486);
nand U14065 (N_14065,N_10519,N_12213);
and U14066 (N_14066,N_12306,N_10428);
nor U14067 (N_14067,N_11577,N_10504);
xnor U14068 (N_14068,N_10584,N_10856);
and U14069 (N_14069,N_10119,N_11181);
nor U14070 (N_14070,N_10558,N_11496);
nor U14071 (N_14071,N_10572,N_10626);
or U14072 (N_14072,N_11104,N_12236);
or U14073 (N_14073,N_10880,N_11804);
nand U14074 (N_14074,N_12489,N_11169);
or U14075 (N_14075,N_10789,N_10332);
nand U14076 (N_14076,N_11655,N_11882);
nand U14077 (N_14077,N_11330,N_12278);
nor U14078 (N_14078,N_10161,N_10875);
and U14079 (N_14079,N_10685,N_12419);
nand U14080 (N_14080,N_11268,N_10185);
or U14081 (N_14081,N_10158,N_10970);
or U14082 (N_14082,N_11314,N_12114);
and U14083 (N_14083,N_11329,N_10393);
or U14084 (N_14084,N_12014,N_11519);
nor U14085 (N_14085,N_10948,N_11369);
nand U14086 (N_14086,N_10936,N_12206);
or U14087 (N_14087,N_11059,N_10325);
or U14088 (N_14088,N_10495,N_10933);
nor U14089 (N_14089,N_10453,N_10530);
nor U14090 (N_14090,N_10278,N_11645);
or U14091 (N_14091,N_10364,N_10255);
xnor U14092 (N_14092,N_12151,N_10760);
nand U14093 (N_14093,N_11783,N_11549);
or U14094 (N_14094,N_10997,N_11060);
nor U14095 (N_14095,N_11778,N_10823);
xnor U14096 (N_14096,N_10410,N_11992);
or U14097 (N_14097,N_12404,N_10141);
nand U14098 (N_14098,N_12287,N_10876);
nor U14099 (N_14099,N_10030,N_10844);
nand U14100 (N_14100,N_10072,N_12398);
nor U14101 (N_14101,N_10756,N_10419);
nor U14102 (N_14102,N_11752,N_11317);
and U14103 (N_14103,N_10631,N_11063);
nor U14104 (N_14104,N_11226,N_10303);
nor U14105 (N_14105,N_12245,N_12183);
or U14106 (N_14106,N_12367,N_11967);
nor U14107 (N_14107,N_10862,N_10304);
nor U14108 (N_14108,N_12190,N_10272);
and U14109 (N_14109,N_12275,N_12392);
nand U14110 (N_14110,N_11022,N_12494);
or U14111 (N_14111,N_12110,N_12452);
nand U14112 (N_14112,N_12291,N_12476);
nor U14113 (N_14113,N_11601,N_11580);
and U14114 (N_14114,N_10098,N_12095);
and U14115 (N_14115,N_12403,N_12231);
and U14116 (N_14116,N_10257,N_11587);
or U14117 (N_14117,N_11576,N_11979);
nor U14118 (N_14118,N_10422,N_11110);
nand U14119 (N_14119,N_10638,N_11977);
nand U14120 (N_14120,N_10236,N_12064);
or U14121 (N_14121,N_11762,N_10335);
or U14122 (N_14122,N_11846,N_11159);
nand U14123 (N_14123,N_10970,N_12028);
xor U14124 (N_14124,N_11808,N_12354);
nor U14125 (N_14125,N_11567,N_11964);
or U14126 (N_14126,N_10315,N_11558);
nor U14127 (N_14127,N_11195,N_11326);
and U14128 (N_14128,N_11053,N_11759);
or U14129 (N_14129,N_10585,N_10896);
nand U14130 (N_14130,N_11080,N_11532);
nor U14131 (N_14131,N_11669,N_10634);
and U14132 (N_14132,N_11571,N_12447);
nand U14133 (N_14133,N_10802,N_11625);
and U14134 (N_14134,N_10459,N_11068);
nand U14135 (N_14135,N_11393,N_11022);
nor U14136 (N_14136,N_11948,N_10016);
or U14137 (N_14137,N_11519,N_10230);
and U14138 (N_14138,N_10866,N_12422);
nor U14139 (N_14139,N_10265,N_11595);
nor U14140 (N_14140,N_10101,N_10585);
and U14141 (N_14141,N_10406,N_10109);
or U14142 (N_14142,N_11824,N_10036);
nand U14143 (N_14143,N_10315,N_12134);
nor U14144 (N_14144,N_10885,N_10200);
and U14145 (N_14145,N_10341,N_12469);
xnor U14146 (N_14146,N_11535,N_12091);
nor U14147 (N_14147,N_11303,N_11451);
or U14148 (N_14148,N_12467,N_12461);
nor U14149 (N_14149,N_10404,N_11485);
nand U14150 (N_14150,N_11960,N_11431);
nand U14151 (N_14151,N_12314,N_11001);
or U14152 (N_14152,N_11848,N_11295);
and U14153 (N_14153,N_11788,N_10349);
and U14154 (N_14154,N_10409,N_12384);
and U14155 (N_14155,N_12268,N_12344);
nand U14156 (N_14156,N_11878,N_10450);
xor U14157 (N_14157,N_11132,N_12478);
and U14158 (N_14158,N_10159,N_10289);
nand U14159 (N_14159,N_12168,N_11070);
xor U14160 (N_14160,N_11520,N_11301);
or U14161 (N_14161,N_11937,N_11775);
or U14162 (N_14162,N_12288,N_12092);
and U14163 (N_14163,N_12390,N_11024);
xnor U14164 (N_14164,N_11897,N_11795);
or U14165 (N_14165,N_12188,N_11865);
or U14166 (N_14166,N_11527,N_12087);
nand U14167 (N_14167,N_10127,N_11187);
nand U14168 (N_14168,N_12008,N_11709);
and U14169 (N_14169,N_11363,N_11665);
nor U14170 (N_14170,N_11623,N_10318);
nor U14171 (N_14171,N_11643,N_11003);
or U14172 (N_14172,N_11485,N_11762);
and U14173 (N_14173,N_11510,N_11699);
or U14174 (N_14174,N_10385,N_10615);
and U14175 (N_14175,N_10537,N_11599);
nor U14176 (N_14176,N_11220,N_12051);
nand U14177 (N_14177,N_10371,N_10949);
nand U14178 (N_14178,N_10755,N_11215);
nand U14179 (N_14179,N_12484,N_10212);
and U14180 (N_14180,N_11093,N_11701);
nor U14181 (N_14181,N_11905,N_11443);
or U14182 (N_14182,N_11638,N_11144);
nor U14183 (N_14183,N_11019,N_11235);
and U14184 (N_14184,N_10205,N_11086);
or U14185 (N_14185,N_11758,N_10607);
nor U14186 (N_14186,N_12412,N_10563);
or U14187 (N_14187,N_10050,N_11079);
or U14188 (N_14188,N_12088,N_11724);
xor U14189 (N_14189,N_10264,N_11804);
nand U14190 (N_14190,N_10884,N_11648);
nand U14191 (N_14191,N_10792,N_11653);
or U14192 (N_14192,N_10081,N_12442);
and U14193 (N_14193,N_11980,N_11900);
nand U14194 (N_14194,N_11026,N_11921);
or U14195 (N_14195,N_10306,N_10517);
nor U14196 (N_14196,N_11116,N_12343);
and U14197 (N_14197,N_10528,N_12164);
and U14198 (N_14198,N_12175,N_11555);
and U14199 (N_14199,N_10869,N_11422);
xnor U14200 (N_14200,N_12360,N_11363);
xor U14201 (N_14201,N_10005,N_11993);
or U14202 (N_14202,N_10059,N_12360);
and U14203 (N_14203,N_12058,N_12386);
nor U14204 (N_14204,N_11109,N_10417);
nand U14205 (N_14205,N_10773,N_10740);
nand U14206 (N_14206,N_11586,N_10163);
and U14207 (N_14207,N_11949,N_11294);
and U14208 (N_14208,N_10247,N_11616);
nand U14209 (N_14209,N_12176,N_10153);
xnor U14210 (N_14210,N_11089,N_11336);
nor U14211 (N_14211,N_11557,N_11628);
or U14212 (N_14212,N_11455,N_10613);
nand U14213 (N_14213,N_11336,N_10168);
or U14214 (N_14214,N_10843,N_10230);
or U14215 (N_14215,N_11555,N_11638);
xor U14216 (N_14216,N_10190,N_10324);
nand U14217 (N_14217,N_11866,N_10127);
or U14218 (N_14218,N_11250,N_12096);
nand U14219 (N_14219,N_12496,N_10683);
and U14220 (N_14220,N_11963,N_12410);
or U14221 (N_14221,N_12370,N_11905);
or U14222 (N_14222,N_11922,N_11147);
nand U14223 (N_14223,N_10767,N_11471);
nor U14224 (N_14224,N_12209,N_11046);
and U14225 (N_14225,N_11927,N_10366);
xor U14226 (N_14226,N_11847,N_10786);
nor U14227 (N_14227,N_10180,N_11322);
or U14228 (N_14228,N_10289,N_12004);
xnor U14229 (N_14229,N_10565,N_12184);
nand U14230 (N_14230,N_11153,N_12372);
nor U14231 (N_14231,N_12393,N_12251);
xnor U14232 (N_14232,N_11523,N_11642);
nor U14233 (N_14233,N_11797,N_10632);
nor U14234 (N_14234,N_12448,N_10610);
nand U14235 (N_14235,N_11493,N_10484);
or U14236 (N_14236,N_12246,N_10497);
xnor U14237 (N_14237,N_11151,N_10951);
nor U14238 (N_14238,N_10462,N_11721);
nand U14239 (N_14239,N_10170,N_10969);
nor U14240 (N_14240,N_10882,N_10374);
and U14241 (N_14241,N_10162,N_10572);
and U14242 (N_14242,N_12187,N_10174);
and U14243 (N_14243,N_10204,N_10007);
nor U14244 (N_14244,N_11408,N_10534);
and U14245 (N_14245,N_10379,N_10535);
nor U14246 (N_14246,N_11156,N_12281);
nor U14247 (N_14247,N_12028,N_10789);
nand U14248 (N_14248,N_10757,N_10529);
or U14249 (N_14249,N_10748,N_11785);
or U14250 (N_14250,N_10138,N_11467);
nor U14251 (N_14251,N_12346,N_11802);
nand U14252 (N_14252,N_10536,N_11275);
or U14253 (N_14253,N_10083,N_10335);
and U14254 (N_14254,N_11950,N_12247);
or U14255 (N_14255,N_11533,N_10119);
and U14256 (N_14256,N_10462,N_10417);
xor U14257 (N_14257,N_10194,N_11511);
or U14258 (N_14258,N_11105,N_12168);
or U14259 (N_14259,N_10183,N_10822);
xnor U14260 (N_14260,N_11073,N_11083);
nor U14261 (N_14261,N_10699,N_11030);
and U14262 (N_14262,N_10799,N_10995);
nor U14263 (N_14263,N_11956,N_10531);
and U14264 (N_14264,N_11605,N_11871);
nor U14265 (N_14265,N_10704,N_10780);
nor U14266 (N_14266,N_10789,N_12039);
nand U14267 (N_14267,N_10631,N_11380);
and U14268 (N_14268,N_12466,N_10509);
nand U14269 (N_14269,N_11890,N_10061);
or U14270 (N_14270,N_12311,N_10040);
nor U14271 (N_14271,N_11290,N_12469);
nor U14272 (N_14272,N_11988,N_12200);
nor U14273 (N_14273,N_11653,N_11414);
nand U14274 (N_14274,N_10059,N_10930);
or U14275 (N_14275,N_10705,N_11976);
and U14276 (N_14276,N_11200,N_10937);
nand U14277 (N_14277,N_11781,N_10319);
nor U14278 (N_14278,N_12435,N_11830);
nor U14279 (N_14279,N_11111,N_12151);
nor U14280 (N_14280,N_10946,N_11412);
nand U14281 (N_14281,N_10213,N_10860);
or U14282 (N_14282,N_12098,N_11466);
and U14283 (N_14283,N_12011,N_11351);
or U14284 (N_14284,N_11538,N_10511);
and U14285 (N_14285,N_10756,N_10758);
nor U14286 (N_14286,N_10395,N_10615);
nand U14287 (N_14287,N_11607,N_10249);
xor U14288 (N_14288,N_12147,N_10977);
nor U14289 (N_14289,N_10890,N_11370);
nor U14290 (N_14290,N_11652,N_12390);
xor U14291 (N_14291,N_11338,N_12165);
nand U14292 (N_14292,N_10922,N_11055);
nand U14293 (N_14293,N_10230,N_11931);
or U14294 (N_14294,N_11746,N_11383);
nor U14295 (N_14295,N_11094,N_10222);
nand U14296 (N_14296,N_10129,N_10636);
xnor U14297 (N_14297,N_11282,N_10038);
or U14298 (N_14298,N_10351,N_10810);
xnor U14299 (N_14299,N_10911,N_11779);
nor U14300 (N_14300,N_11690,N_12467);
and U14301 (N_14301,N_11552,N_11746);
nand U14302 (N_14302,N_12105,N_10580);
and U14303 (N_14303,N_10480,N_11126);
nand U14304 (N_14304,N_10950,N_11869);
nor U14305 (N_14305,N_11891,N_10135);
nor U14306 (N_14306,N_11457,N_11102);
or U14307 (N_14307,N_10547,N_11368);
nand U14308 (N_14308,N_10097,N_10646);
nor U14309 (N_14309,N_12382,N_10898);
nand U14310 (N_14310,N_10465,N_11317);
nand U14311 (N_14311,N_10317,N_10719);
nor U14312 (N_14312,N_11541,N_12439);
or U14313 (N_14313,N_12121,N_11348);
and U14314 (N_14314,N_10736,N_11368);
nor U14315 (N_14315,N_11941,N_10019);
and U14316 (N_14316,N_10225,N_10160);
nor U14317 (N_14317,N_10038,N_10508);
nand U14318 (N_14318,N_11255,N_10382);
and U14319 (N_14319,N_10131,N_12321);
nor U14320 (N_14320,N_12450,N_11552);
nor U14321 (N_14321,N_11008,N_12203);
and U14322 (N_14322,N_10457,N_11164);
or U14323 (N_14323,N_11707,N_11143);
nor U14324 (N_14324,N_10883,N_10798);
or U14325 (N_14325,N_11833,N_11209);
nor U14326 (N_14326,N_10057,N_11687);
nand U14327 (N_14327,N_11998,N_10279);
nor U14328 (N_14328,N_10643,N_11304);
or U14329 (N_14329,N_10884,N_11632);
nand U14330 (N_14330,N_10073,N_11758);
and U14331 (N_14331,N_11261,N_11820);
and U14332 (N_14332,N_11172,N_10621);
nand U14333 (N_14333,N_11952,N_10123);
nand U14334 (N_14334,N_10955,N_10180);
or U14335 (N_14335,N_10360,N_11367);
or U14336 (N_14336,N_10928,N_10180);
nor U14337 (N_14337,N_11345,N_10445);
or U14338 (N_14338,N_11989,N_11646);
nand U14339 (N_14339,N_11699,N_11658);
nor U14340 (N_14340,N_11997,N_10463);
or U14341 (N_14341,N_12307,N_10198);
nand U14342 (N_14342,N_11621,N_11782);
nor U14343 (N_14343,N_10658,N_12274);
nor U14344 (N_14344,N_10738,N_12489);
and U14345 (N_14345,N_10597,N_12121);
xnor U14346 (N_14346,N_10509,N_11409);
and U14347 (N_14347,N_11445,N_11140);
and U14348 (N_14348,N_12078,N_11591);
nand U14349 (N_14349,N_12075,N_12400);
xnor U14350 (N_14350,N_10914,N_10227);
and U14351 (N_14351,N_10568,N_11983);
xor U14352 (N_14352,N_10618,N_10950);
xor U14353 (N_14353,N_11204,N_12057);
nor U14354 (N_14354,N_12132,N_11494);
nand U14355 (N_14355,N_11396,N_11787);
and U14356 (N_14356,N_12231,N_10339);
nor U14357 (N_14357,N_10459,N_10735);
nand U14358 (N_14358,N_10643,N_10005);
xor U14359 (N_14359,N_10050,N_11444);
and U14360 (N_14360,N_11417,N_11227);
or U14361 (N_14361,N_12233,N_10583);
nor U14362 (N_14362,N_11380,N_10366);
nand U14363 (N_14363,N_10188,N_11056);
or U14364 (N_14364,N_11598,N_10156);
nand U14365 (N_14365,N_11712,N_10091);
and U14366 (N_14366,N_10676,N_10738);
nor U14367 (N_14367,N_11601,N_10448);
nor U14368 (N_14368,N_11837,N_10308);
nand U14369 (N_14369,N_11942,N_12061);
xor U14370 (N_14370,N_11244,N_11794);
nand U14371 (N_14371,N_12490,N_12187);
and U14372 (N_14372,N_11567,N_11661);
and U14373 (N_14373,N_11369,N_11551);
nor U14374 (N_14374,N_10975,N_12189);
nor U14375 (N_14375,N_12103,N_10664);
or U14376 (N_14376,N_11475,N_11627);
and U14377 (N_14377,N_11647,N_11494);
and U14378 (N_14378,N_11538,N_10604);
nor U14379 (N_14379,N_10973,N_10272);
nor U14380 (N_14380,N_11387,N_10393);
nand U14381 (N_14381,N_11886,N_12020);
xor U14382 (N_14382,N_11699,N_10951);
or U14383 (N_14383,N_11643,N_11312);
nor U14384 (N_14384,N_12052,N_12119);
nor U14385 (N_14385,N_11512,N_10397);
or U14386 (N_14386,N_11382,N_10857);
nand U14387 (N_14387,N_10825,N_10633);
or U14388 (N_14388,N_10470,N_10827);
nor U14389 (N_14389,N_11387,N_10985);
nor U14390 (N_14390,N_10335,N_12379);
or U14391 (N_14391,N_10775,N_10086);
or U14392 (N_14392,N_11027,N_11374);
nand U14393 (N_14393,N_10028,N_10086);
nand U14394 (N_14394,N_12265,N_10638);
nand U14395 (N_14395,N_10196,N_11218);
and U14396 (N_14396,N_10122,N_12182);
or U14397 (N_14397,N_11010,N_12366);
and U14398 (N_14398,N_10816,N_10421);
nor U14399 (N_14399,N_10627,N_10972);
or U14400 (N_14400,N_10142,N_11107);
and U14401 (N_14401,N_10564,N_11884);
nor U14402 (N_14402,N_10481,N_11784);
or U14403 (N_14403,N_10150,N_10842);
and U14404 (N_14404,N_11945,N_11487);
and U14405 (N_14405,N_12468,N_12288);
nand U14406 (N_14406,N_11394,N_10404);
nor U14407 (N_14407,N_11521,N_12174);
nand U14408 (N_14408,N_10191,N_11825);
and U14409 (N_14409,N_12130,N_10142);
and U14410 (N_14410,N_10364,N_11225);
nand U14411 (N_14411,N_11856,N_11529);
or U14412 (N_14412,N_10014,N_11912);
nor U14413 (N_14413,N_11846,N_10902);
nor U14414 (N_14414,N_10941,N_12062);
nand U14415 (N_14415,N_10413,N_11302);
xor U14416 (N_14416,N_10967,N_10493);
nand U14417 (N_14417,N_10360,N_12484);
nand U14418 (N_14418,N_11917,N_12037);
or U14419 (N_14419,N_11251,N_11283);
and U14420 (N_14420,N_10071,N_11334);
xnor U14421 (N_14421,N_10532,N_11494);
nor U14422 (N_14422,N_10436,N_12260);
and U14423 (N_14423,N_10382,N_11378);
or U14424 (N_14424,N_10273,N_11159);
xor U14425 (N_14425,N_12420,N_10503);
nand U14426 (N_14426,N_11710,N_10613);
or U14427 (N_14427,N_11220,N_11913);
or U14428 (N_14428,N_12180,N_11846);
nand U14429 (N_14429,N_10088,N_10530);
or U14430 (N_14430,N_12266,N_12466);
nand U14431 (N_14431,N_12461,N_12074);
nand U14432 (N_14432,N_10213,N_10701);
and U14433 (N_14433,N_10592,N_10565);
nor U14434 (N_14434,N_11185,N_10561);
and U14435 (N_14435,N_10250,N_10874);
nor U14436 (N_14436,N_11282,N_10747);
or U14437 (N_14437,N_11741,N_10248);
nor U14438 (N_14438,N_10632,N_12011);
or U14439 (N_14439,N_12462,N_12441);
and U14440 (N_14440,N_11275,N_12234);
or U14441 (N_14441,N_11916,N_10913);
nor U14442 (N_14442,N_11589,N_10563);
xor U14443 (N_14443,N_10089,N_11591);
xor U14444 (N_14444,N_11393,N_10061);
nand U14445 (N_14445,N_10041,N_10756);
nand U14446 (N_14446,N_10581,N_11799);
nand U14447 (N_14447,N_11534,N_10606);
and U14448 (N_14448,N_11360,N_10393);
xnor U14449 (N_14449,N_11713,N_11174);
xor U14450 (N_14450,N_10355,N_11860);
or U14451 (N_14451,N_10314,N_12041);
and U14452 (N_14452,N_10568,N_10266);
nand U14453 (N_14453,N_10242,N_11284);
or U14454 (N_14454,N_10853,N_11589);
or U14455 (N_14455,N_12315,N_11029);
nor U14456 (N_14456,N_11740,N_12098);
or U14457 (N_14457,N_11739,N_10926);
or U14458 (N_14458,N_11308,N_11312);
or U14459 (N_14459,N_10118,N_11024);
nor U14460 (N_14460,N_10071,N_10182);
and U14461 (N_14461,N_10213,N_10781);
and U14462 (N_14462,N_12441,N_11463);
or U14463 (N_14463,N_10701,N_12486);
and U14464 (N_14464,N_11605,N_10508);
nand U14465 (N_14465,N_10637,N_12022);
nor U14466 (N_14466,N_12447,N_10664);
and U14467 (N_14467,N_10121,N_10581);
nor U14468 (N_14468,N_11580,N_10500);
nand U14469 (N_14469,N_11677,N_12276);
or U14470 (N_14470,N_12161,N_10900);
xnor U14471 (N_14471,N_11294,N_11342);
and U14472 (N_14472,N_10955,N_11384);
nand U14473 (N_14473,N_12351,N_11745);
and U14474 (N_14474,N_11546,N_12327);
and U14475 (N_14475,N_12353,N_12483);
and U14476 (N_14476,N_10760,N_10610);
nand U14477 (N_14477,N_11346,N_10881);
nand U14478 (N_14478,N_12179,N_12113);
or U14479 (N_14479,N_11183,N_11192);
and U14480 (N_14480,N_11278,N_10034);
and U14481 (N_14481,N_12157,N_12418);
xor U14482 (N_14482,N_10158,N_10780);
or U14483 (N_14483,N_12029,N_11649);
nand U14484 (N_14484,N_11393,N_11844);
nor U14485 (N_14485,N_11857,N_11453);
nand U14486 (N_14486,N_11252,N_11126);
or U14487 (N_14487,N_10060,N_10346);
nor U14488 (N_14488,N_11408,N_10282);
nor U14489 (N_14489,N_12157,N_10627);
xnor U14490 (N_14490,N_10361,N_10883);
nand U14491 (N_14491,N_10071,N_11082);
or U14492 (N_14492,N_11411,N_12285);
and U14493 (N_14493,N_10497,N_12220);
nand U14494 (N_14494,N_11555,N_10769);
and U14495 (N_14495,N_12280,N_10068);
or U14496 (N_14496,N_11901,N_10063);
and U14497 (N_14497,N_11284,N_11905);
and U14498 (N_14498,N_11491,N_10848);
or U14499 (N_14499,N_10931,N_11924);
nand U14500 (N_14500,N_10569,N_10804);
nor U14501 (N_14501,N_11136,N_10301);
and U14502 (N_14502,N_11146,N_11747);
xnor U14503 (N_14503,N_11283,N_11806);
nor U14504 (N_14504,N_10250,N_11229);
nand U14505 (N_14505,N_11544,N_10609);
or U14506 (N_14506,N_11518,N_10955);
or U14507 (N_14507,N_10917,N_10385);
nand U14508 (N_14508,N_10417,N_12223);
nor U14509 (N_14509,N_11956,N_11042);
nor U14510 (N_14510,N_11753,N_12139);
xnor U14511 (N_14511,N_10268,N_10551);
nand U14512 (N_14512,N_10866,N_10645);
nand U14513 (N_14513,N_10707,N_11542);
nand U14514 (N_14514,N_10558,N_10414);
or U14515 (N_14515,N_10532,N_11164);
xor U14516 (N_14516,N_12404,N_10433);
and U14517 (N_14517,N_12158,N_11839);
nand U14518 (N_14518,N_11247,N_10961);
or U14519 (N_14519,N_12210,N_11341);
nand U14520 (N_14520,N_10272,N_12146);
or U14521 (N_14521,N_12353,N_11704);
nor U14522 (N_14522,N_12276,N_10701);
and U14523 (N_14523,N_10080,N_11846);
nand U14524 (N_14524,N_11606,N_11664);
or U14525 (N_14525,N_12015,N_10801);
xnor U14526 (N_14526,N_11084,N_10894);
nand U14527 (N_14527,N_10988,N_12392);
nor U14528 (N_14528,N_10587,N_11751);
nand U14529 (N_14529,N_12130,N_12081);
xnor U14530 (N_14530,N_11755,N_10755);
and U14531 (N_14531,N_10163,N_11889);
or U14532 (N_14532,N_11267,N_10785);
and U14533 (N_14533,N_11671,N_11451);
xor U14534 (N_14534,N_11753,N_12375);
xnor U14535 (N_14535,N_11692,N_11888);
nand U14536 (N_14536,N_11632,N_11394);
xnor U14537 (N_14537,N_10372,N_10917);
and U14538 (N_14538,N_12222,N_10851);
xnor U14539 (N_14539,N_12130,N_12014);
nand U14540 (N_14540,N_11490,N_10086);
nor U14541 (N_14541,N_10660,N_10015);
nor U14542 (N_14542,N_10917,N_11039);
or U14543 (N_14543,N_12176,N_11318);
and U14544 (N_14544,N_10496,N_11695);
nor U14545 (N_14545,N_10919,N_11395);
nand U14546 (N_14546,N_10684,N_10614);
and U14547 (N_14547,N_10431,N_10746);
nand U14548 (N_14548,N_10514,N_11013);
nand U14549 (N_14549,N_10065,N_11752);
or U14550 (N_14550,N_11958,N_11862);
or U14551 (N_14551,N_12158,N_11112);
nor U14552 (N_14552,N_10241,N_12068);
or U14553 (N_14553,N_11799,N_11224);
nand U14554 (N_14554,N_11040,N_10369);
xor U14555 (N_14555,N_10334,N_10983);
and U14556 (N_14556,N_12278,N_11711);
nor U14557 (N_14557,N_11502,N_11081);
nand U14558 (N_14558,N_11375,N_11310);
nor U14559 (N_14559,N_11385,N_10086);
nand U14560 (N_14560,N_12207,N_11393);
or U14561 (N_14561,N_12159,N_12453);
and U14562 (N_14562,N_12060,N_11648);
and U14563 (N_14563,N_12121,N_10547);
nor U14564 (N_14564,N_10364,N_12088);
nand U14565 (N_14565,N_10858,N_12092);
xnor U14566 (N_14566,N_11775,N_11792);
nand U14567 (N_14567,N_11189,N_11576);
and U14568 (N_14568,N_10013,N_10629);
and U14569 (N_14569,N_10666,N_11183);
xnor U14570 (N_14570,N_11278,N_11334);
nand U14571 (N_14571,N_11353,N_11448);
and U14572 (N_14572,N_12492,N_11734);
nand U14573 (N_14573,N_11252,N_11213);
or U14574 (N_14574,N_11769,N_10154);
nand U14575 (N_14575,N_11065,N_10280);
and U14576 (N_14576,N_11501,N_10820);
nor U14577 (N_14577,N_11347,N_10759);
nor U14578 (N_14578,N_11238,N_10808);
and U14579 (N_14579,N_11384,N_12440);
nand U14580 (N_14580,N_11077,N_12015);
nand U14581 (N_14581,N_12267,N_10708);
nor U14582 (N_14582,N_11026,N_11668);
nor U14583 (N_14583,N_10189,N_12228);
xor U14584 (N_14584,N_12123,N_12036);
nand U14585 (N_14585,N_10761,N_12249);
or U14586 (N_14586,N_10308,N_11557);
or U14587 (N_14587,N_11643,N_10280);
or U14588 (N_14588,N_12254,N_11973);
or U14589 (N_14589,N_11542,N_11401);
nor U14590 (N_14590,N_12250,N_11092);
nand U14591 (N_14591,N_11287,N_10350);
nand U14592 (N_14592,N_11188,N_10804);
xnor U14593 (N_14593,N_12341,N_10923);
nand U14594 (N_14594,N_11512,N_10291);
xor U14595 (N_14595,N_10648,N_11363);
nor U14596 (N_14596,N_11736,N_10206);
nor U14597 (N_14597,N_10005,N_10707);
nor U14598 (N_14598,N_12128,N_10999);
nor U14599 (N_14599,N_12457,N_10466);
nor U14600 (N_14600,N_10392,N_10993);
nor U14601 (N_14601,N_10470,N_12473);
or U14602 (N_14602,N_11118,N_10459);
nand U14603 (N_14603,N_10963,N_10923);
or U14604 (N_14604,N_12327,N_11377);
and U14605 (N_14605,N_10058,N_10890);
and U14606 (N_14606,N_11933,N_11672);
nand U14607 (N_14607,N_12426,N_10642);
and U14608 (N_14608,N_12112,N_10736);
xnor U14609 (N_14609,N_10133,N_10143);
nor U14610 (N_14610,N_11598,N_10363);
nand U14611 (N_14611,N_11580,N_10188);
nand U14612 (N_14612,N_11249,N_10815);
and U14613 (N_14613,N_11244,N_11837);
or U14614 (N_14614,N_11503,N_11133);
xor U14615 (N_14615,N_11820,N_11878);
nand U14616 (N_14616,N_11446,N_12464);
nand U14617 (N_14617,N_12254,N_11085);
and U14618 (N_14618,N_11535,N_11369);
nor U14619 (N_14619,N_10451,N_10562);
nand U14620 (N_14620,N_11564,N_10570);
xor U14621 (N_14621,N_11835,N_11002);
nor U14622 (N_14622,N_10385,N_10784);
nor U14623 (N_14623,N_10602,N_11268);
or U14624 (N_14624,N_12100,N_10002);
xnor U14625 (N_14625,N_11483,N_10186);
nand U14626 (N_14626,N_10665,N_10498);
nand U14627 (N_14627,N_12382,N_10304);
nor U14628 (N_14628,N_10852,N_10125);
or U14629 (N_14629,N_11101,N_11373);
nor U14630 (N_14630,N_11148,N_11402);
and U14631 (N_14631,N_12109,N_11846);
xor U14632 (N_14632,N_11752,N_12252);
xor U14633 (N_14633,N_12221,N_11581);
nand U14634 (N_14634,N_10918,N_11302);
and U14635 (N_14635,N_11503,N_10816);
or U14636 (N_14636,N_11325,N_11893);
nand U14637 (N_14637,N_10914,N_11699);
or U14638 (N_14638,N_10871,N_11938);
and U14639 (N_14639,N_10756,N_10130);
and U14640 (N_14640,N_10717,N_11366);
or U14641 (N_14641,N_12275,N_10641);
nand U14642 (N_14642,N_12229,N_11764);
or U14643 (N_14643,N_10659,N_11298);
and U14644 (N_14644,N_11951,N_12339);
nand U14645 (N_14645,N_11147,N_11794);
or U14646 (N_14646,N_10841,N_11211);
nor U14647 (N_14647,N_10499,N_11545);
nand U14648 (N_14648,N_11047,N_12488);
xor U14649 (N_14649,N_12092,N_11648);
nand U14650 (N_14650,N_10643,N_11098);
xnor U14651 (N_14651,N_10321,N_11379);
or U14652 (N_14652,N_11406,N_12156);
or U14653 (N_14653,N_11046,N_10257);
and U14654 (N_14654,N_10056,N_11947);
nand U14655 (N_14655,N_10705,N_10986);
and U14656 (N_14656,N_10239,N_11767);
nor U14657 (N_14657,N_11933,N_12190);
or U14658 (N_14658,N_11326,N_11060);
nor U14659 (N_14659,N_10006,N_11744);
nor U14660 (N_14660,N_12202,N_11728);
and U14661 (N_14661,N_11500,N_12357);
or U14662 (N_14662,N_10013,N_10843);
and U14663 (N_14663,N_12166,N_10815);
and U14664 (N_14664,N_12014,N_10811);
nand U14665 (N_14665,N_11215,N_10941);
and U14666 (N_14666,N_11194,N_10736);
or U14667 (N_14667,N_11216,N_10824);
nand U14668 (N_14668,N_12134,N_10702);
and U14669 (N_14669,N_10358,N_10475);
nor U14670 (N_14670,N_10478,N_11724);
or U14671 (N_14671,N_10177,N_12256);
nor U14672 (N_14672,N_10795,N_12293);
nor U14673 (N_14673,N_10864,N_11802);
and U14674 (N_14674,N_12449,N_11520);
nand U14675 (N_14675,N_11788,N_10143);
nor U14676 (N_14676,N_12013,N_12134);
and U14677 (N_14677,N_11002,N_10318);
and U14678 (N_14678,N_10373,N_12090);
nand U14679 (N_14679,N_10154,N_11021);
nand U14680 (N_14680,N_12056,N_11846);
and U14681 (N_14681,N_11557,N_11624);
nor U14682 (N_14682,N_10453,N_11482);
or U14683 (N_14683,N_12196,N_12033);
xor U14684 (N_14684,N_10746,N_10337);
nand U14685 (N_14685,N_12222,N_10299);
or U14686 (N_14686,N_10670,N_10530);
nor U14687 (N_14687,N_10680,N_11250);
xnor U14688 (N_14688,N_10772,N_11667);
nand U14689 (N_14689,N_12492,N_10138);
and U14690 (N_14690,N_11538,N_12089);
or U14691 (N_14691,N_11129,N_10696);
nand U14692 (N_14692,N_12167,N_10776);
nor U14693 (N_14693,N_12097,N_10320);
xor U14694 (N_14694,N_11799,N_10922);
or U14695 (N_14695,N_10112,N_10220);
nor U14696 (N_14696,N_10295,N_11273);
and U14697 (N_14697,N_11500,N_10307);
nand U14698 (N_14698,N_10934,N_10774);
and U14699 (N_14699,N_11925,N_10213);
nand U14700 (N_14700,N_12179,N_11268);
xnor U14701 (N_14701,N_11578,N_11740);
and U14702 (N_14702,N_12462,N_10488);
nand U14703 (N_14703,N_10470,N_10894);
and U14704 (N_14704,N_10276,N_10204);
or U14705 (N_14705,N_11115,N_10607);
xor U14706 (N_14706,N_11701,N_11940);
and U14707 (N_14707,N_10238,N_12301);
or U14708 (N_14708,N_10552,N_11246);
or U14709 (N_14709,N_10717,N_11954);
or U14710 (N_14710,N_11906,N_10177);
and U14711 (N_14711,N_10521,N_10537);
or U14712 (N_14712,N_11100,N_12417);
and U14713 (N_14713,N_12264,N_10736);
nand U14714 (N_14714,N_12419,N_11019);
nor U14715 (N_14715,N_11761,N_10724);
or U14716 (N_14716,N_11830,N_11020);
xnor U14717 (N_14717,N_11146,N_10873);
and U14718 (N_14718,N_10997,N_11815);
or U14719 (N_14719,N_11587,N_12168);
nand U14720 (N_14720,N_11105,N_12298);
xor U14721 (N_14721,N_10730,N_10186);
nand U14722 (N_14722,N_12186,N_10343);
nand U14723 (N_14723,N_12180,N_11240);
nand U14724 (N_14724,N_11232,N_11868);
nand U14725 (N_14725,N_12096,N_12325);
and U14726 (N_14726,N_11699,N_11982);
or U14727 (N_14727,N_12136,N_12408);
or U14728 (N_14728,N_12199,N_10281);
nand U14729 (N_14729,N_11123,N_12326);
or U14730 (N_14730,N_11014,N_11335);
or U14731 (N_14731,N_11535,N_10997);
or U14732 (N_14732,N_10910,N_12001);
nand U14733 (N_14733,N_11836,N_10677);
or U14734 (N_14734,N_11415,N_10483);
nor U14735 (N_14735,N_10577,N_11914);
nor U14736 (N_14736,N_11632,N_10909);
xor U14737 (N_14737,N_11844,N_10521);
or U14738 (N_14738,N_10455,N_11034);
nor U14739 (N_14739,N_10540,N_11148);
nor U14740 (N_14740,N_10059,N_11990);
nor U14741 (N_14741,N_10675,N_12452);
nand U14742 (N_14742,N_10628,N_11222);
nand U14743 (N_14743,N_10580,N_10830);
or U14744 (N_14744,N_12455,N_10385);
xnor U14745 (N_14745,N_11363,N_10158);
nor U14746 (N_14746,N_12478,N_11457);
or U14747 (N_14747,N_12168,N_10180);
nand U14748 (N_14748,N_11262,N_10180);
and U14749 (N_14749,N_12003,N_10308);
xor U14750 (N_14750,N_11502,N_10160);
or U14751 (N_14751,N_11063,N_10424);
nor U14752 (N_14752,N_12491,N_11776);
and U14753 (N_14753,N_11186,N_12257);
nor U14754 (N_14754,N_10392,N_12401);
nand U14755 (N_14755,N_12110,N_12348);
nor U14756 (N_14756,N_11150,N_10481);
nor U14757 (N_14757,N_10375,N_12447);
nor U14758 (N_14758,N_12348,N_10747);
nand U14759 (N_14759,N_12225,N_11536);
nor U14760 (N_14760,N_12016,N_10284);
nand U14761 (N_14761,N_10790,N_11826);
nor U14762 (N_14762,N_10203,N_12357);
and U14763 (N_14763,N_10046,N_12362);
or U14764 (N_14764,N_10456,N_10917);
or U14765 (N_14765,N_11859,N_11945);
and U14766 (N_14766,N_11273,N_10876);
or U14767 (N_14767,N_12257,N_10069);
nand U14768 (N_14768,N_10006,N_10039);
or U14769 (N_14769,N_12482,N_12234);
or U14770 (N_14770,N_12201,N_12104);
nor U14771 (N_14771,N_11966,N_11472);
and U14772 (N_14772,N_10870,N_12344);
nand U14773 (N_14773,N_11114,N_10119);
nor U14774 (N_14774,N_11940,N_11082);
and U14775 (N_14775,N_11849,N_11020);
nand U14776 (N_14776,N_11575,N_11837);
or U14777 (N_14777,N_11557,N_12272);
or U14778 (N_14778,N_12296,N_10165);
and U14779 (N_14779,N_10666,N_12449);
nor U14780 (N_14780,N_10581,N_11888);
nor U14781 (N_14781,N_12008,N_12286);
and U14782 (N_14782,N_11185,N_11085);
or U14783 (N_14783,N_11436,N_11754);
nor U14784 (N_14784,N_11623,N_12447);
or U14785 (N_14785,N_10103,N_10410);
nand U14786 (N_14786,N_12225,N_11589);
nor U14787 (N_14787,N_11706,N_10228);
nand U14788 (N_14788,N_10018,N_10680);
and U14789 (N_14789,N_10533,N_11115);
nor U14790 (N_14790,N_12226,N_12091);
nor U14791 (N_14791,N_12336,N_10434);
or U14792 (N_14792,N_10162,N_11360);
and U14793 (N_14793,N_12377,N_11627);
xor U14794 (N_14794,N_12402,N_10280);
nand U14795 (N_14795,N_10632,N_12463);
and U14796 (N_14796,N_11279,N_10118);
nand U14797 (N_14797,N_11796,N_10048);
or U14798 (N_14798,N_10859,N_10853);
or U14799 (N_14799,N_10680,N_12269);
nor U14800 (N_14800,N_10147,N_12019);
nor U14801 (N_14801,N_12451,N_10459);
and U14802 (N_14802,N_11645,N_10499);
and U14803 (N_14803,N_12089,N_10752);
nand U14804 (N_14804,N_10557,N_11262);
xnor U14805 (N_14805,N_11940,N_11232);
or U14806 (N_14806,N_11026,N_10898);
or U14807 (N_14807,N_10728,N_10474);
or U14808 (N_14808,N_10716,N_10120);
and U14809 (N_14809,N_11980,N_11870);
or U14810 (N_14810,N_11026,N_11782);
or U14811 (N_14811,N_11574,N_12080);
xor U14812 (N_14812,N_12294,N_11738);
or U14813 (N_14813,N_10300,N_10502);
nand U14814 (N_14814,N_12131,N_10907);
or U14815 (N_14815,N_12353,N_11555);
or U14816 (N_14816,N_12287,N_10161);
xnor U14817 (N_14817,N_11706,N_11983);
nand U14818 (N_14818,N_11474,N_11373);
and U14819 (N_14819,N_10131,N_10526);
and U14820 (N_14820,N_10178,N_12244);
and U14821 (N_14821,N_12123,N_12099);
nor U14822 (N_14822,N_10473,N_11461);
nand U14823 (N_14823,N_10998,N_11450);
nand U14824 (N_14824,N_11711,N_11975);
or U14825 (N_14825,N_11358,N_12464);
and U14826 (N_14826,N_11367,N_11973);
nor U14827 (N_14827,N_12323,N_11553);
xor U14828 (N_14828,N_11857,N_12136);
or U14829 (N_14829,N_11902,N_11439);
xor U14830 (N_14830,N_10053,N_11679);
nor U14831 (N_14831,N_11218,N_11651);
nor U14832 (N_14832,N_11440,N_11704);
nand U14833 (N_14833,N_12463,N_11290);
or U14834 (N_14834,N_10392,N_11564);
or U14835 (N_14835,N_10959,N_10638);
or U14836 (N_14836,N_10862,N_10092);
nand U14837 (N_14837,N_10139,N_10174);
nor U14838 (N_14838,N_10718,N_10111);
and U14839 (N_14839,N_11309,N_11048);
xor U14840 (N_14840,N_11770,N_12390);
nor U14841 (N_14841,N_10268,N_10226);
nand U14842 (N_14842,N_11489,N_12367);
and U14843 (N_14843,N_10085,N_11482);
nand U14844 (N_14844,N_11021,N_12029);
nor U14845 (N_14845,N_10516,N_12094);
nand U14846 (N_14846,N_11134,N_11682);
nor U14847 (N_14847,N_11014,N_11707);
and U14848 (N_14848,N_10799,N_10412);
nor U14849 (N_14849,N_10485,N_11598);
nand U14850 (N_14850,N_10500,N_10116);
nand U14851 (N_14851,N_11641,N_11536);
or U14852 (N_14852,N_10030,N_11504);
or U14853 (N_14853,N_11579,N_11404);
and U14854 (N_14854,N_11036,N_12123);
nand U14855 (N_14855,N_10098,N_10186);
and U14856 (N_14856,N_11471,N_10598);
nor U14857 (N_14857,N_11585,N_11649);
nor U14858 (N_14858,N_11533,N_10982);
nor U14859 (N_14859,N_11856,N_12259);
and U14860 (N_14860,N_11577,N_12392);
or U14861 (N_14861,N_11851,N_11623);
or U14862 (N_14862,N_10149,N_11727);
nand U14863 (N_14863,N_10560,N_12487);
and U14864 (N_14864,N_10088,N_10227);
and U14865 (N_14865,N_10470,N_10903);
and U14866 (N_14866,N_10026,N_12198);
or U14867 (N_14867,N_11479,N_12099);
and U14868 (N_14868,N_11202,N_12198);
xor U14869 (N_14869,N_11532,N_12116);
and U14870 (N_14870,N_12445,N_10015);
nand U14871 (N_14871,N_11382,N_11269);
nand U14872 (N_14872,N_10020,N_10153);
nand U14873 (N_14873,N_10847,N_11016);
or U14874 (N_14874,N_11151,N_10579);
nor U14875 (N_14875,N_12020,N_12471);
or U14876 (N_14876,N_10505,N_11130);
nand U14877 (N_14877,N_11102,N_11471);
nor U14878 (N_14878,N_11276,N_11811);
xnor U14879 (N_14879,N_10608,N_12155);
xnor U14880 (N_14880,N_11207,N_11707);
nor U14881 (N_14881,N_10640,N_11407);
nand U14882 (N_14882,N_10344,N_11593);
nand U14883 (N_14883,N_12496,N_11976);
nand U14884 (N_14884,N_11769,N_12325);
or U14885 (N_14885,N_11945,N_10602);
nor U14886 (N_14886,N_12282,N_11790);
or U14887 (N_14887,N_10925,N_10556);
or U14888 (N_14888,N_12337,N_10882);
and U14889 (N_14889,N_11122,N_12268);
nor U14890 (N_14890,N_10191,N_11557);
and U14891 (N_14891,N_10924,N_12062);
xnor U14892 (N_14892,N_11163,N_10208);
nand U14893 (N_14893,N_10022,N_12226);
nor U14894 (N_14894,N_10258,N_11283);
nand U14895 (N_14895,N_11340,N_11547);
nor U14896 (N_14896,N_10705,N_11994);
and U14897 (N_14897,N_10262,N_10612);
or U14898 (N_14898,N_10329,N_12499);
nand U14899 (N_14899,N_11625,N_11185);
xor U14900 (N_14900,N_11728,N_11461);
nor U14901 (N_14901,N_11676,N_11698);
nor U14902 (N_14902,N_10313,N_10733);
and U14903 (N_14903,N_10062,N_12390);
or U14904 (N_14904,N_11479,N_10876);
nor U14905 (N_14905,N_11215,N_10312);
or U14906 (N_14906,N_10360,N_11817);
or U14907 (N_14907,N_10030,N_11043);
and U14908 (N_14908,N_11590,N_11874);
or U14909 (N_14909,N_11331,N_12310);
xnor U14910 (N_14910,N_10259,N_11203);
xor U14911 (N_14911,N_12047,N_11236);
nand U14912 (N_14912,N_10033,N_10542);
nand U14913 (N_14913,N_10668,N_11419);
or U14914 (N_14914,N_11105,N_12346);
nand U14915 (N_14915,N_12319,N_11645);
and U14916 (N_14916,N_11344,N_11181);
nand U14917 (N_14917,N_12299,N_11936);
and U14918 (N_14918,N_10337,N_10777);
or U14919 (N_14919,N_11708,N_11989);
nand U14920 (N_14920,N_11257,N_11923);
or U14921 (N_14921,N_11524,N_10468);
nor U14922 (N_14922,N_10029,N_10513);
nand U14923 (N_14923,N_11204,N_11441);
and U14924 (N_14924,N_10248,N_11624);
or U14925 (N_14925,N_10693,N_11531);
and U14926 (N_14926,N_12273,N_10685);
nand U14927 (N_14927,N_11181,N_10050);
nor U14928 (N_14928,N_12059,N_10761);
nor U14929 (N_14929,N_10582,N_12102);
nor U14930 (N_14930,N_11606,N_10089);
and U14931 (N_14931,N_12306,N_10246);
and U14932 (N_14932,N_10770,N_10841);
and U14933 (N_14933,N_11206,N_10482);
or U14934 (N_14934,N_12171,N_12275);
nand U14935 (N_14935,N_11850,N_11893);
nor U14936 (N_14936,N_12492,N_11198);
nor U14937 (N_14937,N_11785,N_12436);
or U14938 (N_14938,N_10439,N_12409);
nand U14939 (N_14939,N_10672,N_12159);
nand U14940 (N_14940,N_10941,N_12477);
or U14941 (N_14941,N_11202,N_10168);
and U14942 (N_14942,N_12462,N_10539);
xor U14943 (N_14943,N_11027,N_11905);
nand U14944 (N_14944,N_11574,N_12221);
nand U14945 (N_14945,N_11184,N_10105);
nor U14946 (N_14946,N_12166,N_10371);
or U14947 (N_14947,N_12067,N_10144);
and U14948 (N_14948,N_12290,N_11064);
or U14949 (N_14949,N_10632,N_10202);
nand U14950 (N_14950,N_11999,N_10669);
or U14951 (N_14951,N_10227,N_10146);
nand U14952 (N_14952,N_11410,N_11386);
or U14953 (N_14953,N_12343,N_10661);
and U14954 (N_14954,N_10906,N_10471);
nor U14955 (N_14955,N_10751,N_10428);
nand U14956 (N_14956,N_10064,N_12075);
and U14957 (N_14957,N_10719,N_12295);
and U14958 (N_14958,N_10060,N_11288);
nor U14959 (N_14959,N_11679,N_10182);
xnor U14960 (N_14960,N_10442,N_10218);
nand U14961 (N_14961,N_11221,N_11923);
nor U14962 (N_14962,N_10600,N_11749);
nand U14963 (N_14963,N_12314,N_11863);
nor U14964 (N_14964,N_11062,N_10629);
nand U14965 (N_14965,N_11969,N_12163);
or U14966 (N_14966,N_10465,N_10752);
and U14967 (N_14967,N_10899,N_11761);
nor U14968 (N_14968,N_11409,N_10257);
nor U14969 (N_14969,N_10324,N_12251);
and U14970 (N_14970,N_11275,N_12153);
nand U14971 (N_14971,N_12399,N_10392);
nand U14972 (N_14972,N_10605,N_12309);
xor U14973 (N_14973,N_10315,N_11807);
nor U14974 (N_14974,N_11855,N_11945);
and U14975 (N_14975,N_10703,N_11408);
or U14976 (N_14976,N_10939,N_10484);
or U14977 (N_14977,N_11870,N_10764);
xnor U14978 (N_14978,N_10424,N_10418);
nor U14979 (N_14979,N_11952,N_11436);
nand U14980 (N_14980,N_10880,N_10191);
nor U14981 (N_14981,N_11318,N_10875);
and U14982 (N_14982,N_11080,N_11746);
or U14983 (N_14983,N_11619,N_10089);
nand U14984 (N_14984,N_10169,N_11143);
or U14985 (N_14985,N_10704,N_11330);
nor U14986 (N_14986,N_12416,N_11078);
or U14987 (N_14987,N_10202,N_11192);
nor U14988 (N_14988,N_10576,N_10749);
and U14989 (N_14989,N_12423,N_11154);
nor U14990 (N_14990,N_11544,N_10264);
nand U14991 (N_14991,N_11011,N_10411);
xor U14992 (N_14992,N_11559,N_11236);
xnor U14993 (N_14993,N_12466,N_10010);
nand U14994 (N_14994,N_10340,N_11228);
nand U14995 (N_14995,N_11852,N_12266);
nor U14996 (N_14996,N_12216,N_12164);
xnor U14997 (N_14997,N_11035,N_11641);
nor U14998 (N_14998,N_11949,N_11852);
nand U14999 (N_14999,N_10243,N_11727);
nand U15000 (N_15000,N_13059,N_13776);
and U15001 (N_15001,N_14098,N_12840);
nand U15002 (N_15002,N_13124,N_13727);
nand U15003 (N_15003,N_14709,N_14151);
xnor U15004 (N_15004,N_12947,N_12918);
or U15005 (N_15005,N_13288,N_14786);
nand U15006 (N_15006,N_13627,N_13345);
xor U15007 (N_15007,N_14117,N_12533);
nor U15008 (N_15008,N_13431,N_14582);
and U15009 (N_15009,N_12861,N_14240);
and U15010 (N_15010,N_13144,N_12895);
and U15011 (N_15011,N_13471,N_14630);
and U15012 (N_15012,N_12755,N_12558);
nor U15013 (N_15013,N_13879,N_14453);
nand U15014 (N_15014,N_12700,N_12789);
and U15015 (N_15015,N_13182,N_14733);
nor U15016 (N_15016,N_13433,N_13874);
xor U15017 (N_15017,N_14533,N_14219);
xor U15018 (N_15018,N_14579,N_14134);
nor U15019 (N_15019,N_14947,N_13268);
and U15020 (N_15020,N_13284,N_13725);
nand U15021 (N_15021,N_13826,N_13200);
and U15022 (N_15022,N_14758,N_13617);
and U15023 (N_15023,N_14738,N_13639);
and U15024 (N_15024,N_12961,N_14862);
nand U15025 (N_15025,N_14973,N_14030);
nor U15026 (N_15026,N_13888,N_13326);
nand U15027 (N_15027,N_13738,N_14093);
nand U15028 (N_15028,N_12886,N_13553);
or U15029 (N_15029,N_12848,N_14596);
nand U15030 (N_15030,N_14872,N_14616);
and U15031 (N_15031,N_13536,N_12740);
nand U15032 (N_15032,N_14992,N_13550);
nand U15033 (N_15033,N_12667,N_13171);
nand U15034 (N_15034,N_12715,N_12856);
or U15035 (N_15035,N_13451,N_14879);
nand U15036 (N_15036,N_14585,N_12636);
and U15037 (N_15037,N_14624,N_13159);
nor U15038 (N_15038,N_14346,N_13321);
and U15039 (N_15039,N_13971,N_14819);
or U15040 (N_15040,N_14195,N_14395);
nand U15041 (N_15041,N_12993,N_13744);
nand U15042 (N_15042,N_14713,N_14995);
and U15043 (N_15043,N_12821,N_13071);
xor U15044 (N_15044,N_14405,N_13253);
nand U15045 (N_15045,N_14534,N_14642);
and U15046 (N_15046,N_12726,N_13134);
or U15047 (N_15047,N_14573,N_13614);
and U15048 (N_15048,N_12983,N_13648);
or U15049 (N_15049,N_13298,N_12938);
nand U15050 (N_15050,N_13684,N_13101);
nand U15051 (N_15051,N_13573,N_13166);
or U15052 (N_15052,N_13294,N_14000);
or U15053 (N_15053,N_14291,N_13419);
nand U15054 (N_15054,N_14551,N_13848);
and U15055 (N_15055,N_13031,N_14181);
or U15056 (N_15056,N_12833,N_14442);
and U15057 (N_15057,N_14806,N_13849);
or U15058 (N_15058,N_12600,N_13003);
or U15059 (N_15059,N_13790,N_12772);
nor U15060 (N_15060,N_13440,N_14572);
or U15061 (N_15061,N_14634,N_14594);
or U15062 (N_15062,N_12505,N_13760);
nand U15063 (N_15063,N_14621,N_14179);
or U15064 (N_15064,N_14329,N_14741);
or U15065 (N_15065,N_12682,N_13740);
or U15066 (N_15066,N_13339,N_14892);
nor U15067 (N_15067,N_14787,N_12515);
nor U15068 (N_15068,N_14568,N_14148);
and U15069 (N_15069,N_12501,N_12539);
or U15070 (N_15070,N_14189,N_13198);
and U15071 (N_15071,N_12666,N_14650);
xor U15072 (N_15072,N_12956,N_13683);
xnor U15073 (N_15073,N_14988,N_12550);
or U15074 (N_15074,N_14658,N_14712);
nand U15075 (N_15075,N_14717,N_14601);
and U15076 (N_15076,N_14318,N_13328);
or U15077 (N_15077,N_14206,N_12754);
xor U15078 (N_15078,N_13677,N_12637);
nor U15079 (N_15079,N_13434,N_13518);
nor U15080 (N_15080,N_14505,N_13331);
or U15081 (N_15081,N_14675,N_14818);
nor U15082 (N_15082,N_14916,N_13105);
xnor U15083 (N_15083,N_12770,N_14150);
xor U15084 (N_15084,N_13482,N_13791);
nor U15085 (N_15085,N_12785,N_12508);
nand U15086 (N_15086,N_13396,N_14677);
and U15087 (N_15087,N_14834,N_13370);
xnor U15088 (N_15088,N_14428,N_14792);
nor U15089 (N_15089,N_14767,N_13523);
nand U15090 (N_15090,N_13570,N_13317);
or U15091 (N_15091,N_13155,N_13717);
nand U15092 (N_15092,N_12572,N_14719);
nand U15093 (N_15093,N_14425,N_14183);
xnor U15094 (N_15094,N_12967,N_13384);
and U15095 (N_15095,N_12719,N_13947);
nand U15096 (N_15096,N_13704,N_14293);
and U15097 (N_15097,N_14320,N_13883);
and U15098 (N_15098,N_12589,N_14258);
or U15099 (N_15099,N_13452,N_13530);
nand U15100 (N_15100,N_12899,N_13873);
or U15101 (N_15101,N_14742,N_14218);
nand U15102 (N_15102,N_12880,N_14952);
xor U15103 (N_15103,N_14904,N_14244);
nor U15104 (N_15104,N_14536,N_12894);
nor U15105 (N_15105,N_12592,N_13227);
and U15106 (N_15106,N_13663,N_14454);
and U15107 (N_15107,N_12900,N_13931);
or U15108 (N_15108,N_12520,N_13800);
or U15109 (N_15109,N_13803,N_14427);
nand U15110 (N_15110,N_14580,N_13854);
or U15111 (N_15111,N_14489,N_12858);
nand U15112 (N_15112,N_14790,N_13205);
or U15113 (N_15113,N_14173,N_14625);
or U15114 (N_15114,N_14363,N_14079);
and U15115 (N_15115,N_13807,N_13492);
nor U15116 (N_15116,N_13167,N_12563);
nor U15117 (N_15117,N_12925,N_14822);
nor U15118 (N_15118,N_14914,N_14578);
or U15119 (N_15119,N_13611,N_12642);
nand U15120 (N_15120,N_13732,N_13042);
nor U15121 (N_15121,N_12807,N_14707);
nor U15122 (N_15122,N_14004,N_12962);
or U15123 (N_15123,N_13246,N_14043);
and U15124 (N_15124,N_12885,N_13590);
and U15125 (N_15125,N_13259,N_14070);
xor U15126 (N_15126,N_13325,N_14076);
nand U15127 (N_15127,N_14403,N_14488);
nand U15128 (N_15128,N_13481,N_13232);
nor U15129 (N_15129,N_14492,N_13972);
nor U15130 (N_15130,N_13443,N_13699);
xor U15131 (N_15131,N_14358,N_14276);
nor U15132 (N_15132,N_13464,N_14899);
nor U15133 (N_15133,N_14845,N_14559);
or U15134 (N_15134,N_13587,N_14417);
nand U15135 (N_15135,N_14801,N_14101);
and U15136 (N_15136,N_12676,N_14471);
and U15137 (N_15137,N_12898,N_13889);
or U15138 (N_15138,N_14993,N_12901);
nand U15139 (N_15139,N_14884,N_12929);
or U15140 (N_15140,N_14386,N_13556);
nand U15141 (N_15141,N_14273,N_12613);
nor U15142 (N_15142,N_13568,N_12564);
nand U15143 (N_15143,N_12705,N_13034);
or U15144 (N_15144,N_13912,N_13867);
or U15145 (N_15145,N_12775,N_12619);
or U15146 (N_15146,N_13162,N_12650);
nor U15147 (N_15147,N_14300,N_14754);
or U15148 (N_15148,N_13706,N_12988);
xnor U15149 (N_15149,N_13187,N_14739);
nand U15150 (N_15150,N_14656,N_14774);
nor U15151 (N_15151,N_14635,N_14651);
nor U15152 (N_15152,N_13956,N_14356);
or U15153 (N_15153,N_14722,N_13930);
nor U15154 (N_15154,N_13652,N_13483);
and U15155 (N_15155,N_14521,N_13705);
and U15156 (N_15156,N_14493,N_12949);
nand U15157 (N_15157,N_13884,N_12603);
nand U15158 (N_15158,N_14986,N_12915);
nand U15159 (N_15159,N_14788,N_13675);
nand U15160 (N_15160,N_14322,N_13377);
and U15161 (N_15161,N_13610,N_13851);
or U15162 (N_15162,N_12575,N_12966);
and U15163 (N_15163,N_12826,N_12626);
or U15164 (N_15164,N_13756,N_13881);
or U15165 (N_15165,N_13604,N_14599);
or U15166 (N_15166,N_12679,N_13635);
or U15167 (N_15167,N_13168,N_13479);
nand U15168 (N_15168,N_14216,N_14160);
nor U15169 (N_15169,N_13001,N_14360);
nand U15170 (N_15170,N_13901,N_14750);
nor U15171 (N_15171,N_13835,N_14296);
nand U15172 (N_15172,N_13577,N_14779);
and U15173 (N_15173,N_14543,N_13494);
xor U15174 (N_15174,N_14416,N_14220);
nor U15175 (N_15175,N_12698,N_14145);
and U15176 (N_15176,N_12732,N_13092);
or U15177 (N_15177,N_13117,N_12546);
or U15178 (N_15178,N_13600,N_13358);
xor U15179 (N_15179,N_14752,N_14736);
xor U15180 (N_15180,N_13176,N_13542);
xor U15181 (N_15181,N_14807,N_14950);
or U15182 (N_15182,N_14923,N_14481);
or U15183 (N_15183,N_14254,N_13334);
nand U15184 (N_15184,N_13619,N_14255);
or U15185 (N_15185,N_13714,N_14515);
nand U15186 (N_15186,N_12681,N_14436);
nor U15187 (N_15187,N_13660,N_13084);
and U15188 (N_15188,N_14411,N_12714);
or U15189 (N_15189,N_13329,N_13301);
xor U15190 (N_15190,N_14919,N_12937);
nor U15191 (N_15191,N_12686,N_14497);
or U15192 (N_15192,N_14540,N_14851);
nor U15193 (N_15193,N_14704,N_13593);
nor U15194 (N_15194,N_13389,N_14928);
and U15195 (N_15195,N_12519,N_12979);
xnor U15196 (N_15196,N_13208,N_13422);
nand U15197 (N_15197,N_13313,N_13609);
nor U15198 (N_15198,N_13870,N_13424);
nand U15199 (N_15199,N_13595,N_13073);
nand U15200 (N_15200,N_13104,N_13856);
and U15201 (N_15201,N_13312,N_14180);
nor U15202 (N_15202,N_14940,N_13916);
nand U15203 (N_15203,N_14887,N_13656);
or U15204 (N_15204,N_14144,N_14143);
or U15205 (N_15205,N_13897,N_12517);
nor U15206 (N_15206,N_14924,N_12828);
nor U15207 (N_15207,N_14569,N_13256);
and U15208 (N_15208,N_14031,N_12994);
nand U15209 (N_15209,N_13465,N_14013);
nand U15210 (N_15210,N_14055,N_13747);
or U15211 (N_15211,N_14646,N_14606);
nand U15212 (N_15212,N_13022,N_13946);
nor U15213 (N_15213,N_14100,N_13505);
or U15214 (N_15214,N_12530,N_13302);
or U15215 (N_15215,N_13153,N_14064);
xor U15216 (N_15216,N_14657,N_14597);
and U15217 (N_15217,N_13236,N_14889);
nor U15218 (N_15218,N_14020,N_14462);
nand U15219 (N_15219,N_13707,N_13002);
or U15220 (N_15220,N_14939,N_14825);
or U15221 (N_15221,N_14494,N_14292);
xor U15222 (N_15222,N_13113,N_14035);
nor U15223 (N_15223,N_14708,N_12786);
and U15224 (N_15224,N_13340,N_12713);
nand U15225 (N_15225,N_14567,N_14918);
and U15226 (N_15226,N_12934,N_13172);
and U15227 (N_15227,N_13346,N_12771);
xor U15228 (N_15228,N_14131,N_14396);
or U15229 (N_15229,N_14522,N_12752);
nand U15230 (N_15230,N_14324,N_13276);
nand U15231 (N_15231,N_14350,N_13291);
nand U15232 (N_15232,N_13769,N_14858);
or U15233 (N_15233,N_13527,N_13837);
nor U15234 (N_15234,N_14478,N_14764);
or U15235 (N_15235,N_13669,N_13624);
nand U15236 (N_15236,N_14590,N_14351);
and U15237 (N_15237,N_13336,N_13563);
xnor U15238 (N_15238,N_13403,N_13662);
and U15239 (N_15239,N_13928,N_13372);
and U15240 (N_15240,N_13671,N_13439);
and U15241 (N_15241,N_13043,N_14404);
xnor U15242 (N_15242,N_13202,N_13233);
or U15243 (N_15243,N_13736,N_12616);
or U15244 (N_15244,N_12566,N_14252);
and U15245 (N_15245,N_14877,N_14169);
and U15246 (N_15246,N_14095,N_13546);
and U15247 (N_15247,N_12980,N_13027);
and U15248 (N_15248,N_14009,N_13351);
and U15249 (N_15249,N_12778,N_13668);
nand U15250 (N_15250,N_14999,N_13632);
nor U15251 (N_15251,N_14636,N_13770);
nand U15252 (N_15252,N_12941,N_14105);
and U15253 (N_15253,N_12823,N_14645);
nand U15254 (N_15254,N_14688,N_14935);
nor U15255 (N_15255,N_13123,N_12627);
and U15256 (N_15256,N_12783,N_14384);
or U15257 (N_15257,N_13984,N_14192);
xnor U15258 (N_15258,N_14217,N_13497);
and U15259 (N_15259,N_14723,N_14971);
nand U15260 (N_15260,N_13075,N_14566);
or U15261 (N_15261,N_14469,N_13189);
and U15262 (N_15262,N_13498,N_12832);
and U15263 (N_15263,N_14294,N_14243);
nand U15264 (N_15264,N_12809,N_14452);
nor U15265 (N_15265,N_13753,N_13140);
xnor U15266 (N_15266,N_12647,N_13575);
or U15267 (N_15267,N_14480,N_13132);
xor U15268 (N_15268,N_14513,N_14987);
or U15269 (N_15269,N_13369,N_12534);
or U15270 (N_15270,N_13041,N_14163);
and U15271 (N_15271,N_12521,N_14332);
or U15272 (N_15272,N_13818,N_12974);
xor U15273 (N_15273,N_13701,N_14418);
nand U15274 (N_15274,N_14498,N_13983);
xnor U15275 (N_15275,N_14575,N_14083);
or U15276 (N_15276,N_12877,N_12611);
and U15277 (N_15277,N_13130,N_14647);
and U15278 (N_15278,N_12645,N_13516);
xor U15279 (N_15279,N_14381,N_12535);
nand U15280 (N_15280,N_14519,N_12510);
or U15281 (N_15281,N_14668,N_13539);
nor U15282 (N_15282,N_13967,N_14793);
and U15283 (N_15283,N_13057,N_14593);
and U15284 (N_15284,N_13891,N_12744);
and U15285 (N_15285,N_12986,N_12855);
xnor U15286 (N_15286,N_14387,N_13773);
nand U15287 (N_15287,N_12882,N_13463);
nand U15288 (N_15288,N_13616,N_14054);
and U15289 (N_15289,N_14484,N_13148);
or U15290 (N_15290,N_12818,N_12707);
nand U15291 (N_15291,N_13455,N_14175);
and U15292 (N_15292,N_14201,N_14434);
xnor U15293 (N_15293,N_14854,N_12867);
nand U15294 (N_15294,N_13560,N_13687);
nor U15295 (N_15295,N_14282,N_14262);
nor U15296 (N_15296,N_13921,N_12608);
and U15297 (N_15297,N_14628,N_13250);
or U15298 (N_15298,N_12927,N_13388);
nand U15299 (N_15299,N_13258,N_13924);
nor U15300 (N_15300,N_12850,N_12531);
nand U15301 (N_15301,N_14860,N_14769);
and U15302 (N_15302,N_14018,N_13193);
or U15303 (N_15303,N_13658,N_13833);
xnor U15304 (N_15304,N_13812,N_14001);
and U15305 (N_15305,N_14383,N_14167);
nand U15306 (N_15306,N_14073,N_14831);
nor U15307 (N_15307,N_13605,N_13949);
nor U15308 (N_15308,N_13032,N_13447);
nor U15309 (N_15309,N_14090,N_13295);
nor U15310 (N_15310,N_13238,N_12952);
nor U15311 (N_15311,N_13968,N_13383);
and U15312 (N_15312,N_13741,N_12606);
nand U15313 (N_15313,N_13794,N_14689);
and U15314 (N_15314,N_13661,N_12609);
and U15315 (N_15315,N_14187,N_12528);
nand U15316 (N_15316,N_13531,N_12944);
and U15317 (N_15317,N_14437,N_13508);
nand U15318 (N_15318,N_12796,N_14047);
and U15319 (N_15319,N_14440,N_14391);
and U15320 (N_15320,N_13063,N_13748);
xnor U15321 (N_15321,N_13923,N_12964);
or U15322 (N_15322,N_13493,N_12583);
nor U15323 (N_15323,N_13911,N_14236);
nor U15324 (N_15324,N_14172,N_14191);
and U15325 (N_15325,N_14005,N_12567);
nand U15326 (N_15326,N_13565,N_13810);
nand U15327 (N_15327,N_13350,N_14603);
nand U15328 (N_15328,N_12646,N_12946);
nand U15329 (N_15329,N_14985,N_14334);
or U15330 (N_15330,N_13024,N_14921);
xor U15331 (N_15331,N_14715,N_14925);
and U15332 (N_15332,N_13926,N_12844);
xnor U15333 (N_15333,N_13417,N_13160);
or U15334 (N_15334,N_14174,N_14905);
xnor U15335 (N_15335,N_13708,N_13391);
nor U15336 (N_15336,N_14979,N_14034);
nor U15337 (N_15337,N_13023,N_14552);
and U15338 (N_15338,N_13230,N_13788);
nor U15339 (N_15339,N_14890,N_13653);
nor U15340 (N_15340,N_12893,N_12588);
and U15341 (N_15341,N_13461,N_14902);
nand U15342 (N_15342,N_12921,N_14755);
or U15343 (N_15343,N_14699,N_14591);
xnor U15344 (N_15344,N_12570,N_13460);
nor U15345 (N_15345,N_14837,N_13135);
or U15346 (N_15346,N_14210,N_14288);
or U15347 (N_15347,N_14354,N_14588);
nand U15348 (N_15348,N_13579,N_12825);
nand U15349 (N_15349,N_14479,N_13960);
and U15350 (N_15350,N_14728,N_14913);
or U15351 (N_15351,N_14137,N_12767);
nor U15352 (N_15352,N_13512,N_13185);
nand U15353 (N_15353,N_12725,N_13603);
and U15354 (N_15354,N_14235,N_14949);
nand U15355 (N_15355,N_14659,N_12751);
nand U15356 (N_15356,N_13502,N_14367);
and U15357 (N_15357,N_14313,N_13371);
or U15358 (N_15358,N_14897,N_13175);
and U15359 (N_15359,N_12928,N_13306);
nor U15360 (N_15360,N_12835,N_14937);
xnor U15361 (N_15361,N_13141,N_13183);
nor U15362 (N_15362,N_14125,N_13715);
and U15363 (N_15363,N_13802,N_12730);
xnor U15364 (N_15364,N_14110,N_12795);
or U15365 (N_15365,N_14112,N_14865);
nor U15366 (N_15366,N_13067,N_14412);
and U15367 (N_15367,N_13941,N_13044);
and U15368 (N_15368,N_12958,N_14827);
and U15369 (N_15369,N_13940,N_14065);
and U15370 (N_15370,N_13589,N_14649);
nor U15371 (N_15371,N_13197,N_13423);
and U15372 (N_15372,N_14305,N_14549);
or U15373 (N_15373,N_13836,N_13091);
nor U15374 (N_15374,N_12942,N_14570);
nor U15375 (N_15375,N_14458,N_14103);
nand U15376 (N_15376,N_12935,N_14036);
nor U15377 (N_15377,N_13862,N_14321);
and U15378 (N_15378,N_12869,N_12760);
nand U15379 (N_15379,N_14190,N_13721);
xnor U15380 (N_15380,N_12595,N_14122);
nand U15381 (N_15381,N_12995,N_14640);
xor U15382 (N_15382,N_13861,N_14287);
and U15383 (N_15383,N_13919,N_13737);
nor U15384 (N_15384,N_13585,N_12635);
nor U15385 (N_15385,N_13225,N_13529);
nand U15386 (N_15386,N_14673,N_14718);
and U15387 (N_15387,N_14895,N_14298);
or U15388 (N_15388,N_14177,N_13842);
xnor U15389 (N_15389,N_14355,N_14060);
or U15390 (N_15390,N_13846,N_13735);
nor U15391 (N_15391,N_13780,N_13201);
xnor U15392 (N_15392,N_12577,N_14523);
and U15393 (N_15393,N_13218,N_14003);
nand U15394 (N_15394,N_14422,N_13213);
or U15395 (N_15395,N_13913,N_13866);
or U15396 (N_15396,N_12593,N_14771);
or U15397 (N_15397,N_13535,N_14873);
or U15398 (N_15398,N_13378,N_13910);
and U15399 (N_15399,N_12883,N_12509);
or U15400 (N_15400,N_12594,N_13990);
or U15401 (N_15401,N_12556,N_13927);
and U15402 (N_15402,N_13880,N_13885);
nand U15403 (N_15403,N_13726,N_14770);
or U15404 (N_15404,N_13337,N_14639);
or U15405 (N_15405,N_14086,N_14204);
and U15406 (N_15406,N_13382,N_14108);
xnor U15407 (N_15407,N_14421,N_13248);
nor U15408 (N_15408,N_14022,N_14375);
nand U15409 (N_15409,N_14188,N_14457);
and U15410 (N_15410,N_13933,N_13942);
or U15411 (N_15411,N_14875,N_13999);
and U15412 (N_15412,N_12862,N_14832);
nor U15413 (N_15413,N_14426,N_13980);
nand U15414 (N_15414,N_13532,N_13262);
nor U15415 (N_15415,N_14406,N_14510);
nor U15416 (N_15416,N_14944,N_13338);
nand U15417 (N_15417,N_14517,N_12954);
nand U15418 (N_15418,N_14976,N_13394);
xor U15419 (N_15419,N_13592,N_12663);
nor U15420 (N_15420,N_12507,N_13580);
nor U15421 (N_15421,N_13872,N_13491);
nor U15422 (N_15422,N_14056,N_13107);
nor U15423 (N_15423,N_13362,N_14265);
nor U15424 (N_15424,N_12683,N_14111);
and U15425 (N_15425,N_12881,N_13899);
or U15426 (N_15426,N_14352,N_13380);
or U15427 (N_15427,N_14158,N_14791);
nor U15428 (N_15428,N_13718,N_14664);
or U15429 (N_15429,N_14909,N_13314);
nor U15430 (N_15430,N_13586,N_14932);
nor U15431 (N_15431,N_14042,N_12782);
nand U15432 (N_15432,N_12662,N_13759);
nor U15433 (N_15433,N_14275,N_14808);
nor U15434 (N_15434,N_14142,N_12585);
nor U15435 (N_15435,N_13551,N_14848);
and U15436 (N_15436,N_14655,N_13713);
xor U15437 (N_15437,N_13249,N_13622);
and U15438 (N_15438,N_14866,N_14824);
nand U15439 (N_15439,N_14325,N_13521);
nand U15440 (N_15440,N_14735,N_14882);
nor U15441 (N_15441,N_13642,N_12654);
nor U15442 (N_15442,N_12815,N_14891);
or U15443 (N_15443,N_14555,N_14136);
nand U15444 (N_15444,N_12649,N_12648);
and U15445 (N_15445,N_12708,N_12685);
and U15446 (N_15446,N_12897,N_13108);
nand U15447 (N_15447,N_13817,N_12513);
nand U15448 (N_15448,N_14432,N_13486);
nand U15449 (N_15449,N_13650,N_12748);
and U15450 (N_15450,N_14953,N_13420);
xnor U15451 (N_15451,N_14246,N_12580);
nor U15452 (N_15452,N_14502,N_13381);
nor U15453 (N_15453,N_13435,N_14113);
and U15454 (N_15454,N_12582,N_14828);
or U15455 (N_15455,N_14785,N_13664);
nand U15456 (N_15456,N_13712,N_13543);
and U15457 (N_15457,N_13226,N_13682);
or U15458 (N_15458,N_13547,N_14227);
nand U15459 (N_15459,N_12784,N_13425);
and U15460 (N_15460,N_13178,N_13771);
and U15461 (N_15461,N_14983,N_13915);
nor U15462 (N_15462,N_13511,N_14341);
and U15463 (N_15463,N_14269,N_14205);
nor U15464 (N_15464,N_13961,N_14789);
nand U15465 (N_15465,N_12989,N_12963);
or U15466 (N_15466,N_14941,N_14978);
nand U15467 (N_15467,N_14900,N_13698);
or U15468 (N_15468,N_12658,N_14053);
nand U15469 (N_15469,N_14149,N_13470);
nor U15470 (N_15470,N_14960,N_14251);
nand U15471 (N_15471,N_14681,N_13427);
nor U15472 (N_15472,N_14997,N_12914);
nor U15473 (N_15473,N_13989,N_14700);
nand U15474 (N_15474,N_13877,N_13569);
nor U15475 (N_15475,N_14701,N_14257);
and U15476 (N_15476,N_13305,N_13673);
nand U15477 (N_15477,N_13286,N_13364);
and U15478 (N_15478,N_14456,N_12644);
and U15479 (N_15479,N_13342,N_14982);
or U15480 (N_15480,N_14162,N_12978);
or U15481 (N_15481,N_13557,N_14438);
or U15482 (N_15482,N_13597,N_14958);
nand U15483 (N_15483,N_14278,N_13363);
nand U15484 (N_15484,N_13680,N_12674);
or U15485 (N_15485,N_13029,N_14577);
or U15486 (N_15486,N_13304,N_13475);
or U15487 (N_15487,N_14221,N_12657);
nand U15488 (N_15488,N_13149,N_13804);
or U15489 (N_15489,N_13049,N_14326);
or U15490 (N_15490,N_12617,N_14512);
nor U15491 (N_15491,N_13028,N_14571);
nand U15492 (N_15492,N_13578,N_13036);
nand U15493 (N_15493,N_13315,N_13118);
or U15494 (N_15494,N_12907,N_14685);
nor U15495 (N_15495,N_14135,N_14608);
nand U15496 (N_15496,N_12889,N_13476);
or U15497 (N_15497,N_14643,N_13733);
or U15498 (N_15498,N_13048,N_13405);
xnor U15499 (N_15499,N_12668,N_14763);
nor U15500 (N_15500,N_14015,N_13277);
and U15501 (N_15501,N_12769,N_14379);
or U15502 (N_15502,N_13824,N_13796);
nand U15503 (N_15503,N_13620,N_14980);
nand U15504 (N_15504,N_12830,N_13678);
nor U15505 (N_15505,N_12597,N_14613);
xor U15506 (N_15506,N_12879,N_14525);
xor U15507 (N_15507,N_14361,N_13103);
nand U15508 (N_15508,N_13853,N_12633);
nand U15509 (N_15509,N_12656,N_13181);
and U15510 (N_15510,N_12598,N_12820);
nand U15511 (N_15511,N_13311,N_12702);
nand U15512 (N_15512,N_14336,N_13240);
or U15513 (N_15513,N_13485,N_14450);
nor U15514 (N_15514,N_14678,N_13774);
and U15515 (N_15515,N_13016,N_14676);
nand U15516 (N_15516,N_13265,N_13739);
nor U15517 (N_15517,N_14279,N_12723);
and U15518 (N_15518,N_13909,N_14804);
nor U15519 (N_15519,N_12610,N_14233);
nand U15520 (N_15520,N_14885,N_14063);
and U15521 (N_15521,N_13018,N_12812);
xor U15522 (N_15522,N_13282,N_14680);
xnor U15523 (N_15523,N_14327,N_14753);
or U15524 (N_15524,N_12684,N_14331);
nand U15525 (N_15525,N_13122,N_14281);
or U15526 (N_15526,N_14448,N_13549);
nor U15527 (N_15527,N_13320,N_13190);
nor U15528 (N_15528,N_13052,N_13805);
nand U15529 (N_15529,N_14429,N_13353);
nand U15530 (N_15530,N_14633,N_12743);
nor U15531 (N_15531,N_14961,N_13019);
and U15532 (N_15532,N_13307,N_14695);
and U15533 (N_15533,N_13814,N_13488);
and U15534 (N_15534,N_12688,N_13986);
nand U15535 (N_15535,N_13723,N_13864);
and U15536 (N_15536,N_12851,N_13467);
nand U15537 (N_15537,N_12799,N_14800);
and U15538 (N_15538,N_13283,N_13962);
xnor U15539 (N_15539,N_14441,N_12839);
or U15540 (N_15540,N_13322,N_14473);
and U15541 (N_15541,N_13068,N_14963);
nor U15542 (N_15542,N_13571,N_13011);
and U15543 (N_15543,N_13444,N_13969);
nand U15544 (N_15544,N_13316,N_14330);
nand U15545 (N_15545,N_14099,N_14365);
and U15546 (N_15546,N_13413,N_14562);
xor U15547 (N_15547,N_13293,N_14618);
or U15548 (N_15548,N_13598,N_13845);
xnor U15549 (N_15549,N_12822,N_13349);
nor U15550 (N_15550,N_12892,N_13533);
or U15551 (N_15551,N_12943,N_12924);
xnor U15552 (N_15552,N_12975,N_13468);
nor U15553 (N_15553,N_14007,N_13400);
nor U15554 (N_15554,N_14344,N_12814);
nand U15555 (N_15555,N_12992,N_12866);
nor U15556 (N_15556,N_14969,N_13822);
nand U15557 (N_15557,N_14424,N_13398);
nand U15558 (N_15558,N_13700,N_14337);
xnor U15559 (N_15559,N_13013,N_12607);
nand U15560 (N_15560,N_13374,N_14981);
and U15561 (N_15561,N_13285,N_14554);
nor U15562 (N_15562,N_12931,N_14045);
and U15563 (N_15563,N_14683,N_13142);
nand U15564 (N_15564,N_14674,N_13072);
and U15565 (N_15565,N_13808,N_12950);
or U15566 (N_15566,N_13562,N_14912);
nand U15567 (N_15567,N_13454,N_14072);
nand U15568 (N_15568,N_13469,N_13210);
or U15569 (N_15569,N_14164,N_14783);
nand U15570 (N_15570,N_14920,N_12669);
nor U15571 (N_15571,N_13418,N_13429);
xnor U15572 (N_15572,N_14716,N_13366);
nor U15573 (N_15573,N_13538,N_14156);
xnor U15574 (N_15574,N_12596,N_12991);
or U15575 (N_15575,N_14795,N_12659);
or U15576 (N_15576,N_13310,N_14798);
and U15577 (N_15577,N_12716,N_13655);
or U15578 (N_15578,N_12761,N_13720);
and U15579 (N_15579,N_14694,N_13365);
nor U15580 (N_15580,N_12587,N_12829);
or U15581 (N_15581,N_13206,N_14538);
xor U15582 (N_15582,N_12870,N_13630);
nor U15583 (N_15583,N_14903,N_14527);
and U15584 (N_15584,N_14665,N_14546);
nor U15585 (N_15585,N_13863,N_13188);
or U15586 (N_15586,N_12905,N_13584);
nand U15587 (N_15587,N_14311,N_13147);
xnor U15588 (N_15588,N_13839,N_13868);
or U15589 (N_15589,N_13273,N_14908);
xor U15590 (N_15590,N_14168,N_14215);
or U15591 (N_15591,N_13456,N_13393);
or U15592 (N_15592,N_12843,N_12909);
or U15593 (N_15593,N_13343,N_13158);
and U15594 (N_15594,N_13843,N_12703);
xnor U15595 (N_15595,N_14721,N_14087);
or U15596 (N_15596,N_13125,N_14362);
nand U15597 (N_15597,N_13534,N_13319);
nor U15598 (N_15598,N_14392,N_14508);
or U15599 (N_15599,N_14611,N_14531);
nor U15600 (N_15600,N_14085,N_12912);
or U15601 (N_15601,N_14152,N_12800);
or U15602 (N_15602,N_12571,N_14420);
nand U15603 (N_15603,N_14012,N_12522);
or U15604 (N_15604,N_14316,N_12804);
or U15605 (N_15605,N_14661,N_13047);
and U15606 (N_15606,N_14869,N_13102);
nand U15607 (N_15607,N_13191,N_13830);
nand U15608 (N_15608,N_13015,N_13763);
and U15609 (N_15609,N_13504,N_13106);
and U15610 (N_15610,N_13169,N_14170);
xnor U15611 (N_15611,N_12801,N_14620);
and U15612 (N_15612,N_14023,N_14413);
nor U15613 (N_15613,N_12888,N_13272);
nand U15614 (N_15614,N_13006,N_12661);
xor U15615 (N_15615,N_14499,N_14951);
or U15616 (N_15616,N_13235,N_14990);
nor U15617 (N_15617,N_13278,N_13582);
and U15618 (N_15618,N_13641,N_14127);
or U15619 (N_15619,N_12565,N_14323);
or U15620 (N_15620,N_13170,N_14141);
nand U15621 (N_15621,N_14198,N_12936);
or U15622 (N_15622,N_14974,N_12639);
nor U15623 (N_15623,N_13938,N_13082);
nor U15624 (N_15624,N_13702,N_14263);
nand U15625 (N_15625,N_14019,N_14041);
nor U15626 (N_15626,N_12803,N_12518);
or U15627 (N_15627,N_13545,N_13778);
or U15628 (N_15628,N_13935,N_13007);
nor U15629 (N_15629,N_14766,N_14878);
nand U15630 (N_15630,N_12538,N_14883);
nand U15631 (N_15631,N_12787,N_13689);
nand U15632 (N_15632,N_14917,N_13174);
nor U15633 (N_15633,N_12781,N_14234);
nand U15634 (N_15634,N_14231,N_12602);
nor U15635 (N_15635,N_13459,N_12773);
nor U15636 (N_15636,N_13355,N_12604);
and U15637 (N_15637,N_13466,N_13361);
nor U15638 (N_15638,N_12951,N_13507);
nor U15639 (N_15639,N_13793,N_14509);
nor U15640 (N_15640,N_13876,N_13697);
or U15641 (N_15641,N_14062,N_13347);
and U15642 (N_15642,N_14846,N_12933);
or U15643 (N_15643,N_14040,N_12971);
nor U15644 (N_15644,N_14302,N_14541);
or U15645 (N_15645,N_13428,N_13367);
xor U15646 (N_15646,N_14408,N_12576);
nor U15647 (N_15647,N_12630,N_14277);
nand U15648 (N_15648,N_13000,N_13973);
or U15649 (N_15649,N_14595,N_14225);
xnor U15650 (N_15650,N_12903,N_13895);
nor U15651 (N_15651,N_13445,N_14929);
or U15652 (N_15652,N_12990,N_13416);
nand U15653 (N_15653,N_13795,N_12853);
xnor U15654 (N_15654,N_12792,N_13050);
nand U15655 (N_15655,N_13066,N_13242);
nand U15656 (N_15656,N_14747,N_13537);
or U15657 (N_15657,N_13267,N_14114);
nand U15658 (N_15658,N_12579,N_14025);
xor U15659 (N_15659,N_13955,N_14778);
and U15660 (N_15660,N_13829,N_14933);
xnor U15661 (N_15661,N_14414,N_13821);
and U15662 (N_15662,N_14886,N_14091);
and U15663 (N_15663,N_14826,N_13121);
nor U15664 (N_15664,N_14956,N_13607);
xnor U15665 (N_15665,N_14830,N_13450);
and U15666 (N_15666,N_13878,N_13857);
or U15667 (N_15667,N_13192,N_13670);
nand U15668 (N_15668,N_13615,N_13847);
and U15669 (N_15669,N_13762,N_12523);
or U15670 (N_15670,N_13640,N_13860);
xnor U15671 (N_15671,N_14816,N_13303);
nor U15672 (N_15672,N_14377,N_14373);
nand U15673 (N_15673,N_14915,N_13711);
nand U15674 (N_15674,N_14838,N_14124);
and U15675 (N_15675,N_12777,N_13917);
nand U15676 (N_15676,N_13035,N_14388);
or U15677 (N_15677,N_14046,N_13647);
or U15678 (N_15678,N_14465,N_14815);
nand U15679 (N_15679,N_12581,N_14214);
xnor U15680 (N_15680,N_13964,N_13978);
or U15681 (N_15681,N_14811,N_12976);
nand U15682 (N_15682,N_13239,N_14161);
nand U15683 (N_15683,N_14107,N_13566);
nor U15684 (N_15684,N_13053,N_13462);
or U15685 (N_15685,N_14349,N_12618);
or U15686 (N_15686,N_14433,N_12762);
nand U15687 (N_15687,N_13021,N_12904);
nor U15688 (N_15688,N_13195,N_13506);
nor U15689 (N_15689,N_14814,N_13629);
nor U15690 (N_15690,N_13564,N_14724);
xnor U15691 (N_15691,N_12678,N_13932);
or U15692 (N_15692,N_14711,N_14203);
nor U15693 (N_15693,N_13709,N_14586);
or U15694 (N_15694,N_13514,N_14859);
xnor U15695 (N_15695,N_13009,N_13894);
nor U15696 (N_15696,N_14380,N_14299);
xnor U15697 (N_15697,N_12728,N_13046);
or U15698 (N_15698,N_14096,N_13244);
nor U15699 (N_15699,N_12836,N_13058);
or U15700 (N_15700,N_14542,N_13038);
nand U15701 (N_15701,N_14032,N_13815);
and U15702 (N_15702,N_13691,N_12798);
or U15703 (N_15703,N_13194,N_13561);
nor U15704 (N_15704,N_12729,N_12875);
and U15705 (N_15705,N_12545,N_13308);
nor U15706 (N_15706,N_14833,N_12960);
or U15707 (N_15707,N_14476,N_13222);
or U15708 (N_15708,N_14314,N_13216);
and U15709 (N_15709,N_14506,N_13207);
xnor U15710 (N_15710,N_14486,N_13255);
nand U15711 (N_15711,N_12614,N_14409);
nand U15712 (N_15712,N_13375,N_13890);
xor U15713 (N_15713,N_13060,N_13281);
nand U15714 (N_15714,N_13540,N_13757);
and U15715 (N_15715,N_14583,N_13397);
and U15716 (N_15716,N_14259,N_12849);
and U15717 (N_15717,N_13583,N_13279);
and U15718 (N_15718,N_14328,N_13922);
nand U15719 (N_15719,N_13750,N_13634);
nor U15720 (N_15720,N_14129,N_14667);
and U15721 (N_15721,N_14842,N_12739);
or U15722 (N_15722,N_13300,N_12673);
or U15723 (N_15723,N_14312,N_13816);
nand U15724 (N_15724,N_14061,N_14295);
nand U15725 (N_15725,N_13012,N_13484);
xor U15726 (N_15726,N_13900,N_14451);
or U15727 (N_15727,N_12996,N_13827);
xnor U15728 (N_15728,N_13613,N_14077);
nor U15729 (N_15729,N_14372,N_14600);
and U15730 (N_15730,N_14393,N_14844);
nor U15731 (N_15731,N_13037,N_13892);
or U15732 (N_15732,N_13840,N_13110);
nor U15733 (N_15733,N_13245,N_12779);
nor U15734 (N_15734,N_13165,N_13496);
or U15735 (N_15735,N_13925,N_12511);
nand U15736 (N_15736,N_13402,N_14014);
nor U15737 (N_15737,N_13356,N_13100);
nor U15738 (N_15738,N_13782,N_12834);
nor U15739 (N_15739,N_13644,N_12532);
or U15740 (N_15740,N_12984,N_13832);
or U15741 (N_15741,N_14307,N_13777);
or U15742 (N_15742,N_14955,N_14128);
nor U15743 (N_15743,N_12601,N_13792);
nand U15744 (N_15744,N_13109,N_12873);
and U15745 (N_15745,N_14229,N_14843);
nand U15746 (N_15746,N_13665,N_12788);
or U15747 (N_15747,N_13693,N_12621);
nand U15748 (N_15748,N_13898,N_13936);
nand U15749 (N_15749,N_13798,N_13729);
nor U15750 (N_15750,N_13089,N_13742);
or U15751 (N_15751,N_14563,N_14455);
nand U15752 (N_15752,N_12643,N_14485);
nor U15753 (N_15753,N_12548,N_14638);
and U15754 (N_15754,N_13667,N_13785);
nor U15755 (N_15755,N_13548,N_14520);
nand U15756 (N_15756,N_14679,N_13772);
or U15757 (N_15757,N_14757,N_13177);
or U15758 (N_15758,N_13156,N_14106);
or U15759 (N_15759,N_12733,N_13120);
nor U15760 (N_15760,N_14342,N_13215);
nor U15761 (N_15761,N_14654,N_14057);
nor U15762 (N_15762,N_12745,N_14368);
and U15763 (N_15763,N_14029,N_14648);
or U15764 (N_15764,N_14821,N_12997);
and U15765 (N_15765,N_13591,N_14861);
or U15766 (N_15766,N_13404,N_12512);
nor U15767 (N_15767,N_12859,N_13929);
nor U15768 (N_15768,N_14071,N_13186);
nand U15769 (N_15769,N_13692,N_13975);
xnor U15770 (N_15770,N_13332,N_13229);
nand U15771 (N_15771,N_12884,N_14684);
nor U15772 (N_15772,N_13994,N_13251);
xor U15773 (N_15773,N_14272,N_14871);
xnor U15774 (N_15774,N_13243,N_14690);
or U15775 (N_15775,N_13976,N_12712);
nor U15776 (N_15776,N_14439,N_14548);
or U15777 (N_15777,N_12691,N_13982);
nand U15778 (N_15778,N_12837,N_12776);
or U15779 (N_15779,N_13524,N_14906);
nor U15780 (N_15780,N_14006,N_14102);
nand U15781 (N_15781,N_13775,N_14672);
nor U15782 (N_15782,N_13287,N_13636);
nor U15783 (N_15783,N_12765,N_14490);
or U15784 (N_15784,N_14415,N_13767);
or U15785 (N_15785,N_14178,N_13241);
or U15786 (N_15786,N_12696,N_14423);
and U15787 (N_15787,N_13051,N_13408);
or U15788 (N_15788,N_14930,N_14274);
nor U15789 (N_15789,N_13752,N_14202);
or U15790 (N_15790,N_14430,N_14765);
nor U15791 (N_15791,N_13478,N_14619);
xor U15792 (N_15792,N_14338,N_14853);
xor U15793 (N_15793,N_12675,N_14027);
nand U15794 (N_15794,N_13765,N_12640);
nor U15795 (N_15795,N_12845,N_12756);
nand U15796 (N_15796,N_14706,N_14376);
nand U15797 (N_15797,N_12802,N_14615);
or U15798 (N_15798,N_14176,N_14762);
nand U15799 (N_15799,N_13651,N_13139);
or U15800 (N_15800,N_14431,N_13501);
nand U15801 (N_15801,N_13631,N_14772);
and U15802 (N_15802,N_14461,N_14075);
or U15803 (N_15803,N_12857,N_13055);
xnor U15804 (N_15804,N_12999,N_13859);
nor U15805 (N_15805,N_13406,N_14140);
nand U15806 (N_15806,N_14241,N_14850);
xnor U15807 (N_15807,N_13039,N_13686);
and U15808 (N_15808,N_13086,N_12808);
xor U15809 (N_15809,N_12749,N_12920);
nor U15810 (N_15810,N_14931,N_13412);
nand U15811 (N_15811,N_12553,N_14760);
and U15812 (N_15812,N_13280,N_14315);
nor U15813 (N_15813,N_14547,N_14232);
and U15814 (N_15814,N_14829,N_14666);
or U15815 (N_15815,N_14159,N_12502);
nand U15816 (N_15816,N_13576,N_12638);
or U15817 (N_15817,N_14773,N_13695);
and U15818 (N_15818,N_14984,N_14385);
and U15819 (N_15819,N_14926,N_14078);
nor U15820 (N_15820,N_14589,N_14609);
or U15821 (N_15821,N_14212,N_14970);
xor U15822 (N_15822,N_14400,N_14507);
nand U15823 (N_15823,N_13987,N_14686);
nand U15824 (N_15824,N_12612,N_14592);
nand U15825 (N_15825,N_12655,N_12738);
or U15826 (N_15826,N_14464,N_13074);
nor U15827 (N_15827,N_14226,N_13755);
and U15828 (N_15828,N_12793,N_12634);
and U15829 (N_15829,N_14836,N_14398);
nand U15830 (N_15830,N_14286,N_13173);
nor U15831 (N_15831,N_13087,N_13674);
xor U15832 (N_15832,N_13386,N_14166);
and U15833 (N_15833,N_14026,N_13905);
nor U15834 (N_15834,N_12953,N_13606);
and U15835 (N_15835,N_12816,N_14975);
nand U15836 (N_15836,N_12526,N_14496);
nor U15837 (N_15837,N_13799,N_14193);
nor U15838 (N_15838,N_13659,N_14184);
nor U15839 (N_15839,N_14623,N_14602);
and U15840 (N_15840,N_13231,N_13333);
and U15841 (N_15841,N_12624,N_12860);
nand U15842 (N_15842,N_13449,N_13414);
or U15843 (N_15843,N_12759,N_13261);
nor U15844 (N_15844,N_12972,N_14745);
xnor U15845 (N_15845,N_14335,N_14710);
nand U15846 (N_15846,N_13499,N_13934);
or U15847 (N_15847,N_14823,N_13128);
or U15848 (N_15848,N_14558,N_13761);
nand U15849 (N_15849,N_14898,N_12629);
nor U15850 (N_15850,N_12965,N_13152);
and U15851 (N_15851,N_13722,N_12631);
or U15852 (N_15852,N_12868,N_13623);
nand U15853 (N_15853,N_12537,N_14310);
and U15854 (N_15854,N_12651,N_13330);
and U15855 (N_15855,N_14994,N_14477);
and U15856 (N_15856,N_13399,N_14812);
xnor U15857 (N_15857,N_14289,N_13411);
nor U15858 (N_15858,N_12913,N_13907);
and U15859 (N_15859,N_12810,N_14068);
or U15860 (N_15860,N_13098,N_13126);
nor U15861 (N_15861,N_14781,N_14856);
and U15862 (N_15862,N_14230,N_13054);
and U15863 (N_15863,N_14132,N_14962);
nor U15864 (N_15864,N_12852,N_12910);
nand U15865 (N_15865,N_12559,N_14565);
and U15866 (N_15866,N_13626,N_12516);
and U15867 (N_15867,N_13220,N_12677);
or U15868 (N_15868,N_12872,N_14998);
or U15869 (N_15869,N_14864,N_14500);
or U15870 (N_15870,N_12945,N_13783);
and U15871 (N_15871,N_12506,N_13939);
or U15872 (N_15872,N_13264,N_13871);
nor U15873 (N_15873,N_13525,N_14514);
nand U15874 (N_15874,N_13716,N_13779);
nand U15875 (N_15875,N_14868,N_13998);
or U15876 (N_15876,N_12529,N_13252);
and U15877 (N_15877,N_13266,N_13065);
and U15878 (N_15878,N_12876,N_13490);
or U15879 (N_15879,N_13937,N_14165);
or U15880 (N_15880,N_13040,N_13902);
nand U15881 (N_15881,N_13154,N_14687);
or U15882 (N_15882,N_13541,N_13809);
nand U15883 (N_15883,N_14652,N_13005);
nand U15884 (N_15884,N_13948,N_13503);
nand U15885 (N_15885,N_14084,N_13813);
nand U15886 (N_15886,N_14197,N_13850);
nand U15887 (N_15887,N_13904,N_12549);
and U15888 (N_15888,N_14797,N_13981);
nand U15889 (N_15889,N_13685,N_14248);
and U15890 (N_15890,N_12813,N_14996);
nand U15891 (N_15891,N_13344,N_13688);
or U15892 (N_15892,N_14768,N_14155);
and U15893 (N_15893,N_13151,N_13602);
nand U15894 (N_15894,N_13487,N_13554);
and U15895 (N_15895,N_14092,N_14319);
nand U15896 (N_15896,N_12724,N_13119);
nor U15897 (N_15897,N_14058,N_14968);
xor U15898 (N_15898,N_13544,N_13392);
nor U15899 (N_15899,N_14209,N_12734);
nand U15900 (N_15900,N_14780,N_13212);
nor U15901 (N_15901,N_12981,N_12871);
nor U15902 (N_15902,N_14703,N_13676);
nor U15903 (N_15903,N_13407,N_14120);
xor U15904 (N_15904,N_14249,N_14629);
or U15905 (N_15905,N_14348,N_14714);
nand U15906 (N_15906,N_14839,N_13150);
and U15907 (N_15907,N_14641,N_12922);
and U15908 (N_15908,N_14333,N_14256);
and U15909 (N_15909,N_13269,N_13299);
nor U15910 (N_15910,N_12695,N_14584);
and U15911 (N_15911,N_13437,N_12554);
nand U15912 (N_15912,N_13710,N_14965);
or U15913 (N_15913,N_14339,N_13801);
or U15914 (N_15914,N_14011,N_12838);
or U15915 (N_15915,N_12790,N_13628);
nor U15916 (N_15916,N_14907,N_14016);
nor U15917 (N_15917,N_12704,N_13085);
nor U15918 (N_15918,N_14146,N_13745);
or U15919 (N_15919,N_13430,N_12591);
or U15920 (N_15920,N_14977,N_13247);
nand U15921 (N_15921,N_14447,N_14139);
or U15922 (N_15922,N_14280,N_13965);
or U15923 (N_15923,N_14748,N_14598);
nand U15924 (N_15924,N_12722,N_13811);
or U15925 (N_15925,N_14524,N_13920);
and U15926 (N_15926,N_13690,N_14614);
and U15927 (N_15927,N_12917,N_12706);
and U15928 (N_15928,N_14495,N_12641);
or U15929 (N_15929,N_13080,N_14612);
nand U15930 (N_15930,N_14943,N_14304);
xor U15931 (N_15931,N_14017,N_14967);
nand U15932 (N_15932,N_14366,N_12916);
and U15933 (N_15933,N_13858,N_12717);
nand U15934 (N_15934,N_14115,N_14066);
and U15935 (N_15935,N_14734,N_14270);
and U15936 (N_15936,N_14410,N_13260);
or U15937 (N_15937,N_12864,N_14946);
xnor U15938 (N_15938,N_12919,N_13297);
xor U15939 (N_15939,N_14805,N_14399);
and U15940 (N_15940,N_14130,N_12865);
or U15941 (N_15941,N_13292,N_14239);
or U15942 (N_15942,N_12557,N_13061);
or U15943 (N_15943,N_13360,N_12599);
and U15944 (N_15944,N_13679,N_12697);
xnor U15945 (N_15945,N_13116,N_13638);
nor U15946 (N_15946,N_12969,N_13728);
or U15947 (N_15947,N_13749,N_12878);
and U15948 (N_15948,N_14693,N_12547);
nand U15949 (N_15949,N_14133,N_12753);
or U15950 (N_15950,N_14746,N_13290);
and U15951 (N_15951,N_13004,N_13696);
or U15952 (N_15952,N_14504,N_13457);
nand U15953 (N_15953,N_14357,N_14731);
nand U15954 (N_15954,N_13335,N_14696);
xnor U15955 (N_15955,N_14732,N_13844);
or U15956 (N_15956,N_14038,N_12863);
xnor U15957 (N_15957,N_14532,N_13209);
and U15958 (N_15958,N_13908,N_13161);
or U15959 (N_15959,N_13263,N_13097);
and U15960 (N_15960,N_14775,N_14761);
nor U15961 (N_15961,N_14048,N_14224);
nand U15962 (N_15962,N_12551,N_13633);
nor U15963 (N_15963,N_13008,N_14809);
or U15964 (N_15964,N_12842,N_14740);
xor U15965 (N_15965,N_14052,N_14285);
xor U15966 (N_15966,N_14537,N_14284);
xor U15967 (N_15967,N_13219,N_12560);
nor U15968 (N_15968,N_14345,N_13480);
or U15969 (N_15969,N_14503,N_13196);
nor U15970 (N_15970,N_13997,N_13520);
nand U15971 (N_15971,N_14089,N_12578);
or U15972 (N_15972,N_13217,N_13581);
nand U15973 (N_15973,N_14782,N_12806);
xor U15974 (N_15974,N_13228,N_14945);
nand U15975 (N_15975,N_12970,N_14116);
nor U15976 (N_15976,N_12746,N_13373);
nor U15977 (N_15977,N_13988,N_14556);
and U15978 (N_15978,N_12541,N_14847);
nor U15979 (N_15979,N_12552,N_12959);
and U15980 (N_15980,N_13918,N_14049);
nand U15981 (N_15981,N_13415,N_14550);
or U15982 (N_15982,N_13115,N_13996);
or U15983 (N_15983,N_14989,N_12527);
nor U15984 (N_15984,N_13855,N_14374);
or U15985 (N_15985,N_13730,N_12680);
or U15986 (N_15986,N_13526,N_13954);
and U15987 (N_15987,N_13574,N_14528);
and U15988 (N_15988,N_13064,N_14966);
nor U15989 (N_15989,N_12758,N_13567);
or U15990 (N_15990,N_12797,N_14213);
and U15991 (N_15991,N_12720,N_13896);
nor U15992 (N_15992,N_12831,N_12615);
nor U15993 (N_15993,N_14237,N_12766);
nand U15994 (N_15994,N_14491,N_14881);
nor U15995 (N_15995,N_13974,N_14835);
nand U15996 (N_15996,N_13257,N_12747);
or U15997 (N_15997,N_13081,N_13781);
nand U15998 (N_15998,N_13751,N_13223);
or U15999 (N_15999,N_14737,N_14910);
or U16000 (N_16000,N_14260,N_13164);
and U16001 (N_16001,N_14138,N_13495);
or U16002 (N_16002,N_14863,N_13020);
or U16003 (N_16003,N_12652,N_12817);
nand U16004 (N_16004,N_13180,N_14449);
or U16005 (N_16005,N_14301,N_12985);
nand U16006 (N_16006,N_12939,N_13977);
or U16007 (N_16007,N_12926,N_12757);
and U16008 (N_16008,N_14605,N_14199);
and U16009 (N_16009,N_14849,N_14207);
xnor U16010 (N_16010,N_13099,N_14991);
nand U16011 (N_16011,N_13062,N_13090);
and U16012 (N_16012,N_14729,N_12562);
xor U16013 (N_16013,N_13834,N_13426);
and U16014 (N_16014,N_13966,N_13448);
nand U16015 (N_16015,N_13646,N_13945);
xnor U16016 (N_16016,N_14796,N_13500);
and U16017 (N_16017,N_13076,N_12500);
nor U16018 (N_16018,N_13401,N_12653);
and U16019 (N_16019,N_14487,N_13309);
or U16020 (N_16020,N_14008,N_14283);
xor U16021 (N_16021,N_13970,N_14419);
xnor U16022 (N_16022,N_14662,N_14390);
nand U16023 (N_16023,N_14803,N_14059);
xor U16024 (N_16024,N_12741,N_13093);
xnor U16025 (N_16025,N_12672,N_14353);
and U16026 (N_16026,N_14261,N_14435);
or U16027 (N_16027,N_14669,N_13348);
nor U16028 (N_16028,N_14250,N_13446);
or U16029 (N_16029,N_14957,N_14051);
and U16030 (N_16030,N_13875,N_13489);
and U16031 (N_16031,N_14670,N_14200);
xnor U16032 (N_16032,N_13458,N_14817);
nand U16033 (N_16033,N_14529,N_13806);
nand U16034 (N_16034,N_12625,N_14841);
nor U16035 (N_16035,N_12514,N_14010);
nor U16036 (N_16036,N_12574,N_13992);
nor U16037 (N_16037,N_13643,N_12632);
and U16038 (N_16038,N_13045,N_13079);
nor U16039 (N_16039,N_14446,N_13184);
and U16040 (N_16040,N_13131,N_13387);
and U16041 (N_16041,N_12764,N_14691);
nand U16042 (N_16042,N_13764,N_14460);
nand U16043 (N_16043,N_12750,N_12524);
nor U16044 (N_16044,N_13204,N_13017);
nor U16045 (N_16045,N_13077,N_12692);
and U16046 (N_16046,N_12544,N_14751);
nand U16047 (N_16047,N_14044,N_14698);
nand U16048 (N_16048,N_13224,N_12841);
and U16049 (N_16049,N_14911,N_14264);
nand U16050 (N_16050,N_13136,N_14581);
and U16051 (N_16051,N_14653,N_13819);
nor U16052 (N_16052,N_12573,N_13694);
or U16053 (N_16053,N_14743,N_13841);
and U16054 (N_16054,N_13274,N_14080);
and U16055 (N_16055,N_13914,N_13951);
and U16056 (N_16056,N_14776,N_14389);
nor U16057 (N_16057,N_14626,N_14308);
nor U16058 (N_16058,N_13952,N_13528);
xnor U16059 (N_16059,N_12525,N_13519);
or U16060 (N_16060,N_13601,N_14088);
and U16061 (N_16061,N_12932,N_13323);
or U16062 (N_16062,N_13453,N_12687);
or U16063 (N_16063,N_13509,N_13163);
nor U16064 (N_16064,N_14637,N_13199);
nand U16065 (N_16065,N_12568,N_12689);
and U16066 (N_16066,N_14347,N_14466);
xor U16067 (N_16067,N_14855,N_13786);
and U16068 (N_16068,N_13025,N_12569);
and U16069 (N_16069,N_14720,N_14810);
or U16070 (N_16070,N_13368,N_14253);
and U16071 (N_16071,N_12586,N_12665);
xor U16072 (N_16072,N_14343,N_14813);
and U16073 (N_16073,N_13731,N_14154);
and U16074 (N_16074,N_13327,N_14378);
and U16075 (N_16075,N_14526,N_14934);
or U16076 (N_16076,N_12827,N_12584);
nand U16077 (N_16077,N_14802,N_13743);
and U16078 (N_16078,N_13608,N_14725);
nand U16079 (N_16079,N_12846,N_14697);
or U16080 (N_16080,N_14870,N_13088);
and U16081 (N_16081,N_12811,N_13985);
nand U16082 (N_16082,N_14268,N_14530);
nand U16083 (N_16083,N_13552,N_14028);
nand U16084 (N_16084,N_14474,N_14682);
or U16085 (N_16085,N_13657,N_13473);
nor U16086 (N_16086,N_14482,N_13477);
nor U16087 (N_16087,N_13129,N_12690);
and U16088 (N_16088,N_14021,N_14037);
xor U16089 (N_16089,N_13645,N_13143);
xnor U16090 (N_16090,N_13078,N_14483);
nor U16091 (N_16091,N_14290,N_13513);
nand U16092 (N_16092,N_13275,N_14208);
nand U16093 (N_16093,N_12671,N_14544);
or U16094 (N_16094,N_13906,N_14369);
or U16095 (N_16095,N_12763,N_14364);
nor U16096 (N_16096,N_14744,N_13719);
and U16097 (N_16097,N_13831,N_14157);
and U16098 (N_16098,N_14894,N_14730);
nor U16099 (N_16099,N_13133,N_12908);
nand U16100 (N_16100,N_12896,N_13958);
nand U16101 (N_16101,N_12774,N_13995);
or U16102 (N_16102,N_13703,N_14194);
and U16103 (N_16103,N_14663,N_12736);
or U16104 (N_16104,N_12906,N_14119);
nand U16105 (N_16105,N_14459,N_13828);
xor U16106 (N_16106,N_12718,N_14196);
nor U16107 (N_16107,N_14896,N_13409);
or U16108 (N_16108,N_14756,N_14557);
nor U16109 (N_16109,N_14097,N_14561);
nor U16110 (N_16110,N_13993,N_14118);
nand U16111 (N_16111,N_13797,N_13341);
or U16112 (N_16112,N_13594,N_12791);
and U16113 (N_16113,N_13157,N_13618);
and U16114 (N_16114,N_14705,N_14539);
nor U16115 (N_16115,N_14632,N_13385);
nor U16116 (N_16116,N_13957,N_12605);
and U16117 (N_16117,N_14727,N_12721);
or U16118 (N_16118,N_13588,N_12923);
nor U16119 (N_16119,N_12982,N_13318);
and U16120 (N_16120,N_12973,N_13324);
nor U16121 (N_16121,N_14876,N_14857);
nand U16122 (N_16122,N_13559,N_13096);
or U16123 (N_16123,N_13352,N_14182);
nor U16124 (N_16124,N_13146,N_13436);
or U16125 (N_16125,N_13014,N_13681);
xnor U16126 (N_16126,N_14604,N_14799);
xor U16127 (N_16127,N_12930,N_12955);
nand U16128 (N_16128,N_14081,N_14340);
nand U16129 (N_16129,N_13510,N_14443);
xor U16130 (N_16130,N_14309,N_12911);
nor U16131 (N_16131,N_13515,N_14407);
nand U16132 (N_16132,N_12957,N_13886);
nand U16133 (N_16133,N_14242,N_14574);
xnor U16134 (N_16134,N_14382,N_13111);
and U16135 (N_16135,N_13599,N_12504);
nor U16136 (N_16136,N_12794,N_12694);
or U16137 (N_16137,N_14938,N_13825);
and U16138 (N_16138,N_13296,N_14153);
nand U16139 (N_16139,N_14147,N_14121);
nand U16140 (N_16140,N_14104,N_14545);
or U16141 (N_16141,N_13474,N_12805);
nor U16142 (N_16142,N_13095,N_14475);
nand U16143 (N_16143,N_14759,N_14266);
nor U16144 (N_16144,N_13410,N_14922);
or U16145 (N_16145,N_13214,N_13289);
or U16146 (N_16146,N_14576,N_14564);
or U16147 (N_16147,N_14948,N_13030);
and U16148 (N_16148,N_14039,N_13882);
nor U16149 (N_16149,N_13517,N_13432);
and U16150 (N_16150,N_14726,N_13211);
nand U16151 (N_16151,N_13979,N_13596);
nand U16152 (N_16152,N_14936,N_14223);
and U16153 (N_16153,N_13950,N_14067);
or U16154 (N_16154,N_14820,N_13069);
and U16155 (N_16155,N_14954,N_14171);
and U16156 (N_16156,N_12693,N_14247);
xnor U16157 (N_16157,N_14472,N_12670);
nor U16158 (N_16158,N_14852,N_14501);
nand U16159 (N_16159,N_13237,N_13758);
nand U16160 (N_16160,N_14123,N_13472);
or U16161 (N_16161,N_14245,N_14401);
and U16162 (N_16162,N_12940,N_14371);
nand U16163 (N_16163,N_14033,N_14516);
nand U16164 (N_16164,N_12660,N_13555);
nand U16165 (N_16165,N_13959,N_12902);
nor U16166 (N_16166,N_14069,N_13766);
nor U16167 (N_16167,N_12998,N_13887);
nor U16168 (N_16168,N_14185,N_13637);
nand U16169 (N_16169,N_13666,N_13094);
nor U16170 (N_16170,N_12847,N_12664);
or U16171 (N_16171,N_12987,N_12948);
or U16172 (N_16172,N_12890,N_13724);
or U16173 (N_16173,N_14777,N_13625);
or U16174 (N_16174,N_14397,N_13114);
xor U16175 (N_16175,N_13784,N_14468);
or U16176 (N_16176,N_14560,N_12735);
nor U16177 (N_16177,N_14297,N_13254);
nor U16178 (N_16178,N_12727,N_13621);
nor U16179 (N_16179,N_14303,N_14959);
and U16180 (N_16180,N_12737,N_13865);
xor U16181 (N_16181,N_13820,N_14901);
xnor U16182 (N_16182,N_13203,N_14627);
or U16183 (N_16183,N_14470,N_14267);
xor U16184 (N_16184,N_14402,N_13746);
nor U16185 (N_16185,N_13354,N_13145);
nand U16186 (N_16186,N_13442,N_14082);
or U16187 (N_16187,N_13359,N_12561);
nand U16188 (N_16188,N_13376,N_14186);
xor U16189 (N_16189,N_12887,N_14749);
and U16190 (N_16190,N_14888,N_13390);
or U16191 (N_16191,N_13137,N_13138);
or U16192 (N_16192,N_12891,N_13649);
xnor U16193 (N_16193,N_14617,N_14109);
nor U16194 (N_16194,N_12824,N_13056);
nand U16195 (N_16195,N_14024,N_13789);
and U16196 (N_16196,N_14587,N_14126);
xor U16197 (N_16197,N_13943,N_13395);
or U16198 (N_16198,N_14518,N_13754);
and U16199 (N_16199,N_13026,N_14271);
and U16200 (N_16200,N_13438,N_13033);
nor U16201 (N_16201,N_13522,N_14610);
and U16202 (N_16202,N_12699,N_14535);
nor U16203 (N_16203,N_13010,N_14880);
xor U16204 (N_16204,N_12628,N_13083);
nor U16205 (N_16205,N_13421,N_12536);
and U16206 (N_16206,N_13768,N_13953);
xnor U16207 (N_16207,N_14972,N_13823);
nand U16208 (N_16208,N_14463,N_12542);
nand U16209 (N_16209,N_14607,N_12540);
nand U16210 (N_16210,N_13734,N_14874);
and U16211 (N_16211,N_12555,N_12623);
and U16212 (N_16212,N_14228,N_13221);
or U16213 (N_16213,N_13179,N_13112);
xnor U16214 (N_16214,N_13234,N_13357);
or U16215 (N_16215,N_13270,N_14444);
nand U16216 (N_16216,N_12711,N_14692);
or U16217 (N_16217,N_14840,N_14867);
xor U16218 (N_16218,N_14394,N_14445);
nor U16219 (N_16219,N_14359,N_14660);
nor U16220 (N_16220,N_13572,N_14784);
nand U16221 (N_16221,N_12968,N_12819);
and U16222 (N_16222,N_12874,N_13654);
or U16223 (N_16223,N_13441,N_13070);
nor U16224 (N_16224,N_12543,N_14094);
or U16225 (N_16225,N_13127,N_13558);
or U16226 (N_16226,N_14050,N_13852);
nor U16227 (N_16227,N_13838,N_12854);
and U16228 (N_16228,N_12768,N_14211);
nand U16229 (N_16229,N_14238,N_14702);
nor U16230 (N_16230,N_14222,N_13271);
xnor U16231 (N_16231,N_13991,N_14927);
and U16232 (N_16232,N_14553,N_12780);
and U16233 (N_16233,N_14511,N_12977);
nand U16234 (N_16234,N_12620,N_14794);
nand U16235 (N_16235,N_12622,N_12590);
nand U16236 (N_16236,N_14631,N_14644);
nor U16237 (N_16237,N_14306,N_12503);
xor U16238 (N_16238,N_12742,N_14671);
or U16239 (N_16239,N_14893,N_12709);
and U16240 (N_16240,N_14467,N_13672);
and U16241 (N_16241,N_13787,N_14622);
nor U16242 (N_16242,N_12710,N_12701);
nor U16243 (N_16243,N_12731,N_13963);
and U16244 (N_16244,N_13612,N_13944);
nand U16245 (N_16245,N_14964,N_14317);
or U16246 (N_16246,N_14002,N_13903);
or U16247 (N_16247,N_13379,N_13893);
or U16248 (N_16248,N_14074,N_14370);
and U16249 (N_16249,N_14942,N_13869);
nand U16250 (N_16250,N_14024,N_12630);
and U16251 (N_16251,N_14547,N_13292);
nor U16252 (N_16252,N_13750,N_14446);
nand U16253 (N_16253,N_14064,N_12987);
nor U16254 (N_16254,N_14727,N_14806);
nor U16255 (N_16255,N_12759,N_14688);
nor U16256 (N_16256,N_14139,N_14816);
nor U16257 (N_16257,N_13433,N_14206);
nand U16258 (N_16258,N_13189,N_13377);
and U16259 (N_16259,N_13495,N_14498);
nor U16260 (N_16260,N_14588,N_14185);
or U16261 (N_16261,N_13993,N_12760);
and U16262 (N_16262,N_14833,N_13391);
nand U16263 (N_16263,N_14999,N_14821);
nand U16264 (N_16264,N_12618,N_13523);
nor U16265 (N_16265,N_14497,N_13601);
xnor U16266 (N_16266,N_13152,N_14169);
and U16267 (N_16267,N_14383,N_13855);
nand U16268 (N_16268,N_14156,N_12955);
or U16269 (N_16269,N_14435,N_13776);
and U16270 (N_16270,N_14403,N_14082);
and U16271 (N_16271,N_13229,N_13219);
or U16272 (N_16272,N_13900,N_12579);
and U16273 (N_16273,N_12752,N_14314);
nor U16274 (N_16274,N_14315,N_14514);
nand U16275 (N_16275,N_12580,N_13599);
xor U16276 (N_16276,N_14343,N_12612);
or U16277 (N_16277,N_13703,N_13934);
nor U16278 (N_16278,N_13952,N_14861);
nor U16279 (N_16279,N_13000,N_12921);
and U16280 (N_16280,N_14809,N_13271);
nand U16281 (N_16281,N_13953,N_12981);
nor U16282 (N_16282,N_14991,N_13161);
and U16283 (N_16283,N_14303,N_13746);
xor U16284 (N_16284,N_14195,N_12645);
or U16285 (N_16285,N_14537,N_14674);
or U16286 (N_16286,N_14155,N_14689);
nand U16287 (N_16287,N_13042,N_12846);
nor U16288 (N_16288,N_14271,N_13118);
nand U16289 (N_16289,N_13623,N_14235);
or U16290 (N_16290,N_14838,N_12528);
nand U16291 (N_16291,N_14236,N_14662);
or U16292 (N_16292,N_13493,N_14383);
and U16293 (N_16293,N_12947,N_14719);
or U16294 (N_16294,N_12711,N_13941);
nor U16295 (N_16295,N_14705,N_13483);
nor U16296 (N_16296,N_14422,N_12989);
nor U16297 (N_16297,N_13847,N_12797);
and U16298 (N_16298,N_14304,N_12556);
nand U16299 (N_16299,N_13581,N_14423);
or U16300 (N_16300,N_13440,N_13691);
xor U16301 (N_16301,N_13916,N_14399);
nand U16302 (N_16302,N_13022,N_14752);
and U16303 (N_16303,N_14543,N_12699);
nand U16304 (N_16304,N_14769,N_14531);
nand U16305 (N_16305,N_14345,N_14246);
nor U16306 (N_16306,N_12641,N_13709);
nand U16307 (N_16307,N_12925,N_12712);
or U16308 (N_16308,N_14169,N_14147);
nor U16309 (N_16309,N_13954,N_14899);
nor U16310 (N_16310,N_12832,N_14886);
nor U16311 (N_16311,N_13084,N_14840);
nor U16312 (N_16312,N_13808,N_13330);
xnor U16313 (N_16313,N_12728,N_13386);
nor U16314 (N_16314,N_13527,N_13565);
and U16315 (N_16315,N_12776,N_14556);
or U16316 (N_16316,N_13320,N_13426);
and U16317 (N_16317,N_13420,N_14363);
and U16318 (N_16318,N_12675,N_13811);
nand U16319 (N_16319,N_13462,N_14118);
nand U16320 (N_16320,N_13923,N_13356);
and U16321 (N_16321,N_14245,N_14546);
and U16322 (N_16322,N_12616,N_12954);
or U16323 (N_16323,N_12552,N_13522);
xnor U16324 (N_16324,N_14727,N_13158);
xor U16325 (N_16325,N_13033,N_13483);
nand U16326 (N_16326,N_13517,N_14855);
nor U16327 (N_16327,N_14567,N_14773);
xor U16328 (N_16328,N_13395,N_13473);
and U16329 (N_16329,N_13502,N_14185);
or U16330 (N_16330,N_13755,N_14841);
or U16331 (N_16331,N_12943,N_14228);
nor U16332 (N_16332,N_14482,N_14696);
nand U16333 (N_16333,N_13906,N_13646);
nor U16334 (N_16334,N_14079,N_14825);
and U16335 (N_16335,N_13329,N_14036);
or U16336 (N_16336,N_14619,N_14984);
nor U16337 (N_16337,N_13590,N_13400);
nor U16338 (N_16338,N_12819,N_12770);
and U16339 (N_16339,N_14925,N_14824);
or U16340 (N_16340,N_13396,N_13846);
nand U16341 (N_16341,N_14027,N_13389);
nor U16342 (N_16342,N_14260,N_13373);
nand U16343 (N_16343,N_13054,N_13559);
nand U16344 (N_16344,N_14442,N_13461);
and U16345 (N_16345,N_14408,N_12911);
or U16346 (N_16346,N_13530,N_12642);
nand U16347 (N_16347,N_14323,N_12582);
nor U16348 (N_16348,N_12567,N_12519);
and U16349 (N_16349,N_13241,N_12702);
nor U16350 (N_16350,N_14274,N_14574);
and U16351 (N_16351,N_12851,N_13003);
and U16352 (N_16352,N_13533,N_12561);
nand U16353 (N_16353,N_13969,N_13038);
nor U16354 (N_16354,N_12813,N_13089);
xnor U16355 (N_16355,N_14671,N_14136);
or U16356 (N_16356,N_14414,N_13124);
xor U16357 (N_16357,N_13784,N_14351);
nand U16358 (N_16358,N_14399,N_13982);
nor U16359 (N_16359,N_13090,N_14439);
nor U16360 (N_16360,N_14860,N_13806);
nand U16361 (N_16361,N_14028,N_13707);
nand U16362 (N_16362,N_13528,N_14589);
xnor U16363 (N_16363,N_14911,N_14731);
and U16364 (N_16364,N_13883,N_14463);
nor U16365 (N_16365,N_12678,N_14116);
xor U16366 (N_16366,N_12753,N_14221);
or U16367 (N_16367,N_13106,N_14453);
nor U16368 (N_16368,N_14479,N_14335);
xnor U16369 (N_16369,N_14504,N_12562);
nand U16370 (N_16370,N_13728,N_12636);
and U16371 (N_16371,N_12731,N_14751);
or U16372 (N_16372,N_13185,N_14758);
nand U16373 (N_16373,N_13184,N_12646);
or U16374 (N_16374,N_12936,N_12850);
nor U16375 (N_16375,N_12780,N_12752);
and U16376 (N_16376,N_14088,N_12742);
nor U16377 (N_16377,N_12740,N_12963);
xor U16378 (N_16378,N_14825,N_13862);
and U16379 (N_16379,N_12842,N_12789);
nand U16380 (N_16380,N_12889,N_13260);
or U16381 (N_16381,N_13983,N_13830);
nor U16382 (N_16382,N_14983,N_13761);
nand U16383 (N_16383,N_14928,N_12687);
nor U16384 (N_16384,N_13548,N_14767);
or U16385 (N_16385,N_14656,N_14467);
nand U16386 (N_16386,N_13210,N_12905);
nand U16387 (N_16387,N_14391,N_14436);
xor U16388 (N_16388,N_12790,N_14523);
and U16389 (N_16389,N_14344,N_13074);
and U16390 (N_16390,N_12559,N_13841);
nand U16391 (N_16391,N_14939,N_14970);
nand U16392 (N_16392,N_13976,N_14728);
nor U16393 (N_16393,N_14709,N_13478);
and U16394 (N_16394,N_14963,N_14124);
and U16395 (N_16395,N_13031,N_13041);
and U16396 (N_16396,N_14385,N_13769);
nor U16397 (N_16397,N_14379,N_14244);
and U16398 (N_16398,N_14177,N_12827);
xnor U16399 (N_16399,N_13443,N_14399);
nor U16400 (N_16400,N_13680,N_13324);
and U16401 (N_16401,N_13087,N_13286);
and U16402 (N_16402,N_14839,N_13076);
nand U16403 (N_16403,N_14184,N_14513);
or U16404 (N_16404,N_13878,N_12595);
nand U16405 (N_16405,N_13318,N_14361);
and U16406 (N_16406,N_13806,N_13111);
nand U16407 (N_16407,N_12957,N_13100);
and U16408 (N_16408,N_14996,N_14165);
or U16409 (N_16409,N_14553,N_14052);
nand U16410 (N_16410,N_13106,N_13543);
or U16411 (N_16411,N_14900,N_13355);
or U16412 (N_16412,N_14615,N_13683);
or U16413 (N_16413,N_14330,N_12980);
and U16414 (N_16414,N_14745,N_12706);
nand U16415 (N_16415,N_13442,N_13927);
nor U16416 (N_16416,N_13850,N_12710);
and U16417 (N_16417,N_14399,N_13060);
nand U16418 (N_16418,N_13792,N_12647);
nor U16419 (N_16419,N_14660,N_13314);
and U16420 (N_16420,N_13385,N_14730);
xor U16421 (N_16421,N_12753,N_14406);
nor U16422 (N_16422,N_14533,N_14405);
and U16423 (N_16423,N_12995,N_13954);
nor U16424 (N_16424,N_13561,N_13004);
nor U16425 (N_16425,N_13387,N_14758);
nand U16426 (N_16426,N_12926,N_12604);
nand U16427 (N_16427,N_12860,N_14646);
or U16428 (N_16428,N_14177,N_12819);
or U16429 (N_16429,N_14980,N_14683);
and U16430 (N_16430,N_14644,N_14094);
nand U16431 (N_16431,N_13829,N_14043);
and U16432 (N_16432,N_12841,N_13534);
nor U16433 (N_16433,N_12838,N_14345);
nand U16434 (N_16434,N_14592,N_13912);
nor U16435 (N_16435,N_14565,N_14174);
xor U16436 (N_16436,N_12878,N_13984);
or U16437 (N_16437,N_13312,N_12942);
and U16438 (N_16438,N_13284,N_12532);
and U16439 (N_16439,N_12696,N_14215);
nand U16440 (N_16440,N_14004,N_13621);
nor U16441 (N_16441,N_12670,N_13703);
and U16442 (N_16442,N_14075,N_12876);
or U16443 (N_16443,N_13706,N_14685);
and U16444 (N_16444,N_12773,N_14253);
and U16445 (N_16445,N_13289,N_13385);
and U16446 (N_16446,N_14193,N_13272);
xor U16447 (N_16447,N_13230,N_14233);
nand U16448 (N_16448,N_13655,N_12970);
xor U16449 (N_16449,N_14951,N_12806);
nor U16450 (N_16450,N_13101,N_13364);
nand U16451 (N_16451,N_12613,N_12551);
nand U16452 (N_16452,N_14935,N_14698);
or U16453 (N_16453,N_14201,N_12815);
nor U16454 (N_16454,N_12516,N_13192);
or U16455 (N_16455,N_13383,N_14583);
nand U16456 (N_16456,N_12540,N_14098);
nor U16457 (N_16457,N_14603,N_13505);
nor U16458 (N_16458,N_13374,N_14175);
or U16459 (N_16459,N_13657,N_13415);
and U16460 (N_16460,N_13137,N_12863);
nand U16461 (N_16461,N_13692,N_13343);
nor U16462 (N_16462,N_12524,N_13852);
and U16463 (N_16463,N_14220,N_12752);
or U16464 (N_16464,N_13445,N_13271);
and U16465 (N_16465,N_13112,N_13630);
nand U16466 (N_16466,N_14864,N_13264);
nand U16467 (N_16467,N_14352,N_14472);
nand U16468 (N_16468,N_14854,N_14183);
nand U16469 (N_16469,N_14214,N_14141);
nand U16470 (N_16470,N_13200,N_14432);
nor U16471 (N_16471,N_14593,N_12637);
nor U16472 (N_16472,N_13713,N_14124);
and U16473 (N_16473,N_14546,N_13527);
nor U16474 (N_16474,N_13179,N_14057);
nand U16475 (N_16475,N_14740,N_13229);
and U16476 (N_16476,N_13469,N_14097);
nor U16477 (N_16477,N_13227,N_14489);
nand U16478 (N_16478,N_14160,N_14928);
xnor U16479 (N_16479,N_13328,N_14561);
or U16480 (N_16480,N_12781,N_13150);
nor U16481 (N_16481,N_13245,N_14523);
and U16482 (N_16482,N_12698,N_13207);
or U16483 (N_16483,N_13144,N_12676);
and U16484 (N_16484,N_12911,N_14525);
and U16485 (N_16485,N_12723,N_12791);
or U16486 (N_16486,N_14735,N_14986);
nor U16487 (N_16487,N_13223,N_14333);
and U16488 (N_16488,N_14351,N_12996);
or U16489 (N_16489,N_13122,N_14515);
nor U16490 (N_16490,N_13683,N_14709);
nand U16491 (N_16491,N_13315,N_13982);
or U16492 (N_16492,N_14016,N_12952);
and U16493 (N_16493,N_12954,N_13324);
and U16494 (N_16494,N_13835,N_14680);
and U16495 (N_16495,N_13909,N_14871);
or U16496 (N_16496,N_12648,N_12646);
or U16497 (N_16497,N_13312,N_14726);
or U16498 (N_16498,N_14983,N_13749);
nor U16499 (N_16499,N_14804,N_14441);
or U16500 (N_16500,N_13937,N_14334);
or U16501 (N_16501,N_14833,N_12716);
or U16502 (N_16502,N_12631,N_12852);
nand U16503 (N_16503,N_14078,N_14922);
nand U16504 (N_16504,N_12591,N_14122);
nor U16505 (N_16505,N_13105,N_14649);
nand U16506 (N_16506,N_12826,N_12515);
and U16507 (N_16507,N_13977,N_13786);
and U16508 (N_16508,N_14567,N_14921);
and U16509 (N_16509,N_13604,N_14669);
nand U16510 (N_16510,N_14555,N_13477);
nor U16511 (N_16511,N_12584,N_13247);
and U16512 (N_16512,N_13447,N_12786);
nor U16513 (N_16513,N_13939,N_14003);
or U16514 (N_16514,N_13217,N_14698);
and U16515 (N_16515,N_13159,N_14065);
or U16516 (N_16516,N_12759,N_14419);
nor U16517 (N_16517,N_14431,N_13175);
or U16518 (N_16518,N_13851,N_12746);
or U16519 (N_16519,N_14060,N_12560);
or U16520 (N_16520,N_14874,N_13625);
and U16521 (N_16521,N_12781,N_13469);
and U16522 (N_16522,N_13159,N_12804);
xnor U16523 (N_16523,N_13037,N_14595);
nand U16524 (N_16524,N_14151,N_14676);
or U16525 (N_16525,N_13045,N_13005);
nand U16526 (N_16526,N_14702,N_14679);
nor U16527 (N_16527,N_12579,N_13778);
or U16528 (N_16528,N_14132,N_12893);
nand U16529 (N_16529,N_12909,N_13181);
or U16530 (N_16530,N_14251,N_14651);
xor U16531 (N_16531,N_14814,N_13743);
and U16532 (N_16532,N_13990,N_12658);
nor U16533 (N_16533,N_14973,N_13020);
nor U16534 (N_16534,N_12564,N_13938);
nand U16535 (N_16535,N_14231,N_14722);
nand U16536 (N_16536,N_14077,N_12596);
nor U16537 (N_16537,N_12703,N_13656);
or U16538 (N_16538,N_13147,N_12900);
nand U16539 (N_16539,N_12906,N_14926);
nand U16540 (N_16540,N_14772,N_13514);
nor U16541 (N_16541,N_14386,N_13360);
or U16542 (N_16542,N_13486,N_14968);
and U16543 (N_16543,N_14927,N_14278);
nand U16544 (N_16544,N_12911,N_13235);
nor U16545 (N_16545,N_12940,N_13929);
and U16546 (N_16546,N_14512,N_12527);
xnor U16547 (N_16547,N_13280,N_14124);
and U16548 (N_16548,N_13850,N_14587);
and U16549 (N_16549,N_12713,N_13307);
and U16550 (N_16550,N_13716,N_13611);
nand U16551 (N_16551,N_12649,N_13028);
or U16552 (N_16552,N_14692,N_12665);
or U16553 (N_16553,N_13201,N_13186);
nor U16554 (N_16554,N_14174,N_14757);
nand U16555 (N_16555,N_13266,N_13593);
nand U16556 (N_16556,N_13880,N_14329);
and U16557 (N_16557,N_13932,N_13763);
or U16558 (N_16558,N_14343,N_14986);
and U16559 (N_16559,N_13333,N_14986);
or U16560 (N_16560,N_12601,N_14677);
nand U16561 (N_16561,N_13389,N_14383);
and U16562 (N_16562,N_14528,N_14531);
or U16563 (N_16563,N_13980,N_14712);
nand U16564 (N_16564,N_12682,N_13846);
nor U16565 (N_16565,N_14383,N_13336);
nand U16566 (N_16566,N_13577,N_14895);
and U16567 (N_16567,N_14771,N_14611);
and U16568 (N_16568,N_12744,N_12892);
xor U16569 (N_16569,N_13246,N_13640);
nand U16570 (N_16570,N_12592,N_14544);
nor U16571 (N_16571,N_13153,N_13445);
nor U16572 (N_16572,N_14387,N_14805);
and U16573 (N_16573,N_14343,N_13262);
and U16574 (N_16574,N_13465,N_14651);
xor U16575 (N_16575,N_12953,N_13191);
or U16576 (N_16576,N_12734,N_13640);
xnor U16577 (N_16577,N_12803,N_14399);
nor U16578 (N_16578,N_12580,N_13829);
and U16579 (N_16579,N_14843,N_14511);
nor U16580 (N_16580,N_14895,N_13053);
or U16581 (N_16581,N_13570,N_14651);
nor U16582 (N_16582,N_14734,N_13775);
nor U16583 (N_16583,N_14613,N_13976);
or U16584 (N_16584,N_13550,N_14193);
nor U16585 (N_16585,N_14731,N_14034);
nor U16586 (N_16586,N_14955,N_12951);
and U16587 (N_16587,N_13515,N_13249);
nand U16588 (N_16588,N_13802,N_14608);
nor U16589 (N_16589,N_13505,N_14102);
or U16590 (N_16590,N_14702,N_14651);
xor U16591 (N_16591,N_14063,N_13516);
xnor U16592 (N_16592,N_14598,N_12749);
or U16593 (N_16593,N_13090,N_13236);
or U16594 (N_16594,N_14462,N_13721);
nor U16595 (N_16595,N_12797,N_12910);
nand U16596 (N_16596,N_14744,N_12669);
nand U16597 (N_16597,N_14391,N_13767);
or U16598 (N_16598,N_13853,N_14836);
nand U16599 (N_16599,N_12844,N_13168);
and U16600 (N_16600,N_13485,N_13545);
and U16601 (N_16601,N_13618,N_13609);
xnor U16602 (N_16602,N_14891,N_12879);
or U16603 (N_16603,N_14907,N_12851);
and U16604 (N_16604,N_14926,N_12612);
and U16605 (N_16605,N_13247,N_12514);
nor U16606 (N_16606,N_13364,N_14132);
and U16607 (N_16607,N_14953,N_13473);
nor U16608 (N_16608,N_12566,N_13137);
nor U16609 (N_16609,N_12547,N_12677);
or U16610 (N_16610,N_14775,N_13085);
or U16611 (N_16611,N_12943,N_13064);
and U16612 (N_16612,N_12982,N_13853);
and U16613 (N_16613,N_13013,N_14400);
or U16614 (N_16614,N_13149,N_12923);
or U16615 (N_16615,N_14229,N_13597);
nor U16616 (N_16616,N_14944,N_12932);
or U16617 (N_16617,N_14304,N_14730);
or U16618 (N_16618,N_13901,N_13262);
nor U16619 (N_16619,N_12637,N_14372);
or U16620 (N_16620,N_14159,N_13022);
nand U16621 (N_16621,N_14312,N_12544);
nand U16622 (N_16622,N_13184,N_14080);
nor U16623 (N_16623,N_13453,N_13676);
nor U16624 (N_16624,N_13815,N_12762);
or U16625 (N_16625,N_12982,N_13930);
xor U16626 (N_16626,N_12548,N_14830);
or U16627 (N_16627,N_13532,N_14132);
or U16628 (N_16628,N_13560,N_14199);
nand U16629 (N_16629,N_13302,N_14738);
xnor U16630 (N_16630,N_12954,N_13288);
nor U16631 (N_16631,N_14414,N_13214);
nand U16632 (N_16632,N_14849,N_13953);
and U16633 (N_16633,N_13472,N_13285);
nor U16634 (N_16634,N_12882,N_13303);
nor U16635 (N_16635,N_14677,N_14308);
nor U16636 (N_16636,N_13466,N_14205);
and U16637 (N_16637,N_14081,N_14020);
xor U16638 (N_16638,N_13504,N_14554);
or U16639 (N_16639,N_14024,N_12546);
xor U16640 (N_16640,N_13138,N_13806);
xor U16641 (N_16641,N_13359,N_13107);
and U16642 (N_16642,N_13949,N_14884);
or U16643 (N_16643,N_12918,N_14920);
nand U16644 (N_16644,N_12803,N_12959);
or U16645 (N_16645,N_12587,N_14459);
or U16646 (N_16646,N_14914,N_12562);
nand U16647 (N_16647,N_14100,N_14924);
xor U16648 (N_16648,N_13809,N_13397);
nor U16649 (N_16649,N_13171,N_12793);
nand U16650 (N_16650,N_14243,N_13000);
and U16651 (N_16651,N_13620,N_14825);
and U16652 (N_16652,N_13088,N_13844);
and U16653 (N_16653,N_13224,N_13007);
and U16654 (N_16654,N_13855,N_13544);
nor U16655 (N_16655,N_14061,N_14885);
nand U16656 (N_16656,N_13243,N_13778);
and U16657 (N_16657,N_13622,N_12844);
nand U16658 (N_16658,N_13289,N_13033);
or U16659 (N_16659,N_12751,N_14828);
nand U16660 (N_16660,N_13760,N_14742);
nand U16661 (N_16661,N_14922,N_13941);
or U16662 (N_16662,N_13156,N_14785);
and U16663 (N_16663,N_14073,N_14119);
xor U16664 (N_16664,N_13023,N_14731);
and U16665 (N_16665,N_14253,N_14594);
or U16666 (N_16666,N_14371,N_13675);
or U16667 (N_16667,N_13364,N_14509);
nor U16668 (N_16668,N_13543,N_14590);
and U16669 (N_16669,N_13628,N_14589);
nor U16670 (N_16670,N_12659,N_13986);
nor U16671 (N_16671,N_13189,N_14138);
nand U16672 (N_16672,N_14803,N_13897);
nor U16673 (N_16673,N_13543,N_14388);
or U16674 (N_16674,N_14779,N_13546);
and U16675 (N_16675,N_12763,N_14257);
nor U16676 (N_16676,N_14666,N_12848);
xor U16677 (N_16677,N_13690,N_12611);
xnor U16678 (N_16678,N_14357,N_14256);
nand U16679 (N_16679,N_14952,N_13299);
or U16680 (N_16680,N_14877,N_14836);
nand U16681 (N_16681,N_12844,N_13735);
nand U16682 (N_16682,N_12541,N_12581);
and U16683 (N_16683,N_13973,N_13723);
nand U16684 (N_16684,N_14122,N_14847);
nand U16685 (N_16685,N_14666,N_13728);
and U16686 (N_16686,N_13937,N_13124);
or U16687 (N_16687,N_13048,N_14960);
nand U16688 (N_16688,N_13304,N_14344);
xnor U16689 (N_16689,N_14441,N_14194);
or U16690 (N_16690,N_14271,N_13439);
and U16691 (N_16691,N_13553,N_14036);
xor U16692 (N_16692,N_13089,N_12682);
xor U16693 (N_16693,N_12766,N_12959);
or U16694 (N_16694,N_14020,N_13200);
and U16695 (N_16695,N_13610,N_13036);
or U16696 (N_16696,N_12793,N_14332);
nor U16697 (N_16697,N_14303,N_14617);
xnor U16698 (N_16698,N_13878,N_12707);
nor U16699 (N_16699,N_13528,N_13977);
and U16700 (N_16700,N_14099,N_12992);
and U16701 (N_16701,N_13329,N_12521);
and U16702 (N_16702,N_13951,N_13818);
nor U16703 (N_16703,N_12710,N_13067);
or U16704 (N_16704,N_13375,N_14220);
and U16705 (N_16705,N_12816,N_12741);
and U16706 (N_16706,N_13854,N_14096);
nor U16707 (N_16707,N_14969,N_12810);
and U16708 (N_16708,N_13322,N_13617);
nand U16709 (N_16709,N_13122,N_13509);
and U16710 (N_16710,N_14597,N_13484);
or U16711 (N_16711,N_14921,N_14047);
or U16712 (N_16712,N_14415,N_13554);
nand U16713 (N_16713,N_12629,N_13365);
nand U16714 (N_16714,N_13851,N_13251);
or U16715 (N_16715,N_13450,N_14697);
nor U16716 (N_16716,N_14376,N_14189);
nor U16717 (N_16717,N_14377,N_13731);
nor U16718 (N_16718,N_12712,N_12966);
nand U16719 (N_16719,N_14913,N_13243);
or U16720 (N_16720,N_14587,N_14996);
nand U16721 (N_16721,N_14430,N_13654);
nor U16722 (N_16722,N_12933,N_14781);
or U16723 (N_16723,N_12780,N_14690);
nor U16724 (N_16724,N_14880,N_14079);
or U16725 (N_16725,N_14899,N_14296);
nand U16726 (N_16726,N_13537,N_14250);
or U16727 (N_16727,N_12520,N_14557);
nor U16728 (N_16728,N_14586,N_14013);
nand U16729 (N_16729,N_14085,N_14628);
and U16730 (N_16730,N_14338,N_13288);
and U16731 (N_16731,N_12728,N_14050);
nand U16732 (N_16732,N_14903,N_14359);
nand U16733 (N_16733,N_14866,N_13311);
or U16734 (N_16734,N_13658,N_14561);
and U16735 (N_16735,N_12995,N_14703);
or U16736 (N_16736,N_14684,N_14160);
nand U16737 (N_16737,N_14090,N_13199);
and U16738 (N_16738,N_14416,N_13771);
nand U16739 (N_16739,N_14087,N_14642);
nand U16740 (N_16740,N_13775,N_12653);
or U16741 (N_16741,N_14448,N_12827);
xor U16742 (N_16742,N_13913,N_12590);
or U16743 (N_16743,N_13773,N_14769);
nand U16744 (N_16744,N_14179,N_13670);
and U16745 (N_16745,N_13732,N_13425);
nor U16746 (N_16746,N_12909,N_14928);
and U16747 (N_16747,N_12951,N_13863);
and U16748 (N_16748,N_14915,N_13392);
or U16749 (N_16749,N_14132,N_13265);
nand U16750 (N_16750,N_14011,N_12920);
nor U16751 (N_16751,N_14239,N_12767);
nand U16752 (N_16752,N_12782,N_12972);
nand U16753 (N_16753,N_12620,N_14699);
nand U16754 (N_16754,N_14641,N_14034);
nand U16755 (N_16755,N_14076,N_12629);
nor U16756 (N_16756,N_13157,N_12970);
nand U16757 (N_16757,N_12525,N_14793);
nand U16758 (N_16758,N_14940,N_14076);
nand U16759 (N_16759,N_13475,N_13232);
xnor U16760 (N_16760,N_14504,N_14976);
nand U16761 (N_16761,N_14303,N_14402);
or U16762 (N_16762,N_13041,N_14762);
or U16763 (N_16763,N_14389,N_12704);
and U16764 (N_16764,N_13258,N_14207);
and U16765 (N_16765,N_14170,N_13849);
nand U16766 (N_16766,N_12739,N_14195);
or U16767 (N_16767,N_13496,N_13803);
xnor U16768 (N_16768,N_13669,N_13184);
or U16769 (N_16769,N_13377,N_14410);
nor U16770 (N_16770,N_14982,N_13355);
xor U16771 (N_16771,N_13073,N_14647);
and U16772 (N_16772,N_13728,N_13189);
nand U16773 (N_16773,N_12761,N_13098);
or U16774 (N_16774,N_14736,N_12652);
nor U16775 (N_16775,N_13876,N_12534);
or U16776 (N_16776,N_13658,N_14145);
xnor U16777 (N_16777,N_14469,N_13853);
and U16778 (N_16778,N_13391,N_12823);
or U16779 (N_16779,N_14018,N_13589);
and U16780 (N_16780,N_14162,N_13944);
nand U16781 (N_16781,N_14582,N_13263);
or U16782 (N_16782,N_14330,N_13801);
and U16783 (N_16783,N_14995,N_14045);
nand U16784 (N_16784,N_12542,N_13927);
or U16785 (N_16785,N_13621,N_12763);
nor U16786 (N_16786,N_13995,N_14542);
and U16787 (N_16787,N_13068,N_14741);
nand U16788 (N_16788,N_12517,N_14927);
nor U16789 (N_16789,N_14834,N_14712);
and U16790 (N_16790,N_14265,N_13150);
and U16791 (N_16791,N_13415,N_14061);
xor U16792 (N_16792,N_13882,N_12749);
nand U16793 (N_16793,N_14040,N_12608);
nor U16794 (N_16794,N_14609,N_13870);
nand U16795 (N_16795,N_12636,N_14829);
nand U16796 (N_16796,N_14127,N_12982);
or U16797 (N_16797,N_14791,N_13776);
nand U16798 (N_16798,N_14390,N_12652);
and U16799 (N_16799,N_14128,N_12946);
xor U16800 (N_16800,N_13199,N_13737);
nand U16801 (N_16801,N_12707,N_12888);
nand U16802 (N_16802,N_14516,N_13022);
and U16803 (N_16803,N_13339,N_13032);
and U16804 (N_16804,N_14411,N_13932);
nand U16805 (N_16805,N_14373,N_13906);
nand U16806 (N_16806,N_12718,N_12930);
and U16807 (N_16807,N_12586,N_14557);
or U16808 (N_16808,N_13185,N_12960);
and U16809 (N_16809,N_12824,N_13759);
nand U16810 (N_16810,N_13892,N_12819);
or U16811 (N_16811,N_12582,N_12705);
nand U16812 (N_16812,N_12577,N_12703);
nand U16813 (N_16813,N_13324,N_13975);
and U16814 (N_16814,N_12667,N_13319);
or U16815 (N_16815,N_13739,N_14624);
and U16816 (N_16816,N_13007,N_13488);
or U16817 (N_16817,N_13523,N_14019);
nor U16818 (N_16818,N_12739,N_12839);
or U16819 (N_16819,N_14621,N_13021);
and U16820 (N_16820,N_13986,N_13301);
xnor U16821 (N_16821,N_13890,N_12581);
nand U16822 (N_16822,N_13774,N_14265);
and U16823 (N_16823,N_14964,N_13152);
nand U16824 (N_16824,N_14335,N_13681);
or U16825 (N_16825,N_14321,N_13968);
xnor U16826 (N_16826,N_14128,N_13183);
and U16827 (N_16827,N_14972,N_14204);
xnor U16828 (N_16828,N_14192,N_12552);
nor U16829 (N_16829,N_14811,N_14211);
nor U16830 (N_16830,N_14915,N_13069);
and U16831 (N_16831,N_12657,N_14546);
and U16832 (N_16832,N_13584,N_14486);
or U16833 (N_16833,N_13111,N_12604);
and U16834 (N_16834,N_13970,N_13652);
nor U16835 (N_16835,N_13070,N_14521);
nor U16836 (N_16836,N_12683,N_13626);
xor U16837 (N_16837,N_14458,N_14668);
nand U16838 (N_16838,N_14106,N_12603);
or U16839 (N_16839,N_13440,N_13486);
and U16840 (N_16840,N_12745,N_12648);
nand U16841 (N_16841,N_13976,N_13206);
and U16842 (N_16842,N_13361,N_13554);
nand U16843 (N_16843,N_13156,N_14316);
or U16844 (N_16844,N_13745,N_14289);
xnor U16845 (N_16845,N_13216,N_13774);
and U16846 (N_16846,N_12732,N_14379);
nor U16847 (N_16847,N_13908,N_14634);
nand U16848 (N_16848,N_14498,N_13826);
nand U16849 (N_16849,N_13930,N_14886);
or U16850 (N_16850,N_13891,N_14532);
nand U16851 (N_16851,N_12879,N_12595);
or U16852 (N_16852,N_12555,N_14476);
or U16853 (N_16853,N_14011,N_14982);
nor U16854 (N_16854,N_12720,N_13492);
and U16855 (N_16855,N_14252,N_13593);
and U16856 (N_16856,N_14995,N_12553);
xnor U16857 (N_16857,N_14327,N_12735);
and U16858 (N_16858,N_14992,N_14892);
or U16859 (N_16859,N_14058,N_14162);
nand U16860 (N_16860,N_13424,N_14067);
and U16861 (N_16861,N_12739,N_13719);
or U16862 (N_16862,N_13780,N_13999);
and U16863 (N_16863,N_14400,N_14007);
and U16864 (N_16864,N_14962,N_12777);
nand U16865 (N_16865,N_13091,N_13661);
nand U16866 (N_16866,N_13826,N_14968);
nand U16867 (N_16867,N_12612,N_14314);
and U16868 (N_16868,N_14258,N_14874);
xor U16869 (N_16869,N_13343,N_14711);
nand U16870 (N_16870,N_13961,N_14205);
and U16871 (N_16871,N_14441,N_14995);
nand U16872 (N_16872,N_14565,N_14537);
and U16873 (N_16873,N_14975,N_12650);
and U16874 (N_16874,N_14018,N_13649);
nand U16875 (N_16875,N_14913,N_12515);
and U16876 (N_16876,N_12923,N_13404);
nor U16877 (N_16877,N_14563,N_13869);
or U16878 (N_16878,N_12700,N_13717);
or U16879 (N_16879,N_13820,N_14814);
nand U16880 (N_16880,N_14605,N_13924);
nor U16881 (N_16881,N_13102,N_14978);
or U16882 (N_16882,N_13855,N_12962);
and U16883 (N_16883,N_14074,N_12606);
and U16884 (N_16884,N_13151,N_13034);
or U16885 (N_16885,N_13791,N_13620);
or U16886 (N_16886,N_14459,N_13619);
nand U16887 (N_16887,N_14575,N_14498);
xnor U16888 (N_16888,N_13360,N_12865);
nor U16889 (N_16889,N_13411,N_13607);
or U16890 (N_16890,N_14605,N_14332);
nor U16891 (N_16891,N_13347,N_13320);
and U16892 (N_16892,N_12995,N_13143);
or U16893 (N_16893,N_13673,N_14721);
or U16894 (N_16894,N_12902,N_13239);
xnor U16895 (N_16895,N_14689,N_13112);
nor U16896 (N_16896,N_14692,N_13712);
xor U16897 (N_16897,N_14744,N_12934);
or U16898 (N_16898,N_13561,N_14914);
nand U16899 (N_16899,N_14677,N_14043);
nand U16900 (N_16900,N_14947,N_14343);
xnor U16901 (N_16901,N_14134,N_13421);
xor U16902 (N_16902,N_12721,N_13284);
or U16903 (N_16903,N_14084,N_14622);
nor U16904 (N_16904,N_14111,N_14540);
nor U16905 (N_16905,N_14498,N_12759);
nand U16906 (N_16906,N_13286,N_12777);
nand U16907 (N_16907,N_14072,N_14062);
and U16908 (N_16908,N_14474,N_14840);
and U16909 (N_16909,N_12908,N_14392);
and U16910 (N_16910,N_14561,N_14342);
or U16911 (N_16911,N_14597,N_14828);
and U16912 (N_16912,N_13586,N_13676);
nand U16913 (N_16913,N_12890,N_14834);
nand U16914 (N_16914,N_14282,N_12634);
nor U16915 (N_16915,N_14584,N_14599);
nand U16916 (N_16916,N_12805,N_14392);
xor U16917 (N_16917,N_14443,N_14405);
nor U16918 (N_16918,N_12791,N_12875);
nor U16919 (N_16919,N_13529,N_14879);
or U16920 (N_16920,N_12671,N_14322);
nand U16921 (N_16921,N_14503,N_14565);
or U16922 (N_16922,N_14118,N_14376);
or U16923 (N_16923,N_13019,N_14405);
nor U16924 (N_16924,N_13004,N_14910);
and U16925 (N_16925,N_14750,N_14397);
or U16926 (N_16926,N_12931,N_13805);
and U16927 (N_16927,N_12550,N_12828);
and U16928 (N_16928,N_13266,N_13059);
or U16929 (N_16929,N_14687,N_14682);
and U16930 (N_16930,N_13626,N_14917);
or U16931 (N_16931,N_13908,N_13928);
and U16932 (N_16932,N_13343,N_12583);
nand U16933 (N_16933,N_13836,N_13127);
xnor U16934 (N_16934,N_14040,N_12935);
nor U16935 (N_16935,N_12962,N_12990);
and U16936 (N_16936,N_12725,N_13934);
and U16937 (N_16937,N_14950,N_12830);
nor U16938 (N_16938,N_14034,N_14369);
nand U16939 (N_16939,N_13435,N_13314);
nor U16940 (N_16940,N_13350,N_13035);
xnor U16941 (N_16941,N_13968,N_14968);
and U16942 (N_16942,N_14161,N_13912);
or U16943 (N_16943,N_13914,N_13994);
nor U16944 (N_16944,N_13967,N_14447);
or U16945 (N_16945,N_13701,N_12585);
nor U16946 (N_16946,N_14957,N_14272);
nand U16947 (N_16947,N_13015,N_14702);
and U16948 (N_16948,N_14584,N_13139);
nor U16949 (N_16949,N_13050,N_14265);
nand U16950 (N_16950,N_12916,N_13855);
or U16951 (N_16951,N_12940,N_14515);
xor U16952 (N_16952,N_13900,N_12762);
xnor U16953 (N_16953,N_13682,N_12962);
or U16954 (N_16954,N_13741,N_14358);
and U16955 (N_16955,N_14566,N_12697);
nand U16956 (N_16956,N_14188,N_14254);
or U16957 (N_16957,N_13367,N_13385);
nand U16958 (N_16958,N_13168,N_14442);
and U16959 (N_16959,N_13736,N_13721);
nor U16960 (N_16960,N_14799,N_13457);
nor U16961 (N_16961,N_12847,N_12562);
nand U16962 (N_16962,N_14493,N_12630);
nand U16963 (N_16963,N_13909,N_12802);
nand U16964 (N_16964,N_13639,N_14223);
xor U16965 (N_16965,N_12981,N_13713);
nor U16966 (N_16966,N_13678,N_13312);
xnor U16967 (N_16967,N_13458,N_12932);
nor U16968 (N_16968,N_14828,N_14160);
or U16969 (N_16969,N_13144,N_14071);
nand U16970 (N_16970,N_14116,N_14006);
nand U16971 (N_16971,N_14117,N_12700);
and U16972 (N_16972,N_13015,N_12988);
and U16973 (N_16973,N_14156,N_13971);
or U16974 (N_16974,N_13600,N_12860);
or U16975 (N_16975,N_13441,N_14585);
nor U16976 (N_16976,N_13237,N_12845);
or U16977 (N_16977,N_12596,N_14304);
nand U16978 (N_16978,N_13868,N_14407);
and U16979 (N_16979,N_14691,N_14782);
xor U16980 (N_16980,N_13798,N_12593);
or U16981 (N_16981,N_13836,N_14772);
nor U16982 (N_16982,N_14457,N_13995);
nand U16983 (N_16983,N_14612,N_13760);
and U16984 (N_16984,N_13700,N_14055);
or U16985 (N_16985,N_12543,N_14662);
nor U16986 (N_16986,N_13090,N_14871);
xnor U16987 (N_16987,N_13192,N_12546);
nor U16988 (N_16988,N_14633,N_13072);
or U16989 (N_16989,N_14037,N_14847);
nand U16990 (N_16990,N_13778,N_14412);
or U16991 (N_16991,N_13660,N_12940);
nor U16992 (N_16992,N_12582,N_13950);
xor U16993 (N_16993,N_12727,N_14544);
or U16994 (N_16994,N_14337,N_14954);
xor U16995 (N_16995,N_14871,N_14231);
and U16996 (N_16996,N_14170,N_14173);
nor U16997 (N_16997,N_12857,N_12779);
and U16998 (N_16998,N_12788,N_14470);
or U16999 (N_16999,N_14760,N_12755);
and U17000 (N_17000,N_12503,N_13970);
nand U17001 (N_17001,N_12745,N_14353);
and U17002 (N_17002,N_14133,N_12532);
nand U17003 (N_17003,N_14838,N_13231);
xor U17004 (N_17004,N_13990,N_14636);
or U17005 (N_17005,N_13116,N_13817);
and U17006 (N_17006,N_14090,N_13202);
xnor U17007 (N_17007,N_13293,N_12992);
or U17008 (N_17008,N_13656,N_13947);
xnor U17009 (N_17009,N_13890,N_14831);
and U17010 (N_17010,N_12610,N_13907);
nand U17011 (N_17011,N_14488,N_13368);
or U17012 (N_17012,N_13143,N_13324);
nand U17013 (N_17013,N_14481,N_13676);
or U17014 (N_17014,N_14347,N_14786);
xor U17015 (N_17015,N_14911,N_13519);
nand U17016 (N_17016,N_13363,N_12712);
and U17017 (N_17017,N_12937,N_13050);
xnor U17018 (N_17018,N_14825,N_12843);
and U17019 (N_17019,N_13350,N_14507);
or U17020 (N_17020,N_12916,N_14206);
or U17021 (N_17021,N_13638,N_14259);
nand U17022 (N_17022,N_13289,N_12801);
xnor U17023 (N_17023,N_14552,N_12663);
xnor U17024 (N_17024,N_13436,N_14671);
nor U17025 (N_17025,N_14622,N_14347);
nand U17026 (N_17026,N_13867,N_13723);
nor U17027 (N_17027,N_13740,N_14581);
and U17028 (N_17028,N_13267,N_14391);
or U17029 (N_17029,N_14676,N_14035);
nor U17030 (N_17030,N_13209,N_14990);
nor U17031 (N_17031,N_13636,N_13994);
nand U17032 (N_17032,N_13195,N_14098);
or U17033 (N_17033,N_14027,N_14889);
nor U17034 (N_17034,N_14748,N_14784);
nor U17035 (N_17035,N_14066,N_14310);
xor U17036 (N_17036,N_14441,N_12970);
xor U17037 (N_17037,N_14460,N_13872);
or U17038 (N_17038,N_13416,N_13766);
nor U17039 (N_17039,N_14997,N_12867);
xnor U17040 (N_17040,N_12680,N_13146);
or U17041 (N_17041,N_13192,N_13125);
and U17042 (N_17042,N_14153,N_14547);
xor U17043 (N_17043,N_13770,N_13014);
nor U17044 (N_17044,N_14600,N_12937);
nand U17045 (N_17045,N_13631,N_12674);
nand U17046 (N_17046,N_12800,N_13994);
nor U17047 (N_17047,N_13302,N_13060);
nor U17048 (N_17048,N_13920,N_13887);
nand U17049 (N_17049,N_14863,N_12933);
and U17050 (N_17050,N_14176,N_13442);
nor U17051 (N_17051,N_12893,N_13717);
or U17052 (N_17052,N_13498,N_13364);
nand U17053 (N_17053,N_14357,N_14271);
xor U17054 (N_17054,N_13594,N_13235);
nand U17055 (N_17055,N_14720,N_14097);
nor U17056 (N_17056,N_14433,N_13039);
and U17057 (N_17057,N_12599,N_14247);
and U17058 (N_17058,N_12789,N_14467);
nand U17059 (N_17059,N_12842,N_14005);
nand U17060 (N_17060,N_12919,N_14865);
nand U17061 (N_17061,N_12528,N_14496);
or U17062 (N_17062,N_14480,N_14858);
or U17063 (N_17063,N_13362,N_13085);
or U17064 (N_17064,N_12605,N_14702);
xnor U17065 (N_17065,N_13509,N_13732);
nor U17066 (N_17066,N_12706,N_14851);
nor U17067 (N_17067,N_13838,N_14725);
or U17068 (N_17068,N_13300,N_14311);
nor U17069 (N_17069,N_13012,N_12523);
or U17070 (N_17070,N_14737,N_14048);
and U17071 (N_17071,N_12781,N_13129);
and U17072 (N_17072,N_13669,N_14828);
nor U17073 (N_17073,N_12687,N_14711);
nor U17074 (N_17074,N_14520,N_13998);
and U17075 (N_17075,N_14543,N_13380);
nor U17076 (N_17076,N_13659,N_12517);
and U17077 (N_17077,N_13023,N_14908);
nor U17078 (N_17078,N_14635,N_14736);
and U17079 (N_17079,N_13403,N_14627);
and U17080 (N_17080,N_13696,N_14938);
nor U17081 (N_17081,N_14323,N_12975);
nand U17082 (N_17082,N_12642,N_13222);
or U17083 (N_17083,N_12590,N_14577);
xor U17084 (N_17084,N_14743,N_13460);
or U17085 (N_17085,N_14500,N_14574);
xnor U17086 (N_17086,N_12842,N_13793);
or U17087 (N_17087,N_13257,N_13627);
and U17088 (N_17088,N_14799,N_13348);
xnor U17089 (N_17089,N_13765,N_12940);
or U17090 (N_17090,N_14674,N_14986);
nand U17091 (N_17091,N_14277,N_14159);
and U17092 (N_17092,N_13338,N_13705);
xnor U17093 (N_17093,N_14821,N_14797);
nor U17094 (N_17094,N_14234,N_13679);
xor U17095 (N_17095,N_14693,N_14091);
and U17096 (N_17096,N_14054,N_13470);
and U17097 (N_17097,N_12683,N_13966);
nand U17098 (N_17098,N_14768,N_13910);
nor U17099 (N_17099,N_14311,N_14825);
nand U17100 (N_17100,N_14633,N_13369);
or U17101 (N_17101,N_13205,N_12846);
nor U17102 (N_17102,N_13131,N_14003);
and U17103 (N_17103,N_14277,N_13590);
and U17104 (N_17104,N_12911,N_12859);
or U17105 (N_17105,N_14141,N_14187);
and U17106 (N_17106,N_14984,N_12856);
nor U17107 (N_17107,N_12541,N_14667);
xnor U17108 (N_17108,N_14753,N_14426);
nor U17109 (N_17109,N_13306,N_12567);
nand U17110 (N_17110,N_13106,N_13475);
or U17111 (N_17111,N_13237,N_13394);
nor U17112 (N_17112,N_14010,N_14470);
xnor U17113 (N_17113,N_14235,N_12788);
or U17114 (N_17114,N_13155,N_12951);
or U17115 (N_17115,N_12857,N_14372);
and U17116 (N_17116,N_12794,N_12559);
and U17117 (N_17117,N_14389,N_13153);
and U17118 (N_17118,N_13990,N_14415);
or U17119 (N_17119,N_13932,N_12749);
nand U17120 (N_17120,N_13029,N_14461);
nand U17121 (N_17121,N_13840,N_14699);
nand U17122 (N_17122,N_13833,N_14639);
nor U17123 (N_17123,N_12636,N_14155);
nor U17124 (N_17124,N_12947,N_13889);
nor U17125 (N_17125,N_14431,N_13323);
nor U17126 (N_17126,N_12871,N_12537);
xnor U17127 (N_17127,N_14249,N_14611);
and U17128 (N_17128,N_12586,N_13951);
nand U17129 (N_17129,N_14271,N_12859);
nor U17130 (N_17130,N_14994,N_14680);
or U17131 (N_17131,N_12915,N_13002);
nor U17132 (N_17132,N_13063,N_13908);
nor U17133 (N_17133,N_12967,N_14019);
and U17134 (N_17134,N_12928,N_14549);
nand U17135 (N_17135,N_14228,N_13663);
nor U17136 (N_17136,N_12740,N_12856);
xnor U17137 (N_17137,N_12655,N_12692);
nand U17138 (N_17138,N_13675,N_12652);
and U17139 (N_17139,N_12963,N_14974);
or U17140 (N_17140,N_13861,N_13351);
nor U17141 (N_17141,N_12933,N_13371);
xnor U17142 (N_17142,N_14903,N_14256);
nand U17143 (N_17143,N_14605,N_14574);
or U17144 (N_17144,N_13205,N_13200);
and U17145 (N_17145,N_14856,N_14861);
xor U17146 (N_17146,N_14585,N_12714);
nor U17147 (N_17147,N_13972,N_14184);
nand U17148 (N_17148,N_14177,N_14266);
nand U17149 (N_17149,N_12626,N_12589);
nand U17150 (N_17150,N_14169,N_12764);
nor U17151 (N_17151,N_12877,N_14419);
and U17152 (N_17152,N_13624,N_14528);
nor U17153 (N_17153,N_14490,N_13732);
and U17154 (N_17154,N_13436,N_13313);
nor U17155 (N_17155,N_14733,N_13037);
or U17156 (N_17156,N_14188,N_13662);
and U17157 (N_17157,N_13252,N_12716);
and U17158 (N_17158,N_13580,N_14614);
or U17159 (N_17159,N_14495,N_13667);
and U17160 (N_17160,N_14841,N_14712);
or U17161 (N_17161,N_13671,N_14566);
or U17162 (N_17162,N_14813,N_13633);
nand U17163 (N_17163,N_14480,N_14166);
nand U17164 (N_17164,N_14052,N_14972);
or U17165 (N_17165,N_13211,N_13068);
or U17166 (N_17166,N_14101,N_12621);
or U17167 (N_17167,N_14166,N_13712);
and U17168 (N_17168,N_13868,N_13913);
or U17169 (N_17169,N_13540,N_13179);
or U17170 (N_17170,N_12623,N_14829);
xor U17171 (N_17171,N_13697,N_13488);
nor U17172 (N_17172,N_12979,N_13289);
and U17173 (N_17173,N_14433,N_13203);
and U17174 (N_17174,N_13577,N_14489);
nor U17175 (N_17175,N_14131,N_13943);
nand U17176 (N_17176,N_14775,N_13321);
or U17177 (N_17177,N_12855,N_13331);
nor U17178 (N_17178,N_12743,N_14153);
or U17179 (N_17179,N_13432,N_13817);
xor U17180 (N_17180,N_13255,N_13300);
or U17181 (N_17181,N_14421,N_12776);
and U17182 (N_17182,N_13944,N_14946);
and U17183 (N_17183,N_12753,N_14243);
nand U17184 (N_17184,N_12991,N_13477);
nand U17185 (N_17185,N_14415,N_12512);
nor U17186 (N_17186,N_13814,N_13362);
xor U17187 (N_17187,N_14515,N_13427);
xor U17188 (N_17188,N_14402,N_13423);
nor U17189 (N_17189,N_14531,N_13734);
nand U17190 (N_17190,N_14336,N_14678);
and U17191 (N_17191,N_12641,N_14144);
or U17192 (N_17192,N_13677,N_14470);
nor U17193 (N_17193,N_13689,N_13280);
nand U17194 (N_17194,N_13151,N_13268);
nor U17195 (N_17195,N_13946,N_14554);
nor U17196 (N_17196,N_13143,N_13069);
and U17197 (N_17197,N_14923,N_14098);
or U17198 (N_17198,N_13038,N_13250);
nor U17199 (N_17199,N_14693,N_12745);
and U17200 (N_17200,N_13413,N_14811);
nand U17201 (N_17201,N_13648,N_14179);
or U17202 (N_17202,N_14876,N_13277);
and U17203 (N_17203,N_14470,N_14337);
nor U17204 (N_17204,N_14745,N_14453);
or U17205 (N_17205,N_13267,N_12605);
nand U17206 (N_17206,N_14473,N_14891);
or U17207 (N_17207,N_14055,N_13765);
nor U17208 (N_17208,N_13037,N_13819);
and U17209 (N_17209,N_13552,N_14441);
xor U17210 (N_17210,N_12595,N_12845);
xor U17211 (N_17211,N_12929,N_14801);
nand U17212 (N_17212,N_12692,N_14183);
nor U17213 (N_17213,N_12770,N_13622);
nand U17214 (N_17214,N_12532,N_12697);
and U17215 (N_17215,N_12883,N_14973);
and U17216 (N_17216,N_14343,N_13879);
nand U17217 (N_17217,N_14090,N_12775);
nor U17218 (N_17218,N_14003,N_14815);
nand U17219 (N_17219,N_14096,N_13185);
xor U17220 (N_17220,N_14455,N_14683);
nand U17221 (N_17221,N_13945,N_14643);
nand U17222 (N_17222,N_13966,N_14822);
and U17223 (N_17223,N_13671,N_12523);
or U17224 (N_17224,N_13644,N_12503);
or U17225 (N_17225,N_12960,N_14048);
nand U17226 (N_17226,N_12773,N_13784);
and U17227 (N_17227,N_12727,N_13494);
nor U17228 (N_17228,N_14825,N_13300);
or U17229 (N_17229,N_13982,N_14444);
or U17230 (N_17230,N_13449,N_14317);
and U17231 (N_17231,N_13707,N_14538);
xor U17232 (N_17232,N_13070,N_12619);
nand U17233 (N_17233,N_13673,N_14245);
nand U17234 (N_17234,N_14141,N_14731);
xor U17235 (N_17235,N_14161,N_14517);
nor U17236 (N_17236,N_14962,N_12921);
nand U17237 (N_17237,N_14944,N_12720);
nand U17238 (N_17238,N_14223,N_12531);
nand U17239 (N_17239,N_14178,N_12919);
and U17240 (N_17240,N_13483,N_13678);
xnor U17241 (N_17241,N_14029,N_13421);
or U17242 (N_17242,N_13057,N_13027);
nand U17243 (N_17243,N_13015,N_13659);
or U17244 (N_17244,N_14061,N_13071);
nand U17245 (N_17245,N_14615,N_12863);
nor U17246 (N_17246,N_13772,N_12840);
and U17247 (N_17247,N_14556,N_12645);
or U17248 (N_17248,N_13713,N_12523);
nor U17249 (N_17249,N_12612,N_13876);
or U17250 (N_17250,N_14184,N_13206);
xor U17251 (N_17251,N_13993,N_13397);
or U17252 (N_17252,N_12679,N_14033);
or U17253 (N_17253,N_14935,N_12934);
or U17254 (N_17254,N_12529,N_14062);
and U17255 (N_17255,N_13891,N_13722);
nor U17256 (N_17256,N_14209,N_13617);
and U17257 (N_17257,N_14671,N_14683);
xnor U17258 (N_17258,N_13717,N_13434);
nor U17259 (N_17259,N_14994,N_14734);
or U17260 (N_17260,N_12725,N_14133);
nor U17261 (N_17261,N_14090,N_13227);
and U17262 (N_17262,N_13943,N_14379);
xnor U17263 (N_17263,N_13894,N_13993);
and U17264 (N_17264,N_13630,N_13981);
nor U17265 (N_17265,N_12720,N_13817);
nor U17266 (N_17266,N_13318,N_14217);
or U17267 (N_17267,N_12972,N_14556);
nor U17268 (N_17268,N_14799,N_14318);
or U17269 (N_17269,N_14376,N_14932);
or U17270 (N_17270,N_14390,N_12926);
and U17271 (N_17271,N_14858,N_14207);
xnor U17272 (N_17272,N_12993,N_14252);
and U17273 (N_17273,N_14494,N_14282);
nor U17274 (N_17274,N_13093,N_12730);
and U17275 (N_17275,N_13470,N_13487);
or U17276 (N_17276,N_13351,N_13910);
or U17277 (N_17277,N_14465,N_14935);
nor U17278 (N_17278,N_13507,N_14103);
and U17279 (N_17279,N_14319,N_14266);
nand U17280 (N_17280,N_14657,N_12621);
nor U17281 (N_17281,N_13748,N_14325);
nand U17282 (N_17282,N_14914,N_13740);
and U17283 (N_17283,N_14509,N_12647);
and U17284 (N_17284,N_13686,N_14904);
and U17285 (N_17285,N_13147,N_14586);
nor U17286 (N_17286,N_12645,N_13702);
or U17287 (N_17287,N_14468,N_13982);
or U17288 (N_17288,N_13713,N_14762);
nand U17289 (N_17289,N_14905,N_13373);
and U17290 (N_17290,N_13964,N_14318);
nand U17291 (N_17291,N_12858,N_14968);
nand U17292 (N_17292,N_14269,N_13005);
and U17293 (N_17293,N_12792,N_13270);
nand U17294 (N_17294,N_14803,N_14811);
or U17295 (N_17295,N_13067,N_14203);
xnor U17296 (N_17296,N_13663,N_13421);
nand U17297 (N_17297,N_13037,N_14181);
and U17298 (N_17298,N_12919,N_12816);
nor U17299 (N_17299,N_14698,N_14340);
or U17300 (N_17300,N_12736,N_14430);
and U17301 (N_17301,N_14342,N_13876);
nand U17302 (N_17302,N_14146,N_13820);
nand U17303 (N_17303,N_13209,N_12712);
or U17304 (N_17304,N_13993,N_14012);
or U17305 (N_17305,N_12789,N_14270);
xor U17306 (N_17306,N_14069,N_14136);
nand U17307 (N_17307,N_12644,N_13866);
and U17308 (N_17308,N_14263,N_14959);
and U17309 (N_17309,N_13098,N_14844);
xnor U17310 (N_17310,N_14192,N_14014);
and U17311 (N_17311,N_13069,N_13275);
nand U17312 (N_17312,N_12872,N_12804);
and U17313 (N_17313,N_14804,N_13981);
and U17314 (N_17314,N_14057,N_12930);
nor U17315 (N_17315,N_13788,N_14814);
and U17316 (N_17316,N_14763,N_14662);
or U17317 (N_17317,N_14047,N_14509);
or U17318 (N_17318,N_13579,N_14395);
or U17319 (N_17319,N_13923,N_14326);
and U17320 (N_17320,N_13140,N_12664);
and U17321 (N_17321,N_13358,N_14206);
or U17322 (N_17322,N_13231,N_14312);
nor U17323 (N_17323,N_13192,N_13371);
xor U17324 (N_17324,N_12631,N_13128);
nor U17325 (N_17325,N_14365,N_12998);
nand U17326 (N_17326,N_14060,N_12685);
and U17327 (N_17327,N_14461,N_12715);
nor U17328 (N_17328,N_14897,N_12641);
nor U17329 (N_17329,N_14253,N_14581);
nor U17330 (N_17330,N_12759,N_13889);
nand U17331 (N_17331,N_12687,N_12864);
or U17332 (N_17332,N_13236,N_13782);
nor U17333 (N_17333,N_13626,N_14726);
nand U17334 (N_17334,N_14739,N_13617);
or U17335 (N_17335,N_13742,N_13566);
or U17336 (N_17336,N_12969,N_13928);
nor U17337 (N_17337,N_12695,N_13286);
or U17338 (N_17338,N_13994,N_14908);
and U17339 (N_17339,N_14230,N_12991);
or U17340 (N_17340,N_14851,N_14550);
or U17341 (N_17341,N_13173,N_13148);
and U17342 (N_17342,N_14365,N_12773);
xnor U17343 (N_17343,N_12772,N_13928);
nand U17344 (N_17344,N_14543,N_13046);
nand U17345 (N_17345,N_13514,N_13869);
or U17346 (N_17346,N_13327,N_13985);
and U17347 (N_17347,N_14593,N_13218);
or U17348 (N_17348,N_12945,N_12551);
or U17349 (N_17349,N_14656,N_14665);
nand U17350 (N_17350,N_13890,N_14930);
nor U17351 (N_17351,N_13250,N_13260);
xnor U17352 (N_17352,N_12530,N_12977);
nor U17353 (N_17353,N_14509,N_13250);
nand U17354 (N_17354,N_12660,N_13365);
or U17355 (N_17355,N_14952,N_12769);
or U17356 (N_17356,N_13731,N_12760);
nor U17357 (N_17357,N_14819,N_13820);
nand U17358 (N_17358,N_13746,N_13028);
or U17359 (N_17359,N_13706,N_12651);
nand U17360 (N_17360,N_13080,N_13941);
nand U17361 (N_17361,N_12752,N_14760);
xnor U17362 (N_17362,N_14551,N_14676);
or U17363 (N_17363,N_14391,N_13500);
nor U17364 (N_17364,N_13261,N_14566);
nand U17365 (N_17365,N_14366,N_13633);
nand U17366 (N_17366,N_14013,N_13438);
or U17367 (N_17367,N_14815,N_14283);
and U17368 (N_17368,N_14339,N_12974);
nand U17369 (N_17369,N_14317,N_13484);
or U17370 (N_17370,N_14701,N_14417);
nand U17371 (N_17371,N_13890,N_14590);
nor U17372 (N_17372,N_14602,N_14334);
and U17373 (N_17373,N_12632,N_14016);
nor U17374 (N_17374,N_13515,N_14280);
xor U17375 (N_17375,N_13714,N_14980);
nand U17376 (N_17376,N_13370,N_13839);
nor U17377 (N_17377,N_12695,N_12683);
nand U17378 (N_17378,N_13783,N_14303);
and U17379 (N_17379,N_14353,N_13461);
or U17380 (N_17380,N_14820,N_12961);
nor U17381 (N_17381,N_13276,N_14767);
or U17382 (N_17382,N_14274,N_13220);
nor U17383 (N_17383,N_14424,N_13514);
xor U17384 (N_17384,N_13281,N_12855);
or U17385 (N_17385,N_14748,N_13307);
nor U17386 (N_17386,N_13091,N_13979);
nand U17387 (N_17387,N_12572,N_14813);
and U17388 (N_17388,N_12841,N_14995);
nor U17389 (N_17389,N_14669,N_13391);
and U17390 (N_17390,N_14366,N_14971);
xor U17391 (N_17391,N_14957,N_14356);
nor U17392 (N_17392,N_12751,N_14670);
nor U17393 (N_17393,N_13196,N_12796);
nand U17394 (N_17394,N_12943,N_13264);
nor U17395 (N_17395,N_13847,N_14924);
or U17396 (N_17396,N_13364,N_13518);
or U17397 (N_17397,N_13272,N_14289);
nand U17398 (N_17398,N_12658,N_14166);
nor U17399 (N_17399,N_13821,N_14874);
nor U17400 (N_17400,N_12940,N_12835);
nor U17401 (N_17401,N_12507,N_13465);
nand U17402 (N_17402,N_14721,N_14528);
nor U17403 (N_17403,N_14251,N_12716);
xor U17404 (N_17404,N_12882,N_13435);
nand U17405 (N_17405,N_14910,N_14671);
or U17406 (N_17406,N_14451,N_12779);
nand U17407 (N_17407,N_13073,N_12755);
or U17408 (N_17408,N_14413,N_12962);
or U17409 (N_17409,N_14526,N_13584);
nor U17410 (N_17410,N_13656,N_14544);
nand U17411 (N_17411,N_14996,N_13557);
or U17412 (N_17412,N_13722,N_13668);
xnor U17413 (N_17413,N_13721,N_13992);
and U17414 (N_17414,N_14661,N_14399);
and U17415 (N_17415,N_13048,N_14794);
nor U17416 (N_17416,N_13644,N_13204);
or U17417 (N_17417,N_13033,N_13342);
and U17418 (N_17418,N_14025,N_14098);
or U17419 (N_17419,N_12653,N_14267);
xnor U17420 (N_17420,N_14381,N_14216);
or U17421 (N_17421,N_12810,N_13762);
nor U17422 (N_17422,N_14414,N_13602);
xnor U17423 (N_17423,N_14054,N_12675);
nand U17424 (N_17424,N_14482,N_14886);
or U17425 (N_17425,N_13746,N_12997);
or U17426 (N_17426,N_14402,N_14164);
and U17427 (N_17427,N_13493,N_12975);
nand U17428 (N_17428,N_13445,N_12978);
and U17429 (N_17429,N_12673,N_12786);
nor U17430 (N_17430,N_13996,N_13752);
and U17431 (N_17431,N_14941,N_14320);
and U17432 (N_17432,N_14190,N_12512);
or U17433 (N_17433,N_13482,N_13123);
and U17434 (N_17434,N_12953,N_14893);
and U17435 (N_17435,N_14294,N_12719);
or U17436 (N_17436,N_13866,N_13198);
and U17437 (N_17437,N_14249,N_12509);
nor U17438 (N_17438,N_14923,N_13282);
nor U17439 (N_17439,N_13289,N_13366);
xor U17440 (N_17440,N_13605,N_14512);
or U17441 (N_17441,N_12753,N_14380);
nand U17442 (N_17442,N_12828,N_14034);
or U17443 (N_17443,N_14805,N_14136);
and U17444 (N_17444,N_13866,N_14388);
and U17445 (N_17445,N_13462,N_13534);
and U17446 (N_17446,N_14409,N_13241);
nor U17447 (N_17447,N_12690,N_12798);
and U17448 (N_17448,N_14010,N_14146);
or U17449 (N_17449,N_14338,N_14199);
and U17450 (N_17450,N_14314,N_14379);
or U17451 (N_17451,N_13596,N_13526);
and U17452 (N_17452,N_13618,N_13160);
nand U17453 (N_17453,N_14635,N_14107);
and U17454 (N_17454,N_14964,N_13974);
and U17455 (N_17455,N_13137,N_12725);
nand U17456 (N_17456,N_13467,N_14510);
and U17457 (N_17457,N_14969,N_13931);
and U17458 (N_17458,N_12648,N_13459);
or U17459 (N_17459,N_14954,N_14593);
nor U17460 (N_17460,N_13553,N_12641);
nand U17461 (N_17461,N_14297,N_14728);
or U17462 (N_17462,N_13779,N_14866);
nor U17463 (N_17463,N_13259,N_12813);
and U17464 (N_17464,N_13704,N_14097);
nor U17465 (N_17465,N_14308,N_14379);
nor U17466 (N_17466,N_14564,N_14311);
or U17467 (N_17467,N_13592,N_13151);
nand U17468 (N_17468,N_13860,N_12725);
nand U17469 (N_17469,N_13069,N_12551);
and U17470 (N_17470,N_13579,N_14641);
nor U17471 (N_17471,N_13334,N_13080);
nand U17472 (N_17472,N_12534,N_14802);
nand U17473 (N_17473,N_13742,N_14287);
xor U17474 (N_17474,N_13837,N_14830);
nor U17475 (N_17475,N_14028,N_14079);
nand U17476 (N_17476,N_13519,N_13322);
xnor U17477 (N_17477,N_14669,N_13426);
nand U17478 (N_17478,N_12569,N_14691);
nor U17479 (N_17479,N_14526,N_14832);
nor U17480 (N_17480,N_14665,N_14193);
xnor U17481 (N_17481,N_14551,N_14084);
and U17482 (N_17482,N_14623,N_14289);
or U17483 (N_17483,N_14794,N_13949);
or U17484 (N_17484,N_14556,N_12568);
and U17485 (N_17485,N_13877,N_13032);
nand U17486 (N_17486,N_12791,N_12811);
and U17487 (N_17487,N_13150,N_13946);
nand U17488 (N_17488,N_13686,N_14004);
or U17489 (N_17489,N_12651,N_13691);
nand U17490 (N_17490,N_13033,N_12850);
nor U17491 (N_17491,N_13686,N_14551);
or U17492 (N_17492,N_13018,N_14196);
nor U17493 (N_17493,N_13252,N_13544);
nor U17494 (N_17494,N_13661,N_13404);
and U17495 (N_17495,N_12945,N_14730);
or U17496 (N_17496,N_14506,N_13858);
and U17497 (N_17497,N_13106,N_13673);
xnor U17498 (N_17498,N_13643,N_14974);
nand U17499 (N_17499,N_13844,N_14882);
and U17500 (N_17500,N_15954,N_15265);
nand U17501 (N_17501,N_15592,N_16124);
nor U17502 (N_17502,N_16850,N_15906);
nand U17503 (N_17503,N_16834,N_16161);
and U17504 (N_17504,N_15752,N_17073);
xor U17505 (N_17505,N_16110,N_15358);
nand U17506 (N_17506,N_16919,N_15572);
xor U17507 (N_17507,N_15822,N_15606);
xnor U17508 (N_17508,N_15922,N_17253);
nand U17509 (N_17509,N_16815,N_15749);
nand U17510 (N_17510,N_16804,N_17230);
nor U17511 (N_17511,N_16095,N_15924);
nand U17512 (N_17512,N_15016,N_16399);
nor U17513 (N_17513,N_15722,N_16824);
xor U17514 (N_17514,N_16250,N_15033);
and U17515 (N_17515,N_17374,N_15447);
or U17516 (N_17516,N_17248,N_17267);
nand U17517 (N_17517,N_17141,N_15996);
nor U17518 (N_17518,N_16353,N_16022);
nor U17519 (N_17519,N_15081,N_16163);
and U17520 (N_17520,N_16916,N_15925);
nor U17521 (N_17521,N_15493,N_17499);
nor U17522 (N_17522,N_16092,N_15389);
nor U17523 (N_17523,N_16688,N_15923);
or U17524 (N_17524,N_15931,N_15860);
and U17525 (N_17525,N_15131,N_15176);
nor U17526 (N_17526,N_15266,N_17407);
xnor U17527 (N_17527,N_15742,N_15034);
xor U17528 (N_17528,N_16818,N_16618);
and U17529 (N_17529,N_16287,N_16104);
and U17530 (N_17530,N_15712,N_15657);
or U17531 (N_17531,N_16579,N_16443);
nor U17532 (N_17532,N_15124,N_15834);
nand U17533 (N_17533,N_16917,N_15256);
and U17534 (N_17534,N_17363,N_16844);
nand U17535 (N_17535,N_15472,N_15270);
or U17536 (N_17536,N_15109,N_15616);
nor U17537 (N_17537,N_16224,N_17204);
xor U17538 (N_17538,N_15709,N_17370);
or U17539 (N_17539,N_15073,N_16629);
nor U17540 (N_17540,N_17268,N_16187);
and U17541 (N_17541,N_17325,N_15519);
or U17542 (N_17542,N_15064,N_15324);
nand U17543 (N_17543,N_17453,N_15411);
nor U17544 (N_17544,N_15175,N_15236);
xnor U17545 (N_17545,N_16821,N_17340);
nor U17546 (N_17546,N_16680,N_15121);
xnor U17547 (N_17547,N_17480,N_16617);
or U17548 (N_17548,N_17240,N_15813);
or U17549 (N_17549,N_17378,N_15443);
nor U17550 (N_17550,N_15908,N_16752);
nand U17551 (N_17551,N_15126,N_15174);
xor U17552 (N_17552,N_15505,N_15186);
nand U17553 (N_17553,N_15886,N_17175);
or U17554 (N_17554,N_16165,N_15146);
and U17555 (N_17555,N_16097,N_16217);
and U17556 (N_17556,N_16973,N_15934);
or U17557 (N_17557,N_15071,N_15531);
nor U17558 (N_17558,N_16085,N_17332);
nor U17559 (N_17559,N_16923,N_17170);
nor U17560 (N_17560,N_17390,N_15720);
nand U17561 (N_17561,N_17421,N_16441);
nand U17562 (N_17562,N_17244,N_15963);
and U17563 (N_17563,N_16429,N_17242);
or U17564 (N_17564,N_16662,N_15969);
and U17565 (N_17565,N_17404,N_15998);
nand U17566 (N_17566,N_15697,N_16836);
nor U17567 (N_17567,N_15274,N_15758);
xnor U17568 (N_17568,N_15764,N_15565);
and U17569 (N_17569,N_15306,N_16442);
xor U17570 (N_17570,N_15976,N_15352);
or U17571 (N_17571,N_16706,N_16091);
nor U17572 (N_17572,N_15234,N_16042);
xor U17573 (N_17573,N_15221,N_15046);
or U17574 (N_17574,N_15083,N_17098);
or U17575 (N_17575,N_16690,N_16137);
and U17576 (N_17576,N_16745,N_15248);
nand U17577 (N_17577,N_16342,N_16955);
and U17578 (N_17578,N_16766,N_16920);
xor U17579 (N_17579,N_17142,N_15661);
and U17580 (N_17580,N_15768,N_16265);
or U17581 (N_17581,N_17041,N_15326);
nand U17582 (N_17582,N_15927,N_15485);
nand U17583 (N_17583,N_15757,N_15580);
nor U17584 (N_17584,N_15172,N_16130);
or U17585 (N_17585,N_16587,N_15189);
nor U17586 (N_17586,N_16350,N_17245);
nand U17587 (N_17587,N_15036,N_16545);
or U17588 (N_17588,N_15353,N_16149);
or U17589 (N_17589,N_15714,N_16822);
or U17590 (N_17590,N_17256,N_17473);
or U17591 (N_17591,N_16950,N_17354);
and U17592 (N_17592,N_15308,N_16538);
nand U17593 (N_17593,N_17434,N_16286);
nand U17594 (N_17594,N_16747,N_15384);
nor U17595 (N_17595,N_17420,N_16310);
and U17596 (N_17596,N_16986,N_16479);
nor U17597 (N_17597,N_16174,N_17428);
and U17598 (N_17598,N_17439,N_16112);
nand U17599 (N_17599,N_17058,N_15032);
nand U17600 (N_17600,N_15800,N_15534);
xor U17601 (N_17601,N_17092,N_15433);
or U17602 (N_17602,N_15831,N_16886);
nor U17603 (N_17603,N_15010,N_16450);
and U17604 (N_17604,N_16235,N_17344);
nor U17605 (N_17605,N_15003,N_15008);
or U17606 (N_17606,N_16282,N_17192);
nor U17607 (N_17607,N_15686,N_15390);
nand U17608 (N_17608,N_17020,N_15878);
and U17609 (N_17609,N_15761,N_16832);
xor U17610 (N_17610,N_15669,N_17030);
and U17611 (N_17611,N_16887,N_15862);
or U17612 (N_17612,N_15090,N_15544);
nor U17613 (N_17613,N_16432,N_15475);
xor U17614 (N_17614,N_15244,N_16323);
or U17615 (N_17615,N_15226,N_15844);
nor U17616 (N_17616,N_16400,N_16966);
and U17617 (N_17617,N_15889,N_15483);
nor U17618 (N_17618,N_17101,N_17074);
nor U17619 (N_17619,N_15677,N_16312);
nor U17620 (N_17620,N_17094,N_15211);
nor U17621 (N_17621,N_17087,N_15796);
nor U17622 (N_17622,N_15624,N_16653);
or U17623 (N_17623,N_16623,N_16727);
nor U17624 (N_17624,N_17379,N_15710);
or U17625 (N_17625,N_17444,N_17157);
nand U17626 (N_17626,N_15741,N_17280);
or U17627 (N_17627,N_16155,N_15028);
or U17628 (N_17628,N_15106,N_15594);
or U17629 (N_17629,N_16489,N_16245);
or U17630 (N_17630,N_16697,N_15776);
or U17631 (N_17631,N_17128,N_15070);
xnor U17632 (N_17632,N_16713,N_16214);
and U17633 (N_17633,N_16499,N_16358);
nor U17634 (N_17634,N_16019,N_15639);
nor U17635 (N_17635,N_17111,N_16608);
or U17636 (N_17636,N_17306,N_16748);
xor U17637 (N_17637,N_15943,N_15099);
nor U17638 (N_17638,N_16719,N_17347);
and U17639 (N_17639,N_16811,N_16632);
nor U17640 (N_17640,N_16351,N_15941);
and U17641 (N_17641,N_16267,N_16225);
and U17642 (N_17642,N_15119,N_16613);
or U17643 (N_17643,N_16740,N_16573);
nor U17644 (N_17644,N_16865,N_15209);
nor U17645 (N_17645,N_15903,N_17290);
nand U17646 (N_17646,N_15799,N_16056);
and U17647 (N_17647,N_16581,N_15554);
nor U17648 (N_17648,N_17257,N_16589);
nand U17649 (N_17649,N_15664,N_15314);
nand U17650 (N_17650,N_16256,N_15332);
and U17651 (N_17651,N_16989,N_16561);
or U17652 (N_17652,N_16813,N_17497);
and U17653 (N_17653,N_16689,N_16055);
nor U17654 (N_17654,N_16776,N_16122);
or U17655 (N_17655,N_16728,N_17062);
and U17656 (N_17656,N_17425,N_15744);
or U17657 (N_17657,N_15229,N_16131);
nor U17658 (N_17658,N_17485,N_16507);
or U17659 (N_17659,N_17021,N_17316);
nor U17660 (N_17660,N_15535,N_17266);
and U17661 (N_17661,N_16830,N_16909);
nand U17662 (N_17662,N_17422,N_17326);
nor U17663 (N_17663,N_15995,N_15958);
and U17664 (N_17664,N_15093,N_16810);
and U17665 (N_17665,N_15165,N_15425);
and U17666 (N_17666,N_16251,N_16356);
or U17667 (N_17667,N_15543,N_15279);
or U17668 (N_17668,N_15777,N_17038);
nor U17669 (N_17669,N_16907,N_17229);
or U17670 (N_17670,N_17068,N_16366);
xnor U17671 (N_17671,N_16864,N_15842);
or U17672 (N_17672,N_16714,N_15436);
xnor U17673 (N_17673,N_15492,N_16999);
and U17674 (N_17674,N_16199,N_16164);
nor U17675 (N_17675,N_15467,N_15438);
nor U17676 (N_17676,N_17351,N_15147);
nand U17677 (N_17677,N_16681,N_17317);
nor U17678 (N_17678,N_16597,N_15988);
xor U17679 (N_17679,N_16381,N_15437);
and U17680 (N_17680,N_15557,N_15414);
nand U17681 (N_17681,N_15487,N_16767);
or U17682 (N_17682,N_15548,N_16814);
nand U17683 (N_17683,N_17149,N_16152);
nor U17684 (N_17684,N_16519,N_17125);
nor U17685 (N_17685,N_15006,N_17088);
nor U17686 (N_17686,N_16548,N_15335);
or U17687 (N_17687,N_15238,N_16274);
nor U17688 (N_17688,N_15541,N_16258);
and U17689 (N_17689,N_15788,N_16123);
and U17690 (N_17690,N_16705,N_15104);
and U17691 (N_17691,N_17348,N_17258);
xor U17692 (N_17692,N_17213,N_16153);
or U17693 (N_17693,N_16614,N_17368);
nor U17694 (N_17694,N_17346,N_15169);
xnor U17695 (N_17695,N_15695,N_15625);
xor U17696 (N_17696,N_16178,N_15247);
and U17697 (N_17697,N_17295,N_16357);
nor U17698 (N_17698,N_15972,N_15719);
nand U17699 (N_17699,N_16079,N_15207);
nand U17700 (N_17700,N_17353,N_16223);
xor U17701 (N_17701,N_16228,N_16635);
nor U17702 (N_17702,N_17312,N_16827);
nor U17703 (N_17703,N_17081,N_15944);
nand U17704 (N_17704,N_17022,N_15869);
and U17705 (N_17705,N_16665,N_15739);
and U17706 (N_17706,N_17144,N_15539);
and U17707 (N_17707,N_16168,N_16290);
nor U17708 (N_17708,N_16983,N_15164);
or U17709 (N_17709,N_16263,N_15357);
and U17710 (N_17710,N_17123,N_16445);
nand U17711 (N_17711,N_17493,N_16807);
and U17712 (N_17712,N_15687,N_16504);
nor U17713 (N_17713,N_16615,N_16255);
nor U17714 (N_17714,N_15840,N_15706);
xor U17715 (N_17715,N_15344,N_16718);
nand U17716 (N_17716,N_17061,N_15901);
nand U17717 (N_17717,N_16028,N_17406);
and U17718 (N_17718,N_16652,N_15632);
nor U17719 (N_17719,N_15152,N_15916);
nand U17720 (N_17720,N_16569,N_15865);
nor U17721 (N_17721,N_15649,N_15276);
nor U17722 (N_17722,N_16295,N_17400);
and U17723 (N_17723,N_16749,N_16057);
nor U17724 (N_17724,N_15202,N_15666);
and U17725 (N_17725,N_15213,N_16183);
or U17726 (N_17726,N_15981,N_15452);
or U17727 (N_17727,N_15679,N_17132);
or U17728 (N_17728,N_15382,N_16655);
nor U17729 (N_17729,N_16160,N_16064);
nor U17730 (N_17730,N_16393,N_16763);
and U17731 (N_17731,N_15037,N_15601);
nor U17732 (N_17732,N_16645,N_17148);
and U17733 (N_17733,N_16189,N_15775);
or U17734 (N_17734,N_17090,N_17078);
and U17735 (N_17735,N_15045,N_17051);
nor U17736 (N_17736,N_15614,N_16646);
or U17737 (N_17737,N_15275,N_15428);
nand U17738 (N_17738,N_17286,N_15284);
and U17739 (N_17739,N_15643,N_15082);
or U17740 (N_17740,N_15962,N_16654);
or U17741 (N_17741,N_15792,N_16177);
xor U17742 (N_17742,N_16476,N_15748);
nand U17743 (N_17743,N_16757,N_16630);
or U17744 (N_17744,N_17122,N_16457);
and U17745 (N_17745,N_16799,N_15011);
or U17746 (N_17746,N_15479,N_17430);
and U17747 (N_17747,N_16081,N_15658);
nor U17748 (N_17748,N_15772,N_17104);
and U17749 (N_17749,N_16625,N_15449);
nand U17750 (N_17750,N_16735,N_15937);
nand U17751 (N_17751,N_17152,N_16492);
nand U17752 (N_17752,N_16930,N_16143);
or U17753 (N_17753,N_16634,N_15759);
or U17754 (N_17754,N_16201,N_17262);
nand U17755 (N_17755,N_15451,N_17118);
xnor U17756 (N_17756,N_16150,N_17447);
nor U17757 (N_17757,N_16211,N_16502);
nand U17758 (N_17758,N_15404,N_15065);
nand U17759 (N_17759,N_15835,N_15043);
or U17760 (N_17760,N_16586,N_15930);
nor U17761 (N_17761,N_16965,N_15893);
nor U17762 (N_17762,N_17367,N_16699);
nor U17763 (N_17763,N_15359,N_15114);
xnor U17764 (N_17764,N_17324,N_15385);
nand U17765 (N_17765,N_15012,N_15026);
nand U17766 (N_17766,N_16873,N_15725);
xor U17767 (N_17767,N_17441,N_15586);
and U17768 (N_17768,N_16825,N_17272);
nand U17769 (N_17769,N_15182,N_15219);
and U17770 (N_17770,N_15975,N_17389);
nand U17771 (N_17771,N_17446,N_17357);
nor U17772 (N_17772,N_16991,N_15965);
and U17773 (N_17773,N_16687,N_17130);
or U17774 (N_17774,N_15120,N_15904);
or U17775 (N_17775,N_17080,N_17483);
nand U17776 (N_17776,N_15007,N_16760);
and U17777 (N_17777,N_17408,N_16754);
or U17778 (N_17778,N_17403,N_17381);
and U17779 (N_17779,N_16773,N_16658);
nor U17780 (N_17780,N_15674,N_17172);
and U17781 (N_17781,N_16927,N_17489);
nor U17782 (N_17782,N_15401,N_15086);
nand U17783 (N_17783,N_15646,N_17469);
and U17784 (N_17784,N_16514,N_15349);
nand U17785 (N_17785,N_15481,N_15518);
nand U17786 (N_17786,N_15023,N_15555);
and U17787 (N_17787,N_15292,N_15949);
xnor U17788 (N_17788,N_16099,N_16898);
nand U17789 (N_17789,N_16076,N_16456);
or U17790 (N_17790,N_16451,N_16431);
xor U17791 (N_17791,N_16259,N_16304);
nor U17792 (N_17792,N_16289,N_16877);
nand U17793 (N_17793,N_17435,N_16379);
xnor U17794 (N_17794,N_17259,N_17195);
xor U17795 (N_17795,N_16606,N_16015);
and U17796 (N_17796,N_17458,N_15162);
nor U17797 (N_17797,N_16102,N_17288);
xnor U17798 (N_17798,N_17083,N_16885);
or U17799 (N_17799,N_17216,N_15418);
and U17800 (N_17800,N_17294,N_15599);
or U17801 (N_17801,N_16668,N_15737);
and U17802 (N_17802,N_15637,N_15589);
nor U17803 (N_17803,N_17273,N_16261);
or U17804 (N_17804,N_15057,N_16624);
and U17805 (N_17805,N_17193,N_15148);
nor U17806 (N_17806,N_16861,N_15750);
and U17807 (N_17807,N_15797,N_17487);
nand U17808 (N_17808,N_16820,N_16378);
nor U17809 (N_17809,N_15673,N_15041);
or U17810 (N_17810,N_16862,N_17412);
nor U17811 (N_17811,N_16544,N_16876);
nand U17812 (N_17812,N_15877,N_17089);
nand U17813 (N_17813,N_17084,N_16236);
nand U17814 (N_17814,N_15214,N_15836);
nand U17815 (N_17815,N_16878,N_16895);
xnor U17816 (N_17816,N_16364,N_15612);
or U17817 (N_17817,N_16856,N_16059);
and U17818 (N_17818,N_16349,N_16789);
xnor U17819 (N_17819,N_15511,N_15832);
nor U17820 (N_17820,N_17099,N_16656);
and U17821 (N_17821,N_15939,N_16924);
and U17822 (N_17822,N_15516,N_16897);
or U17823 (N_17823,N_15498,N_15399);
and U17824 (N_17824,N_17300,N_15851);
and U17825 (N_17825,N_16722,N_15833);
or U17826 (N_17826,N_16068,N_15619);
or U17827 (N_17827,N_16583,N_17462);
nand U17828 (N_17828,N_15216,N_17207);
or U17829 (N_17829,N_15859,N_15268);
or U17830 (N_17830,N_15304,N_15682);
nand U17831 (N_17831,N_15473,N_15115);
and U17832 (N_17832,N_15574,N_16248);
or U17833 (N_17833,N_15621,N_17082);
or U17834 (N_17834,N_15956,N_15648);
nand U17835 (N_17835,N_15133,N_16788);
nor U17836 (N_17836,N_17371,N_15559);
xnor U17837 (N_17837,N_16473,N_16002);
or U17838 (N_17838,N_15762,N_16841);
nor U17839 (N_17839,N_15684,N_16087);
and U17840 (N_17840,N_17362,N_16319);
and U17841 (N_17841,N_15774,N_15160);
nor U17842 (N_17842,N_16272,N_15322);
nand U17843 (N_17843,N_16089,N_15784);
xor U17844 (N_17844,N_17241,N_15515);
nand U17845 (N_17845,N_16833,N_16297);
nand U17846 (N_17846,N_17318,N_16014);
or U17847 (N_17847,N_15149,N_15047);
nor U17848 (N_17848,N_16882,N_16227);
nand U17849 (N_17849,N_16711,N_15703);
nand U17850 (N_17850,N_17179,N_15997);
nor U17851 (N_17851,N_17205,N_17310);
or U17852 (N_17852,N_17026,N_15551);
nor U17853 (N_17853,N_16780,N_15435);
and U17854 (N_17854,N_16447,N_15497);
xnor U17855 (N_17855,N_15474,N_15789);
or U17856 (N_17856,N_15463,N_15000);
nand U17857 (N_17857,N_17052,N_16365);
or U17858 (N_17858,N_17431,N_15458);
or U17859 (N_17859,N_15281,N_16459);
nor U17860 (N_17860,N_16128,N_15159);
nor U17861 (N_17861,N_15113,N_17334);
and U17862 (N_17862,N_15538,N_15760);
or U17863 (N_17863,N_16761,N_17464);
nor U17864 (N_17864,N_15478,N_15610);
nand U17865 (N_17865,N_15527,N_15136);
nand U17866 (N_17866,N_16186,N_16559);
nand U17867 (N_17867,N_17498,N_15685);
and U17868 (N_17868,N_15077,N_16208);
or U17869 (N_17869,N_16347,N_15161);
and U17870 (N_17870,N_15504,N_16408);
nand U17871 (N_17871,N_16746,N_16743);
nor U17872 (N_17872,N_17079,N_15873);
or U17873 (N_17873,N_16196,N_15091);
nand U17874 (N_17874,N_16696,N_16077);
nand U17875 (N_17875,N_15400,N_16430);
and U17876 (N_17876,N_16008,N_15864);
nor U17877 (N_17877,N_15263,N_15919);
xor U17878 (N_17878,N_15329,N_17410);
nand U17879 (N_17879,N_15914,N_15343);
or U17880 (N_17880,N_16937,N_16050);
xnor U17881 (N_17881,N_16020,N_15508);
nor U17882 (N_17882,N_15017,N_17131);
or U17883 (N_17883,N_17249,N_16550);
or U17884 (N_17884,N_16866,N_17448);
nor U17885 (N_17885,N_15655,N_16532);
or U17886 (N_17886,N_15421,N_17405);
nand U17887 (N_17887,N_16968,N_15031);
nor U17888 (N_17888,N_16772,N_15578);
nor U17889 (N_17889,N_17113,N_15462);
nand U17890 (N_17890,N_15167,N_16369);
nor U17891 (N_17891,N_16465,N_16226);
xor U17892 (N_17892,N_16009,N_17047);
nor U17893 (N_17893,N_16648,N_16798);
or U17894 (N_17894,N_15320,N_15379);
nand U17895 (N_17895,N_16851,N_15587);
xor U17896 (N_17896,N_16881,N_16275);
nand U17897 (N_17897,N_16232,N_15305);
and U17898 (N_17898,N_17472,N_17222);
and U17899 (N_17899,N_17042,N_15484);
xor U17900 (N_17900,N_16891,N_15361);
nand U17901 (N_17901,N_15122,N_15694);
nand U17902 (N_17902,N_16205,N_16461);
or U17903 (N_17903,N_17440,N_17212);
or U17904 (N_17904,N_16860,N_15080);
nor U17905 (N_17905,N_15579,N_16726);
or U17906 (N_17906,N_16023,N_17279);
and U17907 (N_17907,N_16032,N_16411);
xnor U17908 (N_17908,N_15932,N_15947);
nor U17909 (N_17909,N_17217,N_16552);
nor U17910 (N_17910,N_16691,N_16116);
and U17911 (N_17911,N_16567,N_15547);
xnor U17912 (N_17912,N_15406,N_16280);
and U17913 (N_17913,N_15815,N_16446);
nor U17914 (N_17914,N_15885,N_16333);
and U17915 (N_17915,N_15821,N_15144);
xnor U17916 (N_17916,N_15464,N_15488);
and U17917 (N_17917,N_16120,N_16880);
or U17918 (N_17918,N_15190,N_15921);
and U17919 (N_17919,N_16336,N_16464);
xor U17920 (N_17920,N_15407,N_16636);
nand U17921 (N_17921,N_15460,N_17036);
or U17922 (N_17922,N_15089,N_16739);
nor U17923 (N_17923,N_16555,N_15699);
nand U17924 (N_17924,N_16390,N_15801);
nand U17925 (N_17925,N_17358,N_15662);
nor U17926 (N_17926,N_16854,N_16542);
xnor U17927 (N_17927,N_16281,N_16765);
nand U17928 (N_17928,N_16219,N_15900);
xnor U17929 (N_17929,N_15038,N_17235);
nor U17930 (N_17930,N_17385,N_16375);
nor U17931 (N_17931,N_15667,N_15872);
nor U17932 (N_17932,N_17127,N_16562);
and U17933 (N_17933,N_17046,N_16327);
nand U17934 (N_17934,N_16935,N_17490);
nor U17935 (N_17935,N_15611,N_17278);
and U17936 (N_17936,N_15617,N_15312);
or U17937 (N_17937,N_15005,N_15936);
and U17938 (N_17938,N_16284,N_16101);
nand U17939 (N_17939,N_16669,N_16500);
nor U17940 (N_17940,N_16574,N_16846);
xnor U17941 (N_17941,N_16819,N_16868);
nor U17942 (N_17942,N_16906,N_15968);
and U17943 (N_17943,N_15419,N_16591);
or U17944 (N_17944,N_17488,N_15231);
or U17945 (N_17945,N_17182,N_16065);
or U17946 (N_17946,N_15494,N_15440);
nand U17947 (N_17947,N_16159,N_16285);
and U17948 (N_17948,N_15356,N_16148);
nand U17949 (N_17949,N_16838,N_17387);
and U17950 (N_17950,N_15066,N_17017);
nand U17951 (N_17951,N_16724,N_17337);
or U17952 (N_17952,N_16033,N_16576);
nor U17953 (N_17953,N_16243,N_17292);
nand U17954 (N_17954,N_16721,N_16977);
nor U17955 (N_17955,N_15255,N_15340);
or U17956 (N_17956,N_17121,N_16921);
nand U17957 (N_17957,N_17203,N_16344);
and U17958 (N_17958,N_16318,N_15929);
or U17959 (N_17959,N_15225,N_16115);
nor U17960 (N_17960,N_15261,N_15708);
nand U17961 (N_17961,N_15430,N_17056);
nor U17962 (N_17962,N_17194,N_16816);
or U17963 (N_17963,N_15980,N_15424);
xnor U17964 (N_17964,N_15645,N_17191);
nand U17965 (N_17965,N_15882,N_17289);
nor U17966 (N_17966,N_15564,N_17287);
or U17967 (N_17967,N_15917,N_16449);
and U17968 (N_17968,N_15715,N_16307);
or U17969 (N_17969,N_17178,N_16132);
nor U17970 (N_17970,N_15716,N_16460);
nand U17971 (N_17971,N_15442,N_15432);
nand U17972 (N_17972,N_17236,N_15781);
or U17973 (N_17973,N_16467,N_17187);
nor U17974 (N_17974,N_15393,N_15291);
nor U17975 (N_17975,N_17375,N_16720);
nor U17976 (N_17976,N_17452,N_16515);
nor U17977 (N_17977,N_17014,N_16162);
and U17978 (N_17978,N_16391,N_15856);
or U17979 (N_17979,N_15738,N_16595);
and U17980 (N_17980,N_16170,N_17158);
nor U17981 (N_17981,N_16710,N_15179);
nand U17982 (N_17982,N_17465,N_16271);
and U17983 (N_17983,N_17064,N_16185);
or U17984 (N_17984,N_15055,N_15663);
nand U17985 (N_17985,N_16038,N_15412);
nand U17986 (N_17986,N_15607,N_16401);
nor U17987 (N_17987,N_16412,N_17009);
nand U17988 (N_17988,N_15964,N_17117);
nand U17989 (N_17989,N_17388,N_15985);
nand U17990 (N_17990,N_16436,N_15138);
and U17991 (N_17991,N_15867,N_16478);
nand U17992 (N_17992,N_17200,N_15318);
nor U17993 (N_17993,N_16388,N_16322);
and U17994 (N_17994,N_17395,N_17126);
and U17995 (N_17995,N_16756,N_15260);
nand U17996 (N_17996,N_15523,N_15271);
nand U17997 (N_17997,N_16938,N_17133);
nand U17998 (N_17998,N_15805,N_15307);
xnor U17999 (N_17999,N_15584,N_15140);
or U18000 (N_18000,N_17044,N_16158);
xor U18001 (N_18001,N_16845,N_15913);
nand U18002 (N_18002,N_15942,N_15992);
and U18003 (N_18003,N_16971,N_15946);
nor U18004 (N_18004,N_16229,N_16931);
nand U18005 (N_18005,N_16291,N_15496);
xnor U18006 (N_18006,N_16928,N_17043);
nand U18007 (N_18007,N_17333,N_15783);
and U18008 (N_18008,N_17360,N_15853);
or U18009 (N_18009,N_16034,N_15027);
nand U18010 (N_18010,N_17231,N_17039);
or U18011 (N_18011,N_15187,N_16926);
and U18012 (N_18012,N_15469,N_15367);
or U18013 (N_18013,N_16070,N_16716);
or U18014 (N_18014,N_16188,N_16294);
and U18015 (N_18015,N_16088,N_15210);
nor U18016 (N_18016,N_16406,N_17251);
nand U18017 (N_18017,N_17314,N_15803);
or U18018 (N_18018,N_15651,N_17147);
nor U18019 (N_18019,N_17209,N_15597);
and U18020 (N_18020,N_15938,N_15665);
and U18021 (N_18021,N_15787,N_16676);
and U18022 (N_18022,N_15891,N_15994);
or U18023 (N_18023,N_16485,N_15773);
nand U18024 (N_18024,N_16992,N_15672);
nand U18025 (N_18025,N_15536,N_17169);
and U18026 (N_18026,N_17309,N_17419);
or U18027 (N_18027,N_16321,N_15778);
nor U18028 (N_18028,N_15546,N_17263);
xor U18029 (N_18029,N_15887,N_15371);
and U18030 (N_18030,N_15155,N_16036);
and U18031 (N_18031,N_15294,N_16213);
nand U18032 (N_18032,N_15874,N_16241);
and U18033 (N_18033,N_15638,N_15319);
xor U18034 (N_18034,N_15823,N_15444);
xor U18035 (N_18035,N_15360,N_15987);
nor U18036 (N_18036,N_15520,N_15517);
and U18037 (N_18037,N_16062,N_16744);
nand U18038 (N_18038,N_17075,N_17261);
nand U18039 (N_18039,N_17091,N_17454);
nand U18040 (N_18040,N_15552,N_15567);
xor U18041 (N_18041,N_17029,N_15058);
or U18042 (N_18042,N_16299,N_15239);
and U18043 (N_18043,N_16067,N_17460);
nand U18044 (N_18044,N_16769,N_16797);
nor U18045 (N_18045,N_15628,N_16823);
xor U18046 (N_18046,N_15282,N_17426);
nor U18047 (N_18047,N_15533,N_15670);
nor U18048 (N_18048,N_16433,N_16043);
or U18049 (N_18049,N_15573,N_16270);
xor U18050 (N_18050,N_17033,N_15094);
nor U18051 (N_18051,N_17071,N_16783);
nor U18052 (N_18052,N_15604,N_15782);
and U18053 (N_18053,N_15688,N_16970);
nor U18054 (N_18054,N_15561,N_16260);
nand U18055 (N_18055,N_16407,N_16296);
or U18056 (N_18056,N_15053,N_15883);
and U18057 (N_18057,N_17032,N_16702);
xnor U18058 (N_18058,N_17180,N_16462);
or U18059 (N_18059,N_17341,N_16018);
and U18060 (N_18060,N_15251,N_17461);
or U18061 (N_18061,N_17119,N_17006);
or U18062 (N_18062,N_17449,N_16354);
and U18063 (N_18063,N_15156,N_15056);
xor U18064 (N_18064,N_16602,N_17311);
or U18065 (N_18065,N_16604,N_15890);
xor U18066 (N_18066,N_15092,N_15383);
xnor U18067 (N_18067,N_16497,N_15957);
or U18068 (N_18068,N_16305,N_15491);
or U18069 (N_18069,N_16300,N_15309);
or U18070 (N_18070,N_15747,N_16768);
nand U18071 (N_18071,N_16420,N_15598);
nor U18072 (N_18072,N_15013,N_15653);
nor U18073 (N_18073,N_15814,N_15105);
xnor U18074 (N_18074,N_15272,N_15642);
and U18075 (N_18075,N_15069,N_16389);
or U18076 (N_18076,N_15313,N_15223);
nand U18077 (N_18077,N_15575,N_17383);
or U18078 (N_18078,N_15405,N_16619);
nand U18079 (N_18079,N_15728,N_15581);
or U18080 (N_18080,N_15330,N_17254);
nor U18081 (N_18081,N_16912,N_15659);
nor U18082 (N_18082,N_16979,N_15415);
and U18083 (N_18083,N_16712,N_15137);
xnor U18084 (N_18084,N_15476,N_15641);
and U18085 (N_18085,N_17450,N_15668);
nor U18086 (N_18086,N_17264,N_15429);
nor U18087 (N_18087,N_17211,N_16486);
nor U18088 (N_18088,N_15054,N_16409);
and U18089 (N_18089,N_17027,N_17059);
nand U18090 (N_18090,N_17201,N_16119);
nand U18091 (N_18091,N_16677,N_15325);
nor U18092 (N_18092,N_15163,N_15108);
and U18093 (N_18093,N_16963,N_15249);
or U18094 (N_18094,N_16869,N_15622);
or U18095 (N_18095,N_16339,N_15259);
nand U18096 (N_18096,N_15423,N_15602);
nor U18097 (N_18097,N_16221,N_16892);
nor U18098 (N_18098,N_15218,N_17110);
and U18099 (N_18099,N_15194,N_15327);
xor U18100 (N_18100,N_16564,N_16918);
or U18101 (N_18101,N_17120,N_16448);
nor U18102 (N_18102,N_15450,N_17474);
nand U18103 (N_18103,N_17024,N_17349);
nor U18104 (N_18104,N_16027,N_17398);
xnor U18105 (N_18105,N_16428,N_16421);
or U18106 (N_18106,N_16863,N_15402);
nor U18107 (N_18107,N_15392,N_17150);
or U18108 (N_18108,N_16078,N_17482);
and U18109 (N_18109,N_16539,N_17138);
and U18110 (N_18110,N_16237,N_16771);
xnor U18111 (N_18111,N_15250,N_16670);
or U18112 (N_18112,N_15542,N_15861);
and U18113 (N_18113,N_16549,N_16398);
nor U18114 (N_18114,N_15647,N_17198);
nor U18115 (N_18115,N_15334,N_16352);
nand U18116 (N_18116,N_15328,N_16495);
nor U18117 (N_18117,N_16961,N_16627);
nand U18118 (N_18118,N_16424,N_15087);
nor U18119 (N_18119,N_15740,N_16370);
nor U18120 (N_18120,N_17208,N_15166);
or U18121 (N_18121,N_15241,N_17281);
xor U18122 (N_18122,N_16454,N_17239);
nor U18123 (N_18123,N_16024,N_15317);
xnor U18124 (N_18124,N_15127,N_17114);
or U18125 (N_18125,N_16809,N_17361);
xnor U18126 (N_18126,N_15470,N_17028);
nand U18127 (N_18127,N_15316,N_16069);
or U18128 (N_18128,N_16016,N_15201);
nand U18129 (N_18129,N_16530,N_15600);
or U18130 (N_18130,N_16643,N_15993);
and U18131 (N_18131,N_15403,N_16700);
nand U18132 (N_18132,N_17416,N_16759);
nor U18133 (N_18133,N_16584,N_15550);
or U18134 (N_18134,N_15375,N_16474);
or U18135 (N_18135,N_17072,N_16738);
nor U18136 (N_18136,N_16980,N_15489);
nor U18137 (N_18137,N_16557,N_16778);
or U18138 (N_18138,N_15378,N_16730);
xnor U18139 (N_18139,N_15507,N_17308);
or U18140 (N_18140,N_16175,N_16496);
nand U18141 (N_18141,N_17237,N_16320);
or U18142 (N_18142,N_15499,N_15593);
nor U18143 (N_18143,N_15409,N_16528);
or U18144 (N_18144,N_17345,N_16037);
or U18145 (N_18145,N_16560,N_15269);
nand U18146 (N_18146,N_15459,N_15235);
nand U18147 (N_18147,N_16096,N_16405);
nand U18148 (N_18148,N_15480,N_17457);
and U18149 (N_18149,N_17491,N_16372);
xor U18150 (N_18150,N_15558,N_17399);
and U18151 (N_18151,N_16326,N_16292);
and U18152 (N_18152,N_16180,N_15771);
or U18153 (N_18153,N_17432,N_16546);
and U18154 (N_18154,N_16704,N_16194);
nand U18155 (N_18155,N_16796,N_17188);
nor U18156 (N_18156,N_17005,N_15983);
nor U18157 (N_18157,N_15096,N_15060);
nand U18158 (N_18158,N_15051,N_15217);
or U18159 (N_18159,N_16434,N_17319);
nand U18160 (N_18160,N_16540,N_16684);
xnor U18161 (N_18161,N_16167,N_17129);
or U18162 (N_18162,N_16480,N_15960);
and U18163 (N_18163,N_15455,N_16582);
or U18164 (N_18164,N_15286,N_15339);
and U18165 (N_18165,N_17096,N_17320);
nand U18166 (N_18166,N_17402,N_16874);
xor U18167 (N_18167,N_16596,N_16082);
or U18168 (N_18168,N_16416,N_15145);
nor U18169 (N_18169,N_17276,N_16004);
nand U18170 (N_18170,N_16770,N_17252);
or U18171 (N_18171,N_16506,N_16592);
or U18172 (N_18172,N_15351,N_15953);
nand U18173 (N_18173,N_16621,N_16193);
nor U18174 (N_18174,N_15640,N_15940);
and U18175 (N_18175,N_17219,N_16541);
nand U18176 (N_18176,N_15196,N_15920);
nand U18177 (N_18177,N_15240,N_17107);
and U18178 (N_18178,N_16647,N_16509);
nand U18179 (N_18179,N_15884,N_16698);
nand U18180 (N_18180,N_16419,N_15434);
nand U18181 (N_18181,N_16192,N_17163);
nor U18182 (N_18182,N_16044,N_16142);
xnor U18183 (N_18183,N_16888,N_16639);
or U18184 (N_18184,N_16837,N_15296);
or U18185 (N_18185,N_16975,N_16244);
and U18186 (N_18186,N_16329,N_17226);
nand U18187 (N_18187,N_15465,N_16633);
nor U18188 (N_18188,N_15623,N_15252);
xor U18189 (N_18189,N_15370,N_16870);
or U18190 (N_18190,N_16527,N_16943);
nand U18191 (N_18191,N_17305,N_15978);
or U18192 (N_18192,N_16204,N_16802);
xor U18193 (N_18193,N_16960,N_17108);
and U18194 (N_18194,N_16054,N_15999);
or U18195 (N_18195,N_16673,N_15528);
nand U18196 (N_18196,N_15029,N_16264);
nor U18197 (N_18197,N_15732,N_15585);
and U18198 (N_18198,N_15116,N_15702);
or U18199 (N_18199,N_17065,N_15295);
nor U18200 (N_18200,N_15192,N_16394);
nand U18201 (N_18201,N_17471,N_16751);
nand U18202 (N_18202,N_17481,N_16136);
and U18203 (N_18203,N_17386,N_16910);
nand U18204 (N_18204,N_16253,N_17366);
nand U18205 (N_18205,N_16151,N_15048);
and U18206 (N_18206,N_16571,N_15171);
nand U18207 (N_18207,N_16875,N_15095);
nand U18208 (N_18208,N_16306,N_15354);
nand U18209 (N_18209,N_16513,N_17476);
xnor U18210 (N_18210,N_15021,N_16512);
and U18211 (N_18211,N_16257,N_15928);
nand U18212 (N_18212,N_16949,N_17307);
and U18213 (N_18213,N_16913,N_17409);
nor U18214 (N_18214,N_15644,N_16786);
nand U18215 (N_18215,N_16387,N_15333);
nand U18216 (N_18216,N_17304,N_15982);
nor U18217 (N_18217,N_15388,N_15376);
nand U18218 (N_18218,N_15847,N_16212);
nand U18219 (N_18219,N_16066,N_16106);
xnor U18220 (N_18220,N_17146,N_16568);
or U18221 (N_18221,N_15767,N_15039);
nor U18222 (N_18222,N_15337,N_16517);
and U18223 (N_18223,N_16565,N_15061);
nor U18224 (N_18224,N_15181,N_15377);
nand U18225 (N_18225,N_16040,N_16858);
and U18226 (N_18226,N_16782,N_16605);
or U18227 (N_18227,N_16338,N_15232);
nand U18228 (N_18228,N_16458,N_16607);
nand U18229 (N_18229,N_17173,N_15355);
or U18230 (N_18230,N_17109,N_17164);
nor U18231 (N_18231,N_16903,N_15971);
nand U18232 (N_18232,N_16793,N_15110);
nand U18233 (N_18233,N_15866,N_15150);
or U18234 (N_18234,N_16835,N_17359);
and U18235 (N_18235,N_15961,N_17066);
nor U18236 (N_18236,N_17103,N_16469);
nor U18237 (N_18237,N_16071,N_15075);
and U18238 (N_18238,N_16373,N_17136);
nand U18239 (N_18239,N_15242,N_16731);
nand U18240 (N_18240,N_15532,N_15178);
nand U18241 (N_18241,N_17077,N_15197);
nand U18242 (N_18242,N_17459,N_17183);
xnor U18243 (N_18243,N_17275,N_16997);
nand U18244 (N_18244,N_16551,N_16414);
or U18245 (N_18245,N_16729,N_16840);
nor U18246 (N_18246,N_16335,N_15482);
or U18247 (N_18247,N_17335,N_15128);
or U18248 (N_18248,N_15184,N_17010);
and U18249 (N_18249,N_16334,N_16269);
or U18250 (N_18250,N_17475,N_17265);
or U18251 (N_18251,N_17161,N_16332);
nand U18252 (N_18252,N_16317,N_16107);
xor U18253 (N_18253,N_16976,N_16013);
xnor U18254 (N_18254,N_16182,N_15899);
nor U18255 (N_18255,N_16521,N_16626);
nor U18256 (N_18256,N_15735,N_15386);
xnor U18257 (N_18257,N_15180,N_15678);
nand U18258 (N_18258,N_15366,N_15583);
and U18259 (N_18259,N_16483,N_16794);
and U18260 (N_18260,N_16848,N_16172);
and U18261 (N_18261,N_15170,N_16905);
nor U18262 (N_18262,N_15342,N_17467);
xor U18263 (N_18263,N_15691,N_15510);
or U18264 (N_18264,N_16468,N_16384);
or U18265 (N_18265,N_16138,N_16580);
and U18266 (N_18266,N_17154,N_17466);
and U18267 (N_18267,N_15713,N_16553);
or U18268 (N_18268,N_15154,N_16470);
and U18269 (N_18269,N_15524,N_15157);
or U18270 (N_18270,N_15387,N_15915);
and U18271 (N_18271,N_16534,N_16437);
nand U18272 (N_18272,N_17470,N_15253);
or U18273 (N_18273,N_15825,N_15427);
nand U18274 (N_18274,N_17364,N_15770);
nand U18275 (N_18275,N_16308,N_16817);
nor U18276 (N_18276,N_16969,N_17171);
xor U18277 (N_18277,N_15977,N_15588);
and U18278 (N_18278,N_15117,N_17190);
nand U18279 (N_18279,N_17085,N_16563);
nand U18280 (N_18280,N_15372,N_16651);
and U18281 (N_18281,N_15331,N_16925);
or U18282 (N_18282,N_16276,N_16660);
nor U18283 (N_18283,N_16341,N_16908);
or U18284 (N_18284,N_16755,N_15103);
and U18285 (N_18285,N_16598,N_16857);
or U18286 (N_18286,N_15022,N_15576);
nor U18287 (N_18287,N_15841,N_15262);
nand U18288 (N_18288,N_16139,N_15829);
and U18289 (N_18289,N_15897,N_16795);
or U18290 (N_18290,N_16314,N_17382);
or U18291 (N_18291,N_15618,N_16157);
or U18292 (N_18292,N_15627,N_15854);
or U18293 (N_18293,N_16114,N_16806);
nand U18294 (N_18294,N_15009,N_17492);
xor U18295 (N_18295,N_15683,N_17277);
or U18296 (N_18296,N_15135,N_15613);
and U18297 (N_18297,N_15457,N_15237);
nand U18298 (N_18298,N_15819,N_15951);
nor U18299 (N_18299,N_17283,N_17356);
nand U18300 (N_18300,N_16444,N_16725);
nor U18301 (N_18301,N_16039,N_16266);
and U18302 (N_18302,N_16246,N_17224);
or U18303 (N_18303,N_16048,N_16488);
and U18304 (N_18304,N_16577,N_15134);
or U18305 (N_18305,N_15810,N_16003);
nor U18306 (N_18306,N_16764,N_15025);
and U18307 (N_18307,N_15786,N_15631);
nand U18308 (N_18308,N_17478,N_15363);
nor U18309 (N_18309,N_16953,N_15416);
nor U18310 (N_18310,N_15656,N_16536);
nor U18311 (N_18311,N_15590,N_16641);
xnor U18312 (N_18312,N_15615,N_17159);
nand U18313 (N_18313,N_16247,N_15794);
or U18314 (N_18314,N_15671,N_15790);
and U18315 (N_18315,N_16737,N_15273);
nand U18316 (N_18316,N_17327,N_16316);
nand U18317 (N_18317,N_15301,N_17415);
nand U18318 (N_18318,N_15734,N_16035);
and U18319 (N_18319,N_17145,N_16707);
and U18320 (N_18320,N_16202,N_15173);
nand U18321 (N_18321,N_17214,N_15974);
nor U18322 (N_18322,N_17177,N_17298);
nor U18323 (N_18323,N_16422,N_15870);
or U18324 (N_18324,N_16784,N_15605);
nand U18325 (N_18325,N_17393,N_15537);
and U18326 (N_18326,N_16117,N_17015);
or U18327 (N_18327,N_15102,N_16140);
or U18328 (N_18328,N_16404,N_15785);
xnor U18329 (N_18329,N_16842,N_15293);
and U18330 (N_18330,N_15898,N_16498);
or U18331 (N_18331,N_17093,N_17322);
or U18332 (N_18332,N_16141,N_16061);
nor U18333 (N_18333,N_16554,N_17437);
and U18334 (N_18334,N_16922,N_16510);
and U18335 (N_18335,N_17155,N_15806);
nand U18336 (N_18336,N_15018,N_15721);
nand U18337 (N_18337,N_16611,N_15754);
nand U18338 (N_18338,N_16206,N_16501);
or U18339 (N_18339,N_17369,N_16041);
or U18340 (N_18340,N_15855,N_15751);
or U18341 (N_18341,N_16988,N_17313);
or U18342 (N_18342,N_17329,N_15310);
nand U18343 (N_18343,N_15809,N_17427);
nand U18344 (N_18344,N_16328,N_15692);
nor U18345 (N_18345,N_17302,N_15849);
nand U18346 (N_18346,N_16594,N_15501);
nand U18347 (N_18347,N_16736,N_15690);
xnor U18348 (N_18348,N_16664,N_16826);
nor U18349 (N_18349,N_16238,N_16995);
or U18350 (N_18350,N_15300,N_16694);
or U18351 (N_18351,N_15745,N_16011);
and U18352 (N_18352,N_17269,N_16029);
or U18353 (N_18353,N_16392,N_17166);
or U18354 (N_18354,N_17255,N_15970);
or U18355 (N_18355,N_15338,N_15215);
nor U18356 (N_18356,N_16709,N_15230);
or U18357 (N_18357,N_15084,N_16883);
and U18358 (N_18358,N_16144,N_16025);
nand U18359 (N_18359,N_15212,N_17112);
nor U18360 (N_18360,N_16374,N_16345);
nand U18361 (N_18361,N_15195,N_16750);
nand U18362 (N_18362,N_16785,N_16547);
and U18363 (N_18363,N_16808,N_16998);
or U18364 (N_18364,N_15807,N_15139);
or U18365 (N_18365,N_16649,N_16026);
and U18366 (N_18366,N_15350,N_16418);
or U18367 (N_18367,N_15397,N_16423);
nand U18368 (N_18368,N_16197,N_15290);
xnor U18369 (N_18369,N_16683,N_15912);
and U18370 (N_18370,N_15984,N_15731);
xor U18371 (N_18371,N_17372,N_16031);
and U18372 (N_18372,N_16871,N_15112);
and U18373 (N_18373,N_17423,N_17243);
and U18374 (N_18374,N_15222,N_16340);
nand U18375 (N_18375,N_16529,N_16791);
nor U18376 (N_18376,N_16397,N_16679);
and U18377 (N_18377,N_15299,N_16762);
or U18378 (N_18378,N_16503,N_16100);
and U18379 (N_18379,N_16852,N_15966);
nand U18380 (N_18380,N_16127,N_16805);
nand U18381 (N_18381,N_15506,N_15895);
and U18382 (N_18382,N_15868,N_16505);
or U18383 (N_18383,N_17004,N_15826);
and U18384 (N_18384,N_15074,N_15626);
nand U18385 (N_18385,N_16325,N_15130);
nor U18386 (N_18386,N_17228,N_17225);
nand U18387 (N_18387,N_16944,N_17196);
or U18388 (N_18388,N_15495,N_15509);
nand U18389 (N_18389,N_15315,N_16093);
and U18390 (N_18390,N_15001,N_16964);
nor U18391 (N_18391,N_16661,N_17338);
nand U18392 (N_18392,N_15726,N_15562);
nand U18393 (N_18393,N_15952,N_15633);
and U18394 (N_18394,N_15650,N_16508);
nor U18395 (N_18395,N_17011,N_16049);
or U18396 (N_18396,N_16672,N_15391);
nand U18397 (N_18397,N_15729,N_16482);
and U18398 (N_18398,N_17053,N_16288);
and U18399 (N_18399,N_16904,N_15763);
and U18400 (N_18400,N_16359,N_15680);
nand U18401 (N_18401,N_17391,N_16220);
or U18402 (N_18402,N_15848,N_17003);
xnor U18403 (N_18403,N_17001,N_16703);
and U18404 (N_18404,N_15002,N_16962);
nand U18405 (N_18405,N_16902,N_16134);
and U18406 (N_18406,N_17401,N_15871);
and U18407 (N_18407,N_15321,N_15439);
nor U18408 (N_18408,N_17380,N_16982);
and U18409 (N_18409,N_15228,N_16958);
or U18410 (N_18410,N_16302,N_17377);
nor U18411 (N_18411,N_16146,N_16053);
or U18412 (N_18412,N_16268,N_15044);
and U18413 (N_18413,N_17486,N_17392);
nand U18414 (N_18414,N_15652,N_16933);
or U18415 (N_18415,N_16262,N_16471);
nand U18416 (N_18416,N_16524,N_16075);
nor U18417 (N_18417,N_15812,N_15730);
or U18418 (N_18418,N_15500,N_15446);
and U18419 (N_18419,N_17330,N_16475);
and U18420 (N_18420,N_15004,N_15603);
or U18421 (N_18421,N_15101,N_16590);
nand U18422 (N_18422,N_16839,N_15345);
nand U18423 (N_18423,N_15935,N_17411);
nor U18424 (N_18424,N_15808,N_16831);
or U18425 (N_18425,N_15280,N_16578);
and U18426 (N_18426,N_16893,N_15979);
nand U18427 (N_18427,N_15858,N_15288);
nor U18428 (N_18428,N_16934,N_16899);
nand U18429 (N_18429,N_17040,N_15049);
nor U18430 (N_18430,N_16659,N_16298);
or U18431 (N_18431,N_16453,N_16181);
and U18432 (N_18432,N_15078,N_15346);
nor U18433 (N_18433,N_16526,N_15556);
nand U18434 (N_18434,N_15323,N_15287);
nor U18435 (N_18435,N_15910,N_16593);
nand U18436 (N_18436,N_17350,N_17328);
nor U18437 (N_18437,N_15838,N_15477);
xor U18438 (N_18438,N_17468,N_16051);
or U18439 (N_18439,N_16466,N_16853);
or U18440 (N_18440,N_16073,N_15142);
xor U18441 (N_18441,N_15067,N_16946);
nand U18442 (N_18442,N_17054,N_16301);
and U18443 (N_18443,N_16176,N_17296);
nor U18444 (N_18444,N_15040,N_16556);
nand U18445 (N_18445,N_16585,N_17174);
and U18446 (N_18446,N_17097,N_15035);
or U18447 (N_18447,N_16425,N_17376);
and U18448 (N_18448,N_16440,N_16929);
and U18449 (N_18449,N_16493,N_17185);
nand U18450 (N_18450,N_17477,N_16309);
or U18451 (N_18451,N_15151,N_15705);
nor U18452 (N_18452,N_15502,N_15297);
or U18453 (N_18453,N_16678,N_16435);
nor U18454 (N_18454,N_16210,N_15563);
nand U18455 (N_18455,N_16021,N_17438);
nand U18456 (N_18456,N_17067,N_15123);
or U18457 (N_18457,N_15522,N_16086);
or U18458 (N_18458,N_15267,N_16781);
nor U18459 (N_18459,N_15514,N_17031);
nor U18460 (N_18460,N_17037,N_15718);
xnor U18461 (N_18461,N_16331,N_16692);
nand U18462 (N_18462,N_16427,N_15085);
nand U18463 (N_18463,N_16543,N_15635);
nor U18464 (N_18464,N_16847,N_15911);
or U18465 (N_18465,N_17218,N_15220);
and U18466 (N_18466,N_17168,N_16640);
nand U18467 (N_18467,N_15727,N_15608);
and U18468 (N_18468,N_15208,N_17060);
or U18469 (N_18469,N_15420,N_17424);
nand U18470 (N_18470,N_17215,N_15205);
and U18471 (N_18471,N_16231,N_15068);
or U18472 (N_18472,N_15052,N_15141);
and U18473 (N_18473,N_15193,N_17274);
or U18474 (N_18474,N_15125,N_16494);
or U18475 (N_18475,N_15926,N_16249);
or U18476 (N_18476,N_15245,N_16603);
and U18477 (N_18477,N_15129,N_17197);
xor U18478 (N_18478,N_15277,N_17035);
or U18479 (N_18479,N_15298,N_16981);
or U18480 (N_18480,N_15050,N_17355);
or U18481 (N_18481,N_15199,N_16657);
nor U18482 (N_18482,N_16803,N_15798);
and U18483 (N_18483,N_15701,N_16972);
and U18484 (N_18484,N_15410,N_16386);
nor U18485 (N_18485,N_15019,N_15448);
and U18486 (N_18486,N_16812,N_15177);
and U18487 (N_18487,N_16956,N_16974);
xor U18488 (N_18488,N_15707,N_16911);
and U18489 (N_18489,N_17025,N_16191);
nor U18490 (N_18490,N_16380,N_16715);
or U18491 (N_18491,N_16233,N_16413);
or U18492 (N_18492,N_16012,N_15168);
xnor U18493 (N_18493,N_16717,N_16650);
and U18494 (N_18494,N_16939,N_17049);
nor U18495 (N_18495,N_15634,N_15595);
and U18496 (N_18496,N_16936,N_15206);
nand U18497 (N_18497,N_17293,N_16990);
or U18498 (N_18498,N_15568,N_17184);
and U18499 (N_18499,N_15791,N_17247);
or U18500 (N_18500,N_15630,N_17271);
and U18501 (N_18501,N_17105,N_15059);
or U18502 (N_18502,N_16941,N_15461);
or U18503 (N_18503,N_16535,N_15020);
or U18504 (N_18504,N_15183,N_17321);
and U18505 (N_18505,N_15224,N_17139);
nand U18506 (N_18506,N_17270,N_15227);
nand U18507 (N_18507,N_15503,N_15879);
xor U18508 (N_18508,N_15875,N_15072);
and U18509 (N_18509,N_17057,N_16987);
nor U18510 (N_18510,N_15839,N_17433);
and U18511 (N_18511,N_15724,N_16558);
and U18512 (N_18512,N_16843,N_17023);
or U18513 (N_18513,N_16531,N_16105);
nor U18514 (N_18514,N_16952,N_16113);
nor U18515 (N_18515,N_17143,N_15456);
xnor U18516 (N_18516,N_17299,N_15107);
xnor U18517 (N_18517,N_15736,N_16395);
nand U18518 (N_18518,N_17238,N_16685);
and U18519 (N_18519,N_15062,N_15843);
nand U18520 (N_18520,N_16518,N_16005);
nor U18521 (N_18521,N_16135,N_15374);
nand U18522 (N_18522,N_16121,N_15549);
xor U18523 (N_18523,N_17086,N_16890);
nand U18524 (N_18524,N_15827,N_16452);
nand U18525 (N_18525,N_15566,N_16109);
nand U18526 (N_18526,N_16734,N_15780);
or U18527 (N_18527,N_16575,N_16094);
or U18528 (N_18528,N_15620,N_16222);
nand U18529 (N_18529,N_15698,N_17019);
xnor U18530 (N_18530,N_16516,N_15693);
nor U18531 (N_18531,N_17008,N_15577);
xor U18532 (N_18532,N_15675,N_15560);
nor U18533 (N_18533,N_15381,N_15743);
or U18534 (N_18534,N_16945,N_15254);
nor U18535 (N_18535,N_15990,N_16156);
or U18536 (N_18536,N_16723,N_16994);
nor U18537 (N_18537,N_16774,N_17202);
nor U18538 (N_18538,N_16343,N_15200);
or U18539 (N_18539,N_16984,N_16855);
nor U18540 (N_18540,N_15753,N_17124);
or U18541 (N_18541,N_17246,N_17162);
nand U18542 (N_18542,N_17034,N_15804);
nand U18543 (N_18543,N_17285,N_15824);
nor U18544 (N_18544,N_17233,N_16084);
or U18545 (N_18545,N_16900,N_16315);
and U18546 (N_18546,N_15158,N_16790);
xor U18547 (N_18547,N_15991,N_15365);
and U18548 (N_18548,N_16914,N_16867);
or U18549 (N_18549,N_15933,N_16007);
nor U18550 (N_18550,N_15828,N_15143);
or U18551 (N_18551,N_15445,N_15629);
nand U18552 (N_18552,N_17220,N_17007);
xor U18553 (N_18553,N_16438,N_16209);
nand U18554 (N_18554,N_16363,N_16396);
or U18555 (N_18555,N_16733,N_15850);
or U18556 (N_18556,N_15779,N_16947);
xor U18557 (N_18557,N_16200,N_15188);
nand U18558 (N_18558,N_17284,N_15591);
nand U18559 (N_18559,N_17153,N_16230);
nand U18560 (N_18560,N_17451,N_16533);
and U18561 (N_18561,N_17291,N_17055);
nor U18562 (N_18562,N_15793,N_17076);
nand U18563 (N_18563,N_15098,N_17134);
nor U18564 (N_18564,N_15569,N_17339);
nor U18565 (N_18565,N_15100,N_15989);
and U18566 (N_18566,N_16273,N_16884);
nand U18567 (N_18567,N_15967,N_17484);
or U18568 (N_18568,N_16951,N_17394);
xnor U18569 (N_18569,N_16609,N_15582);
nor U18570 (N_18570,N_16954,N_16777);
nand U18571 (N_18571,N_15820,N_16693);
nand U18572 (N_18572,N_15512,N_15852);
nand U18573 (N_18573,N_15681,N_15204);
xor U18574 (N_18574,N_16894,N_15795);
xor U18575 (N_18575,N_15088,N_16610);
or U18576 (N_18576,N_16058,N_15948);
xor U18577 (N_18577,N_15394,N_17167);
and U18578 (N_18578,N_16410,N_16674);
xnor U18579 (N_18579,N_17137,N_17223);
nand U18580 (N_18580,N_16663,N_17069);
and U18581 (N_18581,N_16520,N_17000);
and U18582 (N_18582,N_16708,N_16252);
nand U18583 (N_18583,N_17045,N_16522);
nor U18584 (N_18584,N_17018,N_15525);
nand U18585 (N_18585,N_16758,N_15243);
or U18586 (N_18586,N_16525,N_16234);
xnor U18587 (N_18587,N_16190,N_16283);
xnor U18588 (N_18588,N_16279,N_16383);
xor U18589 (N_18589,N_17479,N_16889);
nand U18590 (N_18590,N_15571,N_16277);
or U18591 (N_18591,N_17413,N_15863);
and U18592 (N_18592,N_16361,N_16915);
xor U18593 (N_18593,N_16278,N_16145);
nor U18594 (N_18594,N_15676,N_16644);
xor U18595 (N_18595,N_17443,N_16010);
nand U18596 (N_18596,N_16239,N_16620);
xor U18597 (N_18597,N_16741,N_15233);
and U18598 (N_18598,N_17260,N_17002);
and U18599 (N_18599,N_15902,N_17156);
or U18600 (N_18600,N_16173,N_16006);
xor U18601 (N_18601,N_16742,N_16787);
nor U18602 (N_18602,N_16371,N_16601);
nand U18603 (N_18603,N_15746,N_15845);
or U18604 (N_18604,N_17189,N_17232);
and U18605 (N_18605,N_15817,N_15513);
and U18606 (N_18606,N_17495,N_17463);
or U18607 (N_18607,N_15986,N_17210);
or U18608 (N_18608,N_16207,N_15454);
nor U18609 (N_18609,N_16169,N_15441);
nand U18610 (N_18610,N_16362,N_16046);
xor U18611 (N_18611,N_16382,N_16957);
or U18612 (N_18612,N_16511,N_15369);
and U18613 (N_18613,N_15654,N_16701);
nor U18614 (N_18614,N_15453,N_15015);
and U18615 (N_18615,N_16967,N_17429);
nor U18616 (N_18616,N_15816,N_17199);
or U18617 (N_18617,N_16311,N_17297);
or U18618 (N_18618,N_17442,N_16216);
or U18619 (N_18619,N_16052,N_16218);
nand U18620 (N_18620,N_16017,N_17436);
nand U18621 (N_18621,N_16154,N_16215);
nand U18622 (N_18622,N_16849,N_15426);
nor U18623 (N_18623,N_16537,N_17282);
nor U18624 (N_18624,N_15490,N_15526);
and U18625 (N_18625,N_16337,N_15756);
or U18626 (N_18626,N_16198,N_16695);
and U18627 (N_18627,N_15545,N_17227);
nor U18628 (N_18628,N_15881,N_15689);
xor U18629 (N_18629,N_15521,N_15079);
or U18630 (N_18630,N_17135,N_16402);
and U18631 (N_18631,N_16612,N_16932);
nand U18632 (N_18632,N_16566,N_17456);
nor U18633 (N_18633,N_16439,N_16060);
nor U18634 (N_18634,N_16324,N_15468);
nand U18635 (N_18635,N_15636,N_16000);
and U18636 (N_18636,N_17397,N_16490);
nand U18637 (N_18637,N_17384,N_15973);
and U18638 (N_18638,N_15191,N_16628);
nor U18639 (N_18639,N_15530,N_17181);
nor U18640 (N_18640,N_16638,N_16671);
nand U18641 (N_18641,N_17070,N_15609);
or U18642 (N_18642,N_17373,N_16686);
and U18643 (N_18643,N_16570,N_15894);
or U18644 (N_18644,N_16367,N_15892);
and U18645 (N_18645,N_17221,N_15909);
or U18646 (N_18646,N_16631,N_17336);
and U18647 (N_18647,N_16477,N_16303);
or U18648 (N_18648,N_16111,N_15203);
or U18649 (N_18649,N_15570,N_15364);
nand U18650 (N_18650,N_16800,N_17176);
xor U18651 (N_18651,N_15846,N_16996);
nor U18652 (N_18652,N_16572,N_17095);
nor U18653 (N_18653,N_15837,N_16001);
or U18654 (N_18654,N_16242,N_16417);
and U18655 (N_18655,N_16385,N_16330);
nor U18656 (N_18656,N_16355,N_15368);
nor U18657 (N_18657,N_15285,N_15413);
nor U18658 (N_18658,N_15097,N_15907);
nand U18659 (N_18659,N_15486,N_15723);
nor U18660 (N_18660,N_16484,N_15540);
or U18661 (N_18661,N_15704,N_15341);
nand U18662 (N_18662,N_15818,N_15417);
and U18663 (N_18663,N_15030,N_15769);
nor U18664 (N_18664,N_17012,N_17496);
nor U18665 (N_18665,N_16098,N_16667);
nand U18666 (N_18666,N_16376,N_15396);
and U18667 (N_18667,N_17455,N_17100);
and U18668 (N_18668,N_17013,N_15553);
and U18669 (N_18669,N_15132,N_17106);
nor U18670 (N_18670,N_15888,N_16637);
or U18671 (N_18671,N_17102,N_16293);
nor U18672 (N_18672,N_15303,N_15362);
and U18673 (N_18673,N_15395,N_17250);
and U18674 (N_18674,N_15880,N_16948);
xor U18675 (N_18675,N_16377,N_15380);
and U18676 (N_18676,N_16313,N_17186);
nor U18677 (N_18677,N_16872,N_16360);
and U18678 (N_18678,N_16455,N_16616);
or U18679 (N_18679,N_17396,N_15185);
xor U18680 (N_18680,N_15024,N_16348);
and U18681 (N_18681,N_16599,N_15945);
and U18682 (N_18682,N_15596,N_15348);
and U18683 (N_18683,N_16523,N_16166);
nor U18684 (N_18684,N_16103,N_15876);
nand U18685 (N_18685,N_15802,N_16240);
nand U18686 (N_18686,N_16959,N_15042);
or U18687 (N_18687,N_16487,N_15076);
or U18688 (N_18688,N_17365,N_16147);
or U18689 (N_18689,N_16129,N_16588);
xnor U18690 (N_18690,N_15766,N_16829);
and U18691 (N_18691,N_17445,N_15857);
xor U18692 (N_18692,N_16195,N_16045);
nand U18693 (N_18693,N_16074,N_15431);
or U18694 (N_18694,N_16828,N_16184);
nand U18695 (N_18695,N_15198,N_15905);
nor U18696 (N_18696,N_16985,N_17342);
nor U18697 (N_18697,N_16415,N_15373);
nand U18698 (N_18698,N_17301,N_15153);
and U18699 (N_18699,N_15347,N_16108);
nand U18700 (N_18700,N_16942,N_17303);
nand U18701 (N_18701,N_15264,N_16940);
and U18702 (N_18702,N_15311,N_16346);
nand U18703 (N_18703,N_16901,N_16047);
xor U18704 (N_18704,N_17234,N_15696);
nor U18705 (N_18705,N_16368,N_16801);
nand U18706 (N_18706,N_16753,N_15408);
and U18707 (N_18707,N_16030,N_16171);
nor U18708 (N_18708,N_15246,N_16859);
or U18709 (N_18709,N_15717,N_16126);
nor U18710 (N_18710,N_17418,N_16879);
or U18711 (N_18711,N_16133,N_16118);
nor U18712 (N_18712,N_15830,N_15289);
and U18713 (N_18713,N_15422,N_17323);
or U18714 (N_18714,N_16403,N_15918);
nand U18715 (N_18715,N_17414,N_17315);
or U18716 (N_18716,N_17116,N_17343);
and U18717 (N_18717,N_16063,N_15471);
nor U18718 (N_18718,N_16682,N_17140);
nand U18719 (N_18719,N_15529,N_16179);
nand U18720 (N_18720,N_15955,N_15063);
and U18721 (N_18721,N_15733,N_16072);
nand U18722 (N_18722,N_16083,N_16622);
or U18723 (N_18723,N_16642,N_15466);
or U18724 (N_18724,N_17016,N_17417);
nor U18725 (N_18725,N_16481,N_16254);
nand U18726 (N_18726,N_16463,N_17151);
or U18727 (N_18727,N_15111,N_15118);
or U18728 (N_18728,N_15950,N_15711);
nand U18729 (N_18729,N_17206,N_17494);
and U18730 (N_18730,N_16203,N_15283);
nand U18731 (N_18731,N_15660,N_15302);
nor U18732 (N_18732,N_16896,N_16732);
or U18733 (N_18733,N_17160,N_17048);
nor U18734 (N_18734,N_16978,N_16426);
and U18735 (N_18735,N_15765,N_16775);
nand U18736 (N_18736,N_17352,N_16779);
or U18737 (N_18737,N_17063,N_17115);
xnor U18738 (N_18738,N_15257,N_16993);
and U18739 (N_18739,N_17050,N_16792);
nand U18740 (N_18740,N_15896,N_16491);
nand U18741 (N_18741,N_16472,N_15258);
nand U18742 (N_18742,N_15278,N_15336);
and U18743 (N_18743,N_15811,N_15755);
nor U18744 (N_18744,N_16675,N_15700);
nor U18745 (N_18745,N_17331,N_16125);
or U18746 (N_18746,N_16080,N_16666);
nor U18747 (N_18747,N_16600,N_15014);
nor U18748 (N_18748,N_16090,N_15959);
and U18749 (N_18749,N_17165,N_15398);
nor U18750 (N_18750,N_17159,N_15236);
xnor U18751 (N_18751,N_16633,N_16189);
nor U18752 (N_18752,N_16665,N_17365);
and U18753 (N_18753,N_16708,N_16740);
nand U18754 (N_18754,N_17249,N_16268);
and U18755 (N_18755,N_16716,N_16794);
nand U18756 (N_18756,N_17325,N_16689);
nor U18757 (N_18757,N_16161,N_16274);
xnor U18758 (N_18758,N_15237,N_16915);
nor U18759 (N_18759,N_16382,N_15829);
xor U18760 (N_18760,N_16362,N_16115);
nand U18761 (N_18761,N_15512,N_16482);
nor U18762 (N_18762,N_17104,N_16611);
nand U18763 (N_18763,N_16604,N_16147);
nor U18764 (N_18764,N_15252,N_16714);
or U18765 (N_18765,N_15852,N_17030);
or U18766 (N_18766,N_16423,N_15607);
nor U18767 (N_18767,N_15532,N_17151);
or U18768 (N_18768,N_15898,N_15186);
and U18769 (N_18769,N_15966,N_16936);
or U18770 (N_18770,N_17259,N_17424);
or U18771 (N_18771,N_16191,N_17136);
or U18772 (N_18772,N_15805,N_16418);
nand U18773 (N_18773,N_16990,N_16684);
or U18774 (N_18774,N_15685,N_16003);
nand U18775 (N_18775,N_16474,N_16692);
nor U18776 (N_18776,N_15926,N_16955);
nand U18777 (N_18777,N_16520,N_16409);
and U18778 (N_18778,N_16132,N_16882);
or U18779 (N_18779,N_16076,N_16874);
nand U18780 (N_18780,N_15980,N_16269);
or U18781 (N_18781,N_16535,N_15301);
or U18782 (N_18782,N_16765,N_17371);
and U18783 (N_18783,N_15227,N_15507);
nand U18784 (N_18784,N_15996,N_16007);
and U18785 (N_18785,N_16346,N_16983);
and U18786 (N_18786,N_17163,N_16953);
nand U18787 (N_18787,N_15801,N_17416);
and U18788 (N_18788,N_17166,N_17221);
nand U18789 (N_18789,N_16172,N_15916);
nand U18790 (N_18790,N_15060,N_16242);
and U18791 (N_18791,N_15701,N_15534);
nand U18792 (N_18792,N_16054,N_16238);
and U18793 (N_18793,N_17491,N_15340);
and U18794 (N_18794,N_17192,N_16906);
or U18795 (N_18795,N_16023,N_16106);
nand U18796 (N_18796,N_15713,N_16504);
nand U18797 (N_18797,N_16259,N_16363);
nand U18798 (N_18798,N_15433,N_15281);
or U18799 (N_18799,N_16159,N_17201);
and U18800 (N_18800,N_16907,N_15125);
or U18801 (N_18801,N_15409,N_15620);
nand U18802 (N_18802,N_16552,N_15843);
or U18803 (N_18803,N_15771,N_15291);
or U18804 (N_18804,N_15465,N_17246);
or U18805 (N_18805,N_15469,N_16865);
nand U18806 (N_18806,N_17043,N_15809);
nor U18807 (N_18807,N_15203,N_17171);
nand U18808 (N_18808,N_15925,N_17354);
and U18809 (N_18809,N_16293,N_16226);
and U18810 (N_18810,N_15901,N_17093);
and U18811 (N_18811,N_15867,N_15377);
and U18812 (N_18812,N_17214,N_16712);
or U18813 (N_18813,N_16634,N_17334);
and U18814 (N_18814,N_15535,N_16971);
xnor U18815 (N_18815,N_15021,N_16145);
nor U18816 (N_18816,N_16745,N_15179);
and U18817 (N_18817,N_15245,N_16334);
nand U18818 (N_18818,N_16219,N_15930);
and U18819 (N_18819,N_15101,N_16361);
and U18820 (N_18820,N_17235,N_16004);
or U18821 (N_18821,N_15474,N_16876);
xnor U18822 (N_18822,N_16414,N_16578);
xnor U18823 (N_18823,N_16660,N_15859);
nor U18824 (N_18824,N_16311,N_17269);
or U18825 (N_18825,N_16390,N_17148);
nand U18826 (N_18826,N_17016,N_17272);
or U18827 (N_18827,N_16299,N_16791);
nand U18828 (N_18828,N_15471,N_17455);
nand U18829 (N_18829,N_15401,N_16418);
nand U18830 (N_18830,N_15866,N_17367);
and U18831 (N_18831,N_15580,N_15386);
nor U18832 (N_18832,N_17044,N_17389);
nand U18833 (N_18833,N_16838,N_15568);
nor U18834 (N_18834,N_17030,N_17207);
xnor U18835 (N_18835,N_17172,N_17057);
or U18836 (N_18836,N_15249,N_15455);
or U18837 (N_18837,N_15619,N_15533);
and U18838 (N_18838,N_16187,N_16509);
nand U18839 (N_18839,N_17120,N_15646);
nand U18840 (N_18840,N_17012,N_15469);
xnor U18841 (N_18841,N_15487,N_17476);
nand U18842 (N_18842,N_16369,N_16050);
nor U18843 (N_18843,N_16142,N_15151);
nand U18844 (N_18844,N_16534,N_15910);
and U18845 (N_18845,N_15331,N_16251);
nand U18846 (N_18846,N_15220,N_17179);
and U18847 (N_18847,N_15010,N_17057);
xor U18848 (N_18848,N_17498,N_15998);
xnor U18849 (N_18849,N_17170,N_15789);
xnor U18850 (N_18850,N_17483,N_15848);
and U18851 (N_18851,N_16586,N_15054);
and U18852 (N_18852,N_16743,N_15093);
and U18853 (N_18853,N_15025,N_16553);
or U18854 (N_18854,N_17040,N_17261);
or U18855 (N_18855,N_15040,N_16259);
nand U18856 (N_18856,N_16618,N_15543);
nand U18857 (N_18857,N_15080,N_16286);
nor U18858 (N_18858,N_17248,N_16260);
or U18859 (N_18859,N_15912,N_15878);
and U18860 (N_18860,N_15974,N_17028);
xnor U18861 (N_18861,N_17209,N_16232);
nand U18862 (N_18862,N_15434,N_15545);
xor U18863 (N_18863,N_17032,N_16723);
or U18864 (N_18864,N_17162,N_15759);
nand U18865 (N_18865,N_16205,N_15645);
xor U18866 (N_18866,N_16706,N_17237);
nor U18867 (N_18867,N_15968,N_16790);
or U18868 (N_18868,N_16235,N_15415);
and U18869 (N_18869,N_15553,N_16199);
or U18870 (N_18870,N_17467,N_15921);
and U18871 (N_18871,N_17341,N_16713);
and U18872 (N_18872,N_16219,N_16715);
xor U18873 (N_18873,N_16252,N_16726);
nand U18874 (N_18874,N_15305,N_17479);
nor U18875 (N_18875,N_16222,N_15247);
nand U18876 (N_18876,N_16844,N_16156);
or U18877 (N_18877,N_16669,N_15876);
nor U18878 (N_18878,N_15962,N_15234);
xnor U18879 (N_18879,N_15346,N_16502);
or U18880 (N_18880,N_17056,N_15254);
nand U18881 (N_18881,N_17402,N_16615);
or U18882 (N_18882,N_16631,N_16172);
nor U18883 (N_18883,N_15171,N_15795);
and U18884 (N_18884,N_15465,N_16743);
nor U18885 (N_18885,N_15839,N_17276);
nor U18886 (N_18886,N_16573,N_15590);
nor U18887 (N_18887,N_15452,N_15351);
nand U18888 (N_18888,N_17131,N_15895);
and U18889 (N_18889,N_16954,N_16040);
xnor U18890 (N_18890,N_16832,N_16950);
nor U18891 (N_18891,N_16744,N_15737);
nor U18892 (N_18892,N_16460,N_16953);
or U18893 (N_18893,N_16913,N_15335);
or U18894 (N_18894,N_15175,N_16352);
xnor U18895 (N_18895,N_17273,N_16809);
or U18896 (N_18896,N_17495,N_15754);
nand U18897 (N_18897,N_15550,N_16105);
and U18898 (N_18898,N_15055,N_17464);
nor U18899 (N_18899,N_16280,N_15458);
xor U18900 (N_18900,N_17274,N_17452);
and U18901 (N_18901,N_15201,N_16581);
or U18902 (N_18902,N_15482,N_17294);
nor U18903 (N_18903,N_16364,N_16787);
nand U18904 (N_18904,N_15622,N_17358);
or U18905 (N_18905,N_16442,N_15513);
nor U18906 (N_18906,N_16185,N_17412);
nand U18907 (N_18907,N_15150,N_16015);
or U18908 (N_18908,N_16431,N_16249);
nor U18909 (N_18909,N_15354,N_15707);
and U18910 (N_18910,N_15941,N_15338);
and U18911 (N_18911,N_16659,N_15992);
and U18912 (N_18912,N_15059,N_17182);
nand U18913 (N_18913,N_15279,N_17296);
nand U18914 (N_18914,N_16486,N_16882);
xnor U18915 (N_18915,N_16781,N_15375);
or U18916 (N_18916,N_16073,N_16532);
and U18917 (N_18917,N_15128,N_16507);
and U18918 (N_18918,N_17092,N_16920);
nor U18919 (N_18919,N_17174,N_17341);
and U18920 (N_18920,N_15406,N_15050);
nor U18921 (N_18921,N_15769,N_15895);
xnor U18922 (N_18922,N_15448,N_15002);
or U18923 (N_18923,N_17473,N_15062);
nor U18924 (N_18924,N_16436,N_16020);
or U18925 (N_18925,N_17169,N_17239);
and U18926 (N_18926,N_16715,N_15724);
and U18927 (N_18927,N_16245,N_15569);
nand U18928 (N_18928,N_17464,N_15992);
or U18929 (N_18929,N_15401,N_17494);
nand U18930 (N_18930,N_16268,N_17005);
nand U18931 (N_18931,N_16109,N_15500);
xnor U18932 (N_18932,N_15587,N_15265);
nor U18933 (N_18933,N_16343,N_16731);
nand U18934 (N_18934,N_16828,N_16792);
nor U18935 (N_18935,N_16861,N_16858);
and U18936 (N_18936,N_15171,N_15432);
and U18937 (N_18937,N_17351,N_17114);
nand U18938 (N_18938,N_16973,N_15581);
xor U18939 (N_18939,N_15460,N_15539);
nor U18940 (N_18940,N_16596,N_17289);
nand U18941 (N_18941,N_17236,N_15141);
nor U18942 (N_18942,N_16089,N_16734);
nand U18943 (N_18943,N_16661,N_15954);
and U18944 (N_18944,N_16397,N_15727);
or U18945 (N_18945,N_16357,N_15560);
nand U18946 (N_18946,N_15458,N_16188);
and U18947 (N_18947,N_15072,N_16266);
and U18948 (N_18948,N_16809,N_15389);
nor U18949 (N_18949,N_15046,N_15781);
nor U18950 (N_18950,N_17384,N_17204);
or U18951 (N_18951,N_15402,N_16086);
or U18952 (N_18952,N_15747,N_17194);
nand U18953 (N_18953,N_17305,N_17101);
nor U18954 (N_18954,N_17200,N_15841);
nand U18955 (N_18955,N_17260,N_15429);
nor U18956 (N_18956,N_15924,N_16685);
and U18957 (N_18957,N_16808,N_16698);
nor U18958 (N_18958,N_17218,N_15613);
nand U18959 (N_18959,N_15980,N_17072);
nand U18960 (N_18960,N_16543,N_15996);
and U18961 (N_18961,N_15193,N_15977);
and U18962 (N_18962,N_17473,N_15613);
nor U18963 (N_18963,N_15596,N_17419);
nor U18964 (N_18964,N_17362,N_16973);
and U18965 (N_18965,N_17429,N_15378);
or U18966 (N_18966,N_15069,N_15181);
nand U18967 (N_18967,N_15324,N_15649);
nand U18968 (N_18968,N_16922,N_15738);
or U18969 (N_18969,N_16504,N_16260);
nand U18970 (N_18970,N_16292,N_16872);
nand U18971 (N_18971,N_16017,N_16502);
nor U18972 (N_18972,N_16151,N_15543);
or U18973 (N_18973,N_16745,N_16226);
nor U18974 (N_18974,N_17432,N_15059);
nor U18975 (N_18975,N_15335,N_17385);
or U18976 (N_18976,N_15704,N_17442);
or U18977 (N_18977,N_15735,N_16962);
xor U18978 (N_18978,N_16408,N_16951);
nor U18979 (N_18979,N_15949,N_15237);
and U18980 (N_18980,N_15292,N_15981);
and U18981 (N_18981,N_15685,N_16903);
nand U18982 (N_18982,N_15944,N_17154);
or U18983 (N_18983,N_17079,N_16805);
nand U18984 (N_18984,N_16884,N_15130);
or U18985 (N_18985,N_17337,N_16569);
and U18986 (N_18986,N_15099,N_17032);
or U18987 (N_18987,N_16087,N_15444);
nand U18988 (N_18988,N_17317,N_15041);
and U18989 (N_18989,N_17237,N_15084);
nor U18990 (N_18990,N_15936,N_16396);
and U18991 (N_18991,N_17371,N_16760);
nand U18992 (N_18992,N_15952,N_15177);
nand U18993 (N_18993,N_17159,N_17284);
or U18994 (N_18994,N_17007,N_16134);
nor U18995 (N_18995,N_16623,N_16523);
nand U18996 (N_18996,N_17447,N_15844);
nor U18997 (N_18997,N_15741,N_16729);
nor U18998 (N_18998,N_15402,N_16257);
or U18999 (N_18999,N_15766,N_15995);
nor U19000 (N_19000,N_16187,N_17317);
or U19001 (N_19001,N_15071,N_16178);
nor U19002 (N_19002,N_17420,N_15505);
or U19003 (N_19003,N_17250,N_15406);
nor U19004 (N_19004,N_15204,N_15283);
and U19005 (N_19005,N_16701,N_17481);
nor U19006 (N_19006,N_16866,N_17309);
and U19007 (N_19007,N_15364,N_15864);
or U19008 (N_19008,N_16131,N_16612);
or U19009 (N_19009,N_15567,N_16878);
or U19010 (N_19010,N_15862,N_15027);
or U19011 (N_19011,N_15147,N_16757);
and U19012 (N_19012,N_15930,N_16016);
nand U19013 (N_19013,N_16436,N_15230);
and U19014 (N_19014,N_16890,N_15954);
and U19015 (N_19015,N_15142,N_16565);
nor U19016 (N_19016,N_16850,N_17222);
or U19017 (N_19017,N_16351,N_16158);
or U19018 (N_19018,N_16541,N_15624);
and U19019 (N_19019,N_15833,N_15762);
and U19020 (N_19020,N_17353,N_16589);
and U19021 (N_19021,N_15481,N_16878);
or U19022 (N_19022,N_16660,N_16994);
xor U19023 (N_19023,N_15735,N_16011);
and U19024 (N_19024,N_17040,N_16645);
nand U19025 (N_19025,N_17060,N_16379);
and U19026 (N_19026,N_16122,N_16772);
nor U19027 (N_19027,N_15046,N_15511);
nand U19028 (N_19028,N_16034,N_16429);
and U19029 (N_19029,N_17476,N_16477);
and U19030 (N_19030,N_15799,N_15855);
xor U19031 (N_19031,N_15460,N_16946);
and U19032 (N_19032,N_15524,N_16256);
nor U19033 (N_19033,N_16821,N_17446);
nor U19034 (N_19034,N_16659,N_15285);
or U19035 (N_19035,N_15447,N_16606);
or U19036 (N_19036,N_15155,N_15906);
or U19037 (N_19037,N_15671,N_15803);
nand U19038 (N_19038,N_16658,N_17495);
or U19039 (N_19039,N_16364,N_17244);
xor U19040 (N_19040,N_15555,N_15859);
nor U19041 (N_19041,N_17406,N_15016);
nand U19042 (N_19042,N_17268,N_17329);
or U19043 (N_19043,N_15811,N_16672);
xnor U19044 (N_19044,N_17348,N_16587);
or U19045 (N_19045,N_16601,N_17385);
nor U19046 (N_19046,N_15909,N_16773);
nand U19047 (N_19047,N_15218,N_16879);
or U19048 (N_19048,N_15808,N_17168);
nand U19049 (N_19049,N_15956,N_17165);
nand U19050 (N_19050,N_15448,N_15949);
nor U19051 (N_19051,N_17335,N_15113);
and U19052 (N_19052,N_15720,N_15129);
or U19053 (N_19053,N_16348,N_16698);
or U19054 (N_19054,N_16283,N_16210);
or U19055 (N_19055,N_16164,N_15674);
and U19056 (N_19056,N_17328,N_17454);
xor U19057 (N_19057,N_16692,N_17243);
nor U19058 (N_19058,N_16426,N_15113);
or U19059 (N_19059,N_15488,N_15889);
nor U19060 (N_19060,N_15831,N_16336);
or U19061 (N_19061,N_15247,N_16361);
and U19062 (N_19062,N_15199,N_15749);
nor U19063 (N_19063,N_15922,N_16540);
or U19064 (N_19064,N_16635,N_17365);
nand U19065 (N_19065,N_15467,N_17437);
or U19066 (N_19066,N_15567,N_15058);
and U19067 (N_19067,N_16773,N_16733);
nand U19068 (N_19068,N_16450,N_17159);
nand U19069 (N_19069,N_15476,N_16366);
nor U19070 (N_19070,N_15437,N_16811);
xnor U19071 (N_19071,N_16548,N_16892);
and U19072 (N_19072,N_17482,N_16967);
xnor U19073 (N_19073,N_16813,N_15141);
or U19074 (N_19074,N_17232,N_16162);
nand U19075 (N_19075,N_16895,N_16045);
nor U19076 (N_19076,N_16346,N_16500);
nand U19077 (N_19077,N_15747,N_16580);
nor U19078 (N_19078,N_17381,N_15174);
nor U19079 (N_19079,N_17261,N_15783);
nand U19080 (N_19080,N_17252,N_15572);
nor U19081 (N_19081,N_15589,N_15245);
or U19082 (N_19082,N_15972,N_15216);
or U19083 (N_19083,N_15446,N_17126);
xor U19084 (N_19084,N_15882,N_15326);
nor U19085 (N_19085,N_15265,N_15988);
xor U19086 (N_19086,N_17480,N_15049);
and U19087 (N_19087,N_16225,N_17371);
nand U19088 (N_19088,N_15009,N_15652);
or U19089 (N_19089,N_15415,N_16830);
or U19090 (N_19090,N_16291,N_16154);
nor U19091 (N_19091,N_15638,N_16993);
nor U19092 (N_19092,N_16137,N_15792);
and U19093 (N_19093,N_16583,N_15408);
or U19094 (N_19094,N_17039,N_16334);
or U19095 (N_19095,N_16312,N_16792);
and U19096 (N_19096,N_16315,N_16496);
or U19097 (N_19097,N_16430,N_17459);
xor U19098 (N_19098,N_17006,N_16995);
nor U19099 (N_19099,N_16868,N_17429);
nand U19100 (N_19100,N_17286,N_16740);
nand U19101 (N_19101,N_16316,N_15122);
nor U19102 (N_19102,N_15012,N_15540);
nor U19103 (N_19103,N_15958,N_17122);
and U19104 (N_19104,N_16918,N_15590);
nand U19105 (N_19105,N_15991,N_15175);
nor U19106 (N_19106,N_16818,N_16708);
nand U19107 (N_19107,N_15579,N_15694);
nand U19108 (N_19108,N_15543,N_16850);
nand U19109 (N_19109,N_16873,N_15213);
or U19110 (N_19110,N_15291,N_16837);
nor U19111 (N_19111,N_16516,N_15403);
and U19112 (N_19112,N_17079,N_15856);
or U19113 (N_19113,N_15174,N_15588);
and U19114 (N_19114,N_15591,N_15117);
or U19115 (N_19115,N_15357,N_15402);
nor U19116 (N_19116,N_15332,N_15570);
nor U19117 (N_19117,N_15489,N_17099);
and U19118 (N_19118,N_15239,N_17397);
or U19119 (N_19119,N_15575,N_17154);
or U19120 (N_19120,N_16567,N_17477);
nor U19121 (N_19121,N_15680,N_16356);
nand U19122 (N_19122,N_15989,N_16272);
xnor U19123 (N_19123,N_16021,N_16659);
nor U19124 (N_19124,N_15893,N_16298);
nor U19125 (N_19125,N_15625,N_15811);
xor U19126 (N_19126,N_16688,N_16561);
nor U19127 (N_19127,N_16323,N_15412);
nor U19128 (N_19128,N_15276,N_15653);
nor U19129 (N_19129,N_16024,N_17367);
nand U19130 (N_19130,N_15696,N_16297);
nand U19131 (N_19131,N_15330,N_15603);
nand U19132 (N_19132,N_16631,N_16869);
or U19133 (N_19133,N_16171,N_16293);
xnor U19134 (N_19134,N_16749,N_15861);
or U19135 (N_19135,N_15620,N_16985);
nand U19136 (N_19136,N_15284,N_16817);
or U19137 (N_19137,N_15629,N_15327);
nor U19138 (N_19138,N_16134,N_15385);
nand U19139 (N_19139,N_16632,N_16232);
nor U19140 (N_19140,N_15687,N_15291);
or U19141 (N_19141,N_15377,N_16623);
or U19142 (N_19142,N_15416,N_16237);
nand U19143 (N_19143,N_17246,N_15267);
nand U19144 (N_19144,N_16254,N_15469);
xor U19145 (N_19145,N_16426,N_17407);
and U19146 (N_19146,N_17120,N_15267);
nor U19147 (N_19147,N_15740,N_16511);
nand U19148 (N_19148,N_15139,N_15462);
or U19149 (N_19149,N_15980,N_17154);
or U19150 (N_19150,N_16200,N_16752);
nor U19151 (N_19151,N_16108,N_16291);
nor U19152 (N_19152,N_16627,N_15236);
nor U19153 (N_19153,N_16181,N_15642);
nand U19154 (N_19154,N_15706,N_15103);
nor U19155 (N_19155,N_17166,N_16397);
nor U19156 (N_19156,N_17479,N_16894);
or U19157 (N_19157,N_16743,N_15037);
or U19158 (N_19158,N_15567,N_16121);
xnor U19159 (N_19159,N_16958,N_17325);
nand U19160 (N_19160,N_17248,N_15901);
nand U19161 (N_19161,N_16277,N_15847);
nor U19162 (N_19162,N_17047,N_17197);
and U19163 (N_19163,N_17269,N_16593);
and U19164 (N_19164,N_16063,N_15263);
nand U19165 (N_19165,N_17271,N_15422);
or U19166 (N_19166,N_17382,N_15443);
xor U19167 (N_19167,N_15792,N_15368);
nor U19168 (N_19168,N_15682,N_15647);
or U19169 (N_19169,N_16108,N_16393);
nor U19170 (N_19170,N_16530,N_15902);
xnor U19171 (N_19171,N_16801,N_17367);
nand U19172 (N_19172,N_15912,N_16101);
xnor U19173 (N_19173,N_15303,N_15065);
nor U19174 (N_19174,N_16067,N_15997);
xor U19175 (N_19175,N_17168,N_16823);
and U19176 (N_19176,N_16473,N_15420);
nand U19177 (N_19177,N_17078,N_15625);
nor U19178 (N_19178,N_17171,N_17162);
nand U19179 (N_19179,N_16998,N_15301);
or U19180 (N_19180,N_16475,N_16055);
or U19181 (N_19181,N_16153,N_15741);
or U19182 (N_19182,N_15576,N_16233);
xor U19183 (N_19183,N_15487,N_15373);
nand U19184 (N_19184,N_15266,N_15850);
nand U19185 (N_19185,N_15856,N_16891);
nor U19186 (N_19186,N_15192,N_15332);
or U19187 (N_19187,N_16482,N_15215);
or U19188 (N_19188,N_16396,N_17218);
nor U19189 (N_19189,N_15501,N_15622);
and U19190 (N_19190,N_17171,N_16930);
nor U19191 (N_19191,N_17409,N_17179);
or U19192 (N_19192,N_16459,N_16836);
nand U19193 (N_19193,N_17463,N_17457);
nor U19194 (N_19194,N_16115,N_17028);
and U19195 (N_19195,N_17372,N_16765);
and U19196 (N_19196,N_16450,N_15795);
xnor U19197 (N_19197,N_17027,N_17306);
or U19198 (N_19198,N_15158,N_15793);
nor U19199 (N_19199,N_16281,N_16581);
nor U19200 (N_19200,N_15885,N_16862);
nand U19201 (N_19201,N_16747,N_16777);
nand U19202 (N_19202,N_15427,N_16516);
nor U19203 (N_19203,N_16689,N_16043);
and U19204 (N_19204,N_16633,N_16298);
xnor U19205 (N_19205,N_17226,N_16018);
nand U19206 (N_19206,N_17416,N_16580);
or U19207 (N_19207,N_16735,N_17237);
nor U19208 (N_19208,N_15618,N_16239);
or U19209 (N_19209,N_16640,N_17488);
or U19210 (N_19210,N_16569,N_16228);
nor U19211 (N_19211,N_16616,N_16188);
nor U19212 (N_19212,N_17306,N_15704);
or U19213 (N_19213,N_15685,N_16882);
and U19214 (N_19214,N_15818,N_15285);
and U19215 (N_19215,N_16667,N_16695);
nor U19216 (N_19216,N_15597,N_15925);
nand U19217 (N_19217,N_16128,N_17471);
nor U19218 (N_19218,N_15675,N_16499);
nor U19219 (N_19219,N_17101,N_15473);
or U19220 (N_19220,N_15841,N_15495);
xor U19221 (N_19221,N_15733,N_16828);
or U19222 (N_19222,N_15791,N_15096);
or U19223 (N_19223,N_16497,N_15200);
xor U19224 (N_19224,N_16074,N_15350);
nor U19225 (N_19225,N_17372,N_15986);
nor U19226 (N_19226,N_15662,N_16633);
and U19227 (N_19227,N_15356,N_15867);
nand U19228 (N_19228,N_15204,N_15110);
xnor U19229 (N_19229,N_16250,N_16639);
and U19230 (N_19230,N_16371,N_15800);
or U19231 (N_19231,N_16486,N_17156);
nor U19232 (N_19232,N_17338,N_15452);
nand U19233 (N_19233,N_17095,N_17379);
xor U19234 (N_19234,N_17294,N_17124);
nor U19235 (N_19235,N_16465,N_16181);
and U19236 (N_19236,N_16968,N_17333);
and U19237 (N_19237,N_15426,N_16708);
and U19238 (N_19238,N_16697,N_16307);
nand U19239 (N_19239,N_15512,N_15752);
nand U19240 (N_19240,N_15218,N_15062);
xor U19241 (N_19241,N_16811,N_16391);
nand U19242 (N_19242,N_15266,N_17417);
and U19243 (N_19243,N_15603,N_15537);
and U19244 (N_19244,N_15972,N_15068);
and U19245 (N_19245,N_16860,N_15772);
and U19246 (N_19246,N_15301,N_15408);
or U19247 (N_19247,N_15195,N_15493);
nor U19248 (N_19248,N_16763,N_17422);
nand U19249 (N_19249,N_15459,N_15576);
nand U19250 (N_19250,N_15688,N_16166);
xor U19251 (N_19251,N_17367,N_15814);
and U19252 (N_19252,N_17194,N_17477);
and U19253 (N_19253,N_15745,N_16656);
and U19254 (N_19254,N_16381,N_15764);
or U19255 (N_19255,N_15889,N_15374);
nor U19256 (N_19256,N_15546,N_16621);
nor U19257 (N_19257,N_16507,N_15367);
nand U19258 (N_19258,N_16355,N_15383);
nor U19259 (N_19259,N_16225,N_17005);
or U19260 (N_19260,N_16108,N_16879);
or U19261 (N_19261,N_16779,N_16670);
and U19262 (N_19262,N_15874,N_15252);
nand U19263 (N_19263,N_16731,N_15587);
nand U19264 (N_19264,N_16345,N_17440);
and U19265 (N_19265,N_17372,N_17253);
and U19266 (N_19266,N_15609,N_17262);
or U19267 (N_19267,N_16532,N_17450);
nand U19268 (N_19268,N_16578,N_15832);
and U19269 (N_19269,N_15808,N_17431);
or U19270 (N_19270,N_15258,N_15158);
and U19271 (N_19271,N_15307,N_16691);
xnor U19272 (N_19272,N_16473,N_16831);
nor U19273 (N_19273,N_15248,N_15924);
xor U19274 (N_19274,N_17087,N_17007);
or U19275 (N_19275,N_17256,N_16636);
and U19276 (N_19276,N_16853,N_15411);
nand U19277 (N_19277,N_15811,N_16473);
xor U19278 (N_19278,N_15608,N_16838);
nor U19279 (N_19279,N_17412,N_16831);
nor U19280 (N_19280,N_16814,N_16525);
nor U19281 (N_19281,N_17494,N_16692);
xor U19282 (N_19282,N_17009,N_15628);
nor U19283 (N_19283,N_16166,N_16125);
or U19284 (N_19284,N_17401,N_17001);
or U19285 (N_19285,N_17248,N_17088);
xnor U19286 (N_19286,N_17115,N_17034);
or U19287 (N_19287,N_15832,N_15166);
and U19288 (N_19288,N_16406,N_15740);
or U19289 (N_19289,N_15859,N_15936);
xor U19290 (N_19290,N_16863,N_17205);
nor U19291 (N_19291,N_15112,N_16316);
or U19292 (N_19292,N_16066,N_16083);
and U19293 (N_19293,N_15246,N_17108);
nor U19294 (N_19294,N_16918,N_15765);
nand U19295 (N_19295,N_16040,N_16100);
and U19296 (N_19296,N_15704,N_16133);
or U19297 (N_19297,N_16890,N_17384);
nor U19298 (N_19298,N_17470,N_16547);
nand U19299 (N_19299,N_15158,N_15649);
nand U19300 (N_19300,N_15727,N_16286);
nor U19301 (N_19301,N_16986,N_16133);
and U19302 (N_19302,N_16144,N_15738);
and U19303 (N_19303,N_15805,N_17187);
nand U19304 (N_19304,N_15739,N_16307);
and U19305 (N_19305,N_16615,N_15913);
and U19306 (N_19306,N_15716,N_15469);
nand U19307 (N_19307,N_17107,N_17138);
and U19308 (N_19308,N_15950,N_15773);
nor U19309 (N_19309,N_17354,N_17152);
or U19310 (N_19310,N_16218,N_15277);
or U19311 (N_19311,N_16130,N_16372);
and U19312 (N_19312,N_16316,N_16766);
and U19313 (N_19313,N_15208,N_15540);
and U19314 (N_19314,N_15669,N_16074);
nor U19315 (N_19315,N_17499,N_17437);
and U19316 (N_19316,N_15072,N_17230);
nor U19317 (N_19317,N_16609,N_16002);
nor U19318 (N_19318,N_16974,N_15197);
nor U19319 (N_19319,N_16908,N_16905);
nor U19320 (N_19320,N_15994,N_17164);
nor U19321 (N_19321,N_16543,N_16736);
xor U19322 (N_19322,N_17287,N_17025);
nand U19323 (N_19323,N_16295,N_15231);
and U19324 (N_19324,N_17095,N_15203);
nand U19325 (N_19325,N_15625,N_16475);
nand U19326 (N_19326,N_15585,N_16551);
and U19327 (N_19327,N_15042,N_15018);
nor U19328 (N_19328,N_16599,N_15018);
or U19329 (N_19329,N_16830,N_16183);
and U19330 (N_19330,N_16903,N_17372);
and U19331 (N_19331,N_16090,N_15484);
or U19332 (N_19332,N_15492,N_16282);
nand U19333 (N_19333,N_17032,N_16070);
nor U19334 (N_19334,N_15167,N_16920);
and U19335 (N_19335,N_17291,N_15585);
nand U19336 (N_19336,N_17232,N_15769);
or U19337 (N_19337,N_15323,N_17341);
nor U19338 (N_19338,N_16693,N_16304);
or U19339 (N_19339,N_15481,N_16840);
or U19340 (N_19340,N_17176,N_16273);
and U19341 (N_19341,N_15132,N_16694);
or U19342 (N_19342,N_16854,N_15617);
and U19343 (N_19343,N_15706,N_16272);
and U19344 (N_19344,N_16431,N_15809);
nand U19345 (N_19345,N_16425,N_16476);
nor U19346 (N_19346,N_15638,N_17408);
xor U19347 (N_19347,N_16745,N_15232);
nor U19348 (N_19348,N_16686,N_15066);
nor U19349 (N_19349,N_15076,N_15580);
nand U19350 (N_19350,N_15487,N_16484);
or U19351 (N_19351,N_15814,N_16057);
and U19352 (N_19352,N_17122,N_17349);
nand U19353 (N_19353,N_17191,N_17235);
xor U19354 (N_19354,N_16281,N_15429);
nand U19355 (N_19355,N_15000,N_16492);
or U19356 (N_19356,N_15430,N_15104);
nand U19357 (N_19357,N_15390,N_16172);
nand U19358 (N_19358,N_15964,N_17036);
or U19359 (N_19359,N_16665,N_15190);
and U19360 (N_19360,N_17363,N_15130);
or U19361 (N_19361,N_15099,N_15575);
nor U19362 (N_19362,N_17435,N_15373);
nand U19363 (N_19363,N_16425,N_17326);
and U19364 (N_19364,N_16009,N_15751);
and U19365 (N_19365,N_15121,N_16156);
or U19366 (N_19366,N_15173,N_17212);
nor U19367 (N_19367,N_16271,N_17023);
nor U19368 (N_19368,N_16546,N_16901);
or U19369 (N_19369,N_16391,N_16727);
nor U19370 (N_19370,N_16202,N_16873);
or U19371 (N_19371,N_16529,N_17483);
and U19372 (N_19372,N_16418,N_15511);
and U19373 (N_19373,N_16691,N_17236);
and U19374 (N_19374,N_15650,N_16692);
nor U19375 (N_19375,N_17280,N_16038);
nand U19376 (N_19376,N_15317,N_15689);
nor U19377 (N_19377,N_16749,N_16090);
or U19378 (N_19378,N_16029,N_16474);
or U19379 (N_19379,N_15004,N_16772);
nand U19380 (N_19380,N_15489,N_15842);
nor U19381 (N_19381,N_16188,N_16271);
or U19382 (N_19382,N_15709,N_15114);
or U19383 (N_19383,N_15219,N_15762);
or U19384 (N_19384,N_17066,N_15892);
and U19385 (N_19385,N_15792,N_15021);
nor U19386 (N_19386,N_15674,N_16000);
or U19387 (N_19387,N_16414,N_15055);
nor U19388 (N_19388,N_17264,N_16608);
nor U19389 (N_19389,N_16243,N_16548);
and U19390 (N_19390,N_15025,N_16626);
xnor U19391 (N_19391,N_17104,N_16298);
and U19392 (N_19392,N_16679,N_16817);
nand U19393 (N_19393,N_17415,N_16668);
or U19394 (N_19394,N_15094,N_16818);
xnor U19395 (N_19395,N_17028,N_15659);
and U19396 (N_19396,N_15508,N_17010);
nor U19397 (N_19397,N_16676,N_15373);
and U19398 (N_19398,N_15738,N_15160);
nor U19399 (N_19399,N_16695,N_16895);
or U19400 (N_19400,N_15990,N_17101);
nand U19401 (N_19401,N_15647,N_15017);
xnor U19402 (N_19402,N_17159,N_17322);
nand U19403 (N_19403,N_15848,N_16135);
nor U19404 (N_19404,N_16461,N_15430);
nor U19405 (N_19405,N_17197,N_17066);
xor U19406 (N_19406,N_16913,N_17230);
xor U19407 (N_19407,N_16789,N_15764);
nand U19408 (N_19408,N_16247,N_16296);
xnor U19409 (N_19409,N_15875,N_16149);
and U19410 (N_19410,N_16244,N_15623);
and U19411 (N_19411,N_16245,N_16774);
nor U19412 (N_19412,N_15030,N_15611);
nor U19413 (N_19413,N_15576,N_15500);
or U19414 (N_19414,N_16447,N_15634);
nand U19415 (N_19415,N_15583,N_16359);
nor U19416 (N_19416,N_17007,N_17061);
nand U19417 (N_19417,N_16802,N_16706);
or U19418 (N_19418,N_15078,N_17392);
or U19419 (N_19419,N_17257,N_16323);
or U19420 (N_19420,N_15193,N_16305);
xnor U19421 (N_19421,N_16905,N_16873);
nor U19422 (N_19422,N_17142,N_16751);
or U19423 (N_19423,N_16254,N_17089);
or U19424 (N_19424,N_15575,N_16975);
nor U19425 (N_19425,N_15531,N_17024);
or U19426 (N_19426,N_16165,N_15186);
nand U19427 (N_19427,N_15141,N_17479);
and U19428 (N_19428,N_15798,N_16357);
nor U19429 (N_19429,N_16569,N_16919);
nand U19430 (N_19430,N_16863,N_15470);
or U19431 (N_19431,N_17300,N_16385);
nor U19432 (N_19432,N_15603,N_17290);
nand U19433 (N_19433,N_16212,N_16019);
or U19434 (N_19434,N_15954,N_17043);
and U19435 (N_19435,N_15387,N_15969);
nor U19436 (N_19436,N_15434,N_15777);
and U19437 (N_19437,N_17110,N_17007);
nand U19438 (N_19438,N_17234,N_17367);
and U19439 (N_19439,N_15579,N_17179);
nor U19440 (N_19440,N_16222,N_16893);
and U19441 (N_19441,N_15129,N_15685);
xor U19442 (N_19442,N_16311,N_15010);
nor U19443 (N_19443,N_17480,N_16179);
and U19444 (N_19444,N_16996,N_16252);
or U19445 (N_19445,N_16098,N_15106);
and U19446 (N_19446,N_15173,N_15778);
nand U19447 (N_19447,N_17468,N_15259);
and U19448 (N_19448,N_15160,N_16384);
and U19449 (N_19449,N_16923,N_16303);
nor U19450 (N_19450,N_17055,N_16639);
nor U19451 (N_19451,N_15231,N_15483);
xnor U19452 (N_19452,N_15175,N_15184);
and U19453 (N_19453,N_15786,N_17353);
nand U19454 (N_19454,N_15839,N_16463);
and U19455 (N_19455,N_16487,N_15740);
and U19456 (N_19456,N_16630,N_17445);
xnor U19457 (N_19457,N_15507,N_16716);
nor U19458 (N_19458,N_17118,N_16726);
nor U19459 (N_19459,N_16338,N_17433);
nand U19460 (N_19460,N_16698,N_16451);
nand U19461 (N_19461,N_16243,N_17459);
nor U19462 (N_19462,N_16638,N_17010);
xnor U19463 (N_19463,N_17423,N_15331);
and U19464 (N_19464,N_17208,N_16174);
and U19465 (N_19465,N_15848,N_15461);
nor U19466 (N_19466,N_16855,N_16501);
or U19467 (N_19467,N_15849,N_16448);
nor U19468 (N_19468,N_15275,N_16313);
nor U19469 (N_19469,N_17127,N_16134);
or U19470 (N_19470,N_15402,N_17016);
and U19471 (N_19471,N_16595,N_15289);
and U19472 (N_19472,N_16299,N_15342);
nand U19473 (N_19473,N_15978,N_16941);
or U19474 (N_19474,N_15038,N_16497);
nand U19475 (N_19475,N_15618,N_15057);
nor U19476 (N_19476,N_15590,N_16920);
nor U19477 (N_19477,N_17308,N_15749);
and U19478 (N_19478,N_16509,N_16044);
nand U19479 (N_19479,N_17136,N_15737);
nand U19480 (N_19480,N_15090,N_16124);
nand U19481 (N_19481,N_16542,N_16482);
nand U19482 (N_19482,N_16088,N_17026);
or U19483 (N_19483,N_15452,N_15938);
nor U19484 (N_19484,N_15783,N_16497);
nand U19485 (N_19485,N_15738,N_16602);
xor U19486 (N_19486,N_15963,N_16748);
or U19487 (N_19487,N_16786,N_16005);
nand U19488 (N_19488,N_16795,N_15218);
or U19489 (N_19489,N_16503,N_15400);
xor U19490 (N_19490,N_16075,N_16622);
nor U19491 (N_19491,N_15881,N_16656);
nor U19492 (N_19492,N_16165,N_15998);
nor U19493 (N_19493,N_15863,N_16970);
and U19494 (N_19494,N_15040,N_16011);
nand U19495 (N_19495,N_15528,N_15074);
and U19496 (N_19496,N_15900,N_17362);
nor U19497 (N_19497,N_15957,N_17210);
nor U19498 (N_19498,N_16900,N_17419);
nand U19499 (N_19499,N_16460,N_17143);
or U19500 (N_19500,N_15892,N_16644);
nor U19501 (N_19501,N_15763,N_16905);
nand U19502 (N_19502,N_16526,N_16407);
and U19503 (N_19503,N_15800,N_17389);
nor U19504 (N_19504,N_16659,N_17290);
xnor U19505 (N_19505,N_17050,N_16959);
or U19506 (N_19506,N_17345,N_16932);
nand U19507 (N_19507,N_15805,N_17141);
nor U19508 (N_19508,N_16071,N_15717);
xor U19509 (N_19509,N_15252,N_15288);
or U19510 (N_19510,N_16011,N_15353);
xor U19511 (N_19511,N_15024,N_16607);
nand U19512 (N_19512,N_15636,N_16052);
and U19513 (N_19513,N_16830,N_15309);
or U19514 (N_19514,N_16001,N_15189);
and U19515 (N_19515,N_16573,N_17245);
nand U19516 (N_19516,N_16221,N_16213);
or U19517 (N_19517,N_16300,N_16180);
nor U19518 (N_19518,N_16284,N_16226);
nand U19519 (N_19519,N_15058,N_16002);
nor U19520 (N_19520,N_16986,N_16345);
nor U19521 (N_19521,N_16756,N_15961);
or U19522 (N_19522,N_16337,N_16963);
xnor U19523 (N_19523,N_15752,N_16173);
or U19524 (N_19524,N_17025,N_16967);
nor U19525 (N_19525,N_16162,N_16494);
or U19526 (N_19526,N_16743,N_16784);
or U19527 (N_19527,N_15487,N_15620);
nand U19528 (N_19528,N_15419,N_17427);
or U19529 (N_19529,N_16872,N_16983);
nor U19530 (N_19530,N_15026,N_15774);
and U19531 (N_19531,N_15564,N_15447);
or U19532 (N_19532,N_16018,N_17427);
nand U19533 (N_19533,N_17042,N_15208);
nor U19534 (N_19534,N_16430,N_16378);
nand U19535 (N_19535,N_16828,N_16435);
or U19536 (N_19536,N_16187,N_16177);
nand U19537 (N_19537,N_17349,N_17089);
or U19538 (N_19538,N_15565,N_16351);
and U19539 (N_19539,N_16061,N_16004);
and U19540 (N_19540,N_15813,N_15852);
nand U19541 (N_19541,N_15057,N_16545);
nor U19542 (N_19542,N_15887,N_16985);
and U19543 (N_19543,N_15660,N_16429);
and U19544 (N_19544,N_17447,N_17026);
or U19545 (N_19545,N_16913,N_16383);
nand U19546 (N_19546,N_15964,N_15537);
or U19547 (N_19547,N_15411,N_17286);
or U19548 (N_19548,N_15122,N_16651);
and U19549 (N_19549,N_15043,N_15398);
nor U19550 (N_19550,N_17303,N_15897);
xor U19551 (N_19551,N_16895,N_15687);
or U19552 (N_19552,N_16987,N_16401);
nand U19553 (N_19553,N_15310,N_16128);
nor U19554 (N_19554,N_16842,N_16815);
and U19555 (N_19555,N_15287,N_15241);
nand U19556 (N_19556,N_16977,N_16127);
or U19557 (N_19557,N_16213,N_16607);
nand U19558 (N_19558,N_16278,N_15149);
nand U19559 (N_19559,N_15023,N_15592);
or U19560 (N_19560,N_15117,N_17381);
nor U19561 (N_19561,N_16259,N_16920);
nor U19562 (N_19562,N_16467,N_15028);
nor U19563 (N_19563,N_17451,N_15131);
nand U19564 (N_19564,N_15637,N_16488);
nor U19565 (N_19565,N_15002,N_15398);
and U19566 (N_19566,N_15706,N_15571);
or U19567 (N_19567,N_15014,N_16270);
nand U19568 (N_19568,N_16998,N_15837);
nand U19569 (N_19569,N_15939,N_15230);
and U19570 (N_19570,N_15052,N_15766);
xor U19571 (N_19571,N_16791,N_15285);
nand U19572 (N_19572,N_16501,N_15852);
nand U19573 (N_19573,N_17259,N_17491);
and U19574 (N_19574,N_17438,N_15009);
nand U19575 (N_19575,N_15984,N_16177);
and U19576 (N_19576,N_16227,N_16560);
nor U19577 (N_19577,N_15216,N_15994);
xnor U19578 (N_19578,N_15518,N_15279);
and U19579 (N_19579,N_16364,N_16449);
or U19580 (N_19580,N_15274,N_15042);
or U19581 (N_19581,N_15407,N_15570);
nand U19582 (N_19582,N_15819,N_16532);
nor U19583 (N_19583,N_16360,N_16961);
or U19584 (N_19584,N_16679,N_16872);
nand U19585 (N_19585,N_16654,N_15266);
nor U19586 (N_19586,N_17190,N_16126);
and U19587 (N_19587,N_16044,N_16373);
nand U19588 (N_19588,N_16484,N_15917);
xnor U19589 (N_19589,N_17041,N_15754);
nor U19590 (N_19590,N_15475,N_15439);
nand U19591 (N_19591,N_15024,N_17277);
and U19592 (N_19592,N_17340,N_16941);
or U19593 (N_19593,N_16303,N_17123);
xnor U19594 (N_19594,N_16216,N_16493);
and U19595 (N_19595,N_15508,N_15931);
or U19596 (N_19596,N_16025,N_15379);
nand U19597 (N_19597,N_17030,N_17142);
or U19598 (N_19598,N_15069,N_15991);
nor U19599 (N_19599,N_17464,N_16390);
and U19600 (N_19600,N_15108,N_17452);
nand U19601 (N_19601,N_16812,N_16517);
and U19602 (N_19602,N_15865,N_16698);
xor U19603 (N_19603,N_15470,N_15462);
nor U19604 (N_19604,N_16759,N_15185);
or U19605 (N_19605,N_15061,N_16479);
nor U19606 (N_19606,N_15343,N_15734);
nor U19607 (N_19607,N_15741,N_15944);
nand U19608 (N_19608,N_16714,N_15354);
or U19609 (N_19609,N_17098,N_15653);
or U19610 (N_19610,N_16566,N_15733);
nand U19611 (N_19611,N_16903,N_17275);
nand U19612 (N_19612,N_16955,N_17090);
or U19613 (N_19613,N_16967,N_17386);
nand U19614 (N_19614,N_17400,N_17012);
nor U19615 (N_19615,N_16423,N_17206);
nor U19616 (N_19616,N_16798,N_16676);
and U19617 (N_19617,N_17271,N_15864);
and U19618 (N_19618,N_17319,N_15964);
and U19619 (N_19619,N_16744,N_15667);
or U19620 (N_19620,N_15454,N_15510);
xor U19621 (N_19621,N_17223,N_16672);
nand U19622 (N_19622,N_15584,N_17072);
and U19623 (N_19623,N_17466,N_15709);
and U19624 (N_19624,N_16625,N_16081);
nor U19625 (N_19625,N_15712,N_16925);
and U19626 (N_19626,N_15341,N_15116);
nor U19627 (N_19627,N_16809,N_15530);
and U19628 (N_19628,N_15670,N_16146);
nor U19629 (N_19629,N_15136,N_15576);
nor U19630 (N_19630,N_16826,N_16332);
nand U19631 (N_19631,N_16315,N_16969);
xnor U19632 (N_19632,N_15435,N_16195);
nor U19633 (N_19633,N_16331,N_15298);
nor U19634 (N_19634,N_16051,N_16653);
and U19635 (N_19635,N_15957,N_15682);
nor U19636 (N_19636,N_15113,N_15639);
or U19637 (N_19637,N_15966,N_17201);
nor U19638 (N_19638,N_16807,N_15719);
nor U19639 (N_19639,N_16826,N_16034);
nand U19640 (N_19640,N_15815,N_16036);
nor U19641 (N_19641,N_17306,N_15772);
and U19642 (N_19642,N_15339,N_17040);
nor U19643 (N_19643,N_16647,N_16261);
nand U19644 (N_19644,N_16433,N_16033);
and U19645 (N_19645,N_15113,N_16815);
or U19646 (N_19646,N_15524,N_16612);
or U19647 (N_19647,N_17030,N_15993);
or U19648 (N_19648,N_17244,N_16786);
and U19649 (N_19649,N_16957,N_15265);
and U19650 (N_19650,N_17007,N_16855);
nand U19651 (N_19651,N_15021,N_17177);
or U19652 (N_19652,N_15043,N_16966);
and U19653 (N_19653,N_15943,N_17350);
or U19654 (N_19654,N_15159,N_17064);
nor U19655 (N_19655,N_16468,N_16630);
or U19656 (N_19656,N_15228,N_16359);
or U19657 (N_19657,N_15977,N_16918);
or U19658 (N_19658,N_16523,N_16719);
and U19659 (N_19659,N_15455,N_17144);
nor U19660 (N_19660,N_16202,N_17062);
xnor U19661 (N_19661,N_17322,N_16294);
nand U19662 (N_19662,N_17477,N_15202);
nor U19663 (N_19663,N_16101,N_15043);
and U19664 (N_19664,N_15522,N_15255);
or U19665 (N_19665,N_15340,N_17284);
or U19666 (N_19666,N_15170,N_16666);
nand U19667 (N_19667,N_16484,N_15561);
nand U19668 (N_19668,N_16366,N_16300);
or U19669 (N_19669,N_15098,N_15598);
or U19670 (N_19670,N_15447,N_17352);
and U19671 (N_19671,N_17165,N_16070);
or U19672 (N_19672,N_16622,N_17339);
or U19673 (N_19673,N_15764,N_15206);
and U19674 (N_19674,N_17341,N_16237);
nor U19675 (N_19675,N_15863,N_15673);
nand U19676 (N_19676,N_15742,N_15703);
nand U19677 (N_19677,N_15801,N_15187);
nor U19678 (N_19678,N_16445,N_16917);
and U19679 (N_19679,N_17125,N_15587);
and U19680 (N_19680,N_17090,N_16633);
nor U19681 (N_19681,N_17387,N_16308);
nand U19682 (N_19682,N_16450,N_16531);
xnor U19683 (N_19683,N_15773,N_15712);
nor U19684 (N_19684,N_17133,N_17116);
nand U19685 (N_19685,N_15694,N_16240);
and U19686 (N_19686,N_15984,N_17115);
and U19687 (N_19687,N_16916,N_15356);
or U19688 (N_19688,N_17053,N_15020);
or U19689 (N_19689,N_15702,N_16382);
nand U19690 (N_19690,N_16109,N_15009);
or U19691 (N_19691,N_15748,N_17483);
xnor U19692 (N_19692,N_16629,N_15525);
xor U19693 (N_19693,N_15428,N_16553);
and U19694 (N_19694,N_16376,N_15122);
or U19695 (N_19695,N_16006,N_16189);
nand U19696 (N_19696,N_17063,N_16600);
nand U19697 (N_19697,N_17278,N_15537);
nor U19698 (N_19698,N_15396,N_15833);
xnor U19699 (N_19699,N_16065,N_15827);
and U19700 (N_19700,N_15072,N_15774);
and U19701 (N_19701,N_16818,N_15548);
and U19702 (N_19702,N_16783,N_16443);
or U19703 (N_19703,N_17401,N_17465);
and U19704 (N_19704,N_17038,N_15194);
and U19705 (N_19705,N_15257,N_16082);
nor U19706 (N_19706,N_16679,N_15050);
nand U19707 (N_19707,N_17249,N_15439);
nor U19708 (N_19708,N_17455,N_16560);
and U19709 (N_19709,N_17275,N_17144);
nor U19710 (N_19710,N_15928,N_16102);
or U19711 (N_19711,N_16767,N_16333);
nand U19712 (N_19712,N_17049,N_15979);
nand U19713 (N_19713,N_16333,N_17469);
nor U19714 (N_19714,N_16703,N_16003);
or U19715 (N_19715,N_16131,N_16726);
and U19716 (N_19716,N_15376,N_15057);
or U19717 (N_19717,N_15028,N_17469);
xor U19718 (N_19718,N_16824,N_15328);
nor U19719 (N_19719,N_17308,N_15164);
nor U19720 (N_19720,N_15578,N_16203);
xnor U19721 (N_19721,N_16252,N_15501);
nor U19722 (N_19722,N_16319,N_15291);
nor U19723 (N_19723,N_15676,N_16908);
and U19724 (N_19724,N_17463,N_17462);
or U19725 (N_19725,N_15770,N_15999);
nor U19726 (N_19726,N_15714,N_15343);
xnor U19727 (N_19727,N_17187,N_16362);
or U19728 (N_19728,N_17037,N_16107);
nand U19729 (N_19729,N_16968,N_16601);
or U19730 (N_19730,N_16972,N_16218);
nor U19731 (N_19731,N_15033,N_15852);
and U19732 (N_19732,N_17280,N_16419);
or U19733 (N_19733,N_15510,N_15526);
nor U19734 (N_19734,N_15979,N_16172);
nand U19735 (N_19735,N_16112,N_16246);
or U19736 (N_19736,N_15677,N_15713);
and U19737 (N_19737,N_16453,N_16691);
or U19738 (N_19738,N_16300,N_15575);
nand U19739 (N_19739,N_15275,N_15130);
and U19740 (N_19740,N_17059,N_17443);
nor U19741 (N_19741,N_17322,N_16540);
and U19742 (N_19742,N_15678,N_15376);
xnor U19743 (N_19743,N_16281,N_16499);
or U19744 (N_19744,N_16920,N_17027);
or U19745 (N_19745,N_16066,N_15574);
and U19746 (N_19746,N_16217,N_16370);
or U19747 (N_19747,N_16837,N_15775);
and U19748 (N_19748,N_15255,N_15760);
and U19749 (N_19749,N_16461,N_16987);
nor U19750 (N_19750,N_16572,N_16655);
nand U19751 (N_19751,N_15787,N_15595);
nand U19752 (N_19752,N_16522,N_16181);
and U19753 (N_19753,N_15422,N_17204);
or U19754 (N_19754,N_16821,N_15354);
and U19755 (N_19755,N_15518,N_16319);
or U19756 (N_19756,N_15571,N_15119);
xnor U19757 (N_19757,N_16745,N_16068);
nor U19758 (N_19758,N_15381,N_15452);
and U19759 (N_19759,N_17472,N_16303);
nand U19760 (N_19760,N_15984,N_16106);
nand U19761 (N_19761,N_15730,N_16801);
and U19762 (N_19762,N_15951,N_16394);
and U19763 (N_19763,N_17203,N_17210);
and U19764 (N_19764,N_15316,N_16384);
or U19765 (N_19765,N_15749,N_15096);
and U19766 (N_19766,N_17045,N_17362);
or U19767 (N_19767,N_16128,N_15967);
and U19768 (N_19768,N_16141,N_15360);
or U19769 (N_19769,N_17191,N_15988);
nor U19770 (N_19770,N_17010,N_16224);
and U19771 (N_19771,N_15100,N_17157);
and U19772 (N_19772,N_16954,N_16868);
and U19773 (N_19773,N_15627,N_15461);
nor U19774 (N_19774,N_16149,N_15769);
nor U19775 (N_19775,N_17321,N_17332);
and U19776 (N_19776,N_15875,N_16866);
or U19777 (N_19777,N_15440,N_16820);
or U19778 (N_19778,N_15346,N_15667);
nor U19779 (N_19779,N_16618,N_15656);
nor U19780 (N_19780,N_16305,N_15608);
nor U19781 (N_19781,N_16731,N_16284);
xor U19782 (N_19782,N_15350,N_16550);
xor U19783 (N_19783,N_16675,N_17248);
and U19784 (N_19784,N_16515,N_16148);
or U19785 (N_19785,N_15162,N_17205);
nand U19786 (N_19786,N_15526,N_17200);
or U19787 (N_19787,N_17445,N_15864);
xor U19788 (N_19788,N_15568,N_16390);
nand U19789 (N_19789,N_17060,N_17072);
or U19790 (N_19790,N_15775,N_17408);
or U19791 (N_19791,N_17357,N_16635);
xnor U19792 (N_19792,N_15563,N_17129);
and U19793 (N_19793,N_15401,N_17339);
nor U19794 (N_19794,N_16222,N_16825);
xnor U19795 (N_19795,N_15397,N_17321);
xnor U19796 (N_19796,N_15657,N_15986);
nand U19797 (N_19797,N_15641,N_16269);
or U19798 (N_19798,N_15918,N_15004);
nor U19799 (N_19799,N_15312,N_16782);
nand U19800 (N_19800,N_17110,N_15525);
nor U19801 (N_19801,N_15375,N_16311);
or U19802 (N_19802,N_16809,N_16796);
or U19803 (N_19803,N_15287,N_16771);
or U19804 (N_19804,N_15345,N_16817);
or U19805 (N_19805,N_15525,N_16366);
nand U19806 (N_19806,N_16997,N_17462);
nand U19807 (N_19807,N_15742,N_17459);
nor U19808 (N_19808,N_15010,N_16768);
nand U19809 (N_19809,N_15359,N_17119);
nand U19810 (N_19810,N_16862,N_15759);
nand U19811 (N_19811,N_17276,N_16927);
and U19812 (N_19812,N_15508,N_15410);
nor U19813 (N_19813,N_16142,N_16780);
and U19814 (N_19814,N_17483,N_15563);
nor U19815 (N_19815,N_16833,N_16485);
or U19816 (N_19816,N_16613,N_15897);
and U19817 (N_19817,N_17458,N_16802);
and U19818 (N_19818,N_17219,N_15966);
nand U19819 (N_19819,N_17367,N_16243);
or U19820 (N_19820,N_16525,N_16870);
or U19821 (N_19821,N_16196,N_16611);
xnor U19822 (N_19822,N_16378,N_15188);
and U19823 (N_19823,N_15224,N_15290);
or U19824 (N_19824,N_15953,N_15767);
xor U19825 (N_19825,N_15933,N_17187);
nor U19826 (N_19826,N_15392,N_17148);
xor U19827 (N_19827,N_16918,N_16307);
nand U19828 (N_19828,N_17026,N_15884);
and U19829 (N_19829,N_15514,N_15825);
and U19830 (N_19830,N_16912,N_15436);
nand U19831 (N_19831,N_17337,N_15814);
nor U19832 (N_19832,N_15821,N_16149);
nor U19833 (N_19833,N_17276,N_16868);
nor U19834 (N_19834,N_15683,N_17226);
nor U19835 (N_19835,N_15532,N_17385);
xor U19836 (N_19836,N_16043,N_16089);
nand U19837 (N_19837,N_16419,N_15171);
xnor U19838 (N_19838,N_16860,N_15391);
and U19839 (N_19839,N_15884,N_16410);
or U19840 (N_19840,N_16024,N_16117);
nand U19841 (N_19841,N_15146,N_16942);
nand U19842 (N_19842,N_16490,N_16738);
or U19843 (N_19843,N_15335,N_15151);
nor U19844 (N_19844,N_15458,N_17239);
nor U19845 (N_19845,N_15333,N_16715);
nor U19846 (N_19846,N_16029,N_15618);
nor U19847 (N_19847,N_17014,N_15180);
and U19848 (N_19848,N_17374,N_17143);
and U19849 (N_19849,N_15752,N_15313);
or U19850 (N_19850,N_17254,N_16845);
nor U19851 (N_19851,N_17482,N_17179);
nand U19852 (N_19852,N_16276,N_16010);
xor U19853 (N_19853,N_16401,N_16339);
or U19854 (N_19854,N_16112,N_15029);
nand U19855 (N_19855,N_16938,N_15210);
nor U19856 (N_19856,N_16521,N_16881);
or U19857 (N_19857,N_15883,N_16094);
nand U19858 (N_19858,N_15222,N_16349);
and U19859 (N_19859,N_16642,N_17185);
nor U19860 (N_19860,N_15585,N_16034);
nor U19861 (N_19861,N_16385,N_15479);
or U19862 (N_19862,N_15132,N_17333);
and U19863 (N_19863,N_16729,N_15264);
nand U19864 (N_19864,N_15582,N_15185);
and U19865 (N_19865,N_15027,N_15616);
nand U19866 (N_19866,N_16096,N_15443);
and U19867 (N_19867,N_15488,N_15386);
nand U19868 (N_19868,N_17380,N_15848);
nand U19869 (N_19869,N_17410,N_16738);
and U19870 (N_19870,N_15229,N_15155);
nor U19871 (N_19871,N_15708,N_17032);
or U19872 (N_19872,N_15371,N_15363);
or U19873 (N_19873,N_15113,N_15273);
xnor U19874 (N_19874,N_17296,N_16372);
nand U19875 (N_19875,N_16727,N_17141);
nand U19876 (N_19876,N_16374,N_15583);
xnor U19877 (N_19877,N_17376,N_15622);
nand U19878 (N_19878,N_15854,N_17174);
and U19879 (N_19879,N_15746,N_15533);
nor U19880 (N_19880,N_16792,N_15721);
xor U19881 (N_19881,N_17228,N_15108);
and U19882 (N_19882,N_15175,N_15694);
or U19883 (N_19883,N_15351,N_15760);
or U19884 (N_19884,N_17221,N_15175);
nor U19885 (N_19885,N_16287,N_15913);
nor U19886 (N_19886,N_15872,N_15929);
nor U19887 (N_19887,N_16121,N_15424);
nor U19888 (N_19888,N_15400,N_16128);
and U19889 (N_19889,N_17156,N_17132);
or U19890 (N_19890,N_16918,N_16997);
or U19891 (N_19891,N_16261,N_17100);
nand U19892 (N_19892,N_15882,N_15435);
and U19893 (N_19893,N_16625,N_16836);
nor U19894 (N_19894,N_17180,N_15857);
or U19895 (N_19895,N_17020,N_15331);
or U19896 (N_19896,N_17143,N_16079);
or U19897 (N_19897,N_15158,N_15153);
nand U19898 (N_19898,N_16241,N_16469);
nand U19899 (N_19899,N_15155,N_16883);
and U19900 (N_19900,N_17242,N_16177);
and U19901 (N_19901,N_15453,N_16516);
and U19902 (N_19902,N_15300,N_16804);
and U19903 (N_19903,N_17409,N_17369);
nor U19904 (N_19904,N_15594,N_15797);
xor U19905 (N_19905,N_16359,N_15938);
or U19906 (N_19906,N_17321,N_16520);
and U19907 (N_19907,N_15452,N_17490);
nand U19908 (N_19908,N_17393,N_17413);
or U19909 (N_19909,N_16846,N_17381);
or U19910 (N_19910,N_17060,N_16516);
nand U19911 (N_19911,N_15522,N_16124);
xnor U19912 (N_19912,N_15559,N_15233);
nand U19913 (N_19913,N_15619,N_15935);
and U19914 (N_19914,N_15248,N_15440);
or U19915 (N_19915,N_17280,N_17100);
nand U19916 (N_19916,N_16245,N_15378);
nand U19917 (N_19917,N_16821,N_17070);
and U19918 (N_19918,N_16531,N_17140);
nor U19919 (N_19919,N_16655,N_16353);
nand U19920 (N_19920,N_15544,N_17018);
or U19921 (N_19921,N_17013,N_17110);
and U19922 (N_19922,N_16855,N_17408);
xnor U19923 (N_19923,N_17462,N_16240);
and U19924 (N_19924,N_17256,N_17270);
and U19925 (N_19925,N_15908,N_15872);
or U19926 (N_19926,N_16769,N_15797);
nor U19927 (N_19927,N_16901,N_15652);
nor U19928 (N_19928,N_16197,N_16958);
or U19929 (N_19929,N_15321,N_16695);
nor U19930 (N_19930,N_15209,N_15875);
xor U19931 (N_19931,N_15655,N_16630);
or U19932 (N_19932,N_17009,N_16022);
nor U19933 (N_19933,N_15269,N_15463);
nor U19934 (N_19934,N_16498,N_15545);
xnor U19935 (N_19935,N_15266,N_15134);
nand U19936 (N_19936,N_16695,N_17179);
xor U19937 (N_19937,N_16729,N_15676);
nor U19938 (N_19938,N_16654,N_16687);
nor U19939 (N_19939,N_16605,N_15197);
and U19940 (N_19940,N_16930,N_17117);
and U19941 (N_19941,N_16301,N_16150);
xor U19942 (N_19942,N_16737,N_17229);
or U19943 (N_19943,N_15342,N_17062);
and U19944 (N_19944,N_16669,N_15503);
nand U19945 (N_19945,N_15080,N_17227);
nor U19946 (N_19946,N_15735,N_16323);
xnor U19947 (N_19947,N_15625,N_15369);
and U19948 (N_19948,N_16047,N_16556);
and U19949 (N_19949,N_16090,N_15666);
and U19950 (N_19950,N_16248,N_15001);
nor U19951 (N_19951,N_17055,N_16636);
nand U19952 (N_19952,N_16075,N_16477);
nor U19953 (N_19953,N_17431,N_15237);
nor U19954 (N_19954,N_17386,N_15594);
and U19955 (N_19955,N_15654,N_15969);
and U19956 (N_19956,N_15689,N_16947);
and U19957 (N_19957,N_15955,N_16044);
or U19958 (N_19958,N_15344,N_15738);
nor U19959 (N_19959,N_16722,N_16397);
nand U19960 (N_19960,N_16299,N_16311);
nand U19961 (N_19961,N_15439,N_16931);
or U19962 (N_19962,N_17433,N_16821);
and U19963 (N_19963,N_15811,N_15226);
nor U19964 (N_19964,N_15468,N_17488);
or U19965 (N_19965,N_15772,N_15329);
and U19966 (N_19966,N_16104,N_15950);
or U19967 (N_19967,N_16940,N_17255);
and U19968 (N_19968,N_15654,N_17396);
xor U19969 (N_19969,N_15915,N_16432);
or U19970 (N_19970,N_16028,N_16080);
nor U19971 (N_19971,N_17467,N_16093);
or U19972 (N_19972,N_16486,N_17415);
xor U19973 (N_19973,N_16209,N_15595);
or U19974 (N_19974,N_17460,N_17462);
and U19975 (N_19975,N_15816,N_15702);
nor U19976 (N_19976,N_15539,N_16252);
nand U19977 (N_19977,N_16373,N_16631);
and U19978 (N_19978,N_16849,N_15491);
and U19979 (N_19979,N_15226,N_17110);
xnor U19980 (N_19980,N_16601,N_16162);
nor U19981 (N_19981,N_15001,N_15200);
xnor U19982 (N_19982,N_16640,N_17073);
nand U19983 (N_19983,N_17310,N_15412);
and U19984 (N_19984,N_16724,N_15100);
nand U19985 (N_19985,N_15099,N_17134);
nor U19986 (N_19986,N_17229,N_16487);
nand U19987 (N_19987,N_15631,N_15083);
nor U19988 (N_19988,N_15289,N_16524);
nor U19989 (N_19989,N_16048,N_15850);
nand U19990 (N_19990,N_16840,N_15464);
or U19991 (N_19991,N_16584,N_15111);
or U19992 (N_19992,N_15840,N_16224);
and U19993 (N_19993,N_15434,N_17492);
and U19994 (N_19994,N_17265,N_16292);
xnor U19995 (N_19995,N_17131,N_16575);
nor U19996 (N_19996,N_16401,N_16179);
or U19997 (N_19997,N_16970,N_15793);
nor U19998 (N_19998,N_15359,N_15674);
nand U19999 (N_19999,N_15634,N_15887);
and U20000 (N_20000,N_19119,N_18160);
and U20001 (N_20001,N_17569,N_18120);
or U20002 (N_20002,N_19724,N_19994);
and U20003 (N_20003,N_17516,N_18674);
nor U20004 (N_20004,N_18127,N_18647);
or U20005 (N_20005,N_17951,N_18267);
and U20006 (N_20006,N_19149,N_18624);
and U20007 (N_20007,N_17792,N_17953);
nor U20008 (N_20008,N_19627,N_18035);
nand U20009 (N_20009,N_18212,N_18795);
or U20010 (N_20010,N_19676,N_17727);
nor U20011 (N_20011,N_17614,N_19088);
nand U20012 (N_20012,N_18649,N_18416);
nor U20013 (N_20013,N_19282,N_18184);
and U20014 (N_20014,N_18867,N_19963);
nand U20015 (N_20015,N_18700,N_19787);
nand U20016 (N_20016,N_18147,N_18710);
or U20017 (N_20017,N_19421,N_17777);
or U20018 (N_20018,N_19722,N_19038);
or U20019 (N_20019,N_18937,N_19021);
and U20020 (N_20020,N_19017,N_18140);
or U20021 (N_20021,N_17844,N_18450);
and U20022 (N_20022,N_17623,N_18480);
and U20023 (N_20023,N_18492,N_19848);
nor U20024 (N_20024,N_17832,N_18695);
nor U20025 (N_20025,N_17500,N_19650);
and U20026 (N_20026,N_18681,N_18005);
nand U20027 (N_20027,N_18353,N_18866);
nor U20028 (N_20028,N_19438,N_19753);
nand U20029 (N_20029,N_18792,N_18716);
nand U20030 (N_20030,N_18722,N_19492);
or U20031 (N_20031,N_19815,N_17537);
xnor U20032 (N_20032,N_19698,N_18659);
xor U20033 (N_20033,N_17738,N_19425);
nor U20034 (N_20034,N_18664,N_19805);
or U20035 (N_20035,N_18001,N_17863);
nor U20036 (N_20036,N_19285,N_19075);
nand U20037 (N_20037,N_18266,N_19110);
xor U20038 (N_20038,N_17881,N_19095);
nor U20039 (N_20039,N_18972,N_18224);
nor U20040 (N_20040,N_19906,N_19467);
and U20041 (N_20041,N_17575,N_18757);
nand U20042 (N_20042,N_17534,N_18247);
or U20043 (N_20043,N_19346,N_17707);
nor U20044 (N_20044,N_18306,N_17725);
nor U20045 (N_20045,N_19476,N_18406);
xor U20046 (N_20046,N_18167,N_19998);
and U20047 (N_20047,N_18110,N_17719);
or U20048 (N_20048,N_18836,N_18408);
and U20049 (N_20049,N_17542,N_18448);
nor U20050 (N_20050,N_17960,N_19794);
and U20051 (N_20051,N_17914,N_18694);
nand U20052 (N_20052,N_17886,N_19071);
or U20053 (N_20053,N_18025,N_18967);
and U20054 (N_20054,N_18427,N_18029);
and U20055 (N_20055,N_19435,N_18227);
nor U20056 (N_20056,N_19025,N_18785);
or U20057 (N_20057,N_18244,N_17654);
xnor U20058 (N_20058,N_18115,N_18968);
and U20059 (N_20059,N_19675,N_19197);
xor U20060 (N_20060,N_19209,N_18639);
or U20061 (N_20061,N_17539,N_18597);
nor U20062 (N_20062,N_18661,N_17599);
or U20063 (N_20063,N_19696,N_18194);
or U20064 (N_20064,N_19242,N_17814);
nor U20065 (N_20065,N_17984,N_19937);
and U20066 (N_20066,N_19631,N_17928);
nor U20067 (N_20067,N_19389,N_19861);
or U20068 (N_20068,N_19816,N_18189);
and U20069 (N_20069,N_18572,N_17919);
or U20070 (N_20070,N_17970,N_19645);
nor U20071 (N_20071,N_18027,N_18500);
and U20072 (N_20072,N_17821,N_19252);
nor U20073 (N_20073,N_19576,N_19341);
or U20074 (N_20074,N_19719,N_19977);
nand U20075 (N_20075,N_18780,N_18458);
or U20076 (N_20076,N_17664,N_18508);
xnor U20077 (N_20077,N_17962,N_18553);
xor U20078 (N_20078,N_18913,N_18513);
nand U20079 (N_20079,N_19142,N_19103);
nand U20080 (N_20080,N_19016,N_18778);
or U20081 (N_20081,N_18550,N_18761);
and U20082 (N_20082,N_18092,N_17749);
nor U20083 (N_20083,N_19027,N_19161);
xor U20084 (N_20084,N_19683,N_18763);
xor U20085 (N_20085,N_18343,N_19496);
nor U20086 (N_20086,N_18621,N_19889);
and U20087 (N_20087,N_19239,N_18821);
nand U20088 (N_20088,N_18293,N_19536);
nand U20089 (N_20089,N_19508,N_18767);
or U20090 (N_20090,N_19426,N_19751);
and U20091 (N_20091,N_18504,N_17952);
and U20092 (N_20092,N_17801,N_18496);
nand U20093 (N_20093,N_19456,N_19742);
and U20094 (N_20094,N_19063,N_19549);
nor U20095 (N_20095,N_19754,N_17548);
nand U20096 (N_20096,N_18411,N_17948);
nand U20097 (N_20097,N_18667,N_19781);
nand U20098 (N_20098,N_19913,N_18789);
nor U20099 (N_20099,N_17826,N_19824);
or U20100 (N_20100,N_18403,N_19703);
xnor U20101 (N_20101,N_17772,N_18328);
nor U20102 (N_20102,N_19033,N_18552);
and U20103 (N_20103,N_19740,N_18298);
or U20104 (N_20104,N_18180,N_18197);
and U20105 (N_20105,N_19361,N_17865);
and U20106 (N_20106,N_19577,N_18852);
nor U20107 (N_20107,N_17862,N_19424);
and U20108 (N_20108,N_17904,N_18948);
nor U20109 (N_20109,N_19241,N_18861);
xnor U20110 (N_20110,N_18259,N_19287);
and U20111 (N_20111,N_17616,N_19855);
nor U20112 (N_20112,N_19058,N_19592);
or U20113 (N_20113,N_17879,N_18094);
nand U20114 (N_20114,N_19880,N_17934);
and U20115 (N_20115,N_18739,N_18346);
nand U20116 (N_20116,N_17991,N_19362);
xnor U20117 (N_20117,N_17957,N_19466);
and U20118 (N_20118,N_18315,N_18434);
nand U20119 (N_20119,N_18146,N_19166);
or U20120 (N_20120,N_19042,N_19074);
and U20121 (N_20121,N_17732,N_19951);
and U20122 (N_20122,N_18028,N_19158);
or U20123 (N_20123,N_18872,N_17715);
nor U20124 (N_20124,N_17676,N_19756);
nor U20125 (N_20125,N_18507,N_19517);
and U20126 (N_20126,N_17657,N_19180);
nand U20127 (N_20127,N_18466,N_18719);
and U20128 (N_20128,N_18314,N_19495);
nor U20129 (N_20129,N_18039,N_18270);
and U20130 (N_20130,N_17529,N_18240);
and U20131 (N_20131,N_17604,N_19920);
nor U20132 (N_20132,N_18082,N_19313);
or U20133 (N_20133,N_19772,N_18164);
and U20134 (N_20134,N_18165,N_19867);
nor U20135 (N_20135,N_19143,N_18461);
nor U20136 (N_20136,N_19383,N_19544);
or U20137 (N_20137,N_19500,N_18568);
or U20138 (N_20138,N_17742,N_19865);
nand U20139 (N_20139,N_19531,N_19097);
nand U20140 (N_20140,N_19829,N_19597);
nand U20141 (N_20141,N_19538,N_19271);
nand U20142 (N_20142,N_18662,N_19875);
and U20143 (N_20143,N_18295,N_18702);
nand U20144 (N_20144,N_18990,N_19689);
nand U20145 (N_20145,N_19374,N_18171);
and U20146 (N_20146,N_17889,N_18402);
nand U20147 (N_20147,N_19647,N_17563);
or U20148 (N_20148,N_19943,N_18991);
and U20149 (N_20149,N_18633,N_18864);
nand U20150 (N_20150,N_18912,N_19409);
nand U20151 (N_20151,N_19638,N_19641);
or U20152 (N_20152,N_19835,N_18144);
or U20153 (N_20153,N_17840,N_19395);
or U20154 (N_20154,N_18585,N_18311);
and U20155 (N_20155,N_18014,N_17762);
or U20156 (N_20156,N_19316,N_17841);
nand U20157 (N_20157,N_17705,N_19786);
nor U20158 (N_20158,N_18525,N_19553);
and U20159 (N_20159,N_18412,N_18004);
nand U20160 (N_20160,N_19182,N_19800);
xor U20161 (N_20161,N_18846,N_18765);
or U20162 (N_20162,N_18290,N_19376);
or U20163 (N_20163,N_19501,N_18442);
nand U20164 (N_20164,N_19050,N_18181);
nor U20165 (N_20165,N_19858,N_19682);
or U20166 (N_20166,N_19710,N_19454);
nor U20167 (N_20167,N_19939,N_19057);
xnor U20168 (N_20168,N_18997,N_19138);
nand U20169 (N_20169,N_19171,N_19803);
nand U20170 (N_20170,N_19381,N_19955);
and U20171 (N_20171,N_18758,N_18302);
xnor U20172 (N_20172,N_17839,N_18729);
or U20173 (N_20173,N_19486,N_19921);
xnor U20174 (N_20174,N_19814,N_17830);
nor U20175 (N_20175,N_17950,N_18822);
nand U20176 (N_20176,N_18121,N_19744);
or U20177 (N_20177,N_17852,N_17631);
and U20178 (N_20178,N_18620,N_18220);
nor U20179 (N_20179,N_18773,N_18289);
nor U20180 (N_20180,N_19422,N_19594);
and U20181 (N_20181,N_18494,N_19962);
xnor U20182 (N_20182,N_17573,N_19035);
and U20183 (N_20183,N_17905,N_17835);
or U20184 (N_20184,N_17729,N_18611);
xnor U20185 (N_20185,N_19981,N_17627);
or U20186 (N_20186,N_18506,N_18566);
nand U20187 (N_20187,N_19052,N_18177);
nand U20188 (N_20188,N_17975,N_19045);
nor U20189 (N_20189,N_19733,N_19372);
nand U20190 (N_20190,N_19432,N_19193);
nand U20191 (N_20191,N_18687,N_17845);
nand U20192 (N_20192,N_19709,N_18734);
or U20193 (N_20193,N_19768,N_18105);
and U20194 (N_20194,N_18536,N_19692);
xor U20195 (N_20195,N_19916,N_17601);
and U20196 (N_20196,N_18788,N_19928);
or U20197 (N_20197,N_19817,N_18320);
or U20198 (N_20198,N_19225,N_17511);
or U20199 (N_20199,N_19938,N_18210);
nor U20200 (N_20200,N_18455,N_17767);
or U20201 (N_20201,N_19923,N_18892);
and U20202 (N_20202,N_19192,N_19946);
and U20203 (N_20203,N_19819,N_17702);
nor U20204 (N_20204,N_18888,N_17764);
nor U20205 (N_20205,N_19712,N_19279);
nand U20206 (N_20206,N_18697,N_18617);
and U20207 (N_20207,N_17625,N_18996);
nor U20208 (N_20208,N_19202,N_18569);
nand U20209 (N_20209,N_18192,N_17938);
or U20210 (N_20210,N_19877,N_18128);
and U20211 (N_20211,N_19839,N_18663);
nor U20212 (N_20212,N_18034,N_18933);
xnor U20213 (N_20213,N_18631,N_19561);
nor U20214 (N_20214,N_18954,N_19739);
and U20215 (N_20215,N_19067,N_19603);
nand U20216 (N_20216,N_19494,N_19146);
and U20217 (N_20217,N_19465,N_18595);
nor U20218 (N_20218,N_17804,N_17753);
nor U20219 (N_20219,N_19310,N_17704);
nor U20220 (N_20220,N_18045,N_19725);
nand U20221 (N_20221,N_18457,N_19551);
xor U20222 (N_20222,N_19633,N_19613);
and U20223 (N_20223,N_17987,N_17994);
nor U20224 (N_20224,N_19224,N_17783);
nand U20225 (N_20225,N_19121,N_18489);
nand U20226 (N_20226,N_18970,N_18546);
nand U20227 (N_20227,N_18333,N_17535);
nand U20228 (N_20228,N_18243,N_18062);
nor U20229 (N_20229,N_19932,N_17527);
or U20230 (N_20230,N_19655,N_17787);
or U20231 (N_20231,N_18287,N_19303);
nor U20232 (N_20232,N_19284,N_19628);
nand U20233 (N_20233,N_19010,N_19073);
or U20234 (N_20234,N_18759,N_18932);
xor U20235 (N_20235,N_19643,N_18425);
and U20236 (N_20236,N_18648,N_18810);
or U20237 (N_20237,N_17505,N_18474);
or U20238 (N_20238,N_19542,N_19915);
nor U20239 (N_20239,N_17810,N_17680);
xor U20240 (N_20240,N_19713,N_18326);
nor U20241 (N_20241,N_17893,N_18675);
nor U20242 (N_20242,N_17915,N_19231);
xor U20243 (N_20243,N_19559,N_17972);
and U20244 (N_20244,N_18891,N_19608);
nor U20245 (N_20245,N_18006,N_19236);
xnor U20246 (N_20246,N_19838,N_19407);
and U20247 (N_20247,N_17528,N_17565);
or U20248 (N_20248,N_19293,N_18236);
nand U20249 (N_20249,N_19695,N_18635);
nand U20250 (N_20250,N_18584,N_17907);
and U20251 (N_20251,N_18505,N_19799);
nand U20252 (N_20252,N_18252,N_19328);
nor U20253 (N_20253,N_19468,N_18969);
nor U20254 (N_20254,N_18196,N_18993);
nand U20255 (N_20255,N_17901,N_18166);
and U20256 (N_20256,N_19043,N_18741);
and U20257 (N_20257,N_18280,N_19047);
or U20258 (N_20258,N_18469,N_19862);
or U20259 (N_20259,N_18807,N_18735);
nor U20260 (N_20260,N_17926,N_18445);
and U20261 (N_20261,N_18055,N_18652);
nor U20262 (N_20262,N_19081,N_18570);
xor U20263 (N_20263,N_18873,N_19770);
nand U20264 (N_20264,N_19165,N_19782);
or U20265 (N_20265,N_19114,N_17647);
and U20266 (N_20266,N_19404,N_18387);
and U20267 (N_20267,N_17723,N_18379);
or U20268 (N_20268,N_19746,N_18397);
nand U20269 (N_20269,N_18117,N_19415);
nor U20270 (N_20270,N_19579,N_17812);
or U20271 (N_20271,N_17860,N_17793);
nor U20272 (N_20272,N_19318,N_19498);
or U20273 (N_20273,N_17884,N_19723);
or U20274 (N_20274,N_19449,N_19954);
nor U20275 (N_20275,N_18638,N_17946);
xnor U20276 (N_20276,N_18430,N_19154);
or U20277 (N_20277,N_18726,N_18830);
and U20278 (N_20278,N_17559,N_19758);
nand U20279 (N_20279,N_19526,N_17998);
nand U20280 (N_20280,N_19028,N_18798);
nor U20281 (N_20281,N_19995,N_19207);
nand U20282 (N_20282,N_17936,N_18041);
or U20283 (N_20283,N_18129,N_19297);
nand U20284 (N_20284,N_18053,N_17751);
and U20285 (N_20285,N_18883,N_19257);
nor U20286 (N_20286,N_19094,N_18720);
and U20287 (N_20287,N_19054,N_19490);
and U20288 (N_20288,N_19964,N_18254);
and U20289 (N_20289,N_17874,N_18683);
and U20290 (N_20290,N_17791,N_18112);
and U20291 (N_20291,N_18653,N_18470);
and U20292 (N_20292,N_17965,N_19323);
and U20293 (N_20293,N_17518,N_18943);
nor U20294 (N_20294,N_18309,N_18625);
or U20295 (N_20295,N_19775,N_18539);
nor U20296 (N_20296,N_18318,N_18042);
nand U20297 (N_20297,N_18561,N_18389);
or U20298 (N_20298,N_18354,N_18188);
nor U20299 (N_20299,N_18078,N_17993);
and U20300 (N_20300,N_17731,N_18095);
nand U20301 (N_20301,N_17718,N_18876);
nand U20302 (N_20302,N_18900,N_19522);
or U20303 (N_20303,N_17756,N_18960);
or U20304 (N_20304,N_17556,N_19320);
nor U20305 (N_20305,N_19879,N_17825);
or U20306 (N_20306,N_18277,N_18206);
or U20307 (N_20307,N_18145,N_19240);
nor U20308 (N_20308,N_19621,N_18151);
or U20309 (N_20309,N_17591,N_18752);
and U20310 (N_20310,N_17611,N_19200);
or U20311 (N_20311,N_18725,N_18829);
or U20312 (N_20312,N_19760,N_18865);
or U20313 (N_20313,N_17920,N_17925);
nor U20314 (N_20314,N_18911,N_18685);
nand U20315 (N_20315,N_19089,N_19208);
nor U20316 (N_20316,N_19299,N_19774);
xnor U20317 (N_20317,N_19779,N_19777);
or U20318 (N_20318,N_18061,N_17503);
nand U20319 (N_20319,N_18433,N_19262);
or U20320 (N_20320,N_18701,N_18715);
nor U20321 (N_20321,N_18338,N_17512);
or U20322 (N_20322,N_19115,N_19298);
and U20323 (N_20323,N_19809,N_17551);
or U20324 (N_20324,N_18058,N_18400);
and U20325 (N_20325,N_17522,N_18271);
nand U20326 (N_20326,N_18202,N_18258);
or U20327 (N_20327,N_18643,N_17891);
or U20328 (N_20328,N_19974,N_19030);
nand U20329 (N_20329,N_18499,N_18732);
xnor U20330 (N_20330,N_17615,N_18869);
xnor U20331 (N_20331,N_18509,N_18921);
nand U20332 (N_20332,N_19791,N_19872);
nand U20333 (N_20333,N_18362,N_19873);
nand U20334 (N_20334,N_18669,N_18111);
nand U20335 (N_20335,N_17653,N_19321);
nand U20336 (N_20336,N_19223,N_19140);
xor U20337 (N_20337,N_19717,N_18711);
nand U20338 (N_20338,N_19598,N_19525);
nand U20339 (N_20339,N_18564,N_19355);
and U20340 (N_20340,N_18794,N_19895);
nor U20341 (N_20341,N_19375,N_19228);
or U20342 (N_20342,N_19793,N_18626);
nand U20343 (N_20343,N_19111,N_18882);
or U20344 (N_20344,N_19371,N_18574);
or U20345 (N_20345,N_17969,N_17813);
and U20346 (N_20346,N_18918,N_17797);
or U20347 (N_20347,N_19615,N_19132);
nand U20348 (N_20348,N_17917,N_18690);
or U20349 (N_20349,N_19090,N_19445);
or U20350 (N_20350,N_18958,N_19730);
xnor U20351 (N_20351,N_19327,N_19077);
or U20352 (N_20352,N_17586,N_18072);
nand U20353 (N_20353,N_19162,N_19024);
nand U20354 (N_20354,N_17550,N_19976);
nand U20355 (N_20355,N_19181,N_18070);
or U20356 (N_20356,N_17808,N_18345);
nand U20357 (N_20357,N_17638,N_17691);
nor U20358 (N_20358,N_18493,N_19541);
or U20359 (N_20359,N_18590,N_18123);
and U20360 (N_20360,N_19163,N_19459);
nor U20361 (N_20361,N_19272,N_17780);
and U20362 (N_20362,N_19126,N_19993);
and U20363 (N_20363,N_18380,N_17900);
and U20364 (N_20364,N_18530,N_18723);
nand U20365 (N_20365,N_18994,N_17931);
xnor U20366 (N_20366,N_19177,N_18919);
and U20367 (N_20367,N_19452,N_19296);
nor U20368 (N_20368,N_19159,N_18842);
or U20369 (N_20369,N_19899,N_18670);
nor U20370 (N_20370,N_18705,N_19591);
and U20371 (N_20371,N_19892,N_18571);
nand U20372 (N_20372,N_19353,N_17916);
and U20373 (N_20373,N_18949,N_19651);
nand U20374 (N_20374,N_18419,N_19509);
nand U20375 (N_20375,N_19317,N_18407);
and U20376 (N_20376,N_18404,N_18294);
or U20377 (N_20377,N_18424,N_18781);
or U20378 (N_20378,N_18141,N_19385);
and U20379 (N_20379,N_17778,N_19392);
or U20380 (N_20380,N_18714,N_18203);
nand U20381 (N_20381,N_17803,N_18526);
nor U20382 (N_20382,N_19277,N_19635);
and U20383 (N_20383,N_18441,N_19230);
nor U20384 (N_20384,N_19771,N_18490);
or U20385 (N_20385,N_17966,N_17698);
nor U20386 (N_20386,N_18820,N_19155);
nor U20387 (N_20387,N_19741,N_19186);
and U20388 (N_20388,N_19199,N_19267);
nor U20389 (N_20389,N_18335,N_17894);
nand U20390 (N_20390,N_18414,N_18415);
and U20391 (N_20391,N_18340,N_19876);
nand U20392 (N_20392,N_19141,N_19464);
and U20393 (N_20393,N_17538,N_18832);
nand U20394 (N_20394,N_19255,N_19188);
xor U20395 (N_20395,N_18514,N_19965);
xnor U20396 (N_20396,N_19078,N_19792);
or U20397 (N_20397,N_18248,N_18350);
and U20398 (N_20398,N_18109,N_17681);
nor U20399 (N_20399,N_18547,N_19100);
and U20400 (N_20400,N_18986,N_18768);
nand U20401 (N_20401,N_18327,N_18565);
nand U20402 (N_20402,N_19825,N_19380);
or U20403 (N_20403,N_17985,N_19585);
nor U20404 (N_20404,N_18782,N_17906);
and U20405 (N_20405,N_18100,N_19804);
or U20406 (N_20406,N_17903,N_18205);
nor U20407 (N_20407,N_19039,N_19988);
nor U20408 (N_20408,N_18906,N_17560);
and U20409 (N_20409,N_17855,N_18291);
nor U20410 (N_20410,N_18366,N_19480);
xor U20411 (N_20411,N_19607,N_17716);
nand U20412 (N_20412,N_17589,N_19471);
nand U20413 (N_20413,N_18790,N_17520);
xor U20414 (N_20414,N_19416,N_18558);
or U20415 (N_20415,N_19338,N_18106);
xor U20416 (N_20416,N_18049,N_18437);
nand U20417 (N_20417,N_18680,N_17805);
nand U20418 (N_20418,N_19485,N_17622);
or U20419 (N_20419,N_17871,N_18330);
or U20420 (N_20420,N_18541,N_17635);
or U20421 (N_20421,N_18381,N_19684);
and U20422 (N_20422,N_18059,N_18033);
nand U20423 (N_20423,N_17763,N_18791);
nor U20424 (N_20424,N_18760,N_18193);
nor U20425 (N_20425,N_18871,N_18088);
nor U20426 (N_20426,N_18839,N_18334);
nand U20427 (N_20427,N_17571,N_19902);
nand U20428 (N_20428,N_17544,N_18024);
or U20429 (N_20429,N_18962,N_19187);
nand U20430 (N_20430,N_17597,N_19900);
nand U20431 (N_20431,N_19367,N_17566);
and U20432 (N_20432,N_19157,N_18168);
xnor U20433 (N_20433,N_18102,N_19528);
or U20434 (N_20434,N_19442,N_19731);
nor U20435 (N_20435,N_17822,N_19034);
or U20436 (N_20436,N_19344,N_17848);
or U20437 (N_20437,N_18691,N_17922);
or U20438 (N_20438,N_19031,N_17937);
nand U20439 (N_20439,N_18535,N_19391);
nor U20440 (N_20440,N_19798,N_18301);
nand U20441 (N_20441,N_18936,N_17674);
nor U20442 (N_20442,N_17648,N_18162);
nand U20443 (N_20443,N_19311,N_19204);
nand U20444 (N_20444,N_19986,N_18537);
nor U20445 (N_20445,N_18534,N_18071);
and U20446 (N_20446,N_18602,N_19379);
or U20447 (N_20447,N_19649,N_17515);
nor U20448 (N_20448,N_18809,N_18099);
or U20449 (N_20449,N_17927,N_19469);
nand U20450 (N_20450,N_18370,N_19612);
nand U20451 (N_20451,N_19562,N_18651);
nor U20452 (N_20452,N_17935,N_19983);
and U20453 (N_20453,N_19125,N_17782);
nand U20454 (N_20454,N_17743,N_18849);
and U20455 (N_20455,N_17620,N_19840);
nand U20456 (N_20456,N_18800,N_18929);
nand U20457 (N_20457,N_17533,N_18264);
xor U20458 (N_20458,N_17788,N_19563);
or U20459 (N_20459,N_19832,N_17609);
nand U20460 (N_20460,N_18840,N_18805);
and U20461 (N_20461,N_17933,N_18609);
and U20462 (N_20462,N_18952,N_19145);
or U20463 (N_20463,N_17612,N_18737);
or U20464 (N_20464,N_18011,N_19656);
nor U20465 (N_20465,N_18678,N_17532);
nor U20466 (N_20466,N_17567,N_18172);
and U20467 (N_20467,N_18398,N_19854);
nor U20468 (N_20468,N_18031,N_19474);
nor U20469 (N_20469,N_18655,N_19936);
nor U20470 (N_20470,N_19811,N_19686);
nor U20471 (N_20471,N_18879,N_17843);
nand U20472 (N_20472,N_18613,N_19258);
and U20473 (N_20473,N_18783,N_18736);
or U20474 (N_20474,N_17642,N_18485);
nand U20475 (N_20475,N_19661,N_18272);
nand U20476 (N_20476,N_18169,N_19715);
or U20477 (N_20477,N_19360,N_18361);
nor U20478 (N_20478,N_19191,N_18901);
nor U20479 (N_20479,N_17558,N_19663);
nand U20480 (N_20480,N_19634,N_18592);
nand U20481 (N_20481,N_18043,N_19351);
or U20482 (N_20482,N_17695,N_19654);
nor U20483 (N_20483,N_18920,N_19226);
xnor U20484 (N_20484,N_18951,N_19743);
and U20485 (N_20485,N_18351,N_18817);
nand U20486 (N_20486,N_19307,N_18754);
and U20487 (N_20487,N_18373,N_18523);
nor U20488 (N_20488,N_18237,N_18632);
or U20489 (N_20489,N_19716,N_17986);
or U20490 (N_20490,N_19929,N_18325);
nor U20491 (N_20491,N_18671,N_19477);
or U20492 (N_20492,N_17864,N_17944);
nor U20493 (N_20493,N_17728,N_18356);
nor U20494 (N_20494,N_19173,N_18157);
or U20495 (N_20495,N_17711,N_19040);
or U20496 (N_20496,N_18023,N_17572);
and U20497 (N_20497,N_18246,N_18922);
or U20498 (N_20498,N_19680,N_19679);
and U20499 (N_20499,N_19384,N_19958);
nand U20500 (N_20500,N_19336,N_18357);
xnor U20501 (N_20501,N_18423,N_17883);
nor U20502 (N_20502,N_19534,N_19513);
xnor U20503 (N_20503,N_18222,N_19419);
or U20504 (N_20504,N_18015,N_18134);
and U20505 (N_20505,N_17679,N_18728);
nand U20506 (N_20506,N_19605,N_17541);
nor U20507 (N_20507,N_19168,N_17692);
or U20508 (N_20508,N_19018,N_18556);
nor U20509 (N_20509,N_17606,N_19535);
nor U20510 (N_20510,N_18075,N_18375);
nand U20511 (N_20511,N_18984,N_19124);
nor U20512 (N_20512,N_19167,N_19022);
xnor U20513 (N_20513,N_19914,N_18358);
nor U20514 (N_20514,N_18854,N_19053);
or U20515 (N_20515,N_18957,N_19301);
and U20516 (N_20516,N_19588,N_17823);
nor U20517 (N_20517,N_18747,N_18393);
nor U20518 (N_20518,N_19640,N_19062);
xor U20519 (N_20519,N_17675,N_18916);
or U20520 (N_20520,N_18636,N_17699);
nor U20521 (N_20521,N_17690,N_17670);
nor U20522 (N_20522,N_17740,N_17523);
nand U20523 (N_20523,N_18142,N_19108);
or U20524 (N_20524,N_18935,N_17897);
nand U20525 (N_20525,N_18487,N_17771);
and U20526 (N_20526,N_19623,N_18925);
xor U20527 (N_20527,N_18693,N_18743);
or U20528 (N_20528,N_17717,N_19305);
nor U20529 (N_20529,N_19427,N_19762);
and U20530 (N_20530,N_18517,N_19738);
nand U20531 (N_20531,N_19967,N_18159);
nand U20532 (N_20532,N_19084,N_18775);
nor U20533 (N_20533,N_18902,N_18019);
or U20534 (N_20534,N_19769,N_18589);
or U20535 (N_20535,N_19127,N_18646);
nand U20536 (N_20536,N_19941,N_19665);
or U20537 (N_20537,N_18009,N_19339);
nor U20538 (N_20538,N_18395,N_19219);
or U20539 (N_20539,N_19860,N_17685);
and U20540 (N_20540,N_18348,N_18874);
or U20541 (N_20541,N_19514,N_18050);
nand U20542 (N_20542,N_17815,N_18844);
xnor U20543 (N_20543,N_18154,N_18221);
nand U20544 (N_20544,N_18980,N_19748);
nor U20545 (N_20545,N_18831,N_17701);
nor U20546 (N_20546,N_19023,N_17833);
xor U20547 (N_20547,N_18578,N_17673);
or U20548 (N_20548,N_18727,N_19133);
and U20549 (N_20549,N_19315,N_17776);
or U20550 (N_20550,N_18209,N_19413);
or U20551 (N_20551,N_18784,N_19343);
xnor U20552 (N_20552,N_19687,N_19778);
or U20553 (N_20553,N_19253,N_19396);
nand U20554 (N_20554,N_17768,N_17956);
xor U20555 (N_20555,N_19366,N_18813);
nand U20556 (N_20556,N_17689,N_18841);
or U20557 (N_20557,N_17700,N_19831);
nor U20558 (N_20558,N_17759,N_17870);
nor U20559 (N_20559,N_19574,N_19669);
or U20560 (N_20560,N_19430,N_17652);
nand U20561 (N_20561,N_17842,N_17888);
or U20562 (N_20562,N_19953,N_18392);
nand U20563 (N_20563,N_18591,N_19933);
nand U20564 (N_20564,N_17632,N_19348);
or U20565 (N_20565,N_18175,N_18603);
nor U20566 (N_20566,N_18332,N_19763);
nor U20567 (N_20567,N_19288,N_19925);
nand U20568 (N_20568,N_18596,N_17629);
xor U20569 (N_20569,N_19980,N_17868);
nor U20570 (N_20570,N_18204,N_19991);
nor U20571 (N_20571,N_19265,N_19711);
and U20572 (N_20572,N_19457,N_18020);
nor U20573 (N_20573,N_17521,N_19812);
or U20574 (N_20574,N_17847,N_18629);
nor U20575 (N_20575,N_18239,N_17898);
and U20576 (N_20576,N_19044,N_18856);
and U20577 (N_20577,N_18860,N_19079);
xor U20578 (N_20578,N_18532,N_17811);
or U20579 (N_20579,N_19333,N_19985);
nor U20580 (N_20580,N_18606,N_18497);
or U20581 (N_20581,N_18002,N_17861);
nand U20582 (N_20582,N_18668,N_18107);
nand U20583 (N_20583,N_18890,N_17543);
nand U20584 (N_20584,N_17646,N_19493);
nand U20585 (N_20585,N_18322,N_18477);
nand U20586 (N_20586,N_19601,N_18614);
nor U20587 (N_20587,N_17596,N_18017);
nor U20588 (N_20588,N_18527,N_19583);
and U20589 (N_20589,N_18155,N_18420);
nand U20590 (N_20590,N_17828,N_19350);
xnor U20591 (N_20591,N_19358,N_17819);
nand U20592 (N_20592,N_17554,N_17669);
nand U20593 (N_20593,N_19274,N_18273);
and U20594 (N_20594,N_18447,N_18944);
nand U20595 (N_20595,N_19957,N_19606);
or U20596 (N_20596,N_19706,N_18583);
nand U20597 (N_20597,N_19572,N_17605);
or U20598 (N_20598,N_18207,N_18253);
xor U20599 (N_20599,N_19325,N_19102);
nor U20600 (N_20600,N_19620,N_19281);
nand U20601 (N_20601,N_18021,N_18903);
and U20602 (N_20602,N_18413,N_19238);
nor U20603 (N_20603,N_18868,N_19373);
nand U20604 (N_20604,N_18619,N_17800);
nor U20605 (N_20605,N_18241,N_19912);
and U20606 (N_20606,N_19973,N_19826);
and U20607 (N_20607,N_19227,N_17552);
nor U20608 (N_20608,N_19842,N_19475);
xnor U20609 (N_20609,N_19506,N_19662);
xnor U20610 (N_20610,N_18835,N_19554);
or U20611 (N_20611,N_19701,N_18941);
or U20612 (N_20612,N_19629,N_19573);
nor U20613 (N_20613,N_18376,N_18108);
and U20614 (N_20614,N_18915,N_17555);
xnor U20615 (N_20615,N_18699,N_17671);
xor U20616 (N_20616,N_19691,N_19308);
xor U20617 (N_20617,N_18533,N_18201);
nand U20618 (N_20618,N_19304,N_19833);
nand U20619 (N_20619,N_19570,N_17942);
and U20620 (N_20620,N_17524,N_18232);
and U20621 (N_20621,N_18003,N_18097);
nand U20622 (N_20622,N_18217,N_17785);
or U20623 (N_20623,N_18870,N_19497);
xnor U20624 (N_20624,N_19150,N_18047);
nand U20625 (N_20625,N_19418,N_19048);
nor U20626 (N_20626,N_19924,N_18363);
and U20627 (N_20627,N_18905,N_18909);
nand U20628 (N_20628,N_19697,N_19198);
nor U20629 (N_20629,N_19945,N_18156);
nand U20630 (N_20630,N_17857,N_17545);
nor U20631 (N_20631,N_19245,N_18803);
nand U20632 (N_20632,N_18946,N_18278);
and U20633 (N_20633,N_18360,N_19558);
and U20634 (N_20634,N_17747,N_19960);
xnor U20635 (N_20635,N_17990,N_18894);
nor U20636 (N_20636,N_19388,N_19537);
and U20637 (N_20637,N_18101,N_18475);
xnor U20638 (N_20638,N_19003,N_19672);
nor U20639 (N_20639,N_19547,N_18599);
nor U20640 (N_20640,N_19011,N_18850);
nand U20641 (N_20641,N_18618,N_17961);
nor U20642 (N_20642,N_18026,N_19211);
and U20643 (N_20643,N_18623,N_18482);
or U20644 (N_20644,N_19278,N_19319);
and U20645 (N_20645,N_19489,N_18689);
nor U20646 (N_20646,N_19984,N_19856);
nor U20647 (N_20647,N_19764,N_17786);
nand U20648 (N_20648,N_18793,N_18286);
or U20649 (N_20649,N_19604,N_17974);
and U20650 (N_20650,N_17630,N_18310);
nor U20651 (N_20651,N_17943,N_19841);
nand U20652 (N_20652,N_17587,N_17694);
or U20653 (N_20653,N_18284,N_19447);
nand U20654 (N_20654,N_18927,N_18945);
nand U20655 (N_20655,N_18880,N_18979);
nor U20656 (N_20656,N_18703,N_18910);
xor U20657 (N_20657,N_19205,N_19896);
nor U20658 (N_20658,N_17892,N_18543);
or U20659 (N_20659,N_18040,N_17955);
nor U20660 (N_20660,N_18999,N_19734);
xor U20661 (N_20661,N_19670,N_17794);
nand U20662 (N_20662,N_18052,N_19144);
nor U20663 (N_20663,N_19989,N_19164);
nand U20664 (N_20664,N_19796,N_18153);
nor U20665 (N_20665,N_18124,N_18150);
nand U20666 (N_20666,N_17818,N_18531);
nor U20667 (N_20667,N_17941,N_19453);
nand U20668 (N_20668,N_19332,N_18956);
xor U20669 (N_20669,N_17713,N_18484);
nor U20670 (N_20670,N_19708,N_17661);
nand U20671 (N_20671,N_19852,N_19473);
and U20672 (N_20672,N_18551,N_18679);
and U20673 (N_20673,N_18501,N_18746);
or U20674 (N_20674,N_19106,N_19055);
and U20675 (N_20675,N_17504,N_17655);
xor U20676 (N_20676,N_19978,N_18538);
nor U20677 (N_20677,N_18312,N_19847);
nor U20678 (N_20678,N_18304,N_19590);
xnor U20679 (N_20679,N_19148,N_17549);
nor U20680 (N_20680,N_19539,N_17770);
nand U20681 (N_20681,N_19291,N_18751);
and U20682 (N_20682,N_18038,N_18369);
nand U20683 (N_20683,N_17588,N_19690);
nand U20684 (N_20684,N_19091,N_18965);
nor U20685 (N_20685,N_19894,N_18085);
or U20686 (N_20686,N_18630,N_19685);
nand U20687 (N_20687,N_19694,N_19616);
nand U20688 (N_20688,N_17838,N_19503);
and U20689 (N_20689,N_19970,N_17876);
nor U20690 (N_20690,N_17721,N_17981);
and U20691 (N_20691,N_19269,N_18981);
nor U20692 (N_20692,N_18516,N_19637);
xor U20693 (N_20693,N_19324,N_19170);
or U20694 (N_20694,N_18640,N_19472);
nand U20695 (N_20695,N_18262,N_19237);
and U20696 (N_20696,N_18510,N_18223);
xor U20697 (N_20697,N_19206,N_18924);
nor U20698 (N_20698,N_19956,N_19688);
xnor U20699 (N_20699,N_19836,N_19290);
nor U20700 (N_20700,N_18429,N_18359);
nor U20701 (N_20701,N_18382,N_17547);
nand U20702 (N_20702,N_17501,N_18588);
and U20703 (N_20703,N_19444,N_17553);
and U20704 (N_20704,N_19306,N_17686);
nor U20705 (N_20705,N_18907,N_18283);
nor U20706 (N_20706,N_19502,N_17911);
xor U20707 (N_20707,N_18989,N_18992);
and U20708 (N_20708,N_18607,N_18567);
nand U20709 (N_20709,N_18195,N_17706);
nor U20710 (N_20710,N_19636,N_18030);
or U20711 (N_20711,N_18439,N_19926);
nand U20712 (N_20712,N_18176,N_17834);
and U20713 (N_20713,N_18456,N_19234);
and U20714 (N_20714,N_19524,N_19961);
nand U20715 (N_20715,N_17724,N_19334);
xnor U20716 (N_20716,N_17582,N_19314);
nor U20717 (N_20717,N_18481,N_18814);
and U20718 (N_20718,N_18740,N_19565);
nand U20719 (N_20719,N_18051,N_18036);
nor U20720 (N_20720,N_17816,N_18917);
or U20721 (N_20721,N_18093,N_19005);
xnor U20722 (N_20722,N_18656,N_17651);
and U20723 (N_20723,N_18261,N_19195);
xor U20724 (N_20724,N_18770,N_18857);
nor U20725 (N_20725,N_19905,N_19431);
or U20726 (N_20726,N_18463,N_18818);
xor U20727 (N_20727,N_19331,N_19934);
nand U20728 (N_20728,N_17766,N_18113);
and U20729 (N_20729,N_18344,N_18698);
and U20730 (N_20730,N_17958,N_19673);
nand U20731 (N_20731,N_18087,N_19658);
and U20732 (N_20732,N_18562,N_19174);
xnor U20733 (N_20733,N_19671,N_19657);
and U20734 (N_20734,N_18468,N_18601);
nor U20735 (N_20735,N_17709,N_18491);
nand U20736 (N_20736,N_18187,N_17909);
xnor U20737 (N_20737,N_19947,N_18733);
xnor U20738 (N_20738,N_19752,N_17637);
nand U20739 (N_20739,N_19178,N_19548);
nand U20740 (N_20740,N_17683,N_19992);
xor U20741 (N_20741,N_19172,N_19555);
xnor U20742 (N_20742,N_18978,N_18191);
or U20743 (N_20743,N_19660,N_19611);
nor U20744 (N_20744,N_19484,N_18973);
or U20745 (N_20745,N_19593,N_18594);
and U20746 (N_20746,N_19041,N_18384);
xnor U20747 (N_20747,N_17949,N_19190);
xnor U20748 (N_20748,N_18938,N_18214);
or U20749 (N_20749,N_18779,N_18235);
or U20750 (N_20750,N_17895,N_19259);
or U20751 (N_20751,N_19417,N_19300);
or U20752 (N_20752,N_18426,N_19512);
nor U20753 (N_20753,N_18586,N_18418);
nor U20754 (N_20754,N_17737,N_17963);
and U20755 (N_20755,N_19256,N_19584);
nor U20756 (N_20756,N_19569,N_19749);
nand U20757 (N_20757,N_17836,N_19356);
nor U20758 (N_20758,N_19130,N_19911);
and U20759 (N_20759,N_19887,N_18688);
xor U20760 (N_20760,N_19529,N_19273);
nor U20761 (N_20761,N_18961,N_18889);
and U20762 (N_20762,N_18234,N_18642);
and U20763 (N_20763,N_19783,N_19888);
nand U20764 (N_20764,N_18673,N_18213);
nand U20765 (N_20765,N_17912,N_19354);
nand U20766 (N_20766,N_19666,N_18285);
or U20767 (N_20767,N_19013,N_18769);
nor U20768 (N_20768,N_19864,N_17940);
nor U20769 (N_20769,N_19893,N_17799);
or U20770 (N_20770,N_17902,N_19927);
nand U20771 (N_20771,N_18650,N_17636);
nand U20772 (N_20772,N_19411,N_17846);
nand U20773 (N_20773,N_18331,N_19446);
or U20774 (N_20774,N_19720,N_19072);
and U20775 (N_20775,N_18079,N_18063);
nor U20776 (N_20776,N_18119,N_19019);
or U20777 (N_20777,N_17736,N_18483);
xor U20778 (N_20778,N_18478,N_18355);
nor U20779 (N_20779,N_18837,N_17873);
and U20780 (N_20780,N_19378,N_18329);
or U20781 (N_20781,N_18557,N_18473);
nand U20782 (N_20782,N_18016,N_18845);
nand U20783 (N_20783,N_18118,N_18834);
xnor U20784 (N_20784,N_17856,N_19412);
nand U20785 (N_20785,N_18149,N_17656);
or U20786 (N_20786,N_17746,N_19441);
or U20787 (N_20787,N_19530,N_19394);
nand U20788 (N_20788,N_17774,N_18731);
or U20789 (N_20789,N_19196,N_18875);
and U20790 (N_20790,N_19488,N_18251);
nand U20791 (N_20791,N_19294,N_19881);
and U20792 (N_20792,N_17971,N_19082);
and U20793 (N_20793,N_19859,N_18459);
and U20794 (N_20794,N_19292,N_19268);
nor U20795 (N_20795,N_18605,N_18692);
nand U20796 (N_20796,N_19678,N_19568);
and U20797 (N_20797,N_18174,N_19564);
nor U20798 (N_20798,N_19705,N_19677);
nand U20799 (N_20799,N_18116,N_17930);
nor U20800 (N_20800,N_19377,N_19069);
xor U20801 (N_20801,N_18542,N_18064);
nor U20802 (N_20802,N_19909,N_17964);
nor U20803 (N_20803,N_17973,N_19646);
xor U20804 (N_20804,N_19659,N_18037);
or U20805 (N_20805,N_18438,N_18216);
xor U20806 (N_20806,N_17628,N_19105);
and U20807 (N_20807,N_18529,N_19175);
nor U20808 (N_20808,N_19653,N_18610);
or U20809 (N_20809,N_19797,N_19552);
and U20810 (N_20810,N_18498,N_17645);
or U20811 (N_20811,N_18208,N_18833);
and U20812 (N_20812,N_18843,N_18666);
nor U20813 (N_20813,N_19216,N_19959);
or U20814 (N_20814,N_19648,N_19868);
or U20815 (N_20815,N_18914,N_17668);
xnor U20816 (N_20816,N_18801,N_19871);
nor U20817 (N_20817,N_17508,N_18409);
and U20818 (N_20818,N_18686,N_19761);
xor U20819 (N_20819,N_17672,N_18069);
nand U20820 (N_20820,N_18339,N_19184);
and U20821 (N_20821,N_18367,N_19101);
nor U20822 (N_20822,N_18460,N_19667);
or U20823 (N_20823,N_18446,N_19369);
nand U20824 (N_20824,N_19461,N_18815);
nand U20825 (N_20825,N_18634,N_18825);
and U20826 (N_20826,N_19644,N_18066);
nor U20827 (N_20827,N_19059,N_19642);
xnor U20828 (N_20828,N_17667,N_19520);
or U20829 (N_20829,N_17583,N_19107);
or U20830 (N_20830,N_18137,N_19251);
xor U20831 (N_20831,N_17977,N_19618);
nor U20832 (N_20832,N_18000,N_18554);
xor U20833 (N_20833,N_18385,N_18940);
nand U20834 (N_20834,N_18307,N_18265);
or U20835 (N_20835,N_18013,N_17564);
nand U20836 (N_20836,N_18528,N_17570);
nor U20837 (N_20837,N_18096,N_17999);
nand U20838 (N_20838,N_18974,N_18563);
and U20839 (N_20839,N_19014,N_19152);
nand U20840 (N_20840,N_18612,N_19340);
nor U20841 (N_20841,N_18934,N_18130);
nor U20842 (N_20842,N_18684,N_19060);
xor U20843 (N_20843,N_19904,N_18300);
and U20844 (N_20844,N_19134,N_18453);
xnor U20845 (N_20845,N_18032,N_18676);
and U20846 (N_20846,N_18771,N_17744);
nor U20847 (N_20847,N_17996,N_18083);
or U20848 (N_20848,N_19462,N_18229);
or U20849 (N_20849,N_18215,N_18488);
or U20850 (N_20850,N_18495,N_19083);
nor U20851 (N_20851,N_18859,N_18717);
nand U20852 (N_20852,N_18057,N_18862);
nor U20853 (N_20853,N_18440,N_19085);
nor U20854 (N_20854,N_18257,N_18750);
and U20855 (N_20855,N_19580,N_19185);
or U20856 (N_20856,N_19406,N_19364);
and U20857 (N_20857,N_18465,N_18148);
or U20858 (N_20858,N_19015,N_19342);
nor U20859 (N_20859,N_19434,N_18226);
xor U20860 (N_20860,N_17590,N_18084);
nand U20861 (N_20861,N_17945,N_17849);
or U20862 (N_20862,N_19546,N_19365);
and U20863 (N_20863,N_18645,N_19408);
nand U20864 (N_20864,N_17784,N_17607);
and U20865 (N_20865,N_18388,N_18819);
nand U20866 (N_20866,N_19878,N_18250);
or U20867 (N_20867,N_19049,N_18560);
and U20868 (N_20868,N_19232,N_19463);
or U20869 (N_20869,N_19004,N_19732);
or U20870 (N_20870,N_18383,N_18238);
and U20871 (N_20871,N_18512,N_17734);
and U20872 (N_20872,N_18672,N_17619);
and U20873 (N_20873,N_19244,N_19414);
and U20874 (N_20874,N_17750,N_19996);
and U20875 (N_20875,N_19248,N_17745);
nand U20876 (N_20876,N_19747,N_19460);
or U20877 (N_20877,N_18796,N_19221);
or U20878 (N_20878,N_17959,N_19249);
or U20879 (N_20879,N_17584,N_17968);
nand U20880 (N_20880,N_17593,N_18963);
nor U20881 (N_20881,N_19065,N_19112);
or U20882 (N_20882,N_18540,N_19626);
nor U20883 (N_20883,N_17733,N_19922);
and U20884 (N_20884,N_19387,N_17982);
nor U20885 (N_20885,N_19632,N_17714);
and U20886 (N_20886,N_18928,N_19721);
and U20887 (N_20887,N_19704,N_19714);
and U20888 (N_20888,N_17693,N_18549);
or U20889 (N_20889,N_19487,N_18347);
nand U20890 (N_20890,N_17502,N_19851);
xor U20891 (N_20891,N_19610,N_18749);
nand U20892 (N_20892,N_19139,N_17979);
nand U20893 (N_20893,N_18577,N_18098);
nand U20894 (N_20894,N_18545,N_19818);
or U20895 (N_20895,N_17853,N_19302);
and U20896 (N_20896,N_18428,N_17710);
nand U20897 (N_20897,N_18518,N_19329);
and U20898 (N_20898,N_18707,N_18054);
or U20899 (N_20899,N_17877,N_17754);
or U20900 (N_20900,N_17859,N_18143);
or U20901 (N_20901,N_19201,N_17510);
nand U20902 (N_20902,N_18022,N_18242);
nand U20903 (N_20903,N_18744,N_17854);
nand U20904 (N_20904,N_19135,N_18522);
and U20905 (N_20905,N_18296,N_18454);
or U20906 (N_20906,N_18228,N_18365);
xnor U20907 (N_20907,N_19280,N_17517);
and U20908 (N_20908,N_18548,N_18886);
nor U20909 (N_20909,N_19882,N_18377);
xor U20910 (N_20910,N_18893,N_19987);
or U20911 (N_20911,N_17660,N_18709);
xor U20912 (N_20912,N_19214,N_17872);
or U20913 (N_20913,N_19942,N_19619);
xor U20914 (N_20914,N_18158,N_18225);
nor U20915 (N_20915,N_18305,N_18010);
nand U20916 (N_20916,N_19116,N_18580);
nand U20917 (N_20917,N_17851,N_19229);
nand U20918 (N_20918,N_18179,N_17643);
or U20919 (N_20919,N_18988,N_18657);
nor U20920 (N_20920,N_18774,N_17837);
or U20921 (N_20921,N_18263,N_18797);
and U20922 (N_20922,N_19505,N_18136);
or U20923 (N_20923,N_19834,N_19066);
and U20924 (N_20924,N_18256,N_17594);
or U20925 (N_20925,N_19589,N_17858);
xnor U20926 (N_20926,N_17677,N_19639);
xor U20927 (N_20927,N_18368,N_19702);
and U20928 (N_20928,N_17580,N_17682);
or U20929 (N_20929,N_17796,N_17887);
nand U20930 (N_20930,N_19602,N_19693);
nand U20931 (N_20931,N_19969,N_18756);
nand U20932 (N_20932,N_18303,N_18576);
nand U20933 (N_20933,N_19117,N_17678);
nor U20934 (N_20934,N_19420,N_19586);
nor U20935 (N_20935,N_17626,N_19076);
nand U20936 (N_20936,N_18555,N_18337);
or U20937 (N_20937,N_17540,N_18048);
or U20938 (N_20938,N_18007,N_19359);
and U20939 (N_20939,N_18190,N_18163);
nand U20940 (N_20940,N_19056,N_19910);
or U20941 (N_20941,N_19451,N_17639);
nand U20942 (N_20942,N_18628,N_18255);
xnor U20943 (N_20943,N_17992,N_19950);
nor U20944 (N_20944,N_19952,N_18877);
nor U20945 (N_20945,N_19890,N_17748);
nand U20946 (N_20946,N_19169,N_17650);
or U20947 (N_20947,N_18787,N_19122);
nand U20948 (N_20948,N_19789,N_18417);
nand U20949 (N_20949,N_19009,N_18931);
and U20950 (N_20950,N_18391,N_17932);
or U20951 (N_20951,N_19773,N_18987);
and U20952 (N_20952,N_19735,N_18249);
nand U20953 (N_20953,N_18282,N_19807);
nor U20954 (N_20954,N_19863,N_19400);
and U20955 (N_20955,N_18269,N_19813);
and U20956 (N_20956,N_19006,N_18170);
or U20957 (N_20957,N_19515,N_19571);
xor U20958 (N_20958,N_19788,N_19250);
nor U20959 (N_20959,N_19032,N_17509);
nand U20960 (N_20960,N_17574,N_19001);
nand U20961 (N_20961,N_18926,N_18126);
and U20962 (N_20962,N_19147,N_17773);
nor U20963 (N_20963,N_17610,N_19540);
nand U20964 (N_20964,N_18930,N_18755);
or U20965 (N_20965,N_19398,N_17995);
nand U20966 (N_20966,N_18122,N_18616);
and U20967 (N_20967,N_17921,N_19046);
nor U20968 (N_20968,N_19156,N_19940);
and U20969 (N_20969,N_17506,N_18520);
and U20970 (N_20970,N_18544,N_18908);
nor U20971 (N_20971,N_19625,N_17899);
nand U20972 (N_20972,N_17720,N_19246);
nor U20973 (N_20973,N_18371,N_19550);
and U20974 (N_20974,N_19997,N_18776);
or U20975 (N_20975,N_19264,N_19189);
xor U20976 (N_20976,N_18067,N_17536);
and U20977 (N_20977,N_19437,N_18939);
nor U20978 (N_20978,N_17603,N_17913);
and U20979 (N_20979,N_19560,N_19581);
nand U20980 (N_20980,N_18896,N_19393);
and U20981 (N_20981,N_18183,N_19399);
nand U20982 (N_20982,N_17939,N_18851);
nand U20983 (N_20983,N_18953,N_19903);
nand U20984 (N_20984,N_19151,N_19322);
nand U20985 (N_20985,N_19874,N_18738);
nor U20986 (N_20986,N_18231,N_17688);
xnor U20987 (N_20987,N_18503,N_19884);
xnor U20988 (N_20988,N_18135,N_18950);
nand U20989 (N_20989,N_17802,N_18942);
nor U20990 (N_20990,N_17769,N_17600);
and U20991 (N_20991,N_18581,N_19897);
nor U20992 (N_20992,N_19345,N_17757);
nor U20993 (N_20993,N_18995,N_17546);
nor U20994 (N_20994,N_18476,N_19737);
nor U20995 (N_20995,N_18139,N_18677);
or U20996 (N_20996,N_17978,N_18895);
nor U20997 (N_20997,N_17659,N_19759);
and U20998 (N_20998,N_18811,N_19403);
and U20999 (N_20999,N_17866,N_19254);
or U21000 (N_21000,N_18615,N_19566);
and U21001 (N_21001,N_18352,N_19736);
nand U21002 (N_21002,N_18422,N_19099);
nor U21003 (N_21003,N_17598,N_19286);
or U21004 (N_21004,N_18276,N_18827);
or U21005 (N_21005,N_19898,N_17924);
and U21006 (N_21006,N_18341,N_19949);
or U21007 (N_21007,N_18218,N_17775);
nand U21008 (N_21008,N_19160,N_19386);
nand U21009 (N_21009,N_18321,N_18125);
and U21010 (N_21010,N_17576,N_19917);
xnor U21011 (N_21011,N_19533,N_17980);
nand U21012 (N_21012,N_18786,N_18708);
or U21013 (N_21013,N_18076,N_17640);
nand U21014 (N_21014,N_18435,N_18826);
nor U21015 (N_21015,N_19368,N_17896);
nor U21016 (N_21016,N_17608,N_19919);
and U21017 (N_21017,N_19129,N_18977);
and U21018 (N_21018,N_18152,N_19179);
xnor U21019 (N_21019,N_18598,N_18317);
nor U21020 (N_21020,N_18138,N_17666);
nand U21021 (N_21021,N_19532,N_19567);
or U21022 (N_21022,N_18983,N_19776);
and U21023 (N_21023,N_18200,N_18604);
and U21024 (N_21024,N_19037,N_18696);
nor U21025 (N_21025,N_18898,N_19096);
and U21026 (N_21026,N_18274,N_19210);
and U21027 (N_21027,N_19433,N_19483);
and U21028 (N_21028,N_18132,N_17761);
and U21029 (N_21029,N_19853,N_17665);
or U21030 (N_21030,N_18297,N_19845);
and U21031 (N_21031,N_19131,N_17592);
or U21032 (N_21032,N_17730,N_19883);
or U21033 (N_21033,N_19120,N_19401);
nor U21034 (N_21034,N_19087,N_18762);
nand U21035 (N_21035,N_19007,N_19036);
and U21036 (N_21036,N_18268,N_17624);
nor U21037 (N_21037,N_18587,N_17739);
and U21038 (N_21038,N_18559,N_17577);
nor U21039 (N_21039,N_19785,N_17809);
nor U21040 (N_21040,N_17885,N_17827);
nand U21041 (N_21041,N_18724,N_19276);
and U21042 (N_21042,N_19370,N_17760);
or U21043 (N_21043,N_18519,N_18260);
xor U21044 (N_21044,N_18887,N_18374);
nand U21045 (N_21045,N_18046,N_17908);
xnor U21046 (N_21046,N_17882,N_19810);
or U21047 (N_21047,N_19999,N_17918);
xnor U21048 (N_21048,N_18753,N_18479);
and U21049 (N_21049,N_18764,N_17807);
xnor U21050 (N_21050,N_17697,N_18185);
nor U21051 (N_21051,N_19233,N_17561);
or U21052 (N_21052,N_18245,N_19885);
nor U21053 (N_21053,N_18682,N_19363);
or U21054 (N_21054,N_18665,N_19093);
and U21055 (N_21055,N_19519,N_19213);
or U21056 (N_21056,N_19700,N_17850);
nand U21057 (N_21057,N_19699,N_17579);
or U21058 (N_21058,N_19128,N_17989);
nor U21059 (N_21059,N_17712,N_19470);
xor U21060 (N_21060,N_19080,N_19617);
nand U21061 (N_21061,N_17617,N_18451);
nand U21062 (N_21062,N_19870,N_19652);
or U21063 (N_21063,N_17824,N_17708);
and U21064 (N_21064,N_17513,N_17602);
and U21065 (N_21065,N_19137,N_19235);
nor U21066 (N_21066,N_19511,N_18799);
nor U21067 (N_21067,N_17954,N_19504);
and U21068 (N_21068,N_17557,N_18462);
and U21069 (N_21069,N_19624,N_17829);
nand U21070 (N_21070,N_19012,N_19837);
xor U21071 (N_21071,N_17820,N_18658);
or U21072 (N_21072,N_19510,N_18390);
nand U21073 (N_21073,N_17519,N_19869);
nand U21074 (N_21074,N_18060,N_18964);
and U21075 (N_21075,N_19335,N_19784);
and U21076 (N_21076,N_19578,N_18828);
nand U21077 (N_21077,N_18660,N_19260);
nor U21078 (N_21078,N_19347,N_19718);
or U21079 (N_21079,N_17758,N_19008);
and U21080 (N_21080,N_18012,N_17507);
nor U21081 (N_21081,N_19443,N_19668);
nor U21082 (N_21082,N_18018,N_17526);
nor U21083 (N_21083,N_19312,N_18971);
xor U21084 (N_21084,N_18627,N_18881);
nor U21085 (N_21085,N_19061,N_18056);
and U21086 (N_21086,N_19243,N_18742);
nand U21087 (N_21087,N_17568,N_19118);
nand U21088 (N_21088,N_17662,N_17867);
nor U21089 (N_21089,N_18712,N_17531);
nand U21090 (N_21090,N_17585,N_18299);
nand U21091 (N_21091,N_19806,N_18323);
nor U21092 (N_21092,N_18838,N_18316);
and U21093 (N_21093,N_19212,N_17875);
nor U21094 (N_21094,N_18976,N_19971);
or U21095 (N_21095,N_19790,N_18230);
or U21096 (N_21096,N_19630,N_19439);
nand U21097 (N_21097,N_19423,N_18959);
nand U21098 (N_21098,N_18211,N_18449);
nand U21099 (N_21099,N_19029,N_17798);
or U21100 (N_21100,N_19478,N_19557);
and U21101 (N_21101,N_18713,N_18410);
and U21102 (N_21102,N_19765,N_19261);
nand U21103 (N_21103,N_18511,N_18091);
nor U21104 (N_21104,N_19247,N_18133);
and U21105 (N_21105,N_18008,N_17644);
nand U21106 (N_21106,N_18982,N_19390);
or U21107 (N_21107,N_17641,N_18823);
nand U21108 (N_21108,N_17633,N_18467);
xnor U21109 (N_21109,N_19098,N_19614);
or U21110 (N_21110,N_18804,N_18396);
nand U21111 (N_21111,N_18521,N_19820);
nand U21112 (N_21112,N_19827,N_17530);
and U21113 (N_21113,N_18182,N_17997);
nor U21114 (N_21114,N_18812,N_18824);
nand U21115 (N_21115,N_19979,N_18730);
and U21116 (N_21116,N_19516,N_19802);
and U21117 (N_21117,N_19436,N_18378);
nand U21118 (N_21118,N_18848,N_19203);
nand U21119 (N_21119,N_19750,N_19405);
nor U21120 (N_21120,N_18858,N_19935);
xor U21121 (N_21121,N_18077,N_18074);
and U21122 (N_21122,N_19674,N_19846);
and U21123 (N_21123,N_18637,N_18405);
or U21124 (N_21124,N_17649,N_17880);
nand U21125 (N_21125,N_19440,N_19123);
nor U21126 (N_21126,N_19582,N_18816);
or U21127 (N_21127,N_18044,N_19767);
or U21128 (N_21128,N_18899,N_18090);
and U21129 (N_21129,N_19972,N_19821);
and U21130 (N_21130,N_18766,N_17735);
nor U21131 (N_21131,N_18855,N_18998);
xnor U21132 (N_21132,N_18923,N_18104);
nor U21133 (N_21133,N_18575,N_19337);
or U21134 (N_21134,N_17890,N_19215);
nand U21135 (N_21135,N_18443,N_18073);
xor U21136 (N_21136,N_18472,N_17663);
or U21137 (N_21137,N_18080,N_19755);
nor U21138 (N_21138,N_19727,N_17726);
nor U21139 (N_21139,N_19931,N_18718);
or U21140 (N_21140,N_18199,N_18524);
nor U21141 (N_21141,N_19518,N_18114);
and U21142 (N_21142,N_19220,N_18985);
nor U21143 (N_21143,N_18748,N_18081);
nor U21144 (N_21144,N_17806,N_19402);
nor U21145 (N_21145,N_19109,N_19491);
and U21146 (N_21146,N_17613,N_19153);
xor U21147 (N_21147,N_17983,N_19595);
and U21148 (N_21148,N_18399,N_17621);
and U21149 (N_21149,N_18342,N_18313);
nor U21150 (N_21150,N_19545,N_19266);
nor U21151 (N_21151,N_19309,N_19575);
or U21152 (N_21152,N_17755,N_19450);
or U21153 (N_21153,N_19930,N_18745);
or U21154 (N_21154,N_18806,N_19136);
nor U21155 (N_21155,N_19263,N_19975);
nor U21156 (N_21156,N_18897,N_18579);
or U21157 (N_21157,N_18281,N_19176);
nand U21158 (N_21158,N_18275,N_17703);
or U21159 (N_21159,N_19780,N_18186);
nand U21160 (N_21160,N_19822,N_18654);
xnor U21161 (N_21161,N_18161,N_19295);
and U21162 (N_21162,N_18173,N_17790);
xnor U21163 (N_21163,N_19600,N_18444);
nor U21164 (N_21164,N_19757,N_17514);
nor U21165 (N_21165,N_19104,N_18904);
xor U21166 (N_21166,N_19766,N_19455);
or U21167 (N_21167,N_18777,N_18336);
or U21168 (N_21168,N_18065,N_17988);
and U21169 (N_21169,N_18884,N_18863);
or U21170 (N_21170,N_19908,N_19357);
nand U21171 (N_21171,N_19448,N_18372);
nand U21172 (N_21172,N_17687,N_17684);
xnor U21173 (N_21173,N_18622,N_19429);
or U21174 (N_21174,N_17795,N_19051);
or U21175 (N_21175,N_18600,N_17947);
nand U21176 (N_21176,N_19270,N_19726);
nor U21177 (N_21177,N_18068,N_18885);
and U21178 (N_21178,N_19217,N_19918);
xnor U21179 (N_21179,N_19857,N_19352);
or U21180 (N_21180,N_19183,N_19596);
and U21181 (N_21181,N_18431,N_18288);
and U21182 (N_21182,N_19681,N_18878);
nor U21183 (N_21183,N_17869,N_18198);
or U21184 (N_21184,N_17910,N_18178);
nand U21185 (N_21185,N_19458,N_18471);
and U21186 (N_21186,N_17976,N_17525);
nand U21187 (N_21187,N_19326,N_19349);
nand U21188 (N_21188,N_19968,N_19808);
or U21189 (N_21189,N_19527,N_19382);
nand U21190 (N_21190,N_17741,N_19844);
nor U21191 (N_21191,N_18515,N_17634);
xor U21192 (N_21192,N_18131,N_17752);
and U21193 (N_21193,N_19330,N_18947);
nor U21194 (N_21194,N_17562,N_18103);
nand U21195 (N_21195,N_18401,N_18279);
nor U21196 (N_21196,N_17595,N_19070);
xnor U21197 (N_21197,N_18966,N_19707);
or U21198 (N_21198,N_17967,N_19275);
nor U21199 (N_21199,N_19218,N_18847);
nor U21200 (N_21200,N_19397,N_18364);
nor U21201 (N_21201,N_19428,N_19886);
nor U21202 (N_21202,N_17696,N_17658);
xnor U21203 (N_21203,N_19523,N_18706);
nor U21204 (N_21204,N_18308,N_17789);
and U21205 (N_21205,N_18573,N_18608);
or U21206 (N_21206,N_19507,N_19850);
nand U21207 (N_21207,N_19026,N_19113);
nor U21208 (N_21208,N_17765,N_18086);
and U21209 (N_21209,N_19901,N_19948);
or U21210 (N_21210,N_17618,N_19002);
xor U21211 (N_21211,N_18233,N_18394);
or U21212 (N_21212,N_18421,N_19000);
nor U21213 (N_21213,N_19664,N_19479);
or U21214 (N_21214,N_18975,N_19556);
nor U21215 (N_21215,N_19599,N_19481);
nor U21216 (N_21216,N_19729,N_17929);
and U21217 (N_21217,N_18955,N_19020);
nor U21218 (N_21218,N_19990,N_18219);
or U21219 (N_21219,N_19907,N_18721);
nand U21220 (N_21220,N_19728,N_19194);
nand U21221 (N_21221,N_18319,N_17578);
nor U21222 (N_21222,N_18502,N_19068);
nor U21223 (N_21223,N_18089,N_19944);
nor U21224 (N_21224,N_18641,N_17779);
or U21225 (N_21225,N_19283,N_19086);
or U21226 (N_21226,N_18704,N_19866);
xnor U21227 (N_21227,N_17722,N_17581);
nand U21228 (N_21228,N_19499,N_18324);
or U21229 (N_21229,N_18802,N_18452);
and U21230 (N_21230,N_18593,N_19622);
xor U21231 (N_21231,N_19543,N_19982);
xnor U21232 (N_21232,N_19289,N_18853);
or U21233 (N_21233,N_19795,N_18808);
nor U21234 (N_21234,N_19823,N_19064);
or U21235 (N_21235,N_18349,N_18486);
nand U21236 (N_21236,N_18386,N_19521);
and U21237 (N_21237,N_17923,N_19801);
and U21238 (N_21238,N_19587,N_19843);
nand U21239 (N_21239,N_19410,N_18292);
nand U21240 (N_21240,N_19092,N_19745);
nor U21241 (N_21241,N_18464,N_17878);
xor U21242 (N_21242,N_19849,N_19828);
and U21243 (N_21243,N_17817,N_19966);
nor U21244 (N_21244,N_17781,N_19609);
nand U21245 (N_21245,N_19482,N_18436);
nand U21246 (N_21246,N_19830,N_18644);
nor U21247 (N_21247,N_17831,N_18432);
nor U21248 (N_21248,N_19222,N_19891);
and U21249 (N_21249,N_18772,N_18582);
and U21250 (N_21250,N_18915,N_19281);
or U21251 (N_21251,N_18394,N_18089);
nand U21252 (N_21252,N_17727,N_19142);
nand U21253 (N_21253,N_18497,N_17576);
nor U21254 (N_21254,N_19623,N_19070);
and U21255 (N_21255,N_17937,N_17910);
nand U21256 (N_21256,N_18977,N_19757);
nor U21257 (N_21257,N_17638,N_18893);
nor U21258 (N_21258,N_18789,N_19859);
or U21259 (N_21259,N_17863,N_18472);
or U21260 (N_21260,N_19010,N_19955);
or U21261 (N_21261,N_17980,N_18543);
nand U21262 (N_21262,N_19326,N_18006);
nor U21263 (N_21263,N_19275,N_19875);
nand U21264 (N_21264,N_19758,N_18074);
nand U21265 (N_21265,N_19304,N_17596);
or U21266 (N_21266,N_19045,N_17991);
nand U21267 (N_21267,N_18893,N_18520);
and U21268 (N_21268,N_18661,N_18719);
or U21269 (N_21269,N_19940,N_17853);
or U21270 (N_21270,N_19510,N_19345);
or U21271 (N_21271,N_18590,N_19458);
xnor U21272 (N_21272,N_18920,N_19550);
and U21273 (N_21273,N_19127,N_18181);
or U21274 (N_21274,N_19700,N_18232);
and U21275 (N_21275,N_18415,N_19512);
nand U21276 (N_21276,N_19553,N_19388);
nor U21277 (N_21277,N_19111,N_19250);
or U21278 (N_21278,N_18805,N_18198);
nand U21279 (N_21279,N_19596,N_19549);
and U21280 (N_21280,N_19211,N_18319);
or U21281 (N_21281,N_18150,N_18973);
or U21282 (N_21282,N_19868,N_19391);
nor U21283 (N_21283,N_19513,N_18983);
and U21284 (N_21284,N_18461,N_18956);
nor U21285 (N_21285,N_19010,N_19546);
xnor U21286 (N_21286,N_17901,N_19163);
xnor U21287 (N_21287,N_19659,N_19325);
or U21288 (N_21288,N_18227,N_17762);
nand U21289 (N_21289,N_18243,N_19314);
xor U21290 (N_21290,N_19880,N_18573);
nor U21291 (N_21291,N_19559,N_19323);
or U21292 (N_21292,N_19396,N_19530);
or U21293 (N_21293,N_18267,N_19295);
or U21294 (N_21294,N_19276,N_19302);
nand U21295 (N_21295,N_19408,N_18094);
nor U21296 (N_21296,N_17501,N_19907);
and U21297 (N_21297,N_18907,N_19991);
nand U21298 (N_21298,N_18905,N_19856);
and U21299 (N_21299,N_19427,N_18825);
and U21300 (N_21300,N_18975,N_17575);
and U21301 (N_21301,N_19868,N_17944);
and U21302 (N_21302,N_19026,N_18296);
and U21303 (N_21303,N_19237,N_19414);
nor U21304 (N_21304,N_18811,N_19904);
or U21305 (N_21305,N_19763,N_19334);
xnor U21306 (N_21306,N_18029,N_19391);
nand U21307 (N_21307,N_18731,N_19234);
nand U21308 (N_21308,N_19901,N_18053);
nor U21309 (N_21309,N_18537,N_19687);
and U21310 (N_21310,N_18852,N_19426);
and U21311 (N_21311,N_19209,N_17737);
and U21312 (N_21312,N_18969,N_19545);
nor U21313 (N_21313,N_18201,N_18025);
or U21314 (N_21314,N_19459,N_18151);
and U21315 (N_21315,N_19608,N_18845);
xnor U21316 (N_21316,N_19360,N_18533);
nand U21317 (N_21317,N_18525,N_18136);
or U21318 (N_21318,N_18188,N_19959);
or U21319 (N_21319,N_18897,N_17640);
and U21320 (N_21320,N_19980,N_19137);
nand U21321 (N_21321,N_19280,N_19532);
nor U21322 (N_21322,N_18066,N_18218);
or U21323 (N_21323,N_17981,N_19426);
or U21324 (N_21324,N_19166,N_19497);
nand U21325 (N_21325,N_19462,N_19962);
or U21326 (N_21326,N_17940,N_19138);
and U21327 (N_21327,N_18903,N_19064);
nor U21328 (N_21328,N_17528,N_19520);
nor U21329 (N_21329,N_18013,N_19669);
or U21330 (N_21330,N_19224,N_18278);
nand U21331 (N_21331,N_17641,N_18802);
or U21332 (N_21332,N_18601,N_17780);
nand U21333 (N_21333,N_19961,N_18011);
nor U21334 (N_21334,N_19654,N_19386);
nor U21335 (N_21335,N_18134,N_19345);
nor U21336 (N_21336,N_17503,N_19281);
nand U21337 (N_21337,N_18361,N_18282);
xor U21338 (N_21338,N_18682,N_18753);
or U21339 (N_21339,N_19151,N_19825);
nor U21340 (N_21340,N_17685,N_19814);
nor U21341 (N_21341,N_19298,N_18665);
xnor U21342 (N_21342,N_18189,N_19864);
xnor U21343 (N_21343,N_19939,N_18396);
or U21344 (N_21344,N_19772,N_18442);
and U21345 (N_21345,N_19975,N_19214);
nor U21346 (N_21346,N_19178,N_19737);
and U21347 (N_21347,N_19577,N_19704);
nand U21348 (N_21348,N_19033,N_19541);
nand U21349 (N_21349,N_19717,N_17641);
or U21350 (N_21350,N_19426,N_19831);
or U21351 (N_21351,N_17521,N_18221);
nor U21352 (N_21352,N_18756,N_19000);
nor U21353 (N_21353,N_19650,N_17754);
xor U21354 (N_21354,N_18782,N_18033);
and U21355 (N_21355,N_19033,N_17669);
or U21356 (N_21356,N_18856,N_19534);
or U21357 (N_21357,N_19830,N_18163);
or U21358 (N_21358,N_18354,N_17755);
nor U21359 (N_21359,N_17884,N_18367);
or U21360 (N_21360,N_19658,N_18689);
or U21361 (N_21361,N_17683,N_17559);
and U21362 (N_21362,N_17954,N_17590);
nor U21363 (N_21363,N_17617,N_17640);
or U21364 (N_21364,N_19026,N_18381);
or U21365 (N_21365,N_17592,N_19456);
or U21366 (N_21366,N_19222,N_19115);
nor U21367 (N_21367,N_18472,N_18434);
nor U21368 (N_21368,N_18561,N_19675);
and U21369 (N_21369,N_17526,N_18303);
and U21370 (N_21370,N_18198,N_19267);
and U21371 (N_21371,N_19839,N_19399);
or U21372 (N_21372,N_19259,N_19913);
nor U21373 (N_21373,N_19356,N_19102);
or U21374 (N_21374,N_18993,N_19189);
nand U21375 (N_21375,N_17708,N_19842);
or U21376 (N_21376,N_19335,N_17655);
nor U21377 (N_21377,N_18536,N_18210);
and U21378 (N_21378,N_17989,N_19555);
nand U21379 (N_21379,N_18441,N_19964);
or U21380 (N_21380,N_19053,N_17844);
and U21381 (N_21381,N_19534,N_18363);
and U21382 (N_21382,N_19837,N_18269);
nand U21383 (N_21383,N_19196,N_18117);
nor U21384 (N_21384,N_18892,N_19922);
nand U21385 (N_21385,N_18936,N_18492);
nor U21386 (N_21386,N_18934,N_19559);
xnor U21387 (N_21387,N_19065,N_19394);
nand U21388 (N_21388,N_18969,N_19470);
and U21389 (N_21389,N_19767,N_17592);
xor U21390 (N_21390,N_19518,N_19552);
and U21391 (N_21391,N_17843,N_18436);
nor U21392 (N_21392,N_19081,N_19627);
nor U21393 (N_21393,N_18134,N_17598);
nand U21394 (N_21394,N_19505,N_18108);
nand U21395 (N_21395,N_19125,N_19847);
nor U21396 (N_21396,N_17657,N_18970);
nor U21397 (N_21397,N_19159,N_19114);
and U21398 (N_21398,N_18996,N_18991);
nand U21399 (N_21399,N_19580,N_18137);
xor U21400 (N_21400,N_18057,N_19845);
xnor U21401 (N_21401,N_18820,N_18171);
nor U21402 (N_21402,N_19691,N_18604);
nor U21403 (N_21403,N_18328,N_18757);
and U21404 (N_21404,N_19739,N_18191);
and U21405 (N_21405,N_17737,N_18557);
or U21406 (N_21406,N_19322,N_19476);
or U21407 (N_21407,N_18772,N_19531);
nand U21408 (N_21408,N_18427,N_19832);
and U21409 (N_21409,N_17618,N_19216);
and U21410 (N_21410,N_17641,N_19924);
or U21411 (N_21411,N_18773,N_17851);
nor U21412 (N_21412,N_18337,N_17576);
or U21413 (N_21413,N_18778,N_19847);
or U21414 (N_21414,N_18450,N_17693);
nor U21415 (N_21415,N_17503,N_17738);
or U21416 (N_21416,N_19450,N_17642);
or U21417 (N_21417,N_17981,N_17929);
nor U21418 (N_21418,N_19618,N_18030);
nand U21419 (N_21419,N_18000,N_17515);
or U21420 (N_21420,N_17903,N_18940);
or U21421 (N_21421,N_19840,N_18697);
nand U21422 (N_21422,N_18674,N_19634);
or U21423 (N_21423,N_18766,N_17646);
nor U21424 (N_21424,N_18347,N_19311);
or U21425 (N_21425,N_19934,N_18575);
nand U21426 (N_21426,N_17837,N_18448);
and U21427 (N_21427,N_18571,N_18963);
nand U21428 (N_21428,N_18399,N_19515);
and U21429 (N_21429,N_19336,N_19414);
nor U21430 (N_21430,N_17736,N_17681);
or U21431 (N_21431,N_17573,N_17665);
nor U21432 (N_21432,N_17547,N_18393);
nor U21433 (N_21433,N_19505,N_19391);
and U21434 (N_21434,N_18888,N_17695);
nand U21435 (N_21435,N_19004,N_19746);
nand U21436 (N_21436,N_18939,N_17681);
nor U21437 (N_21437,N_18807,N_18910);
nor U21438 (N_21438,N_18910,N_17692);
nor U21439 (N_21439,N_19326,N_18611);
and U21440 (N_21440,N_17645,N_18668);
nand U21441 (N_21441,N_17813,N_19993);
nand U21442 (N_21442,N_18815,N_19392);
or U21443 (N_21443,N_19080,N_19047);
nor U21444 (N_21444,N_18369,N_18253);
nor U21445 (N_21445,N_19573,N_19014);
nor U21446 (N_21446,N_17567,N_17724);
and U21447 (N_21447,N_17645,N_18618);
and U21448 (N_21448,N_19701,N_17914);
or U21449 (N_21449,N_18361,N_18973);
or U21450 (N_21450,N_19509,N_19301);
and U21451 (N_21451,N_17691,N_18736);
xnor U21452 (N_21452,N_17846,N_18902);
or U21453 (N_21453,N_19096,N_19786);
nor U21454 (N_21454,N_18283,N_18744);
xor U21455 (N_21455,N_19652,N_19510);
nand U21456 (N_21456,N_19058,N_18790);
xor U21457 (N_21457,N_17999,N_19817);
and U21458 (N_21458,N_17955,N_18283);
xnor U21459 (N_21459,N_18228,N_19555);
and U21460 (N_21460,N_18553,N_19257);
nand U21461 (N_21461,N_18100,N_18578);
xnor U21462 (N_21462,N_19513,N_18729);
nor U21463 (N_21463,N_18587,N_17584);
nor U21464 (N_21464,N_17796,N_18414);
nand U21465 (N_21465,N_18884,N_18297);
nand U21466 (N_21466,N_18129,N_18347);
or U21467 (N_21467,N_18688,N_19268);
nand U21468 (N_21468,N_19411,N_17740);
and U21469 (N_21469,N_17626,N_19292);
and U21470 (N_21470,N_19729,N_19421);
xnor U21471 (N_21471,N_18066,N_18964);
nor U21472 (N_21472,N_19060,N_18284);
nor U21473 (N_21473,N_18618,N_19092);
xor U21474 (N_21474,N_19690,N_19116);
nand U21475 (N_21475,N_19956,N_19652);
or U21476 (N_21476,N_19191,N_18820);
or U21477 (N_21477,N_18386,N_19987);
nor U21478 (N_21478,N_18174,N_19922);
nor U21479 (N_21479,N_19632,N_18230);
nor U21480 (N_21480,N_18095,N_19401);
nor U21481 (N_21481,N_19044,N_18587);
nor U21482 (N_21482,N_18694,N_19928);
nor U21483 (N_21483,N_18156,N_18581);
nand U21484 (N_21484,N_19274,N_18284);
nand U21485 (N_21485,N_18587,N_19586);
nor U21486 (N_21486,N_18481,N_18313);
nor U21487 (N_21487,N_17514,N_18595);
nand U21488 (N_21488,N_18654,N_18879);
nand U21489 (N_21489,N_18715,N_19250);
xor U21490 (N_21490,N_19257,N_18067);
nor U21491 (N_21491,N_19353,N_17665);
or U21492 (N_21492,N_19975,N_19867);
and U21493 (N_21493,N_18525,N_18681);
and U21494 (N_21494,N_18457,N_19237);
nand U21495 (N_21495,N_17527,N_18353);
nand U21496 (N_21496,N_17611,N_19525);
xor U21497 (N_21497,N_18098,N_18960);
or U21498 (N_21498,N_18320,N_17683);
nor U21499 (N_21499,N_18848,N_19620);
nand U21500 (N_21500,N_17949,N_19106);
nor U21501 (N_21501,N_17594,N_19917);
nor U21502 (N_21502,N_18607,N_19780);
nor U21503 (N_21503,N_18749,N_19675);
nor U21504 (N_21504,N_18671,N_19774);
and U21505 (N_21505,N_17678,N_19109);
or U21506 (N_21506,N_18868,N_18391);
nor U21507 (N_21507,N_18154,N_19966);
nand U21508 (N_21508,N_18576,N_19069);
nor U21509 (N_21509,N_18368,N_18499);
nand U21510 (N_21510,N_17885,N_18605);
and U21511 (N_21511,N_18526,N_19627);
or U21512 (N_21512,N_19222,N_19973);
xnor U21513 (N_21513,N_17558,N_18531);
xnor U21514 (N_21514,N_19070,N_17509);
and U21515 (N_21515,N_18358,N_19060);
or U21516 (N_21516,N_17695,N_17767);
nor U21517 (N_21517,N_18577,N_19971);
and U21518 (N_21518,N_19430,N_17896);
nor U21519 (N_21519,N_19496,N_17511);
and U21520 (N_21520,N_18147,N_19766);
and U21521 (N_21521,N_18202,N_18421);
or U21522 (N_21522,N_18502,N_17575);
or U21523 (N_21523,N_19596,N_19302);
or U21524 (N_21524,N_19568,N_18625);
and U21525 (N_21525,N_19836,N_19093);
xor U21526 (N_21526,N_18628,N_18430);
or U21527 (N_21527,N_17901,N_18719);
nor U21528 (N_21528,N_18620,N_17566);
and U21529 (N_21529,N_17835,N_19839);
nor U21530 (N_21530,N_19317,N_18951);
and U21531 (N_21531,N_17708,N_18282);
nor U21532 (N_21532,N_19646,N_18539);
nand U21533 (N_21533,N_19135,N_19219);
nor U21534 (N_21534,N_17581,N_17733);
and U21535 (N_21535,N_18208,N_18693);
and U21536 (N_21536,N_18893,N_19844);
and U21537 (N_21537,N_19197,N_17681);
nand U21538 (N_21538,N_17510,N_18787);
nor U21539 (N_21539,N_17942,N_17917);
nand U21540 (N_21540,N_18268,N_17759);
or U21541 (N_21541,N_17517,N_18856);
xor U21542 (N_21542,N_17917,N_17710);
nor U21543 (N_21543,N_18047,N_18120);
nor U21544 (N_21544,N_18169,N_17752);
or U21545 (N_21545,N_19815,N_18486);
nor U21546 (N_21546,N_19105,N_19546);
and U21547 (N_21547,N_18448,N_17943);
and U21548 (N_21548,N_19139,N_19743);
and U21549 (N_21549,N_17571,N_17539);
nand U21550 (N_21550,N_18155,N_18492);
nor U21551 (N_21551,N_18196,N_18023);
and U21552 (N_21552,N_18570,N_18456);
nand U21553 (N_21553,N_19970,N_19834);
nor U21554 (N_21554,N_18150,N_19270);
and U21555 (N_21555,N_17782,N_19374);
or U21556 (N_21556,N_18279,N_17855);
nor U21557 (N_21557,N_18598,N_17606);
or U21558 (N_21558,N_17786,N_19285);
or U21559 (N_21559,N_18826,N_18799);
nand U21560 (N_21560,N_18875,N_19050);
and U21561 (N_21561,N_17944,N_17649);
nor U21562 (N_21562,N_18605,N_19095);
and U21563 (N_21563,N_18504,N_18434);
or U21564 (N_21564,N_19821,N_17614);
or U21565 (N_21565,N_17809,N_18783);
and U21566 (N_21566,N_18639,N_17705);
or U21567 (N_21567,N_19742,N_18039);
and U21568 (N_21568,N_18627,N_17925);
nand U21569 (N_21569,N_19056,N_19284);
and U21570 (N_21570,N_19694,N_19817);
nand U21571 (N_21571,N_18149,N_18074);
nor U21572 (N_21572,N_19782,N_19189);
or U21573 (N_21573,N_17792,N_19425);
or U21574 (N_21574,N_19199,N_18114);
xnor U21575 (N_21575,N_19317,N_18752);
nor U21576 (N_21576,N_17650,N_18892);
or U21577 (N_21577,N_17991,N_18615);
or U21578 (N_21578,N_19669,N_18174);
nor U21579 (N_21579,N_19750,N_19377);
or U21580 (N_21580,N_17809,N_19354);
or U21581 (N_21581,N_19470,N_18512);
and U21582 (N_21582,N_17944,N_19639);
and U21583 (N_21583,N_19748,N_19998);
nand U21584 (N_21584,N_17954,N_17512);
nand U21585 (N_21585,N_18093,N_18415);
and U21586 (N_21586,N_19259,N_19246);
nand U21587 (N_21587,N_18341,N_18214);
nand U21588 (N_21588,N_18590,N_18359);
xnor U21589 (N_21589,N_18175,N_18615);
or U21590 (N_21590,N_19266,N_17622);
nand U21591 (N_21591,N_19084,N_18934);
or U21592 (N_21592,N_18453,N_19444);
nor U21593 (N_21593,N_17564,N_18833);
and U21594 (N_21594,N_17892,N_19171);
and U21595 (N_21595,N_17896,N_17835);
nor U21596 (N_21596,N_18283,N_17583);
and U21597 (N_21597,N_17785,N_18261);
nor U21598 (N_21598,N_18299,N_19551);
nor U21599 (N_21599,N_19719,N_17527);
and U21600 (N_21600,N_18522,N_18245);
and U21601 (N_21601,N_19117,N_17914);
and U21602 (N_21602,N_18863,N_17970);
nor U21603 (N_21603,N_19004,N_18255);
nor U21604 (N_21604,N_17835,N_18725);
and U21605 (N_21605,N_19829,N_19615);
nand U21606 (N_21606,N_17787,N_17874);
nand U21607 (N_21607,N_19405,N_18347);
and U21608 (N_21608,N_18517,N_19158);
nor U21609 (N_21609,N_19765,N_19058);
nor U21610 (N_21610,N_18745,N_18411);
or U21611 (N_21611,N_18588,N_19546);
nor U21612 (N_21612,N_17956,N_18586);
nand U21613 (N_21613,N_19805,N_18249);
or U21614 (N_21614,N_17951,N_17786);
xor U21615 (N_21615,N_19409,N_19523);
nor U21616 (N_21616,N_17594,N_19849);
and U21617 (N_21617,N_18011,N_18009);
and U21618 (N_21618,N_18214,N_18486);
nor U21619 (N_21619,N_17806,N_19299);
nand U21620 (N_21620,N_19194,N_18829);
and U21621 (N_21621,N_18425,N_19366);
and U21622 (N_21622,N_18891,N_18241);
and U21623 (N_21623,N_18473,N_18624);
nor U21624 (N_21624,N_18731,N_18262);
or U21625 (N_21625,N_18958,N_19332);
nand U21626 (N_21626,N_18162,N_19524);
and U21627 (N_21627,N_19452,N_19016);
nand U21628 (N_21628,N_18148,N_19713);
and U21629 (N_21629,N_17685,N_17992);
and U21630 (N_21630,N_18559,N_19357);
nand U21631 (N_21631,N_18827,N_17616);
and U21632 (N_21632,N_18037,N_19874);
or U21633 (N_21633,N_18735,N_19026);
nor U21634 (N_21634,N_19543,N_18127);
nand U21635 (N_21635,N_19255,N_18092);
or U21636 (N_21636,N_19876,N_19757);
or U21637 (N_21637,N_18958,N_17904);
nand U21638 (N_21638,N_18460,N_19967);
nor U21639 (N_21639,N_17501,N_19395);
nand U21640 (N_21640,N_17616,N_19692);
and U21641 (N_21641,N_18382,N_17518);
or U21642 (N_21642,N_18895,N_17986);
nor U21643 (N_21643,N_19310,N_17536);
xnor U21644 (N_21644,N_19859,N_19991);
or U21645 (N_21645,N_18180,N_19354);
xor U21646 (N_21646,N_18064,N_17803);
or U21647 (N_21647,N_19079,N_17658);
nor U21648 (N_21648,N_17993,N_19750);
nand U21649 (N_21649,N_18388,N_18012);
xor U21650 (N_21650,N_19023,N_18920);
nand U21651 (N_21651,N_18014,N_18090);
xor U21652 (N_21652,N_19327,N_19234);
or U21653 (N_21653,N_19074,N_18441);
or U21654 (N_21654,N_18320,N_17707);
xor U21655 (N_21655,N_19162,N_18941);
or U21656 (N_21656,N_18528,N_18319);
and U21657 (N_21657,N_17852,N_18273);
nor U21658 (N_21658,N_17735,N_19111);
nor U21659 (N_21659,N_17781,N_18867);
nand U21660 (N_21660,N_19164,N_19604);
or U21661 (N_21661,N_17649,N_17518);
nor U21662 (N_21662,N_19042,N_18429);
xnor U21663 (N_21663,N_18091,N_19602);
or U21664 (N_21664,N_19984,N_18000);
xor U21665 (N_21665,N_18578,N_18910);
or U21666 (N_21666,N_18623,N_19829);
nand U21667 (N_21667,N_18283,N_17881);
nor U21668 (N_21668,N_19622,N_18660);
nand U21669 (N_21669,N_19946,N_18950);
nand U21670 (N_21670,N_19743,N_19044);
or U21671 (N_21671,N_17667,N_18321);
nor U21672 (N_21672,N_19898,N_18605);
nor U21673 (N_21673,N_18146,N_17905);
nand U21674 (N_21674,N_19822,N_19952);
nor U21675 (N_21675,N_18563,N_17695);
or U21676 (N_21676,N_19999,N_17579);
xnor U21677 (N_21677,N_19896,N_19489);
xnor U21678 (N_21678,N_18716,N_19433);
or U21679 (N_21679,N_18063,N_17831);
nand U21680 (N_21680,N_19408,N_19139);
and U21681 (N_21681,N_17968,N_18879);
or U21682 (N_21682,N_17805,N_18695);
xnor U21683 (N_21683,N_17663,N_18428);
xor U21684 (N_21684,N_18264,N_18047);
nor U21685 (N_21685,N_19112,N_19064);
nand U21686 (N_21686,N_17581,N_18551);
nor U21687 (N_21687,N_19293,N_19166);
and U21688 (N_21688,N_19965,N_18436);
nor U21689 (N_21689,N_18730,N_17923);
and U21690 (N_21690,N_19051,N_18005);
xnor U21691 (N_21691,N_19305,N_18784);
and U21692 (N_21692,N_19538,N_18912);
or U21693 (N_21693,N_19847,N_18348);
xnor U21694 (N_21694,N_18925,N_17500);
or U21695 (N_21695,N_19113,N_19684);
or U21696 (N_21696,N_19414,N_17830);
nor U21697 (N_21697,N_19482,N_18443);
nor U21698 (N_21698,N_17924,N_18480);
nand U21699 (N_21699,N_19068,N_19935);
nand U21700 (N_21700,N_18845,N_17981);
and U21701 (N_21701,N_17929,N_19069);
nand U21702 (N_21702,N_19278,N_19562);
or U21703 (N_21703,N_18571,N_19193);
and U21704 (N_21704,N_18650,N_18130);
nor U21705 (N_21705,N_18362,N_17608);
and U21706 (N_21706,N_17772,N_18969);
or U21707 (N_21707,N_19071,N_19552);
or U21708 (N_21708,N_19838,N_17910);
and U21709 (N_21709,N_18984,N_17990);
and U21710 (N_21710,N_19375,N_18034);
nor U21711 (N_21711,N_19925,N_18218);
and U21712 (N_21712,N_17581,N_17951);
xor U21713 (N_21713,N_17999,N_18200);
or U21714 (N_21714,N_19868,N_17539);
or U21715 (N_21715,N_19289,N_18868);
nand U21716 (N_21716,N_18670,N_18503);
nor U21717 (N_21717,N_18356,N_19238);
nor U21718 (N_21718,N_18567,N_17685);
and U21719 (N_21719,N_18316,N_19018);
nand U21720 (N_21720,N_19905,N_19912);
nand U21721 (N_21721,N_18700,N_19588);
nor U21722 (N_21722,N_19238,N_18102);
nand U21723 (N_21723,N_19130,N_18763);
or U21724 (N_21724,N_19619,N_19013);
nand U21725 (N_21725,N_18006,N_18715);
and U21726 (N_21726,N_17873,N_17933);
and U21727 (N_21727,N_18014,N_17915);
nor U21728 (N_21728,N_19262,N_17572);
nand U21729 (N_21729,N_19247,N_18854);
nand U21730 (N_21730,N_18301,N_19573);
and U21731 (N_21731,N_19004,N_18985);
nor U21732 (N_21732,N_19290,N_19407);
and U21733 (N_21733,N_19763,N_18159);
nor U21734 (N_21734,N_19078,N_17526);
nor U21735 (N_21735,N_17772,N_17853);
xnor U21736 (N_21736,N_18452,N_17885);
nand U21737 (N_21737,N_19050,N_18259);
nand U21738 (N_21738,N_19119,N_18445);
nor U21739 (N_21739,N_17642,N_18914);
xor U21740 (N_21740,N_18898,N_19958);
nand U21741 (N_21741,N_19227,N_18507);
and U21742 (N_21742,N_18761,N_17586);
nand U21743 (N_21743,N_19876,N_19587);
nor U21744 (N_21744,N_18962,N_17562);
and U21745 (N_21745,N_18557,N_18267);
nand U21746 (N_21746,N_18693,N_18099);
nor U21747 (N_21747,N_18585,N_19757);
nand U21748 (N_21748,N_19154,N_19920);
and U21749 (N_21749,N_19375,N_19648);
nor U21750 (N_21750,N_18129,N_19538);
nand U21751 (N_21751,N_19708,N_19228);
and U21752 (N_21752,N_19695,N_17937);
nor U21753 (N_21753,N_19429,N_18545);
nand U21754 (N_21754,N_17779,N_19643);
nand U21755 (N_21755,N_18012,N_17653);
nand U21756 (N_21756,N_18180,N_19982);
or U21757 (N_21757,N_19192,N_18357);
nand U21758 (N_21758,N_18709,N_19428);
or U21759 (N_21759,N_17520,N_18395);
xor U21760 (N_21760,N_19930,N_18147);
xnor U21761 (N_21761,N_18305,N_17727);
nand U21762 (N_21762,N_19861,N_18557);
nand U21763 (N_21763,N_18008,N_19978);
nand U21764 (N_21764,N_19143,N_18205);
xnor U21765 (N_21765,N_18978,N_18486);
nand U21766 (N_21766,N_19994,N_17811);
and U21767 (N_21767,N_19000,N_19508);
nand U21768 (N_21768,N_19387,N_19345);
nor U21769 (N_21769,N_19064,N_19947);
xor U21770 (N_21770,N_17766,N_18882);
and U21771 (N_21771,N_19076,N_19190);
and U21772 (N_21772,N_17572,N_17812);
xnor U21773 (N_21773,N_19606,N_19949);
nor U21774 (N_21774,N_19310,N_18910);
or U21775 (N_21775,N_18851,N_18687);
nand U21776 (N_21776,N_19278,N_19984);
or U21777 (N_21777,N_19550,N_18046);
nor U21778 (N_21778,N_18747,N_19896);
and U21779 (N_21779,N_19530,N_19423);
and U21780 (N_21780,N_18462,N_17861);
nand U21781 (N_21781,N_18692,N_19107);
nand U21782 (N_21782,N_19703,N_17940);
and U21783 (N_21783,N_17829,N_19482);
and U21784 (N_21784,N_17714,N_18035);
or U21785 (N_21785,N_17719,N_17732);
or U21786 (N_21786,N_18140,N_18124);
nand U21787 (N_21787,N_17949,N_19216);
nand U21788 (N_21788,N_18661,N_17582);
xnor U21789 (N_21789,N_19474,N_17845);
nor U21790 (N_21790,N_18352,N_17523);
and U21791 (N_21791,N_18937,N_18505);
xor U21792 (N_21792,N_18718,N_18483);
nand U21793 (N_21793,N_19377,N_18323);
nand U21794 (N_21794,N_18886,N_17883);
or U21795 (N_21795,N_17545,N_19235);
or U21796 (N_21796,N_19074,N_18750);
nor U21797 (N_21797,N_18741,N_18485);
or U21798 (N_21798,N_18223,N_18169);
xnor U21799 (N_21799,N_18615,N_17930);
or U21800 (N_21800,N_17522,N_19199);
xor U21801 (N_21801,N_17626,N_19829);
nor U21802 (N_21802,N_18524,N_19448);
nor U21803 (N_21803,N_18308,N_18435);
and U21804 (N_21804,N_17583,N_18783);
nand U21805 (N_21805,N_18695,N_17572);
xor U21806 (N_21806,N_17986,N_18433);
nand U21807 (N_21807,N_17648,N_18196);
nand U21808 (N_21808,N_18929,N_19119);
and U21809 (N_21809,N_18262,N_17550);
nand U21810 (N_21810,N_18281,N_17798);
xor U21811 (N_21811,N_18806,N_19984);
or U21812 (N_21812,N_18787,N_18580);
or U21813 (N_21813,N_19400,N_17650);
or U21814 (N_21814,N_17828,N_19868);
nor U21815 (N_21815,N_17960,N_18453);
nand U21816 (N_21816,N_19118,N_18537);
and U21817 (N_21817,N_17582,N_18735);
nand U21818 (N_21818,N_18619,N_18112);
and U21819 (N_21819,N_19948,N_19302);
nand U21820 (N_21820,N_18362,N_17712);
nor U21821 (N_21821,N_18760,N_19142);
or U21822 (N_21822,N_19915,N_18495);
nor U21823 (N_21823,N_18791,N_19317);
or U21824 (N_21824,N_18589,N_19658);
and U21825 (N_21825,N_19132,N_18478);
or U21826 (N_21826,N_18224,N_17785);
and U21827 (N_21827,N_18575,N_17568);
or U21828 (N_21828,N_19891,N_18654);
or U21829 (N_21829,N_17683,N_18852);
nor U21830 (N_21830,N_18682,N_19845);
xnor U21831 (N_21831,N_17870,N_18937);
or U21832 (N_21832,N_18287,N_18429);
nand U21833 (N_21833,N_18585,N_17764);
xor U21834 (N_21834,N_19377,N_17999);
or U21835 (N_21835,N_17705,N_17840);
nand U21836 (N_21836,N_17974,N_19876);
nand U21837 (N_21837,N_18638,N_18168);
nor U21838 (N_21838,N_17946,N_17888);
xor U21839 (N_21839,N_19741,N_19997);
nor U21840 (N_21840,N_17698,N_18283);
and U21841 (N_21841,N_17536,N_19977);
or U21842 (N_21842,N_18644,N_17856);
and U21843 (N_21843,N_18701,N_18230);
and U21844 (N_21844,N_17736,N_18821);
and U21845 (N_21845,N_19439,N_17590);
nand U21846 (N_21846,N_19747,N_19161);
or U21847 (N_21847,N_18660,N_19288);
or U21848 (N_21848,N_19788,N_18861);
nor U21849 (N_21849,N_19202,N_17831);
xor U21850 (N_21850,N_18457,N_17526);
and U21851 (N_21851,N_18565,N_18218);
or U21852 (N_21852,N_19924,N_19102);
nor U21853 (N_21853,N_19673,N_19080);
nand U21854 (N_21854,N_19551,N_17927);
or U21855 (N_21855,N_18795,N_19130);
and U21856 (N_21856,N_19751,N_17777);
nand U21857 (N_21857,N_18021,N_18953);
nand U21858 (N_21858,N_18733,N_18955);
nand U21859 (N_21859,N_18984,N_18166);
nor U21860 (N_21860,N_17790,N_18570);
xor U21861 (N_21861,N_19859,N_18514);
xnor U21862 (N_21862,N_18710,N_17779);
xor U21863 (N_21863,N_18948,N_18527);
nor U21864 (N_21864,N_17564,N_17579);
nor U21865 (N_21865,N_19874,N_18639);
and U21866 (N_21866,N_18232,N_19650);
and U21867 (N_21867,N_18228,N_19696);
xor U21868 (N_21868,N_18893,N_18710);
xor U21869 (N_21869,N_19746,N_18220);
nor U21870 (N_21870,N_18514,N_18352);
nor U21871 (N_21871,N_18913,N_19898);
and U21872 (N_21872,N_19440,N_19829);
xnor U21873 (N_21873,N_18780,N_19270);
or U21874 (N_21874,N_17940,N_19781);
and U21875 (N_21875,N_18779,N_19104);
or U21876 (N_21876,N_18303,N_19926);
nand U21877 (N_21877,N_18817,N_18656);
nor U21878 (N_21878,N_19921,N_18475);
nand U21879 (N_21879,N_17999,N_18706);
nor U21880 (N_21880,N_18532,N_18077);
and U21881 (N_21881,N_19606,N_19127);
and U21882 (N_21882,N_19169,N_17573);
nor U21883 (N_21883,N_19018,N_19074);
nand U21884 (N_21884,N_17516,N_19262);
xor U21885 (N_21885,N_18633,N_19488);
nor U21886 (N_21886,N_18330,N_18649);
or U21887 (N_21887,N_18453,N_18810);
nand U21888 (N_21888,N_18486,N_17789);
nand U21889 (N_21889,N_17543,N_18603);
nand U21890 (N_21890,N_19043,N_19416);
nand U21891 (N_21891,N_17892,N_18042);
nor U21892 (N_21892,N_18979,N_19591);
and U21893 (N_21893,N_17544,N_18334);
nor U21894 (N_21894,N_19933,N_18780);
or U21895 (N_21895,N_18624,N_17865);
or U21896 (N_21896,N_19410,N_18894);
nor U21897 (N_21897,N_19413,N_18334);
nand U21898 (N_21898,N_18773,N_19698);
nand U21899 (N_21899,N_17955,N_17591);
nand U21900 (N_21900,N_18073,N_17827);
nand U21901 (N_21901,N_18671,N_19020);
or U21902 (N_21902,N_19927,N_17597);
or U21903 (N_21903,N_17520,N_19067);
xor U21904 (N_21904,N_18433,N_17915);
or U21905 (N_21905,N_18192,N_18872);
and U21906 (N_21906,N_18108,N_19613);
nand U21907 (N_21907,N_18399,N_18682);
nand U21908 (N_21908,N_18429,N_17863);
and U21909 (N_21909,N_19957,N_18043);
xnor U21910 (N_21910,N_19513,N_18986);
and U21911 (N_21911,N_19020,N_17799);
or U21912 (N_21912,N_19691,N_18929);
xnor U21913 (N_21913,N_19490,N_17754);
xnor U21914 (N_21914,N_18927,N_17708);
nor U21915 (N_21915,N_17772,N_17625);
or U21916 (N_21916,N_18278,N_18388);
or U21917 (N_21917,N_17557,N_18406);
nand U21918 (N_21918,N_18249,N_19609);
nand U21919 (N_21919,N_19046,N_17620);
nor U21920 (N_21920,N_19119,N_19749);
and U21921 (N_21921,N_18096,N_17559);
and U21922 (N_21922,N_18267,N_19721);
and U21923 (N_21923,N_19875,N_17753);
and U21924 (N_21924,N_19155,N_18882);
xnor U21925 (N_21925,N_18852,N_19843);
or U21926 (N_21926,N_18463,N_17681);
nand U21927 (N_21927,N_18752,N_19821);
nand U21928 (N_21928,N_19164,N_19718);
xor U21929 (N_21929,N_19325,N_19821);
xor U21930 (N_21930,N_18095,N_19233);
or U21931 (N_21931,N_18350,N_19064);
nor U21932 (N_21932,N_18279,N_17911);
nand U21933 (N_21933,N_17561,N_19050);
nand U21934 (N_21934,N_19351,N_18696);
and U21935 (N_21935,N_18050,N_18093);
nand U21936 (N_21936,N_18162,N_19280);
nor U21937 (N_21937,N_18333,N_18144);
and U21938 (N_21938,N_19956,N_19258);
nor U21939 (N_21939,N_18401,N_19924);
nand U21940 (N_21940,N_18080,N_18140);
and U21941 (N_21941,N_18634,N_18300);
or U21942 (N_21942,N_18034,N_19499);
nor U21943 (N_21943,N_18188,N_19403);
or U21944 (N_21944,N_18171,N_18383);
or U21945 (N_21945,N_19334,N_19045);
and U21946 (N_21946,N_18539,N_17833);
nand U21947 (N_21947,N_19023,N_18972);
or U21948 (N_21948,N_18891,N_18212);
and U21949 (N_21949,N_19538,N_18725);
and U21950 (N_21950,N_18290,N_17569);
xnor U21951 (N_21951,N_18762,N_19750);
xnor U21952 (N_21952,N_18725,N_17682);
nor U21953 (N_21953,N_19087,N_18330);
or U21954 (N_21954,N_18742,N_19390);
and U21955 (N_21955,N_17837,N_19331);
and U21956 (N_21956,N_18239,N_19387);
and U21957 (N_21957,N_18088,N_19247);
nand U21958 (N_21958,N_18889,N_18208);
nor U21959 (N_21959,N_18483,N_18171);
and U21960 (N_21960,N_18935,N_18286);
nor U21961 (N_21961,N_17889,N_18203);
nor U21962 (N_21962,N_18713,N_18384);
nor U21963 (N_21963,N_18080,N_19260);
or U21964 (N_21964,N_17585,N_19649);
nand U21965 (N_21965,N_18499,N_18647);
and U21966 (N_21966,N_18474,N_17557);
or U21967 (N_21967,N_18284,N_18510);
nand U21968 (N_21968,N_18583,N_19458);
nor U21969 (N_21969,N_19955,N_19343);
and U21970 (N_21970,N_19021,N_19974);
xor U21971 (N_21971,N_19086,N_18785);
or U21972 (N_21972,N_18395,N_18439);
nor U21973 (N_21973,N_18852,N_18300);
and U21974 (N_21974,N_19695,N_17917);
and U21975 (N_21975,N_17920,N_17593);
nor U21976 (N_21976,N_17776,N_18727);
nand U21977 (N_21977,N_17793,N_18329);
and U21978 (N_21978,N_19113,N_18306);
and U21979 (N_21979,N_17939,N_19183);
or U21980 (N_21980,N_17659,N_19100);
nand U21981 (N_21981,N_19648,N_18129);
and U21982 (N_21982,N_19598,N_19519);
nor U21983 (N_21983,N_18148,N_19735);
nand U21984 (N_21984,N_17901,N_18034);
and U21985 (N_21985,N_19477,N_18889);
nor U21986 (N_21986,N_19651,N_19219);
and U21987 (N_21987,N_19375,N_18685);
nor U21988 (N_21988,N_19994,N_19830);
nor U21989 (N_21989,N_18284,N_18015);
nor U21990 (N_21990,N_17656,N_18181);
xor U21991 (N_21991,N_19177,N_17750);
xnor U21992 (N_21992,N_17835,N_18851);
nor U21993 (N_21993,N_17983,N_19959);
nand U21994 (N_21994,N_18763,N_19292);
xnor U21995 (N_21995,N_17518,N_19122);
and U21996 (N_21996,N_18259,N_19318);
and U21997 (N_21997,N_17948,N_19312);
or U21998 (N_21998,N_17924,N_19474);
nand U21999 (N_21999,N_18146,N_19691);
nand U22000 (N_22000,N_18589,N_18953);
nor U22001 (N_22001,N_18492,N_18635);
xor U22002 (N_22002,N_17718,N_18015);
xnor U22003 (N_22003,N_19807,N_18030);
nor U22004 (N_22004,N_18151,N_19062);
xnor U22005 (N_22005,N_19467,N_19082);
nand U22006 (N_22006,N_17851,N_18176);
nand U22007 (N_22007,N_18780,N_18493);
or U22008 (N_22008,N_18439,N_19765);
nor U22009 (N_22009,N_18375,N_18215);
nor U22010 (N_22010,N_19687,N_17932);
nor U22011 (N_22011,N_19605,N_19400);
and U22012 (N_22012,N_19083,N_18118);
or U22013 (N_22013,N_19076,N_17586);
nor U22014 (N_22014,N_19811,N_18546);
nand U22015 (N_22015,N_18068,N_18688);
nand U22016 (N_22016,N_18158,N_18170);
and U22017 (N_22017,N_19667,N_18749);
nor U22018 (N_22018,N_19006,N_19905);
xor U22019 (N_22019,N_19699,N_19786);
nand U22020 (N_22020,N_18711,N_18638);
or U22021 (N_22021,N_17983,N_18625);
and U22022 (N_22022,N_18622,N_19523);
or U22023 (N_22023,N_19837,N_18578);
nand U22024 (N_22024,N_18161,N_17607);
nand U22025 (N_22025,N_17790,N_18755);
and U22026 (N_22026,N_17929,N_18997);
nor U22027 (N_22027,N_18525,N_19310);
xnor U22028 (N_22028,N_19060,N_19475);
and U22029 (N_22029,N_18164,N_18777);
xnor U22030 (N_22030,N_19578,N_18181);
nand U22031 (N_22031,N_19407,N_19307);
nand U22032 (N_22032,N_17666,N_18753);
nand U22033 (N_22033,N_17845,N_18012);
nor U22034 (N_22034,N_19794,N_19934);
and U22035 (N_22035,N_19813,N_17754);
nor U22036 (N_22036,N_18276,N_18136);
nor U22037 (N_22037,N_17915,N_17942);
xnor U22038 (N_22038,N_17816,N_18360);
nand U22039 (N_22039,N_18045,N_19465);
nand U22040 (N_22040,N_18437,N_17947);
and U22041 (N_22041,N_18657,N_17758);
and U22042 (N_22042,N_18308,N_18160);
xor U22043 (N_22043,N_19640,N_18365);
and U22044 (N_22044,N_18388,N_19757);
or U22045 (N_22045,N_18590,N_19765);
nand U22046 (N_22046,N_19447,N_18434);
nor U22047 (N_22047,N_19709,N_17551);
nor U22048 (N_22048,N_19286,N_18056);
nor U22049 (N_22049,N_18175,N_18605);
or U22050 (N_22050,N_19634,N_18291);
and U22051 (N_22051,N_17934,N_19332);
nor U22052 (N_22052,N_17595,N_18502);
nand U22053 (N_22053,N_17736,N_17827);
nand U22054 (N_22054,N_19749,N_19011);
nor U22055 (N_22055,N_19467,N_19377);
nor U22056 (N_22056,N_19900,N_19624);
nor U22057 (N_22057,N_19791,N_17566);
nor U22058 (N_22058,N_18090,N_19396);
xor U22059 (N_22059,N_17620,N_18437);
nor U22060 (N_22060,N_19543,N_19493);
nand U22061 (N_22061,N_18304,N_18288);
or U22062 (N_22062,N_18412,N_19210);
nand U22063 (N_22063,N_18934,N_18690);
or U22064 (N_22064,N_18593,N_18621);
nand U22065 (N_22065,N_18254,N_18672);
xor U22066 (N_22066,N_18272,N_19480);
and U22067 (N_22067,N_19833,N_18332);
xor U22068 (N_22068,N_18202,N_17865);
xor U22069 (N_22069,N_17556,N_17932);
or U22070 (N_22070,N_18112,N_17914);
or U22071 (N_22071,N_18655,N_18387);
nand U22072 (N_22072,N_19960,N_19674);
or U22073 (N_22073,N_18627,N_18922);
xnor U22074 (N_22074,N_19150,N_19762);
or U22075 (N_22075,N_19975,N_19804);
nand U22076 (N_22076,N_19630,N_19253);
or U22077 (N_22077,N_19891,N_18728);
nand U22078 (N_22078,N_17740,N_19473);
or U22079 (N_22079,N_18878,N_18153);
nand U22080 (N_22080,N_17985,N_18832);
or U22081 (N_22081,N_18592,N_17837);
xnor U22082 (N_22082,N_17947,N_18793);
and U22083 (N_22083,N_17636,N_18892);
nand U22084 (N_22084,N_19272,N_18284);
xnor U22085 (N_22085,N_19204,N_18398);
nand U22086 (N_22086,N_19693,N_19970);
nor U22087 (N_22087,N_17717,N_18138);
or U22088 (N_22088,N_18032,N_18300);
xor U22089 (N_22089,N_18100,N_18119);
nor U22090 (N_22090,N_18797,N_19866);
nand U22091 (N_22091,N_19183,N_19474);
xnor U22092 (N_22092,N_19586,N_19464);
nor U22093 (N_22093,N_17665,N_17817);
nor U22094 (N_22094,N_18667,N_18066);
or U22095 (N_22095,N_19187,N_19287);
and U22096 (N_22096,N_19747,N_18623);
and U22097 (N_22097,N_17928,N_19382);
or U22098 (N_22098,N_17998,N_18186);
xor U22099 (N_22099,N_18231,N_18259);
xor U22100 (N_22100,N_18352,N_19668);
nand U22101 (N_22101,N_18823,N_18590);
and U22102 (N_22102,N_18866,N_18334);
or U22103 (N_22103,N_17556,N_17637);
nor U22104 (N_22104,N_19887,N_18371);
and U22105 (N_22105,N_17930,N_19971);
or U22106 (N_22106,N_18123,N_18579);
nor U22107 (N_22107,N_18308,N_18830);
xor U22108 (N_22108,N_19182,N_18429);
nor U22109 (N_22109,N_19770,N_19284);
nand U22110 (N_22110,N_17807,N_18136);
and U22111 (N_22111,N_18210,N_18589);
or U22112 (N_22112,N_19598,N_18258);
nor U22113 (N_22113,N_17501,N_18968);
and U22114 (N_22114,N_17878,N_18432);
nand U22115 (N_22115,N_19162,N_18960);
xor U22116 (N_22116,N_19312,N_18954);
nor U22117 (N_22117,N_18043,N_18750);
and U22118 (N_22118,N_17568,N_19632);
nor U22119 (N_22119,N_18836,N_19816);
or U22120 (N_22120,N_19994,N_18299);
and U22121 (N_22121,N_18420,N_18036);
nor U22122 (N_22122,N_18197,N_19119);
and U22123 (N_22123,N_19588,N_18210);
or U22124 (N_22124,N_18997,N_19980);
nand U22125 (N_22125,N_17646,N_17981);
or U22126 (N_22126,N_17780,N_19873);
and U22127 (N_22127,N_17981,N_18589);
xor U22128 (N_22128,N_19237,N_18377);
nor U22129 (N_22129,N_19900,N_17601);
nand U22130 (N_22130,N_18215,N_18412);
nor U22131 (N_22131,N_17828,N_17957);
nand U22132 (N_22132,N_18468,N_17749);
nor U22133 (N_22133,N_19200,N_18177);
nand U22134 (N_22134,N_18928,N_18057);
nand U22135 (N_22135,N_18442,N_18934);
and U22136 (N_22136,N_19093,N_18686);
nor U22137 (N_22137,N_18012,N_18264);
nor U22138 (N_22138,N_18465,N_18663);
or U22139 (N_22139,N_17519,N_17608);
and U22140 (N_22140,N_18382,N_18326);
nand U22141 (N_22141,N_19315,N_18474);
and U22142 (N_22142,N_17813,N_19270);
nand U22143 (N_22143,N_19318,N_19107);
nand U22144 (N_22144,N_19513,N_17618);
nor U22145 (N_22145,N_18782,N_18358);
nor U22146 (N_22146,N_18001,N_18301);
and U22147 (N_22147,N_18735,N_19808);
xnor U22148 (N_22148,N_19984,N_18409);
and U22149 (N_22149,N_18129,N_19375);
nor U22150 (N_22150,N_17952,N_17841);
nand U22151 (N_22151,N_17693,N_18556);
xnor U22152 (N_22152,N_19843,N_19355);
and U22153 (N_22153,N_17548,N_19765);
or U22154 (N_22154,N_18595,N_18665);
and U22155 (N_22155,N_18439,N_19351);
nor U22156 (N_22156,N_19491,N_18879);
and U22157 (N_22157,N_19637,N_19755);
or U22158 (N_22158,N_18504,N_17689);
and U22159 (N_22159,N_19880,N_19928);
and U22160 (N_22160,N_19655,N_17928);
or U22161 (N_22161,N_19180,N_17918);
xor U22162 (N_22162,N_19433,N_18663);
and U22163 (N_22163,N_18269,N_18181);
xnor U22164 (N_22164,N_17850,N_18320);
and U22165 (N_22165,N_19383,N_17790);
nor U22166 (N_22166,N_19132,N_18742);
nand U22167 (N_22167,N_17541,N_19811);
nand U22168 (N_22168,N_17528,N_17944);
or U22169 (N_22169,N_18339,N_18029);
nand U22170 (N_22170,N_18484,N_19673);
and U22171 (N_22171,N_17701,N_19845);
and U22172 (N_22172,N_18890,N_18447);
and U22173 (N_22173,N_19909,N_19953);
xor U22174 (N_22174,N_19071,N_19917);
and U22175 (N_22175,N_17760,N_19121);
nand U22176 (N_22176,N_19174,N_17798);
xnor U22177 (N_22177,N_19796,N_18216);
nand U22178 (N_22178,N_18837,N_19645);
and U22179 (N_22179,N_19499,N_18505);
or U22180 (N_22180,N_17526,N_18239);
nor U22181 (N_22181,N_19709,N_18008);
xor U22182 (N_22182,N_19232,N_19351);
nor U22183 (N_22183,N_18345,N_18016);
nor U22184 (N_22184,N_18927,N_18779);
and U22185 (N_22185,N_18936,N_17854);
and U22186 (N_22186,N_17500,N_19948);
or U22187 (N_22187,N_18678,N_17945);
xnor U22188 (N_22188,N_18138,N_18876);
or U22189 (N_22189,N_18383,N_18617);
nor U22190 (N_22190,N_18477,N_17933);
or U22191 (N_22191,N_19993,N_19590);
and U22192 (N_22192,N_19998,N_19855);
or U22193 (N_22193,N_19987,N_18943);
or U22194 (N_22194,N_19571,N_19793);
and U22195 (N_22195,N_17750,N_17730);
xnor U22196 (N_22196,N_19307,N_18424);
and U22197 (N_22197,N_18183,N_18842);
and U22198 (N_22198,N_17827,N_19330);
and U22199 (N_22199,N_17502,N_19716);
xor U22200 (N_22200,N_17904,N_19207);
nand U22201 (N_22201,N_17643,N_19850);
or U22202 (N_22202,N_18329,N_19523);
or U22203 (N_22203,N_19110,N_17573);
or U22204 (N_22204,N_18690,N_19348);
and U22205 (N_22205,N_17583,N_19599);
nand U22206 (N_22206,N_19421,N_19225);
or U22207 (N_22207,N_19782,N_19990);
and U22208 (N_22208,N_18652,N_17518);
or U22209 (N_22209,N_19282,N_18387);
and U22210 (N_22210,N_19919,N_18694);
nor U22211 (N_22211,N_19605,N_17568);
or U22212 (N_22212,N_19646,N_19320);
nor U22213 (N_22213,N_19257,N_18097);
or U22214 (N_22214,N_19302,N_19184);
nor U22215 (N_22215,N_18585,N_17927);
or U22216 (N_22216,N_18109,N_17820);
xor U22217 (N_22217,N_18002,N_18285);
nor U22218 (N_22218,N_17846,N_18284);
or U22219 (N_22219,N_18213,N_19068);
nor U22220 (N_22220,N_18982,N_19925);
nor U22221 (N_22221,N_18068,N_18058);
or U22222 (N_22222,N_19976,N_19287);
and U22223 (N_22223,N_18087,N_17823);
nor U22224 (N_22224,N_18674,N_18333);
and U22225 (N_22225,N_18046,N_19839);
xnor U22226 (N_22226,N_18189,N_19152);
nor U22227 (N_22227,N_17767,N_19427);
nor U22228 (N_22228,N_19699,N_18801);
xnor U22229 (N_22229,N_19108,N_18773);
nand U22230 (N_22230,N_19009,N_18612);
and U22231 (N_22231,N_19481,N_19419);
and U22232 (N_22232,N_19294,N_19774);
nand U22233 (N_22233,N_18244,N_19984);
nand U22234 (N_22234,N_17659,N_18443);
nand U22235 (N_22235,N_17732,N_19853);
xnor U22236 (N_22236,N_17805,N_19491);
or U22237 (N_22237,N_19477,N_19620);
xor U22238 (N_22238,N_17522,N_18719);
and U22239 (N_22239,N_18462,N_19822);
xnor U22240 (N_22240,N_19739,N_18162);
and U22241 (N_22241,N_19054,N_18597);
or U22242 (N_22242,N_17528,N_19480);
and U22243 (N_22243,N_19331,N_18272);
xnor U22244 (N_22244,N_18010,N_18221);
nor U22245 (N_22245,N_19942,N_17854);
nand U22246 (N_22246,N_19579,N_19643);
and U22247 (N_22247,N_19217,N_19001);
nor U22248 (N_22248,N_18560,N_18445);
nor U22249 (N_22249,N_19034,N_17679);
and U22250 (N_22250,N_19798,N_18325);
and U22251 (N_22251,N_18105,N_18521);
or U22252 (N_22252,N_18479,N_17710);
xnor U22253 (N_22253,N_18685,N_18298);
and U22254 (N_22254,N_19867,N_19620);
or U22255 (N_22255,N_18594,N_18233);
and U22256 (N_22256,N_17655,N_19576);
nor U22257 (N_22257,N_18332,N_19187);
nand U22258 (N_22258,N_18632,N_18169);
and U22259 (N_22259,N_17525,N_18742);
and U22260 (N_22260,N_18067,N_18118);
nand U22261 (N_22261,N_18054,N_18806);
and U22262 (N_22262,N_18044,N_18569);
nand U22263 (N_22263,N_17739,N_19353);
or U22264 (N_22264,N_17951,N_19157);
nor U22265 (N_22265,N_19486,N_17736);
nor U22266 (N_22266,N_18387,N_18852);
nand U22267 (N_22267,N_18999,N_18374);
or U22268 (N_22268,N_19621,N_19412);
nand U22269 (N_22269,N_18687,N_19427);
xor U22270 (N_22270,N_18434,N_19309);
nor U22271 (N_22271,N_19190,N_19172);
nand U22272 (N_22272,N_19493,N_18749);
and U22273 (N_22273,N_17691,N_19469);
or U22274 (N_22274,N_18930,N_18486);
or U22275 (N_22275,N_19837,N_18847);
nor U22276 (N_22276,N_18554,N_19312);
nor U22277 (N_22277,N_19907,N_18208);
and U22278 (N_22278,N_17676,N_19545);
and U22279 (N_22279,N_18671,N_17836);
and U22280 (N_22280,N_18467,N_17597);
nand U22281 (N_22281,N_18474,N_18967);
nor U22282 (N_22282,N_19131,N_19498);
and U22283 (N_22283,N_19909,N_19282);
xnor U22284 (N_22284,N_17541,N_19869);
nand U22285 (N_22285,N_18618,N_19740);
and U22286 (N_22286,N_18027,N_19699);
or U22287 (N_22287,N_19310,N_17584);
nand U22288 (N_22288,N_19621,N_19417);
and U22289 (N_22289,N_17881,N_18799);
or U22290 (N_22290,N_19733,N_18462);
nand U22291 (N_22291,N_17778,N_19766);
and U22292 (N_22292,N_19199,N_18594);
xnor U22293 (N_22293,N_19804,N_18492);
or U22294 (N_22294,N_19582,N_17801);
and U22295 (N_22295,N_18139,N_17812);
and U22296 (N_22296,N_19717,N_19366);
xnor U22297 (N_22297,N_19571,N_17982);
nand U22298 (N_22298,N_19577,N_19980);
nand U22299 (N_22299,N_19030,N_18855);
nor U22300 (N_22300,N_18584,N_18055);
xor U22301 (N_22301,N_18503,N_19910);
xor U22302 (N_22302,N_18556,N_18726);
nand U22303 (N_22303,N_18755,N_19517);
xnor U22304 (N_22304,N_19325,N_17608);
and U22305 (N_22305,N_19115,N_19116);
and U22306 (N_22306,N_19672,N_18781);
nand U22307 (N_22307,N_18625,N_19663);
and U22308 (N_22308,N_17923,N_19802);
or U22309 (N_22309,N_18149,N_18030);
and U22310 (N_22310,N_17874,N_19409);
xor U22311 (N_22311,N_19808,N_17845);
xor U22312 (N_22312,N_18911,N_18195);
xor U22313 (N_22313,N_18815,N_19012);
or U22314 (N_22314,N_19193,N_18144);
nand U22315 (N_22315,N_18920,N_17756);
nand U22316 (N_22316,N_17909,N_17583);
and U22317 (N_22317,N_19307,N_19460);
and U22318 (N_22318,N_18708,N_18602);
nor U22319 (N_22319,N_19553,N_18876);
and U22320 (N_22320,N_19995,N_18236);
or U22321 (N_22321,N_18995,N_19384);
nor U22322 (N_22322,N_19979,N_18487);
nor U22323 (N_22323,N_18878,N_17987);
nand U22324 (N_22324,N_19163,N_19642);
and U22325 (N_22325,N_19509,N_17793);
or U22326 (N_22326,N_19687,N_19206);
nand U22327 (N_22327,N_19421,N_18784);
nor U22328 (N_22328,N_19615,N_17747);
and U22329 (N_22329,N_18648,N_19423);
nor U22330 (N_22330,N_18673,N_18635);
nor U22331 (N_22331,N_19610,N_19437);
nand U22332 (N_22332,N_17856,N_17702);
nand U22333 (N_22333,N_18384,N_19439);
and U22334 (N_22334,N_18897,N_19151);
or U22335 (N_22335,N_18197,N_17865);
or U22336 (N_22336,N_18838,N_17588);
nor U22337 (N_22337,N_18808,N_19413);
nor U22338 (N_22338,N_19650,N_17975);
or U22339 (N_22339,N_19221,N_19616);
nor U22340 (N_22340,N_19149,N_19132);
nand U22341 (N_22341,N_19005,N_19906);
and U22342 (N_22342,N_18939,N_19830);
and U22343 (N_22343,N_17619,N_19502);
nand U22344 (N_22344,N_19940,N_18583);
or U22345 (N_22345,N_18993,N_18771);
xnor U22346 (N_22346,N_17844,N_18225);
or U22347 (N_22347,N_18279,N_19295);
nor U22348 (N_22348,N_18035,N_19760);
nor U22349 (N_22349,N_19895,N_18606);
and U22350 (N_22350,N_18530,N_17627);
nor U22351 (N_22351,N_17788,N_18976);
nor U22352 (N_22352,N_19619,N_18177);
nand U22353 (N_22353,N_18935,N_17581);
or U22354 (N_22354,N_19774,N_19182);
or U22355 (N_22355,N_17852,N_17799);
xnor U22356 (N_22356,N_18357,N_19069);
or U22357 (N_22357,N_19016,N_19460);
or U22358 (N_22358,N_19946,N_18220);
nor U22359 (N_22359,N_18861,N_18671);
nor U22360 (N_22360,N_18777,N_18094);
nor U22361 (N_22361,N_17947,N_19450);
nor U22362 (N_22362,N_19430,N_18623);
or U22363 (N_22363,N_19548,N_18595);
nor U22364 (N_22364,N_17850,N_18851);
nor U22365 (N_22365,N_18876,N_18096);
nand U22366 (N_22366,N_18638,N_18586);
xnor U22367 (N_22367,N_19146,N_17823);
nand U22368 (N_22368,N_17959,N_19741);
and U22369 (N_22369,N_17519,N_19565);
and U22370 (N_22370,N_19880,N_18112);
nor U22371 (N_22371,N_18220,N_18368);
nor U22372 (N_22372,N_19726,N_18670);
xor U22373 (N_22373,N_19081,N_19748);
nand U22374 (N_22374,N_18271,N_19110);
and U22375 (N_22375,N_19825,N_19424);
nand U22376 (N_22376,N_19993,N_19669);
nand U22377 (N_22377,N_19468,N_19494);
nor U22378 (N_22378,N_17859,N_18923);
nand U22379 (N_22379,N_18099,N_19675);
nor U22380 (N_22380,N_18997,N_17809);
or U22381 (N_22381,N_18684,N_18034);
nor U22382 (N_22382,N_19307,N_19105);
nand U22383 (N_22383,N_17582,N_18574);
or U22384 (N_22384,N_17609,N_19011);
nand U22385 (N_22385,N_18121,N_19635);
nand U22386 (N_22386,N_18867,N_19072);
or U22387 (N_22387,N_19558,N_19773);
or U22388 (N_22388,N_17768,N_17960);
and U22389 (N_22389,N_19337,N_19488);
nand U22390 (N_22390,N_19622,N_19375);
or U22391 (N_22391,N_19666,N_19259);
nand U22392 (N_22392,N_18588,N_19447);
nand U22393 (N_22393,N_18661,N_18662);
or U22394 (N_22394,N_18823,N_17880);
or U22395 (N_22395,N_17601,N_18537);
and U22396 (N_22396,N_19773,N_19702);
or U22397 (N_22397,N_19832,N_19761);
or U22398 (N_22398,N_19419,N_19773);
nand U22399 (N_22399,N_18444,N_18526);
or U22400 (N_22400,N_19531,N_19558);
nand U22401 (N_22401,N_19736,N_19579);
nand U22402 (N_22402,N_19318,N_17997);
or U22403 (N_22403,N_17900,N_17653);
nand U22404 (N_22404,N_18209,N_17559);
and U22405 (N_22405,N_18858,N_17932);
nand U22406 (N_22406,N_17950,N_19861);
nand U22407 (N_22407,N_18024,N_19607);
nor U22408 (N_22408,N_19452,N_17594);
and U22409 (N_22409,N_18095,N_19063);
nand U22410 (N_22410,N_18040,N_19895);
or U22411 (N_22411,N_19389,N_19779);
xnor U22412 (N_22412,N_18626,N_18681);
or U22413 (N_22413,N_19482,N_19129);
nor U22414 (N_22414,N_19552,N_19137);
or U22415 (N_22415,N_18760,N_18822);
or U22416 (N_22416,N_18205,N_17627);
nand U22417 (N_22417,N_19663,N_19587);
or U22418 (N_22418,N_17721,N_18161);
or U22419 (N_22419,N_18726,N_17706);
xnor U22420 (N_22420,N_18120,N_19974);
and U22421 (N_22421,N_18349,N_18496);
nor U22422 (N_22422,N_19589,N_19016);
and U22423 (N_22423,N_18257,N_19611);
nor U22424 (N_22424,N_18748,N_18703);
and U22425 (N_22425,N_19474,N_18927);
xnor U22426 (N_22426,N_19019,N_19334);
or U22427 (N_22427,N_18221,N_19726);
and U22428 (N_22428,N_19377,N_19056);
or U22429 (N_22429,N_18605,N_19396);
and U22430 (N_22430,N_19170,N_19931);
nor U22431 (N_22431,N_18070,N_18873);
and U22432 (N_22432,N_19507,N_19394);
and U22433 (N_22433,N_18229,N_17783);
xor U22434 (N_22434,N_17692,N_17619);
nor U22435 (N_22435,N_18008,N_19222);
and U22436 (N_22436,N_18527,N_18779);
nor U22437 (N_22437,N_19280,N_17932);
and U22438 (N_22438,N_17599,N_19913);
and U22439 (N_22439,N_18037,N_18837);
nor U22440 (N_22440,N_17780,N_17608);
nand U22441 (N_22441,N_18927,N_18006);
nor U22442 (N_22442,N_19620,N_18558);
or U22443 (N_22443,N_19588,N_18779);
nor U22444 (N_22444,N_18400,N_18761);
and U22445 (N_22445,N_18228,N_17633);
nand U22446 (N_22446,N_17931,N_17737);
and U22447 (N_22447,N_19129,N_19779);
nor U22448 (N_22448,N_18230,N_19287);
and U22449 (N_22449,N_18977,N_18454);
and U22450 (N_22450,N_18207,N_19954);
or U22451 (N_22451,N_19364,N_19466);
or U22452 (N_22452,N_18759,N_17614);
or U22453 (N_22453,N_18359,N_17659);
nor U22454 (N_22454,N_18053,N_17856);
and U22455 (N_22455,N_19185,N_18595);
nor U22456 (N_22456,N_19718,N_17896);
nor U22457 (N_22457,N_18454,N_17519);
nor U22458 (N_22458,N_18045,N_19573);
and U22459 (N_22459,N_18057,N_19497);
nor U22460 (N_22460,N_18521,N_19252);
or U22461 (N_22461,N_18654,N_19968);
xnor U22462 (N_22462,N_18246,N_18213);
and U22463 (N_22463,N_17622,N_18285);
and U22464 (N_22464,N_18568,N_19067);
xnor U22465 (N_22465,N_19715,N_17517);
nor U22466 (N_22466,N_18531,N_17895);
xnor U22467 (N_22467,N_18045,N_17979);
xnor U22468 (N_22468,N_17957,N_17808);
nor U22469 (N_22469,N_19998,N_17993);
xnor U22470 (N_22470,N_19515,N_18219);
nand U22471 (N_22471,N_18688,N_18215);
and U22472 (N_22472,N_18024,N_17507);
xnor U22473 (N_22473,N_18596,N_18453);
nand U22474 (N_22474,N_18433,N_17791);
nor U22475 (N_22475,N_18851,N_19331);
and U22476 (N_22476,N_19864,N_18178);
nor U22477 (N_22477,N_17962,N_17536);
or U22478 (N_22478,N_18353,N_19955);
and U22479 (N_22479,N_18213,N_19336);
nand U22480 (N_22480,N_19678,N_18223);
nor U22481 (N_22481,N_18140,N_19961);
and U22482 (N_22482,N_18677,N_17582);
and U22483 (N_22483,N_19565,N_19310);
xor U22484 (N_22484,N_19873,N_19460);
nor U22485 (N_22485,N_19071,N_19914);
nand U22486 (N_22486,N_18590,N_18528);
and U22487 (N_22487,N_18827,N_18260);
xor U22488 (N_22488,N_18258,N_17625);
xnor U22489 (N_22489,N_18584,N_19150);
nand U22490 (N_22490,N_18581,N_19585);
nor U22491 (N_22491,N_19548,N_18678);
and U22492 (N_22492,N_19965,N_19403);
nor U22493 (N_22493,N_19212,N_18137);
nor U22494 (N_22494,N_18553,N_19444);
nand U22495 (N_22495,N_19387,N_19629);
nand U22496 (N_22496,N_18275,N_19303);
and U22497 (N_22497,N_17578,N_19514);
and U22498 (N_22498,N_19330,N_19752);
nor U22499 (N_22499,N_18500,N_18280);
nand U22500 (N_22500,N_21416,N_20835);
xnor U22501 (N_22501,N_22239,N_21362);
nor U22502 (N_22502,N_20479,N_21344);
nand U22503 (N_22503,N_21163,N_20018);
xnor U22504 (N_22504,N_20546,N_20350);
nand U22505 (N_22505,N_22476,N_21969);
nor U22506 (N_22506,N_21276,N_20888);
or U22507 (N_22507,N_20948,N_21300);
nand U22508 (N_22508,N_20199,N_21766);
nor U22509 (N_22509,N_21378,N_21595);
nor U22510 (N_22510,N_21026,N_21626);
nand U22511 (N_22511,N_21236,N_21289);
nor U22512 (N_22512,N_20234,N_20300);
nand U22513 (N_22513,N_20067,N_20415);
or U22514 (N_22514,N_22477,N_22464);
nand U22515 (N_22515,N_21352,N_21886);
nor U22516 (N_22516,N_20397,N_21423);
xnor U22517 (N_22517,N_20187,N_21814);
nand U22518 (N_22518,N_20190,N_21000);
and U22519 (N_22519,N_20308,N_21082);
nor U22520 (N_22520,N_21979,N_21386);
nand U22521 (N_22521,N_20060,N_20727);
nand U22522 (N_22522,N_22409,N_22350);
nand U22523 (N_22523,N_20609,N_20878);
nand U22524 (N_22524,N_22018,N_22094);
nand U22525 (N_22525,N_20864,N_20023);
xnor U22526 (N_22526,N_20443,N_21197);
xor U22527 (N_22527,N_21327,N_20445);
or U22528 (N_22528,N_22147,N_21575);
xnor U22529 (N_22529,N_21133,N_20163);
nand U22530 (N_22530,N_21643,N_20162);
and U22531 (N_22531,N_20282,N_20976);
nand U22532 (N_22532,N_20395,N_21436);
and U22533 (N_22533,N_21426,N_20161);
and U22534 (N_22534,N_22376,N_22057);
nand U22535 (N_22535,N_21737,N_20891);
or U22536 (N_22536,N_21865,N_20863);
nand U22537 (N_22537,N_20555,N_22141);
or U22538 (N_22538,N_22280,N_21347);
nor U22539 (N_22539,N_20268,N_21278);
and U22540 (N_22540,N_21847,N_20184);
xnor U22541 (N_22541,N_21075,N_20764);
and U22542 (N_22542,N_20689,N_20450);
nand U22543 (N_22543,N_21809,N_21369);
nand U22544 (N_22544,N_20077,N_21356);
nand U22545 (N_22545,N_20478,N_20579);
or U22546 (N_22546,N_21337,N_22438);
or U22547 (N_22547,N_21898,N_22312);
xnor U22548 (N_22548,N_20514,N_20344);
nand U22549 (N_22549,N_21741,N_21852);
or U22550 (N_22550,N_20877,N_20881);
or U22551 (N_22551,N_20797,N_22112);
and U22552 (N_22552,N_20492,N_20916);
xnor U22553 (N_22553,N_20226,N_20735);
and U22554 (N_22554,N_21102,N_20982);
and U22555 (N_22555,N_21259,N_20611);
nand U22556 (N_22556,N_20346,N_20964);
or U22557 (N_22557,N_20848,N_20588);
nand U22558 (N_22558,N_21660,N_21552);
nand U22559 (N_22559,N_21962,N_22049);
or U22560 (N_22560,N_22213,N_20885);
xnor U22561 (N_22561,N_22490,N_20311);
and U22562 (N_22562,N_20527,N_20124);
or U22563 (N_22563,N_22260,N_21535);
or U22564 (N_22564,N_20194,N_20994);
or U22565 (N_22565,N_20010,N_22048);
and U22566 (N_22566,N_21353,N_22287);
nor U22567 (N_22567,N_20151,N_22053);
and U22568 (N_22568,N_20560,N_21345);
nand U22569 (N_22569,N_22098,N_21086);
and U22570 (N_22570,N_21183,N_22027);
nor U22571 (N_22571,N_20818,N_21717);
nor U22572 (N_22572,N_20203,N_22069);
and U22573 (N_22573,N_20025,N_20592);
nand U22574 (N_22574,N_21946,N_20690);
nand U22575 (N_22575,N_22468,N_20629);
nand U22576 (N_22576,N_20080,N_21406);
and U22577 (N_22577,N_21457,N_22430);
nand U22578 (N_22578,N_20271,N_21387);
xnor U22579 (N_22579,N_22116,N_21617);
nand U22580 (N_22580,N_20167,N_21682);
nand U22581 (N_22581,N_20286,N_21905);
nor U22582 (N_22582,N_22181,N_22104);
nand U22583 (N_22583,N_21128,N_22082);
and U22584 (N_22584,N_20854,N_20128);
nand U22585 (N_22585,N_21718,N_21733);
nor U22586 (N_22586,N_20558,N_21155);
or U22587 (N_22587,N_22066,N_22336);
or U22588 (N_22588,N_21107,N_20784);
or U22589 (N_22589,N_21459,N_20157);
and U22590 (N_22590,N_22404,N_22257);
nor U22591 (N_22591,N_20660,N_21885);
xnor U22592 (N_22592,N_20298,N_21937);
and U22593 (N_22593,N_21392,N_21448);
and U22594 (N_22594,N_21869,N_21250);
and U22595 (N_22595,N_20971,N_20534);
and U22596 (N_22596,N_21669,N_22361);
or U22597 (N_22597,N_21631,N_21950);
or U22598 (N_22598,N_20827,N_22209);
nor U22599 (N_22599,N_20383,N_22444);
nor U22600 (N_22600,N_22122,N_22331);
nand U22601 (N_22601,N_21523,N_22422);
nor U22602 (N_22602,N_20375,N_22414);
and U22603 (N_22603,N_20024,N_22394);
nor U22604 (N_22604,N_20378,N_21980);
or U22605 (N_22605,N_21228,N_21999);
and U22606 (N_22606,N_20637,N_22222);
and U22607 (N_22607,N_22272,N_20561);
xnor U22608 (N_22608,N_21934,N_21903);
or U22609 (N_22609,N_20084,N_20035);
nor U22610 (N_22610,N_22005,N_22443);
nor U22611 (N_22611,N_21433,N_21062);
nand U22612 (N_22612,N_20762,N_22183);
nand U22613 (N_22613,N_20063,N_22292);
nand U22614 (N_22614,N_22378,N_22220);
and U22615 (N_22615,N_22145,N_20713);
nand U22616 (N_22616,N_21602,N_22470);
xnor U22617 (N_22617,N_20135,N_22172);
or U22618 (N_22618,N_21654,N_22363);
or U22619 (N_22619,N_21394,N_20321);
and U22620 (N_22620,N_21398,N_20123);
nor U22621 (N_22621,N_22229,N_20759);
nor U22622 (N_22622,N_20153,N_20086);
and U22623 (N_22623,N_22319,N_21634);
and U22624 (N_22624,N_22396,N_22189);
nor U22625 (N_22625,N_22389,N_22129);
xnor U22626 (N_22626,N_20515,N_22061);
nor U22627 (N_22627,N_22111,N_21720);
nor U22628 (N_22628,N_20334,N_20800);
or U22629 (N_22629,N_21877,N_21312);
nand U22630 (N_22630,N_21685,N_20511);
nand U22631 (N_22631,N_22461,N_21712);
or U22632 (N_22632,N_20285,N_20239);
and U22633 (N_22633,N_20704,N_20869);
nor U22634 (N_22634,N_20246,N_21042);
nand U22635 (N_22635,N_21794,N_22177);
nand U22636 (N_22636,N_20997,N_21373);
and U22637 (N_22637,N_20129,N_20834);
nand U22638 (N_22638,N_20882,N_21543);
or U22639 (N_22639,N_20504,N_20955);
nor U22640 (N_22640,N_21301,N_22352);
nand U22641 (N_22641,N_20512,N_21213);
and U22642 (N_22642,N_21243,N_21853);
or U22643 (N_22643,N_20741,N_21451);
nor U22644 (N_22644,N_20033,N_20027);
or U22645 (N_22645,N_20752,N_21405);
or U22646 (N_22646,N_22277,N_22339);
or U22647 (N_22647,N_21145,N_22424);
xnor U22648 (N_22648,N_21058,N_20493);
and U22649 (N_22649,N_20614,N_20975);
nor U22650 (N_22650,N_22089,N_20461);
or U22651 (N_22651,N_22371,N_20076);
nand U22652 (N_22652,N_21695,N_22279);
or U22653 (N_22653,N_22403,N_21256);
and U22654 (N_22654,N_20841,N_20968);
and U22655 (N_22655,N_21791,N_22499);
or U22656 (N_22656,N_21568,N_22046);
and U22657 (N_22657,N_22263,N_21430);
or U22658 (N_22658,N_20926,N_21648);
nand U22659 (N_22659,N_20826,N_21103);
or U22660 (N_22660,N_22191,N_21828);
and U22661 (N_22661,N_20409,N_22271);
and U22662 (N_22662,N_21551,N_22010);
nor U22663 (N_22663,N_20840,N_22140);
nand U22664 (N_22664,N_21330,N_20915);
or U22665 (N_22665,N_20543,N_20989);
nor U22666 (N_22666,N_21024,N_20932);
nor U22667 (N_22667,N_21715,N_21917);
nand U22668 (N_22668,N_20216,N_20455);
nor U22669 (N_22669,N_20981,N_22273);
nand U22670 (N_22670,N_20739,N_21558);
and U22671 (N_22671,N_21269,N_22332);
nand U22672 (N_22672,N_21901,N_20481);
and U22673 (N_22673,N_21341,N_20627);
nand U22674 (N_22674,N_20570,N_20571);
nand U22675 (N_22675,N_20541,N_21578);
nor U22676 (N_22676,N_20936,N_21131);
nand U22677 (N_22677,N_20717,N_20638);
xor U22678 (N_22678,N_21659,N_20255);
and U22679 (N_22679,N_22455,N_22096);
nor U22680 (N_22680,N_20348,N_21808);
nand U22681 (N_22681,N_22103,N_21870);
nand U22682 (N_22682,N_22206,N_22025);
nor U22683 (N_22683,N_21252,N_21196);
nor U22684 (N_22684,N_21144,N_20567);
and U22685 (N_22685,N_21235,N_21326);
or U22686 (N_22686,N_20209,N_21125);
and U22687 (N_22687,N_22131,N_21759);
or U22688 (N_22688,N_21566,N_20978);
nor U22689 (N_22689,N_20520,N_20715);
nand U22690 (N_22690,N_20486,N_21015);
and U22691 (N_22691,N_22083,N_20391);
and U22692 (N_22692,N_21921,N_21149);
or U22693 (N_22693,N_20488,N_20559);
or U22694 (N_22694,N_22058,N_20657);
nor U22695 (N_22695,N_21271,N_20783);
nand U22696 (N_22696,N_20171,N_20829);
or U22697 (N_22697,N_20808,N_21105);
nor U22698 (N_22698,N_21052,N_20725);
and U22699 (N_22699,N_20116,N_22199);
and U22700 (N_22700,N_21773,N_20751);
or U22701 (N_22701,N_21306,N_21399);
nor U22702 (N_22702,N_21478,N_20273);
nor U22703 (N_22703,N_20332,N_21764);
xnor U22704 (N_22704,N_21468,N_20695);
nor U22705 (N_22705,N_20089,N_20069);
and U22706 (N_22706,N_21630,N_21233);
nor U22707 (N_22707,N_21684,N_21806);
or U22708 (N_22708,N_22202,N_21624);
nor U22709 (N_22709,N_22134,N_21040);
nand U22710 (N_22710,N_22020,N_20448);
or U22711 (N_22711,N_22054,N_22442);
or U22712 (N_22712,N_20257,N_22024);
nor U22713 (N_22713,N_22495,N_21424);
nand U22714 (N_22714,N_21198,N_20687);
xnor U22715 (N_22715,N_21751,N_22415);
or U22716 (N_22716,N_20770,N_20112);
xnor U22717 (N_22717,N_22268,N_20471);
nand U22718 (N_22718,N_22086,N_22227);
nor U22719 (N_22719,N_21428,N_20718);
and U22720 (N_22720,N_22360,N_21588);
nand U22721 (N_22721,N_20954,N_21091);
nand U22722 (N_22722,N_22395,N_22317);
nor U22723 (N_22723,N_20529,N_22467);
and U22724 (N_22724,N_21221,N_20453);
nor U22725 (N_22725,N_21444,N_21382);
and U22726 (N_22726,N_21829,N_22356);
nand U22727 (N_22727,N_20533,N_21364);
nand U22728 (N_22728,N_21132,N_21953);
or U22729 (N_22729,N_21411,N_22076);
xor U22730 (N_22730,N_21612,N_20156);
and U22731 (N_22731,N_20091,N_21332);
nor U22732 (N_22732,N_21704,N_21971);
nor U22733 (N_22733,N_21227,N_21517);
nand U22734 (N_22734,N_20223,N_22168);
nand U22735 (N_22735,N_22454,N_20736);
nor U22736 (N_22736,N_20798,N_20327);
nand U22737 (N_22737,N_20889,N_21959);
and U22738 (N_22738,N_20367,N_20436);
nand U22739 (N_22739,N_22347,N_21212);
and U22740 (N_22740,N_20711,N_21796);
or U22741 (N_22741,N_21201,N_20119);
and U22742 (N_22742,N_20118,N_22327);
or U22743 (N_22743,N_22100,N_20786);
nor U22744 (N_22744,N_21846,N_21435);
xnor U22745 (N_22745,N_22377,N_21524);
and U22746 (N_22746,N_20110,N_21570);
nor U22747 (N_22747,N_21175,N_20137);
and U22748 (N_22748,N_20940,N_22426);
and U22749 (N_22749,N_22380,N_21887);
or U22750 (N_22750,N_20422,N_21838);
xor U22751 (N_22751,N_22250,N_21122);
xnor U22752 (N_22752,N_20056,N_21936);
or U22753 (N_22753,N_21943,N_22472);
and U22754 (N_22754,N_21319,N_21801);
or U22755 (N_22755,N_20993,N_20211);
xnor U22756 (N_22756,N_20340,N_21622);
and U22757 (N_22757,N_20355,N_22407);
or U22758 (N_22758,N_21134,N_21765);
or U22759 (N_22759,N_20399,N_21786);
nand U22760 (N_22760,N_20779,N_21117);
or U22761 (N_22761,N_21172,N_22249);
or U22762 (N_22762,N_21991,N_20122);
nor U22763 (N_22763,N_21963,N_22451);
or U22764 (N_22764,N_22235,N_21391);
nand U22765 (N_22765,N_20961,N_21967);
xnor U22766 (N_22766,N_20210,N_22487);
or U22767 (N_22767,N_21047,N_20856);
and U22768 (N_22768,N_21005,N_22037);
and U22769 (N_22769,N_22298,N_21013);
nand U22770 (N_22770,N_21264,N_21830);
nor U22771 (N_22771,N_22119,N_20754);
nor U22772 (N_22772,N_22182,N_20291);
and U22773 (N_22773,N_20011,N_21672);
nand U22774 (N_22774,N_21204,N_20523);
nor U22775 (N_22775,N_21006,N_20883);
or U22776 (N_22776,N_20101,N_21135);
nor U22777 (N_22777,N_21842,N_22022);
and U22778 (N_22778,N_22445,N_20031);
xor U22779 (N_22779,N_21510,N_21483);
or U22780 (N_22780,N_22346,N_20790);
or U22781 (N_22781,N_21057,N_21036);
nor U22782 (N_22782,N_21409,N_21789);
nand U22783 (N_22783,N_21372,N_21035);
or U22784 (N_22784,N_21475,N_21257);
nand U22785 (N_22785,N_22408,N_20668);
xnor U22786 (N_22786,N_20359,N_20740);
xor U22787 (N_22787,N_22033,N_20463);
or U22788 (N_22788,N_21965,N_22391);
and U22789 (N_22789,N_21313,N_20960);
nor U22790 (N_22790,N_20302,N_21489);
nand U22791 (N_22791,N_21318,N_22078);
or U22792 (N_22792,N_22435,N_20061);
or U22793 (N_22793,N_21835,N_21431);
nor U22794 (N_22794,N_21249,N_21787);
and U22795 (N_22795,N_21707,N_20671);
and U22796 (N_22796,N_22198,N_21792);
nand U22797 (N_22797,N_21066,N_22091);
and U22798 (N_22798,N_21731,N_20979);
nand U22799 (N_22799,N_22106,N_20905);
or U22800 (N_22800,N_21855,N_21195);
nor U22801 (N_22801,N_21650,N_21742);
xor U22802 (N_22802,N_21390,N_21627);
or U22803 (N_22803,N_20237,N_20143);
xnor U22804 (N_22804,N_20097,N_20102);
nand U22805 (N_22805,N_20900,N_20678);
or U22806 (N_22806,N_21490,N_21701);
xnor U22807 (N_22807,N_22232,N_22234);
nor U22808 (N_22808,N_21140,N_22115);
and U22809 (N_22809,N_21929,N_20828);
nand U22810 (N_22810,N_21713,N_22265);
nand U22811 (N_22811,N_20674,N_20966);
nand U22812 (N_22812,N_20303,N_22335);
and U22813 (N_22813,N_21586,N_22255);
xnor U22814 (N_22814,N_21214,N_20701);
nand U22815 (N_22815,N_21079,N_20049);
or U22816 (N_22816,N_22252,N_20871);
and U22817 (N_22817,N_20662,N_21290);
and U22818 (N_22818,N_21048,N_21008);
nor U22819 (N_22819,N_20029,N_21802);
nand U22820 (N_22820,N_21606,N_21994);
nand U22821 (N_22821,N_20221,N_20326);
xor U22822 (N_22822,N_20501,N_20707);
and U22823 (N_22823,N_20050,N_21819);
nor U22824 (N_22824,N_21536,N_21442);
nor U22825 (N_22825,N_21506,N_21826);
and U22826 (N_22826,N_21260,N_21790);
nor U22827 (N_22827,N_21644,N_20503);
or U22828 (N_22828,N_20051,N_20824);
or U22829 (N_22829,N_20601,N_20890);
nand U22830 (N_22830,N_21261,N_20604);
or U22831 (N_22831,N_22275,N_20476);
and U22832 (N_22832,N_20850,N_21844);
nor U22833 (N_22833,N_21480,N_22351);
and U22834 (N_22834,N_21652,N_21094);
nor U22835 (N_22835,N_21817,N_20676);
nor U22836 (N_22836,N_22294,N_21174);
nand U22837 (N_22837,N_21966,N_20653);
or U22838 (N_22838,N_20912,N_20973);
nand U22839 (N_22839,N_20250,N_22028);
and U22840 (N_22840,N_21600,N_21605);
or U22841 (N_22841,N_21031,N_21771);
nor U22842 (N_22842,N_20530,N_20763);
nand U22843 (N_22843,N_21297,N_20289);
nand U22844 (N_22844,N_22215,N_21618);
nor U22845 (N_22845,N_21653,N_21975);
and U22846 (N_22846,N_21232,N_20939);
and U22847 (N_22847,N_22488,N_22450);
nand U22848 (N_22848,N_20694,N_20219);
nand U22849 (N_22849,N_20313,N_21774);
or U22850 (N_22850,N_22449,N_22063);
nor U22851 (N_22851,N_21841,N_21218);
nand U22852 (N_22852,N_20109,N_22055);
or U22853 (N_22853,N_22469,N_21349);
and U22854 (N_22854,N_20917,N_21001);
nand U22855 (N_22855,N_20908,N_21358);
or U22856 (N_22856,N_20158,N_22186);
xnor U22857 (N_22857,N_21793,N_20988);
nand U22858 (N_22858,N_21284,N_22418);
or U22859 (N_22859,N_22211,N_21178);
or U22860 (N_22860,N_21460,N_21656);
or U22861 (N_22861,N_21189,N_21299);
xor U22862 (N_22862,N_21585,N_21990);
or U22863 (N_22863,N_21242,N_20618);
nand U22864 (N_22864,N_20130,N_22301);
or U22865 (N_22865,N_20758,N_22300);
or U22866 (N_22866,N_22125,N_20147);
and U22867 (N_22867,N_21873,N_21686);
xnor U22868 (N_22868,N_21651,N_21871);
and U22869 (N_22869,N_21880,N_21158);
or U22870 (N_22870,N_21286,N_21157);
xor U22871 (N_22871,N_21797,N_21170);
nand U22872 (N_22872,N_20342,N_21938);
or U22873 (N_22873,N_20283,N_21893);
nand U22874 (N_22874,N_22355,N_21099);
nor U22875 (N_22875,N_20489,N_22192);
and U22876 (N_22876,N_21488,N_22373);
nand U22877 (N_22877,N_21674,N_20572);
and U22878 (N_22878,N_22493,N_20120);
nand U22879 (N_22879,N_22475,N_21499);
and U22880 (N_22880,N_22353,N_20983);
and U22881 (N_22881,N_21033,N_21926);
nor U22882 (N_22882,N_21804,N_21217);
or U22883 (N_22883,N_21646,N_21940);
xnor U22884 (N_22884,N_21528,N_22074);
nor U22885 (N_22885,N_22153,N_22099);
nand U22886 (N_22886,N_22052,N_21714);
nor U22887 (N_22887,N_21445,N_21987);
or U22888 (N_22888,N_21721,N_20262);
or U22889 (N_22889,N_20716,N_21508);
and U22890 (N_22890,N_20996,N_20886);
nor U22891 (N_22891,N_21825,N_21609);
xnor U22892 (N_22892,N_20269,N_20505);
nor U22893 (N_22893,N_21692,N_20875);
nand U22894 (N_22894,N_22204,N_21710);
and U22895 (N_22895,N_20942,N_20938);
or U22896 (N_22896,N_22108,N_22245);
nand U22897 (N_22897,N_21941,N_20995);
or U22898 (N_22898,N_20336,N_20483);
or U22899 (N_22899,N_20466,N_21813);
nand U22900 (N_22900,N_20057,N_21758);
and U22901 (N_22901,N_20853,N_20460);
nand U22902 (N_22902,N_21064,N_20215);
and U22903 (N_22903,N_21205,N_20584);
or U22904 (N_22904,N_21760,N_21018);
and U22905 (N_22905,N_21884,N_22474);
nand U22906 (N_22906,N_20360,N_20406);
nor U22907 (N_22907,N_20594,N_22297);
nor U22908 (N_22908,N_21171,N_21509);
and U22909 (N_22909,N_21756,N_21348);
nand U22910 (N_22910,N_20901,N_21114);
xnor U22911 (N_22911,N_20004,N_22023);
and U22912 (N_22912,N_20170,N_21619);
or U22913 (N_22913,N_22374,N_21121);
nor U22914 (N_22914,N_20799,N_20785);
and U22915 (N_22915,N_21918,N_21060);
nor U22916 (N_22916,N_21223,N_20266);
and U22917 (N_22917,N_20094,N_20418);
nand U22918 (N_22918,N_20108,N_20910);
nand U22919 (N_22919,N_21632,N_20183);
and U22920 (N_22920,N_21550,N_22453);
and U22921 (N_22921,N_22440,N_21541);
or U22922 (N_22922,N_22233,N_20892);
nand U22923 (N_22923,N_22486,N_22276);
nand U22924 (N_22924,N_20107,N_22345);
xor U22925 (N_22925,N_21723,N_20794);
nor U22926 (N_22926,N_20849,N_20791);
and U22927 (N_22927,N_22228,N_21303);
and U22928 (N_22928,N_21988,N_22207);
nand U22929 (N_22929,N_20615,N_20923);
nor U22930 (N_22930,N_20034,N_20003);
nand U22931 (N_22931,N_21857,N_21845);
xnor U22932 (N_22932,N_21913,N_21661);
and U22933 (N_22933,N_21727,N_21474);
nor U22934 (N_22934,N_20692,N_20398);
or U22935 (N_22935,N_20087,N_21415);
or U22936 (N_22936,N_21194,N_20263);
nor U22937 (N_22937,N_20722,N_21978);
or U22938 (N_22938,N_20251,N_20729);
nand U22939 (N_22939,N_21241,N_21580);
and U22940 (N_22940,N_20253,N_21851);
or U22941 (N_22941,N_22341,N_21417);
nor U22942 (N_22942,N_21287,N_20607);
and U22943 (N_22943,N_22175,N_20986);
nor U22944 (N_22944,N_21366,N_20175);
and U22945 (N_22945,N_20059,N_21203);
nand U22946 (N_22946,N_21533,N_22458);
nand U22947 (N_22947,N_20085,N_20401);
nand U22948 (N_22948,N_20768,N_20258);
or U22949 (N_22949,N_21788,N_20793);
or U22950 (N_22950,N_21004,N_20956);
nor U22951 (N_22951,N_21583,N_22081);
nor U22952 (N_22952,N_20081,N_22375);
and U22953 (N_22953,N_20281,N_20805);
and U22954 (N_22954,N_20887,N_20549);
nand U22955 (N_22955,N_21699,N_21812);
xor U22956 (N_22956,N_20773,N_22372);
or U22957 (N_22957,N_20036,N_22496);
nor U22958 (N_22958,N_20371,N_21803);
nor U22959 (N_22959,N_22225,N_20345);
and U22960 (N_22960,N_20817,N_20329);
nor U22961 (N_22961,N_20434,N_22230);
and U22962 (N_22962,N_20999,N_21253);
nor U22963 (N_22963,N_20366,N_21747);
or U22964 (N_22964,N_21996,N_21447);
nor U22965 (N_22965,N_20306,N_20620);
or U22966 (N_22966,N_21820,N_20895);
nand U22967 (N_22967,N_22330,N_20760);
nand U22968 (N_22968,N_20240,N_21432);
or U22969 (N_22969,N_22219,N_20491);
nand U22970 (N_22970,N_21534,N_21437);
nor U22971 (N_22971,N_20022,N_21557);
nand U22972 (N_22972,N_20179,N_20945);
and U22973 (N_22973,N_21467,N_22073);
and U22974 (N_22974,N_20622,N_20231);
xnor U22975 (N_22975,N_21384,N_20602);
or U22976 (N_22976,N_20680,N_20054);
nand U22977 (N_22977,N_21729,N_21649);
or U22978 (N_22978,N_20696,N_20899);
nand U22979 (N_22979,N_21702,N_21662);
and U22980 (N_22980,N_20655,N_21821);
xnor U22981 (N_22981,N_20613,N_20953);
and U22982 (N_22982,N_22483,N_22379);
and U22983 (N_22983,N_20047,N_20082);
xnor U22984 (N_22984,N_20586,N_20628);
nand U22985 (N_22985,N_21968,N_21401);
and U22986 (N_22986,N_22328,N_20104);
and U22987 (N_22987,N_22165,N_21106);
nor U22988 (N_22988,N_20749,N_20508);
xnor U22989 (N_22989,N_21207,N_21574);
nand U22990 (N_22990,N_21565,N_22214);
and U22991 (N_22991,N_22002,N_20113);
and U22992 (N_22992,N_21562,N_20860);
or U22993 (N_22993,N_21573,N_21899);
nor U22994 (N_22994,N_21932,N_20064);
and U22995 (N_22995,N_20806,N_20426);
nor U22996 (N_22996,N_21584,N_20164);
nor U22997 (N_22997,N_20845,N_21051);
nor U22998 (N_22998,N_22405,N_20669);
or U22999 (N_22999,N_21897,N_20139);
and U23000 (N_23000,N_20407,N_22288);
xor U23001 (N_23001,N_22001,N_20623);
nand U23002 (N_23002,N_21407,N_21027);
and U23003 (N_23003,N_20771,N_20733);
nand U23004 (N_23004,N_20893,N_21500);
nor U23005 (N_23005,N_21097,N_20152);
or U23006 (N_23006,N_20468,N_21531);
and U23007 (N_23007,N_21141,N_20985);
or U23008 (N_23008,N_20042,N_20804);
xnor U23009 (N_23009,N_22421,N_21683);
or U23010 (N_23010,N_20847,N_21434);
and U23011 (N_23011,N_22065,N_20545);
or U23012 (N_23012,N_20103,N_21768);
or U23013 (N_23013,N_21315,N_22067);
and U23014 (N_23014,N_20232,N_20755);
nand U23015 (N_23015,N_20127,N_20384);
nor U23016 (N_23016,N_21603,N_21334);
and U23017 (N_23017,N_21663,N_22036);
nand U23018 (N_23018,N_20382,N_21538);
and U23019 (N_23019,N_20838,N_22386);
nor U23020 (N_23020,N_20233,N_22492);
nor U23021 (N_23021,N_21350,N_22325);
xor U23022 (N_23022,N_21961,N_21449);
and U23023 (N_23023,N_20719,N_21539);
and U23024 (N_23024,N_22237,N_20980);
nand U23025 (N_23025,N_21059,N_20666);
xor U23026 (N_23026,N_21211,N_20098);
or U23027 (N_23027,N_22132,N_22253);
or U23028 (N_23028,N_22236,N_21705);
nor U23029 (N_23029,N_20709,N_21440);
nor U23030 (N_23030,N_20922,N_21069);
nand U23031 (N_23031,N_20169,N_21516);
nor U23032 (N_23032,N_21115,N_20159);
nor U23033 (N_23033,N_22243,N_21696);
and U23034 (N_23034,N_20410,N_20521);
or U23035 (N_23035,N_21043,N_20987);
nand U23036 (N_23036,N_21738,N_20354);
or U23037 (N_23037,N_20575,N_22307);
xnor U23038 (N_23038,N_20208,N_21637);
nand U23039 (N_23039,N_22029,N_20788);
or U23040 (N_23040,N_20325,N_22208);
nor U23041 (N_23041,N_20580,N_20747);
xor U23042 (N_23042,N_21778,N_22437);
and U23043 (N_23043,N_22417,N_21493);
or U23044 (N_23044,N_20020,N_21945);
nand U23045 (N_23045,N_20447,N_20884);
xnor U23046 (N_23046,N_20402,N_21486);
nand U23047 (N_23047,N_20017,N_22254);
or U23048 (N_23048,N_21180,N_22357);
nor U23049 (N_23049,N_20634,N_20862);
nand U23050 (N_23050,N_22196,N_21840);
and U23051 (N_23051,N_20991,N_20055);
and U23052 (N_23052,N_21017,N_21666);
and U23053 (N_23053,N_22342,N_22427);
nand U23054 (N_23054,N_20337,N_20778);
and U23055 (N_23055,N_20928,N_20392);
and U23056 (N_23056,N_21776,N_20930);
nor U23057 (N_23057,N_21782,N_20259);
nand U23058 (N_23058,N_22171,N_20941);
nand U23059 (N_23059,N_20145,N_21670);
nand U23060 (N_23060,N_21636,N_20013);
nand U23061 (N_23061,N_21507,N_22462);
and U23062 (N_23062,N_21225,N_20723);
nand U23063 (N_23063,N_21272,N_22318);
nand U23064 (N_23064,N_21339,N_21138);
nand U23065 (N_23065,N_20698,N_22008);
nor U23066 (N_23066,N_20509,N_20554);
or U23067 (N_23067,N_20338,N_20001);
or U23068 (N_23068,N_20472,N_21564);
nor U23069 (N_23069,N_21555,N_22340);
or U23070 (N_23070,N_20278,N_20720);
or U23071 (N_23071,N_22152,N_22216);
nand U23072 (N_23072,N_21657,N_21267);
and U23073 (N_23073,N_20526,N_20525);
or U23074 (N_23074,N_20168,N_22185);
or U23075 (N_23075,N_20477,N_21623);
nor U23076 (N_23076,N_22241,N_21034);
and U23077 (N_23077,N_20537,N_22013);
nor U23078 (N_23078,N_21504,N_20368);
nor U23079 (N_23079,N_21268,N_21162);
and U23080 (N_23080,N_21719,N_20173);
or U23081 (N_23081,N_21995,N_21532);
nor U23082 (N_23082,N_21161,N_20815);
xnor U23083 (N_23083,N_22267,N_21323);
nand U23084 (N_23084,N_20149,N_21410);
nand U23085 (N_23085,N_20195,N_20897);
or U23086 (N_23086,N_20552,N_22436);
and U23087 (N_23087,N_20358,N_20812);
and U23088 (N_23088,N_21379,N_21951);
nor U23089 (N_23089,N_21755,N_20777);
or U23090 (N_23090,N_22343,N_20576);
or U23091 (N_23091,N_21544,N_21496);
nand U23092 (N_23092,N_20229,N_22393);
nor U23093 (N_23093,N_20174,N_20556);
and U23094 (N_23094,N_21216,N_20444);
or U23095 (N_23095,N_20879,N_22428);
xor U23096 (N_23096,N_22047,N_22366);
nor U23097 (N_23097,N_20645,N_21724);
or U23098 (N_23098,N_20413,N_20248);
or U23099 (N_23099,N_21815,N_20469);
and U23100 (N_23100,N_22359,N_20825);
xor U23101 (N_23101,N_21693,N_22126);
or U23102 (N_23102,N_20353,N_21044);
nor U23103 (N_23103,N_20438,N_21354);
nand U23104 (N_23104,N_21481,N_21009);
nor U23105 (N_23105,N_21126,N_21942);
xor U23106 (N_23106,N_20731,N_20374);
xnor U23107 (N_23107,N_21346,N_21479);
and U23108 (N_23108,N_22401,N_20304);
nor U23109 (N_23109,N_21482,N_21933);
xnor U23110 (N_23110,N_20074,N_21716);
and U23111 (N_23111,N_20290,N_20131);
xor U23112 (N_23112,N_20624,N_20925);
or U23113 (N_23113,N_20693,N_20949);
nand U23114 (N_23114,N_20324,N_21050);
xor U23115 (N_23115,N_20212,N_20563);
nand U23116 (N_23116,N_22247,N_21084);
and U23117 (N_23117,N_21924,N_21441);
nor U23118 (N_23118,N_21862,N_20030);
nand U23119 (N_23119,N_20934,N_22446);
nand U23120 (N_23120,N_21070,N_21836);
nor U23121 (N_23121,N_21664,N_22261);
nand U23122 (N_23122,N_20317,N_20792);
or U23123 (N_23123,N_21329,N_22156);
nand U23124 (N_23124,N_22210,N_21087);
or U23125 (N_23125,N_20380,N_20920);
nand U23126 (N_23126,N_22167,N_21615);
or U23127 (N_23127,N_21956,N_21484);
and U23128 (N_23128,N_22419,N_20487);
or U23129 (N_23129,N_22051,N_22090);
or U23130 (N_23130,N_21827,N_20045);
nand U23131 (N_23131,N_20507,N_20721);
or U23132 (N_23132,N_20593,N_20408);
and U23133 (N_23133,N_21039,N_20836);
nor U23134 (N_23134,N_22200,N_21244);
nand U23135 (N_23135,N_21054,N_20454);
and U23136 (N_23136,N_20083,N_20432);
or U23137 (N_23137,N_20032,N_20921);
and U23138 (N_23138,N_21298,N_21931);
and U23139 (N_23139,N_20333,N_22071);
nand U23140 (N_23140,N_20522,N_21689);
nor U23141 (N_23141,N_20439,N_22246);
nand U23142 (N_23142,N_21472,N_21331);
nor U23143 (N_23143,N_21156,N_22040);
nand U23144 (N_23144,N_20160,N_20414);
nor U23145 (N_23145,N_21761,N_20946);
and U23146 (N_23146,N_20417,N_21202);
nor U23147 (N_23147,N_21307,N_22296);
xor U23148 (N_23148,N_20814,N_21032);
and U23149 (N_23149,N_22075,N_21757);
nand U23150 (N_23150,N_20274,N_21295);
nand U23151 (N_23151,N_22097,N_20114);
or U23152 (N_23152,N_21143,N_21964);
nand U23153 (N_23153,N_20037,N_20117);
nand U23154 (N_23154,N_21335,N_20428);
xnor U23155 (N_23155,N_21370,N_20535);
or U23156 (N_23156,N_20021,N_20902);
or U23157 (N_23157,N_20066,N_22079);
and U23158 (N_23158,N_21188,N_21518);
or U23159 (N_23159,N_20608,N_21120);
nor U23160 (N_23160,N_20241,N_22240);
nand U23161 (N_23161,N_21016,N_21209);
nor U23162 (N_23162,N_21960,N_20557);
nor U23163 (N_23163,N_22161,N_21549);
nand U23164 (N_23164,N_21316,N_20518);
nand U23165 (N_23165,N_21446,N_20654);
and U23166 (N_23166,N_20485,N_21123);
or U23167 (N_23167,N_20217,N_20379);
nor U23168 (N_23168,N_20640,N_21860);
nand U23169 (N_23169,N_20710,N_21698);
nor U23170 (N_23170,N_21743,N_22334);
nand U23171 (N_23171,N_22491,N_21864);
nand U23172 (N_23172,N_20765,N_21007);
nand U23173 (N_23173,N_22323,N_21781);
and U23174 (N_23174,N_21165,N_21735);
or U23175 (N_23175,N_21101,N_22251);
and U23176 (N_23176,N_22149,N_21292);
nor U23177 (N_23177,N_20482,N_20296);
and U23178 (N_23178,N_21169,N_20458);
nand U23179 (N_23179,N_22085,N_22148);
nand U23180 (N_23180,N_20756,N_22441);
or U23181 (N_23181,N_20363,N_20992);
nor U23182 (N_23182,N_22142,N_22479);
nor U23183 (N_23183,N_21904,N_21511);
and U23184 (N_23184,N_20649,N_20430);
nor U23185 (N_23185,N_20318,N_20356);
or U23186 (N_23186,N_21638,N_21067);
and U23187 (N_23187,N_20207,N_20681);
and U23188 (N_23188,N_21546,N_21772);
nand U23189 (N_23189,N_20284,N_20644);
and U23190 (N_23190,N_21582,N_21908);
and U23191 (N_23191,N_21856,N_21041);
and U23192 (N_23192,N_20347,N_22173);
and U23193 (N_23193,N_21746,N_20568);
or U23194 (N_23194,N_22068,N_22315);
nand U23195 (N_23195,N_21336,N_20236);
nor U23196 (N_23196,N_21667,N_21697);
xor U23197 (N_23197,N_22130,N_20490);
nor U23198 (N_23198,N_21779,N_21080);
and U23199 (N_23199,N_20548,N_21675);
nor U23200 (N_23200,N_21247,N_22390);
and U23201 (N_23201,N_20155,N_21073);
and U23202 (N_23202,N_22270,N_22056);
nor U23203 (N_23203,N_20831,N_22195);
nor U23204 (N_23204,N_22184,N_20706);
xor U23205 (N_23205,N_21258,N_21984);
nor U23206 (N_23206,N_20277,N_20287);
nor U23207 (N_23207,N_20730,N_21593);
nand U23208 (N_23208,N_20365,N_22144);
nand U23209 (N_23209,N_21763,N_22447);
and U23210 (N_23210,N_21265,N_21192);
nor U23211 (N_23211,N_21262,N_21400);
and U23212 (N_23212,N_21234,N_20636);
and U23213 (N_23213,N_20685,N_20364);
nor U23214 (N_23214,N_20039,N_20907);
nand U23215 (N_23215,N_20743,N_21030);
nand U23216 (N_23216,N_21679,N_21308);
or U23217 (N_23217,N_21240,N_20630);
xor U23218 (N_23218,N_20197,N_21892);
xnor U23219 (N_23219,N_22381,N_22118);
nor U23220 (N_23220,N_20264,N_21708);
or U23221 (N_23221,N_21403,N_21875);
xnor U23222 (N_23222,N_20191,N_21833);
xnor U23223 (N_23223,N_20802,N_20144);
xor U23224 (N_23224,N_21461,N_22362);
or U23225 (N_23225,N_21397,N_21063);
or U23226 (N_23226,N_22163,N_21022);
xor U23227 (N_23227,N_20830,N_21777);
nand U23228 (N_23228,N_21726,N_20242);
and U23229 (N_23229,N_20990,N_22226);
nor U23230 (N_23230,N_21906,N_20598);
nor U23231 (N_23231,N_22434,N_21497);
or U23232 (N_23232,N_20610,N_20857);
nor U23233 (N_23233,N_22411,N_21302);
nand U23234 (N_23234,N_22157,N_20591);
or U23235 (N_23235,N_20058,N_20564);
nor U23236 (N_23236,N_22050,N_20309);
nor U23237 (N_23237,N_22320,N_20235);
nor U23238 (N_23238,N_20820,N_21754);
or U23239 (N_23239,N_21872,N_20539);
xnor U23240 (N_23240,N_20352,N_20377);
nand U23241 (N_23241,N_20038,N_20244);
or U23242 (N_23242,N_20046,N_20651);
or U23243 (N_23243,N_20876,N_21150);
and U23244 (N_23244,N_20294,N_21952);
or U23245 (N_23245,N_21112,N_21849);
and U23246 (N_23246,N_22032,N_21658);
and U23247 (N_23247,N_21111,N_20553);
nand U23248 (N_23248,N_22481,N_21834);
xor U23249 (N_23249,N_21396,N_20832);
nand U23250 (N_23250,N_21750,N_21368);
and U23251 (N_23251,N_21088,N_20252);
or U23252 (N_23252,N_22017,N_22439);
nor U23253 (N_23253,N_21206,N_21891);
nor U23254 (N_23254,N_21492,N_21910);
and U23255 (N_23255,N_20464,N_22031);
nand U23256 (N_23256,N_21973,N_21071);
and U23257 (N_23257,N_20293,N_21547);
or U23258 (N_23258,N_21986,N_20435);
or U23259 (N_23259,N_21635,N_21277);
or U23260 (N_23260,N_22087,N_20612);
nand U23261 (N_23261,N_22258,N_20019);
nor U23262 (N_23262,N_20373,N_20880);
and U23263 (N_23263,N_20524,N_20679);
or U23264 (N_23264,N_20858,N_20686);
nor U23265 (N_23265,N_20467,N_21883);
and U23266 (N_23266,N_21049,N_21061);
xor U23267 (N_23267,N_22035,N_21404);
nor U23268 (N_23268,N_20677,N_22262);
and U23269 (N_23269,N_20811,N_22399);
nor U23270 (N_23270,N_21839,N_20617);
or U23271 (N_23271,N_21744,N_20427);
nand U23272 (N_23272,N_22162,N_22045);
nand U23273 (N_23273,N_22242,N_21311);
nand U23274 (N_23274,N_21160,N_20133);
or U23275 (N_23275,N_20578,N_20673);
xor U23276 (N_23276,N_22041,N_20852);
xnor U23277 (N_23277,N_20952,N_20204);
or U23278 (N_23278,N_20270,N_22433);
and U23279 (N_23279,N_21911,N_22107);
nor U23280 (N_23280,N_21173,N_20937);
nand U23281 (N_23281,N_22093,N_21456);
and U23282 (N_23282,N_20459,N_20813);
or U23283 (N_23283,N_22224,N_21473);
and U23284 (N_23284,N_21520,N_20044);
nor U23285 (N_23285,N_21191,N_20642);
and U23286 (N_23286,N_21927,N_20214);
nand U23287 (N_23287,N_22011,N_21273);
nor U23288 (N_23288,N_22194,N_22305);
or U23289 (N_23289,N_20699,N_21616);
xor U23290 (N_23290,N_20652,N_20513);
nor U23291 (N_23291,N_22478,N_20166);
or U23292 (N_23292,N_21894,N_21137);
nand U23293 (N_23293,N_20411,N_20670);
or U23294 (N_23294,N_20606,N_22402);
xnor U23295 (N_23295,N_20106,N_20096);
or U23296 (N_23296,N_21909,N_21208);
xor U23297 (N_23297,N_20913,N_20984);
and U23298 (N_23298,N_21421,N_21611);
and U23299 (N_23299,N_20181,N_20138);
and U23300 (N_23300,N_20070,N_22084);
nand U23301 (N_23301,N_20935,N_21282);
and U23302 (N_23302,N_20265,N_20600);
nor U23303 (N_23303,N_20807,N_20972);
or U23304 (N_23304,N_22248,N_21882);
nand U23305 (N_23305,N_21739,N_22324);
or U23306 (N_23306,N_21427,N_20684);
nor U23307 (N_23307,N_21935,N_22193);
nand U23308 (N_23308,N_21554,N_21589);
nand U23309 (N_23309,N_20000,N_20744);
nor U23310 (N_23310,N_20009,N_20967);
nor U23311 (N_23311,N_22310,N_21923);
or U23312 (N_23312,N_20040,N_21255);
nor U23313 (N_23313,N_20335,N_21525);
and U23314 (N_23314,N_20100,N_21385);
nand U23315 (N_23315,N_21279,N_21930);
nand U23316 (N_23316,N_20998,N_21805);
or U23317 (N_23317,N_22269,N_22266);
nor U23318 (N_23318,N_21056,N_21981);
nand U23319 (N_23319,N_21453,N_21238);
nor U23320 (N_23320,N_21333,N_21377);
nand U23321 (N_23321,N_20574,N_20500);
nand U23322 (N_23322,N_20172,N_21571);
xor U23323 (N_23323,N_20279,N_21823);
and U23324 (N_23324,N_21816,N_21109);
and U23325 (N_23325,N_20566,N_21083);
nor U23326 (N_23326,N_20842,N_22400);
or U23327 (N_23327,N_22303,N_22088);
and U23328 (N_23328,N_21465,N_22314);
and U23329 (N_23329,N_20431,N_20769);
and U23330 (N_23330,N_21176,N_21357);
or U23331 (N_23331,N_21889,N_20498);
nand U23332 (N_23332,N_21068,N_20648);
and U23333 (N_23333,N_20349,N_21328);
nand U23334 (N_23334,N_22019,N_21182);
nor U23335 (N_23335,N_20341,N_21868);
or U23336 (N_23336,N_21597,N_21246);
or U23337 (N_23337,N_21854,N_21861);
nor U23338 (N_23338,N_20947,N_22121);
and U23339 (N_23339,N_20243,N_20750);
and U23340 (N_23340,N_20542,N_20712);
or U23341 (N_23341,N_22413,N_21470);
and U23342 (N_23342,N_21576,N_20519);
nand U23343 (N_23343,N_21230,N_20596);
or U23344 (N_23344,N_21668,N_21462);
and U23345 (N_23345,N_20538,N_20833);
and U23346 (N_23346,N_20218,N_22466);
or U23347 (N_23347,N_21003,N_21389);
xnor U23348 (N_23348,N_22109,N_20772);
and U23349 (N_23349,N_20577,N_21874);
nor U23350 (N_23350,N_21028,N_21136);
xnor U23351 (N_23351,N_21916,N_22416);
xor U23352 (N_23352,N_22264,N_21559);
and U23353 (N_23353,N_20105,N_21985);
or U23354 (N_23354,N_22170,N_22497);
or U23355 (N_23355,N_20416,N_21494);
nand U23356 (N_23356,N_22030,N_22034);
xnor U23357 (N_23357,N_21179,N_22286);
and U23358 (N_23358,N_21505,N_21915);
or U23359 (N_23359,N_22009,N_21038);
xnor U23360 (N_23360,N_21159,N_20599);
nor U23361 (N_23361,N_20536,N_21914);
nor U23362 (N_23362,N_21187,N_20738);
nand U23363 (N_23363,N_21503,N_21338);
and U23364 (N_23364,N_21512,N_21414);
nand U23365 (N_23365,N_21947,N_22062);
or U23366 (N_23366,N_21477,N_21784);
nand U23367 (N_23367,N_22465,N_21438);
or U23368 (N_23368,N_20230,N_21498);
nor U23369 (N_23369,N_22006,N_20774);
nor U23370 (N_23370,N_21529,N_20705);
nor U23371 (N_23371,N_21540,N_21285);
or U23372 (N_23372,N_22484,N_21633);
and U23373 (N_23373,N_21530,N_21591);
or U23374 (N_23374,N_20906,N_21976);
nand U23375 (N_23375,N_21799,N_20370);
nand U23376 (N_23376,N_20496,N_20299);
nand U23377 (N_23377,N_20177,N_20048);
or U23378 (N_23378,N_21037,N_21219);
or U23379 (N_23379,N_22365,N_22480);
nor U23380 (N_23380,N_21355,N_22448);
nor U23381 (N_23381,N_22155,N_22187);
and U23382 (N_23382,N_22482,N_21193);
nor U23383 (N_23383,N_20068,N_21100);
nor U23384 (N_23384,N_21422,N_22221);
or U23385 (N_23385,N_20126,N_21519);
nor U23386 (N_23386,N_21725,N_20095);
or U23387 (N_23387,N_21972,N_22159);
nand U23388 (N_23388,N_20361,N_21526);
nor U23389 (N_23389,N_20595,N_21837);
nand U23390 (N_23390,N_20136,N_20667);
and U23391 (N_23391,N_21081,N_20664);
or U23392 (N_23392,N_21139,N_20745);
and U23393 (N_23393,N_20247,N_22151);
and U23394 (N_23394,N_22080,N_20641);
and U23395 (N_23395,N_20272,N_22038);
nor U23396 (N_23396,N_21890,N_20261);
nor U23397 (N_23397,N_21604,N_20866);
and U23398 (N_23398,N_20851,N_21625);
and U23399 (N_23399,N_21740,N_21210);
nor U23400 (N_23400,N_22289,N_22000);
nand U23401 (N_23401,N_22043,N_20470);
nor U23402 (N_23402,N_20062,N_20728);
and U23403 (N_23403,N_21997,N_22095);
nand U23404 (N_23404,N_20053,N_21454);
nor U23405 (N_23405,N_22398,N_21110);
nor U23406 (N_23406,N_20517,N_22321);
nor U23407 (N_23407,N_22128,N_20688);
nor U23408 (N_23408,N_21395,N_21610);
nor U23409 (N_23409,N_21222,N_20732);
and U23410 (N_23410,N_21376,N_21581);
or U23411 (N_23411,N_21304,N_20859);
and U23412 (N_23412,N_21167,N_20154);
or U23413 (N_23413,N_21367,N_20502);
and U23414 (N_23414,N_21795,N_20550);
or U23415 (N_23415,N_20977,N_21800);
nor U23416 (N_23416,N_22117,N_20659);
nand U23417 (N_23417,N_21895,N_21263);
or U23418 (N_23418,N_22042,N_22281);
nand U23419 (N_23419,N_20702,N_20006);
or U23420 (N_23420,N_21859,N_22498);
nor U23421 (N_23421,N_20801,N_20675);
or U23422 (N_23422,N_22494,N_21010);
nand U23423 (N_23423,N_20809,N_21629);
nand U23424 (N_23424,N_22178,N_21055);
or U23425 (N_23425,N_21501,N_21275);
nand U23426 (N_23426,N_22367,N_21983);
nand U23427 (N_23427,N_22007,N_20803);
nor U23428 (N_23428,N_21639,N_20310);
or U23429 (N_23429,N_20950,N_21599);
nand U23430 (N_23430,N_21020,N_21919);
nor U23431 (N_23431,N_20597,N_20632);
and U23432 (N_23432,N_22309,N_20267);
nor U23433 (N_23433,N_21745,N_20192);
nor U23434 (N_23434,N_20079,N_20510);
nand U23435 (N_23435,N_22044,N_20369);
nor U23436 (N_23436,N_21977,N_22014);
nor U23437 (N_23437,N_21749,N_21681);
nor U23438 (N_23438,N_22420,N_22308);
nand U23439 (N_23439,N_20362,N_22369);
nor U23440 (N_23440,N_21647,N_21955);
and U23441 (N_23441,N_20656,N_20822);
and U23442 (N_23442,N_22201,N_22383);
nor U23443 (N_23443,N_21146,N_22285);
nand U23444 (N_23444,N_22384,N_20437);
and U23445 (N_23445,N_21767,N_20846);
and U23446 (N_23446,N_22299,N_22133);
nor U23447 (N_23447,N_20746,N_21464);
nand U23448 (N_23448,N_20714,N_22137);
or U23449 (N_23449,N_21881,N_21119);
nand U23450 (N_23450,N_21822,N_22124);
nand U23451 (N_23451,N_21577,N_21608);
nand U23452 (N_23452,N_21957,N_20442);
or U23453 (N_23453,N_20420,N_21455);
and U23454 (N_23454,N_22290,N_21108);
or U23455 (N_23455,N_21614,N_20451);
xor U23456 (N_23456,N_21888,N_20449);
nor U23457 (N_23457,N_21770,N_22203);
or U23458 (N_23458,N_22410,N_21025);
and U23459 (N_23459,N_20506,N_21381);
or U23460 (N_23460,N_21553,N_20621);
nand U23461 (N_23461,N_21579,N_20691);
or U23462 (N_23462,N_21709,N_21998);
nand U23463 (N_23463,N_21736,N_20931);
and U23464 (N_23464,N_22101,N_21762);
and U23465 (N_23465,N_21185,N_20625);
nand U23466 (N_23466,N_21867,N_21113);
nor U23467 (N_23467,N_20182,N_20959);
xnor U23468 (N_23468,N_20433,N_20148);
nand U23469 (N_23469,N_20180,N_21452);
nand U23470 (N_23470,N_22021,N_20073);
nand U23471 (N_23471,N_21491,N_22382);
or U23472 (N_23472,N_20249,N_20874);
nand U23473 (N_23473,N_20475,N_22135);
or U23474 (N_23474,N_20323,N_20844);
nand U23475 (N_23475,N_20605,N_20394);
nand U23476 (N_23476,N_21730,N_21878);
xor U23477 (N_23477,N_20288,N_20795);
nand U23478 (N_23478,N_22316,N_21690);
or U23479 (N_23479,N_21371,N_21363);
nor U23480 (N_23480,N_20090,N_20134);
nor U23481 (N_23481,N_22138,N_22003);
nand U23482 (N_23482,N_21848,N_20626);
and U23483 (N_23483,N_21215,N_20929);
nand U23484 (N_23484,N_21466,N_22123);
or U23485 (N_23485,N_20452,N_20484);
nand U23486 (N_23486,N_20041,N_20462);
and U23487 (N_23487,N_21340,N_20071);
or U23488 (N_23488,N_20682,N_20473);
xor U23489 (N_23489,N_20140,N_22166);
xor U23490 (N_23490,N_22169,N_22349);
nand U23491 (N_23491,N_20425,N_21393);
nor U23492 (N_23492,N_21556,N_22485);
nor U23493 (N_23493,N_21732,N_20423);
and U23494 (N_23494,N_20547,N_22274);
nor U23495 (N_23495,N_21342,N_21116);
xnor U23496 (N_23496,N_21294,N_21722);
and U23497 (N_23497,N_21095,N_20532);
nand U23498 (N_23498,N_21753,N_21463);
nor U23499 (N_23499,N_22120,N_20185);
xor U23500 (N_23500,N_21325,N_21974);
xor U23501 (N_23501,N_21425,N_20569);
or U23502 (N_23502,N_20665,N_21184);
and U23503 (N_23503,N_20305,N_21691);
and U23504 (N_23504,N_21587,N_21527);
nand U23505 (N_23505,N_21177,N_21537);
or U23506 (N_23506,N_21266,N_21850);
nand U23507 (N_23507,N_22238,N_21607);
or U23508 (N_23508,N_20092,N_22016);
or U23509 (N_23509,N_22231,N_20753);
nand U23510 (N_23510,N_21687,N_21148);
nor U23511 (N_23511,N_20495,N_20224);
and U23512 (N_23512,N_20819,N_21831);
nor U23513 (N_23513,N_20189,N_20297);
nand U23514 (N_23514,N_20150,N_22429);
and U23515 (N_23515,N_22143,N_20870);
or U23516 (N_23516,N_20810,N_22197);
nand U23517 (N_23517,N_20319,N_22385);
nand U23518 (N_23518,N_22139,N_21092);
or U23519 (N_23519,N_22282,N_20587);
and U23520 (N_23520,N_21166,N_20099);
nor U23521 (N_23521,N_22146,N_20962);
or U23522 (N_23522,N_21748,N_22459);
nor U23523 (N_23523,N_21688,N_20386);
nor U23524 (N_23524,N_20742,N_22431);
nand U23525 (N_23525,N_20176,N_21014);
or U23526 (N_23526,N_20005,N_20909);
xor U23527 (N_23527,N_21072,N_20724);
or U23528 (N_23528,N_22304,N_21958);
and U23529 (N_23529,N_20295,N_21545);
and U23530 (N_23530,N_20581,N_20301);
or U23531 (N_23531,N_20002,N_20075);
or U23532 (N_23532,N_21640,N_20016);
and U23533 (N_23533,N_21601,N_21359);
or U23534 (N_23534,N_21089,N_20782);
and U23535 (N_23535,N_21514,N_20603);
nand U23536 (N_23536,N_22256,N_20315);
and U23537 (N_23537,N_21925,N_20708);
and U23538 (N_23538,N_21810,N_22259);
or U23539 (N_23539,N_21310,N_21769);
xor U23540 (N_23540,N_21305,N_20065);
and U23541 (N_23541,N_21077,N_21314);
nand U23542 (N_23542,N_22114,N_21439);
and U23543 (N_23543,N_20499,N_21469);
and U23544 (N_23544,N_20918,N_21413);
nor U23545 (N_23545,N_21944,N_22337);
or U23546 (N_23546,N_21053,N_21487);
and U23547 (N_23547,N_22070,N_21181);
and U23548 (N_23548,N_21096,N_22364);
and U23549 (N_23549,N_21734,N_20465);
or U23550 (N_23550,N_21907,N_21374);
nand U23551 (N_23551,N_21321,N_20944);
and U23552 (N_23552,N_21798,N_20343);
or U23553 (N_23553,N_20132,N_22333);
xnor U23554 (N_23554,N_20419,N_21129);
nand U23555 (N_23555,N_20658,N_20861);
xor U23556 (N_23556,N_20429,N_20590);
and U23557 (N_23557,N_22358,N_22489);
nor U23558 (N_23558,N_21186,N_22244);
nor U23559 (N_23559,N_21154,N_21542);
and U23560 (N_23560,N_21928,N_21513);
and U23561 (N_23561,N_22113,N_21628);
xor U23562 (N_23562,N_20974,N_21291);
or U23563 (N_23563,N_21863,N_20312);
nand U23564 (N_23564,N_22306,N_20121);
nand U23565 (N_23565,N_22217,N_21866);
nand U23566 (N_23566,N_21164,N_21563);
and U23567 (N_23567,N_22218,N_21343);
nor U23568 (N_23568,N_21224,N_21807);
nand U23569 (N_23569,N_20388,N_20903);
xnor U23570 (N_23570,N_20331,N_21515);
nor U23571 (N_23571,N_21680,N_20837);
and U23572 (N_23572,N_21598,N_20582);
and U23573 (N_23573,N_20222,N_21920);
or U23574 (N_23574,N_21676,N_20043);
nor U23575 (N_23575,N_20254,N_20737);
or U23576 (N_23576,N_22059,N_20213);
or U23577 (N_23577,N_21780,N_21380);
nor U23578 (N_23578,N_21694,N_21147);
xnor U23579 (N_23579,N_22092,N_20396);
or U23580 (N_23580,N_21076,N_20372);
nor U23581 (N_23581,N_20256,N_20894);
nor U23582 (N_23582,N_21561,N_21645);
or U23583 (N_23583,N_22326,N_21098);
or U23584 (N_23584,N_22370,N_20766);
xnor U23585 (N_23585,N_20014,N_20446);
and U23586 (N_23586,N_20316,N_20573);
nor U23587 (N_23587,N_21085,N_21783);
nand U23588 (N_23588,N_21641,N_20872);
nand U23589 (N_23589,N_22397,N_20400);
nand U23590 (N_23590,N_22278,N_20421);
xor U23591 (N_23591,N_21858,N_21992);
or U23592 (N_23592,N_20619,N_21700);
and U23593 (N_23593,N_20072,N_20700);
and U23594 (N_23594,N_20924,N_22452);
nor U23595 (N_23595,N_21502,N_21251);
nand U23596 (N_23596,N_21365,N_20404);
and U23597 (N_23597,N_21420,N_21029);
or U23598 (N_23598,N_21642,N_20015);
xnor U23599 (N_23599,N_20412,N_22190);
nand U23600 (N_23600,N_21104,N_22039);
and U23601 (N_23601,N_20424,N_21281);
or U23602 (N_23602,N_21412,N_21093);
nand U23603 (N_23603,N_22110,N_22127);
or U23604 (N_23604,N_22077,N_20474);
xor U23605 (N_23605,N_21843,N_22072);
or U23606 (N_23606,N_21248,N_21245);
xnor U23607 (N_23607,N_22102,N_21019);
and U23608 (N_23608,N_21408,N_20007);
or U23609 (N_23609,N_21045,N_21569);
nand U23610 (N_23610,N_21142,N_21752);
and U23611 (N_23611,N_20919,N_22302);
nor U23612 (N_23612,N_20963,N_20275);
nand U23613 (N_23613,N_21785,N_20198);
nand U23614 (N_23614,N_20647,N_21993);
nand U23615 (N_23615,N_21151,N_21949);
or U23616 (N_23616,N_20201,N_20008);
xor U23617 (N_23617,N_20823,N_20757);
and U23618 (N_23618,N_20186,N_21592);
and U23619 (N_23619,N_21450,N_21620);
and U23620 (N_23620,N_20650,N_21879);
and U23621 (N_23621,N_21402,N_22311);
nor U23622 (N_23622,N_20440,N_21485);
or U23623 (N_23623,N_22205,N_22313);
xnor U23624 (N_23624,N_21190,N_22188);
nand U23625 (N_23625,N_20865,N_21296);
and U23626 (N_23626,N_20911,N_20672);
or U23627 (N_23627,N_21124,N_20205);
and U23628 (N_23628,N_20585,N_21896);
nor U23629 (N_23629,N_20873,N_20540);
and U23630 (N_23630,N_21168,N_21074);
and U23631 (N_23631,N_22026,N_20178);
nand U23632 (N_23632,N_22154,N_20292);
nand U23633 (N_23633,N_22460,N_20683);
nand U23634 (N_23634,N_22136,N_21231);
nor U23635 (N_23635,N_21522,N_20562);
nand U23636 (N_23636,N_20896,N_20748);
nand U23637 (N_23637,N_20775,N_21900);
and U23638 (N_23638,N_20238,N_20497);
xnor U23639 (N_23639,N_20028,N_21324);
nor U23640 (N_23640,N_21127,N_20320);
nor U23641 (N_23641,N_21317,N_20357);
and U23642 (N_23642,N_21011,N_20781);
nor U23643 (N_23643,N_20957,N_21811);
and U23644 (N_23644,N_21254,N_21152);
or U23645 (N_23645,N_20142,N_22432);
nand U23646 (N_23646,N_22212,N_20796);
nand U23647 (N_23647,N_21237,N_21226);
and U23648 (N_23648,N_21229,N_21948);
or U23649 (N_23649,N_22368,N_20387);
or U23650 (N_23650,N_21655,N_21706);
xnor U23651 (N_23651,N_20965,N_20322);
and U23652 (N_23652,N_21495,N_21521);
and U23653 (N_23653,N_20093,N_20381);
nor U23654 (N_23654,N_21118,N_22160);
nor U23655 (N_23655,N_20958,N_22283);
nor U23656 (N_23656,N_20385,N_20531);
nor U23657 (N_23657,N_20193,N_21351);
or U23658 (N_23658,N_22293,N_21419);
and U23659 (N_23659,N_20225,N_20165);
or U23660 (N_23660,N_20867,N_20544);
nand U23661 (N_23661,N_22463,N_20821);
nor U23662 (N_23662,N_20734,N_22180);
or U23663 (N_23663,N_22176,N_20789);
nand U23664 (N_23664,N_22158,N_21320);
nand U23665 (N_23665,N_21876,N_20393);
nand U23666 (N_23666,N_20551,N_21824);
and U23667 (N_23667,N_22348,N_21388);
nor U23668 (N_23668,N_20111,N_21283);
xor U23669 (N_23669,N_21678,N_21274);
nand U23670 (N_23670,N_20787,N_21902);
or U23671 (N_23671,N_22387,N_20146);
nand U23672 (N_23672,N_20351,N_22105);
nand U23673 (N_23673,N_22284,N_22064);
and U23674 (N_23674,N_20227,N_22473);
and U23675 (N_23675,N_20125,N_21594);
or U23676 (N_23676,N_22425,N_21775);
and U23677 (N_23677,N_21982,N_21429);
nor U23678 (N_23678,N_21153,N_21078);
and U23679 (N_23679,N_20276,N_20583);
and U23680 (N_23680,N_21939,N_20202);
nor U23681 (N_23681,N_20228,N_21002);
or U23682 (N_23682,N_20661,N_22322);
xnor U23683 (N_23683,N_21280,N_21270);
and U23684 (N_23684,N_20403,N_21613);
xnor U23685 (N_23685,N_20390,N_21309);
and U23686 (N_23686,N_20643,N_20245);
xor U23687 (N_23687,N_20761,N_21677);
or U23688 (N_23688,N_20405,N_20012);
and U23689 (N_23689,N_21090,N_21590);
nor U23690 (N_23690,N_21970,N_20330);
nand U23691 (N_23691,N_20280,N_20951);
and U23692 (N_23692,N_22344,N_20441);
nand U23693 (N_23693,N_20646,N_20663);
and U23694 (N_23694,N_20457,N_21360);
xnor U23695 (N_23695,N_22338,N_21572);
and U23696 (N_23696,N_20816,N_20780);
nor U23697 (N_23697,N_20703,N_21200);
nor U23698 (N_23698,N_20633,N_20026);
xnor U23699 (N_23699,N_20456,N_20516);
and U23700 (N_23700,N_22457,N_22291);
nand U23701 (N_23701,N_21703,N_22150);
nand U23702 (N_23702,N_22060,N_20839);
nor U23703 (N_23703,N_20565,N_22295);
and U23704 (N_23704,N_22456,N_20898);
or U23705 (N_23705,N_21989,N_21065);
nor U23706 (N_23706,N_20843,N_20078);
and U23707 (N_23707,N_20943,N_21322);
nor U23708 (N_23708,N_21012,N_20339);
and U23709 (N_23709,N_22004,N_22406);
and U23710 (N_23710,N_21471,N_22015);
nor U23711 (N_23711,N_20196,N_22179);
nor U23712 (N_23712,N_20904,N_20970);
nand U23713 (N_23713,N_20480,N_21560);
nand U23714 (N_23714,N_22174,N_20088);
and U23715 (N_23715,N_20927,N_21596);
xnor U23716 (N_23716,N_20631,N_22354);
or U23717 (N_23717,N_20188,N_21818);
and U23718 (N_23718,N_20141,N_21199);
nand U23719 (N_23719,N_21912,N_21130);
nand U23720 (N_23720,N_20206,N_22329);
nor U23721 (N_23721,N_20052,N_21220);
and U23722 (N_23722,N_20528,N_21383);
nand U23723 (N_23723,N_22412,N_20639);
or U23724 (N_23724,N_20328,N_21922);
and U23725 (N_23725,N_20933,N_21711);
or U23726 (N_23726,N_21671,N_20307);
nand U23727 (N_23727,N_20776,N_21021);
nand U23728 (N_23728,N_20220,N_20494);
and U23729 (N_23729,N_20635,N_21728);
nand U23730 (N_23730,N_21418,N_22388);
and U23731 (N_23731,N_21239,N_21046);
xor U23732 (N_23732,N_21023,N_20389);
nor U23733 (N_23733,N_21548,N_22471);
nor U23734 (N_23734,N_20697,N_20855);
nand U23735 (N_23735,N_22392,N_21375);
xor U23736 (N_23736,N_21361,N_21673);
and U23737 (N_23737,N_20314,N_21293);
xor U23738 (N_23738,N_21567,N_20589);
nand U23739 (N_23739,N_22423,N_21832);
nor U23740 (N_23740,N_20969,N_21954);
or U23741 (N_23741,N_20200,N_21458);
and U23742 (N_23742,N_21288,N_20726);
nor U23743 (N_23743,N_21621,N_20260);
and U23744 (N_23744,N_20376,N_22164);
xor U23745 (N_23745,N_20616,N_20868);
nand U23746 (N_23746,N_22223,N_22012);
and U23747 (N_23747,N_20115,N_20767);
and U23748 (N_23748,N_21665,N_20914);
or U23749 (N_23749,N_21476,N_21443);
and U23750 (N_23750,N_21088,N_20621);
and U23751 (N_23751,N_20083,N_20160);
xnor U23752 (N_23752,N_20574,N_20689);
nand U23753 (N_23753,N_20826,N_20494);
nor U23754 (N_23754,N_20717,N_20237);
nand U23755 (N_23755,N_21951,N_20931);
and U23756 (N_23756,N_22234,N_21113);
nor U23757 (N_23757,N_20905,N_20131);
nand U23758 (N_23758,N_20364,N_20769);
nor U23759 (N_23759,N_21822,N_21869);
and U23760 (N_23760,N_20197,N_20099);
and U23761 (N_23761,N_20074,N_20172);
nand U23762 (N_23762,N_21244,N_21076);
nor U23763 (N_23763,N_20372,N_20147);
or U23764 (N_23764,N_20191,N_22282);
or U23765 (N_23765,N_21061,N_20463);
nor U23766 (N_23766,N_20545,N_21381);
or U23767 (N_23767,N_21733,N_20390);
or U23768 (N_23768,N_20649,N_22413);
and U23769 (N_23769,N_21044,N_20916);
nand U23770 (N_23770,N_21044,N_20191);
nand U23771 (N_23771,N_21662,N_21622);
xnor U23772 (N_23772,N_21533,N_20547);
nand U23773 (N_23773,N_22050,N_21429);
xnor U23774 (N_23774,N_22135,N_20459);
xnor U23775 (N_23775,N_20739,N_22401);
nor U23776 (N_23776,N_21304,N_20995);
nand U23777 (N_23777,N_22157,N_20547);
nor U23778 (N_23778,N_21927,N_20944);
nor U23779 (N_23779,N_21727,N_21808);
nor U23780 (N_23780,N_21073,N_21402);
nand U23781 (N_23781,N_21772,N_22102);
or U23782 (N_23782,N_20244,N_20717);
nor U23783 (N_23783,N_21944,N_21249);
xor U23784 (N_23784,N_20854,N_22021);
nor U23785 (N_23785,N_21792,N_20314);
xor U23786 (N_23786,N_22104,N_20645);
or U23787 (N_23787,N_22235,N_21815);
nand U23788 (N_23788,N_20655,N_20300);
nor U23789 (N_23789,N_20148,N_20790);
nand U23790 (N_23790,N_21953,N_20197);
nor U23791 (N_23791,N_22047,N_22461);
or U23792 (N_23792,N_21663,N_20713);
or U23793 (N_23793,N_21329,N_20557);
or U23794 (N_23794,N_20229,N_21502);
or U23795 (N_23795,N_22005,N_20493);
nand U23796 (N_23796,N_21336,N_22298);
nor U23797 (N_23797,N_22166,N_22249);
nor U23798 (N_23798,N_22448,N_21175);
nand U23799 (N_23799,N_21844,N_21125);
nand U23800 (N_23800,N_20117,N_22402);
and U23801 (N_23801,N_20401,N_20533);
and U23802 (N_23802,N_21490,N_21480);
nand U23803 (N_23803,N_20888,N_21901);
nand U23804 (N_23804,N_21203,N_21615);
or U23805 (N_23805,N_21701,N_20793);
xor U23806 (N_23806,N_20702,N_22166);
nand U23807 (N_23807,N_22135,N_21722);
nor U23808 (N_23808,N_20724,N_21066);
nand U23809 (N_23809,N_22281,N_22395);
or U23810 (N_23810,N_20969,N_20088);
nor U23811 (N_23811,N_20833,N_21824);
or U23812 (N_23812,N_20542,N_21071);
or U23813 (N_23813,N_21764,N_21934);
nand U23814 (N_23814,N_20038,N_22157);
and U23815 (N_23815,N_20358,N_20370);
or U23816 (N_23816,N_21210,N_20759);
nand U23817 (N_23817,N_20457,N_21679);
nand U23818 (N_23818,N_21187,N_22029);
nor U23819 (N_23819,N_21495,N_20746);
xnor U23820 (N_23820,N_20778,N_21515);
nor U23821 (N_23821,N_20562,N_22431);
nor U23822 (N_23822,N_21123,N_20866);
or U23823 (N_23823,N_21327,N_21861);
nand U23824 (N_23824,N_22120,N_21482);
xnor U23825 (N_23825,N_20923,N_20011);
xor U23826 (N_23826,N_21912,N_20556);
nand U23827 (N_23827,N_22443,N_20472);
nand U23828 (N_23828,N_22428,N_22346);
xor U23829 (N_23829,N_20327,N_21741);
nor U23830 (N_23830,N_20507,N_21377);
nor U23831 (N_23831,N_22454,N_22176);
or U23832 (N_23832,N_20218,N_22380);
nand U23833 (N_23833,N_21549,N_20144);
nand U23834 (N_23834,N_21203,N_21394);
and U23835 (N_23835,N_22022,N_20252);
nor U23836 (N_23836,N_21388,N_22389);
nand U23837 (N_23837,N_22085,N_22408);
nor U23838 (N_23838,N_22257,N_22344);
xnor U23839 (N_23839,N_22460,N_20756);
nor U23840 (N_23840,N_20884,N_21815);
xnor U23841 (N_23841,N_21008,N_20273);
and U23842 (N_23842,N_21375,N_20894);
and U23843 (N_23843,N_21073,N_21010);
and U23844 (N_23844,N_20254,N_21527);
or U23845 (N_23845,N_20995,N_20628);
or U23846 (N_23846,N_22118,N_21634);
nand U23847 (N_23847,N_22441,N_20725);
and U23848 (N_23848,N_21780,N_21673);
nor U23849 (N_23849,N_20095,N_20692);
nand U23850 (N_23850,N_21176,N_21917);
nor U23851 (N_23851,N_21427,N_21315);
xor U23852 (N_23852,N_22211,N_21018);
and U23853 (N_23853,N_20816,N_21646);
and U23854 (N_23854,N_20533,N_20629);
nor U23855 (N_23855,N_21301,N_21855);
nand U23856 (N_23856,N_20749,N_21362);
nor U23857 (N_23857,N_20152,N_22406);
xnor U23858 (N_23858,N_20998,N_20465);
or U23859 (N_23859,N_21930,N_21510);
nand U23860 (N_23860,N_20665,N_21867);
and U23861 (N_23861,N_21056,N_21556);
nand U23862 (N_23862,N_22337,N_21010);
nand U23863 (N_23863,N_21107,N_21043);
and U23864 (N_23864,N_22423,N_20476);
or U23865 (N_23865,N_20208,N_21567);
and U23866 (N_23866,N_20164,N_21716);
or U23867 (N_23867,N_22022,N_20232);
nand U23868 (N_23868,N_21595,N_22379);
nand U23869 (N_23869,N_21533,N_21313);
xnor U23870 (N_23870,N_22087,N_22480);
and U23871 (N_23871,N_21480,N_20440);
nor U23872 (N_23872,N_20548,N_21349);
nor U23873 (N_23873,N_21359,N_20960);
or U23874 (N_23874,N_21944,N_22000);
xnor U23875 (N_23875,N_22298,N_21801);
nor U23876 (N_23876,N_21374,N_22352);
nand U23877 (N_23877,N_20520,N_21061);
nand U23878 (N_23878,N_20797,N_21391);
or U23879 (N_23879,N_20168,N_21833);
and U23880 (N_23880,N_20013,N_20106);
and U23881 (N_23881,N_20971,N_20159);
and U23882 (N_23882,N_21511,N_22144);
and U23883 (N_23883,N_22020,N_20150);
nor U23884 (N_23884,N_20792,N_20553);
nand U23885 (N_23885,N_21098,N_21442);
nor U23886 (N_23886,N_21466,N_22020);
nor U23887 (N_23887,N_21543,N_20324);
and U23888 (N_23888,N_20673,N_21078);
nand U23889 (N_23889,N_22248,N_22173);
or U23890 (N_23890,N_20255,N_20478);
xnor U23891 (N_23891,N_20991,N_20875);
and U23892 (N_23892,N_22097,N_20635);
and U23893 (N_23893,N_21926,N_21483);
nand U23894 (N_23894,N_21104,N_22216);
nand U23895 (N_23895,N_21689,N_21653);
nor U23896 (N_23896,N_20910,N_20921);
or U23897 (N_23897,N_21980,N_20653);
nand U23898 (N_23898,N_21983,N_22355);
and U23899 (N_23899,N_20253,N_20164);
or U23900 (N_23900,N_21660,N_20425);
and U23901 (N_23901,N_20222,N_21739);
nor U23902 (N_23902,N_21163,N_21478);
nand U23903 (N_23903,N_20390,N_21094);
or U23904 (N_23904,N_20995,N_20434);
and U23905 (N_23905,N_20113,N_21914);
or U23906 (N_23906,N_22047,N_21786);
nor U23907 (N_23907,N_20007,N_20336);
nor U23908 (N_23908,N_20268,N_22431);
and U23909 (N_23909,N_21696,N_22250);
or U23910 (N_23910,N_20401,N_22370);
nor U23911 (N_23911,N_21051,N_21068);
or U23912 (N_23912,N_20071,N_20385);
nand U23913 (N_23913,N_21481,N_20143);
or U23914 (N_23914,N_20381,N_22107);
and U23915 (N_23915,N_20608,N_22005);
nor U23916 (N_23916,N_20161,N_22066);
or U23917 (N_23917,N_21307,N_20026);
xor U23918 (N_23918,N_20414,N_22282);
and U23919 (N_23919,N_22149,N_21191);
or U23920 (N_23920,N_21396,N_20976);
nand U23921 (N_23921,N_21383,N_20382);
xnor U23922 (N_23922,N_21421,N_21383);
nor U23923 (N_23923,N_21331,N_21314);
nor U23924 (N_23924,N_21603,N_22426);
and U23925 (N_23925,N_20798,N_21010);
or U23926 (N_23926,N_20781,N_20851);
nor U23927 (N_23927,N_21023,N_21245);
nor U23928 (N_23928,N_20468,N_20116);
and U23929 (N_23929,N_20864,N_20450);
nand U23930 (N_23930,N_20025,N_21814);
nor U23931 (N_23931,N_20867,N_21472);
and U23932 (N_23932,N_21981,N_20291);
or U23933 (N_23933,N_20515,N_22169);
nand U23934 (N_23934,N_22224,N_21678);
xor U23935 (N_23935,N_21348,N_21953);
and U23936 (N_23936,N_20250,N_21369);
or U23937 (N_23937,N_21313,N_20039);
and U23938 (N_23938,N_21935,N_21215);
and U23939 (N_23939,N_22014,N_21691);
nand U23940 (N_23940,N_22267,N_22378);
nand U23941 (N_23941,N_21220,N_20399);
nand U23942 (N_23942,N_22201,N_20177);
and U23943 (N_23943,N_22142,N_21764);
xnor U23944 (N_23944,N_20083,N_20270);
or U23945 (N_23945,N_21954,N_20913);
and U23946 (N_23946,N_20434,N_20986);
nand U23947 (N_23947,N_22003,N_22155);
and U23948 (N_23948,N_21223,N_22110);
nor U23949 (N_23949,N_20324,N_20858);
nand U23950 (N_23950,N_20399,N_21773);
xnor U23951 (N_23951,N_21881,N_22057);
nor U23952 (N_23952,N_20277,N_21843);
or U23953 (N_23953,N_20223,N_21467);
xnor U23954 (N_23954,N_20044,N_21446);
or U23955 (N_23955,N_22141,N_20990);
or U23956 (N_23956,N_22307,N_20153);
nor U23957 (N_23957,N_20065,N_22482);
and U23958 (N_23958,N_21920,N_20676);
nand U23959 (N_23959,N_22184,N_20251);
or U23960 (N_23960,N_21230,N_21417);
nor U23961 (N_23961,N_20549,N_21446);
or U23962 (N_23962,N_20390,N_20054);
or U23963 (N_23963,N_22157,N_20615);
and U23964 (N_23964,N_21771,N_20496);
and U23965 (N_23965,N_22393,N_22316);
nor U23966 (N_23966,N_21050,N_21663);
or U23967 (N_23967,N_20726,N_20241);
nor U23968 (N_23968,N_22045,N_22268);
nor U23969 (N_23969,N_20156,N_22337);
nor U23970 (N_23970,N_22382,N_20642);
nand U23971 (N_23971,N_21982,N_22146);
and U23972 (N_23972,N_20424,N_20724);
nor U23973 (N_23973,N_21020,N_20416);
nand U23974 (N_23974,N_21061,N_22471);
or U23975 (N_23975,N_21024,N_21576);
nand U23976 (N_23976,N_20176,N_22081);
nand U23977 (N_23977,N_20642,N_21967);
or U23978 (N_23978,N_21230,N_21883);
nand U23979 (N_23979,N_20564,N_20491);
or U23980 (N_23980,N_22413,N_22457);
nor U23981 (N_23981,N_22371,N_20986);
or U23982 (N_23982,N_21124,N_22174);
nor U23983 (N_23983,N_20412,N_22311);
nor U23984 (N_23984,N_20063,N_20440);
nand U23985 (N_23985,N_21744,N_21434);
and U23986 (N_23986,N_21837,N_20350);
nand U23987 (N_23987,N_21585,N_21776);
nand U23988 (N_23988,N_20152,N_20678);
and U23989 (N_23989,N_21249,N_20865);
xor U23990 (N_23990,N_21191,N_21436);
and U23991 (N_23991,N_20193,N_20174);
nor U23992 (N_23992,N_21127,N_20437);
and U23993 (N_23993,N_20081,N_20369);
nand U23994 (N_23994,N_22223,N_20283);
or U23995 (N_23995,N_21524,N_21156);
nor U23996 (N_23996,N_20808,N_21425);
xor U23997 (N_23997,N_22371,N_20180);
and U23998 (N_23998,N_21800,N_21888);
or U23999 (N_23999,N_20142,N_20070);
nand U24000 (N_24000,N_20589,N_20424);
nand U24001 (N_24001,N_20231,N_21920);
nor U24002 (N_24002,N_21979,N_20235);
nor U24003 (N_24003,N_20702,N_21494);
nor U24004 (N_24004,N_22142,N_20489);
or U24005 (N_24005,N_20791,N_20012);
nor U24006 (N_24006,N_22227,N_21236);
and U24007 (N_24007,N_22295,N_21461);
nor U24008 (N_24008,N_21616,N_20958);
nand U24009 (N_24009,N_21626,N_20509);
nand U24010 (N_24010,N_20673,N_21630);
and U24011 (N_24011,N_20894,N_21278);
nand U24012 (N_24012,N_21118,N_21863);
xor U24013 (N_24013,N_21477,N_20570);
or U24014 (N_24014,N_20372,N_20169);
nor U24015 (N_24015,N_21257,N_21252);
or U24016 (N_24016,N_21104,N_22384);
nor U24017 (N_24017,N_20781,N_21573);
and U24018 (N_24018,N_22449,N_20795);
nand U24019 (N_24019,N_21062,N_21448);
and U24020 (N_24020,N_21206,N_20100);
or U24021 (N_24021,N_22431,N_22142);
nor U24022 (N_24022,N_21856,N_21762);
xor U24023 (N_24023,N_20062,N_22037);
and U24024 (N_24024,N_21151,N_20595);
or U24025 (N_24025,N_20148,N_21792);
and U24026 (N_24026,N_20886,N_21483);
and U24027 (N_24027,N_21585,N_21927);
or U24028 (N_24028,N_20607,N_20624);
or U24029 (N_24029,N_22257,N_20974);
and U24030 (N_24030,N_21474,N_20865);
xnor U24031 (N_24031,N_20134,N_20047);
nor U24032 (N_24032,N_22438,N_22114);
and U24033 (N_24033,N_21187,N_22181);
nand U24034 (N_24034,N_20260,N_20752);
or U24035 (N_24035,N_22318,N_21928);
nand U24036 (N_24036,N_20238,N_21554);
nor U24037 (N_24037,N_20254,N_21288);
or U24038 (N_24038,N_21167,N_21917);
or U24039 (N_24039,N_20512,N_20347);
nand U24040 (N_24040,N_22215,N_21374);
nor U24041 (N_24041,N_21204,N_20965);
or U24042 (N_24042,N_21735,N_21141);
nor U24043 (N_24043,N_20357,N_22172);
or U24044 (N_24044,N_20796,N_20913);
and U24045 (N_24045,N_20379,N_22409);
and U24046 (N_24046,N_20802,N_21694);
and U24047 (N_24047,N_21478,N_21675);
and U24048 (N_24048,N_20396,N_20053);
nand U24049 (N_24049,N_20711,N_21113);
or U24050 (N_24050,N_22062,N_22207);
nand U24051 (N_24051,N_21776,N_21923);
and U24052 (N_24052,N_20661,N_20876);
xnor U24053 (N_24053,N_21798,N_21037);
nand U24054 (N_24054,N_20436,N_21761);
or U24055 (N_24055,N_21722,N_21457);
nand U24056 (N_24056,N_22320,N_21285);
nand U24057 (N_24057,N_21153,N_20033);
or U24058 (N_24058,N_21085,N_20998);
nand U24059 (N_24059,N_21526,N_21348);
xor U24060 (N_24060,N_21696,N_20229);
nand U24061 (N_24061,N_21449,N_20332);
or U24062 (N_24062,N_21620,N_20704);
nand U24063 (N_24063,N_22491,N_20332);
nor U24064 (N_24064,N_22016,N_21498);
and U24065 (N_24065,N_20047,N_21518);
nor U24066 (N_24066,N_21508,N_21609);
nand U24067 (N_24067,N_20980,N_22361);
and U24068 (N_24068,N_21865,N_21329);
nand U24069 (N_24069,N_20688,N_21081);
xnor U24070 (N_24070,N_20775,N_20920);
and U24071 (N_24071,N_20168,N_22217);
xnor U24072 (N_24072,N_21015,N_21456);
nand U24073 (N_24073,N_21478,N_20793);
nor U24074 (N_24074,N_20257,N_21689);
xor U24075 (N_24075,N_21389,N_21943);
nor U24076 (N_24076,N_21946,N_20110);
xor U24077 (N_24077,N_21412,N_20706);
and U24078 (N_24078,N_20021,N_21453);
nand U24079 (N_24079,N_22149,N_21268);
and U24080 (N_24080,N_21228,N_22246);
or U24081 (N_24081,N_21561,N_20372);
and U24082 (N_24082,N_21140,N_20352);
and U24083 (N_24083,N_21614,N_21972);
nor U24084 (N_24084,N_21380,N_21234);
or U24085 (N_24085,N_22176,N_21862);
and U24086 (N_24086,N_21870,N_21487);
and U24087 (N_24087,N_20477,N_21810);
nor U24088 (N_24088,N_21678,N_21125);
and U24089 (N_24089,N_20910,N_22280);
and U24090 (N_24090,N_22286,N_20903);
and U24091 (N_24091,N_20842,N_22398);
or U24092 (N_24092,N_20683,N_20658);
or U24093 (N_24093,N_20794,N_21338);
or U24094 (N_24094,N_21209,N_21538);
nor U24095 (N_24095,N_20563,N_21742);
nand U24096 (N_24096,N_20479,N_21250);
nor U24097 (N_24097,N_20981,N_22045);
or U24098 (N_24098,N_21218,N_20578);
and U24099 (N_24099,N_22399,N_21204);
nand U24100 (N_24100,N_22496,N_20775);
or U24101 (N_24101,N_20246,N_21459);
xor U24102 (N_24102,N_21533,N_20107);
nand U24103 (N_24103,N_22006,N_20846);
or U24104 (N_24104,N_20075,N_21845);
nor U24105 (N_24105,N_22407,N_21585);
and U24106 (N_24106,N_20844,N_20108);
and U24107 (N_24107,N_21313,N_21053);
xor U24108 (N_24108,N_22094,N_21164);
or U24109 (N_24109,N_21779,N_21418);
nand U24110 (N_24110,N_21468,N_20793);
or U24111 (N_24111,N_21345,N_21839);
or U24112 (N_24112,N_20314,N_21657);
nor U24113 (N_24113,N_21189,N_22167);
nand U24114 (N_24114,N_22359,N_21523);
xor U24115 (N_24115,N_21837,N_20108);
nand U24116 (N_24116,N_21429,N_20586);
and U24117 (N_24117,N_20631,N_22368);
nor U24118 (N_24118,N_21742,N_22426);
nand U24119 (N_24119,N_20004,N_20978);
nand U24120 (N_24120,N_20416,N_20572);
xor U24121 (N_24121,N_21477,N_21042);
xnor U24122 (N_24122,N_21089,N_20999);
nor U24123 (N_24123,N_21739,N_22460);
and U24124 (N_24124,N_21645,N_20089);
and U24125 (N_24125,N_22237,N_22128);
and U24126 (N_24126,N_21601,N_20332);
nor U24127 (N_24127,N_21475,N_21821);
nand U24128 (N_24128,N_22186,N_20380);
or U24129 (N_24129,N_22310,N_20397);
nand U24130 (N_24130,N_20642,N_21712);
or U24131 (N_24131,N_20970,N_22371);
and U24132 (N_24132,N_20489,N_20881);
and U24133 (N_24133,N_22395,N_21569);
nor U24134 (N_24134,N_21094,N_21883);
and U24135 (N_24135,N_22274,N_20433);
nor U24136 (N_24136,N_21834,N_21128);
xnor U24137 (N_24137,N_20343,N_20153);
or U24138 (N_24138,N_21789,N_21726);
nor U24139 (N_24139,N_21745,N_21634);
nand U24140 (N_24140,N_20352,N_20220);
nor U24141 (N_24141,N_20273,N_20601);
nand U24142 (N_24142,N_21663,N_20462);
nor U24143 (N_24143,N_21837,N_22206);
nand U24144 (N_24144,N_20182,N_21467);
and U24145 (N_24145,N_20563,N_20746);
nor U24146 (N_24146,N_21571,N_21644);
and U24147 (N_24147,N_22465,N_21714);
and U24148 (N_24148,N_20011,N_20309);
or U24149 (N_24149,N_20531,N_20957);
xnor U24150 (N_24150,N_22413,N_22104);
or U24151 (N_24151,N_22465,N_21125);
nor U24152 (N_24152,N_20846,N_20377);
or U24153 (N_24153,N_22467,N_21892);
nor U24154 (N_24154,N_22047,N_20033);
nand U24155 (N_24155,N_20368,N_21059);
and U24156 (N_24156,N_20483,N_20512);
nand U24157 (N_24157,N_21045,N_21148);
nand U24158 (N_24158,N_21768,N_21829);
and U24159 (N_24159,N_22369,N_22270);
nand U24160 (N_24160,N_21303,N_22193);
and U24161 (N_24161,N_22183,N_20923);
nor U24162 (N_24162,N_22406,N_20450);
nor U24163 (N_24163,N_20824,N_20130);
and U24164 (N_24164,N_20199,N_20405);
nor U24165 (N_24165,N_22140,N_22319);
nor U24166 (N_24166,N_20601,N_22201);
or U24167 (N_24167,N_20510,N_20278);
nor U24168 (N_24168,N_21649,N_21552);
nor U24169 (N_24169,N_22062,N_21937);
and U24170 (N_24170,N_20909,N_21413);
or U24171 (N_24171,N_21648,N_21664);
or U24172 (N_24172,N_20752,N_21540);
and U24173 (N_24173,N_21176,N_22113);
or U24174 (N_24174,N_21720,N_20662);
nand U24175 (N_24175,N_21212,N_22069);
xnor U24176 (N_24176,N_20921,N_21783);
or U24177 (N_24177,N_20749,N_21474);
nand U24178 (N_24178,N_20826,N_22442);
nor U24179 (N_24179,N_22346,N_20614);
and U24180 (N_24180,N_20402,N_21094);
and U24181 (N_24181,N_21075,N_20331);
and U24182 (N_24182,N_21048,N_20785);
nand U24183 (N_24183,N_21191,N_20190);
nand U24184 (N_24184,N_21715,N_20495);
or U24185 (N_24185,N_20173,N_20218);
nor U24186 (N_24186,N_21709,N_21118);
and U24187 (N_24187,N_20528,N_20716);
or U24188 (N_24188,N_20360,N_20323);
or U24189 (N_24189,N_20134,N_21861);
or U24190 (N_24190,N_21052,N_21176);
nand U24191 (N_24191,N_22428,N_20148);
and U24192 (N_24192,N_20678,N_21546);
or U24193 (N_24193,N_20449,N_21570);
or U24194 (N_24194,N_20555,N_20662);
nand U24195 (N_24195,N_20740,N_22171);
nand U24196 (N_24196,N_20615,N_20551);
xor U24197 (N_24197,N_20730,N_20912);
nand U24198 (N_24198,N_20895,N_20614);
and U24199 (N_24199,N_22070,N_20827);
xor U24200 (N_24200,N_20895,N_20494);
or U24201 (N_24201,N_21216,N_20437);
nor U24202 (N_24202,N_21738,N_20851);
and U24203 (N_24203,N_21679,N_21800);
or U24204 (N_24204,N_20642,N_20304);
nor U24205 (N_24205,N_21174,N_20228);
nor U24206 (N_24206,N_20827,N_21192);
nor U24207 (N_24207,N_21670,N_21397);
nor U24208 (N_24208,N_21315,N_21148);
nand U24209 (N_24209,N_22356,N_20978);
and U24210 (N_24210,N_22415,N_20530);
nor U24211 (N_24211,N_21531,N_22499);
nor U24212 (N_24212,N_21740,N_20971);
and U24213 (N_24213,N_20647,N_21137);
nand U24214 (N_24214,N_21962,N_21611);
or U24215 (N_24215,N_21811,N_20858);
nand U24216 (N_24216,N_20975,N_21311);
and U24217 (N_24217,N_22431,N_22384);
xor U24218 (N_24218,N_20885,N_20425);
or U24219 (N_24219,N_22461,N_20313);
and U24220 (N_24220,N_21065,N_21098);
and U24221 (N_24221,N_21322,N_20130);
xor U24222 (N_24222,N_22488,N_21671);
nor U24223 (N_24223,N_20571,N_21981);
nor U24224 (N_24224,N_20401,N_22269);
and U24225 (N_24225,N_21220,N_22398);
nor U24226 (N_24226,N_21185,N_20899);
and U24227 (N_24227,N_22359,N_20300);
and U24228 (N_24228,N_21404,N_22064);
xor U24229 (N_24229,N_20991,N_21356);
nand U24230 (N_24230,N_21298,N_21598);
nand U24231 (N_24231,N_22252,N_22445);
or U24232 (N_24232,N_20817,N_21259);
or U24233 (N_24233,N_20573,N_20170);
xnor U24234 (N_24234,N_21733,N_21735);
or U24235 (N_24235,N_20143,N_21110);
and U24236 (N_24236,N_21191,N_21287);
nor U24237 (N_24237,N_21450,N_21718);
or U24238 (N_24238,N_21987,N_21028);
nand U24239 (N_24239,N_21368,N_21046);
and U24240 (N_24240,N_21467,N_21032);
nor U24241 (N_24241,N_20816,N_21262);
and U24242 (N_24242,N_21292,N_22222);
or U24243 (N_24243,N_22122,N_20103);
and U24244 (N_24244,N_22304,N_22424);
and U24245 (N_24245,N_20802,N_21993);
or U24246 (N_24246,N_20935,N_20190);
nor U24247 (N_24247,N_20907,N_22416);
nor U24248 (N_24248,N_20383,N_21729);
and U24249 (N_24249,N_21907,N_20871);
or U24250 (N_24250,N_20007,N_20282);
nor U24251 (N_24251,N_20592,N_22003);
nor U24252 (N_24252,N_22435,N_22244);
or U24253 (N_24253,N_22041,N_20219);
or U24254 (N_24254,N_21756,N_20619);
and U24255 (N_24255,N_20561,N_20752);
nor U24256 (N_24256,N_20213,N_22189);
nand U24257 (N_24257,N_21307,N_20703);
or U24258 (N_24258,N_22409,N_20066);
nor U24259 (N_24259,N_21670,N_21238);
nand U24260 (N_24260,N_20427,N_22204);
and U24261 (N_24261,N_20772,N_20199);
nand U24262 (N_24262,N_20643,N_22310);
nand U24263 (N_24263,N_21769,N_21639);
or U24264 (N_24264,N_22065,N_20414);
nor U24265 (N_24265,N_22379,N_22243);
nand U24266 (N_24266,N_20368,N_20921);
nor U24267 (N_24267,N_21229,N_20754);
or U24268 (N_24268,N_20679,N_22194);
and U24269 (N_24269,N_22379,N_20826);
and U24270 (N_24270,N_20934,N_21285);
nand U24271 (N_24271,N_21786,N_21575);
or U24272 (N_24272,N_21235,N_21266);
nand U24273 (N_24273,N_20529,N_22088);
or U24274 (N_24274,N_20045,N_20709);
nand U24275 (N_24275,N_20702,N_21435);
xor U24276 (N_24276,N_21592,N_20801);
or U24277 (N_24277,N_21450,N_20935);
nor U24278 (N_24278,N_20288,N_20051);
nor U24279 (N_24279,N_21291,N_22481);
or U24280 (N_24280,N_21522,N_21390);
nand U24281 (N_24281,N_21996,N_20951);
nand U24282 (N_24282,N_20011,N_21855);
nand U24283 (N_24283,N_20519,N_20052);
and U24284 (N_24284,N_20665,N_21769);
and U24285 (N_24285,N_21150,N_20899);
or U24286 (N_24286,N_20783,N_22149);
and U24287 (N_24287,N_20500,N_21208);
nand U24288 (N_24288,N_21500,N_20530);
and U24289 (N_24289,N_22124,N_21670);
or U24290 (N_24290,N_20323,N_21986);
and U24291 (N_24291,N_21445,N_21041);
nor U24292 (N_24292,N_20563,N_20728);
or U24293 (N_24293,N_21321,N_22442);
nand U24294 (N_24294,N_20289,N_20326);
xnor U24295 (N_24295,N_20879,N_22016);
nand U24296 (N_24296,N_21050,N_22344);
or U24297 (N_24297,N_20805,N_21454);
nand U24298 (N_24298,N_21179,N_20504);
xor U24299 (N_24299,N_21631,N_22482);
and U24300 (N_24300,N_20830,N_20597);
nor U24301 (N_24301,N_20219,N_22439);
xnor U24302 (N_24302,N_21957,N_21548);
or U24303 (N_24303,N_21617,N_20239);
or U24304 (N_24304,N_20160,N_21389);
xnor U24305 (N_24305,N_22161,N_21224);
nand U24306 (N_24306,N_20272,N_20013);
and U24307 (N_24307,N_21480,N_21618);
nor U24308 (N_24308,N_21260,N_21240);
and U24309 (N_24309,N_20441,N_20275);
nor U24310 (N_24310,N_20483,N_21441);
xnor U24311 (N_24311,N_20456,N_20373);
nand U24312 (N_24312,N_20978,N_20233);
and U24313 (N_24313,N_20363,N_20349);
xnor U24314 (N_24314,N_22364,N_21775);
or U24315 (N_24315,N_21652,N_20052);
nand U24316 (N_24316,N_21173,N_20315);
nor U24317 (N_24317,N_20081,N_20682);
nor U24318 (N_24318,N_22252,N_22139);
nand U24319 (N_24319,N_21887,N_21916);
xnor U24320 (N_24320,N_21660,N_20131);
xor U24321 (N_24321,N_20181,N_21781);
nand U24322 (N_24322,N_20172,N_20103);
and U24323 (N_24323,N_21427,N_20288);
or U24324 (N_24324,N_21453,N_22058);
nor U24325 (N_24325,N_22329,N_21966);
nand U24326 (N_24326,N_20983,N_20019);
or U24327 (N_24327,N_22411,N_20814);
nand U24328 (N_24328,N_21541,N_21730);
nand U24329 (N_24329,N_21705,N_20915);
nor U24330 (N_24330,N_21148,N_20977);
and U24331 (N_24331,N_20718,N_21597);
and U24332 (N_24332,N_22031,N_21065);
nand U24333 (N_24333,N_21287,N_20080);
and U24334 (N_24334,N_20712,N_22150);
and U24335 (N_24335,N_21958,N_20868);
xnor U24336 (N_24336,N_20603,N_21301);
or U24337 (N_24337,N_20636,N_22255);
nand U24338 (N_24338,N_20432,N_21185);
and U24339 (N_24339,N_20771,N_20905);
or U24340 (N_24340,N_21177,N_20130);
nand U24341 (N_24341,N_20290,N_22321);
nor U24342 (N_24342,N_21415,N_21744);
and U24343 (N_24343,N_21938,N_20486);
and U24344 (N_24344,N_22040,N_22366);
nand U24345 (N_24345,N_20922,N_22444);
or U24346 (N_24346,N_20597,N_22273);
xnor U24347 (N_24347,N_21843,N_20386);
and U24348 (N_24348,N_22431,N_21383);
nand U24349 (N_24349,N_22025,N_20064);
or U24350 (N_24350,N_21321,N_22388);
or U24351 (N_24351,N_21563,N_21750);
and U24352 (N_24352,N_22425,N_20748);
nand U24353 (N_24353,N_20903,N_21430);
nand U24354 (N_24354,N_20174,N_21514);
and U24355 (N_24355,N_20008,N_21291);
nor U24356 (N_24356,N_20131,N_22181);
nand U24357 (N_24357,N_20684,N_22449);
nand U24358 (N_24358,N_20935,N_22348);
nand U24359 (N_24359,N_20861,N_22488);
nand U24360 (N_24360,N_20284,N_20152);
and U24361 (N_24361,N_20218,N_21586);
or U24362 (N_24362,N_21913,N_20175);
or U24363 (N_24363,N_21674,N_21183);
and U24364 (N_24364,N_20768,N_22131);
nand U24365 (N_24365,N_21044,N_21135);
xnor U24366 (N_24366,N_20320,N_20668);
and U24367 (N_24367,N_20720,N_20162);
and U24368 (N_24368,N_22170,N_20079);
nand U24369 (N_24369,N_22390,N_20600);
and U24370 (N_24370,N_21026,N_21541);
or U24371 (N_24371,N_22377,N_22310);
and U24372 (N_24372,N_22009,N_20991);
and U24373 (N_24373,N_20490,N_21362);
or U24374 (N_24374,N_20818,N_21647);
and U24375 (N_24375,N_21992,N_20048);
or U24376 (N_24376,N_20836,N_21029);
nor U24377 (N_24377,N_21363,N_20710);
xor U24378 (N_24378,N_22230,N_20478);
nand U24379 (N_24379,N_20469,N_22364);
or U24380 (N_24380,N_20208,N_20969);
nand U24381 (N_24381,N_20689,N_21024);
and U24382 (N_24382,N_20350,N_20986);
nor U24383 (N_24383,N_21414,N_21058);
and U24384 (N_24384,N_21263,N_20861);
nor U24385 (N_24385,N_20917,N_21796);
nor U24386 (N_24386,N_21524,N_21945);
and U24387 (N_24387,N_20889,N_22121);
nor U24388 (N_24388,N_20870,N_20564);
nor U24389 (N_24389,N_20885,N_20546);
and U24390 (N_24390,N_21097,N_21881);
nand U24391 (N_24391,N_20962,N_21825);
nor U24392 (N_24392,N_21330,N_21423);
or U24393 (N_24393,N_20399,N_22216);
and U24394 (N_24394,N_20859,N_21141);
xor U24395 (N_24395,N_22065,N_22231);
nand U24396 (N_24396,N_21529,N_21457);
nand U24397 (N_24397,N_21596,N_20155);
xnor U24398 (N_24398,N_21014,N_20840);
or U24399 (N_24399,N_21249,N_20992);
nor U24400 (N_24400,N_21606,N_20636);
and U24401 (N_24401,N_20398,N_21880);
and U24402 (N_24402,N_20673,N_20096);
nand U24403 (N_24403,N_22178,N_21780);
or U24404 (N_24404,N_20029,N_21843);
nand U24405 (N_24405,N_22058,N_20981);
nor U24406 (N_24406,N_22440,N_21661);
nor U24407 (N_24407,N_21716,N_21044);
or U24408 (N_24408,N_21683,N_21081);
nor U24409 (N_24409,N_21921,N_21108);
and U24410 (N_24410,N_21139,N_20299);
or U24411 (N_24411,N_21283,N_22205);
xor U24412 (N_24412,N_21341,N_20774);
xnor U24413 (N_24413,N_20031,N_21772);
nand U24414 (N_24414,N_22350,N_21896);
or U24415 (N_24415,N_20421,N_20314);
and U24416 (N_24416,N_22153,N_21158);
nor U24417 (N_24417,N_21036,N_20298);
or U24418 (N_24418,N_21216,N_21662);
xnor U24419 (N_24419,N_20640,N_22171);
nor U24420 (N_24420,N_20258,N_21626);
xor U24421 (N_24421,N_22469,N_21088);
nor U24422 (N_24422,N_21233,N_22315);
xnor U24423 (N_24423,N_21611,N_20149);
or U24424 (N_24424,N_21046,N_20537);
and U24425 (N_24425,N_21253,N_22014);
and U24426 (N_24426,N_21263,N_21264);
or U24427 (N_24427,N_21082,N_21828);
xnor U24428 (N_24428,N_20327,N_20442);
nor U24429 (N_24429,N_20078,N_21942);
xnor U24430 (N_24430,N_20086,N_21967);
xor U24431 (N_24431,N_21341,N_20585);
nor U24432 (N_24432,N_21156,N_21370);
xor U24433 (N_24433,N_21627,N_20018);
nand U24434 (N_24434,N_20657,N_22149);
nor U24435 (N_24435,N_21982,N_22076);
or U24436 (N_24436,N_21754,N_20103);
and U24437 (N_24437,N_21128,N_20819);
xor U24438 (N_24438,N_22346,N_21515);
nor U24439 (N_24439,N_21969,N_21710);
and U24440 (N_24440,N_20763,N_20960);
nor U24441 (N_24441,N_22311,N_21625);
or U24442 (N_24442,N_22140,N_20756);
nor U24443 (N_24443,N_20693,N_20444);
nand U24444 (N_24444,N_20978,N_21058);
nand U24445 (N_24445,N_20936,N_20599);
or U24446 (N_24446,N_21905,N_20603);
or U24447 (N_24447,N_20855,N_21716);
nand U24448 (N_24448,N_21020,N_22450);
nor U24449 (N_24449,N_20349,N_21936);
nand U24450 (N_24450,N_22362,N_20768);
nand U24451 (N_24451,N_20947,N_21111);
or U24452 (N_24452,N_22470,N_21302);
nor U24453 (N_24453,N_21994,N_20937);
xnor U24454 (N_24454,N_20242,N_21050);
or U24455 (N_24455,N_22024,N_21957);
and U24456 (N_24456,N_20738,N_21259);
xnor U24457 (N_24457,N_21876,N_20192);
nor U24458 (N_24458,N_21015,N_20546);
and U24459 (N_24459,N_20535,N_21621);
nor U24460 (N_24460,N_21319,N_22194);
or U24461 (N_24461,N_22350,N_21253);
nor U24462 (N_24462,N_21329,N_20012);
or U24463 (N_24463,N_20266,N_20395);
and U24464 (N_24464,N_20933,N_21928);
or U24465 (N_24465,N_21798,N_22440);
or U24466 (N_24466,N_22149,N_20418);
and U24467 (N_24467,N_22181,N_22324);
nand U24468 (N_24468,N_22022,N_20013);
and U24469 (N_24469,N_20763,N_21290);
or U24470 (N_24470,N_21207,N_21548);
and U24471 (N_24471,N_20441,N_22406);
nand U24472 (N_24472,N_22053,N_22443);
or U24473 (N_24473,N_21112,N_22406);
and U24474 (N_24474,N_20110,N_21894);
nand U24475 (N_24475,N_20561,N_22143);
or U24476 (N_24476,N_22274,N_21724);
nand U24477 (N_24477,N_21062,N_20829);
and U24478 (N_24478,N_21903,N_21425);
or U24479 (N_24479,N_21379,N_21805);
and U24480 (N_24480,N_20310,N_20705);
and U24481 (N_24481,N_20557,N_20017);
or U24482 (N_24482,N_21712,N_20425);
or U24483 (N_24483,N_22288,N_20810);
or U24484 (N_24484,N_21418,N_21359);
nor U24485 (N_24485,N_21656,N_20689);
and U24486 (N_24486,N_22329,N_21771);
or U24487 (N_24487,N_22285,N_20618);
nand U24488 (N_24488,N_21276,N_21507);
nor U24489 (N_24489,N_21725,N_20337);
xnor U24490 (N_24490,N_20595,N_21018);
or U24491 (N_24491,N_20586,N_20932);
or U24492 (N_24492,N_21938,N_20728);
nand U24493 (N_24493,N_21394,N_22004);
nand U24494 (N_24494,N_20726,N_20081);
or U24495 (N_24495,N_20657,N_20505);
nand U24496 (N_24496,N_20930,N_20447);
and U24497 (N_24497,N_20245,N_21305);
or U24498 (N_24498,N_20539,N_20757);
and U24499 (N_24499,N_21483,N_21280);
nand U24500 (N_24500,N_20319,N_20932);
and U24501 (N_24501,N_21550,N_22014);
nor U24502 (N_24502,N_21213,N_20286);
nor U24503 (N_24503,N_22371,N_22487);
and U24504 (N_24504,N_20038,N_20114);
nor U24505 (N_24505,N_21243,N_21881);
nor U24506 (N_24506,N_21463,N_20846);
and U24507 (N_24507,N_20547,N_21469);
or U24508 (N_24508,N_20020,N_20460);
nor U24509 (N_24509,N_20920,N_21101);
nand U24510 (N_24510,N_20359,N_22475);
nand U24511 (N_24511,N_20144,N_22296);
or U24512 (N_24512,N_21763,N_21803);
xnor U24513 (N_24513,N_20072,N_21334);
and U24514 (N_24514,N_20545,N_20651);
or U24515 (N_24515,N_21100,N_22056);
nor U24516 (N_24516,N_21569,N_20567);
nor U24517 (N_24517,N_22055,N_20209);
nand U24518 (N_24518,N_20398,N_20436);
or U24519 (N_24519,N_21207,N_20927);
xnor U24520 (N_24520,N_20419,N_21244);
nand U24521 (N_24521,N_22166,N_20972);
nand U24522 (N_24522,N_21813,N_20681);
or U24523 (N_24523,N_20448,N_20254);
nand U24524 (N_24524,N_21429,N_21117);
nor U24525 (N_24525,N_21543,N_21027);
nor U24526 (N_24526,N_20882,N_22257);
nand U24527 (N_24527,N_21116,N_20953);
xnor U24528 (N_24528,N_20350,N_20891);
nand U24529 (N_24529,N_20574,N_21241);
and U24530 (N_24530,N_22289,N_21476);
or U24531 (N_24531,N_21456,N_20085);
nand U24532 (N_24532,N_22059,N_20920);
nand U24533 (N_24533,N_22025,N_21246);
or U24534 (N_24534,N_20180,N_21679);
nand U24535 (N_24535,N_20155,N_20074);
nor U24536 (N_24536,N_22376,N_22010);
or U24537 (N_24537,N_21894,N_20817);
xor U24538 (N_24538,N_22063,N_22450);
nand U24539 (N_24539,N_20232,N_20872);
nand U24540 (N_24540,N_20088,N_21005);
or U24541 (N_24541,N_20999,N_20557);
or U24542 (N_24542,N_20594,N_21737);
nor U24543 (N_24543,N_20593,N_21011);
nand U24544 (N_24544,N_21996,N_20025);
and U24545 (N_24545,N_22312,N_20168);
nand U24546 (N_24546,N_22133,N_20686);
nor U24547 (N_24547,N_22253,N_20702);
nor U24548 (N_24548,N_20454,N_20926);
and U24549 (N_24549,N_21529,N_21824);
and U24550 (N_24550,N_22064,N_21426);
nand U24551 (N_24551,N_22208,N_20328);
nor U24552 (N_24552,N_20866,N_20768);
nor U24553 (N_24553,N_20807,N_21976);
and U24554 (N_24554,N_22388,N_21186);
nor U24555 (N_24555,N_21018,N_22179);
nand U24556 (N_24556,N_22036,N_20772);
nand U24557 (N_24557,N_21875,N_22148);
and U24558 (N_24558,N_20219,N_22226);
or U24559 (N_24559,N_20925,N_20535);
nor U24560 (N_24560,N_20751,N_20649);
xor U24561 (N_24561,N_21560,N_20162);
nand U24562 (N_24562,N_22032,N_21361);
and U24563 (N_24563,N_21760,N_21186);
or U24564 (N_24564,N_20244,N_21903);
or U24565 (N_24565,N_20424,N_21757);
or U24566 (N_24566,N_20053,N_20195);
or U24567 (N_24567,N_21759,N_21301);
nand U24568 (N_24568,N_21449,N_21898);
xnor U24569 (N_24569,N_20571,N_21519);
xor U24570 (N_24570,N_21367,N_21013);
or U24571 (N_24571,N_21459,N_20103);
and U24572 (N_24572,N_21438,N_20561);
and U24573 (N_24573,N_21136,N_22203);
nand U24574 (N_24574,N_20157,N_21740);
or U24575 (N_24575,N_21819,N_22051);
and U24576 (N_24576,N_21588,N_21757);
or U24577 (N_24577,N_21893,N_22115);
nor U24578 (N_24578,N_20638,N_20510);
or U24579 (N_24579,N_20782,N_20375);
or U24580 (N_24580,N_22137,N_20246);
and U24581 (N_24581,N_20727,N_20358);
xor U24582 (N_24582,N_20205,N_21283);
or U24583 (N_24583,N_22388,N_20430);
nor U24584 (N_24584,N_22238,N_21440);
nor U24585 (N_24585,N_21804,N_22320);
or U24586 (N_24586,N_20872,N_21190);
nor U24587 (N_24587,N_20548,N_21641);
nand U24588 (N_24588,N_22294,N_21408);
nor U24589 (N_24589,N_22136,N_21764);
nand U24590 (N_24590,N_22280,N_21655);
or U24591 (N_24591,N_21861,N_20217);
nor U24592 (N_24592,N_21888,N_21142);
nand U24593 (N_24593,N_21388,N_21612);
and U24594 (N_24594,N_20837,N_20753);
or U24595 (N_24595,N_22186,N_22283);
or U24596 (N_24596,N_22448,N_21652);
nor U24597 (N_24597,N_21048,N_21976);
nand U24598 (N_24598,N_20836,N_20366);
or U24599 (N_24599,N_20889,N_22309);
or U24600 (N_24600,N_20137,N_21227);
and U24601 (N_24601,N_20299,N_21882);
xnor U24602 (N_24602,N_20754,N_20054);
and U24603 (N_24603,N_22457,N_20101);
nor U24604 (N_24604,N_21108,N_21442);
or U24605 (N_24605,N_22445,N_21463);
xnor U24606 (N_24606,N_20150,N_20103);
or U24607 (N_24607,N_21324,N_21840);
or U24608 (N_24608,N_20871,N_20332);
nor U24609 (N_24609,N_21975,N_21960);
nand U24610 (N_24610,N_21276,N_21322);
or U24611 (N_24611,N_21477,N_21807);
or U24612 (N_24612,N_20976,N_20126);
nor U24613 (N_24613,N_21813,N_22087);
and U24614 (N_24614,N_21935,N_22379);
and U24615 (N_24615,N_20092,N_20863);
or U24616 (N_24616,N_22425,N_21117);
nor U24617 (N_24617,N_20236,N_20649);
or U24618 (N_24618,N_22451,N_21854);
nor U24619 (N_24619,N_20070,N_21232);
nor U24620 (N_24620,N_20232,N_22211);
or U24621 (N_24621,N_22411,N_20658);
nor U24622 (N_24622,N_21880,N_21421);
or U24623 (N_24623,N_21936,N_22421);
nand U24624 (N_24624,N_20624,N_20332);
nand U24625 (N_24625,N_22245,N_21479);
and U24626 (N_24626,N_21028,N_20298);
nor U24627 (N_24627,N_22005,N_22057);
nor U24628 (N_24628,N_20084,N_21370);
or U24629 (N_24629,N_20355,N_22359);
and U24630 (N_24630,N_22137,N_21162);
or U24631 (N_24631,N_21978,N_20913);
and U24632 (N_24632,N_20260,N_20202);
nor U24633 (N_24633,N_21692,N_20908);
or U24634 (N_24634,N_20896,N_21867);
and U24635 (N_24635,N_20383,N_21637);
nand U24636 (N_24636,N_20408,N_21790);
or U24637 (N_24637,N_22303,N_22149);
nor U24638 (N_24638,N_20089,N_21502);
and U24639 (N_24639,N_21238,N_22428);
nor U24640 (N_24640,N_21124,N_21492);
nand U24641 (N_24641,N_22427,N_22173);
or U24642 (N_24642,N_22432,N_20896);
or U24643 (N_24643,N_22209,N_21988);
nand U24644 (N_24644,N_20019,N_21397);
xnor U24645 (N_24645,N_21074,N_22415);
nand U24646 (N_24646,N_20768,N_21419);
nor U24647 (N_24647,N_20439,N_21802);
or U24648 (N_24648,N_22439,N_20491);
or U24649 (N_24649,N_21461,N_20862);
xnor U24650 (N_24650,N_21459,N_20087);
nor U24651 (N_24651,N_22232,N_21782);
or U24652 (N_24652,N_20081,N_22087);
nor U24653 (N_24653,N_21190,N_22307);
and U24654 (N_24654,N_21126,N_21945);
xnor U24655 (N_24655,N_21566,N_22318);
nor U24656 (N_24656,N_21237,N_20318);
and U24657 (N_24657,N_22088,N_20317);
nand U24658 (N_24658,N_20140,N_22361);
xnor U24659 (N_24659,N_20914,N_20808);
nor U24660 (N_24660,N_21308,N_20123);
nor U24661 (N_24661,N_21405,N_20275);
nand U24662 (N_24662,N_22109,N_20080);
and U24663 (N_24663,N_21245,N_21591);
or U24664 (N_24664,N_20047,N_22154);
nor U24665 (N_24665,N_21359,N_21341);
nand U24666 (N_24666,N_20711,N_21534);
nand U24667 (N_24667,N_22229,N_21129);
nand U24668 (N_24668,N_20064,N_20986);
nand U24669 (N_24669,N_21926,N_22156);
or U24670 (N_24670,N_20430,N_22064);
or U24671 (N_24671,N_20461,N_21238);
nor U24672 (N_24672,N_22365,N_22499);
nor U24673 (N_24673,N_20894,N_21434);
or U24674 (N_24674,N_22218,N_22424);
and U24675 (N_24675,N_22167,N_20994);
nand U24676 (N_24676,N_20101,N_21631);
and U24677 (N_24677,N_21092,N_20956);
or U24678 (N_24678,N_21952,N_20289);
or U24679 (N_24679,N_21987,N_22209);
and U24680 (N_24680,N_20987,N_21949);
and U24681 (N_24681,N_20705,N_20982);
nand U24682 (N_24682,N_20723,N_20064);
and U24683 (N_24683,N_20478,N_22048);
nand U24684 (N_24684,N_22262,N_20217);
and U24685 (N_24685,N_21351,N_20831);
nor U24686 (N_24686,N_20435,N_22456);
nand U24687 (N_24687,N_21778,N_22424);
nor U24688 (N_24688,N_22380,N_20455);
or U24689 (N_24689,N_22215,N_20676);
nand U24690 (N_24690,N_20431,N_21994);
nor U24691 (N_24691,N_22187,N_20764);
nand U24692 (N_24692,N_20718,N_21497);
nor U24693 (N_24693,N_21375,N_20092);
or U24694 (N_24694,N_21114,N_22409);
or U24695 (N_24695,N_20630,N_20171);
nor U24696 (N_24696,N_20907,N_21788);
nand U24697 (N_24697,N_21476,N_20586);
nand U24698 (N_24698,N_21387,N_21696);
nor U24699 (N_24699,N_21749,N_21493);
and U24700 (N_24700,N_20408,N_20042);
nor U24701 (N_24701,N_21019,N_21398);
or U24702 (N_24702,N_20856,N_22181);
and U24703 (N_24703,N_20668,N_21570);
and U24704 (N_24704,N_21610,N_21723);
or U24705 (N_24705,N_21377,N_20279);
nor U24706 (N_24706,N_20087,N_21558);
nand U24707 (N_24707,N_21511,N_21887);
nor U24708 (N_24708,N_21579,N_21583);
nand U24709 (N_24709,N_20341,N_21533);
and U24710 (N_24710,N_22103,N_20631);
or U24711 (N_24711,N_21148,N_21525);
or U24712 (N_24712,N_21503,N_20859);
and U24713 (N_24713,N_20312,N_20374);
and U24714 (N_24714,N_22196,N_22497);
nor U24715 (N_24715,N_21033,N_20874);
and U24716 (N_24716,N_20961,N_21984);
nor U24717 (N_24717,N_22230,N_21667);
xnor U24718 (N_24718,N_20433,N_20099);
and U24719 (N_24719,N_21733,N_20221);
or U24720 (N_24720,N_22204,N_22302);
nor U24721 (N_24721,N_22239,N_22110);
and U24722 (N_24722,N_21869,N_21349);
nand U24723 (N_24723,N_20451,N_20581);
and U24724 (N_24724,N_20510,N_22251);
or U24725 (N_24725,N_22288,N_20275);
and U24726 (N_24726,N_21600,N_20379);
and U24727 (N_24727,N_22301,N_21703);
or U24728 (N_24728,N_20332,N_21045);
and U24729 (N_24729,N_21859,N_21895);
or U24730 (N_24730,N_20939,N_21105);
nor U24731 (N_24731,N_21565,N_22049);
nor U24732 (N_24732,N_21382,N_20324);
and U24733 (N_24733,N_20745,N_20908);
xor U24734 (N_24734,N_20976,N_21875);
or U24735 (N_24735,N_20904,N_20401);
xor U24736 (N_24736,N_21036,N_22412);
nand U24737 (N_24737,N_20607,N_22307);
or U24738 (N_24738,N_20734,N_21236);
nand U24739 (N_24739,N_22056,N_20187);
nand U24740 (N_24740,N_20216,N_21992);
and U24741 (N_24741,N_20186,N_21216);
nor U24742 (N_24742,N_21734,N_21187);
or U24743 (N_24743,N_20788,N_22372);
nand U24744 (N_24744,N_22291,N_22350);
or U24745 (N_24745,N_22265,N_22242);
or U24746 (N_24746,N_20977,N_20693);
nor U24747 (N_24747,N_20246,N_21252);
and U24748 (N_24748,N_22153,N_21608);
or U24749 (N_24749,N_21162,N_21872);
nor U24750 (N_24750,N_20205,N_21655);
nor U24751 (N_24751,N_22263,N_20803);
and U24752 (N_24752,N_22049,N_21116);
xnor U24753 (N_24753,N_22083,N_20849);
nand U24754 (N_24754,N_20978,N_22138);
nand U24755 (N_24755,N_20167,N_20216);
or U24756 (N_24756,N_20569,N_22162);
nand U24757 (N_24757,N_20019,N_21570);
or U24758 (N_24758,N_21075,N_21313);
and U24759 (N_24759,N_22351,N_20581);
nand U24760 (N_24760,N_20895,N_22230);
nor U24761 (N_24761,N_21992,N_20409);
nand U24762 (N_24762,N_21843,N_21131);
nand U24763 (N_24763,N_21713,N_21439);
nand U24764 (N_24764,N_22314,N_22038);
nand U24765 (N_24765,N_20068,N_21917);
or U24766 (N_24766,N_22235,N_21223);
xor U24767 (N_24767,N_20338,N_22192);
or U24768 (N_24768,N_21367,N_21280);
or U24769 (N_24769,N_20355,N_21620);
xor U24770 (N_24770,N_21685,N_21397);
nand U24771 (N_24771,N_20935,N_20081);
or U24772 (N_24772,N_21403,N_22438);
nor U24773 (N_24773,N_20596,N_20302);
xnor U24774 (N_24774,N_20681,N_20828);
or U24775 (N_24775,N_20305,N_22020);
nor U24776 (N_24776,N_20083,N_20282);
nand U24777 (N_24777,N_21582,N_22035);
nor U24778 (N_24778,N_20171,N_22094);
or U24779 (N_24779,N_20887,N_22115);
or U24780 (N_24780,N_22295,N_20040);
nand U24781 (N_24781,N_20879,N_21727);
nand U24782 (N_24782,N_21048,N_21440);
nand U24783 (N_24783,N_21656,N_20108);
nor U24784 (N_24784,N_20234,N_20940);
nor U24785 (N_24785,N_21191,N_20799);
nor U24786 (N_24786,N_21172,N_20058);
and U24787 (N_24787,N_22023,N_20453);
nor U24788 (N_24788,N_22324,N_21443);
and U24789 (N_24789,N_21174,N_20106);
nand U24790 (N_24790,N_22170,N_20602);
nor U24791 (N_24791,N_20182,N_22152);
nor U24792 (N_24792,N_20906,N_20599);
nor U24793 (N_24793,N_20654,N_21233);
or U24794 (N_24794,N_21390,N_22243);
xor U24795 (N_24795,N_20993,N_20141);
or U24796 (N_24796,N_20483,N_20952);
nor U24797 (N_24797,N_21471,N_21977);
nand U24798 (N_24798,N_20459,N_20380);
and U24799 (N_24799,N_22290,N_21814);
and U24800 (N_24800,N_21847,N_20211);
nand U24801 (N_24801,N_20515,N_21669);
and U24802 (N_24802,N_20760,N_22348);
nor U24803 (N_24803,N_20045,N_21022);
nand U24804 (N_24804,N_21027,N_21130);
or U24805 (N_24805,N_20182,N_20557);
nor U24806 (N_24806,N_20885,N_21186);
nor U24807 (N_24807,N_20518,N_20448);
or U24808 (N_24808,N_20497,N_21556);
nor U24809 (N_24809,N_21832,N_20782);
nand U24810 (N_24810,N_21802,N_20317);
nand U24811 (N_24811,N_22085,N_21508);
nand U24812 (N_24812,N_21075,N_21557);
or U24813 (N_24813,N_20244,N_21013);
xnor U24814 (N_24814,N_21499,N_21000);
or U24815 (N_24815,N_21519,N_20631);
and U24816 (N_24816,N_22259,N_20522);
or U24817 (N_24817,N_21949,N_21278);
or U24818 (N_24818,N_21283,N_21611);
or U24819 (N_24819,N_20102,N_20504);
or U24820 (N_24820,N_20644,N_22423);
nand U24821 (N_24821,N_21179,N_21118);
or U24822 (N_24822,N_20772,N_20776);
nor U24823 (N_24823,N_21845,N_21878);
nand U24824 (N_24824,N_20284,N_20155);
nor U24825 (N_24825,N_21318,N_20452);
or U24826 (N_24826,N_20170,N_21278);
nor U24827 (N_24827,N_20728,N_22339);
nor U24828 (N_24828,N_20643,N_20618);
nor U24829 (N_24829,N_22294,N_21336);
or U24830 (N_24830,N_21847,N_22478);
nor U24831 (N_24831,N_22187,N_20004);
nand U24832 (N_24832,N_20629,N_20546);
and U24833 (N_24833,N_22165,N_21959);
xor U24834 (N_24834,N_21727,N_20825);
or U24835 (N_24835,N_21116,N_20312);
nor U24836 (N_24836,N_20339,N_20552);
xor U24837 (N_24837,N_21859,N_21925);
nor U24838 (N_24838,N_21884,N_21713);
or U24839 (N_24839,N_21322,N_21346);
nand U24840 (N_24840,N_20120,N_20709);
or U24841 (N_24841,N_21727,N_22200);
nor U24842 (N_24842,N_20162,N_22129);
or U24843 (N_24843,N_20666,N_20552);
xnor U24844 (N_24844,N_20463,N_21573);
nand U24845 (N_24845,N_20100,N_21528);
or U24846 (N_24846,N_20906,N_21558);
or U24847 (N_24847,N_20883,N_21055);
or U24848 (N_24848,N_22221,N_21268);
nor U24849 (N_24849,N_20811,N_20781);
xor U24850 (N_24850,N_22352,N_22227);
nor U24851 (N_24851,N_21654,N_22137);
xor U24852 (N_24852,N_21546,N_22129);
nor U24853 (N_24853,N_22198,N_20123);
and U24854 (N_24854,N_21331,N_22229);
and U24855 (N_24855,N_21358,N_20142);
xnor U24856 (N_24856,N_20619,N_22335);
and U24857 (N_24857,N_21746,N_21420);
nand U24858 (N_24858,N_20974,N_22172);
xnor U24859 (N_24859,N_22389,N_21735);
or U24860 (N_24860,N_20601,N_20749);
and U24861 (N_24861,N_20437,N_20408);
nor U24862 (N_24862,N_20338,N_20063);
nand U24863 (N_24863,N_22287,N_22136);
nand U24864 (N_24864,N_21595,N_21053);
or U24865 (N_24865,N_20486,N_22421);
nor U24866 (N_24866,N_20900,N_20340);
and U24867 (N_24867,N_22345,N_21065);
and U24868 (N_24868,N_21901,N_20142);
or U24869 (N_24869,N_22293,N_21088);
and U24870 (N_24870,N_20300,N_22100);
or U24871 (N_24871,N_20723,N_22291);
and U24872 (N_24872,N_22090,N_21994);
or U24873 (N_24873,N_20645,N_20372);
nand U24874 (N_24874,N_22468,N_20887);
nand U24875 (N_24875,N_22249,N_22376);
and U24876 (N_24876,N_22126,N_20981);
or U24877 (N_24877,N_20091,N_22386);
nand U24878 (N_24878,N_21620,N_20329);
nor U24879 (N_24879,N_22237,N_20879);
nand U24880 (N_24880,N_21409,N_20803);
nand U24881 (N_24881,N_21581,N_20600);
nand U24882 (N_24882,N_20546,N_20021);
or U24883 (N_24883,N_22456,N_22180);
and U24884 (N_24884,N_22473,N_20367);
or U24885 (N_24885,N_21964,N_21590);
nor U24886 (N_24886,N_20774,N_21694);
or U24887 (N_24887,N_21202,N_21091);
and U24888 (N_24888,N_21458,N_21857);
and U24889 (N_24889,N_20380,N_21219);
nor U24890 (N_24890,N_22189,N_20236);
nand U24891 (N_24891,N_20740,N_21760);
and U24892 (N_24892,N_21683,N_20411);
or U24893 (N_24893,N_20087,N_21736);
or U24894 (N_24894,N_20400,N_22294);
nand U24895 (N_24895,N_20023,N_22023);
or U24896 (N_24896,N_21919,N_20256);
and U24897 (N_24897,N_21200,N_20859);
or U24898 (N_24898,N_20319,N_20601);
or U24899 (N_24899,N_20064,N_20975);
and U24900 (N_24900,N_20910,N_21219);
xor U24901 (N_24901,N_20345,N_20217);
and U24902 (N_24902,N_21976,N_21158);
or U24903 (N_24903,N_21162,N_21897);
or U24904 (N_24904,N_21748,N_21024);
or U24905 (N_24905,N_20924,N_22040);
nand U24906 (N_24906,N_21256,N_22133);
nand U24907 (N_24907,N_22092,N_21948);
or U24908 (N_24908,N_22073,N_22349);
nor U24909 (N_24909,N_21454,N_21662);
and U24910 (N_24910,N_20835,N_20510);
nand U24911 (N_24911,N_20325,N_21103);
and U24912 (N_24912,N_20095,N_21284);
nand U24913 (N_24913,N_20744,N_20433);
or U24914 (N_24914,N_20768,N_22008);
nand U24915 (N_24915,N_22368,N_21623);
nor U24916 (N_24916,N_21303,N_21892);
nand U24917 (N_24917,N_21762,N_22195);
nor U24918 (N_24918,N_22366,N_22023);
nand U24919 (N_24919,N_20094,N_22084);
or U24920 (N_24920,N_20257,N_20320);
and U24921 (N_24921,N_20286,N_20791);
nand U24922 (N_24922,N_22129,N_20397);
or U24923 (N_24923,N_21661,N_20399);
nor U24924 (N_24924,N_22092,N_20783);
nor U24925 (N_24925,N_21675,N_22392);
and U24926 (N_24926,N_20149,N_21320);
and U24927 (N_24927,N_21884,N_21685);
xnor U24928 (N_24928,N_21239,N_20259);
and U24929 (N_24929,N_20679,N_20660);
or U24930 (N_24930,N_20757,N_22321);
nand U24931 (N_24931,N_21381,N_21739);
or U24932 (N_24932,N_22075,N_21978);
nand U24933 (N_24933,N_21645,N_22335);
and U24934 (N_24934,N_20037,N_22152);
nor U24935 (N_24935,N_21991,N_21211);
xor U24936 (N_24936,N_21752,N_20873);
nor U24937 (N_24937,N_21083,N_21058);
and U24938 (N_24938,N_20227,N_20590);
nand U24939 (N_24939,N_22109,N_22180);
nand U24940 (N_24940,N_20682,N_22311);
or U24941 (N_24941,N_21016,N_21026);
and U24942 (N_24942,N_20893,N_21312);
or U24943 (N_24943,N_20514,N_21896);
and U24944 (N_24944,N_21687,N_21186);
nand U24945 (N_24945,N_21633,N_20604);
and U24946 (N_24946,N_20146,N_22111);
or U24947 (N_24947,N_21110,N_21184);
nand U24948 (N_24948,N_22322,N_22112);
and U24949 (N_24949,N_20495,N_20426);
nand U24950 (N_24950,N_21261,N_20651);
or U24951 (N_24951,N_20336,N_20109);
nor U24952 (N_24952,N_20077,N_21886);
nor U24953 (N_24953,N_20135,N_21701);
and U24954 (N_24954,N_21080,N_21665);
or U24955 (N_24955,N_21014,N_20758);
and U24956 (N_24956,N_20516,N_22252);
nand U24957 (N_24957,N_21610,N_21642);
nand U24958 (N_24958,N_20596,N_22195);
and U24959 (N_24959,N_20482,N_21082);
nor U24960 (N_24960,N_21845,N_22089);
or U24961 (N_24961,N_22172,N_21309);
nor U24962 (N_24962,N_21537,N_20159);
nand U24963 (N_24963,N_21495,N_20724);
nor U24964 (N_24964,N_20292,N_22196);
and U24965 (N_24965,N_21975,N_21458);
xnor U24966 (N_24966,N_21099,N_20144);
or U24967 (N_24967,N_21913,N_20545);
nor U24968 (N_24968,N_21002,N_20710);
or U24969 (N_24969,N_20201,N_20791);
or U24970 (N_24970,N_22200,N_22077);
nand U24971 (N_24971,N_22243,N_21889);
nand U24972 (N_24972,N_21967,N_21937);
or U24973 (N_24973,N_21642,N_21441);
nand U24974 (N_24974,N_21977,N_20677);
nand U24975 (N_24975,N_20808,N_22290);
nor U24976 (N_24976,N_20557,N_20423);
nand U24977 (N_24977,N_22204,N_22133);
or U24978 (N_24978,N_20163,N_21010);
nor U24979 (N_24979,N_21206,N_20167);
nand U24980 (N_24980,N_21303,N_20255);
nor U24981 (N_24981,N_21750,N_20942);
nand U24982 (N_24982,N_21287,N_22286);
nor U24983 (N_24983,N_22093,N_22196);
and U24984 (N_24984,N_22185,N_20986);
nor U24985 (N_24985,N_20692,N_22390);
nand U24986 (N_24986,N_21808,N_20622);
nor U24987 (N_24987,N_20252,N_21888);
nand U24988 (N_24988,N_20735,N_21926);
nand U24989 (N_24989,N_21581,N_21663);
or U24990 (N_24990,N_22155,N_22023);
and U24991 (N_24991,N_21736,N_21561);
nor U24992 (N_24992,N_20583,N_20518);
or U24993 (N_24993,N_22432,N_22330);
nand U24994 (N_24994,N_21156,N_21079);
nor U24995 (N_24995,N_21965,N_21214);
nand U24996 (N_24996,N_21588,N_20765);
nand U24997 (N_24997,N_20917,N_21087);
and U24998 (N_24998,N_20060,N_20619);
or U24999 (N_24999,N_21621,N_20082);
nand UO_0 (O_0,N_22766,N_22700);
and UO_1 (O_1,N_24524,N_24766);
or UO_2 (O_2,N_24367,N_23618);
or UO_3 (O_3,N_24362,N_22997);
xor UO_4 (O_4,N_23249,N_24381);
xnor UO_5 (O_5,N_23104,N_23099);
or UO_6 (O_6,N_22882,N_23125);
and UO_7 (O_7,N_23741,N_24620);
or UO_8 (O_8,N_24857,N_22652);
nand UO_9 (O_9,N_24452,N_23160);
and UO_10 (O_10,N_22611,N_23807);
xor UO_11 (O_11,N_24983,N_22547);
or UO_12 (O_12,N_23823,N_24944);
nand UO_13 (O_13,N_22800,N_22826);
xnor UO_14 (O_14,N_22591,N_24667);
or UO_15 (O_15,N_24969,N_24276);
or UO_16 (O_16,N_23431,N_22880);
nor UO_17 (O_17,N_24936,N_24744);
nand UO_18 (O_18,N_24267,N_24904);
or UO_19 (O_19,N_24769,N_24218);
nand UO_20 (O_20,N_24094,N_24601);
and UO_21 (O_21,N_23810,N_23712);
nand UO_22 (O_22,N_23566,N_24864);
nor UO_23 (O_23,N_24184,N_23325);
nand UO_24 (O_24,N_24631,N_22802);
xor UO_25 (O_25,N_22956,N_24914);
or UO_26 (O_26,N_23707,N_23265);
nor UO_27 (O_27,N_23784,N_24471);
and UO_28 (O_28,N_22955,N_23571);
nand UO_29 (O_29,N_23413,N_24164);
nor UO_30 (O_30,N_24485,N_24678);
and UO_31 (O_31,N_23455,N_23281);
or UO_32 (O_32,N_22847,N_22746);
xnor UO_33 (O_33,N_23392,N_24491);
xor UO_34 (O_34,N_23052,N_23449);
or UO_35 (O_35,N_23148,N_23498);
or UO_36 (O_36,N_22731,N_24968);
and UO_37 (O_37,N_24728,N_22825);
nor UO_38 (O_38,N_23865,N_24836);
nand UO_39 (O_39,N_24210,N_23108);
and UO_40 (O_40,N_22723,N_22674);
xnor UO_41 (O_41,N_23997,N_24294);
or UO_42 (O_42,N_23307,N_24919);
xnor UO_43 (O_43,N_23068,N_22959);
or UO_44 (O_44,N_23857,N_23523);
nor UO_45 (O_45,N_23284,N_24392);
nand UO_46 (O_46,N_23527,N_22508);
and UO_47 (O_47,N_24292,N_24319);
and UO_48 (O_48,N_24438,N_23377);
nand UO_49 (O_49,N_22695,N_22720);
nand UO_50 (O_50,N_24799,N_22898);
or UO_51 (O_51,N_23187,N_24053);
and UO_52 (O_52,N_24913,N_24074);
nand UO_53 (O_53,N_23410,N_23841);
xnor UO_54 (O_54,N_24931,N_23429);
and UO_55 (O_55,N_24802,N_23619);
or UO_56 (O_56,N_22984,N_24593);
or UO_57 (O_57,N_23579,N_24318);
or UO_58 (O_58,N_24693,N_22663);
nor UO_59 (O_59,N_24301,N_22849);
or UO_60 (O_60,N_24499,N_23756);
nor UO_61 (O_61,N_24175,N_23942);
nand UO_62 (O_62,N_24461,N_23897);
or UO_63 (O_63,N_24216,N_23558);
xnor UO_64 (O_64,N_23631,N_23822);
or UO_65 (O_65,N_22922,N_22797);
or UO_66 (O_66,N_24364,N_24529);
nor UO_67 (O_67,N_24776,N_23808);
and UO_68 (O_68,N_23555,N_23594);
and UO_69 (O_69,N_23799,N_22869);
nand UO_70 (O_70,N_22530,N_24596);
and UO_71 (O_71,N_23359,N_24657);
xor UO_72 (O_72,N_24980,N_23920);
or UO_73 (O_73,N_23968,N_24662);
nand UO_74 (O_74,N_23882,N_23507);
and UO_75 (O_75,N_23112,N_22538);
nand UO_76 (O_76,N_23173,N_22706);
and UO_77 (O_77,N_23201,N_23578);
nor UO_78 (O_78,N_24571,N_23445);
nand UO_79 (O_79,N_23022,N_23263);
nand UO_80 (O_80,N_23627,N_24553);
xnor UO_81 (O_81,N_24285,N_23067);
nand UO_82 (O_82,N_22933,N_23870);
nor UO_83 (O_83,N_23460,N_24729);
or UO_84 (O_84,N_22698,N_24345);
or UO_85 (O_85,N_24323,N_23760);
nor UO_86 (O_86,N_24201,N_24955);
and UO_87 (O_87,N_24967,N_22550);
nand UO_88 (O_88,N_23800,N_23098);
nand UO_89 (O_89,N_22954,N_23121);
and UO_90 (O_90,N_24670,N_24421);
nor UO_91 (O_91,N_23157,N_22627);
or UO_92 (O_92,N_24163,N_23257);
and UO_93 (O_93,N_24712,N_23216);
nor UO_94 (O_94,N_23039,N_22743);
nor UO_95 (O_95,N_23399,N_23617);
nand UO_96 (O_96,N_24506,N_23178);
nand UO_97 (O_97,N_22668,N_23541);
and UO_98 (O_98,N_22820,N_24705);
nand UO_99 (O_99,N_23419,N_23574);
or UO_100 (O_100,N_24613,N_24543);
and UO_101 (O_101,N_23341,N_23130);
or UO_102 (O_102,N_23670,N_22981);
and UO_103 (O_103,N_24663,N_24911);
nand UO_104 (O_104,N_24972,N_24756);
nand UO_105 (O_105,N_23412,N_24997);
nor UO_106 (O_106,N_24719,N_24498);
xor UO_107 (O_107,N_23615,N_23169);
nor UO_108 (O_108,N_23418,N_23691);
nor UO_109 (O_109,N_24798,N_22803);
nor UO_110 (O_110,N_24668,N_23451);
and UO_111 (O_111,N_23535,N_23883);
nand UO_112 (O_112,N_24054,N_24055);
and UO_113 (O_113,N_24896,N_22588);
or UO_114 (O_114,N_22564,N_24797);
and UO_115 (O_115,N_24343,N_24040);
nor UO_116 (O_116,N_24658,N_24125);
or UO_117 (O_117,N_23006,N_23759);
and UO_118 (O_118,N_22541,N_24328);
nor UO_119 (O_119,N_22560,N_22514);
and UO_120 (O_120,N_22689,N_23790);
nand UO_121 (O_121,N_22761,N_24628);
nand UO_122 (O_122,N_23363,N_24770);
nor UO_123 (O_123,N_23016,N_22991);
nor UO_124 (O_124,N_24420,N_24469);
and UO_125 (O_125,N_23300,N_24066);
nand UO_126 (O_126,N_23466,N_23013);
nand UO_127 (O_127,N_24274,N_23980);
and UO_128 (O_128,N_24189,N_24107);
or UO_129 (O_129,N_24299,N_24023);
or UO_130 (O_130,N_24653,N_24611);
nand UO_131 (O_131,N_22865,N_24166);
nor UO_132 (O_132,N_24260,N_22783);
and UO_133 (O_133,N_23329,N_23755);
nand UO_134 (O_134,N_24211,N_23547);
or UO_135 (O_135,N_23672,N_22604);
nor UO_136 (O_136,N_23398,N_24355);
nor UO_137 (O_137,N_23671,N_23908);
and UO_138 (O_138,N_24500,N_23308);
nand UO_139 (O_139,N_24960,N_23040);
xnor UO_140 (O_140,N_22905,N_23516);
xor UO_141 (O_141,N_22819,N_23838);
nand UO_142 (O_142,N_24924,N_24807);
and UO_143 (O_143,N_23389,N_24632);
nor UO_144 (O_144,N_24140,N_22975);
nand UO_145 (O_145,N_24818,N_22918);
and UO_146 (O_146,N_24856,N_23322);
nand UO_147 (O_147,N_23351,N_24196);
and UO_148 (O_148,N_24929,N_24002);
nand UO_149 (O_149,N_22691,N_22754);
xnor UO_150 (O_150,N_23888,N_23261);
nand UO_151 (O_151,N_24158,N_23681);
xor UO_152 (O_152,N_23368,N_23060);
or UO_153 (O_153,N_23030,N_24021);
or UO_154 (O_154,N_22597,N_23312);
and UO_155 (O_155,N_23791,N_23331);
nor UO_156 (O_156,N_24519,N_23306);
nand UO_157 (O_157,N_22718,N_24338);
xor UO_158 (O_158,N_23590,N_23962);
and UO_159 (O_159,N_22598,N_23628);
or UO_160 (O_160,N_24441,N_24949);
nor UO_161 (O_161,N_24081,N_22528);
or UO_162 (O_162,N_23131,N_22777);
or UO_163 (O_163,N_23669,N_22586);
and UO_164 (O_164,N_23752,N_24759);
xnor UO_165 (O_165,N_23051,N_23666);
nor UO_166 (O_166,N_24775,N_23115);
nor UO_167 (O_167,N_24677,N_23745);
nand UO_168 (O_168,N_24999,N_23927);
nand UO_169 (O_169,N_23336,N_24783);
xor UO_170 (O_170,N_24224,N_23236);
nand UO_171 (O_171,N_23544,N_23387);
nor UO_172 (O_172,N_22793,N_23995);
or UO_173 (O_173,N_22733,N_24892);
and UO_174 (O_174,N_22737,N_23711);
nand UO_175 (O_175,N_23821,N_24534);
nand UO_176 (O_176,N_24626,N_23373);
and UO_177 (O_177,N_24730,N_22934);
and UO_178 (O_178,N_24116,N_23630);
nand UO_179 (O_179,N_24872,N_23948);
nor UO_180 (O_180,N_23901,N_24724);
nand UO_181 (O_181,N_24089,N_23285);
and UO_182 (O_182,N_23436,N_24223);
or UO_183 (O_183,N_24808,N_23459);
or UO_184 (O_184,N_24935,N_23798);
nand UO_185 (O_185,N_22928,N_22549);
or UO_186 (O_186,N_23520,N_22705);
and UO_187 (O_187,N_24739,N_23975);
xnor UO_188 (O_188,N_23018,N_24246);
nor UO_189 (O_189,N_24429,N_24098);
nand UO_190 (O_190,N_23046,N_22608);
nand UO_191 (O_191,N_24105,N_24225);
and UO_192 (O_192,N_24878,N_24120);
nor UO_193 (O_193,N_23082,N_24778);
nor UO_194 (O_194,N_24639,N_23254);
or UO_195 (O_195,N_23977,N_23710);
and UO_196 (O_196,N_24346,N_22730);
nand UO_197 (O_197,N_22799,N_24995);
nor UO_198 (O_198,N_23999,N_23182);
or UO_199 (O_199,N_24974,N_22864);
and UO_200 (O_200,N_24630,N_24638);
and UO_201 (O_201,N_23369,N_23251);
and UO_202 (O_202,N_24232,N_23550);
nor UO_203 (O_203,N_23945,N_23388);
or UO_204 (O_204,N_24956,N_23003);
xor UO_205 (O_205,N_24520,N_23963);
xor UO_206 (O_206,N_24834,N_23593);
and UO_207 (O_207,N_24597,N_23526);
xnor UO_208 (O_208,N_23514,N_23483);
and UO_209 (O_209,N_23071,N_24684);
nand UO_210 (O_210,N_22949,N_24170);
nand UO_211 (O_211,N_22707,N_23867);
nand UO_212 (O_212,N_24689,N_24333);
or UO_213 (O_213,N_23044,N_24371);
nand UO_214 (O_214,N_23026,N_24265);
and UO_215 (O_215,N_24503,N_24888);
nand UO_216 (O_216,N_23836,N_23873);
nand UO_217 (O_217,N_22909,N_24350);
or UO_218 (O_218,N_23894,N_24548);
xnor UO_219 (O_219,N_23402,N_22632);
nor UO_220 (O_220,N_24028,N_24061);
nor UO_221 (O_221,N_24194,N_22908);
nor UO_222 (O_222,N_22522,N_23480);
nor UO_223 (O_223,N_23849,N_23645);
nor UO_224 (O_224,N_22995,N_23903);
nand UO_225 (O_225,N_24942,N_24477);
nor UO_226 (O_226,N_24005,N_22937);
and UO_227 (O_227,N_22584,N_24372);
and UO_228 (O_228,N_24239,N_23657);
or UO_229 (O_229,N_23253,N_24157);
and UO_230 (O_230,N_23358,N_22839);
or UO_231 (O_231,N_24365,N_22968);
nand UO_232 (O_232,N_23879,N_24727);
or UO_233 (O_233,N_22545,N_22506);
nand UO_234 (O_234,N_23232,N_24281);
nand UO_235 (O_235,N_22626,N_23311);
and UO_236 (O_236,N_23946,N_24137);
and UO_237 (O_237,N_22688,N_23802);
and UO_238 (O_238,N_23585,N_24533);
nand UO_239 (O_239,N_24736,N_23910);
nor UO_240 (O_240,N_24746,N_24505);
or UO_241 (O_241,N_22989,N_24191);
nand UO_242 (O_242,N_24612,N_23912);
nand UO_243 (O_243,N_22844,N_24457);
nand UO_244 (O_244,N_24110,N_23083);
and UO_245 (O_245,N_24099,N_23215);
nor UO_246 (O_246,N_24743,N_23106);
nand UO_247 (O_247,N_23620,N_23172);
nor UO_248 (O_248,N_24868,N_23699);
and UO_249 (O_249,N_23180,N_23592);
nor UO_250 (O_250,N_24045,N_23159);
and UO_251 (O_251,N_23393,N_24255);
and UO_252 (O_252,N_24261,N_24322);
and UO_253 (O_253,N_24288,N_23993);
and UO_254 (O_254,N_24873,N_24947);
and UO_255 (O_255,N_24212,N_23414);
and UO_256 (O_256,N_22690,N_24447);
or UO_257 (O_257,N_22916,N_23610);
xor UO_258 (O_258,N_23260,N_23496);
nor UO_259 (O_259,N_23063,N_24829);
or UO_260 (O_260,N_24656,N_24444);
nor UO_261 (O_261,N_24027,N_23887);
xnor UO_262 (O_262,N_23646,N_23080);
nand UO_263 (O_263,N_24101,N_24207);
nand UO_264 (O_264,N_23549,N_24111);
nor UO_265 (O_265,N_24794,N_23509);
nand UO_266 (O_266,N_22500,N_24400);
nor UO_267 (O_267,N_24235,N_23890);
and UO_268 (O_268,N_22517,N_23581);
nor UO_269 (O_269,N_24310,N_23056);
and UO_270 (O_270,N_24877,N_23066);
nand UO_271 (O_271,N_23685,N_24708);
nand UO_272 (O_272,N_23538,N_23757);
or UO_273 (O_273,N_22576,N_24238);
nand UO_274 (O_274,N_24011,N_23939);
nor UO_275 (O_275,N_23833,N_24710);
nor UO_276 (O_276,N_24483,N_23575);
or UO_277 (O_277,N_24900,N_23835);
and UO_278 (O_278,N_23220,N_22906);
xor UO_279 (O_279,N_23270,N_23851);
xor UO_280 (O_280,N_23047,N_22829);
nor UO_281 (O_281,N_24419,N_23837);
or UO_282 (O_282,N_23881,N_24046);
nor UO_283 (O_283,N_23844,N_24915);
nand UO_284 (O_284,N_23668,N_23729);
nand UO_285 (O_285,N_24965,N_23421);
or UO_286 (O_286,N_22902,N_23828);
and UO_287 (O_287,N_23111,N_23053);
nor UO_288 (O_288,N_22628,N_23622);
and UO_289 (O_289,N_24633,N_24622);
or UO_290 (O_290,N_22926,N_23295);
or UO_291 (O_291,N_24380,N_23097);
and UO_292 (O_292,N_23806,N_23477);
or UO_293 (O_293,N_24556,N_23102);
nor UO_294 (O_294,N_22570,N_24405);
nand UO_295 (O_295,N_23124,N_23994);
or UO_296 (O_296,N_24298,N_23689);
nand UO_297 (O_297,N_24898,N_24792);
and UO_298 (O_298,N_22780,N_24476);
and UO_299 (O_299,N_23986,N_23139);
nor UO_300 (O_300,N_22866,N_24479);
nor UO_301 (O_301,N_22927,N_24474);
or UO_302 (O_302,N_22610,N_22595);
or UO_303 (O_303,N_23726,N_24314);
and UO_304 (O_304,N_23580,N_22838);
and UO_305 (O_305,N_22919,N_24145);
nor UO_306 (O_306,N_23568,N_22810);
nand UO_307 (O_307,N_23156,N_23588);
nand UO_308 (O_308,N_23788,N_23589);
and UO_309 (O_309,N_22562,N_22816);
nor UO_310 (O_310,N_23120,N_22646);
and UO_311 (O_311,N_24160,N_24817);
xnor UO_312 (O_312,N_23562,N_24984);
or UO_313 (O_313,N_22603,N_24773);
and UO_314 (O_314,N_23551,N_24609);
and UO_315 (O_315,N_22682,N_22563);
or UO_316 (O_316,N_24991,N_24713);
and UO_317 (O_317,N_23057,N_23599);
nor UO_318 (O_318,N_24692,N_24490);
and UO_319 (O_319,N_23330,N_22565);
nor UO_320 (O_320,N_23352,N_24927);
nor UO_321 (O_321,N_24825,N_22684);
nor UO_322 (O_322,N_24197,N_24654);
and UO_323 (O_323,N_24777,N_24020);
nor UO_324 (O_324,N_23787,N_24006);
nor UO_325 (O_325,N_23292,N_23983);
and UO_326 (O_326,N_24414,N_24340);
or UO_327 (O_327,N_23676,N_24425);
and UO_328 (O_328,N_23227,N_22813);
and UO_329 (O_329,N_23815,N_22579);
nor UO_330 (O_330,N_24015,N_24574);
xor UO_331 (O_331,N_23248,N_22913);
or UO_332 (O_332,N_23716,N_23383);
nor UO_333 (O_333,N_24665,N_24180);
nor UO_334 (O_334,N_22873,N_22917);
nor UO_335 (O_335,N_23959,N_23635);
and UO_336 (O_336,N_22868,N_24789);
nor UO_337 (O_337,N_24649,N_22791);
or UO_338 (O_338,N_24354,N_22987);
and UO_339 (O_339,N_23442,N_22725);
nor UO_340 (O_340,N_24208,N_23332);
nor UO_341 (O_341,N_23043,N_24375);
and UO_342 (O_342,N_22701,N_24680);
xor UO_343 (O_343,N_23033,N_24215);
or UO_344 (O_344,N_24567,N_24791);
and UO_345 (O_345,N_23456,N_24268);
or UO_346 (O_346,N_24643,N_23258);
or UO_347 (O_347,N_23843,N_24455);
nor UO_348 (O_348,N_24240,N_23259);
nand UO_349 (O_349,N_23817,N_22834);
or UO_350 (O_350,N_23397,N_23048);
nor UO_351 (O_351,N_22967,N_22654);
or UO_352 (O_352,N_23086,N_22711);
and UO_353 (O_353,N_23448,N_23665);
or UO_354 (O_354,N_24565,N_24008);
or UO_355 (O_355,N_24738,N_23170);
or UO_356 (O_356,N_22828,N_24645);
xor UO_357 (O_357,N_24859,N_22601);
nor UO_358 (O_358,N_22687,N_24587);
xor UO_359 (O_359,N_24547,N_23722);
and UO_360 (O_360,N_23636,N_22861);
or UO_361 (O_361,N_24109,N_24026);
nor UO_362 (O_362,N_23167,N_23205);
or UO_363 (O_363,N_23548,N_24104);
and UO_364 (O_364,N_24417,N_23027);
and UO_365 (O_365,N_24122,N_23423);
nor UO_366 (O_366,N_23395,N_23639);
and UO_367 (O_367,N_24183,N_23437);
and UO_368 (O_368,N_24249,N_22534);
xor UO_369 (O_369,N_23471,N_23877);
nor UO_370 (O_370,N_24150,N_22750);
and UO_371 (O_371,N_22693,N_24161);
or UO_372 (O_372,N_23805,N_24386);
or UO_373 (O_373,N_24233,N_24466);
xnor UO_374 (O_374,N_22719,N_23545);
nand UO_375 (O_375,N_24714,N_24056);
or UO_376 (O_376,N_23014,N_23853);
nand UO_377 (O_377,N_24932,N_24361);
or UO_378 (O_378,N_23749,N_24711);
or UO_379 (O_379,N_24787,N_22842);
nor UO_380 (O_380,N_24703,N_23296);
or UO_381 (O_381,N_23797,N_22501);
nand UO_382 (O_382,N_24939,N_24404);
nor UO_383 (O_383,N_22726,N_23528);
nand UO_384 (O_384,N_23382,N_23113);
nand UO_385 (O_385,N_24732,N_23486);
nor UO_386 (O_386,N_24749,N_23206);
nand UO_387 (O_387,N_23793,N_24229);
xor UO_388 (O_388,N_24895,N_22557);
nor UO_389 (O_389,N_24492,N_23958);
or UO_390 (O_390,N_24273,N_24774);
or UO_391 (O_391,N_22827,N_23441);
xnor UO_392 (O_392,N_23064,N_23290);
or UO_393 (O_393,N_23081,N_24300);
or UO_394 (O_394,N_22655,N_24092);
and UO_395 (O_395,N_23702,N_24443);
or UO_396 (O_396,N_24848,N_23354);
nor UO_397 (O_397,N_23557,N_23366);
xor UO_398 (O_398,N_23282,N_24847);
and UO_399 (O_399,N_24606,N_23976);
or UO_400 (O_400,N_24540,N_23655);
and UO_401 (O_401,N_23225,N_23416);
nand UO_402 (O_402,N_23433,N_23467);
or UO_403 (O_403,N_23381,N_22516);
and UO_404 (O_404,N_24188,N_23374);
nor UO_405 (O_405,N_23342,N_23186);
nand UO_406 (O_406,N_23758,N_23250);
or UO_407 (O_407,N_23061,N_24874);
nand UO_408 (O_408,N_24644,N_23476);
xnor UO_409 (O_409,N_22985,N_24494);
or UO_410 (O_410,N_24031,N_22753);
and UO_411 (O_411,N_23177,N_23280);
nor UO_412 (O_412,N_23001,N_23109);
and UO_413 (O_413,N_23733,N_24963);
and UO_414 (O_414,N_22769,N_24961);
xor UO_415 (O_415,N_24673,N_24341);
xnor UO_416 (O_416,N_22872,N_24866);
and UO_417 (O_417,N_22596,N_24854);
nor UO_418 (O_418,N_24504,N_23629);
nor UO_419 (O_419,N_24394,N_22554);
nand UO_420 (O_420,N_24979,N_24403);
nor UO_421 (O_421,N_22992,N_24259);
and UO_422 (O_422,N_24190,N_24342);
nor UO_423 (O_423,N_24128,N_22823);
xor UO_424 (O_424,N_24762,N_23244);
nand UO_425 (O_425,N_24366,N_24432);
nand UO_426 (O_426,N_23361,N_24379);
or UO_427 (O_427,N_23319,N_23973);
nor UO_428 (O_428,N_23192,N_23041);
and UO_429 (O_429,N_22551,N_22912);
nor UO_430 (O_430,N_23776,N_23337);
xor UO_431 (O_431,N_24785,N_23773);
nor UO_432 (O_432,N_23531,N_24538);
nor UO_433 (O_433,N_24688,N_24112);
nand UO_434 (O_434,N_23482,N_22634);
and UO_435 (O_435,N_23904,N_24509);
and UO_436 (O_436,N_23967,N_24025);
xnor UO_437 (O_437,N_23819,N_22644);
nand UO_438 (O_438,N_22676,N_22870);
and UO_439 (O_439,N_24508,N_23735);
and UO_440 (O_440,N_23700,N_23534);
or UO_441 (O_441,N_22589,N_24831);
and UO_442 (O_442,N_23885,N_23871);
nor UO_443 (O_443,N_22573,N_24347);
nand UO_444 (O_444,N_24735,N_22567);
or UO_445 (O_445,N_24659,N_24861);
and UO_446 (O_446,N_24754,N_23786);
and UO_447 (O_447,N_24209,N_23469);
nor UO_448 (O_448,N_24182,N_22910);
and UO_449 (O_449,N_23789,N_24591);
nor UO_450 (O_450,N_22890,N_23969);
or UO_451 (O_451,N_23166,N_23780);
nor UO_452 (O_452,N_22856,N_24162);
nor UO_453 (O_453,N_24399,N_23911);
xor UO_454 (O_454,N_24839,N_22858);
nand UO_455 (O_455,N_22936,N_23211);
or UO_456 (O_456,N_24069,N_22637);
and UO_457 (O_457,N_23002,N_24852);
nor UO_458 (O_458,N_22831,N_22709);
nor UO_459 (O_459,N_24132,N_23502);
and UO_460 (O_460,N_23847,N_22854);
nand UO_461 (O_461,N_23127,N_24875);
and UO_462 (O_462,N_23091,N_23443);
xnor UO_463 (O_463,N_24842,N_24472);
nand UO_464 (O_464,N_24072,N_24153);
nor UO_465 (O_465,N_24683,N_24022);
xnor UO_466 (O_466,N_23134,N_23661);
nor UO_467 (O_467,N_22548,N_22620);
nand UO_468 (O_468,N_24515,N_23597);
or UO_469 (O_469,N_22921,N_23537);
or UO_470 (O_470,N_23077,N_23126);
or UO_471 (O_471,N_23649,N_22607);
or UO_472 (O_472,N_22886,N_24755);
nand UO_473 (O_473,N_22785,N_23768);
xor UO_474 (O_474,N_22511,N_24855);
and UO_475 (O_475,N_22990,N_24369);
and UO_476 (O_476,N_24058,N_24812);
or UO_477 (O_477,N_23154,N_23829);
nor UO_478 (O_478,N_24236,N_22961);
and UO_479 (O_479,N_24635,N_23659);
nor UO_480 (O_480,N_22901,N_23899);
and UO_481 (O_481,N_24652,N_24248);
nand UO_482 (O_482,N_23428,N_23898);
nor UO_483 (O_483,N_23000,N_23567);
nand UO_484 (O_484,N_23379,N_24998);
or UO_485 (O_485,N_22680,N_24966);
and UO_486 (O_486,N_22845,N_23652);
nor UO_487 (O_487,N_24199,N_22764);
nand UO_488 (O_488,N_23637,N_24819);
nor UO_489 (O_489,N_24569,N_24747);
and UO_490 (O_490,N_23065,N_24115);
nand UO_491 (O_491,N_24167,N_22679);
nor UO_492 (O_492,N_24370,N_22657);
nand UO_493 (O_493,N_22848,N_23987);
and UO_494 (O_494,N_23695,N_24204);
nand UO_495 (O_495,N_23454,N_23078);
or UO_496 (O_496,N_24296,N_22630);
nor UO_497 (O_497,N_24992,N_23328);
and UO_498 (O_498,N_22945,N_24390);
nor UO_499 (O_499,N_24526,N_22840);
nor UO_500 (O_500,N_22552,N_24741);
and UO_501 (O_501,N_23090,N_22553);
or UO_502 (O_502,N_22738,N_22837);
nor UO_503 (O_503,N_23444,N_24679);
or UO_504 (O_504,N_24742,N_24496);
nor UO_505 (O_505,N_22786,N_22580);
and UO_506 (O_506,N_24846,N_24493);
nor UO_507 (O_507,N_24971,N_22804);
nand UO_508 (O_508,N_23075,N_23050);
nor UO_509 (O_509,N_23662,N_22772);
nor UO_510 (O_510,N_24784,N_23434);
and UO_511 (O_511,N_24975,N_24993);
xnor UO_512 (O_512,N_24087,N_24605);
xor UO_513 (O_513,N_24962,N_24412);
nand UO_514 (O_514,N_22867,N_24849);
nand UO_515 (O_515,N_23029,N_23407);
and UO_516 (O_516,N_23918,N_24687);
nor UO_517 (O_517,N_22675,N_22544);
nor UO_518 (O_518,N_23188,N_24303);
nor UO_519 (O_519,N_23651,N_24253);
nor UO_520 (O_520,N_24725,N_22556);
nand UO_521 (O_521,N_23974,N_24803);
nor UO_522 (O_522,N_23252,N_23136);
and UO_523 (O_523,N_23561,N_24697);
and UO_524 (O_524,N_23680,N_24353);
nor UO_525 (O_525,N_24213,N_24720);
nor UO_526 (O_526,N_24907,N_22980);
or UO_527 (O_527,N_24007,N_24287);
nor UO_528 (O_528,N_23852,N_23876);
or UO_529 (O_529,N_24095,N_24332);
or UO_530 (O_530,N_22685,N_24518);
nor UO_531 (O_531,N_23915,N_24431);
nor UO_532 (O_532,N_24804,N_22817);
nor UO_533 (O_533,N_23404,N_23922);
nand UO_534 (O_534,N_23005,N_22796);
and UO_535 (O_535,N_23219,N_24060);
and UO_536 (O_536,N_24275,N_24758);
or UO_537 (O_537,N_24449,N_23742);
and UO_538 (O_538,N_24573,N_24726);
nor UO_539 (O_539,N_23706,N_24013);
nand UO_540 (O_540,N_24651,N_24378);
and UO_541 (O_541,N_23036,N_24717);
or UO_542 (O_542,N_23769,N_24306);
nand UO_543 (O_543,N_24464,N_24114);
nor UO_544 (O_544,N_24507,N_24393);
nor UO_545 (O_545,N_23990,N_22943);
nor UO_546 (O_546,N_24925,N_24460);
nor UO_547 (O_547,N_22852,N_24634);
or UO_548 (O_548,N_24138,N_22636);
and UO_549 (O_549,N_23274,N_23334);
nor UO_550 (O_550,N_24359,N_24897);
nor UO_551 (O_551,N_23357,N_23644);
or UO_552 (O_552,N_23465,N_24594);
nand UO_553 (O_553,N_22510,N_23724);
nor UO_554 (O_554,N_23647,N_24793);
xor UO_555 (O_555,N_23656,N_24551);
nor UO_556 (O_556,N_24241,N_22649);
and UO_557 (O_557,N_22794,N_22892);
nor UO_558 (O_558,N_23826,N_24416);
or UO_559 (O_559,N_22950,N_22536);
nand UO_560 (O_560,N_24172,N_24484);
nor UO_561 (O_561,N_23582,N_24149);
nand UO_562 (O_562,N_24090,N_24871);
nor UO_563 (O_563,N_23554,N_24753);
nor UO_564 (O_564,N_24675,N_23155);
and UO_565 (O_565,N_24771,N_22694);
nand UO_566 (O_566,N_24428,N_23504);
xnor UO_567 (O_567,N_24462,N_22960);
nor UO_568 (O_568,N_23966,N_23746);
or UO_569 (O_569,N_23648,N_22749);
nand UO_570 (O_570,N_24602,N_22645);
nand UO_571 (O_571,N_22914,N_23577);
nand UO_572 (O_572,N_24168,N_24501);
nor UO_573 (O_573,N_23088,N_24280);
xnor UO_574 (O_574,N_24445,N_23035);
and UO_575 (O_575,N_22763,N_24179);
and UO_576 (O_576,N_23770,N_24243);
or UO_577 (O_577,N_24050,N_23505);
xnor UO_578 (O_578,N_22519,N_24134);
xor UO_579 (O_579,N_22899,N_23430);
or UO_580 (O_580,N_23623,N_24311);
xor UO_581 (O_581,N_23089,N_23074);
nor UO_582 (O_582,N_22824,N_22535);
xnor UO_583 (O_583,N_24699,N_23982);
or UO_584 (O_584,N_24262,N_24901);
and UO_585 (O_585,N_24603,N_23117);
nor UO_586 (O_586,N_24822,N_23279);
nand UO_587 (O_587,N_23344,N_24256);
or UO_588 (O_588,N_23930,N_23426);
nor UO_589 (O_589,N_24143,N_23693);
nor UO_590 (O_590,N_23417,N_23264);
or UO_591 (O_591,N_23149,N_24977);
xnor UO_592 (O_592,N_23608,N_22953);
and UO_593 (O_593,N_23586,N_23150);
nand UO_594 (O_594,N_23730,N_23923);
or UO_595 (O_595,N_24850,N_23750);
nand UO_596 (O_596,N_23391,N_23515);
or UO_597 (O_597,N_24790,N_23935);
and UO_598 (O_598,N_22665,N_24250);
or UO_599 (O_599,N_23521,N_23940);
nand UO_600 (O_600,N_22504,N_24254);
nand UO_601 (O_601,N_22613,N_23390);
or UO_602 (O_602,N_23493,N_23869);
and UO_603 (O_603,N_23019,N_24203);
or UO_604 (O_604,N_23536,N_24044);
xnor UO_605 (O_605,N_24513,N_22559);
or UO_606 (O_606,N_22923,N_22713);
nor UO_607 (O_607,N_23721,N_23909);
or UO_608 (O_608,N_24843,N_24497);
or UO_609 (O_609,N_24557,N_24707);
or UO_610 (O_610,N_24862,N_24813);
nand UO_611 (O_611,N_22821,N_24408);
nand UO_612 (O_612,N_24502,N_24811);
nor UO_613 (O_613,N_24108,N_23985);
and UO_614 (O_614,N_24385,N_23664);
nor UO_615 (O_615,N_23560,N_23801);
nand UO_616 (O_616,N_24851,N_24217);
xor UO_617 (O_617,N_23949,N_22759);
nor UO_618 (O_618,N_22808,N_22656);
and UO_619 (O_619,N_24033,N_23316);
nand UO_620 (O_620,N_22774,N_23553);
or UO_621 (O_621,N_24302,N_22715);
nor UO_622 (O_622,N_23093,N_22893);
xnor UO_623 (O_623,N_23591,N_23473);
and UO_624 (O_624,N_23937,N_23289);
nor UO_625 (O_625,N_24478,N_23234);
and UO_626 (O_626,N_24820,N_23525);
nor UO_627 (O_627,N_22686,N_24934);
nor UO_628 (O_628,N_23424,N_24616);
nor UO_629 (O_629,N_23287,N_22702);
nand UO_630 (O_630,N_24159,N_23860);
nor UO_631 (O_631,N_23011,N_23291);
xnor UO_632 (O_632,N_23440,N_23778);
or UO_633 (O_633,N_24660,N_24142);
nor UO_634 (O_634,N_22736,N_23340);
xnor UO_635 (O_635,N_24827,N_24946);
nand UO_636 (O_636,N_22879,N_24139);
nor UO_637 (O_637,N_23116,N_24070);
or UO_638 (O_638,N_24706,N_24899);
or UO_639 (O_639,N_24097,N_23438);
or UO_640 (O_640,N_24981,N_23499);
or UO_641 (O_641,N_23100,N_24357);
and UO_642 (O_642,N_23501,N_23223);
xnor UO_643 (O_643,N_23427,N_23497);
and UO_644 (O_644,N_23638,N_24650);
or UO_645 (O_645,N_24124,N_24082);
or UO_646 (O_646,N_22537,N_23954);
or UO_647 (O_647,N_22904,N_24989);
or UO_648 (O_648,N_23032,N_22907);
and UO_649 (O_649,N_23266,N_23191);
xnor UO_650 (O_650,N_22734,N_24959);
or UO_651 (O_651,N_24721,N_23552);
or UO_652 (O_652,N_23235,N_24470);
or UO_653 (O_653,N_22818,N_24376);
and UO_654 (O_654,N_24051,N_23133);
and UO_655 (O_655,N_23846,N_22582);
nor UO_656 (O_656,N_23642,N_24075);
nor UO_657 (O_657,N_22957,N_24331);
and UO_658 (O_658,N_23380,N_22739);
and UO_659 (O_659,N_23479,N_23513);
nor UO_660 (O_660,N_23703,N_22973);
or UO_661 (O_661,N_23231,N_23240);
and UO_662 (O_662,N_24102,N_24589);
nand UO_663 (O_663,N_24186,N_24251);
nand UO_664 (O_664,N_22599,N_23105);
or UO_665 (O_665,N_23868,N_23247);
nand UO_666 (O_666,N_22640,N_24561);
and UO_667 (O_667,N_23612,N_23489);
nor UO_668 (O_668,N_23813,N_24284);
nand UO_669 (O_669,N_24468,N_22729);
xor UO_670 (O_670,N_23293,N_24800);
nand UO_671 (O_671,N_23613,N_23401);
nand UO_672 (O_672,N_24828,N_24398);
nand UO_673 (O_673,N_24387,N_24550);
or UO_674 (O_674,N_24325,N_23095);
and UO_675 (O_675,N_24305,N_22875);
nor UO_676 (O_676,N_23228,N_23796);
nor UO_677 (O_677,N_23570,N_22585);
or UO_678 (O_678,N_24448,N_24313);
or UO_679 (O_679,N_24751,N_22716);
or UO_680 (O_680,N_23195,N_24442);
nand UO_681 (O_681,N_22895,N_24317);
nor UO_682 (O_682,N_22658,N_23348);
or UO_683 (O_683,N_23378,N_23272);
or UO_684 (O_684,N_23811,N_24948);
xnor UO_685 (O_685,N_23971,N_22773);
and UO_686 (O_686,N_24978,N_22767);
or UO_687 (O_687,N_24903,N_24205);
nor UO_688 (O_688,N_23171,N_24568);
nor UO_689 (O_689,N_23422,N_24908);
nor UO_690 (O_690,N_23326,N_22938);
or UO_691 (O_691,N_24352,N_23917);
or UO_692 (O_692,N_23572,N_23267);
or UO_693 (O_693,N_23238,N_22851);
or UO_694 (O_694,N_23094,N_23174);
and UO_695 (O_695,N_23569,N_22946);
xor UO_696 (O_696,N_24001,N_23732);
nor UO_697 (O_697,N_24024,N_24552);
and UO_698 (O_698,N_24067,N_24655);
and UO_699 (O_699,N_24244,N_23007);
and UO_700 (O_700,N_24018,N_24185);
or UO_701 (O_701,N_24277,N_24032);
or UO_702 (O_702,N_23185,N_22647);
or UO_703 (O_703,N_22801,N_23543);
or UO_704 (O_704,N_23747,N_24129);
and UO_705 (O_705,N_24330,N_24113);
or UO_706 (O_706,N_22653,N_23744);
and UO_707 (O_707,N_23305,N_23394);
xnor UO_708 (O_708,N_23533,N_23861);
or UO_709 (O_709,N_24321,N_24702);
nand UO_710 (O_710,N_24360,N_24590);
nor UO_711 (O_711,N_24278,N_23302);
nor UO_712 (O_712,N_24544,N_24401);
nand UO_713 (O_713,N_23928,N_23643);
and UO_714 (O_714,N_23667,N_24835);
and UO_715 (O_715,N_23884,N_23435);
nand UO_716 (O_716,N_24976,N_23362);
or UO_717 (O_717,N_23951,N_23425);
or UO_718 (O_718,N_22815,N_23978);
xnor UO_719 (O_719,N_23199,N_24402);
or UO_720 (O_720,N_22742,N_22859);
or UO_721 (O_721,N_24079,N_23965);
nand UO_722 (O_722,N_24648,N_24943);
or UO_723 (O_723,N_24062,N_24853);
nor UO_724 (O_724,N_23283,N_24384);
or UO_725 (O_725,N_22569,N_23848);
nand UO_726 (O_726,N_24614,N_23938);
nor UO_727 (O_727,N_22670,N_24272);
and UO_728 (O_728,N_22533,N_22941);
and UO_729 (O_729,N_23529,N_23237);
and UO_730 (O_730,N_24495,N_23010);
or UO_731 (O_731,N_23107,N_22571);
nor UO_732 (O_732,N_23468,N_23481);
xnor UO_733 (O_733,N_22692,N_23677);
xnor UO_734 (O_734,N_24076,N_22677);
nand UO_735 (O_735,N_23210,N_23370);
and UO_736 (O_736,N_23346,N_22546);
nand UO_737 (O_737,N_23564,N_24564);
or UO_738 (O_738,N_23137,N_22770);
or UO_739 (O_739,N_23145,N_23122);
and UO_740 (O_740,N_23840,N_23487);
or UO_741 (O_741,N_22789,N_24902);
nand UO_742 (O_742,N_24063,N_23988);
nor UO_743 (O_743,N_24865,N_22661);
and UO_744 (O_744,N_23317,N_24566);
nand UO_745 (O_745,N_23653,N_23017);
nand UO_746 (O_746,N_23415,N_22724);
xnor UO_747 (O_747,N_23488,N_23246);
and UO_748 (O_748,N_24234,N_23886);
nand UO_749 (O_749,N_24765,N_24237);
nand UO_750 (O_750,N_23992,N_24135);
nor UO_751 (O_751,N_23510,N_24917);
and UO_752 (O_752,N_24320,N_23165);
nor UO_753 (O_753,N_23834,N_24572);
or UO_754 (O_754,N_22965,N_24734);
nand UO_755 (O_755,N_24465,N_22830);
nand UO_756 (O_756,N_24779,N_23762);
xnor UO_757 (O_757,N_24487,N_24481);
or UO_758 (O_758,N_23197,N_23614);
nor UO_759 (O_759,N_24423,N_24422);
or UO_760 (O_760,N_22807,N_22540);
nor UO_761 (O_761,N_22521,N_23304);
nor UO_762 (O_762,N_23384,N_22524);
xor UO_763 (O_763,N_24126,N_24270);
and UO_764 (O_764,N_24964,N_24970);
and UO_765 (O_765,N_23385,N_24782);
nor UO_766 (O_766,N_22853,N_22699);
or UO_767 (O_767,N_24723,N_22983);
xnor UO_768 (O_768,N_22986,N_24748);
xor UO_769 (O_769,N_24312,N_22578);
or UO_770 (O_770,N_24869,N_23129);
nand UO_771 (O_771,N_23748,N_23632);
nor UO_772 (O_772,N_24815,N_22678);
or UO_773 (O_773,N_24148,N_22812);
nand UO_774 (O_774,N_23073,N_24672);
or UO_775 (O_775,N_23921,N_23950);
or UO_776 (O_776,N_23004,N_24480);
and UO_777 (O_777,N_23872,N_24951);
nand UO_778 (O_778,N_22811,N_24867);
nor UO_779 (O_779,N_23506,N_24909);
and UO_780 (O_780,N_24539,N_22708);
nor UO_781 (O_781,N_24772,N_23952);
nand UO_782 (O_782,N_23364,N_24467);
nor UO_783 (O_783,N_24068,N_22728);
or UO_784 (O_784,N_24953,N_24629);
or UO_785 (O_785,N_22884,N_24844);
nor UO_786 (O_786,N_22681,N_24617);
xnor UO_787 (O_787,N_24435,N_24041);
xnor UO_788 (O_788,N_23054,N_23832);
and UO_789 (O_789,N_23049,N_24100);
and UO_790 (O_790,N_23714,N_24894);
and UO_791 (O_791,N_23690,N_23889);
nand UO_792 (O_792,N_24034,N_24562);
or UO_793 (O_793,N_22860,N_22523);
nor UO_794 (O_794,N_24433,N_22897);
nor UO_795 (O_795,N_23603,N_23069);
xnor UO_796 (O_796,N_23222,N_24003);
nand UO_797 (O_797,N_22778,N_24763);
nor UO_798 (O_798,N_23715,N_22740);
nor UO_799 (O_799,N_24415,N_23058);
nor UO_800 (O_800,N_24592,N_22755);
and UO_801 (O_801,N_24676,N_23725);
nand UO_802 (O_802,N_24740,N_23179);
nand UO_803 (O_803,N_22744,N_23855);
or UO_804 (O_804,N_23275,N_23727);
or UO_805 (O_805,N_22574,N_23794);
xnor UO_806 (O_806,N_23151,N_22911);
nand UO_807 (O_807,N_24119,N_23850);
and UO_808 (O_808,N_24696,N_24221);
nand UO_809 (O_809,N_23464,N_24531);
and UO_810 (O_810,N_22714,N_23485);
nor UO_811 (O_811,N_24788,N_24334);
and UO_812 (O_812,N_24080,N_23255);
nand UO_813 (O_813,N_24921,N_24377);
nor UO_814 (O_814,N_24030,N_23919);
and UO_815 (O_815,N_23654,N_24860);
or UO_816 (O_816,N_23916,N_22572);
or UO_817 (O_817,N_22809,N_23371);
nand UO_818 (O_818,N_23218,N_24155);
xor UO_819 (O_819,N_24722,N_24271);
or UO_820 (O_820,N_24220,N_23360);
and UO_821 (O_821,N_24088,N_22651);
nor UO_822 (O_822,N_24286,N_22735);
or UO_823 (O_823,N_23704,N_22788);
nor UO_824 (O_824,N_24832,N_24337);
nor UO_825 (O_825,N_24558,N_23914);
or UO_826 (O_826,N_22512,N_23181);
or UO_827 (O_827,N_24816,N_23891);
nor UO_828 (O_828,N_24957,N_22614);
or UO_829 (O_829,N_23737,N_24473);
nand UO_830 (O_830,N_24938,N_24192);
or UO_831 (O_831,N_22758,N_22924);
nand UO_832 (O_832,N_23025,N_22600);
or UO_833 (O_833,N_23692,N_23084);
xor UO_834 (O_834,N_24152,N_24545);
or UO_835 (O_835,N_22532,N_24780);
or UO_836 (O_836,N_23587,N_24181);
nand UO_837 (O_837,N_22741,N_23862);
nor UO_838 (O_838,N_24293,N_24701);
or UO_839 (O_839,N_23602,N_24563);
xnor UO_840 (O_840,N_24882,N_24488);
nand UO_841 (O_841,N_24598,N_24621);
xnor UO_842 (O_842,N_23009,N_22776);
nand UO_843 (O_843,N_22638,N_23208);
nor UO_844 (O_844,N_23142,N_22979);
nand UO_845 (O_845,N_23262,N_23960);
nand UO_846 (O_846,N_24757,N_22625);
nand UO_847 (O_847,N_23101,N_24017);
nor UO_848 (O_848,N_24009,N_24646);
and UO_849 (O_849,N_24640,N_24940);
and UO_850 (O_850,N_24996,N_23321);
nand UO_851 (O_851,N_24413,N_23408);
nor UO_852 (O_852,N_24881,N_24133);
and UO_853 (O_853,N_24910,N_23633);
nand UO_854 (O_854,N_23446,N_24517);
nor UO_855 (O_855,N_22969,N_22672);
or UO_856 (O_856,N_24669,N_22633);
and UO_857 (O_857,N_23511,N_22590);
and UO_858 (O_858,N_24833,N_23583);
or UO_859 (O_859,N_23518,N_23241);
and UO_860 (O_860,N_22998,N_24863);
nand UO_861 (O_861,N_23028,N_23143);
nand UO_862 (O_862,N_23299,N_24388);
nor UO_863 (O_863,N_24339,N_23777);
nor UO_864 (O_864,N_22888,N_23020);
nor UO_865 (O_865,N_23863,N_22727);
or UO_866 (O_866,N_23701,N_23462);
and UO_867 (O_867,N_23761,N_23256);
nor UO_868 (O_868,N_23288,N_24926);
nand UO_869 (O_869,N_23375,N_23447);
nand UO_870 (O_870,N_23309,N_24806);
or UO_871 (O_871,N_23964,N_24588);
and UO_872 (O_872,N_24437,N_24581);
xnor UO_873 (O_873,N_23376,N_23517);
and UO_874 (O_874,N_23301,N_24579);
nand UO_875 (O_875,N_22612,N_23781);
or UO_876 (O_876,N_22539,N_23439);
or UO_877 (O_877,N_23979,N_23697);
nand UO_878 (O_878,N_23313,N_23213);
or UO_879 (O_879,N_23771,N_22964);
xor UO_880 (O_880,N_22889,N_24131);
or UO_881 (O_881,N_24389,N_23559);
nor UO_882 (O_882,N_22894,N_23673);
and UO_883 (O_883,N_22843,N_23634);
nand UO_884 (O_884,N_24463,N_24522);
nand UO_885 (O_885,N_24154,N_22850);
nor UO_886 (O_886,N_23675,N_24283);
nor UO_887 (O_887,N_23042,N_24039);
or UO_888 (O_888,N_24690,N_23119);
and UO_889 (O_889,N_23168,N_23403);
nor UO_890 (O_890,N_23859,N_24549);
and UO_891 (O_891,N_24893,N_23062);
or UO_892 (O_892,N_23763,N_24014);
nor UO_893 (O_893,N_24890,N_23400);
nand UO_894 (O_894,N_22878,N_24037);
or UO_895 (O_895,N_23782,N_23717);
nor UO_896 (O_896,N_23765,N_23338);
or UO_897 (O_897,N_23696,N_22900);
xor UO_898 (O_898,N_22667,N_23345);
xnor UO_899 (O_899,N_23820,N_24391);
nand UO_900 (O_900,N_22515,N_23683);
or UO_901 (O_901,N_22732,N_24356);
nand UO_902 (O_902,N_22932,N_23214);
nor UO_903 (O_903,N_23687,N_23457);
and UO_904 (O_904,N_24512,N_22568);
nor UO_905 (O_905,N_24786,N_24542);
nor UO_906 (O_906,N_23409,N_24920);
or UO_907 (O_907,N_24242,N_22618);
nor UO_908 (O_908,N_23827,N_23941);
xor UO_909 (O_909,N_23984,N_22748);
nand UO_910 (O_910,N_24704,N_24266);
or UO_911 (O_911,N_24700,N_23273);
nand UO_912 (O_912,N_24887,N_24595);
and UO_913 (O_913,N_24745,N_22948);
nand UO_914 (O_914,N_24406,N_22781);
or UO_915 (O_915,N_23406,N_22507);
xnor UO_916 (O_916,N_23576,N_24383);
or UO_917 (O_917,N_24173,N_24666);
nor UO_918 (O_918,N_22660,N_24329);
nor UO_919 (O_919,N_24103,N_23008);
and UO_920 (O_920,N_24165,N_23573);
nor UO_921 (O_921,N_23396,N_24694);
nor UO_922 (O_922,N_23663,N_24876);
nor UO_923 (O_923,N_23405,N_23118);
and UO_924 (O_924,N_23512,N_24269);
nor UO_925 (O_925,N_23494,N_23450);
nand UO_926 (O_926,N_22624,N_24912);
and UO_927 (O_927,N_23556,N_23563);
and UO_928 (O_928,N_24307,N_24584);
nor UO_929 (O_929,N_23347,N_22855);
or UO_930 (O_930,N_23152,N_24123);
and UO_931 (O_931,N_24042,N_22757);
nor UO_932 (O_932,N_22903,N_23079);
nand UO_933 (O_933,N_24824,N_24554);
nand UO_934 (O_934,N_23141,N_24019);
nor UO_935 (O_935,N_23153,N_23432);
nand UO_936 (O_936,N_23864,N_22602);
nor UO_937 (O_937,N_24222,N_24363);
nor UO_938 (O_938,N_23972,N_24575);
nor UO_939 (O_939,N_22782,N_24309);
or UO_940 (O_940,N_24886,N_24826);
and UO_941 (O_941,N_24560,N_24570);
nand UO_942 (O_942,N_23601,N_24546);
nand UO_943 (O_943,N_23135,N_24247);
nand UO_944 (O_944,N_23947,N_22721);
xnor UO_945 (O_945,N_24930,N_22669);
or UO_946 (O_946,N_23686,N_24073);
and UO_947 (O_947,N_22629,N_23804);
nor UO_948 (O_948,N_23845,N_24716);
or UO_949 (O_949,N_24446,N_24230);
and UO_950 (O_950,N_24559,N_23315);
and UO_951 (O_951,N_24219,N_23508);
and UO_952 (O_952,N_24809,N_22760);
or UO_953 (O_953,N_22982,N_23718);
or UO_954 (O_954,N_24527,N_24986);
nand UO_955 (O_955,N_23684,N_24297);
nand UO_956 (O_956,N_22593,N_22896);
xnor UO_957 (O_957,N_24171,N_23103);
or UO_958 (O_958,N_23268,N_24737);
xnor UO_959 (O_959,N_24324,N_23738);
or UO_960 (O_960,N_24475,N_24528);
xor UO_961 (O_961,N_24174,N_24282);
nand UO_962 (O_962,N_22993,N_22951);
nand UO_963 (O_963,N_23226,N_23339);
nor UO_964 (O_964,N_22587,N_23709);
nor UO_965 (O_965,N_24682,N_23059);
and UO_966 (O_966,N_23221,N_23892);
nor UO_967 (O_967,N_22616,N_24176);
and UO_968 (O_968,N_24316,N_23818);
nand UO_969 (O_969,N_24536,N_23998);
and UO_970 (O_970,N_24373,N_24382);
or UO_971 (O_971,N_24973,N_23905);
nand UO_972 (O_972,N_23303,N_23327);
xor UO_973 (O_973,N_23926,N_23475);
and UO_974 (O_974,N_24841,N_24290);
and UO_975 (O_975,N_24661,N_24781);
nand UO_976 (O_976,N_23500,N_22768);
nand UO_977 (O_977,N_23229,N_23458);
or UO_978 (O_978,N_24615,N_23070);
and UO_979 (O_979,N_23764,N_23624);
or UO_980 (O_980,N_24077,N_23766);
nor UO_981 (O_981,N_22915,N_24555);
nand UO_982 (O_982,N_23708,N_24336);
nor UO_983 (O_983,N_23278,N_22958);
or UO_984 (O_984,N_24586,N_22833);
xnor UO_985 (O_985,N_24958,N_24228);
nand UO_986 (O_986,N_23297,N_24004);
nor UO_987 (O_987,N_23194,N_24928);
and UO_988 (O_988,N_22696,N_24200);
and UO_989 (O_989,N_24604,N_24625);
and UO_990 (O_990,N_24624,N_24858);
nand UO_991 (O_991,N_23224,N_24440);
nand UO_992 (O_992,N_23034,N_24681);
and UO_993 (O_993,N_22531,N_22971);
or UO_994 (O_994,N_24837,N_24805);
nor UO_995 (O_995,N_24870,N_22683);
nand UO_996 (O_996,N_24906,N_22621);
or UO_997 (O_997,N_24395,N_22606);
nor UO_998 (O_998,N_23981,N_23350);
xor UO_999 (O_999,N_24396,N_22662);
or UO_1000 (O_1000,N_24454,N_22561);
nand UO_1001 (O_1001,N_24106,N_24291);
or UO_1002 (O_1002,N_23294,N_24486);
nor UO_1003 (O_1003,N_23698,N_23728);
nor UO_1004 (O_1004,N_22666,N_23925);
nand UO_1005 (O_1005,N_23021,N_23193);
or UO_1006 (O_1006,N_24430,N_23754);
nand UO_1007 (O_1007,N_23678,N_22639);
or UO_1008 (O_1008,N_24918,N_23816);
nand UO_1009 (O_1009,N_22877,N_23616);
nor UO_1010 (O_1010,N_22972,N_24151);
nand UO_1011 (O_1011,N_22822,N_24752);
nor UO_1012 (O_1012,N_23606,N_24439);
nand UO_1013 (O_1013,N_24523,N_23989);
xor UO_1014 (O_1014,N_22970,N_22963);
and UO_1015 (O_1015,N_22887,N_23189);
or UO_1016 (O_1016,N_24144,N_23906);
or UO_1017 (O_1017,N_22712,N_22974);
and UO_1018 (O_1018,N_23212,N_22976);
and UO_1019 (O_1019,N_23207,N_23830);
or UO_1020 (O_1020,N_23731,N_23452);
nor UO_1021 (O_1021,N_24641,N_23957);
nor UO_1022 (O_1022,N_23854,N_23739);
nor UO_1023 (O_1023,N_24086,N_23679);
nor UO_1024 (O_1024,N_24016,N_23072);
or UO_1025 (O_1025,N_23243,N_23814);
and UO_1026 (O_1026,N_22642,N_23184);
nand UO_1027 (O_1027,N_22929,N_24583);
nand UO_1028 (O_1028,N_23539,N_23641);
or UO_1029 (O_1029,N_23933,N_23783);
and UO_1030 (O_1030,N_24537,N_24418);
and UO_1031 (O_1031,N_23196,N_24600);
and UO_1032 (O_1032,N_23318,N_24685);
or UO_1033 (O_1033,N_23239,N_23146);
xor UO_1034 (O_1034,N_23365,N_23031);
and UO_1035 (O_1035,N_24764,N_22526);
and UO_1036 (O_1036,N_23542,N_24838);
and UO_1037 (O_1037,N_24671,N_23565);
xnor UO_1038 (O_1038,N_24202,N_24731);
and UO_1039 (O_1039,N_23878,N_24178);
and UO_1040 (O_1040,N_23824,N_24047);
nor UO_1041 (O_1041,N_23076,N_24304);
and UO_1042 (O_1042,N_22566,N_24424);
and UO_1043 (O_1043,N_23600,N_24760);
nor UO_1044 (O_1044,N_22525,N_22717);
or UO_1045 (O_1045,N_24450,N_24036);
nor UO_1046 (O_1046,N_22994,N_24245);
or UO_1047 (O_1047,N_23320,N_22920);
or UO_1048 (O_1048,N_23037,N_24141);
nand UO_1049 (O_1049,N_24750,N_24987);
or UO_1050 (O_1050,N_23138,N_22520);
and UO_1051 (O_1051,N_24636,N_23924);
nand UO_1052 (O_1052,N_24043,N_24482);
nor UO_1053 (O_1053,N_23713,N_23372);
nor UO_1054 (O_1054,N_22558,N_23931);
and UO_1055 (O_1055,N_24227,N_24093);
nor UO_1056 (O_1056,N_24698,N_23955);
and UO_1057 (O_1057,N_24922,N_23277);
xnor UO_1058 (O_1058,N_23809,N_23660);
and UO_1059 (O_1059,N_24801,N_22609);
nand UO_1060 (O_1060,N_23162,N_23110);
nor UO_1061 (O_1061,N_22631,N_24990);
xnor UO_1062 (O_1062,N_24407,N_23803);
nand UO_1063 (O_1063,N_22940,N_24674);
and UO_1064 (O_1064,N_22747,N_23519);
or UO_1065 (O_1065,N_23743,N_22751);
or UO_1066 (O_1066,N_23785,N_23530);
or UO_1067 (O_1067,N_22806,N_22792);
or UO_1068 (O_1068,N_22978,N_24580);
and UO_1069 (O_1069,N_24637,N_22671);
and UO_1070 (O_1070,N_22862,N_24136);
nor UO_1071 (O_1071,N_24012,N_24096);
nand UO_1072 (O_1072,N_23492,N_22931);
xnor UO_1073 (O_1073,N_23024,N_23812);
nor UO_1074 (O_1074,N_23038,N_23720);
nand UO_1075 (O_1075,N_24718,N_24279);
and UO_1076 (O_1076,N_22876,N_24796);
and UO_1077 (O_1077,N_23190,N_23276);
nor UO_1078 (O_1078,N_23900,N_24733);
xnor UO_1079 (O_1079,N_24169,N_22814);
nor UO_1080 (O_1080,N_23478,N_23286);
or UO_1081 (O_1081,N_23023,N_23598);
and UO_1082 (O_1082,N_23015,N_23751);
nor UO_1083 (O_1083,N_23163,N_23495);
nand UO_1084 (O_1084,N_24147,N_24427);
nor UO_1085 (O_1085,N_23604,N_22752);
or UO_1086 (O_1086,N_23902,N_24952);
and UO_1087 (O_1087,N_23158,N_22659);
and UO_1088 (O_1088,N_24156,N_23694);
and UO_1089 (O_1089,N_22502,N_24607);
nand UO_1090 (O_1090,N_24426,N_24891);
nand UO_1091 (O_1091,N_24117,N_23779);
or UO_1092 (O_1092,N_24941,N_22617);
or UO_1093 (O_1093,N_24933,N_24057);
or UO_1094 (O_1094,N_24830,N_23767);
xnor UO_1095 (O_1095,N_24577,N_24585);
or UO_1096 (O_1096,N_24889,N_22939);
xnor UO_1097 (O_1097,N_22592,N_23474);
or UO_1098 (O_1098,N_22775,N_24623);
and UO_1099 (O_1099,N_24252,N_22529);
or UO_1100 (O_1100,N_24767,N_24599);
nor UO_1101 (O_1101,N_23096,N_23123);
nor UO_1102 (O_1102,N_24458,N_22581);
nand UO_1103 (O_1103,N_22762,N_23175);
or UO_1104 (O_1104,N_22503,N_22673);
xnor UO_1105 (O_1105,N_22543,N_24525);
and UO_1106 (O_1106,N_23204,N_23335);
or UO_1107 (O_1107,N_24451,N_23893);
nand UO_1108 (O_1108,N_24038,N_22841);
or UO_1109 (O_1109,N_23605,N_23896);
xor UO_1110 (O_1110,N_23128,N_22605);
or UO_1111 (O_1111,N_23349,N_22883);
and UO_1112 (O_1112,N_23202,N_23595);
and UO_1113 (O_1113,N_23333,N_23943);
nor UO_1114 (O_1114,N_22874,N_24823);
or UO_1115 (O_1115,N_24686,N_23625);
and UO_1116 (O_1116,N_24883,N_24071);
or UO_1117 (O_1117,N_24619,N_23472);
or UO_1118 (O_1118,N_24206,N_23453);
and UO_1119 (O_1119,N_24532,N_22542);
or UO_1120 (O_1120,N_24436,N_24879);
nor UO_1121 (O_1121,N_22999,N_24411);
xor UO_1122 (O_1122,N_23411,N_24884);
nand UO_1123 (O_1123,N_24814,N_22505);
nand UO_1124 (O_1124,N_22509,N_22925);
nand UO_1125 (O_1125,N_23907,N_22756);
or UO_1126 (O_1126,N_22704,N_23461);
and UO_1127 (O_1127,N_23650,N_23524);
nand UO_1128 (O_1128,N_24397,N_22765);
or UO_1129 (O_1129,N_24048,N_23626);
and UO_1130 (O_1130,N_23956,N_23609);
or UO_1131 (O_1131,N_24691,N_24374);
or UO_1132 (O_1132,N_22881,N_23420);
nand UO_1133 (O_1133,N_23688,N_22771);
nand UO_1134 (O_1134,N_23611,N_23944);
nor UO_1135 (O_1135,N_24514,N_24198);
nand UO_1136 (O_1136,N_22745,N_23842);
nor UO_1137 (O_1137,N_22635,N_22947);
nor UO_1138 (O_1138,N_23164,N_24795);
or UO_1139 (O_1139,N_24084,N_23970);
or UO_1140 (O_1140,N_24845,N_22722);
or UO_1141 (O_1141,N_24035,N_24905);
nor UO_1142 (O_1142,N_22996,N_22513);
or UO_1143 (O_1143,N_24091,N_24950);
nand UO_1144 (O_1144,N_24937,N_24916);
and UO_1145 (O_1145,N_24118,N_24368);
xor UO_1146 (O_1146,N_22594,N_23858);
nor UO_1147 (O_1147,N_24511,N_23209);
nor UO_1148 (O_1148,N_23132,N_24664);
nand UO_1149 (O_1149,N_23740,N_24289);
and UO_1150 (O_1150,N_23463,N_24085);
or UO_1151 (O_1151,N_22575,N_24029);
nand UO_1152 (O_1152,N_24349,N_24177);
nor UO_1153 (O_1153,N_22664,N_23792);
or UO_1154 (O_1154,N_23996,N_23658);
nand UO_1155 (O_1155,N_23503,N_24335);
nand UO_1156 (O_1156,N_23875,N_24052);
nor UO_1157 (O_1157,N_22836,N_22623);
or UO_1158 (O_1158,N_24127,N_24982);
nand UO_1159 (O_1159,N_24308,N_23540);
xor UO_1160 (O_1160,N_24582,N_24010);
nor UO_1161 (O_1161,N_24000,N_24195);
nand UO_1162 (O_1162,N_22648,N_22935);
or UO_1163 (O_1163,N_24121,N_23271);
nor UO_1164 (O_1164,N_23522,N_23880);
nor UO_1165 (O_1165,N_23772,N_24541);
and UO_1166 (O_1166,N_22846,N_23723);
nand UO_1167 (O_1167,N_23343,N_23055);
nand UO_1168 (O_1168,N_24358,N_23607);
nand UO_1169 (O_1169,N_24642,N_24988);
or UO_1170 (O_1170,N_23200,N_23161);
and UO_1171 (O_1171,N_24459,N_23705);
and UO_1172 (O_1172,N_24510,N_23147);
or UO_1173 (O_1173,N_23176,N_23233);
nand UO_1174 (O_1174,N_23355,N_24456);
nand UO_1175 (O_1175,N_23087,N_22871);
and UO_1176 (O_1176,N_24214,N_22962);
nand UO_1177 (O_1177,N_23217,N_24521);
nand UO_1178 (O_1178,N_23353,N_23198);
and UO_1179 (O_1179,N_24576,N_24257);
and UO_1180 (O_1180,N_23596,N_23825);
nand UO_1181 (O_1181,N_24263,N_22944);
nor UO_1182 (O_1182,N_23674,N_23314);
nor UO_1183 (O_1183,N_23012,N_22703);
nor UO_1184 (O_1184,N_22641,N_23269);
and UO_1185 (O_1185,N_23682,N_22798);
nand UO_1186 (O_1186,N_23774,N_22795);
nand UO_1187 (O_1187,N_23546,N_22710);
nor UO_1188 (O_1188,N_23932,N_24489);
nor UO_1189 (O_1189,N_23839,N_24768);
nand UO_1190 (O_1190,N_22835,N_22832);
or UO_1191 (O_1191,N_23866,N_24709);
nor UO_1192 (O_1192,N_24327,N_23734);
or UO_1193 (O_1193,N_24049,N_23775);
and UO_1194 (O_1194,N_22988,N_23936);
nand UO_1195 (O_1195,N_22891,N_23245);
and UO_1196 (O_1196,N_22697,N_23736);
xnor UO_1197 (O_1197,N_24348,N_24994);
nor UO_1198 (O_1198,N_24226,N_22977);
or UO_1199 (O_1199,N_24064,N_23831);
nand UO_1200 (O_1200,N_22555,N_22518);
nor UO_1201 (O_1201,N_24535,N_24821);
or UO_1202 (O_1202,N_23621,N_24885);
nor UO_1203 (O_1203,N_22885,N_24695);
or UO_1204 (O_1204,N_24647,N_22619);
nor UO_1205 (O_1205,N_22643,N_24344);
and UO_1206 (O_1206,N_22930,N_24608);
and UO_1207 (O_1207,N_23640,N_22863);
and UO_1208 (O_1208,N_22527,N_24840);
and UO_1209 (O_1209,N_22790,N_23584);
nor UO_1210 (O_1210,N_23140,N_22952);
or UO_1211 (O_1211,N_24130,N_24410);
nand UO_1212 (O_1212,N_24187,N_24315);
and UO_1213 (O_1213,N_24610,N_22784);
nor UO_1214 (O_1214,N_23356,N_23719);
xnor UO_1215 (O_1215,N_23092,N_23532);
or UO_1216 (O_1216,N_23045,N_24453);
nor UO_1217 (O_1217,N_22857,N_24434);
and UO_1218 (O_1218,N_24954,N_24627);
xnor UO_1219 (O_1219,N_23386,N_23085);
xnor UO_1220 (O_1220,N_23491,N_23310);
nand UO_1221 (O_1221,N_24193,N_24880);
and UO_1222 (O_1222,N_24295,N_22650);
or UO_1223 (O_1223,N_23183,N_24516);
or UO_1224 (O_1224,N_24231,N_23323);
nand UO_1225 (O_1225,N_23114,N_22615);
or UO_1226 (O_1226,N_23929,N_22622);
xnor UO_1227 (O_1227,N_24078,N_23753);
and UO_1228 (O_1228,N_23470,N_22787);
or UO_1229 (O_1229,N_24258,N_23991);
nor UO_1230 (O_1230,N_23144,N_22583);
nor UO_1231 (O_1231,N_22805,N_24264);
nand UO_1232 (O_1232,N_23230,N_23324);
and UO_1233 (O_1233,N_23874,N_24985);
nand UO_1234 (O_1234,N_22577,N_22942);
nand UO_1235 (O_1235,N_23367,N_24065);
or UO_1236 (O_1236,N_24715,N_24146);
and UO_1237 (O_1237,N_24059,N_22966);
or UO_1238 (O_1238,N_23856,N_23913);
or UO_1239 (O_1239,N_24530,N_22779);
or UO_1240 (O_1240,N_23895,N_23484);
nand UO_1241 (O_1241,N_24083,N_24578);
nor UO_1242 (O_1242,N_24945,N_24326);
or UO_1243 (O_1243,N_23490,N_24923);
and UO_1244 (O_1244,N_23203,N_24409);
nand UO_1245 (O_1245,N_24351,N_23961);
or UO_1246 (O_1246,N_23242,N_23953);
nand UO_1247 (O_1247,N_23298,N_24761);
or UO_1248 (O_1248,N_24810,N_23934);
nor UO_1249 (O_1249,N_24618,N_23795);
xnor UO_1250 (O_1250,N_23298,N_23099);
nor UO_1251 (O_1251,N_23350,N_24290);
nand UO_1252 (O_1252,N_24410,N_24637);
nor UO_1253 (O_1253,N_23041,N_23718);
and UO_1254 (O_1254,N_23306,N_24190);
or UO_1255 (O_1255,N_23658,N_24064);
and UO_1256 (O_1256,N_23478,N_22932);
or UO_1257 (O_1257,N_24906,N_22999);
nand UO_1258 (O_1258,N_24765,N_23017);
or UO_1259 (O_1259,N_24419,N_24422);
nand UO_1260 (O_1260,N_23297,N_24642);
nand UO_1261 (O_1261,N_24831,N_23895);
nor UO_1262 (O_1262,N_23038,N_23104);
nand UO_1263 (O_1263,N_24607,N_24388);
nand UO_1264 (O_1264,N_22932,N_23657);
and UO_1265 (O_1265,N_23087,N_24130);
xnor UO_1266 (O_1266,N_24264,N_23215);
and UO_1267 (O_1267,N_23349,N_24955);
xor UO_1268 (O_1268,N_24587,N_24343);
nand UO_1269 (O_1269,N_23657,N_24440);
nand UO_1270 (O_1270,N_23909,N_24139);
nand UO_1271 (O_1271,N_23214,N_23062);
and UO_1272 (O_1272,N_23915,N_23152);
or UO_1273 (O_1273,N_22827,N_24912);
nand UO_1274 (O_1274,N_23787,N_23725);
or UO_1275 (O_1275,N_24814,N_24811);
nor UO_1276 (O_1276,N_23876,N_23813);
xor UO_1277 (O_1277,N_22558,N_23169);
nand UO_1278 (O_1278,N_22560,N_23539);
nor UO_1279 (O_1279,N_24600,N_22959);
or UO_1280 (O_1280,N_22612,N_24478);
nor UO_1281 (O_1281,N_24840,N_24520);
and UO_1282 (O_1282,N_23724,N_23194);
and UO_1283 (O_1283,N_24752,N_24857);
nand UO_1284 (O_1284,N_22549,N_23245);
nor UO_1285 (O_1285,N_24175,N_23333);
nand UO_1286 (O_1286,N_24742,N_23255);
nor UO_1287 (O_1287,N_24104,N_24714);
and UO_1288 (O_1288,N_24008,N_24892);
xor UO_1289 (O_1289,N_24657,N_23423);
and UO_1290 (O_1290,N_22843,N_23773);
xor UO_1291 (O_1291,N_24277,N_24652);
or UO_1292 (O_1292,N_23479,N_22885);
and UO_1293 (O_1293,N_24097,N_23165);
and UO_1294 (O_1294,N_23349,N_22843);
xnor UO_1295 (O_1295,N_22623,N_24861);
and UO_1296 (O_1296,N_23557,N_24158);
nand UO_1297 (O_1297,N_24910,N_24814);
and UO_1298 (O_1298,N_22629,N_22579);
and UO_1299 (O_1299,N_24791,N_22933);
or UO_1300 (O_1300,N_23921,N_24173);
or UO_1301 (O_1301,N_24238,N_23878);
or UO_1302 (O_1302,N_24398,N_24835);
or UO_1303 (O_1303,N_24071,N_22814);
xnor UO_1304 (O_1304,N_23147,N_22757);
nand UO_1305 (O_1305,N_24765,N_24592);
and UO_1306 (O_1306,N_23580,N_23747);
nand UO_1307 (O_1307,N_22916,N_24375);
or UO_1308 (O_1308,N_23855,N_23592);
or UO_1309 (O_1309,N_23463,N_24738);
nand UO_1310 (O_1310,N_24761,N_24656);
nand UO_1311 (O_1311,N_24453,N_24523);
or UO_1312 (O_1312,N_24139,N_24566);
nor UO_1313 (O_1313,N_23066,N_23221);
nand UO_1314 (O_1314,N_23409,N_24683);
or UO_1315 (O_1315,N_22895,N_24460);
or UO_1316 (O_1316,N_23056,N_23892);
or UO_1317 (O_1317,N_23531,N_23124);
or UO_1318 (O_1318,N_22581,N_23962);
and UO_1319 (O_1319,N_22661,N_23306);
nand UO_1320 (O_1320,N_24580,N_24151);
nand UO_1321 (O_1321,N_24583,N_24073);
and UO_1322 (O_1322,N_22984,N_24387);
nor UO_1323 (O_1323,N_24071,N_23207);
and UO_1324 (O_1324,N_24489,N_24831);
and UO_1325 (O_1325,N_24471,N_24468);
or UO_1326 (O_1326,N_23079,N_22990);
and UO_1327 (O_1327,N_24703,N_23095);
nand UO_1328 (O_1328,N_23833,N_24309);
and UO_1329 (O_1329,N_23061,N_23327);
and UO_1330 (O_1330,N_23210,N_24827);
xor UO_1331 (O_1331,N_24740,N_24588);
nor UO_1332 (O_1332,N_24558,N_23204);
nand UO_1333 (O_1333,N_24584,N_24352);
nand UO_1334 (O_1334,N_24879,N_24503);
xor UO_1335 (O_1335,N_24231,N_23926);
and UO_1336 (O_1336,N_24439,N_23755);
and UO_1337 (O_1337,N_23237,N_23899);
xor UO_1338 (O_1338,N_23578,N_22804);
nand UO_1339 (O_1339,N_24349,N_24371);
nand UO_1340 (O_1340,N_22988,N_23129);
nor UO_1341 (O_1341,N_22626,N_22985);
and UO_1342 (O_1342,N_22764,N_24781);
or UO_1343 (O_1343,N_24670,N_23359);
and UO_1344 (O_1344,N_23846,N_23969);
or UO_1345 (O_1345,N_24252,N_23134);
or UO_1346 (O_1346,N_23746,N_24469);
or UO_1347 (O_1347,N_24707,N_24466);
or UO_1348 (O_1348,N_24837,N_23117);
nand UO_1349 (O_1349,N_24676,N_23116);
nor UO_1350 (O_1350,N_23216,N_23763);
nand UO_1351 (O_1351,N_24945,N_24045);
nor UO_1352 (O_1352,N_23675,N_24140);
and UO_1353 (O_1353,N_24128,N_22614);
or UO_1354 (O_1354,N_24772,N_24170);
nand UO_1355 (O_1355,N_23885,N_22966);
nor UO_1356 (O_1356,N_23784,N_23802);
nor UO_1357 (O_1357,N_24886,N_23682);
nor UO_1358 (O_1358,N_22593,N_22979);
nand UO_1359 (O_1359,N_24243,N_24683);
nand UO_1360 (O_1360,N_23367,N_22538);
nand UO_1361 (O_1361,N_24093,N_24129);
nand UO_1362 (O_1362,N_24192,N_23672);
nor UO_1363 (O_1363,N_23671,N_23968);
nand UO_1364 (O_1364,N_23884,N_23392);
nor UO_1365 (O_1365,N_22842,N_24696);
nor UO_1366 (O_1366,N_22621,N_23579);
nand UO_1367 (O_1367,N_24359,N_23346);
nor UO_1368 (O_1368,N_23983,N_22521);
or UO_1369 (O_1369,N_22525,N_22570);
nor UO_1370 (O_1370,N_23461,N_24186);
and UO_1371 (O_1371,N_23255,N_22624);
or UO_1372 (O_1372,N_23263,N_23716);
nor UO_1373 (O_1373,N_23982,N_24225);
nor UO_1374 (O_1374,N_23126,N_22834);
and UO_1375 (O_1375,N_23350,N_23936);
xor UO_1376 (O_1376,N_23560,N_24202);
nand UO_1377 (O_1377,N_24488,N_23706);
or UO_1378 (O_1378,N_23694,N_23991);
nand UO_1379 (O_1379,N_24057,N_24152);
nand UO_1380 (O_1380,N_23169,N_23860);
and UO_1381 (O_1381,N_23610,N_23824);
and UO_1382 (O_1382,N_24676,N_24346);
or UO_1383 (O_1383,N_22592,N_23841);
or UO_1384 (O_1384,N_24634,N_22526);
nand UO_1385 (O_1385,N_23407,N_24496);
and UO_1386 (O_1386,N_24394,N_23839);
and UO_1387 (O_1387,N_22773,N_24573);
xnor UO_1388 (O_1388,N_24142,N_24752);
nor UO_1389 (O_1389,N_24907,N_22659);
xnor UO_1390 (O_1390,N_22993,N_23376);
nor UO_1391 (O_1391,N_24680,N_23949);
nor UO_1392 (O_1392,N_23677,N_24082);
xor UO_1393 (O_1393,N_24726,N_23104);
nor UO_1394 (O_1394,N_24669,N_22551);
and UO_1395 (O_1395,N_23451,N_24533);
and UO_1396 (O_1396,N_24294,N_22594);
or UO_1397 (O_1397,N_22602,N_23193);
nor UO_1398 (O_1398,N_23409,N_24971);
or UO_1399 (O_1399,N_23145,N_22676);
or UO_1400 (O_1400,N_23011,N_24515);
and UO_1401 (O_1401,N_23637,N_22602);
nor UO_1402 (O_1402,N_22644,N_23526);
nor UO_1403 (O_1403,N_22655,N_24916);
or UO_1404 (O_1404,N_23277,N_23894);
nand UO_1405 (O_1405,N_23374,N_24767);
or UO_1406 (O_1406,N_23407,N_22927);
or UO_1407 (O_1407,N_23984,N_24142);
or UO_1408 (O_1408,N_24932,N_23205);
and UO_1409 (O_1409,N_24511,N_23455);
or UO_1410 (O_1410,N_23602,N_22536);
nand UO_1411 (O_1411,N_22957,N_23146);
nand UO_1412 (O_1412,N_22988,N_23256);
or UO_1413 (O_1413,N_24206,N_24202);
or UO_1414 (O_1414,N_23599,N_22619);
nand UO_1415 (O_1415,N_24538,N_23772);
xor UO_1416 (O_1416,N_24685,N_24706);
xnor UO_1417 (O_1417,N_22845,N_24394);
xnor UO_1418 (O_1418,N_23882,N_24368);
nand UO_1419 (O_1419,N_23814,N_23605);
or UO_1420 (O_1420,N_22660,N_23950);
nand UO_1421 (O_1421,N_22732,N_22913);
nor UO_1422 (O_1422,N_23960,N_24387);
nor UO_1423 (O_1423,N_24901,N_22931);
and UO_1424 (O_1424,N_23917,N_23995);
and UO_1425 (O_1425,N_22565,N_24669);
nor UO_1426 (O_1426,N_24664,N_22668);
xnor UO_1427 (O_1427,N_24248,N_23240);
and UO_1428 (O_1428,N_23826,N_22672);
or UO_1429 (O_1429,N_24325,N_24682);
and UO_1430 (O_1430,N_22780,N_24109);
and UO_1431 (O_1431,N_24220,N_23009);
nor UO_1432 (O_1432,N_24958,N_24896);
or UO_1433 (O_1433,N_22834,N_23293);
xnor UO_1434 (O_1434,N_23686,N_24355);
nor UO_1435 (O_1435,N_23842,N_23253);
nor UO_1436 (O_1436,N_24783,N_24371);
and UO_1437 (O_1437,N_23932,N_22766);
nand UO_1438 (O_1438,N_23565,N_23863);
nor UO_1439 (O_1439,N_22709,N_24880);
or UO_1440 (O_1440,N_24241,N_23233);
and UO_1441 (O_1441,N_22864,N_23069);
nor UO_1442 (O_1442,N_22845,N_23030);
nand UO_1443 (O_1443,N_24340,N_24831);
or UO_1444 (O_1444,N_24087,N_24366);
or UO_1445 (O_1445,N_24889,N_23261);
and UO_1446 (O_1446,N_24561,N_23644);
and UO_1447 (O_1447,N_23964,N_23003);
nand UO_1448 (O_1448,N_23431,N_23791);
nor UO_1449 (O_1449,N_23183,N_24638);
xor UO_1450 (O_1450,N_24582,N_24783);
and UO_1451 (O_1451,N_23160,N_24648);
or UO_1452 (O_1452,N_23087,N_24771);
nand UO_1453 (O_1453,N_24445,N_22605);
nor UO_1454 (O_1454,N_22590,N_23222);
nand UO_1455 (O_1455,N_23232,N_22768);
nand UO_1456 (O_1456,N_24979,N_23235);
or UO_1457 (O_1457,N_24500,N_23655);
and UO_1458 (O_1458,N_24949,N_24149);
nor UO_1459 (O_1459,N_24973,N_23646);
and UO_1460 (O_1460,N_23575,N_24542);
nor UO_1461 (O_1461,N_23034,N_23004);
nor UO_1462 (O_1462,N_24491,N_24283);
xor UO_1463 (O_1463,N_24043,N_23520);
nor UO_1464 (O_1464,N_22810,N_24804);
and UO_1465 (O_1465,N_24918,N_23694);
and UO_1466 (O_1466,N_24692,N_22583);
nand UO_1467 (O_1467,N_23511,N_22683);
xnor UO_1468 (O_1468,N_24605,N_22883);
xnor UO_1469 (O_1469,N_24749,N_24557);
xor UO_1470 (O_1470,N_22621,N_24748);
nor UO_1471 (O_1471,N_23528,N_23048);
nand UO_1472 (O_1472,N_24261,N_22841);
or UO_1473 (O_1473,N_22713,N_24466);
or UO_1474 (O_1474,N_24891,N_22855);
and UO_1475 (O_1475,N_24229,N_23999);
or UO_1476 (O_1476,N_23928,N_24596);
and UO_1477 (O_1477,N_23968,N_24243);
xnor UO_1478 (O_1478,N_24846,N_22836);
or UO_1479 (O_1479,N_24521,N_24777);
nor UO_1480 (O_1480,N_22965,N_23950);
nand UO_1481 (O_1481,N_23439,N_24255);
nor UO_1482 (O_1482,N_24477,N_24467);
or UO_1483 (O_1483,N_24640,N_23810);
or UO_1484 (O_1484,N_23279,N_24742);
nor UO_1485 (O_1485,N_22868,N_24754);
or UO_1486 (O_1486,N_23204,N_24120);
nor UO_1487 (O_1487,N_24410,N_24720);
xor UO_1488 (O_1488,N_23716,N_23137);
nor UO_1489 (O_1489,N_24111,N_23262);
or UO_1490 (O_1490,N_23520,N_23438);
nor UO_1491 (O_1491,N_23471,N_22931);
nor UO_1492 (O_1492,N_23494,N_23106);
nand UO_1493 (O_1493,N_23997,N_23827);
nor UO_1494 (O_1494,N_23640,N_24517);
xor UO_1495 (O_1495,N_24308,N_22633);
nor UO_1496 (O_1496,N_24758,N_22706);
or UO_1497 (O_1497,N_22517,N_24297);
nor UO_1498 (O_1498,N_24807,N_24792);
and UO_1499 (O_1499,N_24861,N_24470);
nand UO_1500 (O_1500,N_23170,N_24876);
nor UO_1501 (O_1501,N_24843,N_23423);
and UO_1502 (O_1502,N_23957,N_24924);
nand UO_1503 (O_1503,N_24051,N_23292);
xor UO_1504 (O_1504,N_23754,N_23182);
nor UO_1505 (O_1505,N_24578,N_24701);
and UO_1506 (O_1506,N_24394,N_23710);
or UO_1507 (O_1507,N_23469,N_24422);
and UO_1508 (O_1508,N_24724,N_24265);
nand UO_1509 (O_1509,N_23263,N_24676);
and UO_1510 (O_1510,N_24510,N_22866);
or UO_1511 (O_1511,N_23003,N_23260);
or UO_1512 (O_1512,N_24207,N_23303);
xnor UO_1513 (O_1513,N_24445,N_23466);
and UO_1514 (O_1514,N_24666,N_24573);
and UO_1515 (O_1515,N_24065,N_22570);
nand UO_1516 (O_1516,N_23616,N_24059);
nand UO_1517 (O_1517,N_24060,N_23379);
nor UO_1518 (O_1518,N_23581,N_23886);
nor UO_1519 (O_1519,N_24800,N_22812);
nor UO_1520 (O_1520,N_22659,N_24633);
xor UO_1521 (O_1521,N_24175,N_23750);
and UO_1522 (O_1522,N_22789,N_24195);
nor UO_1523 (O_1523,N_23969,N_22818);
or UO_1524 (O_1524,N_22504,N_24169);
nor UO_1525 (O_1525,N_22842,N_23375);
nor UO_1526 (O_1526,N_22863,N_24300);
and UO_1527 (O_1527,N_24408,N_22957);
xor UO_1528 (O_1528,N_24939,N_23734);
and UO_1529 (O_1529,N_23637,N_23497);
nand UO_1530 (O_1530,N_24541,N_24898);
or UO_1531 (O_1531,N_24901,N_23257);
nand UO_1532 (O_1532,N_24821,N_24178);
nand UO_1533 (O_1533,N_24441,N_22720);
nor UO_1534 (O_1534,N_24951,N_23619);
or UO_1535 (O_1535,N_23396,N_24883);
nand UO_1536 (O_1536,N_24251,N_23966);
and UO_1537 (O_1537,N_24899,N_24430);
and UO_1538 (O_1538,N_22669,N_24951);
nor UO_1539 (O_1539,N_22631,N_23064);
and UO_1540 (O_1540,N_23251,N_23263);
nand UO_1541 (O_1541,N_24477,N_22965);
or UO_1542 (O_1542,N_23274,N_23072);
nand UO_1543 (O_1543,N_22887,N_24143);
nand UO_1544 (O_1544,N_24506,N_23869);
nand UO_1545 (O_1545,N_23630,N_23330);
and UO_1546 (O_1546,N_24790,N_22618);
and UO_1547 (O_1547,N_24727,N_23572);
nor UO_1548 (O_1548,N_23340,N_24158);
xor UO_1549 (O_1549,N_22629,N_24593);
or UO_1550 (O_1550,N_23655,N_22823);
or UO_1551 (O_1551,N_24044,N_22666);
or UO_1552 (O_1552,N_24018,N_22846);
nor UO_1553 (O_1553,N_23734,N_22994);
and UO_1554 (O_1554,N_24527,N_24239);
and UO_1555 (O_1555,N_24104,N_23053);
nor UO_1556 (O_1556,N_24849,N_23415);
and UO_1557 (O_1557,N_23719,N_23949);
or UO_1558 (O_1558,N_23039,N_24556);
nand UO_1559 (O_1559,N_24436,N_24071);
nor UO_1560 (O_1560,N_24169,N_22766);
and UO_1561 (O_1561,N_24649,N_23221);
or UO_1562 (O_1562,N_23972,N_22738);
nand UO_1563 (O_1563,N_24325,N_22999);
and UO_1564 (O_1564,N_22626,N_22953);
xor UO_1565 (O_1565,N_24365,N_23258);
and UO_1566 (O_1566,N_24147,N_23468);
nor UO_1567 (O_1567,N_23672,N_24046);
xor UO_1568 (O_1568,N_23247,N_24476);
nand UO_1569 (O_1569,N_23724,N_24014);
or UO_1570 (O_1570,N_23375,N_24137);
or UO_1571 (O_1571,N_23396,N_23813);
nor UO_1572 (O_1572,N_22966,N_22592);
nand UO_1573 (O_1573,N_24164,N_24086);
nor UO_1574 (O_1574,N_23058,N_24086);
and UO_1575 (O_1575,N_24105,N_23650);
or UO_1576 (O_1576,N_23575,N_24569);
nor UO_1577 (O_1577,N_22975,N_22789);
or UO_1578 (O_1578,N_22566,N_22772);
nor UO_1579 (O_1579,N_24697,N_23621);
nor UO_1580 (O_1580,N_23799,N_23909);
or UO_1581 (O_1581,N_23335,N_23180);
nand UO_1582 (O_1582,N_22603,N_23201);
nor UO_1583 (O_1583,N_23781,N_24889);
and UO_1584 (O_1584,N_23468,N_24272);
nand UO_1585 (O_1585,N_23147,N_24451);
nor UO_1586 (O_1586,N_24540,N_23713);
nand UO_1587 (O_1587,N_23154,N_23512);
or UO_1588 (O_1588,N_23511,N_23195);
and UO_1589 (O_1589,N_22817,N_23743);
or UO_1590 (O_1590,N_23169,N_23901);
nor UO_1591 (O_1591,N_24154,N_22725);
nand UO_1592 (O_1592,N_22992,N_23952);
or UO_1593 (O_1593,N_23684,N_22601);
nand UO_1594 (O_1594,N_22513,N_24482);
nand UO_1595 (O_1595,N_22850,N_24733);
nor UO_1596 (O_1596,N_24490,N_24169);
xnor UO_1597 (O_1597,N_24104,N_23029);
and UO_1598 (O_1598,N_22968,N_22684);
and UO_1599 (O_1599,N_24541,N_24363);
and UO_1600 (O_1600,N_22884,N_23424);
xor UO_1601 (O_1601,N_22990,N_24533);
or UO_1602 (O_1602,N_22744,N_23247);
or UO_1603 (O_1603,N_24079,N_22997);
xor UO_1604 (O_1604,N_23221,N_23517);
and UO_1605 (O_1605,N_24004,N_23254);
xnor UO_1606 (O_1606,N_22508,N_24042);
nand UO_1607 (O_1607,N_24535,N_24737);
nor UO_1608 (O_1608,N_23753,N_24094);
and UO_1609 (O_1609,N_22810,N_23119);
and UO_1610 (O_1610,N_22886,N_23042);
nand UO_1611 (O_1611,N_24009,N_23645);
nor UO_1612 (O_1612,N_24265,N_23546);
xor UO_1613 (O_1613,N_23915,N_23044);
and UO_1614 (O_1614,N_24992,N_22662);
nand UO_1615 (O_1615,N_22721,N_24806);
and UO_1616 (O_1616,N_22814,N_23541);
and UO_1617 (O_1617,N_23467,N_23271);
nor UO_1618 (O_1618,N_22529,N_22594);
nand UO_1619 (O_1619,N_22988,N_24561);
or UO_1620 (O_1620,N_23556,N_23820);
nor UO_1621 (O_1621,N_24030,N_24513);
nand UO_1622 (O_1622,N_24733,N_23751);
or UO_1623 (O_1623,N_24519,N_23252);
or UO_1624 (O_1624,N_22625,N_22989);
xnor UO_1625 (O_1625,N_23456,N_23182);
nand UO_1626 (O_1626,N_24163,N_24068);
and UO_1627 (O_1627,N_24928,N_22787);
nand UO_1628 (O_1628,N_22911,N_23571);
or UO_1629 (O_1629,N_23394,N_23642);
xnor UO_1630 (O_1630,N_23826,N_24847);
or UO_1631 (O_1631,N_23951,N_24239);
nand UO_1632 (O_1632,N_24861,N_23291);
nand UO_1633 (O_1633,N_24056,N_24897);
xor UO_1634 (O_1634,N_23712,N_24570);
nor UO_1635 (O_1635,N_24473,N_24567);
nand UO_1636 (O_1636,N_22743,N_24953);
xnor UO_1637 (O_1637,N_22663,N_23940);
nand UO_1638 (O_1638,N_22905,N_23404);
or UO_1639 (O_1639,N_24157,N_23127);
nand UO_1640 (O_1640,N_24092,N_23221);
nand UO_1641 (O_1641,N_23780,N_24904);
and UO_1642 (O_1642,N_23322,N_24079);
nor UO_1643 (O_1643,N_24608,N_23883);
nand UO_1644 (O_1644,N_23364,N_22729);
nor UO_1645 (O_1645,N_23218,N_23213);
nor UO_1646 (O_1646,N_23483,N_22657);
nor UO_1647 (O_1647,N_23206,N_24074);
nand UO_1648 (O_1648,N_24458,N_23387);
and UO_1649 (O_1649,N_24107,N_24853);
nand UO_1650 (O_1650,N_22809,N_24988);
and UO_1651 (O_1651,N_22611,N_23710);
nor UO_1652 (O_1652,N_24659,N_24172);
or UO_1653 (O_1653,N_24742,N_24029);
nor UO_1654 (O_1654,N_23674,N_22625);
nor UO_1655 (O_1655,N_24814,N_23608);
nand UO_1656 (O_1656,N_24410,N_23265);
xor UO_1657 (O_1657,N_22994,N_23604);
and UO_1658 (O_1658,N_22743,N_23808);
xor UO_1659 (O_1659,N_24242,N_23927);
or UO_1660 (O_1660,N_23965,N_23890);
nand UO_1661 (O_1661,N_23194,N_23390);
nand UO_1662 (O_1662,N_24044,N_22851);
or UO_1663 (O_1663,N_22890,N_22636);
or UO_1664 (O_1664,N_23225,N_23658);
or UO_1665 (O_1665,N_23731,N_23348);
and UO_1666 (O_1666,N_23978,N_23328);
or UO_1667 (O_1667,N_23874,N_22616);
xnor UO_1668 (O_1668,N_23284,N_24448);
and UO_1669 (O_1669,N_24089,N_24157);
nand UO_1670 (O_1670,N_23657,N_24014);
nand UO_1671 (O_1671,N_23850,N_23877);
nor UO_1672 (O_1672,N_22668,N_24297);
or UO_1673 (O_1673,N_22992,N_24917);
nand UO_1674 (O_1674,N_23543,N_23888);
nand UO_1675 (O_1675,N_23558,N_22650);
and UO_1676 (O_1676,N_23327,N_23562);
and UO_1677 (O_1677,N_23501,N_24157);
or UO_1678 (O_1678,N_22680,N_24604);
or UO_1679 (O_1679,N_22540,N_24441);
nor UO_1680 (O_1680,N_23095,N_23056);
xor UO_1681 (O_1681,N_24197,N_23857);
nand UO_1682 (O_1682,N_23178,N_24392);
xnor UO_1683 (O_1683,N_23230,N_22553);
nor UO_1684 (O_1684,N_24090,N_22643);
and UO_1685 (O_1685,N_23464,N_23084);
or UO_1686 (O_1686,N_23972,N_22828);
and UO_1687 (O_1687,N_23801,N_23711);
nand UO_1688 (O_1688,N_23657,N_23476);
nor UO_1689 (O_1689,N_23314,N_23912);
and UO_1690 (O_1690,N_24966,N_24243);
and UO_1691 (O_1691,N_24327,N_22686);
or UO_1692 (O_1692,N_23876,N_24665);
and UO_1693 (O_1693,N_22670,N_24022);
nor UO_1694 (O_1694,N_24165,N_24511);
or UO_1695 (O_1695,N_23760,N_23570);
and UO_1696 (O_1696,N_24601,N_22789);
or UO_1697 (O_1697,N_23737,N_24236);
or UO_1698 (O_1698,N_22963,N_24945);
nand UO_1699 (O_1699,N_24154,N_24985);
nand UO_1700 (O_1700,N_23988,N_24133);
or UO_1701 (O_1701,N_24976,N_24076);
or UO_1702 (O_1702,N_24893,N_24724);
or UO_1703 (O_1703,N_22760,N_23309);
and UO_1704 (O_1704,N_24261,N_24000);
nor UO_1705 (O_1705,N_24901,N_24679);
or UO_1706 (O_1706,N_24876,N_24890);
nand UO_1707 (O_1707,N_24355,N_23269);
or UO_1708 (O_1708,N_23817,N_23636);
and UO_1709 (O_1709,N_23347,N_24022);
nand UO_1710 (O_1710,N_22541,N_24390);
nor UO_1711 (O_1711,N_22540,N_23760);
or UO_1712 (O_1712,N_23393,N_24548);
or UO_1713 (O_1713,N_22528,N_24213);
or UO_1714 (O_1714,N_24126,N_23279);
nand UO_1715 (O_1715,N_23687,N_24334);
nand UO_1716 (O_1716,N_23504,N_24924);
or UO_1717 (O_1717,N_24093,N_23786);
nor UO_1718 (O_1718,N_23953,N_24090);
and UO_1719 (O_1719,N_24003,N_23528);
nor UO_1720 (O_1720,N_24578,N_22796);
xor UO_1721 (O_1721,N_22633,N_24411);
xor UO_1722 (O_1722,N_23066,N_23921);
nand UO_1723 (O_1723,N_23581,N_24635);
and UO_1724 (O_1724,N_22651,N_22684);
or UO_1725 (O_1725,N_22725,N_23404);
nor UO_1726 (O_1726,N_22701,N_22569);
xnor UO_1727 (O_1727,N_23232,N_24235);
nor UO_1728 (O_1728,N_24219,N_23653);
nand UO_1729 (O_1729,N_24287,N_24081);
xnor UO_1730 (O_1730,N_23756,N_22696);
nand UO_1731 (O_1731,N_23624,N_24868);
nor UO_1732 (O_1732,N_23431,N_24346);
nor UO_1733 (O_1733,N_24989,N_23339);
and UO_1734 (O_1734,N_24966,N_24704);
or UO_1735 (O_1735,N_24060,N_23289);
nor UO_1736 (O_1736,N_22541,N_23412);
nand UO_1737 (O_1737,N_24462,N_23049);
or UO_1738 (O_1738,N_24051,N_22773);
or UO_1739 (O_1739,N_24770,N_23234);
nand UO_1740 (O_1740,N_23914,N_23445);
and UO_1741 (O_1741,N_22839,N_23065);
or UO_1742 (O_1742,N_23630,N_23081);
and UO_1743 (O_1743,N_23974,N_23672);
and UO_1744 (O_1744,N_24047,N_23449);
nand UO_1745 (O_1745,N_22521,N_23863);
or UO_1746 (O_1746,N_23582,N_22895);
or UO_1747 (O_1747,N_23621,N_24441);
and UO_1748 (O_1748,N_23816,N_24096);
xor UO_1749 (O_1749,N_23053,N_24647);
and UO_1750 (O_1750,N_24772,N_23932);
xnor UO_1751 (O_1751,N_23653,N_23862);
nor UO_1752 (O_1752,N_24333,N_23853);
nand UO_1753 (O_1753,N_24999,N_24976);
and UO_1754 (O_1754,N_24595,N_23020);
nand UO_1755 (O_1755,N_22717,N_23669);
and UO_1756 (O_1756,N_22772,N_24128);
and UO_1757 (O_1757,N_22740,N_24627);
nand UO_1758 (O_1758,N_22799,N_22954);
and UO_1759 (O_1759,N_23619,N_24763);
nand UO_1760 (O_1760,N_23399,N_24676);
or UO_1761 (O_1761,N_22804,N_22555);
or UO_1762 (O_1762,N_24109,N_22929);
or UO_1763 (O_1763,N_23773,N_23042);
and UO_1764 (O_1764,N_22654,N_22644);
nor UO_1765 (O_1765,N_24529,N_24421);
or UO_1766 (O_1766,N_24908,N_23709);
or UO_1767 (O_1767,N_22836,N_24747);
nand UO_1768 (O_1768,N_22783,N_24777);
and UO_1769 (O_1769,N_24059,N_22782);
nor UO_1770 (O_1770,N_24914,N_23091);
and UO_1771 (O_1771,N_23199,N_24414);
or UO_1772 (O_1772,N_23741,N_24876);
and UO_1773 (O_1773,N_24380,N_23745);
and UO_1774 (O_1774,N_23534,N_22608);
nor UO_1775 (O_1775,N_22718,N_24312);
or UO_1776 (O_1776,N_23042,N_22957);
or UO_1777 (O_1777,N_24825,N_24363);
nand UO_1778 (O_1778,N_23551,N_23359);
nor UO_1779 (O_1779,N_22750,N_24098);
and UO_1780 (O_1780,N_24423,N_23318);
or UO_1781 (O_1781,N_23894,N_24073);
nor UO_1782 (O_1782,N_24009,N_22760);
nor UO_1783 (O_1783,N_23788,N_24882);
nand UO_1784 (O_1784,N_23813,N_24841);
nor UO_1785 (O_1785,N_22917,N_24200);
or UO_1786 (O_1786,N_23359,N_23337);
or UO_1787 (O_1787,N_23021,N_24090);
and UO_1788 (O_1788,N_23319,N_24919);
nor UO_1789 (O_1789,N_23173,N_24787);
or UO_1790 (O_1790,N_22758,N_24583);
and UO_1791 (O_1791,N_22887,N_23168);
nand UO_1792 (O_1792,N_23293,N_24041);
nor UO_1793 (O_1793,N_23129,N_23023);
and UO_1794 (O_1794,N_22807,N_23393);
xnor UO_1795 (O_1795,N_24016,N_22556);
nand UO_1796 (O_1796,N_24397,N_23470);
or UO_1797 (O_1797,N_24959,N_22887);
nand UO_1798 (O_1798,N_22883,N_22541);
and UO_1799 (O_1799,N_24650,N_24745);
or UO_1800 (O_1800,N_24011,N_23209);
nand UO_1801 (O_1801,N_24965,N_24639);
xnor UO_1802 (O_1802,N_24887,N_23931);
xor UO_1803 (O_1803,N_22678,N_23036);
nor UO_1804 (O_1804,N_23026,N_24242);
nand UO_1805 (O_1805,N_23103,N_23222);
nand UO_1806 (O_1806,N_23424,N_23313);
nand UO_1807 (O_1807,N_22596,N_24965);
xor UO_1808 (O_1808,N_23483,N_22779);
or UO_1809 (O_1809,N_23072,N_24225);
or UO_1810 (O_1810,N_23989,N_22529);
nor UO_1811 (O_1811,N_23070,N_24989);
nand UO_1812 (O_1812,N_24835,N_24739);
nand UO_1813 (O_1813,N_23415,N_22520);
and UO_1814 (O_1814,N_24786,N_23932);
nand UO_1815 (O_1815,N_23047,N_24919);
or UO_1816 (O_1816,N_23554,N_24430);
or UO_1817 (O_1817,N_23377,N_24519);
nor UO_1818 (O_1818,N_23037,N_23495);
nor UO_1819 (O_1819,N_23166,N_23510);
nor UO_1820 (O_1820,N_23105,N_22842);
nand UO_1821 (O_1821,N_24809,N_23770);
nand UO_1822 (O_1822,N_22601,N_23607);
nor UO_1823 (O_1823,N_22561,N_23553);
nor UO_1824 (O_1824,N_24255,N_24432);
nor UO_1825 (O_1825,N_24548,N_24737);
nor UO_1826 (O_1826,N_22510,N_23516);
and UO_1827 (O_1827,N_24507,N_23453);
and UO_1828 (O_1828,N_24985,N_23411);
nor UO_1829 (O_1829,N_24410,N_23219);
nor UO_1830 (O_1830,N_22634,N_23711);
xnor UO_1831 (O_1831,N_24362,N_23222);
or UO_1832 (O_1832,N_22713,N_23936);
and UO_1833 (O_1833,N_23415,N_24054);
and UO_1834 (O_1834,N_24950,N_22736);
nor UO_1835 (O_1835,N_23676,N_24986);
or UO_1836 (O_1836,N_23398,N_22879);
xnor UO_1837 (O_1837,N_24465,N_24129);
nand UO_1838 (O_1838,N_23079,N_24730);
or UO_1839 (O_1839,N_23353,N_24312);
nand UO_1840 (O_1840,N_24938,N_23987);
nor UO_1841 (O_1841,N_24267,N_23972);
or UO_1842 (O_1842,N_24107,N_23886);
nor UO_1843 (O_1843,N_22594,N_24794);
or UO_1844 (O_1844,N_22538,N_22565);
or UO_1845 (O_1845,N_23862,N_22692);
nor UO_1846 (O_1846,N_23933,N_24224);
xnor UO_1847 (O_1847,N_23712,N_22575);
nand UO_1848 (O_1848,N_24141,N_24448);
nand UO_1849 (O_1849,N_23623,N_23160);
xnor UO_1850 (O_1850,N_24510,N_23787);
or UO_1851 (O_1851,N_23801,N_23162);
xor UO_1852 (O_1852,N_24380,N_24796);
or UO_1853 (O_1853,N_24490,N_24377);
nor UO_1854 (O_1854,N_22701,N_22553);
nor UO_1855 (O_1855,N_23542,N_23304);
nand UO_1856 (O_1856,N_22753,N_23483);
or UO_1857 (O_1857,N_24040,N_23723);
xnor UO_1858 (O_1858,N_24827,N_24070);
and UO_1859 (O_1859,N_23104,N_23288);
and UO_1860 (O_1860,N_22520,N_24148);
nand UO_1861 (O_1861,N_23235,N_24472);
and UO_1862 (O_1862,N_22759,N_24509);
and UO_1863 (O_1863,N_23443,N_23988);
and UO_1864 (O_1864,N_22739,N_23128);
xor UO_1865 (O_1865,N_24259,N_23813);
or UO_1866 (O_1866,N_22751,N_23953);
xnor UO_1867 (O_1867,N_23388,N_24598);
nor UO_1868 (O_1868,N_23689,N_23497);
and UO_1869 (O_1869,N_23021,N_24808);
and UO_1870 (O_1870,N_23319,N_22922);
nor UO_1871 (O_1871,N_23160,N_24089);
or UO_1872 (O_1872,N_22724,N_23939);
and UO_1873 (O_1873,N_23570,N_23608);
xnor UO_1874 (O_1874,N_24539,N_23234);
and UO_1875 (O_1875,N_23659,N_23130);
or UO_1876 (O_1876,N_24301,N_24778);
nand UO_1877 (O_1877,N_24722,N_23088);
nand UO_1878 (O_1878,N_23439,N_23929);
or UO_1879 (O_1879,N_24833,N_24538);
or UO_1880 (O_1880,N_22510,N_24157);
nor UO_1881 (O_1881,N_22747,N_23472);
and UO_1882 (O_1882,N_24777,N_23158);
or UO_1883 (O_1883,N_24891,N_24797);
or UO_1884 (O_1884,N_23724,N_22806);
or UO_1885 (O_1885,N_23117,N_24585);
nor UO_1886 (O_1886,N_23519,N_24564);
and UO_1887 (O_1887,N_23510,N_24525);
nand UO_1888 (O_1888,N_23344,N_23568);
nor UO_1889 (O_1889,N_24606,N_23009);
and UO_1890 (O_1890,N_24044,N_22899);
and UO_1891 (O_1891,N_23939,N_23515);
nand UO_1892 (O_1892,N_23265,N_22928);
nand UO_1893 (O_1893,N_23537,N_24256);
or UO_1894 (O_1894,N_24234,N_23902);
and UO_1895 (O_1895,N_23124,N_23437);
nor UO_1896 (O_1896,N_23284,N_24934);
nand UO_1897 (O_1897,N_24043,N_24670);
or UO_1898 (O_1898,N_22638,N_23577);
xor UO_1899 (O_1899,N_24565,N_22644);
and UO_1900 (O_1900,N_24723,N_23861);
or UO_1901 (O_1901,N_24549,N_23286);
and UO_1902 (O_1902,N_24516,N_22514);
nand UO_1903 (O_1903,N_24018,N_24389);
xor UO_1904 (O_1904,N_23909,N_24431);
nand UO_1905 (O_1905,N_23828,N_23071);
xnor UO_1906 (O_1906,N_24746,N_22690);
or UO_1907 (O_1907,N_24861,N_23044);
and UO_1908 (O_1908,N_23613,N_22835);
nand UO_1909 (O_1909,N_24718,N_23994);
and UO_1910 (O_1910,N_23436,N_24981);
or UO_1911 (O_1911,N_23821,N_24289);
xor UO_1912 (O_1912,N_24766,N_22721);
nor UO_1913 (O_1913,N_24218,N_24155);
xor UO_1914 (O_1914,N_24324,N_22595);
or UO_1915 (O_1915,N_22700,N_24241);
nor UO_1916 (O_1916,N_23339,N_23551);
nand UO_1917 (O_1917,N_24288,N_22874);
nand UO_1918 (O_1918,N_23360,N_24625);
or UO_1919 (O_1919,N_23343,N_24863);
or UO_1920 (O_1920,N_24918,N_24034);
xnor UO_1921 (O_1921,N_24703,N_22851);
nor UO_1922 (O_1922,N_24009,N_23657);
xnor UO_1923 (O_1923,N_24131,N_23937);
nor UO_1924 (O_1924,N_24022,N_24451);
nor UO_1925 (O_1925,N_23042,N_22822);
nand UO_1926 (O_1926,N_24864,N_23427);
nor UO_1927 (O_1927,N_23261,N_24380);
and UO_1928 (O_1928,N_22549,N_22534);
and UO_1929 (O_1929,N_24684,N_24437);
nand UO_1930 (O_1930,N_22663,N_24608);
nor UO_1931 (O_1931,N_23675,N_24459);
nand UO_1932 (O_1932,N_24583,N_23354);
nor UO_1933 (O_1933,N_23346,N_24210);
or UO_1934 (O_1934,N_24270,N_22689);
or UO_1935 (O_1935,N_22812,N_23974);
or UO_1936 (O_1936,N_22539,N_23065);
nand UO_1937 (O_1937,N_23396,N_23568);
and UO_1938 (O_1938,N_23042,N_24668);
nor UO_1939 (O_1939,N_23008,N_22788);
nand UO_1940 (O_1940,N_24392,N_22966);
nand UO_1941 (O_1941,N_23215,N_23575);
nand UO_1942 (O_1942,N_24927,N_23216);
and UO_1943 (O_1943,N_23342,N_24450);
and UO_1944 (O_1944,N_23283,N_24938);
nor UO_1945 (O_1945,N_23791,N_23006);
nor UO_1946 (O_1946,N_24726,N_23942);
and UO_1947 (O_1947,N_23353,N_23552);
nor UO_1948 (O_1948,N_24890,N_22758);
and UO_1949 (O_1949,N_24653,N_24708);
and UO_1950 (O_1950,N_23364,N_22734);
or UO_1951 (O_1951,N_24296,N_23158);
nand UO_1952 (O_1952,N_24527,N_22905);
nor UO_1953 (O_1953,N_24297,N_24368);
xor UO_1954 (O_1954,N_24430,N_23143);
nand UO_1955 (O_1955,N_23220,N_23873);
nand UO_1956 (O_1956,N_22776,N_23522);
and UO_1957 (O_1957,N_23137,N_22929);
nor UO_1958 (O_1958,N_24511,N_23797);
nand UO_1959 (O_1959,N_22914,N_23574);
nor UO_1960 (O_1960,N_23632,N_22560);
nor UO_1961 (O_1961,N_24271,N_23437);
and UO_1962 (O_1962,N_24609,N_22812);
or UO_1963 (O_1963,N_24053,N_23267);
and UO_1964 (O_1964,N_23302,N_23024);
and UO_1965 (O_1965,N_23474,N_24867);
nor UO_1966 (O_1966,N_22711,N_23980);
or UO_1967 (O_1967,N_24436,N_23895);
nor UO_1968 (O_1968,N_23200,N_24648);
and UO_1969 (O_1969,N_23219,N_24296);
and UO_1970 (O_1970,N_23779,N_24078);
xnor UO_1971 (O_1971,N_23755,N_23806);
nor UO_1972 (O_1972,N_23076,N_24184);
or UO_1973 (O_1973,N_24927,N_23042);
and UO_1974 (O_1974,N_24387,N_23384);
or UO_1975 (O_1975,N_22699,N_24415);
nor UO_1976 (O_1976,N_23776,N_24672);
xor UO_1977 (O_1977,N_24814,N_24265);
nor UO_1978 (O_1978,N_23447,N_24884);
nor UO_1979 (O_1979,N_23025,N_24486);
nor UO_1980 (O_1980,N_23505,N_24899);
nand UO_1981 (O_1981,N_24960,N_23780);
nand UO_1982 (O_1982,N_22791,N_23939);
or UO_1983 (O_1983,N_23491,N_23565);
or UO_1984 (O_1984,N_24469,N_24261);
and UO_1985 (O_1985,N_24237,N_24876);
nor UO_1986 (O_1986,N_23272,N_23085);
nor UO_1987 (O_1987,N_24323,N_23240);
nor UO_1988 (O_1988,N_24640,N_24313);
nand UO_1989 (O_1989,N_23771,N_23471);
and UO_1990 (O_1990,N_24920,N_23880);
or UO_1991 (O_1991,N_23335,N_23155);
and UO_1992 (O_1992,N_23579,N_22843);
and UO_1993 (O_1993,N_24778,N_23394);
nor UO_1994 (O_1994,N_24046,N_23204);
or UO_1995 (O_1995,N_23498,N_23176);
nand UO_1996 (O_1996,N_24297,N_22914);
nand UO_1997 (O_1997,N_22860,N_23267);
nand UO_1998 (O_1998,N_23494,N_24463);
nor UO_1999 (O_1999,N_23575,N_22702);
or UO_2000 (O_2000,N_23420,N_24832);
or UO_2001 (O_2001,N_23070,N_23157);
and UO_2002 (O_2002,N_24586,N_24406);
or UO_2003 (O_2003,N_23001,N_24840);
and UO_2004 (O_2004,N_23134,N_23891);
nor UO_2005 (O_2005,N_23150,N_23328);
nor UO_2006 (O_2006,N_22718,N_24845);
and UO_2007 (O_2007,N_24948,N_23713);
and UO_2008 (O_2008,N_24808,N_23053);
and UO_2009 (O_2009,N_24083,N_24825);
nor UO_2010 (O_2010,N_23326,N_23440);
nand UO_2011 (O_2011,N_24796,N_24304);
and UO_2012 (O_2012,N_23328,N_24451);
nand UO_2013 (O_2013,N_23890,N_23307);
nand UO_2014 (O_2014,N_23111,N_22612);
and UO_2015 (O_2015,N_23495,N_24801);
and UO_2016 (O_2016,N_22845,N_24091);
xor UO_2017 (O_2017,N_23391,N_22599);
or UO_2018 (O_2018,N_23322,N_23460);
nor UO_2019 (O_2019,N_24113,N_23872);
and UO_2020 (O_2020,N_23242,N_24909);
and UO_2021 (O_2021,N_23639,N_22513);
nor UO_2022 (O_2022,N_23514,N_23986);
and UO_2023 (O_2023,N_23393,N_23206);
or UO_2024 (O_2024,N_22798,N_23639);
nor UO_2025 (O_2025,N_24268,N_23595);
nand UO_2026 (O_2026,N_23002,N_22975);
nand UO_2027 (O_2027,N_24916,N_24929);
nand UO_2028 (O_2028,N_24317,N_24646);
nor UO_2029 (O_2029,N_24908,N_23401);
nor UO_2030 (O_2030,N_24561,N_22814);
nor UO_2031 (O_2031,N_22884,N_23500);
or UO_2032 (O_2032,N_24114,N_24775);
and UO_2033 (O_2033,N_23941,N_23020);
or UO_2034 (O_2034,N_23929,N_24610);
nor UO_2035 (O_2035,N_24135,N_24116);
nand UO_2036 (O_2036,N_22978,N_23348);
nand UO_2037 (O_2037,N_23993,N_22804);
nand UO_2038 (O_2038,N_23671,N_23918);
xnor UO_2039 (O_2039,N_24715,N_22528);
nand UO_2040 (O_2040,N_24701,N_24649);
and UO_2041 (O_2041,N_23274,N_24924);
nand UO_2042 (O_2042,N_24793,N_24663);
nor UO_2043 (O_2043,N_23858,N_23627);
nor UO_2044 (O_2044,N_22974,N_24367);
nand UO_2045 (O_2045,N_22685,N_23110);
nand UO_2046 (O_2046,N_23892,N_23533);
nor UO_2047 (O_2047,N_24059,N_22558);
nand UO_2048 (O_2048,N_22726,N_23385);
nand UO_2049 (O_2049,N_24314,N_22619);
or UO_2050 (O_2050,N_23993,N_24135);
xor UO_2051 (O_2051,N_24118,N_23850);
nor UO_2052 (O_2052,N_23060,N_22665);
or UO_2053 (O_2053,N_22864,N_24703);
nand UO_2054 (O_2054,N_24881,N_24743);
or UO_2055 (O_2055,N_24361,N_22534);
and UO_2056 (O_2056,N_23746,N_24967);
nand UO_2057 (O_2057,N_23955,N_22943);
xor UO_2058 (O_2058,N_23578,N_24333);
nand UO_2059 (O_2059,N_23563,N_24366);
nor UO_2060 (O_2060,N_23027,N_24631);
or UO_2061 (O_2061,N_24683,N_24012);
nand UO_2062 (O_2062,N_22868,N_23616);
and UO_2063 (O_2063,N_23771,N_23300);
or UO_2064 (O_2064,N_23396,N_24979);
nand UO_2065 (O_2065,N_24125,N_24284);
xnor UO_2066 (O_2066,N_24191,N_24226);
and UO_2067 (O_2067,N_23945,N_23347);
or UO_2068 (O_2068,N_24649,N_24571);
nor UO_2069 (O_2069,N_23057,N_23281);
nand UO_2070 (O_2070,N_24819,N_24795);
nand UO_2071 (O_2071,N_23038,N_23320);
or UO_2072 (O_2072,N_23896,N_24006);
nand UO_2073 (O_2073,N_22731,N_24322);
nor UO_2074 (O_2074,N_24016,N_23330);
nor UO_2075 (O_2075,N_22659,N_22665);
nor UO_2076 (O_2076,N_23572,N_22817);
and UO_2077 (O_2077,N_22791,N_24917);
nor UO_2078 (O_2078,N_22915,N_23041);
nand UO_2079 (O_2079,N_24809,N_24153);
xor UO_2080 (O_2080,N_23215,N_23467);
nor UO_2081 (O_2081,N_24520,N_22602);
nor UO_2082 (O_2082,N_24704,N_24174);
xnor UO_2083 (O_2083,N_24915,N_24454);
nand UO_2084 (O_2084,N_23626,N_24329);
nor UO_2085 (O_2085,N_22876,N_24937);
and UO_2086 (O_2086,N_23184,N_24762);
nor UO_2087 (O_2087,N_24698,N_24054);
and UO_2088 (O_2088,N_22623,N_23253);
or UO_2089 (O_2089,N_23309,N_24720);
nand UO_2090 (O_2090,N_22871,N_24844);
and UO_2091 (O_2091,N_22652,N_22910);
nand UO_2092 (O_2092,N_22539,N_23549);
nand UO_2093 (O_2093,N_23009,N_24391);
or UO_2094 (O_2094,N_24038,N_22600);
nor UO_2095 (O_2095,N_23171,N_23457);
nor UO_2096 (O_2096,N_22506,N_23662);
and UO_2097 (O_2097,N_24775,N_23145);
nor UO_2098 (O_2098,N_22762,N_22989);
nor UO_2099 (O_2099,N_23683,N_22649);
nor UO_2100 (O_2100,N_24974,N_23812);
and UO_2101 (O_2101,N_22502,N_22665);
nand UO_2102 (O_2102,N_22907,N_23275);
or UO_2103 (O_2103,N_23375,N_24792);
nand UO_2104 (O_2104,N_23525,N_22699);
nand UO_2105 (O_2105,N_23000,N_23827);
nand UO_2106 (O_2106,N_23641,N_22769);
nand UO_2107 (O_2107,N_22941,N_24627);
or UO_2108 (O_2108,N_22962,N_22743);
or UO_2109 (O_2109,N_24158,N_23024);
nand UO_2110 (O_2110,N_23612,N_24862);
xnor UO_2111 (O_2111,N_23280,N_24741);
or UO_2112 (O_2112,N_23326,N_24482);
and UO_2113 (O_2113,N_22756,N_24779);
xor UO_2114 (O_2114,N_24954,N_23204);
nor UO_2115 (O_2115,N_24753,N_23929);
nand UO_2116 (O_2116,N_23793,N_23707);
nand UO_2117 (O_2117,N_24307,N_23714);
and UO_2118 (O_2118,N_24363,N_24934);
or UO_2119 (O_2119,N_24908,N_23420);
nor UO_2120 (O_2120,N_24455,N_23853);
nand UO_2121 (O_2121,N_24157,N_24915);
nor UO_2122 (O_2122,N_24116,N_23361);
nor UO_2123 (O_2123,N_23512,N_24470);
xor UO_2124 (O_2124,N_22592,N_24287);
or UO_2125 (O_2125,N_24915,N_24189);
or UO_2126 (O_2126,N_22796,N_23333);
nand UO_2127 (O_2127,N_24290,N_23346);
and UO_2128 (O_2128,N_23653,N_24790);
nand UO_2129 (O_2129,N_23684,N_22874);
nand UO_2130 (O_2130,N_23198,N_23643);
nor UO_2131 (O_2131,N_23445,N_24029);
nand UO_2132 (O_2132,N_24074,N_24699);
and UO_2133 (O_2133,N_23257,N_22958);
nand UO_2134 (O_2134,N_23506,N_23582);
xnor UO_2135 (O_2135,N_23994,N_23304);
or UO_2136 (O_2136,N_23839,N_23070);
and UO_2137 (O_2137,N_24655,N_24260);
or UO_2138 (O_2138,N_23480,N_24746);
nor UO_2139 (O_2139,N_24615,N_24572);
nand UO_2140 (O_2140,N_22617,N_24955);
nand UO_2141 (O_2141,N_22633,N_24221);
and UO_2142 (O_2142,N_23696,N_22893);
and UO_2143 (O_2143,N_23035,N_22796);
nand UO_2144 (O_2144,N_22626,N_22517);
xor UO_2145 (O_2145,N_24943,N_24851);
or UO_2146 (O_2146,N_23473,N_24634);
and UO_2147 (O_2147,N_22667,N_24555);
nand UO_2148 (O_2148,N_24040,N_22971);
or UO_2149 (O_2149,N_24153,N_22864);
nor UO_2150 (O_2150,N_24540,N_24899);
or UO_2151 (O_2151,N_23357,N_23139);
and UO_2152 (O_2152,N_24271,N_23401);
xor UO_2153 (O_2153,N_24841,N_23297);
nand UO_2154 (O_2154,N_24319,N_22945);
or UO_2155 (O_2155,N_24364,N_24592);
and UO_2156 (O_2156,N_22657,N_24710);
and UO_2157 (O_2157,N_24881,N_23868);
nor UO_2158 (O_2158,N_24092,N_24024);
nor UO_2159 (O_2159,N_23066,N_24668);
or UO_2160 (O_2160,N_24209,N_24862);
or UO_2161 (O_2161,N_23795,N_22631);
or UO_2162 (O_2162,N_22959,N_24970);
and UO_2163 (O_2163,N_24255,N_23848);
or UO_2164 (O_2164,N_22959,N_23691);
nand UO_2165 (O_2165,N_22761,N_22751);
or UO_2166 (O_2166,N_24249,N_24944);
nor UO_2167 (O_2167,N_23606,N_23404);
nor UO_2168 (O_2168,N_23683,N_22758);
nor UO_2169 (O_2169,N_23190,N_23209);
nor UO_2170 (O_2170,N_23583,N_23068);
or UO_2171 (O_2171,N_22999,N_23352);
or UO_2172 (O_2172,N_24410,N_23805);
nand UO_2173 (O_2173,N_24948,N_23048);
and UO_2174 (O_2174,N_24167,N_24429);
or UO_2175 (O_2175,N_24528,N_23937);
nor UO_2176 (O_2176,N_23228,N_22766);
nor UO_2177 (O_2177,N_23323,N_24103);
and UO_2178 (O_2178,N_24760,N_23788);
and UO_2179 (O_2179,N_22847,N_23614);
nor UO_2180 (O_2180,N_23425,N_24882);
nand UO_2181 (O_2181,N_22558,N_23715);
nand UO_2182 (O_2182,N_24966,N_24618);
nand UO_2183 (O_2183,N_23496,N_23611);
and UO_2184 (O_2184,N_22549,N_24295);
nor UO_2185 (O_2185,N_22632,N_23145);
nand UO_2186 (O_2186,N_24522,N_24714);
and UO_2187 (O_2187,N_22529,N_24702);
and UO_2188 (O_2188,N_23945,N_24284);
or UO_2189 (O_2189,N_24220,N_23858);
and UO_2190 (O_2190,N_23925,N_22948);
or UO_2191 (O_2191,N_23295,N_23748);
nor UO_2192 (O_2192,N_23486,N_24982);
and UO_2193 (O_2193,N_23754,N_24586);
and UO_2194 (O_2194,N_24014,N_24165);
nand UO_2195 (O_2195,N_22565,N_24171);
nor UO_2196 (O_2196,N_24845,N_23382);
or UO_2197 (O_2197,N_23042,N_22977);
or UO_2198 (O_2198,N_24111,N_22718);
or UO_2199 (O_2199,N_22808,N_23390);
xnor UO_2200 (O_2200,N_22944,N_24594);
nor UO_2201 (O_2201,N_22633,N_23722);
nor UO_2202 (O_2202,N_22901,N_24809);
and UO_2203 (O_2203,N_23077,N_23934);
nor UO_2204 (O_2204,N_23887,N_22596);
and UO_2205 (O_2205,N_23039,N_22565);
and UO_2206 (O_2206,N_23561,N_23985);
and UO_2207 (O_2207,N_24757,N_24180);
or UO_2208 (O_2208,N_22786,N_22719);
nand UO_2209 (O_2209,N_24899,N_23013);
nand UO_2210 (O_2210,N_22969,N_23575);
xor UO_2211 (O_2211,N_24407,N_24919);
xnor UO_2212 (O_2212,N_24281,N_23059);
nand UO_2213 (O_2213,N_24453,N_24950);
or UO_2214 (O_2214,N_24270,N_24428);
and UO_2215 (O_2215,N_23478,N_24920);
or UO_2216 (O_2216,N_22654,N_23694);
and UO_2217 (O_2217,N_23544,N_24594);
or UO_2218 (O_2218,N_24382,N_24391);
nand UO_2219 (O_2219,N_23403,N_23184);
or UO_2220 (O_2220,N_22549,N_22536);
nand UO_2221 (O_2221,N_23834,N_24852);
xnor UO_2222 (O_2222,N_23653,N_24249);
and UO_2223 (O_2223,N_23957,N_24313);
or UO_2224 (O_2224,N_23564,N_22995);
or UO_2225 (O_2225,N_23987,N_23723);
nand UO_2226 (O_2226,N_24539,N_22911);
nor UO_2227 (O_2227,N_23338,N_22755);
nor UO_2228 (O_2228,N_22603,N_23202);
nor UO_2229 (O_2229,N_22888,N_22821);
xnor UO_2230 (O_2230,N_24166,N_24287);
and UO_2231 (O_2231,N_24164,N_23371);
and UO_2232 (O_2232,N_22777,N_23345);
nor UO_2233 (O_2233,N_23578,N_23738);
nand UO_2234 (O_2234,N_24826,N_24965);
nor UO_2235 (O_2235,N_24916,N_23141);
nand UO_2236 (O_2236,N_24252,N_22595);
nor UO_2237 (O_2237,N_24817,N_24317);
and UO_2238 (O_2238,N_22986,N_22524);
xnor UO_2239 (O_2239,N_23628,N_23769);
or UO_2240 (O_2240,N_24196,N_23036);
and UO_2241 (O_2241,N_24932,N_22823);
or UO_2242 (O_2242,N_23879,N_24206);
or UO_2243 (O_2243,N_22815,N_24507);
and UO_2244 (O_2244,N_23217,N_23039);
nor UO_2245 (O_2245,N_23976,N_23828);
or UO_2246 (O_2246,N_24661,N_24245);
nand UO_2247 (O_2247,N_22712,N_23207);
nor UO_2248 (O_2248,N_23916,N_24814);
nand UO_2249 (O_2249,N_23546,N_23961);
and UO_2250 (O_2250,N_22759,N_22546);
or UO_2251 (O_2251,N_24042,N_24697);
or UO_2252 (O_2252,N_22589,N_22980);
nand UO_2253 (O_2253,N_24071,N_23632);
or UO_2254 (O_2254,N_24944,N_23936);
or UO_2255 (O_2255,N_22583,N_22904);
nor UO_2256 (O_2256,N_22833,N_24407);
or UO_2257 (O_2257,N_22626,N_22964);
nor UO_2258 (O_2258,N_24521,N_24700);
nor UO_2259 (O_2259,N_24605,N_22956);
or UO_2260 (O_2260,N_24003,N_23698);
nand UO_2261 (O_2261,N_22548,N_23901);
nor UO_2262 (O_2262,N_23903,N_23628);
or UO_2263 (O_2263,N_22556,N_24598);
xor UO_2264 (O_2264,N_23219,N_22818);
nand UO_2265 (O_2265,N_23070,N_24646);
and UO_2266 (O_2266,N_23317,N_24619);
xnor UO_2267 (O_2267,N_24821,N_23424);
and UO_2268 (O_2268,N_23755,N_22545);
xnor UO_2269 (O_2269,N_24956,N_24620);
nor UO_2270 (O_2270,N_22801,N_23227);
nand UO_2271 (O_2271,N_24632,N_24559);
nand UO_2272 (O_2272,N_24653,N_24777);
or UO_2273 (O_2273,N_24470,N_22691);
or UO_2274 (O_2274,N_24466,N_23927);
xor UO_2275 (O_2275,N_24033,N_24952);
and UO_2276 (O_2276,N_22611,N_24388);
nor UO_2277 (O_2277,N_23053,N_24750);
xnor UO_2278 (O_2278,N_24048,N_24441);
nand UO_2279 (O_2279,N_24094,N_22579);
xnor UO_2280 (O_2280,N_22841,N_23770);
and UO_2281 (O_2281,N_24902,N_23977);
or UO_2282 (O_2282,N_24702,N_23584);
nor UO_2283 (O_2283,N_24840,N_23776);
nand UO_2284 (O_2284,N_23890,N_24402);
or UO_2285 (O_2285,N_23572,N_23220);
nand UO_2286 (O_2286,N_24378,N_23347);
nand UO_2287 (O_2287,N_24701,N_23072);
nand UO_2288 (O_2288,N_23396,N_24141);
xnor UO_2289 (O_2289,N_23130,N_23845);
or UO_2290 (O_2290,N_23943,N_22844);
xnor UO_2291 (O_2291,N_23696,N_23557);
nor UO_2292 (O_2292,N_23776,N_22896);
and UO_2293 (O_2293,N_23475,N_22545);
nor UO_2294 (O_2294,N_24055,N_24523);
nand UO_2295 (O_2295,N_24926,N_23394);
and UO_2296 (O_2296,N_24407,N_24082);
or UO_2297 (O_2297,N_23133,N_24643);
xor UO_2298 (O_2298,N_23044,N_23658);
nor UO_2299 (O_2299,N_23002,N_24832);
or UO_2300 (O_2300,N_24909,N_23248);
nor UO_2301 (O_2301,N_24238,N_24815);
or UO_2302 (O_2302,N_23561,N_22652);
or UO_2303 (O_2303,N_24657,N_24715);
nand UO_2304 (O_2304,N_22566,N_24425);
nand UO_2305 (O_2305,N_23451,N_22611);
or UO_2306 (O_2306,N_23171,N_24240);
and UO_2307 (O_2307,N_23822,N_24201);
nor UO_2308 (O_2308,N_23964,N_24821);
nand UO_2309 (O_2309,N_24455,N_24245);
and UO_2310 (O_2310,N_22838,N_24805);
nand UO_2311 (O_2311,N_24077,N_23694);
nor UO_2312 (O_2312,N_23724,N_24417);
or UO_2313 (O_2313,N_24047,N_24221);
nand UO_2314 (O_2314,N_24600,N_23554);
or UO_2315 (O_2315,N_23814,N_23009);
nor UO_2316 (O_2316,N_24689,N_23360);
nor UO_2317 (O_2317,N_24879,N_22607);
or UO_2318 (O_2318,N_24691,N_24478);
nor UO_2319 (O_2319,N_22728,N_22538);
nand UO_2320 (O_2320,N_24518,N_23438);
nand UO_2321 (O_2321,N_22656,N_24353);
and UO_2322 (O_2322,N_23940,N_22602);
nand UO_2323 (O_2323,N_23074,N_23872);
nor UO_2324 (O_2324,N_24431,N_22891);
nor UO_2325 (O_2325,N_22519,N_22588);
xnor UO_2326 (O_2326,N_23460,N_23168);
and UO_2327 (O_2327,N_22787,N_23775);
nor UO_2328 (O_2328,N_23971,N_24601);
nor UO_2329 (O_2329,N_24599,N_22760);
nor UO_2330 (O_2330,N_22717,N_23851);
and UO_2331 (O_2331,N_23817,N_24729);
nand UO_2332 (O_2332,N_24603,N_22663);
nor UO_2333 (O_2333,N_24624,N_24371);
xnor UO_2334 (O_2334,N_24670,N_24702);
nand UO_2335 (O_2335,N_22697,N_22997);
nand UO_2336 (O_2336,N_23989,N_22948);
nand UO_2337 (O_2337,N_24964,N_23988);
and UO_2338 (O_2338,N_23438,N_24954);
xor UO_2339 (O_2339,N_22503,N_22509);
nand UO_2340 (O_2340,N_23689,N_22888);
nand UO_2341 (O_2341,N_24874,N_22977);
and UO_2342 (O_2342,N_23414,N_24012);
and UO_2343 (O_2343,N_22585,N_24966);
nor UO_2344 (O_2344,N_22545,N_23749);
nand UO_2345 (O_2345,N_23641,N_24354);
nor UO_2346 (O_2346,N_24785,N_24583);
or UO_2347 (O_2347,N_22623,N_24223);
or UO_2348 (O_2348,N_23540,N_23359);
or UO_2349 (O_2349,N_24728,N_22851);
nor UO_2350 (O_2350,N_22573,N_23568);
or UO_2351 (O_2351,N_24866,N_24265);
or UO_2352 (O_2352,N_24780,N_24988);
nand UO_2353 (O_2353,N_24953,N_24117);
and UO_2354 (O_2354,N_23285,N_22994);
or UO_2355 (O_2355,N_22968,N_24194);
and UO_2356 (O_2356,N_22842,N_24171);
nor UO_2357 (O_2357,N_24423,N_24753);
nor UO_2358 (O_2358,N_24664,N_23659);
or UO_2359 (O_2359,N_24742,N_24011);
and UO_2360 (O_2360,N_23185,N_22552);
and UO_2361 (O_2361,N_24496,N_22860);
or UO_2362 (O_2362,N_24763,N_24676);
or UO_2363 (O_2363,N_24464,N_24813);
nor UO_2364 (O_2364,N_24099,N_22913);
nor UO_2365 (O_2365,N_24680,N_22581);
nor UO_2366 (O_2366,N_23242,N_23059);
and UO_2367 (O_2367,N_24488,N_23413);
and UO_2368 (O_2368,N_23238,N_24738);
or UO_2369 (O_2369,N_24158,N_24374);
nand UO_2370 (O_2370,N_24876,N_22931);
nor UO_2371 (O_2371,N_24792,N_24052);
and UO_2372 (O_2372,N_24330,N_23056);
and UO_2373 (O_2373,N_23893,N_23576);
or UO_2374 (O_2374,N_24985,N_24269);
or UO_2375 (O_2375,N_22800,N_24864);
nand UO_2376 (O_2376,N_23550,N_23720);
nand UO_2377 (O_2377,N_22918,N_22599);
or UO_2378 (O_2378,N_22792,N_23208);
nor UO_2379 (O_2379,N_24248,N_23095);
nand UO_2380 (O_2380,N_24263,N_23066);
nand UO_2381 (O_2381,N_23547,N_24464);
or UO_2382 (O_2382,N_22568,N_24382);
and UO_2383 (O_2383,N_23018,N_22933);
nor UO_2384 (O_2384,N_22930,N_22703);
xor UO_2385 (O_2385,N_23049,N_23704);
nand UO_2386 (O_2386,N_24864,N_22903);
or UO_2387 (O_2387,N_22684,N_23684);
nor UO_2388 (O_2388,N_24710,N_23722);
nand UO_2389 (O_2389,N_24140,N_23992);
nor UO_2390 (O_2390,N_24191,N_22561);
nand UO_2391 (O_2391,N_23694,N_22547);
nand UO_2392 (O_2392,N_24500,N_24753);
nor UO_2393 (O_2393,N_23967,N_23860);
xor UO_2394 (O_2394,N_22600,N_23183);
nor UO_2395 (O_2395,N_23290,N_23720);
nor UO_2396 (O_2396,N_23450,N_24604);
and UO_2397 (O_2397,N_23917,N_24476);
and UO_2398 (O_2398,N_22992,N_23901);
or UO_2399 (O_2399,N_23607,N_24842);
or UO_2400 (O_2400,N_23395,N_22997);
and UO_2401 (O_2401,N_23588,N_22509);
nor UO_2402 (O_2402,N_24182,N_24425);
and UO_2403 (O_2403,N_23175,N_24713);
nand UO_2404 (O_2404,N_23927,N_22709);
and UO_2405 (O_2405,N_22584,N_24220);
and UO_2406 (O_2406,N_24123,N_23085);
nand UO_2407 (O_2407,N_23625,N_23535);
and UO_2408 (O_2408,N_24344,N_24820);
xor UO_2409 (O_2409,N_23529,N_23820);
and UO_2410 (O_2410,N_23148,N_24346);
nand UO_2411 (O_2411,N_24824,N_22791);
and UO_2412 (O_2412,N_24797,N_24056);
and UO_2413 (O_2413,N_24818,N_24214);
nor UO_2414 (O_2414,N_23303,N_23618);
nand UO_2415 (O_2415,N_23590,N_22824);
or UO_2416 (O_2416,N_23336,N_23798);
nor UO_2417 (O_2417,N_22756,N_22740);
nand UO_2418 (O_2418,N_24043,N_22509);
nand UO_2419 (O_2419,N_22806,N_22531);
nor UO_2420 (O_2420,N_23644,N_22799);
or UO_2421 (O_2421,N_24784,N_24643);
xnor UO_2422 (O_2422,N_24924,N_24005);
and UO_2423 (O_2423,N_24128,N_22660);
or UO_2424 (O_2424,N_24269,N_23528);
and UO_2425 (O_2425,N_24101,N_24960);
nand UO_2426 (O_2426,N_23782,N_22894);
and UO_2427 (O_2427,N_23150,N_23679);
and UO_2428 (O_2428,N_24729,N_23924);
and UO_2429 (O_2429,N_23693,N_24409);
nor UO_2430 (O_2430,N_24549,N_24853);
and UO_2431 (O_2431,N_23735,N_23094);
xor UO_2432 (O_2432,N_24994,N_23526);
and UO_2433 (O_2433,N_24462,N_24986);
and UO_2434 (O_2434,N_24296,N_23920);
nand UO_2435 (O_2435,N_24803,N_23657);
or UO_2436 (O_2436,N_23544,N_22873);
or UO_2437 (O_2437,N_24328,N_24279);
and UO_2438 (O_2438,N_22990,N_23994);
nor UO_2439 (O_2439,N_23831,N_23575);
xor UO_2440 (O_2440,N_23435,N_23729);
or UO_2441 (O_2441,N_23013,N_24794);
and UO_2442 (O_2442,N_23394,N_24393);
or UO_2443 (O_2443,N_22697,N_23118);
and UO_2444 (O_2444,N_22577,N_23057);
and UO_2445 (O_2445,N_24171,N_23592);
nor UO_2446 (O_2446,N_22866,N_24936);
or UO_2447 (O_2447,N_22704,N_23560);
nor UO_2448 (O_2448,N_22645,N_24988);
and UO_2449 (O_2449,N_23458,N_22583);
and UO_2450 (O_2450,N_22548,N_24322);
and UO_2451 (O_2451,N_24265,N_24235);
xor UO_2452 (O_2452,N_23367,N_24356);
nor UO_2453 (O_2453,N_24903,N_23734);
xor UO_2454 (O_2454,N_22733,N_23931);
nor UO_2455 (O_2455,N_23754,N_22997);
nand UO_2456 (O_2456,N_24289,N_24519);
nor UO_2457 (O_2457,N_22738,N_23254);
nand UO_2458 (O_2458,N_24511,N_24970);
xnor UO_2459 (O_2459,N_24341,N_24787);
or UO_2460 (O_2460,N_24634,N_24473);
or UO_2461 (O_2461,N_24899,N_24334);
xor UO_2462 (O_2462,N_24707,N_23130);
nor UO_2463 (O_2463,N_23433,N_23829);
nor UO_2464 (O_2464,N_24340,N_22712);
nand UO_2465 (O_2465,N_23206,N_23098);
nor UO_2466 (O_2466,N_24974,N_22582);
and UO_2467 (O_2467,N_24724,N_23367);
or UO_2468 (O_2468,N_24730,N_23243);
nor UO_2469 (O_2469,N_23238,N_22658);
nor UO_2470 (O_2470,N_23319,N_22527);
and UO_2471 (O_2471,N_23445,N_24948);
and UO_2472 (O_2472,N_24787,N_24135);
nor UO_2473 (O_2473,N_23635,N_23949);
nor UO_2474 (O_2474,N_23867,N_23121);
nand UO_2475 (O_2475,N_23388,N_23596);
nand UO_2476 (O_2476,N_24606,N_22623);
nand UO_2477 (O_2477,N_23331,N_22749);
nand UO_2478 (O_2478,N_23804,N_23244);
xnor UO_2479 (O_2479,N_24138,N_23965);
xnor UO_2480 (O_2480,N_23445,N_23723);
or UO_2481 (O_2481,N_23134,N_24679);
nand UO_2482 (O_2482,N_23910,N_22682);
nor UO_2483 (O_2483,N_22898,N_23297);
or UO_2484 (O_2484,N_24264,N_23534);
xor UO_2485 (O_2485,N_23346,N_24519);
nor UO_2486 (O_2486,N_24765,N_22697);
nand UO_2487 (O_2487,N_23815,N_23671);
and UO_2488 (O_2488,N_24868,N_24960);
or UO_2489 (O_2489,N_22928,N_23298);
nor UO_2490 (O_2490,N_23662,N_24152);
or UO_2491 (O_2491,N_23451,N_22628);
nand UO_2492 (O_2492,N_24789,N_23989);
and UO_2493 (O_2493,N_22775,N_22970);
nor UO_2494 (O_2494,N_24944,N_23907);
and UO_2495 (O_2495,N_23656,N_24861);
and UO_2496 (O_2496,N_22502,N_24689);
and UO_2497 (O_2497,N_23019,N_24628);
or UO_2498 (O_2498,N_22781,N_23729);
and UO_2499 (O_2499,N_23267,N_23542);
or UO_2500 (O_2500,N_24741,N_24117);
xor UO_2501 (O_2501,N_24660,N_23427);
or UO_2502 (O_2502,N_23009,N_24899);
xor UO_2503 (O_2503,N_22870,N_23148);
or UO_2504 (O_2504,N_24783,N_24092);
nand UO_2505 (O_2505,N_24560,N_24734);
and UO_2506 (O_2506,N_23666,N_23524);
or UO_2507 (O_2507,N_22556,N_24422);
nor UO_2508 (O_2508,N_23523,N_23494);
nor UO_2509 (O_2509,N_23257,N_23266);
or UO_2510 (O_2510,N_24339,N_23870);
nand UO_2511 (O_2511,N_23150,N_22538);
xor UO_2512 (O_2512,N_24290,N_23856);
nand UO_2513 (O_2513,N_24379,N_23470);
nand UO_2514 (O_2514,N_23627,N_22637);
nor UO_2515 (O_2515,N_23157,N_23894);
and UO_2516 (O_2516,N_24444,N_24839);
and UO_2517 (O_2517,N_24024,N_22578);
and UO_2518 (O_2518,N_23113,N_23059);
or UO_2519 (O_2519,N_24894,N_23944);
nor UO_2520 (O_2520,N_23394,N_24766);
and UO_2521 (O_2521,N_24401,N_23612);
nand UO_2522 (O_2522,N_24412,N_23431);
or UO_2523 (O_2523,N_23008,N_23847);
xnor UO_2524 (O_2524,N_22771,N_23259);
nand UO_2525 (O_2525,N_23455,N_23467);
nand UO_2526 (O_2526,N_23907,N_24687);
or UO_2527 (O_2527,N_24460,N_24574);
or UO_2528 (O_2528,N_23859,N_24924);
or UO_2529 (O_2529,N_23300,N_23116);
and UO_2530 (O_2530,N_23281,N_23857);
and UO_2531 (O_2531,N_23708,N_22591);
and UO_2532 (O_2532,N_24688,N_24031);
and UO_2533 (O_2533,N_22645,N_23962);
or UO_2534 (O_2534,N_24228,N_22787);
and UO_2535 (O_2535,N_24019,N_24756);
xor UO_2536 (O_2536,N_24184,N_22747);
and UO_2537 (O_2537,N_23835,N_24832);
xor UO_2538 (O_2538,N_24669,N_24136);
or UO_2539 (O_2539,N_23461,N_23758);
nor UO_2540 (O_2540,N_24550,N_24726);
and UO_2541 (O_2541,N_23245,N_24668);
or UO_2542 (O_2542,N_24102,N_23187);
nor UO_2543 (O_2543,N_23790,N_23658);
and UO_2544 (O_2544,N_23189,N_24571);
nand UO_2545 (O_2545,N_24039,N_23355);
or UO_2546 (O_2546,N_24511,N_23610);
and UO_2547 (O_2547,N_24120,N_23642);
nor UO_2548 (O_2548,N_22541,N_24104);
nand UO_2549 (O_2549,N_23874,N_23774);
and UO_2550 (O_2550,N_24018,N_23025);
nand UO_2551 (O_2551,N_24283,N_22941);
nand UO_2552 (O_2552,N_23229,N_22818);
xor UO_2553 (O_2553,N_23507,N_24380);
and UO_2554 (O_2554,N_23782,N_23692);
and UO_2555 (O_2555,N_23900,N_24896);
nand UO_2556 (O_2556,N_24838,N_22511);
or UO_2557 (O_2557,N_24126,N_24401);
nand UO_2558 (O_2558,N_24011,N_24248);
nand UO_2559 (O_2559,N_23242,N_23153);
nand UO_2560 (O_2560,N_24057,N_24782);
nor UO_2561 (O_2561,N_23012,N_24296);
xnor UO_2562 (O_2562,N_23820,N_23823);
and UO_2563 (O_2563,N_24793,N_23814);
or UO_2564 (O_2564,N_23426,N_22972);
nor UO_2565 (O_2565,N_22561,N_24221);
xor UO_2566 (O_2566,N_23769,N_23481);
nor UO_2567 (O_2567,N_23264,N_23789);
nand UO_2568 (O_2568,N_24560,N_24914);
or UO_2569 (O_2569,N_23319,N_23140);
nor UO_2570 (O_2570,N_23844,N_22872);
or UO_2571 (O_2571,N_24168,N_24103);
nand UO_2572 (O_2572,N_23302,N_22777);
nand UO_2573 (O_2573,N_22748,N_23732);
and UO_2574 (O_2574,N_24332,N_24725);
nand UO_2575 (O_2575,N_23061,N_24524);
and UO_2576 (O_2576,N_24249,N_22782);
nor UO_2577 (O_2577,N_24271,N_23952);
and UO_2578 (O_2578,N_23393,N_24010);
nor UO_2579 (O_2579,N_23327,N_23656);
nor UO_2580 (O_2580,N_22863,N_23707);
nand UO_2581 (O_2581,N_24375,N_24262);
and UO_2582 (O_2582,N_24569,N_24581);
or UO_2583 (O_2583,N_22967,N_23675);
or UO_2584 (O_2584,N_24388,N_23710);
xor UO_2585 (O_2585,N_23785,N_23383);
or UO_2586 (O_2586,N_24938,N_22850);
xnor UO_2587 (O_2587,N_22594,N_24665);
and UO_2588 (O_2588,N_22606,N_23466);
or UO_2589 (O_2589,N_24315,N_24562);
and UO_2590 (O_2590,N_23639,N_24279);
nor UO_2591 (O_2591,N_23280,N_22575);
or UO_2592 (O_2592,N_23271,N_22993);
or UO_2593 (O_2593,N_24071,N_24912);
nand UO_2594 (O_2594,N_24885,N_22569);
nor UO_2595 (O_2595,N_23413,N_24061);
and UO_2596 (O_2596,N_22868,N_23689);
and UO_2597 (O_2597,N_23282,N_23048);
nor UO_2598 (O_2598,N_23547,N_23610);
nor UO_2599 (O_2599,N_22537,N_24377);
nand UO_2600 (O_2600,N_24909,N_22917);
or UO_2601 (O_2601,N_23471,N_23425);
xor UO_2602 (O_2602,N_23029,N_23616);
nand UO_2603 (O_2603,N_22789,N_23230);
nor UO_2604 (O_2604,N_23058,N_23295);
nor UO_2605 (O_2605,N_23800,N_22748);
xnor UO_2606 (O_2606,N_22528,N_24085);
and UO_2607 (O_2607,N_24062,N_24329);
and UO_2608 (O_2608,N_22563,N_23388);
nor UO_2609 (O_2609,N_22999,N_24768);
nor UO_2610 (O_2610,N_24420,N_24615);
nor UO_2611 (O_2611,N_24671,N_23215);
nor UO_2612 (O_2612,N_24633,N_23818);
xnor UO_2613 (O_2613,N_24824,N_24871);
nand UO_2614 (O_2614,N_23733,N_23967);
nand UO_2615 (O_2615,N_24529,N_24562);
or UO_2616 (O_2616,N_23965,N_23075);
and UO_2617 (O_2617,N_23664,N_24878);
or UO_2618 (O_2618,N_23455,N_23567);
or UO_2619 (O_2619,N_24085,N_24643);
nand UO_2620 (O_2620,N_23459,N_22727);
and UO_2621 (O_2621,N_24226,N_24878);
or UO_2622 (O_2622,N_22530,N_23489);
nor UO_2623 (O_2623,N_24040,N_23231);
nand UO_2624 (O_2624,N_24794,N_22897);
or UO_2625 (O_2625,N_22620,N_22715);
nand UO_2626 (O_2626,N_24101,N_22987);
or UO_2627 (O_2627,N_24759,N_23378);
and UO_2628 (O_2628,N_23087,N_22883);
xnor UO_2629 (O_2629,N_24634,N_23659);
xnor UO_2630 (O_2630,N_23152,N_23074);
nor UO_2631 (O_2631,N_23030,N_23361);
and UO_2632 (O_2632,N_23680,N_23432);
xor UO_2633 (O_2633,N_23354,N_24581);
and UO_2634 (O_2634,N_24634,N_23862);
and UO_2635 (O_2635,N_23007,N_24432);
nand UO_2636 (O_2636,N_24428,N_22562);
nand UO_2637 (O_2637,N_22565,N_24306);
or UO_2638 (O_2638,N_23322,N_23669);
or UO_2639 (O_2639,N_24911,N_23942);
and UO_2640 (O_2640,N_23582,N_23567);
and UO_2641 (O_2641,N_23875,N_23547);
nor UO_2642 (O_2642,N_24426,N_22818);
and UO_2643 (O_2643,N_24538,N_23501);
xnor UO_2644 (O_2644,N_23009,N_23258);
or UO_2645 (O_2645,N_23639,N_24923);
nand UO_2646 (O_2646,N_22695,N_23550);
nand UO_2647 (O_2647,N_22522,N_24980);
nor UO_2648 (O_2648,N_22987,N_23008);
xnor UO_2649 (O_2649,N_22862,N_22515);
and UO_2650 (O_2650,N_24451,N_24027);
and UO_2651 (O_2651,N_23062,N_22557);
xnor UO_2652 (O_2652,N_22512,N_23106);
nor UO_2653 (O_2653,N_23893,N_24956);
nor UO_2654 (O_2654,N_22576,N_24467);
xnor UO_2655 (O_2655,N_23411,N_24360);
and UO_2656 (O_2656,N_22796,N_23362);
or UO_2657 (O_2657,N_22628,N_23595);
or UO_2658 (O_2658,N_22802,N_24384);
or UO_2659 (O_2659,N_22670,N_24399);
or UO_2660 (O_2660,N_23689,N_23362);
nand UO_2661 (O_2661,N_24262,N_24642);
xnor UO_2662 (O_2662,N_24714,N_22519);
nor UO_2663 (O_2663,N_23901,N_22570);
nand UO_2664 (O_2664,N_22884,N_23196);
or UO_2665 (O_2665,N_24688,N_24673);
and UO_2666 (O_2666,N_24374,N_23770);
xnor UO_2667 (O_2667,N_23098,N_24245);
nand UO_2668 (O_2668,N_23302,N_23398);
nand UO_2669 (O_2669,N_23991,N_23092);
and UO_2670 (O_2670,N_23530,N_24185);
nand UO_2671 (O_2671,N_24372,N_24845);
nand UO_2672 (O_2672,N_24865,N_24703);
nand UO_2673 (O_2673,N_23797,N_23809);
nand UO_2674 (O_2674,N_24038,N_24681);
nand UO_2675 (O_2675,N_22830,N_23010);
and UO_2676 (O_2676,N_22865,N_22697);
nand UO_2677 (O_2677,N_23639,N_24054);
nand UO_2678 (O_2678,N_23750,N_22786);
nand UO_2679 (O_2679,N_24509,N_23528);
xor UO_2680 (O_2680,N_23606,N_24194);
nor UO_2681 (O_2681,N_24908,N_23626);
nor UO_2682 (O_2682,N_23283,N_22637);
nand UO_2683 (O_2683,N_23103,N_24895);
and UO_2684 (O_2684,N_23553,N_23295);
and UO_2685 (O_2685,N_22845,N_23752);
nand UO_2686 (O_2686,N_23072,N_22519);
nand UO_2687 (O_2687,N_22929,N_22827);
nand UO_2688 (O_2688,N_23131,N_23536);
and UO_2689 (O_2689,N_24349,N_22953);
and UO_2690 (O_2690,N_22850,N_23217);
nand UO_2691 (O_2691,N_23897,N_22974);
nor UO_2692 (O_2692,N_24878,N_22549);
xnor UO_2693 (O_2693,N_24555,N_23920);
and UO_2694 (O_2694,N_22562,N_23789);
or UO_2695 (O_2695,N_22743,N_22610);
or UO_2696 (O_2696,N_23130,N_23708);
nor UO_2697 (O_2697,N_22623,N_22699);
and UO_2698 (O_2698,N_24742,N_24933);
or UO_2699 (O_2699,N_23050,N_23476);
or UO_2700 (O_2700,N_22762,N_23634);
xnor UO_2701 (O_2701,N_24059,N_24831);
and UO_2702 (O_2702,N_23585,N_24082);
nor UO_2703 (O_2703,N_23031,N_23492);
nand UO_2704 (O_2704,N_24130,N_23671);
nor UO_2705 (O_2705,N_22929,N_24096);
or UO_2706 (O_2706,N_22909,N_23727);
nor UO_2707 (O_2707,N_23976,N_23677);
or UO_2708 (O_2708,N_24392,N_23933);
nand UO_2709 (O_2709,N_23674,N_24626);
nor UO_2710 (O_2710,N_24582,N_23151);
nand UO_2711 (O_2711,N_23023,N_24339);
and UO_2712 (O_2712,N_24106,N_23431);
nand UO_2713 (O_2713,N_24418,N_23173);
or UO_2714 (O_2714,N_24248,N_22504);
and UO_2715 (O_2715,N_23246,N_24035);
and UO_2716 (O_2716,N_23912,N_22949);
xnor UO_2717 (O_2717,N_23867,N_23953);
nand UO_2718 (O_2718,N_24559,N_23054);
nor UO_2719 (O_2719,N_23195,N_24886);
or UO_2720 (O_2720,N_23376,N_24279);
nand UO_2721 (O_2721,N_24321,N_23344);
nand UO_2722 (O_2722,N_24607,N_22657);
nand UO_2723 (O_2723,N_23575,N_22856);
and UO_2724 (O_2724,N_23450,N_24153);
or UO_2725 (O_2725,N_23398,N_24357);
or UO_2726 (O_2726,N_23598,N_23858);
and UO_2727 (O_2727,N_24189,N_24151);
and UO_2728 (O_2728,N_24447,N_23985);
and UO_2729 (O_2729,N_23659,N_22537);
and UO_2730 (O_2730,N_24879,N_23754);
nand UO_2731 (O_2731,N_22975,N_23322);
and UO_2732 (O_2732,N_23597,N_22830);
or UO_2733 (O_2733,N_24297,N_24402);
nand UO_2734 (O_2734,N_24827,N_22777);
nand UO_2735 (O_2735,N_23856,N_23146);
nor UO_2736 (O_2736,N_24581,N_23804);
nand UO_2737 (O_2737,N_22589,N_23829);
nand UO_2738 (O_2738,N_22516,N_22887);
or UO_2739 (O_2739,N_24541,N_24918);
nor UO_2740 (O_2740,N_23801,N_23139);
and UO_2741 (O_2741,N_22633,N_22529);
and UO_2742 (O_2742,N_22555,N_22883);
nand UO_2743 (O_2743,N_22861,N_24742);
nand UO_2744 (O_2744,N_24000,N_22999);
nand UO_2745 (O_2745,N_24527,N_24048);
or UO_2746 (O_2746,N_24782,N_23076);
nand UO_2747 (O_2747,N_22691,N_23294);
nand UO_2748 (O_2748,N_23522,N_24308);
xor UO_2749 (O_2749,N_22875,N_22731);
or UO_2750 (O_2750,N_23386,N_23999);
nand UO_2751 (O_2751,N_24745,N_22941);
nand UO_2752 (O_2752,N_24883,N_24161);
or UO_2753 (O_2753,N_23752,N_23922);
and UO_2754 (O_2754,N_22679,N_24960);
or UO_2755 (O_2755,N_23640,N_24304);
nand UO_2756 (O_2756,N_24412,N_23763);
or UO_2757 (O_2757,N_24002,N_23142);
nand UO_2758 (O_2758,N_23856,N_24293);
nand UO_2759 (O_2759,N_23328,N_24651);
xnor UO_2760 (O_2760,N_22978,N_22996);
nor UO_2761 (O_2761,N_23524,N_24492);
nand UO_2762 (O_2762,N_24174,N_22558);
xor UO_2763 (O_2763,N_24644,N_24538);
nor UO_2764 (O_2764,N_24959,N_24491);
nand UO_2765 (O_2765,N_23438,N_23063);
nor UO_2766 (O_2766,N_24445,N_22546);
nand UO_2767 (O_2767,N_23685,N_24400);
nand UO_2768 (O_2768,N_22976,N_23461);
nor UO_2769 (O_2769,N_24183,N_23557);
nor UO_2770 (O_2770,N_24920,N_24077);
nand UO_2771 (O_2771,N_23948,N_24078);
xnor UO_2772 (O_2772,N_23149,N_24060);
nor UO_2773 (O_2773,N_23478,N_23483);
nor UO_2774 (O_2774,N_23427,N_24777);
nor UO_2775 (O_2775,N_24340,N_23767);
or UO_2776 (O_2776,N_23564,N_24219);
or UO_2777 (O_2777,N_23440,N_23606);
nand UO_2778 (O_2778,N_24252,N_24080);
xor UO_2779 (O_2779,N_22725,N_23612);
or UO_2780 (O_2780,N_24979,N_22626);
nand UO_2781 (O_2781,N_22941,N_23423);
nand UO_2782 (O_2782,N_24461,N_23269);
xnor UO_2783 (O_2783,N_24253,N_24295);
and UO_2784 (O_2784,N_24912,N_22992);
and UO_2785 (O_2785,N_23628,N_24382);
xor UO_2786 (O_2786,N_23940,N_23022);
nand UO_2787 (O_2787,N_22602,N_24057);
nand UO_2788 (O_2788,N_23163,N_24611);
nor UO_2789 (O_2789,N_23393,N_22808);
xor UO_2790 (O_2790,N_24091,N_24445);
nand UO_2791 (O_2791,N_24389,N_24976);
or UO_2792 (O_2792,N_24962,N_24614);
or UO_2793 (O_2793,N_24234,N_23947);
or UO_2794 (O_2794,N_24858,N_24417);
xor UO_2795 (O_2795,N_23156,N_22867);
or UO_2796 (O_2796,N_23747,N_24818);
nand UO_2797 (O_2797,N_24349,N_23832);
or UO_2798 (O_2798,N_24158,N_24989);
and UO_2799 (O_2799,N_23717,N_24021);
nor UO_2800 (O_2800,N_23598,N_23142);
nand UO_2801 (O_2801,N_22803,N_24236);
or UO_2802 (O_2802,N_23313,N_23301);
nand UO_2803 (O_2803,N_24515,N_22927);
or UO_2804 (O_2804,N_23078,N_24205);
nand UO_2805 (O_2805,N_23921,N_24293);
or UO_2806 (O_2806,N_23306,N_23797);
xor UO_2807 (O_2807,N_24104,N_24527);
or UO_2808 (O_2808,N_23660,N_24198);
nor UO_2809 (O_2809,N_24018,N_23884);
xor UO_2810 (O_2810,N_24926,N_22603);
nand UO_2811 (O_2811,N_24488,N_23122);
nor UO_2812 (O_2812,N_24113,N_23770);
and UO_2813 (O_2813,N_22693,N_22819);
nand UO_2814 (O_2814,N_24332,N_24541);
nand UO_2815 (O_2815,N_23479,N_23260);
nor UO_2816 (O_2816,N_22556,N_23758);
and UO_2817 (O_2817,N_22788,N_23866);
and UO_2818 (O_2818,N_23634,N_24350);
nand UO_2819 (O_2819,N_22965,N_24215);
nand UO_2820 (O_2820,N_22664,N_24039);
or UO_2821 (O_2821,N_23253,N_24041);
xor UO_2822 (O_2822,N_24769,N_23951);
or UO_2823 (O_2823,N_24921,N_24438);
and UO_2824 (O_2824,N_22830,N_24066);
nor UO_2825 (O_2825,N_24932,N_22649);
or UO_2826 (O_2826,N_22979,N_24163);
or UO_2827 (O_2827,N_22965,N_24333);
nand UO_2828 (O_2828,N_24945,N_23308);
and UO_2829 (O_2829,N_22713,N_24729);
nor UO_2830 (O_2830,N_22586,N_23819);
nor UO_2831 (O_2831,N_24835,N_24520);
nor UO_2832 (O_2832,N_23128,N_22571);
or UO_2833 (O_2833,N_24129,N_24210);
nand UO_2834 (O_2834,N_22613,N_24777);
or UO_2835 (O_2835,N_24992,N_23163);
nand UO_2836 (O_2836,N_22838,N_24180);
nand UO_2837 (O_2837,N_22645,N_23544);
xor UO_2838 (O_2838,N_22751,N_22508);
nor UO_2839 (O_2839,N_24941,N_23622);
nand UO_2840 (O_2840,N_24464,N_24139);
nor UO_2841 (O_2841,N_22955,N_24461);
xnor UO_2842 (O_2842,N_22621,N_24373);
or UO_2843 (O_2843,N_23413,N_24352);
nor UO_2844 (O_2844,N_22560,N_23441);
and UO_2845 (O_2845,N_24069,N_24724);
or UO_2846 (O_2846,N_24312,N_24976);
and UO_2847 (O_2847,N_24856,N_24536);
or UO_2848 (O_2848,N_22527,N_24706);
xnor UO_2849 (O_2849,N_23733,N_24579);
nor UO_2850 (O_2850,N_23832,N_23727);
and UO_2851 (O_2851,N_23986,N_24037);
and UO_2852 (O_2852,N_24080,N_23574);
or UO_2853 (O_2853,N_22986,N_23459);
nor UO_2854 (O_2854,N_23798,N_24352);
or UO_2855 (O_2855,N_23481,N_23353);
and UO_2856 (O_2856,N_23687,N_23413);
or UO_2857 (O_2857,N_24292,N_23060);
and UO_2858 (O_2858,N_24915,N_22505);
nor UO_2859 (O_2859,N_22721,N_23687);
nor UO_2860 (O_2860,N_22637,N_23537);
or UO_2861 (O_2861,N_23373,N_23291);
xnor UO_2862 (O_2862,N_24647,N_24240);
or UO_2863 (O_2863,N_23900,N_24601);
nor UO_2864 (O_2864,N_23796,N_22535);
or UO_2865 (O_2865,N_24942,N_23458);
xor UO_2866 (O_2866,N_23266,N_24216);
or UO_2867 (O_2867,N_24483,N_24127);
nor UO_2868 (O_2868,N_23730,N_22943);
nand UO_2869 (O_2869,N_23259,N_24223);
nor UO_2870 (O_2870,N_24646,N_22819);
or UO_2871 (O_2871,N_23046,N_23949);
nand UO_2872 (O_2872,N_24679,N_24932);
nand UO_2873 (O_2873,N_24855,N_22810);
and UO_2874 (O_2874,N_22536,N_22728);
nand UO_2875 (O_2875,N_24559,N_24800);
and UO_2876 (O_2876,N_24508,N_23301);
nor UO_2877 (O_2877,N_24967,N_24525);
or UO_2878 (O_2878,N_22944,N_23982);
or UO_2879 (O_2879,N_23833,N_24813);
xnor UO_2880 (O_2880,N_24877,N_22930);
or UO_2881 (O_2881,N_23077,N_24533);
nor UO_2882 (O_2882,N_23939,N_23677);
or UO_2883 (O_2883,N_23292,N_24152);
nor UO_2884 (O_2884,N_24585,N_22977);
or UO_2885 (O_2885,N_22510,N_22915);
xnor UO_2886 (O_2886,N_23971,N_23676);
or UO_2887 (O_2887,N_23959,N_23933);
nand UO_2888 (O_2888,N_24721,N_24269);
or UO_2889 (O_2889,N_24923,N_23480);
or UO_2890 (O_2890,N_24417,N_23505);
and UO_2891 (O_2891,N_22797,N_23096);
and UO_2892 (O_2892,N_22653,N_24694);
or UO_2893 (O_2893,N_23244,N_23452);
or UO_2894 (O_2894,N_24497,N_23415);
or UO_2895 (O_2895,N_22719,N_24547);
nand UO_2896 (O_2896,N_23568,N_23677);
nor UO_2897 (O_2897,N_24866,N_24026);
nand UO_2898 (O_2898,N_23813,N_22938);
nor UO_2899 (O_2899,N_23318,N_22774);
nand UO_2900 (O_2900,N_24837,N_23863);
or UO_2901 (O_2901,N_24898,N_24999);
nand UO_2902 (O_2902,N_22879,N_24352);
xnor UO_2903 (O_2903,N_22613,N_22697);
nor UO_2904 (O_2904,N_23109,N_22817);
and UO_2905 (O_2905,N_23600,N_24926);
or UO_2906 (O_2906,N_23769,N_24938);
nor UO_2907 (O_2907,N_24172,N_23551);
nand UO_2908 (O_2908,N_24824,N_24972);
and UO_2909 (O_2909,N_23160,N_22854);
xor UO_2910 (O_2910,N_22588,N_23629);
and UO_2911 (O_2911,N_22747,N_24649);
xor UO_2912 (O_2912,N_24872,N_24492);
xnor UO_2913 (O_2913,N_24874,N_24404);
nand UO_2914 (O_2914,N_24939,N_23851);
nor UO_2915 (O_2915,N_24166,N_23300);
nor UO_2916 (O_2916,N_23587,N_23025);
nor UO_2917 (O_2917,N_22551,N_24253);
or UO_2918 (O_2918,N_23590,N_24735);
nor UO_2919 (O_2919,N_23082,N_23529);
and UO_2920 (O_2920,N_23846,N_24963);
nand UO_2921 (O_2921,N_23326,N_23764);
nor UO_2922 (O_2922,N_24477,N_23659);
or UO_2923 (O_2923,N_22668,N_24464);
or UO_2924 (O_2924,N_24550,N_23771);
or UO_2925 (O_2925,N_24324,N_22749);
nor UO_2926 (O_2926,N_23728,N_24032);
nor UO_2927 (O_2927,N_22591,N_23519);
nor UO_2928 (O_2928,N_24578,N_23702);
and UO_2929 (O_2929,N_24555,N_22949);
nor UO_2930 (O_2930,N_22794,N_23111);
nand UO_2931 (O_2931,N_24079,N_23673);
or UO_2932 (O_2932,N_22877,N_24060);
and UO_2933 (O_2933,N_23483,N_22715);
nor UO_2934 (O_2934,N_24680,N_22630);
or UO_2935 (O_2935,N_23040,N_23267);
and UO_2936 (O_2936,N_23413,N_23764);
and UO_2937 (O_2937,N_23829,N_23787);
nand UO_2938 (O_2938,N_23620,N_23773);
and UO_2939 (O_2939,N_23642,N_22577);
or UO_2940 (O_2940,N_22992,N_22791);
and UO_2941 (O_2941,N_23937,N_23465);
or UO_2942 (O_2942,N_22688,N_23718);
nor UO_2943 (O_2943,N_24408,N_24886);
and UO_2944 (O_2944,N_24126,N_24546);
nor UO_2945 (O_2945,N_24172,N_24394);
and UO_2946 (O_2946,N_22551,N_23315);
and UO_2947 (O_2947,N_24120,N_23257);
nand UO_2948 (O_2948,N_24486,N_23519);
nor UO_2949 (O_2949,N_22914,N_24559);
or UO_2950 (O_2950,N_22836,N_24652);
nand UO_2951 (O_2951,N_23522,N_24852);
and UO_2952 (O_2952,N_23478,N_24926);
nor UO_2953 (O_2953,N_23796,N_22890);
or UO_2954 (O_2954,N_24731,N_22698);
and UO_2955 (O_2955,N_24822,N_22982);
or UO_2956 (O_2956,N_24953,N_24934);
or UO_2957 (O_2957,N_24797,N_23248);
nor UO_2958 (O_2958,N_23983,N_22603);
or UO_2959 (O_2959,N_23375,N_24028);
nand UO_2960 (O_2960,N_24083,N_23664);
or UO_2961 (O_2961,N_22855,N_24481);
nand UO_2962 (O_2962,N_23319,N_23135);
and UO_2963 (O_2963,N_23177,N_24040);
nor UO_2964 (O_2964,N_24363,N_23281);
nand UO_2965 (O_2965,N_22960,N_23835);
or UO_2966 (O_2966,N_24232,N_24870);
nand UO_2967 (O_2967,N_23134,N_23008);
nand UO_2968 (O_2968,N_24087,N_24476);
nand UO_2969 (O_2969,N_23617,N_23674);
nor UO_2970 (O_2970,N_24593,N_23717);
nand UO_2971 (O_2971,N_23372,N_23326);
or UO_2972 (O_2972,N_23234,N_23719);
xnor UO_2973 (O_2973,N_24026,N_24828);
and UO_2974 (O_2974,N_23319,N_24080);
nor UO_2975 (O_2975,N_23309,N_23896);
nor UO_2976 (O_2976,N_23674,N_24147);
nand UO_2977 (O_2977,N_23948,N_24024);
nor UO_2978 (O_2978,N_22612,N_22944);
nor UO_2979 (O_2979,N_24581,N_23833);
and UO_2980 (O_2980,N_23493,N_22692);
or UO_2981 (O_2981,N_23304,N_24228);
xor UO_2982 (O_2982,N_24025,N_23303);
or UO_2983 (O_2983,N_22608,N_24563);
and UO_2984 (O_2984,N_24699,N_23516);
and UO_2985 (O_2985,N_24716,N_24519);
nand UO_2986 (O_2986,N_22963,N_23604);
nor UO_2987 (O_2987,N_22946,N_24857);
nor UO_2988 (O_2988,N_24334,N_24103);
nor UO_2989 (O_2989,N_23031,N_23342);
nand UO_2990 (O_2990,N_22571,N_24855);
and UO_2991 (O_2991,N_22728,N_24155);
and UO_2992 (O_2992,N_24601,N_23290);
and UO_2993 (O_2993,N_22561,N_24374);
nand UO_2994 (O_2994,N_24924,N_23392);
or UO_2995 (O_2995,N_22610,N_22811);
or UO_2996 (O_2996,N_23527,N_23551);
nand UO_2997 (O_2997,N_24402,N_22768);
and UO_2998 (O_2998,N_22857,N_23405);
xnor UO_2999 (O_2999,N_22919,N_22725);
endmodule