module basic_2000_20000_2500_20_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_524,In_369);
or U1 (N_1,In_209,In_1146);
nand U2 (N_2,In_1048,In_1788);
nand U3 (N_3,In_408,In_304);
nand U4 (N_4,In_47,In_980);
xnor U5 (N_5,In_814,In_453);
or U6 (N_6,In_1630,In_1815);
or U7 (N_7,In_997,In_40);
nor U8 (N_8,In_225,In_1879);
nor U9 (N_9,In_538,In_1076);
nor U10 (N_10,In_1626,In_574);
or U11 (N_11,In_3,In_1827);
nor U12 (N_12,In_1,In_398);
and U13 (N_13,In_1047,In_1571);
xor U14 (N_14,In_728,In_1331);
and U15 (N_15,In_1316,In_1245);
and U16 (N_16,In_1195,In_1727);
nor U17 (N_17,In_45,In_1337);
xnor U18 (N_18,In_698,In_833);
and U19 (N_19,In_745,In_1575);
nand U20 (N_20,In_1540,In_509);
and U21 (N_21,In_106,In_135);
nor U22 (N_22,In_709,In_1443);
and U23 (N_23,In_703,In_1394);
nor U24 (N_24,In_1028,In_542);
and U25 (N_25,In_1738,In_1233);
xnor U26 (N_26,In_1003,In_971);
and U27 (N_27,In_1825,In_314);
xor U28 (N_28,In_1932,In_400);
xor U29 (N_29,In_216,In_1034);
nor U30 (N_30,In_1545,In_1618);
nand U31 (N_31,In_361,In_1105);
or U32 (N_32,In_245,In_534);
nor U33 (N_33,In_1033,In_390);
or U34 (N_34,In_202,In_769);
xor U35 (N_35,In_1787,In_994);
and U36 (N_36,In_802,In_1186);
nand U37 (N_37,In_1160,In_562);
nand U38 (N_38,In_374,In_1933);
and U39 (N_39,In_146,In_322);
xor U40 (N_40,In_131,In_1396);
xnor U41 (N_41,In_1684,In_179);
nand U42 (N_42,In_1696,In_1771);
xor U43 (N_43,In_778,In_1949);
nand U44 (N_44,In_1361,In_142);
nand U45 (N_45,In_1594,In_1353);
nor U46 (N_46,In_1658,In_662);
nor U47 (N_47,In_1145,In_1728);
xnor U48 (N_48,In_63,In_1835);
nand U49 (N_49,In_485,In_1668);
nand U50 (N_50,In_1107,In_1050);
nand U51 (N_51,In_439,In_244);
nand U52 (N_52,In_960,In_46);
nand U53 (N_53,In_1924,In_1633);
xnor U54 (N_54,In_850,In_1081);
or U55 (N_55,In_53,In_1373);
or U56 (N_56,In_1561,In_1487);
or U57 (N_57,In_1600,In_729);
nor U58 (N_58,In_672,In_354);
and U59 (N_59,In_78,In_760);
xnor U60 (N_60,In_1972,In_1855);
and U61 (N_61,In_176,In_868);
and U62 (N_62,In_1467,In_804);
xor U63 (N_63,In_1976,In_1007);
nand U64 (N_64,In_1072,In_861);
xnor U65 (N_65,In_305,In_1357);
and U66 (N_66,In_811,In_1180);
and U67 (N_67,In_1139,In_1411);
nor U68 (N_68,In_325,In_221);
and U69 (N_69,In_1015,In_1438);
xor U70 (N_70,In_1816,In_1168);
nor U71 (N_71,In_704,In_264);
and U72 (N_72,In_742,In_1413);
xnor U73 (N_73,In_1100,In_1277);
nand U74 (N_74,In_1650,In_955);
or U75 (N_75,In_123,In_270);
and U76 (N_76,In_1629,In_535);
nand U77 (N_77,In_829,In_1836);
xor U78 (N_78,In_90,In_883);
and U79 (N_79,In_675,In_1150);
and U80 (N_80,In_1884,In_1780);
nand U81 (N_81,In_1607,In_1395);
nor U82 (N_82,In_1334,In_519);
xnor U83 (N_83,In_1243,In_824);
or U84 (N_84,In_681,In_1442);
nor U85 (N_85,In_1420,In_1310);
xor U86 (N_86,In_413,In_251);
xor U87 (N_87,In_1799,In_483);
or U88 (N_88,In_1124,In_281);
nand U89 (N_89,In_1235,In_191);
and U90 (N_90,In_347,In_855);
and U91 (N_91,In_1843,In_284);
and U92 (N_92,In_273,In_472);
nand U93 (N_93,In_1197,In_1426);
and U94 (N_94,In_1770,In_1225);
xnor U95 (N_95,In_1640,In_492);
xor U96 (N_96,In_1117,In_1409);
and U97 (N_97,In_1616,In_197);
nor U98 (N_98,In_1376,In_1000);
xor U99 (N_99,In_88,In_1120);
and U100 (N_100,In_114,In_421);
xnor U101 (N_101,In_1911,In_1522);
nand U102 (N_102,In_1742,In_1937);
xor U103 (N_103,In_302,In_1489);
nand U104 (N_104,In_531,In_1380);
or U105 (N_105,In_838,In_1868);
xnor U106 (N_106,In_1385,In_1130);
nand U107 (N_107,In_1639,In_89);
xor U108 (N_108,In_1214,In_1682);
xor U109 (N_109,In_882,In_185);
nor U110 (N_110,In_1109,In_1758);
or U111 (N_111,In_1590,In_1716);
xor U112 (N_112,In_1326,In_1404);
nand U113 (N_113,In_1025,In_324);
nor U114 (N_114,In_661,In_194);
xnor U115 (N_115,In_1427,In_169);
nor U116 (N_116,In_461,In_1917);
and U117 (N_117,In_611,In_1991);
or U118 (N_118,In_490,In_671);
and U119 (N_119,In_864,In_1269);
xnor U120 (N_120,In_1024,In_1756);
or U121 (N_121,In_514,In_207);
or U122 (N_122,In_392,In_1469);
or U123 (N_123,In_1656,In_344);
xor U124 (N_124,In_523,In_388);
nand U125 (N_125,In_1667,In_1169);
nand U126 (N_126,In_712,In_1273);
xor U127 (N_127,In_1906,In_77);
xor U128 (N_128,In_101,In_1244);
or U129 (N_129,In_1603,In_1913);
or U130 (N_130,In_1206,In_1803);
and U131 (N_131,In_1191,In_1448);
xor U132 (N_132,In_904,In_1903);
and U133 (N_133,In_692,In_628);
and U134 (N_134,In_283,In_480);
nor U135 (N_135,In_1986,In_899);
and U136 (N_136,In_617,In_504);
or U137 (N_137,In_370,In_1615);
and U138 (N_138,In_890,In_260);
nor U139 (N_139,In_342,In_177);
and U140 (N_140,In_637,In_580);
xnor U141 (N_141,In_1637,In_409);
and U142 (N_142,In_1905,In_1088);
or U143 (N_143,In_1265,In_1506);
nor U144 (N_144,In_1956,In_913);
or U145 (N_145,In_642,In_685);
nor U146 (N_146,In_1773,In_1829);
or U147 (N_147,In_1959,In_20);
xor U148 (N_148,In_67,In_1013);
xnor U149 (N_149,In_764,In_1445);
or U150 (N_150,In_276,In_426);
xnor U151 (N_151,In_639,In_998);
or U152 (N_152,In_1189,In_1256);
xnor U153 (N_153,In_1355,In_189);
xnor U154 (N_154,In_740,In_856);
xnor U155 (N_155,In_640,In_964);
and U156 (N_156,In_1020,In_1444);
and U157 (N_157,In_350,In_834);
and U158 (N_158,In_863,In_1468);
and U159 (N_159,In_1203,In_290);
nor U160 (N_160,In_502,In_820);
or U161 (N_161,In_911,In_1270);
and U162 (N_162,In_1695,In_1094);
nand U163 (N_163,In_567,In_1705);
nor U164 (N_164,In_1982,In_756);
or U165 (N_165,In_1557,In_1926);
and U166 (N_166,In_1565,In_1812);
or U167 (N_167,In_239,In_102);
nand U168 (N_168,In_719,In_551);
nand U169 (N_169,In_262,In_86);
xor U170 (N_170,In_946,In_404);
and U171 (N_171,In_1838,In_1957);
xor U172 (N_172,In_233,In_690);
nand U173 (N_173,In_99,In_240);
or U174 (N_174,In_847,In_109);
nor U175 (N_175,In_291,In_635);
and U176 (N_176,In_1674,In_1625);
and U177 (N_177,In_859,In_633);
and U178 (N_178,In_1934,In_949);
or U179 (N_179,In_795,In_593);
or U180 (N_180,In_1889,In_156);
xnor U181 (N_181,In_487,In_1818);
nand U182 (N_182,In_407,In_30);
nor U183 (N_183,In_1927,In_1649);
and U184 (N_184,In_1017,In_765);
or U185 (N_185,In_1001,In_235);
nor U186 (N_186,In_1741,In_1176);
or U187 (N_187,In_926,In_1069);
nand U188 (N_188,In_1755,In_1258);
xor U189 (N_189,In_560,In_1623);
nand U190 (N_190,In_1832,In_1499);
nor U191 (N_191,In_1211,In_1401);
nand U192 (N_192,In_1526,In_296);
nor U193 (N_193,In_1285,In_1782);
and U194 (N_194,In_1200,In_668);
and U195 (N_195,In_1046,In_1645);
xor U196 (N_196,In_1450,In_1582);
or U197 (N_197,In_1447,In_1089);
nor U198 (N_198,In_1227,In_1481);
nor U199 (N_199,In_1054,In_1188);
nand U200 (N_200,In_1282,In_1946);
and U201 (N_201,In_1052,In_1480);
nor U202 (N_202,In_1463,In_153);
or U203 (N_203,In_1477,In_585);
nor U204 (N_204,In_351,In_813);
nand U205 (N_205,In_1091,In_1987);
xnor U206 (N_206,In_1019,In_1599);
or U207 (N_207,In_320,In_190);
and U208 (N_208,In_13,In_1605);
nand U209 (N_209,In_992,In_103);
or U210 (N_210,In_1318,In_973);
xor U211 (N_211,In_1457,In_584);
or U212 (N_212,In_237,In_696);
xor U213 (N_213,In_410,In_1267);
xnor U214 (N_214,In_1985,In_1407);
nand U215 (N_215,In_918,In_718);
xnor U216 (N_216,In_880,In_1722);
or U217 (N_217,In_1171,In_770);
and U218 (N_218,In_1440,In_1979);
and U219 (N_219,In_1711,In_1657);
nor U220 (N_220,In_282,In_1164);
nand U221 (N_221,In_601,In_910);
nor U222 (N_222,In_462,In_348);
xor U223 (N_223,In_817,In_674);
xnor U224 (N_224,In_1663,In_766);
nor U225 (N_225,In_916,In_945);
nor U226 (N_226,In_1056,In_876);
or U227 (N_227,In_1064,In_1205);
nand U228 (N_228,In_1627,In_878);
xor U229 (N_229,In_1786,In_921);
and U230 (N_230,In_822,In_371);
or U231 (N_231,In_943,In_1939);
nand U232 (N_232,In_1867,In_697);
nor U233 (N_233,In_1184,In_749);
and U234 (N_234,In_902,In_211);
and U235 (N_235,In_775,In_1037);
nand U236 (N_236,In_1199,In_938);
xor U237 (N_237,In_1286,In_1390);
nand U238 (N_238,In_1495,In_1482);
nand U239 (N_239,In_29,In_139);
nor U240 (N_240,In_184,In_1324);
or U241 (N_241,In_160,In_446);
nand U242 (N_242,In_1043,In_615);
nor U243 (N_243,In_1701,In_653);
nor U244 (N_244,In_1769,In_612);
xor U245 (N_245,In_75,In_1366);
and U246 (N_246,In_1909,In_1814);
nand U247 (N_247,In_1485,In_1356);
and U248 (N_248,In_1430,In_1058);
and U249 (N_249,In_631,In_1521);
and U250 (N_250,In_482,In_35);
or U251 (N_251,In_17,In_1178);
nand U252 (N_252,In_1008,In_1121);
and U253 (N_253,In_693,In_1789);
nand U254 (N_254,In_1309,In_269);
xnor U255 (N_255,In_571,In_1740);
xnor U256 (N_256,In_605,In_118);
and U257 (N_257,In_1938,In_1219);
or U258 (N_258,In_489,In_725);
nand U259 (N_259,In_1071,In_1347);
nand U260 (N_260,In_1067,In_1510);
and U261 (N_261,In_708,In_1408);
nor U262 (N_262,In_816,In_1116);
or U263 (N_263,In_1023,In_893);
nand U264 (N_264,In_66,In_1079);
nor U265 (N_265,In_1614,In_1768);
xnor U266 (N_266,In_117,In_1317);
nand U267 (N_267,In_223,In_1472);
and U268 (N_268,In_10,In_1876);
xor U269 (N_269,In_23,In_985);
xnor U270 (N_270,In_1719,In_1846);
and U271 (N_271,In_1149,In_111);
nor U272 (N_272,In_1735,In_217);
or U273 (N_273,In_331,In_944);
or U274 (N_274,In_572,In_843);
xor U275 (N_275,In_1830,In_1399);
xor U276 (N_276,In_1453,In_1004);
nor U277 (N_277,In_1246,In_437);
and U278 (N_278,In_1950,In_832);
or U279 (N_279,In_157,In_430);
and U280 (N_280,In_345,In_638);
and U281 (N_281,In_4,In_48);
xor U282 (N_282,In_1672,In_1988);
and U283 (N_283,In_1921,In_1563);
xor U284 (N_284,In_1496,In_214);
or U285 (N_285,In_552,In_199);
nor U286 (N_286,In_1881,In_137);
and U287 (N_287,In_1371,In_1275);
nand U288 (N_288,In_108,In_1305);
nand U289 (N_289,In_181,In_588);
nor U290 (N_290,In_508,In_312);
and U291 (N_291,In_475,In_1170);
or U292 (N_292,In_1055,In_1210);
or U293 (N_293,In_1307,In_1288);
or U294 (N_294,In_1204,In_313);
nor U295 (N_295,In_752,In_1570);
xor U296 (N_296,In_730,In_866);
or U297 (N_297,In_397,In_620);
nand U298 (N_298,In_734,In_1009);
and U299 (N_299,In_839,In_1652);
and U300 (N_300,In_983,In_1462);
xnor U301 (N_301,In_555,In_546);
xnor U302 (N_302,In_1250,In_1359);
or U303 (N_303,In_1961,In_1473);
xnor U304 (N_304,In_791,In_1382);
or U305 (N_305,In_301,In_1147);
nor U306 (N_306,In_1429,In_138);
xnor U307 (N_307,In_19,In_321);
nand U308 (N_308,In_1108,In_1029);
and U309 (N_309,In_815,In_1777);
or U310 (N_310,In_423,In_1391);
or U311 (N_311,In_254,In_606);
nor U312 (N_312,In_1389,In_1894);
or U313 (N_313,In_1266,In_1923);
or U314 (N_314,In_129,In_933);
nor U315 (N_315,In_1252,In_96);
nor U316 (N_316,In_540,In_989);
or U317 (N_317,In_846,In_557);
nand U318 (N_318,In_1676,In_1002);
or U319 (N_319,In_196,In_170);
nor U320 (N_320,In_471,In_999);
nand U321 (N_321,In_1084,In_330);
nor U322 (N_322,In_647,In_929);
nor U323 (N_323,In_623,In_424);
or U324 (N_324,In_1706,In_1759);
or U325 (N_325,In_800,In_544);
nor U326 (N_326,In_587,In_496);
or U327 (N_327,In_333,In_84);
nor U328 (N_328,In_1405,In_1951);
nor U329 (N_329,In_925,In_1700);
and U330 (N_330,In_1474,In_659);
nand U331 (N_331,In_293,In_1778);
nand U332 (N_332,In_1744,In_287);
and U333 (N_333,In_1367,In_1928);
nand U334 (N_334,In_1503,In_1588);
nand U335 (N_335,In_1388,In_1751);
nand U336 (N_336,In_1237,In_1151);
and U337 (N_337,In_144,In_449);
nor U338 (N_338,In_1370,In_1833);
nor U339 (N_339,In_468,In_578);
xnor U340 (N_340,In_1461,In_256);
nand U341 (N_341,In_55,In_1978);
nand U342 (N_342,In_1350,In_649);
xor U343 (N_343,In_627,In_1022);
or U344 (N_344,In_1507,In_1709);
xnor U345 (N_345,In_11,In_812);
and U346 (N_346,In_1196,In_1332);
and U347 (N_347,In_1998,In_1704);
or U348 (N_348,In_722,In_629);
nand U349 (N_349,In_1584,In_1729);
and U350 (N_350,In_70,In_429);
nor U351 (N_351,In_227,In_1654);
or U352 (N_352,In_1862,In_1659);
and U353 (N_353,In_869,In_625);
and U354 (N_354,In_1912,In_226);
nand U355 (N_355,In_897,In_1240);
nor U356 (N_356,In_1733,In_1213);
xor U357 (N_357,In_234,In_255);
and U358 (N_358,In_852,In_1559);
or U359 (N_359,In_1795,In_1045);
nor U360 (N_360,In_1997,In_1864);
and U361 (N_361,In_710,In_62);
nand U362 (N_362,In_495,In_1544);
and U363 (N_363,In_1026,In_317);
nor U364 (N_364,In_1297,In_79);
nand U365 (N_365,In_715,In_394);
nand U366 (N_366,In_941,In_1060);
nor U367 (N_367,In_210,In_1737);
or U368 (N_368,In_511,In_59);
nor U369 (N_369,In_1721,In_173);
xnor U370 (N_370,In_72,In_1621);
nand U371 (N_371,In_726,In_1333);
and U372 (N_372,In_414,In_1552);
and U373 (N_373,In_521,In_1336);
and U374 (N_374,In_69,In_1574);
nand U375 (N_375,In_1980,In_984);
nor U376 (N_376,In_976,In_100);
and U377 (N_377,In_1752,In_874);
xnor U378 (N_378,In_1994,In_65);
nand U379 (N_379,In_143,In_1920);
and U380 (N_380,In_1774,In_1484);
xnor U381 (N_381,In_357,In_713);
or U382 (N_382,In_596,In_1890);
nor U383 (N_383,In_888,In_677);
nand U384 (N_384,In_591,In_1749);
or U385 (N_385,In_434,In_1454);
and U386 (N_386,In_387,In_168);
nand U387 (N_387,In_1323,In_1878);
and U388 (N_388,In_474,In_41);
nand U389 (N_389,In_961,In_1152);
or U390 (N_390,In_478,In_711);
nor U391 (N_391,In_566,In_954);
xor U392 (N_392,In_942,In_1166);
nor U393 (N_393,In_835,In_700);
nand U394 (N_394,In_1187,In_507);
xnor U395 (N_395,In_608,In_1478);
xnor U396 (N_396,In_1655,In_127);
nor U397 (N_397,In_598,In_188);
and U398 (N_398,In_292,In_1785);
and U399 (N_399,In_366,In_917);
nand U400 (N_400,In_297,In_1791);
nand U401 (N_401,In_1710,In_927);
or U402 (N_402,In_786,In_1611);
xor U403 (N_403,In_1549,In_375);
nor U404 (N_404,In_553,In_1345);
xor U405 (N_405,In_1748,In_879);
xor U406 (N_406,In_599,In_1142);
and U407 (N_407,In_1538,In_1712);
xnor U408 (N_408,In_252,In_242);
and U409 (N_409,In_308,In_907);
nand U410 (N_410,In_1126,In_134);
nor U411 (N_411,In_1811,In_948);
or U412 (N_412,In_1841,In_1280);
nand U413 (N_413,In_1844,In_1042);
and U414 (N_414,In_438,In_182);
xor U415 (N_415,In_1494,In_1794);
nand U416 (N_416,In_1073,In_1595);
nor U417 (N_417,In_274,In_1372);
or U418 (N_418,In_1952,In_493);
nand U419 (N_419,In_780,In_459);
nand U420 (N_420,In_646,In_1964);
nor U421 (N_421,In_218,In_1466);
nand U422 (N_422,In_1820,In_1346);
xnor U423 (N_423,In_975,In_898);
and U424 (N_424,In_425,In_1486);
xor U425 (N_425,In_845,In_757);
or U426 (N_426,In_405,In_586);
and U427 (N_427,In_386,In_1352);
xnor U428 (N_428,In_1051,In_1074);
and U429 (N_429,In_1129,In_164);
nor U430 (N_430,In_1446,In_1518);
xor U431 (N_431,In_319,In_1690);
nor U432 (N_432,In_148,In_1810);
nor U433 (N_433,In_643,In_1031);
xor U434 (N_434,In_1261,In_323);
nor U435 (N_435,In_1059,In_126);
or U436 (N_436,In_1941,In_315);
and U437 (N_437,In_1805,In_1101);
xnor U438 (N_438,In_1673,In_727);
nor U439 (N_439,In_1296,In_705);
nand U440 (N_440,In_806,In_1585);
or U441 (N_441,In_1419,In_1433);
and U442 (N_442,In_368,In_559);
nor U443 (N_443,In_1036,In_230);
or U444 (N_444,In_1449,In_1167);
and U445 (N_445,In_1271,In_150);
xor U446 (N_446,In_1732,In_1343);
xnor U447 (N_447,In_432,In_1492);
xnor U448 (N_448,In_1974,In_561);
or U449 (N_449,In_92,In_1006);
and U450 (N_450,In_363,In_1291);
or U451 (N_451,In_974,In_300);
or U452 (N_452,In_327,In_827);
or U453 (N_453,In_1757,In_636);
or U454 (N_454,In_130,In_1831);
or U455 (N_455,In_1198,In_1725);
xnor U456 (N_456,In_630,In_161);
xnor U457 (N_457,In_1312,In_435);
nand U458 (N_458,In_125,In_1702);
and U459 (N_459,In_1502,In_953);
nor U460 (N_460,In_1190,In_1093);
and U461 (N_461,In_1948,In_1403);
or U462 (N_462,In_1547,In_990);
or U463 (N_463,In_683,In_1908);
and U464 (N_464,In_1414,In_966);
and U465 (N_465,In_746,In_785);
and U466 (N_466,In_1935,In_667);
and U467 (N_467,In_1736,In_1513);
xor U468 (N_468,In_844,In_909);
or U469 (N_469,In_1726,In_448);
nor U470 (N_470,In_774,In_141);
nand U471 (N_471,In_583,In_1604);
and U472 (N_472,In_1524,In_1287);
and U473 (N_473,In_840,In_1764);
nand U474 (N_474,In_826,In_1975);
and U475 (N_475,In_34,In_1992);
nand U476 (N_476,In_1344,In_1410);
nor U477 (N_477,In_1272,In_378);
nor U478 (N_478,In_1080,In_959);
or U479 (N_479,In_1775,In_1378);
xor U480 (N_480,In_204,In_1807);
and U481 (N_481,In_470,In_894);
and U482 (N_482,In_520,In_1085);
nor U483 (N_483,In_676,In_1379);
xor U484 (N_484,In_1493,In_1122);
nand U485 (N_485,In_794,In_258);
nor U486 (N_486,In_1593,In_1417);
nor U487 (N_487,In_494,In_1892);
and U488 (N_488,In_121,In_406);
xor U489 (N_489,In_522,In_809);
nand U490 (N_490,In_481,In_1863);
or U491 (N_491,In_1035,In_1895);
nor U492 (N_492,In_1781,In_1644);
or U493 (N_493,In_1292,In_1731);
or U494 (N_494,In_1229,In_1698);
or U495 (N_495,In_600,In_1962);
xor U496 (N_496,In_1157,In_1531);
nor U497 (N_497,In_349,In_1536);
xor U498 (N_498,In_213,In_497);
nand U499 (N_499,In_1251,In_1958);
and U500 (N_500,In_1851,In_577);
nor U501 (N_501,In_286,In_875);
xnor U502 (N_502,In_27,In_1943);
nand U503 (N_503,In_1707,In_1854);
nand U504 (N_504,In_98,In_517);
xnor U505 (N_505,In_1498,In_848);
xnor U506 (N_506,In_871,In_782);
nor U507 (N_507,In_1681,In_837);
and U508 (N_508,In_219,In_1061);
or U509 (N_509,In_603,In_687);
or U510 (N_510,In_743,In_1509);
nand U511 (N_511,In_526,In_246);
and U512 (N_512,In_503,In_965);
nor U513 (N_513,In_1515,In_166);
xnor U514 (N_514,In_590,In_988);
xor U515 (N_515,In_1207,In_1885);
and U516 (N_516,In_393,In_1910);
xor U517 (N_517,In_915,In_1944);
xnor U518 (N_518,In_74,In_1718);
nand U519 (N_519,In_1628,In_1338);
or U520 (N_520,In_550,In_842);
and U521 (N_521,In_762,In_1421);
or U522 (N_522,In_1806,In_1848);
or U523 (N_523,In_1428,In_1476);
and U524 (N_524,In_1102,In_525);
or U525 (N_525,In_1893,In_720);
or U526 (N_526,In_1104,In_1753);
nor U527 (N_527,In_248,In_547);
nor U528 (N_528,In_796,In_1387);
nand U529 (N_529,In_1247,In_1459);
and U530 (N_530,In_1159,In_1564);
or U531 (N_531,In_208,In_957);
nand U532 (N_532,In_340,In_1821);
nand U533 (N_533,In_1439,In_1264);
xnor U534 (N_534,In_1216,In_1222);
nor U535 (N_535,In_58,In_192);
nand U536 (N_536,In_1301,In_1669);
or U537 (N_537,In_607,In_1098);
or U538 (N_538,In_236,In_651);
nor U539 (N_539,In_680,In_1165);
xor U540 (N_540,In_310,In_1041);
nand U541 (N_541,In_1808,In_777);
or U542 (N_542,In_477,In_335);
xnor U543 (N_543,In_174,In_932);
or U544 (N_544,In_365,In_1715);
or U545 (N_545,In_1537,In_554);
xnor U546 (N_546,In_367,In_568);
and U547 (N_547,In_250,In_819);
or U548 (N_548,In_402,In_978);
or U549 (N_549,In_950,In_979);
nand U550 (N_550,In_444,In_136);
xor U551 (N_551,In_1268,In_889);
or U552 (N_552,In_1548,In_1406);
nand U553 (N_553,In_773,In_1723);
or U554 (N_554,In_1720,In_1796);
nor U555 (N_555,In_515,In_1936);
and U556 (N_556,In_12,In_865);
xor U557 (N_557,In_1110,In_1488);
or U558 (N_558,In_220,In_318);
nand U559 (N_559,In_1929,In_1527);
or U560 (N_560,In_433,In_1620);
and U561 (N_561,In_247,In_912);
nor U562 (N_562,In_42,In_1746);
and U563 (N_563,In_790,In_1598);
or U564 (N_564,In_267,In_1314);
xnor U565 (N_565,In_655,In_268);
nand U566 (N_566,In_499,In_1320);
xnor U567 (N_567,In_104,In_754);
nand U568 (N_568,In_1896,In_1981);
nand U569 (N_569,In_1813,In_1156);
xnor U570 (N_570,In_1075,In_1888);
or U571 (N_571,In_299,In_1377);
nand U572 (N_572,In_1221,In_648);
or U573 (N_573,In_825,In_154);
xor U574 (N_574,In_716,In_1248);
nor U575 (N_575,In_277,In_224);
or U576 (N_576,In_717,In_699);
xor U577 (N_577,In_1274,In_857);
or U578 (N_578,In_231,In_1422);
and U579 (N_579,In_1784,In_1685);
xor U580 (N_580,In_1689,In_1989);
xnor U581 (N_581,In_1973,In_50);
or U582 (N_582,In_1032,In_1381);
and U583 (N_583,In_25,In_228);
nor U584 (N_584,In_1747,In_1290);
xor U585 (N_585,In_26,In_678);
nand U586 (N_586,In_1143,In_1231);
or U587 (N_587,In_1651,In_1193);
or U588 (N_588,In_1632,In_1458);
nor U589 (N_589,In_1612,In_372);
nand U590 (N_590,In_91,In_1714);
xor U591 (N_591,In_1115,In_1678);
nand U592 (N_592,In_731,In_1249);
xor U593 (N_593,In_253,In_1897);
nand U594 (N_594,In_1900,In_1602);
or U595 (N_595,In_249,In_1675);
xor U596 (N_596,In_201,In_1730);
and U597 (N_597,In_1354,In_80);
and U598 (N_598,In_991,In_1546);
nor U599 (N_599,In_1383,In_1362);
nand U600 (N_600,In_1471,In_215);
or U601 (N_601,In_518,In_1541);
and U602 (N_602,In_779,In_232);
nor U603 (N_603,In_549,In_851);
nand U604 (N_604,In_1572,In_147);
nand U605 (N_605,In_582,In_1232);
nand U606 (N_606,In_886,In_1610);
or U607 (N_607,In_1849,In_905);
and U608 (N_608,In_1078,In_1284);
nor U609 (N_609,In_682,In_1315);
nor U610 (N_610,In_1455,In_924);
and U611 (N_611,In_1431,In_416);
xnor U612 (N_612,In_1497,In_263);
and U613 (N_613,In_691,In_71);
nor U614 (N_614,In_947,In_922);
xor U615 (N_615,In_83,In_1226);
or U616 (N_616,In_1375,In_1576);
or U617 (N_617,In_1857,In_1797);
nand U618 (N_618,In_1798,In_56);
xnor U619 (N_619,In_1342,In_1970);
nand U620 (N_620,In_391,In_632);
xnor U621 (N_621,In_383,In_346);
nor U622 (N_622,In_1606,In_930);
and U623 (N_623,In_928,In_1647);
and U624 (N_624,In_1907,In_1083);
xnor U625 (N_625,In_418,In_1930);
xnor U626 (N_626,In_831,In_442);
nand U627 (N_627,In_466,In_1329);
or U628 (N_628,In_541,In_380);
nor U629 (N_629,In_172,In_328);
nand U630 (N_630,In_1724,In_1947);
or U631 (N_631,In_1823,In_1553);
nor U632 (N_632,In_1209,In_1853);
and U633 (N_633,In_993,In_76);
and U634 (N_634,In_931,In_1306);
nand U635 (N_635,In_1153,In_229);
or U636 (N_636,In_1111,In_309);
nand U637 (N_637,In_162,In_958);
and U638 (N_638,In_33,In_622);
xor U639 (N_639,In_1348,In_1898);
nor U640 (N_640,In_1542,In_1062);
nor U641 (N_641,In_457,In_570);
xor U642 (N_642,In_896,In_1136);
xor U643 (N_643,In_1456,In_32);
or U644 (N_644,In_689,In_1302);
or U645 (N_645,In_900,In_658);
nand U646 (N_646,In_1694,In_565);
xnor U647 (N_647,In_787,In_463);
xor U648 (N_648,In_61,In_1162);
nand U649 (N_649,In_163,In_1734);
and U650 (N_650,In_1591,In_1341);
nand U651 (N_651,In_1535,In_995);
and U652 (N_652,In_1412,In_1955);
nor U653 (N_653,In_364,In_1824);
or U654 (N_654,In_934,In_1648);
nand U655 (N_655,In_1745,In_54);
xor U656 (N_656,In_1750,In_1132);
xnor U657 (N_657,In_1817,In_1259);
nor U658 (N_658,In_597,In_1114);
and U659 (N_659,In_455,In_967);
or U660 (N_660,In_624,In_1766);
nand U661 (N_661,In_1183,In_498);
nand U662 (N_662,In_384,In_1330);
nand U663 (N_663,In_1452,In_1703);
nor U664 (N_664,In_288,In_1915);
nor U665 (N_665,In_1925,In_401);
and U666 (N_666,In_1762,In_666);
and U667 (N_667,In_1569,In_1077);
nor U668 (N_668,In_1783,In_1465);
nand U669 (N_669,In_1112,In_920);
xor U670 (N_670,In_1692,In_891);
xnor U671 (N_671,In_1802,In_751);
and U672 (N_672,In_152,In_1158);
and U673 (N_673,In_1969,In_533);
or U674 (N_674,In_1708,In_68);
xnor U675 (N_675,In_362,In_171);
xnor U676 (N_676,In_569,In_1234);
nor U677 (N_677,In_721,In_1573);
nor U678 (N_678,In_151,In_5);
or U679 (N_679,In_379,In_536);
nand U680 (N_680,In_1954,In_28);
nand U681 (N_681,In_1525,In_1579);
and U682 (N_682,In_694,In_1294);
or U683 (N_683,In_1179,In_529);
or U684 (N_684,In_1613,In_1066);
or U685 (N_685,In_1687,In_473);
and U686 (N_686,In_1163,In_1967);
nor U687 (N_687,In_458,In_52);
nand U688 (N_688,In_97,In_1514);
and U689 (N_689,In_298,In_1919);
nand U690 (N_690,In_1519,In_1761);
nand U691 (N_691,In_501,In_119);
nor U692 (N_692,In_986,In_604);
or U693 (N_693,In_1971,In_1368);
nand U694 (N_694,In_1622,In_969);
or U695 (N_695,In_1470,In_1587);
nor U696 (N_696,In_1086,In_1804);
or U697 (N_697,In_1119,In_706);
or U698 (N_698,In_1369,In_702);
xnor U699 (N_699,In_1568,In_1217);
nor U700 (N_700,In_1220,In_1942);
xor U701 (N_701,In_1697,In_1635);
or U702 (N_702,In_422,In_1859);
nor U703 (N_703,In_1865,In_1516);
nor U704 (N_704,In_39,In_1837);
nor U705 (N_705,In_792,In_212);
nand U706 (N_706,In_107,In_1436);
xnor U707 (N_707,In_732,In_1828);
nand U708 (N_708,In_95,In_1532);
xor U709 (N_709,In_1281,In_1090);
nor U710 (N_710,In_1899,In_750);
nor U711 (N_711,In_187,In_919);
nand U712 (N_712,In_873,In_1154);
or U713 (N_713,In_1739,In_36);
or U714 (N_714,In_1852,In_884);
and U715 (N_715,In_1118,In_530);
or U716 (N_716,In_1138,In_1977);
or U717 (N_717,In_595,In_1671);
xnor U718 (N_718,In_1262,In_707);
xnor U719 (N_719,In_479,In_1228);
nand U720 (N_720,In_329,In_279);
xor U721 (N_721,In_1551,In_1662);
and U722 (N_722,In_564,In_830);
nor U723 (N_723,In_1087,In_688);
xnor U724 (N_724,In_1842,In_1279);
nand U725 (N_725,In_903,In_452);
and U726 (N_726,In_339,In_303);
and U727 (N_727,In_1850,In_1608);
nand U728 (N_728,In_1360,In_0);
nor U729 (N_729,In_1014,In_1363);
or U730 (N_730,In_935,In_1174);
or U731 (N_731,In_1239,In_1530);
nand U732 (N_732,In_1902,In_467);
nand U733 (N_733,In_1416,In_1617);
and U734 (N_734,In_1276,In_1904);
nor U735 (N_735,In_1049,In_488);
nor U736 (N_736,In_16,In_1634);
nand U737 (N_737,In_1882,In_539);
nand U738 (N_738,In_1887,In_951);
xor U739 (N_739,In_1177,In_1555);
or U740 (N_740,In_1953,In_51);
nor U741 (N_741,In_613,In_970);
and U742 (N_742,In_805,In_1095);
nand U743 (N_743,In_165,In_781);
and U744 (N_744,In_1691,In_120);
nand U745 (N_745,In_1155,In_356);
and U746 (N_746,In_265,In_1779);
or U747 (N_747,In_112,In_1464);
nor U748 (N_748,In_952,In_788);
or U749 (N_749,In_1520,In_403);
or U750 (N_750,In_609,In_1298);
nand U751 (N_751,In_167,In_1295);
xnor U752 (N_752,In_1144,In_1283);
nand U753 (N_753,In_1140,In_558);
xnor U754 (N_754,In_914,In_451);
and U755 (N_755,In_1339,In_133);
nand U756 (N_756,In_1011,In_1858);
nor U757 (N_757,In_1308,In_1212);
nor U758 (N_758,In_1255,In_443);
nor U759 (N_759,In_373,In_1963);
nor U760 (N_760,In_739,In_469);
xor U761 (N_761,In_2,In_1586);
nor U762 (N_762,In_1125,In_440);
or U763 (N_763,In_1068,In_110);
xor U764 (N_764,In_644,In_1601);
and U765 (N_765,In_1103,In_1260);
or U766 (N_766,In_343,In_1398);
nor U767 (N_767,In_1875,In_1965);
xor U768 (N_768,In_355,In_664);
nor U769 (N_769,In_1960,In_456);
and U770 (N_770,In_1460,In_24);
xnor U771 (N_771,In_1743,In_619);
nand U772 (N_772,In_1208,In_1358);
and U773 (N_773,In_1664,In_1392);
and U774 (N_774,In_735,In_1512);
xnor U775 (N_775,In_1425,In_589);
and U776 (N_776,In_1558,In_1475);
xor U777 (N_777,In_257,In_1192);
xor U778 (N_778,In_431,In_877);
xor U779 (N_779,In_537,In_1533);
or U780 (N_780,In_1082,In_1918);
or U781 (N_781,In_798,In_1713);
nand U782 (N_782,In_1236,In_1018);
nor U783 (N_783,In_641,In_1242);
nand U784 (N_784,In_272,In_1822);
and U785 (N_785,In_1760,In_1631);
nand U786 (N_786,In_399,In_1010);
nand U787 (N_787,In_867,In_464);
or U788 (N_788,In_1860,In_1263);
xnor U789 (N_789,In_1097,In_818);
or U790 (N_790,In_532,In_1238);
or U791 (N_791,In_43,In_316);
xnor U792 (N_792,In_1319,In_491);
nand U793 (N_793,In_747,In_241);
nand U794 (N_794,In_460,In_737);
or U795 (N_795,In_506,In_1517);
nor U796 (N_796,In_744,In_271);
or U797 (N_797,In_155,In_38);
nor U798 (N_798,In_360,In_1670);
and U799 (N_799,In_510,In_1792);
xnor U800 (N_800,In_1683,In_441);
or U801 (N_801,In_1096,In_280);
and U802 (N_802,In_1311,In_1434);
nor U803 (N_803,In_1175,In_1534);
xor U804 (N_804,In_1223,In_1638);
xor U805 (N_805,In_936,In_500);
xnor U806 (N_806,In_1999,In_736);
nand U807 (N_807,In_783,In_793);
and U808 (N_808,In_21,In_419);
nand U809 (N_809,In_1218,In_1423);
or U810 (N_810,In_396,In_684);
nand U811 (N_811,In_881,In_516);
and U812 (N_812,In_175,In_759);
nor U813 (N_813,In_1374,In_1754);
nand U814 (N_814,In_180,In_1856);
nor U815 (N_815,In_1325,In_1224);
nand U816 (N_816,In_186,In_113);
xor U817 (N_817,In_1257,In_122);
or U818 (N_818,In_1215,In_669);
xnor U819 (N_819,In_1901,In_1241);
or U820 (N_820,In_1560,In_1990);
and U821 (N_821,In_1340,In_738);
or U822 (N_822,In_266,In_1914);
xnor U823 (N_823,In_1646,In_1641);
nand U824 (N_824,In_1996,In_1578);
or U825 (N_825,In_841,In_1609);
nor U826 (N_826,In_1686,In_326);
nor U827 (N_827,In_198,In_37);
xor U828 (N_828,In_295,In_592);
or U829 (N_829,In_512,In_1044);
xnor U830 (N_830,In_656,In_836);
nor U831 (N_831,In_908,In_85);
or U832 (N_832,In_670,In_1834);
nand U833 (N_833,In_772,In_1303);
nor U834 (N_834,In_673,In_1931);
nand U835 (N_835,In_1677,In_823);
or U836 (N_836,In_1511,In_527);
and U837 (N_837,In_724,In_1021);
xor U838 (N_838,In_1767,In_1660);
nor U839 (N_839,In_602,In_1230);
and U840 (N_840,In_972,In_803);
xor U841 (N_841,In_1113,In_1016);
nand U842 (N_842,In_359,In_178);
xor U843 (N_843,In_808,In_15);
xnor U844 (N_844,In_1131,In_1254);
or U845 (N_845,In_1030,In_1012);
nand U846 (N_846,In_206,In_203);
nand U847 (N_847,In_849,In_337);
or U848 (N_848,In_887,In_1128);
and U849 (N_849,In_450,In_1491);
xor U850 (N_850,In_1397,In_610);
or U851 (N_851,In_1300,In_1583);
nand U852 (N_852,In_1133,In_505);
xor U853 (N_853,In_149,In_1181);
and U854 (N_854,In_1137,In_1968);
nor U855 (N_855,In_311,In_1384);
or U856 (N_856,In_755,In_1508);
nor U857 (N_857,In_307,In_1554);
or U858 (N_858,In_1027,In_14);
nor U859 (N_859,In_428,In_758);
or U860 (N_860,In_81,In_1793);
or U861 (N_861,In_1099,In_1293);
xnor U862 (N_862,In_22,In_977);
nand U863 (N_863,In_797,In_1717);
and U864 (N_864,In_205,In_767);
and U865 (N_865,In_1819,In_686);
xor U866 (N_866,In_513,In_1581);
nor U867 (N_867,In_1966,In_634);
or U868 (N_868,In_556,In_1201);
xor U869 (N_869,In_581,In_436);
xnor U870 (N_870,In_1845,In_1321);
nor U871 (N_871,In_1543,In_334);
and U872 (N_872,In_376,In_714);
nand U873 (N_873,In_870,In_701);
nand U874 (N_874,In_789,In_892);
and U875 (N_875,In_1580,In_860);
or U876 (N_876,In_158,In_901);
or U877 (N_877,In_652,In_1070);
xor U878 (N_878,In_1328,In_810);
and U879 (N_879,In_937,In_563);
and U880 (N_880,In_906,In_1173);
nor U881 (N_881,In_801,In_259);
and U882 (N_882,In_1809,In_1589);
nor U883 (N_883,In_594,In_1665);
or U884 (N_884,In_1800,In_853);
or U885 (N_885,In_411,In_238);
nand U886 (N_886,In_57,In_1500);
nor U887 (N_887,In_1872,In_828);
xnor U888 (N_888,In_1182,In_44);
nor U889 (N_889,In_956,In_895);
nor U890 (N_890,In_454,In_1365);
xnor U891 (N_891,In_31,In_1504);
or U892 (N_892,In_996,In_885);
nand U893 (N_893,In_575,In_1983);
xor U894 (N_894,In_1877,In_1289);
nor U895 (N_895,In_1505,In_1866);
and U896 (N_896,In_579,In_862);
xor U897 (N_897,In_377,In_1619);
nor U898 (N_898,In_82,In_1666);
or U899 (N_899,In_723,In_1776);
nor U900 (N_900,In_1451,In_771);
and U901 (N_901,In_60,In_1304);
nor U902 (N_902,In_1597,In_748);
nand U903 (N_903,In_445,In_1880);
or U904 (N_904,In_1869,In_1065);
or U905 (N_905,In_64,In_768);
nand U906 (N_906,In_1415,In_1313);
nand U907 (N_907,In_1483,In_1437);
and U908 (N_908,In_807,In_963);
or U909 (N_909,In_1763,In_1123);
nand U910 (N_910,In_1940,In_761);
and U911 (N_911,In_733,In_621);
nand U912 (N_912,In_1039,In_465);
nand U913 (N_913,In_1886,In_1479);
or U914 (N_914,In_353,In_1092);
or U915 (N_915,In_115,In_1202);
nand U916 (N_916,In_1490,In_395);
or U917 (N_917,In_1688,In_1038);
xnor U918 (N_918,In_1873,In_939);
xnor U919 (N_919,In_382,In_1874);
nand U920 (N_920,In_1636,In_1418);
xnor U921 (N_921,In_159,In_381);
or U922 (N_922,In_332,In_294);
xnor U923 (N_923,In_1826,In_657);
or U924 (N_924,In_336,In_1253);
xor U925 (N_925,In_486,In_776);
xor U926 (N_926,In_1922,In_275);
xnor U927 (N_927,In_1501,In_1364);
nor U928 (N_928,In_1679,In_618);
xnor U929 (N_929,In_614,In_1528);
xor U930 (N_930,In_358,In_1523);
xnor U931 (N_931,In_412,In_128);
or U932 (N_932,In_1995,In_1322);
xnor U933 (N_933,In_49,In_9);
or U934 (N_934,In_195,In_1040);
nand U935 (N_935,In_1172,In_94);
xor U936 (N_936,In_545,In_1435);
and U937 (N_937,In_1550,In_183);
and U938 (N_938,In_417,In_1772);
and U939 (N_939,In_1566,In_548);
xnor U940 (N_940,In_1393,In_1891);
or U941 (N_941,In_1765,In_858);
and U942 (N_942,In_665,In_763);
xnor U943 (N_943,In_695,In_285);
or U944 (N_944,In_940,In_222);
or U945 (N_945,In_193,In_1057);
xor U946 (N_946,In_626,In_660);
nor U947 (N_947,In_243,In_654);
or U948 (N_948,In_528,In_200);
or U949 (N_949,In_1699,In_854);
and U950 (N_950,In_1299,In_1840);
or U951 (N_951,In_1993,In_576);
and U952 (N_952,In_1063,In_1653);
or U953 (N_953,In_1539,In_663);
or U954 (N_954,In_1127,In_1871);
nor U955 (N_955,In_132,In_616);
xnor U956 (N_956,In_1661,In_415);
and U957 (N_957,In_753,In_962);
nand U958 (N_958,In_1556,In_8);
nor U959 (N_959,In_341,In_1562);
and U960 (N_960,In_821,In_1349);
xnor U961 (N_961,In_987,In_1596);
nand U962 (N_962,In_1432,In_1424);
and U963 (N_963,In_1567,In_645);
or U964 (N_964,In_741,In_1161);
or U965 (N_965,In_116,In_1402);
or U966 (N_966,In_145,In_1327);
xor U967 (N_967,In_1386,In_389);
and U968 (N_968,In_1134,In_1278);
nand U969 (N_969,In_7,In_1400);
and U970 (N_970,In_573,In_1141);
and U971 (N_971,In_1643,In_338);
nand U972 (N_972,In_278,In_1441);
or U973 (N_973,In_447,In_1790);
nand U974 (N_974,In_140,In_1861);
nor U975 (N_975,In_105,In_87);
and U976 (N_976,In_543,In_1642);
and U977 (N_977,In_385,In_1529);
xnor U978 (N_978,In_1148,In_1053);
and U979 (N_979,In_799,In_981);
or U980 (N_980,In_1351,In_1185);
xor U981 (N_981,In_1984,In_1194);
nor U982 (N_982,In_784,In_73);
xor U983 (N_983,In_923,In_1916);
nor U984 (N_984,In_650,In_1883);
nor U985 (N_985,In_1624,In_476);
nand U986 (N_986,In_124,In_982);
and U987 (N_987,In_261,In_1135);
and U988 (N_988,In_1335,In_306);
xor U989 (N_989,In_6,In_1592);
nand U990 (N_990,In_872,In_679);
xnor U991 (N_991,In_93,In_289);
nand U992 (N_992,In_427,In_1801);
or U993 (N_993,In_1005,In_1945);
nor U994 (N_994,In_1847,In_1106);
nand U995 (N_995,In_1693,In_18);
xor U996 (N_996,In_1839,In_484);
or U997 (N_997,In_968,In_1577);
nor U998 (N_998,In_1680,In_1870);
nand U999 (N_999,In_420,In_352);
and U1000 (N_1000,N_979,N_778);
or U1001 (N_1001,N_493,N_460);
and U1002 (N_1002,N_264,N_513);
nand U1003 (N_1003,N_422,N_914);
nand U1004 (N_1004,N_93,N_94);
and U1005 (N_1005,N_964,N_705);
nor U1006 (N_1006,N_576,N_865);
nor U1007 (N_1007,N_52,N_282);
or U1008 (N_1008,N_90,N_198);
and U1009 (N_1009,N_251,N_389);
nand U1010 (N_1010,N_306,N_845);
nor U1011 (N_1011,N_445,N_428);
nand U1012 (N_1012,N_372,N_215);
xor U1013 (N_1013,N_167,N_483);
xnor U1014 (N_1014,N_492,N_578);
xor U1015 (N_1015,N_788,N_846);
and U1016 (N_1016,N_47,N_785);
nand U1017 (N_1017,N_606,N_337);
and U1018 (N_1018,N_291,N_388);
nor U1019 (N_1019,N_943,N_512);
or U1020 (N_1020,N_43,N_396);
and U1021 (N_1021,N_408,N_987);
xor U1022 (N_1022,N_6,N_640);
nor U1023 (N_1023,N_991,N_590);
nand U1024 (N_1024,N_104,N_234);
xor U1025 (N_1025,N_651,N_83);
nand U1026 (N_1026,N_133,N_536);
nor U1027 (N_1027,N_541,N_848);
nor U1028 (N_1028,N_325,N_581);
or U1029 (N_1029,N_672,N_294);
xnor U1030 (N_1030,N_745,N_89);
nand U1031 (N_1031,N_711,N_270);
and U1032 (N_1032,N_718,N_447);
nor U1033 (N_1033,N_1,N_425);
or U1034 (N_1034,N_28,N_277);
nand U1035 (N_1035,N_164,N_438);
and U1036 (N_1036,N_456,N_201);
and U1037 (N_1037,N_615,N_176);
xor U1038 (N_1038,N_693,N_764);
nor U1039 (N_1039,N_310,N_111);
nand U1040 (N_1040,N_811,N_508);
or U1041 (N_1041,N_161,N_582);
and U1042 (N_1042,N_65,N_527);
nor U1043 (N_1043,N_947,N_91);
and U1044 (N_1044,N_165,N_714);
nand U1045 (N_1045,N_568,N_468);
nand U1046 (N_1046,N_398,N_222);
xnor U1047 (N_1047,N_269,N_548);
nor U1048 (N_1048,N_765,N_95);
xor U1049 (N_1049,N_860,N_108);
and U1050 (N_1050,N_587,N_669);
or U1051 (N_1051,N_287,N_800);
nand U1052 (N_1052,N_480,N_288);
nand U1053 (N_1053,N_96,N_376);
and U1054 (N_1054,N_427,N_815);
xnor U1055 (N_1055,N_982,N_183);
or U1056 (N_1056,N_78,N_175);
nand U1057 (N_1057,N_791,N_908);
or U1058 (N_1058,N_974,N_442);
xnor U1059 (N_1059,N_97,N_35);
xnor U1060 (N_1060,N_851,N_237);
nor U1061 (N_1061,N_132,N_598);
nand U1062 (N_1062,N_965,N_329);
or U1063 (N_1063,N_944,N_896);
or U1064 (N_1064,N_124,N_595);
nand U1065 (N_1065,N_546,N_904);
and U1066 (N_1066,N_743,N_903);
nor U1067 (N_1067,N_448,N_603);
nor U1068 (N_1068,N_289,N_967);
nor U1069 (N_1069,N_935,N_121);
or U1070 (N_1070,N_881,N_430);
and U1071 (N_1071,N_510,N_457);
nand U1072 (N_1072,N_324,N_81);
and U1073 (N_1073,N_208,N_130);
and U1074 (N_1074,N_709,N_730);
and U1075 (N_1075,N_423,N_687);
and U1076 (N_1076,N_781,N_195);
nand U1077 (N_1077,N_411,N_638);
and U1078 (N_1078,N_7,N_763);
or U1079 (N_1079,N_283,N_112);
nor U1080 (N_1080,N_879,N_774);
nand U1081 (N_1081,N_117,N_88);
and U1082 (N_1082,N_679,N_464);
xnor U1083 (N_1083,N_959,N_140);
or U1084 (N_1084,N_857,N_924);
or U1085 (N_1085,N_362,N_761);
nand U1086 (N_1086,N_821,N_301);
nand U1087 (N_1087,N_627,N_917);
xor U1088 (N_1088,N_565,N_837);
nand U1089 (N_1089,N_70,N_534);
xnor U1090 (N_1090,N_690,N_487);
nor U1091 (N_1091,N_106,N_169);
nand U1092 (N_1092,N_713,N_542);
xor U1093 (N_1093,N_544,N_831);
nand U1094 (N_1094,N_953,N_549);
nor U1095 (N_1095,N_892,N_580);
or U1096 (N_1096,N_484,N_474);
nand U1097 (N_1097,N_911,N_424);
nor U1098 (N_1098,N_998,N_521);
nor U1099 (N_1099,N_12,N_62);
nand U1100 (N_1100,N_275,N_27);
nor U1101 (N_1101,N_537,N_725);
nor U1102 (N_1102,N_734,N_807);
nor U1103 (N_1103,N_179,N_993);
nor U1104 (N_1104,N_42,N_916);
nand U1105 (N_1105,N_401,N_387);
or U1106 (N_1106,N_212,N_503);
nor U1107 (N_1107,N_805,N_342);
or U1108 (N_1108,N_153,N_583);
nor U1109 (N_1109,N_671,N_359);
and U1110 (N_1110,N_790,N_824);
and U1111 (N_1111,N_796,N_962);
and U1112 (N_1112,N_748,N_789);
xnor U1113 (N_1113,N_685,N_999);
and U1114 (N_1114,N_902,N_73);
or U1115 (N_1115,N_566,N_557);
or U1116 (N_1116,N_189,N_375);
xor U1117 (N_1117,N_279,N_192);
or U1118 (N_1118,N_23,N_155);
xnor U1119 (N_1119,N_531,N_946);
nor U1120 (N_1120,N_631,N_225);
nand U1121 (N_1121,N_190,N_966);
nand U1122 (N_1122,N_381,N_120);
xnor U1123 (N_1123,N_86,N_514);
or U1124 (N_1124,N_773,N_56);
and U1125 (N_1125,N_4,N_769);
xnor U1126 (N_1126,N_741,N_303);
or U1127 (N_1127,N_654,N_639);
and U1128 (N_1128,N_658,N_731);
nand U1129 (N_1129,N_650,N_775);
nand U1130 (N_1130,N_443,N_285);
and U1131 (N_1131,N_616,N_783);
xor U1132 (N_1132,N_641,N_613);
nor U1133 (N_1133,N_258,N_300);
and U1134 (N_1134,N_797,N_753);
xnor U1135 (N_1135,N_632,N_702);
xnor U1136 (N_1136,N_992,N_18);
or U1137 (N_1137,N_819,N_556);
xnor U1138 (N_1138,N_137,N_187);
and U1139 (N_1139,N_852,N_353);
nand U1140 (N_1140,N_662,N_202);
nand U1141 (N_1141,N_226,N_642);
nand U1142 (N_1142,N_913,N_437);
or U1143 (N_1143,N_333,N_945);
or U1144 (N_1144,N_171,N_382);
nand U1145 (N_1145,N_593,N_107);
or U1146 (N_1146,N_507,N_115);
xnor U1147 (N_1147,N_772,N_612);
and U1148 (N_1148,N_410,N_143);
nor U1149 (N_1149,N_216,N_957);
or U1150 (N_1150,N_838,N_569);
nor U1151 (N_1151,N_116,N_59);
nand U1152 (N_1152,N_900,N_77);
nand U1153 (N_1153,N_136,N_147);
or U1154 (N_1154,N_159,N_770);
and U1155 (N_1155,N_166,N_417);
nor U1156 (N_1156,N_610,N_496);
nor U1157 (N_1157,N_884,N_625);
nand U1158 (N_1158,N_379,N_304);
or U1159 (N_1159,N_439,N_470);
nor U1160 (N_1160,N_689,N_564);
or U1161 (N_1161,N_936,N_145);
or U1162 (N_1162,N_954,N_717);
xor U1163 (N_1163,N_758,N_491);
xnor U1164 (N_1164,N_604,N_204);
xor U1165 (N_1165,N_0,N_256);
xor U1166 (N_1166,N_82,N_971);
or U1167 (N_1167,N_346,N_69);
or U1168 (N_1168,N_330,N_281);
or U1169 (N_1169,N_706,N_795);
xor U1170 (N_1170,N_461,N_955);
xor U1171 (N_1171,N_901,N_397);
and U1172 (N_1172,N_859,N_485);
nor U1173 (N_1173,N_218,N_996);
xnor U1174 (N_1174,N_643,N_19);
nand U1175 (N_1175,N_682,N_877);
xnor U1176 (N_1176,N_539,N_554);
xor U1177 (N_1177,N_181,N_67);
or U1178 (N_1178,N_55,N_799);
nand U1179 (N_1179,N_343,N_828);
and U1180 (N_1180,N_421,N_605);
or U1181 (N_1181,N_888,N_697);
and U1182 (N_1182,N_61,N_691);
xnor U1183 (N_1183,N_871,N_313);
and U1184 (N_1184,N_400,N_332);
and U1185 (N_1185,N_928,N_316);
xnor U1186 (N_1186,N_280,N_298);
or U1187 (N_1187,N_191,N_688);
and U1188 (N_1188,N_453,N_829);
nor U1189 (N_1189,N_633,N_599);
and U1190 (N_1190,N_227,N_596);
and U1191 (N_1191,N_60,N_407);
nor U1192 (N_1192,N_634,N_926);
nor U1193 (N_1193,N_571,N_657);
and U1194 (N_1194,N_522,N_182);
nand U1195 (N_1195,N_168,N_645);
xnor U1196 (N_1196,N_668,N_247);
nor U1197 (N_1197,N_336,N_3);
nor U1198 (N_1198,N_648,N_245);
and U1199 (N_1199,N_868,N_273);
or U1200 (N_1200,N_498,N_296);
xnor U1201 (N_1201,N_572,N_980);
nand U1202 (N_1202,N_488,N_994);
and U1203 (N_1203,N_751,N_843);
or U1204 (N_1204,N_33,N_733);
nand U1205 (N_1205,N_114,N_494);
nand U1206 (N_1206,N_656,N_601);
nor U1207 (N_1207,N_715,N_894);
nor U1208 (N_1208,N_319,N_950);
nor U1209 (N_1209,N_738,N_463);
or U1210 (N_1210,N_579,N_525);
nor U1211 (N_1211,N_684,N_899);
xor U1212 (N_1212,N_479,N_38);
nor U1213 (N_1213,N_655,N_981);
and U1214 (N_1214,N_371,N_529);
and U1215 (N_1215,N_855,N_434);
or U1216 (N_1216,N_727,N_406);
nand U1217 (N_1217,N_213,N_197);
nand U1218 (N_1218,N_577,N_249);
or U1219 (N_1219,N_31,N_767);
nor U1220 (N_1220,N_497,N_158);
or U1221 (N_1221,N_261,N_762);
or U1222 (N_1222,N_162,N_482);
nor U1223 (N_1223,N_57,N_635);
or U1224 (N_1224,N_368,N_518);
xor U1225 (N_1225,N_649,N_150);
nor U1226 (N_1226,N_551,N_72);
nand U1227 (N_1227,N_873,N_808);
xnor U1228 (N_1228,N_813,N_412);
xor U1229 (N_1229,N_141,N_302);
nand U1230 (N_1230,N_351,N_87);
and U1231 (N_1231,N_874,N_490);
xnor U1232 (N_1232,N_708,N_110);
and U1233 (N_1233,N_320,N_784);
nand U1234 (N_1234,N_413,N_890);
nand U1235 (N_1235,N_624,N_547);
or U1236 (N_1236,N_930,N_870);
or U1237 (N_1237,N_779,N_918);
or U1238 (N_1238,N_937,N_698);
nand U1239 (N_1239,N_597,N_157);
and U1240 (N_1240,N_517,N_622);
nand U1241 (N_1241,N_887,N_128);
or U1242 (N_1242,N_348,N_794);
xnor U1243 (N_1243,N_895,N_76);
or U1244 (N_1244,N_36,N_502);
nand U1245 (N_1245,N_469,N_103);
or U1246 (N_1246,N_365,N_328);
nor U1247 (N_1247,N_100,N_126);
xor U1248 (N_1248,N_229,N_560);
nand U1249 (N_1249,N_630,N_976);
or U1250 (N_1250,N_17,N_205);
or U1251 (N_1251,N_520,N_653);
and U1252 (N_1252,N_472,N_252);
nor U1253 (N_1253,N_984,N_823);
nor U1254 (N_1254,N_370,N_308);
and U1255 (N_1255,N_575,N_739);
xor U1256 (N_1256,N_942,N_724);
nor U1257 (N_1257,N_803,N_321);
xnor U1258 (N_1258,N_265,N_312);
or U1259 (N_1259,N_737,N_98);
nor U1260 (N_1260,N_240,N_670);
nand U1261 (N_1261,N_809,N_259);
and U1262 (N_1262,N_403,N_969);
nand U1263 (N_1263,N_747,N_905);
xor U1264 (N_1264,N_501,N_804);
nor U1265 (N_1265,N_486,N_722);
and U1266 (N_1266,N_854,N_184);
and U1267 (N_1267,N_699,N_193);
nand U1268 (N_1268,N_864,N_125);
nand U1269 (N_1269,N_290,N_543);
nor U1270 (N_1270,N_552,N_466);
or U1271 (N_1271,N_680,N_210);
or U1272 (N_1272,N_263,N_151);
and U1273 (N_1273,N_146,N_678);
xnor U1274 (N_1274,N_573,N_465);
nor U1275 (N_1275,N_723,N_736);
xnor U1276 (N_1276,N_752,N_444);
nor U1277 (N_1277,N_390,N_34);
nand U1278 (N_1278,N_923,N_742);
or U1279 (N_1279,N_271,N_951);
nor U1280 (N_1280,N_886,N_891);
xor U1281 (N_1281,N_825,N_172);
xnor U1282 (N_1282,N_44,N_335);
nand U1283 (N_1283,N_677,N_39);
nor U1284 (N_1284,N_354,N_883);
nand U1285 (N_1285,N_500,N_611);
or U1286 (N_1286,N_710,N_449);
xor U1287 (N_1287,N_284,N_414);
nand U1288 (N_1288,N_667,N_200);
and U1289 (N_1289,N_949,N_822);
nand U1290 (N_1290,N_160,N_960);
and U1291 (N_1291,N_152,N_344);
and U1292 (N_1292,N_418,N_318);
nor U1293 (N_1293,N_415,N_455);
nand U1294 (N_1294,N_118,N_307);
xnor U1295 (N_1295,N_636,N_614);
and U1296 (N_1296,N_939,N_872);
xnor U1297 (N_1297,N_139,N_909);
or U1298 (N_1298,N_432,N_272);
nand U1299 (N_1299,N_626,N_801);
and U1300 (N_1300,N_459,N_473);
nor U1301 (N_1301,N_63,N_906);
xor U1302 (N_1302,N_694,N_760);
nand U1303 (N_1303,N_757,N_163);
or U1304 (N_1304,N_221,N_224);
nand U1305 (N_1305,N_637,N_833);
nand U1306 (N_1306,N_173,N_339);
xor U1307 (N_1307,N_239,N_102);
and U1308 (N_1308,N_749,N_58);
and U1309 (N_1309,N_921,N_454);
and U1310 (N_1310,N_602,N_948);
xnor U1311 (N_1311,N_985,N_207);
or U1312 (N_1312,N_24,N_910);
nand U1313 (N_1313,N_509,N_440);
nor U1314 (N_1314,N_41,N_740);
xor U1315 (N_1315,N_666,N_219);
xor U1316 (N_1316,N_334,N_681);
nor U1317 (N_1317,N_920,N_628);
xor U1318 (N_1318,N_9,N_374);
and U1319 (N_1319,N_322,N_853);
nor U1320 (N_1320,N_898,N_591);
nor U1321 (N_1321,N_814,N_253);
xor U1322 (N_1322,N_178,N_968);
nand U1323 (N_1323,N_471,N_360);
and U1324 (N_1324,N_402,N_609);
nand U1325 (N_1325,N_409,N_476);
nor U1326 (N_1326,N_478,N_732);
xor U1327 (N_1327,N_786,N_40);
and U1328 (N_1328,N_92,N_119);
and U1329 (N_1329,N_257,N_812);
and U1330 (N_1330,N_26,N_570);
or U1331 (N_1331,N_726,N_934);
nor U1332 (N_1332,N_878,N_350);
and U1333 (N_1333,N_506,N_882);
xor U1334 (N_1334,N_676,N_720);
nand U1335 (N_1335,N_391,N_806);
or U1336 (N_1336,N_826,N_866);
nor U1337 (N_1337,N_893,N_188);
and U1338 (N_1338,N_32,N_429);
or U1339 (N_1339,N_278,N_426);
nand U1340 (N_1340,N_297,N_131);
xor U1341 (N_1341,N_663,N_220);
or U1342 (N_1342,N_975,N_925);
or U1343 (N_1343,N_399,N_528);
xor U1344 (N_1344,N_912,N_553);
or U1345 (N_1345,N_735,N_719);
nor U1346 (N_1346,N_712,N_276);
nand U1347 (N_1347,N_50,N_293);
nand U1348 (N_1348,N_559,N_927);
nand U1349 (N_1349,N_880,N_323);
xnor U1350 (N_1350,N_952,N_516);
nor U1351 (N_1351,N_700,N_394);
xor U1352 (N_1352,N_532,N_744);
or U1353 (N_1353,N_135,N_842);
nand U1354 (N_1354,N_589,N_317);
nand U1355 (N_1355,N_262,N_832);
xor U1356 (N_1356,N_780,N_885);
nor U1357 (N_1357,N_51,N_66);
or U1358 (N_1358,N_84,N_309);
nor U1359 (N_1359,N_787,N_244);
and U1360 (N_1360,N_793,N_246);
or U1361 (N_1361,N_477,N_170);
xnor U1362 (N_1362,N_11,N_958);
or U1363 (N_1363,N_995,N_267);
and U1364 (N_1364,N_695,N_535);
nand U1365 (N_1365,N_361,N_327);
nand U1366 (N_1366,N_526,N_123);
nand U1367 (N_1367,N_850,N_863);
and U1368 (N_1368,N_433,N_274);
nand U1369 (N_1369,N_567,N_144);
xnor U1370 (N_1370,N_431,N_840);
xnor U1371 (N_1371,N_802,N_356);
or U1372 (N_1372,N_305,N_292);
nand U1373 (N_1373,N_756,N_30);
and U1374 (N_1374,N_326,N_254);
xnor U1375 (N_1375,N_938,N_810);
or U1376 (N_1376,N_983,N_835);
or U1377 (N_1377,N_363,N_686);
and U1378 (N_1378,N_369,N_236);
nand U1379 (N_1379,N_85,N_538);
nor U1380 (N_1380,N_74,N_386);
nor U1381 (N_1381,N_436,N_209);
and U1382 (N_1382,N_177,N_562);
and U1383 (N_1383,N_592,N_963);
nor U1384 (N_1384,N_675,N_420);
nor U1385 (N_1385,N_989,N_174);
nor U1386 (N_1386,N_268,N_10);
and U1387 (N_1387,N_707,N_203);
nor U1388 (N_1388,N_766,N_841);
and U1389 (N_1389,N_515,N_238);
and U1390 (N_1390,N_798,N_315);
and U1391 (N_1391,N_644,N_782);
nand U1392 (N_1392,N_467,N_231);
nor U1393 (N_1393,N_341,N_355);
nand U1394 (N_1394,N_349,N_232);
xor U1395 (N_1395,N_149,N_661);
xor U1396 (N_1396,N_48,N_419);
nor U1397 (N_1397,N_378,N_338);
nand U1398 (N_1398,N_523,N_199);
nor U1399 (N_1399,N_915,N_776);
xor U1400 (N_1400,N_617,N_875);
and U1401 (N_1401,N_266,N_357);
or U1402 (N_1402,N_393,N_836);
nor U1403 (N_1403,N_750,N_729);
nand U1404 (N_1404,N_366,N_223);
or U1405 (N_1405,N_345,N_25);
nor U1406 (N_1406,N_816,N_988);
nand U1407 (N_1407,N_29,N_352);
xnor U1408 (N_1408,N_862,N_858);
and U1409 (N_1409,N_754,N_818);
and U1410 (N_1410,N_235,N_834);
or U1411 (N_1411,N_156,N_839);
nand U1412 (N_1412,N_495,N_986);
nand U1413 (N_1413,N_629,N_489);
nor U1414 (N_1414,N_768,N_997);
nand U1415 (N_1415,N_561,N_620);
nor U1416 (N_1416,N_230,N_673);
xor U1417 (N_1417,N_652,N_383);
and U1418 (N_1418,N_385,N_180);
nor U1419 (N_1419,N_206,N_558);
nor U1420 (N_1420,N_458,N_5);
nor U1421 (N_1421,N_540,N_594);
or U1422 (N_1422,N_475,N_533);
and U1423 (N_1423,N_555,N_109);
nand U1424 (N_1424,N_196,N_827);
nand U1425 (N_1425,N_75,N_703);
nor U1426 (N_1426,N_395,N_659);
nand U1427 (N_1427,N_435,N_416);
and U1428 (N_1428,N_99,N_664);
xnor U1429 (N_1429,N_746,N_142);
xnor U1430 (N_1430,N_941,N_792);
and U1431 (N_1431,N_665,N_68);
or U1432 (N_1432,N_978,N_907);
nor U1433 (N_1433,N_897,N_856);
or U1434 (N_1434,N_817,N_519);
nand U1435 (N_1435,N_820,N_15);
or U1436 (N_1436,N_45,N_990);
or U1437 (N_1437,N_377,N_940);
or U1438 (N_1438,N_755,N_550);
xor U1439 (N_1439,N_340,N_194);
and U1440 (N_1440,N_574,N_311);
and U1441 (N_1441,N_830,N_692);
nor U1442 (N_1442,N_13,N_255);
and U1443 (N_1443,N_134,N_608);
nand U1444 (N_1444,N_122,N_716);
xor U1445 (N_1445,N_16,N_563);
nor U1446 (N_1446,N_49,N_364);
or U1447 (N_1447,N_241,N_20);
xor U1448 (N_1448,N_113,N_380);
nand U1449 (N_1449,N_481,N_704);
and U1450 (N_1450,N_154,N_721);
nor U1451 (N_1451,N_71,N_623);
or U1452 (N_1452,N_367,N_932);
nand U1453 (N_1453,N_505,N_931);
xnor U1454 (N_1454,N_2,N_530);
and U1455 (N_1455,N_405,N_80);
and U1456 (N_1456,N_889,N_867);
nand U1457 (N_1457,N_511,N_347);
xnor U1458 (N_1458,N_211,N_585);
xor U1459 (N_1459,N_14,N_8);
nand U1460 (N_1460,N_446,N_248);
or U1461 (N_1461,N_37,N_777);
nand U1462 (N_1462,N_646,N_452);
nand U1463 (N_1463,N_250,N_970);
and U1464 (N_1464,N_127,N_358);
nand U1465 (N_1465,N_392,N_404);
nor U1466 (N_1466,N_972,N_586);
xor U1467 (N_1467,N_701,N_977);
or U1468 (N_1468,N_22,N_217);
and U1469 (N_1469,N_647,N_101);
nor U1470 (N_1470,N_847,N_524);
nor U1471 (N_1471,N_607,N_728);
nand U1472 (N_1472,N_973,N_64);
nand U1473 (N_1473,N_295,N_619);
xnor U1474 (N_1474,N_683,N_869);
and U1475 (N_1475,N_618,N_922);
xor U1476 (N_1476,N_660,N_233);
nor U1477 (N_1477,N_504,N_441);
xnor U1478 (N_1478,N_674,N_228);
and U1479 (N_1479,N_771,N_588);
xor U1480 (N_1480,N_499,N_876);
and U1481 (N_1481,N_105,N_138);
nor U1482 (N_1482,N_621,N_450);
nor U1483 (N_1483,N_286,N_384);
xor U1484 (N_1484,N_54,N_373);
nor U1485 (N_1485,N_919,N_129);
or U1486 (N_1486,N_53,N_956);
nor U1487 (N_1487,N_961,N_545);
and U1488 (N_1488,N_46,N_314);
or U1489 (N_1489,N_696,N_600);
nand U1490 (N_1490,N_260,N_331);
nand U1491 (N_1491,N_299,N_584);
and U1492 (N_1492,N_242,N_79);
nand U1493 (N_1493,N_243,N_844);
nor U1494 (N_1494,N_929,N_186);
or U1495 (N_1495,N_933,N_214);
nand U1496 (N_1496,N_759,N_462);
nand U1497 (N_1497,N_21,N_185);
nand U1498 (N_1498,N_451,N_849);
nor U1499 (N_1499,N_861,N_148);
and U1500 (N_1500,N_679,N_225);
nand U1501 (N_1501,N_491,N_422);
nor U1502 (N_1502,N_999,N_312);
nor U1503 (N_1503,N_488,N_783);
xnor U1504 (N_1504,N_169,N_79);
and U1505 (N_1505,N_448,N_765);
nand U1506 (N_1506,N_188,N_198);
nor U1507 (N_1507,N_878,N_972);
xor U1508 (N_1508,N_3,N_554);
xnor U1509 (N_1509,N_224,N_980);
xnor U1510 (N_1510,N_712,N_649);
or U1511 (N_1511,N_642,N_700);
nand U1512 (N_1512,N_651,N_120);
xor U1513 (N_1513,N_984,N_667);
nand U1514 (N_1514,N_198,N_241);
or U1515 (N_1515,N_41,N_677);
nor U1516 (N_1516,N_84,N_141);
and U1517 (N_1517,N_785,N_539);
nor U1518 (N_1518,N_41,N_725);
nand U1519 (N_1519,N_57,N_478);
nand U1520 (N_1520,N_731,N_147);
xor U1521 (N_1521,N_531,N_112);
nor U1522 (N_1522,N_480,N_750);
nor U1523 (N_1523,N_599,N_622);
xor U1524 (N_1524,N_143,N_657);
xor U1525 (N_1525,N_232,N_223);
nor U1526 (N_1526,N_287,N_922);
nand U1527 (N_1527,N_509,N_121);
xor U1528 (N_1528,N_214,N_219);
nor U1529 (N_1529,N_653,N_699);
and U1530 (N_1530,N_345,N_115);
nand U1531 (N_1531,N_936,N_416);
nor U1532 (N_1532,N_278,N_530);
xor U1533 (N_1533,N_955,N_254);
nor U1534 (N_1534,N_616,N_517);
or U1535 (N_1535,N_637,N_53);
and U1536 (N_1536,N_34,N_621);
nand U1537 (N_1537,N_693,N_824);
nand U1538 (N_1538,N_458,N_401);
xnor U1539 (N_1539,N_659,N_241);
xnor U1540 (N_1540,N_350,N_443);
nor U1541 (N_1541,N_51,N_799);
or U1542 (N_1542,N_935,N_735);
xnor U1543 (N_1543,N_922,N_127);
and U1544 (N_1544,N_823,N_390);
xnor U1545 (N_1545,N_205,N_821);
or U1546 (N_1546,N_551,N_500);
xnor U1547 (N_1547,N_841,N_598);
nand U1548 (N_1548,N_960,N_822);
and U1549 (N_1549,N_473,N_129);
xnor U1550 (N_1550,N_468,N_500);
or U1551 (N_1551,N_133,N_389);
or U1552 (N_1552,N_270,N_89);
and U1553 (N_1553,N_331,N_356);
and U1554 (N_1554,N_562,N_388);
nand U1555 (N_1555,N_967,N_750);
and U1556 (N_1556,N_802,N_141);
nand U1557 (N_1557,N_290,N_238);
nand U1558 (N_1558,N_497,N_984);
nand U1559 (N_1559,N_202,N_786);
xor U1560 (N_1560,N_486,N_45);
and U1561 (N_1561,N_473,N_648);
nor U1562 (N_1562,N_494,N_631);
xor U1563 (N_1563,N_80,N_792);
nand U1564 (N_1564,N_785,N_572);
nand U1565 (N_1565,N_658,N_301);
xnor U1566 (N_1566,N_240,N_669);
xor U1567 (N_1567,N_107,N_902);
nor U1568 (N_1568,N_195,N_469);
and U1569 (N_1569,N_666,N_280);
nor U1570 (N_1570,N_704,N_654);
nor U1571 (N_1571,N_178,N_210);
nand U1572 (N_1572,N_168,N_164);
or U1573 (N_1573,N_568,N_189);
xor U1574 (N_1574,N_401,N_839);
or U1575 (N_1575,N_954,N_772);
and U1576 (N_1576,N_465,N_427);
nand U1577 (N_1577,N_884,N_105);
or U1578 (N_1578,N_244,N_278);
and U1579 (N_1579,N_623,N_284);
and U1580 (N_1580,N_572,N_874);
xnor U1581 (N_1581,N_227,N_545);
nand U1582 (N_1582,N_862,N_663);
xnor U1583 (N_1583,N_650,N_1);
xnor U1584 (N_1584,N_962,N_426);
or U1585 (N_1585,N_67,N_541);
or U1586 (N_1586,N_915,N_676);
and U1587 (N_1587,N_13,N_98);
and U1588 (N_1588,N_632,N_126);
nor U1589 (N_1589,N_397,N_790);
xnor U1590 (N_1590,N_639,N_680);
and U1591 (N_1591,N_534,N_794);
or U1592 (N_1592,N_27,N_387);
or U1593 (N_1593,N_423,N_195);
nand U1594 (N_1594,N_504,N_591);
or U1595 (N_1595,N_857,N_464);
and U1596 (N_1596,N_244,N_570);
nand U1597 (N_1597,N_724,N_790);
and U1598 (N_1598,N_239,N_123);
and U1599 (N_1599,N_675,N_240);
xor U1600 (N_1600,N_327,N_761);
xor U1601 (N_1601,N_726,N_500);
and U1602 (N_1602,N_247,N_600);
nor U1603 (N_1603,N_127,N_688);
xor U1604 (N_1604,N_626,N_308);
xnor U1605 (N_1605,N_625,N_781);
nand U1606 (N_1606,N_554,N_416);
xor U1607 (N_1607,N_179,N_346);
nand U1608 (N_1608,N_137,N_713);
xnor U1609 (N_1609,N_156,N_970);
nand U1610 (N_1610,N_539,N_88);
nand U1611 (N_1611,N_232,N_561);
nand U1612 (N_1612,N_185,N_762);
or U1613 (N_1613,N_458,N_408);
xnor U1614 (N_1614,N_557,N_998);
nand U1615 (N_1615,N_785,N_698);
xnor U1616 (N_1616,N_302,N_600);
nand U1617 (N_1617,N_382,N_746);
nor U1618 (N_1618,N_170,N_662);
nand U1619 (N_1619,N_814,N_958);
nand U1620 (N_1620,N_116,N_396);
xor U1621 (N_1621,N_902,N_589);
nand U1622 (N_1622,N_860,N_982);
xnor U1623 (N_1623,N_101,N_509);
nand U1624 (N_1624,N_114,N_122);
and U1625 (N_1625,N_838,N_370);
or U1626 (N_1626,N_263,N_215);
or U1627 (N_1627,N_663,N_184);
nor U1628 (N_1628,N_867,N_588);
nor U1629 (N_1629,N_158,N_978);
and U1630 (N_1630,N_159,N_355);
and U1631 (N_1631,N_353,N_475);
and U1632 (N_1632,N_599,N_568);
or U1633 (N_1633,N_904,N_709);
nor U1634 (N_1634,N_865,N_117);
nor U1635 (N_1635,N_986,N_936);
xor U1636 (N_1636,N_5,N_42);
nand U1637 (N_1637,N_422,N_360);
nand U1638 (N_1638,N_783,N_38);
xnor U1639 (N_1639,N_980,N_998);
nor U1640 (N_1640,N_233,N_64);
or U1641 (N_1641,N_290,N_671);
nand U1642 (N_1642,N_631,N_260);
and U1643 (N_1643,N_805,N_906);
xnor U1644 (N_1644,N_819,N_340);
nor U1645 (N_1645,N_455,N_216);
and U1646 (N_1646,N_865,N_238);
xor U1647 (N_1647,N_474,N_593);
xor U1648 (N_1648,N_304,N_771);
and U1649 (N_1649,N_370,N_984);
nor U1650 (N_1650,N_368,N_994);
and U1651 (N_1651,N_354,N_86);
and U1652 (N_1652,N_453,N_368);
and U1653 (N_1653,N_800,N_947);
nor U1654 (N_1654,N_351,N_37);
xor U1655 (N_1655,N_388,N_766);
nand U1656 (N_1656,N_560,N_513);
nand U1657 (N_1657,N_426,N_492);
or U1658 (N_1658,N_164,N_616);
nor U1659 (N_1659,N_223,N_899);
or U1660 (N_1660,N_843,N_356);
or U1661 (N_1661,N_199,N_780);
or U1662 (N_1662,N_177,N_785);
nor U1663 (N_1663,N_750,N_462);
nand U1664 (N_1664,N_749,N_480);
nand U1665 (N_1665,N_139,N_73);
and U1666 (N_1666,N_545,N_669);
and U1667 (N_1667,N_184,N_873);
xor U1668 (N_1668,N_36,N_68);
xor U1669 (N_1669,N_968,N_442);
and U1670 (N_1670,N_634,N_318);
nor U1671 (N_1671,N_340,N_992);
nor U1672 (N_1672,N_720,N_312);
or U1673 (N_1673,N_551,N_872);
or U1674 (N_1674,N_42,N_940);
nand U1675 (N_1675,N_766,N_405);
xnor U1676 (N_1676,N_909,N_780);
and U1677 (N_1677,N_358,N_248);
xnor U1678 (N_1678,N_693,N_596);
and U1679 (N_1679,N_951,N_347);
nand U1680 (N_1680,N_358,N_697);
nor U1681 (N_1681,N_963,N_863);
or U1682 (N_1682,N_934,N_330);
or U1683 (N_1683,N_196,N_143);
and U1684 (N_1684,N_312,N_762);
nand U1685 (N_1685,N_385,N_138);
xnor U1686 (N_1686,N_159,N_17);
nand U1687 (N_1687,N_703,N_5);
nor U1688 (N_1688,N_972,N_436);
or U1689 (N_1689,N_931,N_868);
xor U1690 (N_1690,N_18,N_955);
nor U1691 (N_1691,N_363,N_335);
nor U1692 (N_1692,N_301,N_119);
or U1693 (N_1693,N_331,N_355);
xor U1694 (N_1694,N_761,N_32);
xor U1695 (N_1695,N_204,N_617);
and U1696 (N_1696,N_975,N_842);
xnor U1697 (N_1697,N_237,N_131);
nand U1698 (N_1698,N_790,N_434);
nor U1699 (N_1699,N_743,N_282);
xor U1700 (N_1700,N_865,N_535);
xnor U1701 (N_1701,N_461,N_277);
nand U1702 (N_1702,N_540,N_553);
or U1703 (N_1703,N_664,N_17);
and U1704 (N_1704,N_216,N_497);
nand U1705 (N_1705,N_997,N_715);
nor U1706 (N_1706,N_561,N_68);
and U1707 (N_1707,N_169,N_973);
or U1708 (N_1708,N_250,N_689);
and U1709 (N_1709,N_954,N_585);
nand U1710 (N_1710,N_450,N_355);
nand U1711 (N_1711,N_768,N_944);
nand U1712 (N_1712,N_199,N_426);
nor U1713 (N_1713,N_252,N_97);
or U1714 (N_1714,N_609,N_250);
and U1715 (N_1715,N_943,N_725);
and U1716 (N_1716,N_681,N_63);
nor U1717 (N_1717,N_972,N_378);
xnor U1718 (N_1718,N_81,N_731);
nand U1719 (N_1719,N_623,N_82);
or U1720 (N_1720,N_208,N_205);
xnor U1721 (N_1721,N_941,N_870);
and U1722 (N_1722,N_99,N_695);
and U1723 (N_1723,N_967,N_147);
and U1724 (N_1724,N_270,N_442);
and U1725 (N_1725,N_212,N_799);
or U1726 (N_1726,N_677,N_570);
and U1727 (N_1727,N_729,N_357);
nor U1728 (N_1728,N_168,N_122);
nand U1729 (N_1729,N_215,N_678);
xnor U1730 (N_1730,N_854,N_983);
and U1731 (N_1731,N_343,N_355);
nand U1732 (N_1732,N_813,N_773);
xor U1733 (N_1733,N_16,N_950);
and U1734 (N_1734,N_169,N_461);
xnor U1735 (N_1735,N_41,N_63);
nand U1736 (N_1736,N_44,N_529);
and U1737 (N_1737,N_471,N_730);
and U1738 (N_1738,N_71,N_21);
or U1739 (N_1739,N_663,N_340);
nor U1740 (N_1740,N_901,N_52);
nand U1741 (N_1741,N_860,N_106);
or U1742 (N_1742,N_2,N_27);
nand U1743 (N_1743,N_222,N_303);
or U1744 (N_1744,N_327,N_545);
and U1745 (N_1745,N_970,N_808);
or U1746 (N_1746,N_912,N_146);
and U1747 (N_1747,N_541,N_77);
nor U1748 (N_1748,N_273,N_271);
or U1749 (N_1749,N_205,N_905);
nand U1750 (N_1750,N_144,N_688);
or U1751 (N_1751,N_321,N_677);
and U1752 (N_1752,N_3,N_203);
xnor U1753 (N_1753,N_659,N_800);
nand U1754 (N_1754,N_135,N_199);
nor U1755 (N_1755,N_513,N_44);
nor U1756 (N_1756,N_623,N_334);
nand U1757 (N_1757,N_65,N_163);
xnor U1758 (N_1758,N_260,N_194);
xor U1759 (N_1759,N_862,N_874);
and U1760 (N_1760,N_190,N_662);
and U1761 (N_1761,N_158,N_911);
xnor U1762 (N_1762,N_209,N_23);
or U1763 (N_1763,N_748,N_198);
and U1764 (N_1764,N_794,N_813);
nor U1765 (N_1765,N_253,N_258);
nor U1766 (N_1766,N_969,N_121);
xnor U1767 (N_1767,N_572,N_474);
or U1768 (N_1768,N_448,N_707);
and U1769 (N_1769,N_306,N_204);
xnor U1770 (N_1770,N_990,N_563);
nand U1771 (N_1771,N_889,N_167);
nand U1772 (N_1772,N_763,N_742);
nand U1773 (N_1773,N_272,N_352);
or U1774 (N_1774,N_365,N_707);
nand U1775 (N_1775,N_293,N_39);
or U1776 (N_1776,N_560,N_571);
nand U1777 (N_1777,N_967,N_36);
nor U1778 (N_1778,N_722,N_429);
nand U1779 (N_1779,N_838,N_836);
nand U1780 (N_1780,N_547,N_653);
nor U1781 (N_1781,N_166,N_59);
nor U1782 (N_1782,N_197,N_434);
nor U1783 (N_1783,N_910,N_143);
nor U1784 (N_1784,N_947,N_639);
or U1785 (N_1785,N_258,N_43);
nor U1786 (N_1786,N_437,N_857);
nor U1787 (N_1787,N_307,N_861);
xnor U1788 (N_1788,N_779,N_458);
nand U1789 (N_1789,N_723,N_848);
or U1790 (N_1790,N_437,N_42);
or U1791 (N_1791,N_897,N_88);
nor U1792 (N_1792,N_798,N_353);
and U1793 (N_1793,N_802,N_827);
nor U1794 (N_1794,N_754,N_767);
nor U1795 (N_1795,N_580,N_127);
xor U1796 (N_1796,N_262,N_193);
nor U1797 (N_1797,N_324,N_753);
nand U1798 (N_1798,N_217,N_230);
and U1799 (N_1799,N_242,N_116);
and U1800 (N_1800,N_684,N_396);
nor U1801 (N_1801,N_340,N_969);
and U1802 (N_1802,N_936,N_222);
and U1803 (N_1803,N_445,N_810);
nor U1804 (N_1804,N_302,N_592);
nand U1805 (N_1805,N_551,N_676);
nor U1806 (N_1806,N_488,N_376);
nand U1807 (N_1807,N_599,N_830);
or U1808 (N_1808,N_816,N_822);
nor U1809 (N_1809,N_517,N_7);
or U1810 (N_1810,N_100,N_699);
nand U1811 (N_1811,N_200,N_509);
or U1812 (N_1812,N_741,N_107);
and U1813 (N_1813,N_66,N_949);
xnor U1814 (N_1814,N_937,N_105);
and U1815 (N_1815,N_610,N_856);
nor U1816 (N_1816,N_660,N_472);
nand U1817 (N_1817,N_21,N_131);
or U1818 (N_1818,N_460,N_444);
nand U1819 (N_1819,N_638,N_247);
nand U1820 (N_1820,N_587,N_931);
nand U1821 (N_1821,N_15,N_641);
and U1822 (N_1822,N_802,N_689);
xor U1823 (N_1823,N_2,N_762);
xor U1824 (N_1824,N_785,N_457);
or U1825 (N_1825,N_556,N_813);
and U1826 (N_1826,N_554,N_522);
xnor U1827 (N_1827,N_849,N_379);
and U1828 (N_1828,N_0,N_887);
nor U1829 (N_1829,N_634,N_792);
and U1830 (N_1830,N_98,N_513);
nand U1831 (N_1831,N_933,N_592);
nor U1832 (N_1832,N_903,N_98);
nor U1833 (N_1833,N_456,N_191);
or U1834 (N_1834,N_800,N_132);
xnor U1835 (N_1835,N_41,N_678);
nor U1836 (N_1836,N_976,N_370);
nand U1837 (N_1837,N_51,N_945);
nor U1838 (N_1838,N_225,N_778);
and U1839 (N_1839,N_222,N_271);
and U1840 (N_1840,N_716,N_592);
nor U1841 (N_1841,N_995,N_327);
or U1842 (N_1842,N_155,N_615);
or U1843 (N_1843,N_643,N_866);
or U1844 (N_1844,N_946,N_630);
nand U1845 (N_1845,N_888,N_549);
xor U1846 (N_1846,N_498,N_97);
or U1847 (N_1847,N_368,N_571);
nor U1848 (N_1848,N_673,N_247);
or U1849 (N_1849,N_439,N_665);
nand U1850 (N_1850,N_136,N_736);
nand U1851 (N_1851,N_145,N_608);
or U1852 (N_1852,N_173,N_855);
and U1853 (N_1853,N_237,N_970);
nand U1854 (N_1854,N_478,N_925);
or U1855 (N_1855,N_597,N_272);
and U1856 (N_1856,N_871,N_435);
nor U1857 (N_1857,N_625,N_414);
and U1858 (N_1858,N_372,N_566);
or U1859 (N_1859,N_764,N_443);
xor U1860 (N_1860,N_633,N_970);
nor U1861 (N_1861,N_655,N_176);
xor U1862 (N_1862,N_576,N_23);
xor U1863 (N_1863,N_25,N_992);
or U1864 (N_1864,N_170,N_415);
nor U1865 (N_1865,N_333,N_20);
and U1866 (N_1866,N_843,N_163);
and U1867 (N_1867,N_809,N_379);
nor U1868 (N_1868,N_457,N_821);
nor U1869 (N_1869,N_883,N_785);
and U1870 (N_1870,N_348,N_182);
and U1871 (N_1871,N_512,N_623);
and U1872 (N_1872,N_439,N_310);
nor U1873 (N_1873,N_140,N_321);
or U1874 (N_1874,N_779,N_816);
xor U1875 (N_1875,N_38,N_867);
or U1876 (N_1876,N_638,N_273);
xnor U1877 (N_1877,N_364,N_851);
nand U1878 (N_1878,N_228,N_994);
nand U1879 (N_1879,N_813,N_208);
nand U1880 (N_1880,N_380,N_625);
nand U1881 (N_1881,N_833,N_189);
nor U1882 (N_1882,N_603,N_98);
nor U1883 (N_1883,N_858,N_341);
nor U1884 (N_1884,N_407,N_961);
nand U1885 (N_1885,N_382,N_4);
nor U1886 (N_1886,N_283,N_21);
and U1887 (N_1887,N_521,N_942);
nor U1888 (N_1888,N_149,N_146);
or U1889 (N_1889,N_209,N_917);
xor U1890 (N_1890,N_150,N_628);
nand U1891 (N_1891,N_70,N_230);
xnor U1892 (N_1892,N_722,N_462);
nand U1893 (N_1893,N_675,N_315);
or U1894 (N_1894,N_504,N_673);
xor U1895 (N_1895,N_462,N_194);
nor U1896 (N_1896,N_853,N_469);
xor U1897 (N_1897,N_856,N_960);
or U1898 (N_1898,N_432,N_490);
nor U1899 (N_1899,N_81,N_739);
or U1900 (N_1900,N_220,N_490);
nor U1901 (N_1901,N_599,N_919);
xor U1902 (N_1902,N_453,N_708);
and U1903 (N_1903,N_368,N_173);
nand U1904 (N_1904,N_296,N_811);
xnor U1905 (N_1905,N_74,N_482);
xor U1906 (N_1906,N_585,N_490);
nand U1907 (N_1907,N_778,N_842);
nor U1908 (N_1908,N_215,N_232);
nor U1909 (N_1909,N_469,N_676);
nand U1910 (N_1910,N_683,N_231);
and U1911 (N_1911,N_775,N_574);
xnor U1912 (N_1912,N_101,N_227);
and U1913 (N_1913,N_54,N_991);
nor U1914 (N_1914,N_659,N_57);
nand U1915 (N_1915,N_342,N_536);
nor U1916 (N_1916,N_605,N_597);
or U1917 (N_1917,N_197,N_835);
nand U1918 (N_1918,N_883,N_615);
or U1919 (N_1919,N_9,N_777);
or U1920 (N_1920,N_344,N_215);
nor U1921 (N_1921,N_834,N_940);
nor U1922 (N_1922,N_292,N_634);
nor U1923 (N_1923,N_757,N_215);
xnor U1924 (N_1924,N_192,N_384);
or U1925 (N_1925,N_533,N_846);
nand U1926 (N_1926,N_983,N_884);
nand U1927 (N_1927,N_276,N_256);
nor U1928 (N_1928,N_879,N_448);
nor U1929 (N_1929,N_97,N_883);
or U1930 (N_1930,N_734,N_885);
xor U1931 (N_1931,N_561,N_376);
and U1932 (N_1932,N_637,N_248);
xnor U1933 (N_1933,N_714,N_897);
xnor U1934 (N_1934,N_738,N_871);
nand U1935 (N_1935,N_270,N_727);
xnor U1936 (N_1936,N_217,N_513);
and U1937 (N_1937,N_604,N_546);
xor U1938 (N_1938,N_359,N_294);
nor U1939 (N_1939,N_793,N_254);
xor U1940 (N_1940,N_765,N_392);
xor U1941 (N_1941,N_153,N_590);
or U1942 (N_1942,N_89,N_616);
xor U1943 (N_1943,N_811,N_734);
or U1944 (N_1944,N_10,N_454);
or U1945 (N_1945,N_186,N_217);
and U1946 (N_1946,N_49,N_394);
xor U1947 (N_1947,N_520,N_218);
and U1948 (N_1948,N_597,N_148);
or U1949 (N_1949,N_293,N_562);
xor U1950 (N_1950,N_61,N_247);
or U1951 (N_1951,N_675,N_425);
xor U1952 (N_1952,N_495,N_788);
nand U1953 (N_1953,N_987,N_454);
xor U1954 (N_1954,N_501,N_807);
xor U1955 (N_1955,N_886,N_582);
nor U1956 (N_1956,N_801,N_346);
xor U1957 (N_1957,N_912,N_258);
nor U1958 (N_1958,N_714,N_558);
nand U1959 (N_1959,N_204,N_250);
and U1960 (N_1960,N_371,N_108);
nand U1961 (N_1961,N_237,N_43);
xnor U1962 (N_1962,N_510,N_545);
xnor U1963 (N_1963,N_598,N_394);
nor U1964 (N_1964,N_68,N_572);
or U1965 (N_1965,N_751,N_102);
or U1966 (N_1966,N_846,N_532);
or U1967 (N_1967,N_929,N_301);
or U1968 (N_1968,N_666,N_975);
or U1969 (N_1969,N_665,N_493);
nor U1970 (N_1970,N_243,N_779);
and U1971 (N_1971,N_213,N_324);
xnor U1972 (N_1972,N_33,N_193);
xnor U1973 (N_1973,N_727,N_16);
or U1974 (N_1974,N_71,N_503);
nand U1975 (N_1975,N_464,N_484);
xnor U1976 (N_1976,N_562,N_729);
or U1977 (N_1977,N_636,N_251);
nand U1978 (N_1978,N_560,N_303);
nor U1979 (N_1979,N_780,N_778);
nor U1980 (N_1980,N_291,N_187);
and U1981 (N_1981,N_269,N_557);
xnor U1982 (N_1982,N_599,N_714);
or U1983 (N_1983,N_97,N_901);
or U1984 (N_1984,N_574,N_952);
or U1985 (N_1985,N_314,N_407);
and U1986 (N_1986,N_473,N_24);
xor U1987 (N_1987,N_883,N_578);
nand U1988 (N_1988,N_78,N_11);
nor U1989 (N_1989,N_994,N_755);
nand U1990 (N_1990,N_385,N_426);
nor U1991 (N_1991,N_98,N_959);
and U1992 (N_1992,N_914,N_709);
and U1993 (N_1993,N_577,N_708);
and U1994 (N_1994,N_446,N_330);
nand U1995 (N_1995,N_895,N_659);
xnor U1996 (N_1996,N_757,N_36);
and U1997 (N_1997,N_318,N_70);
or U1998 (N_1998,N_692,N_951);
or U1999 (N_1999,N_242,N_598);
nand U2000 (N_2000,N_1758,N_1502);
xnor U2001 (N_2001,N_1936,N_1759);
and U2002 (N_2002,N_1580,N_1333);
nand U2003 (N_2003,N_1428,N_1357);
nor U2004 (N_2004,N_1078,N_1185);
xnor U2005 (N_2005,N_1953,N_1760);
nand U2006 (N_2006,N_1343,N_1263);
nor U2007 (N_2007,N_1354,N_1103);
xor U2008 (N_2008,N_1996,N_1269);
nand U2009 (N_2009,N_1014,N_1607);
nand U2010 (N_2010,N_1605,N_1823);
or U2011 (N_2011,N_1283,N_1739);
xor U2012 (N_2012,N_1179,N_1683);
or U2013 (N_2013,N_1437,N_1167);
and U2014 (N_2014,N_1470,N_1472);
and U2015 (N_2015,N_1433,N_1136);
nand U2016 (N_2016,N_1853,N_1532);
nor U2017 (N_2017,N_1616,N_1315);
and U2018 (N_2018,N_1553,N_1714);
or U2019 (N_2019,N_1864,N_1304);
and U2020 (N_2020,N_1265,N_1647);
and U2021 (N_2021,N_1541,N_1915);
and U2022 (N_2022,N_1126,N_1220);
xor U2023 (N_2023,N_1518,N_1694);
or U2024 (N_2024,N_1319,N_1260);
and U2025 (N_2025,N_1109,N_1379);
xor U2026 (N_2026,N_1296,N_1848);
nand U2027 (N_2027,N_1091,N_1908);
xnor U2028 (N_2028,N_1123,N_1106);
nand U2029 (N_2029,N_1350,N_1652);
or U2030 (N_2030,N_1514,N_1599);
and U2031 (N_2031,N_1799,N_1337);
nand U2032 (N_2032,N_1551,N_1496);
nor U2033 (N_2033,N_1271,N_1400);
and U2034 (N_2034,N_1798,N_1554);
or U2035 (N_2035,N_1802,N_1197);
or U2036 (N_2036,N_1373,N_1385);
or U2037 (N_2037,N_1279,N_1439);
and U2038 (N_2038,N_1979,N_1672);
nor U2039 (N_2039,N_1305,N_1447);
nor U2040 (N_2040,N_1187,N_1827);
xor U2041 (N_2041,N_1468,N_1158);
or U2042 (N_2042,N_1483,N_1028);
xnor U2043 (N_2043,N_1509,N_1576);
xnor U2044 (N_2044,N_1199,N_1239);
and U2045 (N_2045,N_1035,N_1222);
or U2046 (N_2046,N_1963,N_1741);
or U2047 (N_2047,N_1013,N_1837);
or U2048 (N_2048,N_1768,N_1678);
nor U2049 (N_2049,N_1087,N_1648);
nand U2050 (N_2050,N_1570,N_1467);
and U2051 (N_2051,N_1590,N_1019);
nor U2052 (N_2052,N_1773,N_1165);
or U2053 (N_2053,N_1724,N_1191);
nor U2054 (N_2054,N_1670,N_1164);
or U2055 (N_2055,N_1059,N_1726);
or U2056 (N_2056,N_1620,N_1940);
or U2057 (N_2057,N_1662,N_1029);
or U2058 (N_2058,N_1568,N_1392);
and U2059 (N_2059,N_1588,N_1493);
or U2060 (N_2060,N_1812,N_1521);
nor U2061 (N_2061,N_1184,N_1905);
nor U2062 (N_2062,N_1077,N_1891);
or U2063 (N_2063,N_1453,N_1317);
and U2064 (N_2064,N_1805,N_1828);
xor U2065 (N_2065,N_1387,N_1107);
xor U2066 (N_2066,N_1204,N_1881);
nor U2067 (N_2067,N_1644,N_1376);
xnor U2068 (N_2068,N_1489,N_1162);
or U2069 (N_2069,N_1064,N_1847);
nor U2070 (N_2070,N_1398,N_1173);
nor U2071 (N_2071,N_1135,N_1210);
xor U2072 (N_2072,N_1024,N_1093);
and U2073 (N_2073,N_1508,N_1564);
and U2074 (N_2074,N_1976,N_1414);
nor U2075 (N_2075,N_1461,N_1095);
nand U2076 (N_2076,N_1657,N_1249);
or U2077 (N_2077,N_1443,N_1270);
nor U2078 (N_2078,N_1840,N_1170);
nor U2079 (N_2079,N_1535,N_1854);
xor U2080 (N_2080,N_1193,N_1182);
and U2081 (N_2081,N_1355,N_1870);
nor U2082 (N_2082,N_1094,N_1448);
and U2083 (N_2083,N_1693,N_1757);
xnor U2084 (N_2084,N_1410,N_1115);
xor U2085 (N_2085,N_1866,N_1331);
nand U2086 (N_2086,N_1506,N_1890);
nor U2087 (N_2087,N_1838,N_1415);
and U2088 (N_2088,N_1120,N_1086);
nand U2089 (N_2089,N_1937,N_1227);
nor U2090 (N_2090,N_1688,N_1190);
and U2091 (N_2091,N_1313,N_1674);
xnor U2092 (N_2092,N_1062,N_1749);
nand U2093 (N_2093,N_1995,N_1946);
nand U2094 (N_2094,N_1863,N_1036);
and U2095 (N_2095,N_1214,N_1237);
xnor U2096 (N_2096,N_1650,N_1743);
or U2097 (N_2097,N_1980,N_1617);
and U2098 (N_2098,N_1351,N_1619);
and U2099 (N_2099,N_1292,N_1441);
xor U2100 (N_2100,N_1941,N_1865);
xnor U2101 (N_2101,N_1732,N_1056);
xor U2102 (N_2102,N_1321,N_1733);
nor U2103 (N_2103,N_1073,N_1485);
xnor U2104 (N_2104,N_1593,N_1851);
or U2105 (N_2105,N_1667,N_1690);
nor U2106 (N_2106,N_1904,N_1744);
nand U2107 (N_2107,N_1556,N_1500);
xnor U2108 (N_2108,N_1044,N_1618);
nor U2109 (N_2109,N_1329,N_1407);
and U2110 (N_2110,N_1591,N_1018);
xnor U2111 (N_2111,N_1640,N_1037);
or U2112 (N_2112,N_1386,N_1278);
xor U2113 (N_2113,N_1643,N_1814);
nor U2114 (N_2114,N_1302,N_1651);
and U2115 (N_2115,N_1228,N_1318);
and U2116 (N_2116,N_1806,N_1686);
nor U2117 (N_2117,N_1572,N_1677);
xnor U2118 (N_2118,N_1346,N_1801);
and U2119 (N_2119,N_1928,N_1931);
or U2120 (N_2120,N_1314,N_1188);
nor U2121 (N_2121,N_1026,N_1703);
or U2122 (N_2122,N_1253,N_1082);
or U2123 (N_2123,N_1586,N_1034);
xor U2124 (N_2124,N_1911,N_1236);
nor U2125 (N_2125,N_1010,N_1923);
nand U2126 (N_2126,N_1324,N_1510);
and U2127 (N_2127,N_1702,N_1339);
or U2128 (N_2128,N_1246,N_1396);
nand U2129 (N_2129,N_1665,N_1032);
and U2130 (N_2130,N_1965,N_1810);
or U2131 (N_2131,N_1559,N_1008);
nand U2132 (N_2132,N_1110,N_1245);
or U2133 (N_2133,N_1133,N_1431);
or U2134 (N_2134,N_1708,N_1765);
and U2135 (N_2135,N_1862,N_1074);
xnor U2136 (N_2136,N_1178,N_1452);
xnor U2137 (N_2137,N_1762,N_1574);
nand U2138 (N_2138,N_1132,N_1338);
and U2139 (N_2139,N_1131,N_1161);
or U2140 (N_2140,N_1927,N_1836);
nand U2141 (N_2141,N_1769,N_1705);
and U2142 (N_2142,N_1503,N_1168);
xor U2143 (N_2143,N_1088,N_1456);
nor U2144 (N_2144,N_1918,N_1846);
nand U2145 (N_2145,N_1780,N_1139);
nand U2146 (N_2146,N_1886,N_1458);
or U2147 (N_2147,N_1982,N_1994);
nand U2148 (N_2148,N_1868,N_1839);
nand U2149 (N_2149,N_1406,N_1740);
nand U2150 (N_2150,N_1203,N_1397);
xnor U2151 (N_2151,N_1235,N_1303);
nor U2152 (N_2152,N_1015,N_1171);
or U2153 (N_2153,N_1877,N_1912);
and U2154 (N_2154,N_1910,N_1804);
and U2155 (N_2155,N_1573,N_1033);
xor U2156 (N_2156,N_1790,N_1924);
and U2157 (N_2157,N_1858,N_1875);
nor U2158 (N_2158,N_1763,N_1540);
xor U2159 (N_2159,N_1516,N_1920);
nand U2160 (N_2160,N_1523,N_1603);
xnor U2161 (N_2161,N_1205,N_1089);
nand U2162 (N_2162,N_1613,N_1309);
nand U2163 (N_2163,N_1311,N_1080);
nand U2164 (N_2164,N_1718,N_1772);
and U2165 (N_2165,N_1697,N_1796);
and U2166 (N_2166,N_1720,N_1916);
nand U2167 (N_2167,N_1990,N_1753);
or U2168 (N_2168,N_1819,N_1345);
or U2169 (N_2169,N_1577,N_1887);
xnor U2170 (N_2170,N_1943,N_1102);
nor U2171 (N_2171,N_1975,N_1104);
nand U2172 (N_2172,N_1567,N_1186);
nor U2173 (N_2173,N_1889,N_1435);
or U2174 (N_2174,N_1874,N_1192);
and U2175 (N_2175,N_1378,N_1566);
or U2176 (N_2176,N_1709,N_1584);
and U2177 (N_2177,N_1861,N_1215);
or U2178 (N_2178,N_1207,N_1009);
and U2179 (N_2179,N_1334,N_1427);
nor U2180 (N_2180,N_1101,N_1180);
nor U2181 (N_2181,N_1999,N_1728);
nor U2182 (N_2182,N_1002,N_1970);
nand U2183 (N_2183,N_1692,N_1942);
nand U2184 (N_2184,N_1229,N_1820);
and U2185 (N_2185,N_1706,N_1112);
nand U2186 (N_2186,N_1884,N_1153);
nand U2187 (N_2187,N_1234,N_1972);
and U2188 (N_2188,N_1842,N_1770);
or U2189 (N_2189,N_1710,N_1646);
and U2190 (N_2190,N_1835,N_1582);
nand U2191 (N_2191,N_1156,N_1715);
nor U2192 (N_2192,N_1154,N_1257);
nor U2193 (N_2193,N_1140,N_1707);
nand U2194 (N_2194,N_1501,N_1625);
nor U2195 (N_2195,N_1731,N_1680);
nand U2196 (N_2196,N_1174,N_1543);
nand U2197 (N_2197,N_1370,N_1108);
nand U2198 (N_2198,N_1211,N_1206);
or U2199 (N_2199,N_1536,N_1785);
and U2200 (N_2200,N_1849,N_1627);
and U2201 (N_2201,N_1114,N_1560);
nor U2202 (N_2202,N_1469,N_1954);
xnor U2203 (N_2203,N_1713,N_1579);
nand U2204 (N_2204,N_1267,N_1668);
xor U2205 (N_2205,N_1117,N_1711);
xor U2206 (N_2206,N_1575,N_1699);
nand U2207 (N_2207,N_1050,N_1383);
and U2208 (N_2208,N_1360,N_1546);
xnor U2209 (N_2209,N_1494,N_1423);
or U2210 (N_2210,N_1226,N_1783);
and U2211 (N_2211,N_1020,N_1045);
nand U2212 (N_2212,N_1833,N_1090);
or U2213 (N_2213,N_1634,N_1127);
and U2214 (N_2214,N_1907,N_1476);
and U2215 (N_2215,N_1888,N_1826);
nor U2216 (N_2216,N_1611,N_1098);
xor U2217 (N_2217,N_1150,N_1202);
nor U2218 (N_2218,N_1176,N_1764);
xnor U2219 (N_2219,N_1442,N_1776);
nor U2220 (N_2220,N_1460,N_1636);
nand U2221 (N_2221,N_1602,N_1654);
and U2222 (N_2222,N_1121,N_1388);
nand U2223 (N_2223,N_1793,N_1195);
xnor U2224 (N_2224,N_1834,N_1285);
xnor U2225 (N_2225,N_1957,N_1487);
and U2226 (N_2226,N_1007,N_1061);
or U2227 (N_2227,N_1601,N_1983);
and U2228 (N_2228,N_1375,N_1198);
or U2229 (N_2229,N_1438,N_1233);
nand U2230 (N_2230,N_1981,N_1216);
xnor U2231 (N_2231,N_1716,N_1779);
nand U2232 (N_2232,N_1374,N_1641);
nor U2233 (N_2233,N_1615,N_1621);
nand U2234 (N_2234,N_1399,N_1977);
or U2235 (N_2235,N_1522,N_1259);
or U2236 (N_2236,N_1001,N_1561);
xor U2237 (N_2237,N_1956,N_1592);
nor U2238 (N_2238,N_1539,N_1276);
nand U2239 (N_2239,N_1172,N_1721);
or U2240 (N_2240,N_1053,N_1196);
nor U2241 (N_2241,N_1538,N_1160);
or U2242 (N_2242,N_1390,N_1791);
xor U2243 (N_2243,N_1991,N_1633);
nor U2244 (N_2244,N_1017,N_1049);
and U2245 (N_2245,N_1282,N_1902);
and U2246 (N_2246,N_1882,N_1655);
and U2247 (N_2247,N_1571,N_1581);
nor U2248 (N_2248,N_1352,N_1288);
nand U2249 (N_2249,N_1722,N_1040);
nor U2250 (N_2250,N_1039,N_1134);
xor U2251 (N_2251,N_1065,N_1903);
nor U2252 (N_2252,N_1395,N_1482);
and U2253 (N_2253,N_1047,N_1097);
or U2254 (N_2254,N_1926,N_1052);
xnor U2255 (N_2255,N_1252,N_1585);
nor U2256 (N_2256,N_1012,N_1307);
xor U2257 (N_2257,N_1830,N_1752);
nor U2258 (N_2258,N_1027,N_1816);
nand U2259 (N_2259,N_1878,N_1023);
and U2260 (N_2260,N_1664,N_1869);
nor U2261 (N_2261,N_1434,N_1921);
nor U2262 (N_2262,N_1898,N_1076);
or U2263 (N_2263,N_1929,N_1671);
nor U2264 (N_2264,N_1661,N_1320);
xor U2265 (N_2265,N_1681,N_1043);
xor U2266 (N_2266,N_1843,N_1003);
nor U2267 (N_2267,N_1578,N_1358);
xor U2268 (N_2268,N_1105,N_1380);
or U2269 (N_2269,N_1030,N_1323);
and U2270 (N_2270,N_1143,N_1159);
nor U2271 (N_2271,N_1359,N_1058);
or U2272 (N_2272,N_1209,N_1057);
nand U2273 (N_2273,N_1381,N_1701);
xor U2274 (N_2274,N_1529,N_1232);
and U2275 (N_2275,N_1455,N_1416);
nand U2276 (N_2276,N_1829,N_1860);
nor U2277 (N_2277,N_1961,N_1958);
or U2278 (N_2278,N_1771,N_1526);
or U2279 (N_2279,N_1124,N_1436);
nand U2280 (N_2280,N_1565,N_1213);
xor U2281 (N_2281,N_1988,N_1348);
or U2282 (N_2282,N_1212,N_1258);
or U2283 (N_2283,N_1254,N_1629);
nand U2284 (N_2284,N_1746,N_1642);
xnor U2285 (N_2285,N_1925,N_1275);
xnor U2286 (N_2286,N_1281,N_1507);
or U2287 (N_2287,N_1939,N_1660);
xnor U2288 (N_2288,N_1984,N_1729);
nand U2289 (N_2289,N_1060,N_1445);
or U2290 (N_2290,N_1291,N_1363);
and U2291 (N_2291,N_1788,N_1069);
or U2292 (N_2292,N_1967,N_1264);
or U2293 (N_2293,N_1824,N_1429);
nor U2294 (N_2294,N_1774,N_1473);
and U2295 (N_2295,N_1492,N_1474);
or U2296 (N_2296,N_1063,N_1300);
xnor U2297 (N_2297,N_1649,N_1755);
or U2298 (N_2298,N_1084,N_1832);
xor U2299 (N_2299,N_1504,N_1085);
and U2300 (N_2300,N_1223,N_1969);
nor U2301 (N_2301,N_1730,N_1340);
and U2302 (N_2302,N_1287,N_1597);
nor U2303 (N_2303,N_1369,N_1653);
xor U2304 (N_2304,N_1673,N_1335);
or U2305 (N_2305,N_1895,N_1738);
nor U2306 (N_2306,N_1238,N_1480);
and U2307 (N_2307,N_1808,N_1450);
xor U2308 (N_2308,N_1778,N_1964);
nand U2309 (N_2309,N_1517,N_1725);
and U2310 (N_2310,N_1596,N_1815);
nor U2311 (N_2311,N_1747,N_1952);
and U2312 (N_2312,N_1623,N_1850);
or U2313 (N_2313,N_1119,N_1817);
or U2314 (N_2314,N_1736,N_1189);
xor U2315 (N_2315,N_1530,N_1682);
nand U2316 (N_2316,N_1499,N_1217);
nand U2317 (N_2317,N_1831,N_1691);
xor U2318 (N_2318,N_1368,N_1297);
xor U2319 (N_2319,N_1389,N_1930);
nor U2320 (N_2320,N_1457,N_1242);
nor U2321 (N_2321,N_1951,N_1147);
nor U2322 (N_2322,N_1322,N_1118);
nand U2323 (N_2323,N_1872,N_1513);
nor U2324 (N_2324,N_1344,N_1308);
nand U2325 (N_2325,N_1221,N_1481);
nor U2326 (N_2326,N_1745,N_1272);
and U2327 (N_2327,N_1966,N_1631);
nand U2328 (N_2328,N_1251,N_1520);
nor U2329 (N_2329,N_1989,N_1372);
nor U2330 (N_2330,N_1695,N_1645);
nand U2331 (N_2331,N_1255,N_1301);
and U2332 (N_2332,N_1800,N_1262);
and U2333 (N_2333,N_1971,N_1250);
or U2334 (N_2334,N_1004,N_1933);
or U2335 (N_2335,N_1675,N_1825);
nand U2336 (N_2336,N_1484,N_1054);
xnor U2337 (N_2337,N_1949,N_1512);
nand U2338 (N_2338,N_1316,N_1782);
and U2339 (N_2339,N_1985,N_1491);
and U2340 (N_2340,N_1997,N_1341);
or U2341 (N_2341,N_1632,N_1148);
xnor U2342 (N_2342,N_1444,N_1737);
xnor U2343 (N_2343,N_1356,N_1751);
xnor U2344 (N_2344,N_1552,N_1856);
and U2345 (N_2345,N_1626,N_1622);
xnor U2346 (N_2346,N_1734,N_1754);
xnor U2347 (N_2347,N_1948,N_1595);
nor U2348 (N_2348,N_1426,N_1679);
or U2349 (N_2349,N_1353,N_1116);
and U2350 (N_2350,N_1766,N_1349);
nand U2351 (N_2351,N_1486,N_1382);
and U2352 (N_2352,N_1181,N_1273);
xnor U2353 (N_2353,N_1256,N_1896);
or U2354 (N_2354,N_1364,N_1944);
nand U2355 (N_2355,N_1548,N_1163);
and U2356 (N_2356,N_1261,N_1157);
nand U2357 (N_2357,N_1775,N_1465);
xor U2358 (N_2358,N_1310,N_1841);
xnor U2359 (N_2359,N_1284,N_1628);
and U2360 (N_2360,N_1748,N_1247);
nor U2361 (N_2361,N_1562,N_1422);
nand U2362 (N_2362,N_1042,N_1330);
nor U2363 (N_2363,N_1717,N_1612);
or U2364 (N_2364,N_1528,N_1240);
and U2365 (N_2365,N_1208,N_1614);
or U2366 (N_2366,N_1096,N_1700);
and U2367 (N_2367,N_1479,N_1130);
and U2368 (N_2368,N_1630,N_1542);
nand U2369 (N_2369,N_1876,N_1488);
and U2370 (N_2370,N_1813,N_1224);
or U2371 (N_2371,N_1795,N_1462);
nand U2372 (N_2372,N_1125,N_1637);
or U2373 (N_2373,N_1742,N_1879);
or U2374 (N_2374,N_1867,N_1071);
xnor U2375 (N_2375,N_1031,N_1006);
xor U2376 (N_2376,N_1000,N_1295);
or U2377 (N_2377,N_1885,N_1459);
and U2378 (N_2378,N_1550,N_1786);
nand U2379 (N_2379,N_1454,N_1490);
and U2380 (N_2380,N_1347,N_1973);
nor U2381 (N_2381,N_1471,N_1384);
or U2382 (N_2382,N_1402,N_1883);
nor U2383 (N_2383,N_1658,N_1803);
or U2384 (N_2384,N_1151,N_1294);
xor U2385 (N_2385,N_1478,N_1998);
xor U2386 (N_2386,N_1950,N_1421);
nand U2387 (N_2387,N_1524,N_1892);
nor U2388 (N_2388,N_1547,N_1361);
xor U2389 (N_2389,N_1231,N_1070);
or U2390 (N_2390,N_1475,N_1587);
or U2391 (N_2391,N_1141,N_1934);
and U2392 (N_2392,N_1306,N_1968);
or U2393 (N_2393,N_1945,N_1777);
and U2394 (N_2394,N_1391,N_1146);
nor U2395 (N_2395,N_1451,N_1327);
nand U2396 (N_2396,N_1298,N_1377);
nor U2397 (N_2397,N_1767,N_1067);
nor U2398 (N_2398,N_1598,N_1818);
xnor U2399 (N_2399,N_1635,N_1083);
nand U2400 (N_2400,N_1293,N_1420);
xnor U2401 (N_2401,N_1545,N_1604);
xnor U2402 (N_2402,N_1676,N_1336);
nand U2403 (N_2403,N_1225,N_1404);
or U2404 (N_2404,N_1122,N_1544);
nor U2405 (N_2405,N_1312,N_1075);
or U2406 (N_2406,N_1873,N_1917);
or U2407 (N_2407,N_1366,N_1684);
xnor U2408 (N_2408,N_1092,N_1978);
nand U2409 (N_2409,N_1326,N_1609);
xor U2410 (N_2410,N_1408,N_1663);
nor U2411 (N_2411,N_1155,N_1797);
and U2412 (N_2412,N_1589,N_1325);
nand U2413 (N_2413,N_1145,N_1413);
and U2414 (N_2414,N_1608,N_1072);
nor U2415 (N_2415,N_1913,N_1498);
nand U2416 (N_2416,N_1248,N_1932);
or U2417 (N_2417,N_1328,N_1138);
and U2418 (N_2418,N_1807,N_1394);
nor U2419 (N_2419,N_1505,N_1811);
xnor U2420 (N_2420,N_1955,N_1393);
or U2421 (N_2421,N_1549,N_1129);
and U2422 (N_2422,N_1497,N_1792);
nor U2423 (N_2423,N_1880,N_1696);
nor U2424 (N_2424,N_1241,N_1669);
xor U2425 (N_2425,N_1666,N_1449);
xnor U2426 (N_2426,N_1639,N_1638);
or U2427 (N_2427,N_1723,N_1794);
and U2428 (N_2428,N_1822,N_1855);
nand U2429 (N_2429,N_1149,N_1342);
nor U2430 (N_2430,N_1424,N_1569);
xor U2431 (N_2431,N_1600,N_1477);
nand U2432 (N_2432,N_1405,N_1986);
or U2433 (N_2433,N_1974,N_1463);
nor U2434 (N_2434,N_1169,N_1787);
or U2435 (N_2435,N_1685,N_1403);
nor U2436 (N_2436,N_1362,N_1750);
or U2437 (N_2437,N_1280,N_1142);
and U2438 (N_2438,N_1519,N_1055);
xor U2439 (N_2439,N_1906,N_1659);
or U2440 (N_2440,N_1068,N_1011);
nor U2441 (N_2441,N_1809,N_1038);
and U2442 (N_2442,N_1789,N_1515);
and U2443 (N_2443,N_1993,N_1610);
or U2444 (N_2444,N_1893,N_1111);
nand U2445 (N_2445,N_1409,N_1914);
or U2446 (N_2446,N_1852,N_1289);
or U2447 (N_2447,N_1299,N_1016);
nor U2448 (N_2448,N_1845,N_1099);
xor U2449 (N_2449,N_1784,N_1922);
xor U2450 (N_2450,N_1960,N_1137);
and U2451 (N_2451,N_1527,N_1332);
or U2452 (N_2452,N_1735,N_1425);
or U2453 (N_2453,N_1243,N_1277);
xnor U2454 (N_2454,N_1200,N_1606);
xnor U2455 (N_2455,N_1367,N_1081);
nand U2456 (N_2456,N_1537,N_1201);
or U2457 (N_2457,N_1079,N_1901);
nand U2458 (N_2458,N_1113,N_1557);
or U2459 (N_2459,N_1177,N_1511);
nand U2460 (N_2460,N_1418,N_1021);
and U2461 (N_2461,N_1051,N_1218);
nand U2462 (N_2462,N_1417,N_1268);
nor U2463 (N_2463,N_1594,N_1290);
xor U2464 (N_2464,N_1022,N_1781);
and U2465 (N_2465,N_1992,N_1025);
xor U2466 (N_2466,N_1041,N_1432);
and U2467 (N_2467,N_1947,N_1066);
and U2468 (N_2468,N_1687,N_1919);
or U2469 (N_2469,N_1464,N_1656);
or U2470 (N_2470,N_1899,N_1555);
and U2471 (N_2471,N_1274,N_1761);
xor U2472 (N_2472,N_1365,N_1401);
and U2473 (N_2473,N_1144,N_1712);
and U2474 (N_2474,N_1495,N_1821);
nor U2475 (N_2475,N_1533,N_1183);
nor U2476 (N_2476,N_1531,N_1563);
nor U2477 (N_2477,N_1525,N_1244);
nor U2478 (N_2478,N_1166,N_1152);
xnor U2479 (N_2479,N_1859,N_1719);
or U2480 (N_2480,N_1230,N_1046);
or U2481 (N_2481,N_1175,N_1430);
and U2482 (N_2482,N_1371,N_1959);
or U2483 (N_2483,N_1897,N_1857);
nand U2484 (N_2484,N_1583,N_1894);
and U2485 (N_2485,N_1624,N_1286);
xnor U2486 (N_2486,N_1871,N_1689);
and U2487 (N_2487,N_1128,N_1266);
nand U2488 (N_2488,N_1935,N_1962);
nand U2489 (N_2489,N_1987,N_1558);
nor U2490 (N_2490,N_1534,N_1412);
nor U2491 (N_2491,N_1900,N_1194);
xor U2492 (N_2492,N_1100,N_1219);
nor U2493 (N_2493,N_1419,N_1411);
nand U2494 (N_2494,N_1466,N_1005);
or U2495 (N_2495,N_1704,N_1938);
nor U2496 (N_2496,N_1048,N_1756);
nand U2497 (N_2497,N_1844,N_1909);
and U2498 (N_2498,N_1727,N_1440);
nor U2499 (N_2499,N_1446,N_1698);
nor U2500 (N_2500,N_1079,N_1515);
nor U2501 (N_2501,N_1960,N_1701);
and U2502 (N_2502,N_1007,N_1233);
nand U2503 (N_2503,N_1620,N_1165);
xor U2504 (N_2504,N_1245,N_1570);
or U2505 (N_2505,N_1784,N_1964);
nand U2506 (N_2506,N_1946,N_1273);
or U2507 (N_2507,N_1600,N_1793);
nand U2508 (N_2508,N_1829,N_1710);
xnor U2509 (N_2509,N_1677,N_1790);
nor U2510 (N_2510,N_1685,N_1589);
nor U2511 (N_2511,N_1159,N_1251);
or U2512 (N_2512,N_1860,N_1176);
nor U2513 (N_2513,N_1015,N_1398);
or U2514 (N_2514,N_1329,N_1520);
xnor U2515 (N_2515,N_1357,N_1870);
and U2516 (N_2516,N_1708,N_1278);
nor U2517 (N_2517,N_1129,N_1330);
xnor U2518 (N_2518,N_1862,N_1503);
and U2519 (N_2519,N_1819,N_1936);
or U2520 (N_2520,N_1252,N_1836);
xor U2521 (N_2521,N_1992,N_1133);
xnor U2522 (N_2522,N_1423,N_1823);
nand U2523 (N_2523,N_1504,N_1892);
xor U2524 (N_2524,N_1318,N_1022);
nand U2525 (N_2525,N_1822,N_1955);
xor U2526 (N_2526,N_1014,N_1863);
xor U2527 (N_2527,N_1591,N_1391);
xor U2528 (N_2528,N_1928,N_1226);
xor U2529 (N_2529,N_1950,N_1502);
xnor U2530 (N_2530,N_1839,N_1581);
nand U2531 (N_2531,N_1237,N_1174);
or U2532 (N_2532,N_1222,N_1819);
nand U2533 (N_2533,N_1151,N_1789);
nand U2534 (N_2534,N_1625,N_1830);
and U2535 (N_2535,N_1953,N_1349);
nor U2536 (N_2536,N_1001,N_1224);
nand U2537 (N_2537,N_1783,N_1876);
nand U2538 (N_2538,N_1359,N_1858);
nor U2539 (N_2539,N_1700,N_1709);
and U2540 (N_2540,N_1762,N_1599);
and U2541 (N_2541,N_1548,N_1028);
nand U2542 (N_2542,N_1950,N_1899);
nor U2543 (N_2543,N_1155,N_1452);
or U2544 (N_2544,N_1391,N_1743);
xnor U2545 (N_2545,N_1246,N_1248);
nor U2546 (N_2546,N_1879,N_1386);
nor U2547 (N_2547,N_1324,N_1174);
nor U2548 (N_2548,N_1439,N_1834);
or U2549 (N_2549,N_1532,N_1914);
xnor U2550 (N_2550,N_1206,N_1128);
and U2551 (N_2551,N_1064,N_1846);
and U2552 (N_2552,N_1432,N_1851);
or U2553 (N_2553,N_1741,N_1533);
nand U2554 (N_2554,N_1342,N_1264);
nand U2555 (N_2555,N_1448,N_1471);
nor U2556 (N_2556,N_1040,N_1208);
nand U2557 (N_2557,N_1406,N_1704);
nand U2558 (N_2558,N_1485,N_1673);
nand U2559 (N_2559,N_1762,N_1723);
and U2560 (N_2560,N_1817,N_1416);
and U2561 (N_2561,N_1665,N_1794);
nor U2562 (N_2562,N_1927,N_1068);
xnor U2563 (N_2563,N_1820,N_1973);
and U2564 (N_2564,N_1725,N_1113);
and U2565 (N_2565,N_1557,N_1469);
and U2566 (N_2566,N_1001,N_1325);
nor U2567 (N_2567,N_1016,N_1699);
nand U2568 (N_2568,N_1948,N_1807);
or U2569 (N_2569,N_1037,N_1811);
xnor U2570 (N_2570,N_1222,N_1593);
xnor U2571 (N_2571,N_1756,N_1607);
nand U2572 (N_2572,N_1653,N_1367);
and U2573 (N_2573,N_1637,N_1429);
xnor U2574 (N_2574,N_1725,N_1147);
xnor U2575 (N_2575,N_1291,N_1697);
xnor U2576 (N_2576,N_1401,N_1800);
or U2577 (N_2577,N_1060,N_1849);
nor U2578 (N_2578,N_1467,N_1353);
xor U2579 (N_2579,N_1476,N_1426);
or U2580 (N_2580,N_1417,N_1114);
nor U2581 (N_2581,N_1611,N_1809);
and U2582 (N_2582,N_1359,N_1397);
or U2583 (N_2583,N_1885,N_1184);
nor U2584 (N_2584,N_1856,N_1366);
and U2585 (N_2585,N_1101,N_1149);
nor U2586 (N_2586,N_1716,N_1274);
xnor U2587 (N_2587,N_1597,N_1196);
nand U2588 (N_2588,N_1422,N_1827);
nand U2589 (N_2589,N_1614,N_1342);
nand U2590 (N_2590,N_1767,N_1670);
xnor U2591 (N_2591,N_1906,N_1856);
nor U2592 (N_2592,N_1562,N_1520);
nand U2593 (N_2593,N_1680,N_1311);
and U2594 (N_2594,N_1410,N_1302);
nor U2595 (N_2595,N_1819,N_1217);
nor U2596 (N_2596,N_1656,N_1897);
and U2597 (N_2597,N_1915,N_1995);
or U2598 (N_2598,N_1378,N_1324);
or U2599 (N_2599,N_1194,N_1984);
and U2600 (N_2600,N_1420,N_1485);
and U2601 (N_2601,N_1257,N_1522);
nand U2602 (N_2602,N_1209,N_1534);
nand U2603 (N_2603,N_1982,N_1179);
nand U2604 (N_2604,N_1394,N_1020);
xor U2605 (N_2605,N_1413,N_1086);
or U2606 (N_2606,N_1507,N_1372);
nand U2607 (N_2607,N_1088,N_1403);
xor U2608 (N_2608,N_1295,N_1598);
xnor U2609 (N_2609,N_1592,N_1940);
xor U2610 (N_2610,N_1598,N_1607);
nor U2611 (N_2611,N_1478,N_1519);
nand U2612 (N_2612,N_1523,N_1391);
and U2613 (N_2613,N_1430,N_1722);
nand U2614 (N_2614,N_1339,N_1960);
and U2615 (N_2615,N_1448,N_1773);
xor U2616 (N_2616,N_1255,N_1406);
xnor U2617 (N_2617,N_1595,N_1219);
nor U2618 (N_2618,N_1655,N_1148);
xnor U2619 (N_2619,N_1407,N_1435);
or U2620 (N_2620,N_1816,N_1065);
xnor U2621 (N_2621,N_1718,N_1818);
nor U2622 (N_2622,N_1417,N_1129);
and U2623 (N_2623,N_1942,N_1557);
or U2624 (N_2624,N_1908,N_1295);
or U2625 (N_2625,N_1552,N_1559);
nand U2626 (N_2626,N_1600,N_1806);
and U2627 (N_2627,N_1330,N_1599);
nand U2628 (N_2628,N_1801,N_1934);
nand U2629 (N_2629,N_1428,N_1175);
nand U2630 (N_2630,N_1890,N_1255);
nor U2631 (N_2631,N_1763,N_1946);
and U2632 (N_2632,N_1641,N_1783);
and U2633 (N_2633,N_1314,N_1964);
or U2634 (N_2634,N_1927,N_1839);
nor U2635 (N_2635,N_1879,N_1903);
and U2636 (N_2636,N_1368,N_1262);
and U2637 (N_2637,N_1812,N_1685);
or U2638 (N_2638,N_1949,N_1185);
nor U2639 (N_2639,N_1461,N_1986);
nor U2640 (N_2640,N_1095,N_1375);
and U2641 (N_2641,N_1542,N_1726);
or U2642 (N_2642,N_1534,N_1128);
and U2643 (N_2643,N_1687,N_1769);
xnor U2644 (N_2644,N_1452,N_1788);
nor U2645 (N_2645,N_1836,N_1529);
nand U2646 (N_2646,N_1339,N_1334);
xnor U2647 (N_2647,N_1625,N_1664);
nor U2648 (N_2648,N_1715,N_1593);
nand U2649 (N_2649,N_1442,N_1084);
nor U2650 (N_2650,N_1427,N_1149);
or U2651 (N_2651,N_1937,N_1323);
nor U2652 (N_2652,N_1783,N_1958);
or U2653 (N_2653,N_1731,N_1716);
and U2654 (N_2654,N_1017,N_1417);
and U2655 (N_2655,N_1884,N_1935);
nor U2656 (N_2656,N_1837,N_1246);
nor U2657 (N_2657,N_1647,N_1644);
xor U2658 (N_2658,N_1439,N_1410);
xor U2659 (N_2659,N_1089,N_1400);
and U2660 (N_2660,N_1482,N_1402);
and U2661 (N_2661,N_1413,N_1201);
nor U2662 (N_2662,N_1831,N_1860);
xor U2663 (N_2663,N_1102,N_1262);
nor U2664 (N_2664,N_1227,N_1269);
nand U2665 (N_2665,N_1972,N_1031);
and U2666 (N_2666,N_1125,N_1684);
nor U2667 (N_2667,N_1521,N_1209);
and U2668 (N_2668,N_1836,N_1800);
or U2669 (N_2669,N_1568,N_1462);
or U2670 (N_2670,N_1503,N_1856);
or U2671 (N_2671,N_1702,N_1392);
or U2672 (N_2672,N_1203,N_1491);
xnor U2673 (N_2673,N_1118,N_1063);
nor U2674 (N_2674,N_1017,N_1630);
nor U2675 (N_2675,N_1345,N_1908);
nor U2676 (N_2676,N_1272,N_1610);
xor U2677 (N_2677,N_1860,N_1819);
and U2678 (N_2678,N_1357,N_1318);
xor U2679 (N_2679,N_1675,N_1061);
xnor U2680 (N_2680,N_1774,N_1476);
and U2681 (N_2681,N_1713,N_1273);
nor U2682 (N_2682,N_1829,N_1928);
nor U2683 (N_2683,N_1054,N_1889);
nand U2684 (N_2684,N_1320,N_1285);
nand U2685 (N_2685,N_1323,N_1716);
or U2686 (N_2686,N_1043,N_1254);
nor U2687 (N_2687,N_1362,N_1090);
nor U2688 (N_2688,N_1276,N_1705);
and U2689 (N_2689,N_1324,N_1783);
xor U2690 (N_2690,N_1164,N_1390);
nor U2691 (N_2691,N_1774,N_1091);
nor U2692 (N_2692,N_1783,N_1130);
nand U2693 (N_2693,N_1178,N_1698);
nor U2694 (N_2694,N_1229,N_1327);
or U2695 (N_2695,N_1688,N_1466);
or U2696 (N_2696,N_1119,N_1673);
xor U2697 (N_2697,N_1147,N_1918);
or U2698 (N_2698,N_1858,N_1362);
or U2699 (N_2699,N_1576,N_1943);
nand U2700 (N_2700,N_1784,N_1057);
xor U2701 (N_2701,N_1129,N_1203);
xnor U2702 (N_2702,N_1104,N_1499);
nand U2703 (N_2703,N_1071,N_1383);
nand U2704 (N_2704,N_1535,N_1620);
xnor U2705 (N_2705,N_1596,N_1093);
or U2706 (N_2706,N_1215,N_1815);
nand U2707 (N_2707,N_1644,N_1650);
nor U2708 (N_2708,N_1335,N_1679);
or U2709 (N_2709,N_1487,N_1406);
or U2710 (N_2710,N_1844,N_1253);
and U2711 (N_2711,N_1257,N_1371);
or U2712 (N_2712,N_1013,N_1085);
xor U2713 (N_2713,N_1652,N_1427);
xor U2714 (N_2714,N_1122,N_1599);
and U2715 (N_2715,N_1414,N_1127);
or U2716 (N_2716,N_1305,N_1747);
and U2717 (N_2717,N_1569,N_1046);
xor U2718 (N_2718,N_1540,N_1698);
and U2719 (N_2719,N_1645,N_1913);
nand U2720 (N_2720,N_1038,N_1047);
or U2721 (N_2721,N_1874,N_1520);
nand U2722 (N_2722,N_1926,N_1196);
nand U2723 (N_2723,N_1401,N_1981);
or U2724 (N_2724,N_1060,N_1385);
or U2725 (N_2725,N_1250,N_1696);
and U2726 (N_2726,N_1474,N_1988);
nor U2727 (N_2727,N_1212,N_1657);
xor U2728 (N_2728,N_1689,N_1698);
and U2729 (N_2729,N_1872,N_1490);
nor U2730 (N_2730,N_1555,N_1370);
nand U2731 (N_2731,N_1137,N_1424);
nor U2732 (N_2732,N_1312,N_1384);
or U2733 (N_2733,N_1780,N_1995);
nand U2734 (N_2734,N_1224,N_1466);
nor U2735 (N_2735,N_1699,N_1232);
and U2736 (N_2736,N_1717,N_1407);
and U2737 (N_2737,N_1575,N_1463);
and U2738 (N_2738,N_1586,N_1473);
xor U2739 (N_2739,N_1405,N_1870);
or U2740 (N_2740,N_1918,N_1116);
xor U2741 (N_2741,N_1565,N_1483);
nand U2742 (N_2742,N_1833,N_1375);
or U2743 (N_2743,N_1466,N_1415);
xnor U2744 (N_2744,N_1606,N_1290);
xor U2745 (N_2745,N_1460,N_1373);
and U2746 (N_2746,N_1107,N_1928);
or U2747 (N_2747,N_1005,N_1655);
nand U2748 (N_2748,N_1293,N_1262);
or U2749 (N_2749,N_1859,N_1502);
and U2750 (N_2750,N_1151,N_1363);
nand U2751 (N_2751,N_1382,N_1186);
and U2752 (N_2752,N_1297,N_1298);
or U2753 (N_2753,N_1795,N_1365);
nand U2754 (N_2754,N_1124,N_1728);
and U2755 (N_2755,N_1708,N_1237);
and U2756 (N_2756,N_1538,N_1449);
and U2757 (N_2757,N_1009,N_1708);
nor U2758 (N_2758,N_1857,N_1337);
nor U2759 (N_2759,N_1989,N_1171);
and U2760 (N_2760,N_1860,N_1888);
or U2761 (N_2761,N_1114,N_1986);
xnor U2762 (N_2762,N_1237,N_1952);
xor U2763 (N_2763,N_1254,N_1845);
nor U2764 (N_2764,N_1569,N_1485);
xor U2765 (N_2765,N_1761,N_1642);
nand U2766 (N_2766,N_1481,N_1151);
nor U2767 (N_2767,N_1503,N_1264);
nor U2768 (N_2768,N_1576,N_1339);
nand U2769 (N_2769,N_1666,N_1103);
nor U2770 (N_2770,N_1039,N_1364);
and U2771 (N_2771,N_1238,N_1946);
or U2772 (N_2772,N_1416,N_1271);
and U2773 (N_2773,N_1460,N_1087);
nor U2774 (N_2774,N_1256,N_1722);
nand U2775 (N_2775,N_1031,N_1738);
and U2776 (N_2776,N_1137,N_1596);
nand U2777 (N_2777,N_1590,N_1731);
and U2778 (N_2778,N_1836,N_1182);
or U2779 (N_2779,N_1483,N_1684);
nor U2780 (N_2780,N_1857,N_1159);
nand U2781 (N_2781,N_1138,N_1136);
nor U2782 (N_2782,N_1450,N_1096);
nand U2783 (N_2783,N_1293,N_1811);
nor U2784 (N_2784,N_1222,N_1732);
xnor U2785 (N_2785,N_1723,N_1055);
xnor U2786 (N_2786,N_1642,N_1448);
xor U2787 (N_2787,N_1010,N_1191);
nand U2788 (N_2788,N_1938,N_1999);
and U2789 (N_2789,N_1824,N_1270);
nor U2790 (N_2790,N_1571,N_1303);
xor U2791 (N_2791,N_1884,N_1663);
nand U2792 (N_2792,N_1164,N_1791);
xnor U2793 (N_2793,N_1015,N_1020);
nand U2794 (N_2794,N_1815,N_1338);
xnor U2795 (N_2795,N_1914,N_1554);
xor U2796 (N_2796,N_1074,N_1661);
or U2797 (N_2797,N_1263,N_1044);
xnor U2798 (N_2798,N_1079,N_1910);
or U2799 (N_2799,N_1452,N_1607);
or U2800 (N_2800,N_1089,N_1267);
nor U2801 (N_2801,N_1875,N_1688);
xnor U2802 (N_2802,N_1537,N_1105);
and U2803 (N_2803,N_1469,N_1346);
or U2804 (N_2804,N_1247,N_1634);
or U2805 (N_2805,N_1227,N_1757);
and U2806 (N_2806,N_1925,N_1686);
nand U2807 (N_2807,N_1516,N_1889);
xor U2808 (N_2808,N_1829,N_1850);
and U2809 (N_2809,N_1259,N_1247);
nor U2810 (N_2810,N_1769,N_1592);
xor U2811 (N_2811,N_1861,N_1414);
or U2812 (N_2812,N_1844,N_1511);
nor U2813 (N_2813,N_1221,N_1694);
xor U2814 (N_2814,N_1573,N_1811);
nand U2815 (N_2815,N_1016,N_1382);
xnor U2816 (N_2816,N_1884,N_1721);
nor U2817 (N_2817,N_1099,N_1694);
and U2818 (N_2818,N_1016,N_1094);
and U2819 (N_2819,N_1997,N_1584);
nand U2820 (N_2820,N_1442,N_1293);
or U2821 (N_2821,N_1232,N_1216);
or U2822 (N_2822,N_1610,N_1595);
xor U2823 (N_2823,N_1838,N_1067);
xnor U2824 (N_2824,N_1794,N_1973);
xor U2825 (N_2825,N_1792,N_1999);
and U2826 (N_2826,N_1335,N_1867);
nor U2827 (N_2827,N_1960,N_1489);
xor U2828 (N_2828,N_1697,N_1899);
nand U2829 (N_2829,N_1173,N_1139);
or U2830 (N_2830,N_1673,N_1092);
xnor U2831 (N_2831,N_1827,N_1577);
nand U2832 (N_2832,N_1817,N_1121);
nor U2833 (N_2833,N_1378,N_1710);
and U2834 (N_2834,N_1050,N_1151);
or U2835 (N_2835,N_1139,N_1802);
nand U2836 (N_2836,N_1074,N_1426);
xor U2837 (N_2837,N_1194,N_1991);
nand U2838 (N_2838,N_1448,N_1569);
nand U2839 (N_2839,N_1408,N_1274);
xor U2840 (N_2840,N_1570,N_1822);
or U2841 (N_2841,N_1649,N_1272);
or U2842 (N_2842,N_1228,N_1233);
or U2843 (N_2843,N_1466,N_1619);
nand U2844 (N_2844,N_1533,N_1222);
xnor U2845 (N_2845,N_1115,N_1282);
nand U2846 (N_2846,N_1250,N_1098);
or U2847 (N_2847,N_1931,N_1944);
and U2848 (N_2848,N_1053,N_1591);
nand U2849 (N_2849,N_1058,N_1395);
nand U2850 (N_2850,N_1215,N_1140);
or U2851 (N_2851,N_1989,N_1235);
or U2852 (N_2852,N_1829,N_1315);
nand U2853 (N_2853,N_1948,N_1382);
nand U2854 (N_2854,N_1115,N_1864);
or U2855 (N_2855,N_1747,N_1116);
or U2856 (N_2856,N_1018,N_1732);
xnor U2857 (N_2857,N_1787,N_1811);
or U2858 (N_2858,N_1724,N_1233);
and U2859 (N_2859,N_1438,N_1304);
nor U2860 (N_2860,N_1516,N_1896);
and U2861 (N_2861,N_1530,N_1754);
nand U2862 (N_2862,N_1508,N_1775);
xor U2863 (N_2863,N_1573,N_1475);
xor U2864 (N_2864,N_1283,N_1821);
nor U2865 (N_2865,N_1342,N_1566);
nor U2866 (N_2866,N_1523,N_1272);
nand U2867 (N_2867,N_1289,N_1797);
nor U2868 (N_2868,N_1140,N_1647);
nor U2869 (N_2869,N_1223,N_1204);
nor U2870 (N_2870,N_1961,N_1025);
xor U2871 (N_2871,N_1398,N_1204);
nor U2872 (N_2872,N_1701,N_1462);
or U2873 (N_2873,N_1208,N_1266);
and U2874 (N_2874,N_1281,N_1972);
nor U2875 (N_2875,N_1509,N_1890);
xor U2876 (N_2876,N_1743,N_1918);
nand U2877 (N_2877,N_1996,N_1928);
xnor U2878 (N_2878,N_1327,N_1994);
or U2879 (N_2879,N_1006,N_1760);
nand U2880 (N_2880,N_1591,N_1138);
or U2881 (N_2881,N_1989,N_1975);
nor U2882 (N_2882,N_1302,N_1553);
or U2883 (N_2883,N_1281,N_1197);
nor U2884 (N_2884,N_1339,N_1792);
or U2885 (N_2885,N_1072,N_1305);
or U2886 (N_2886,N_1417,N_1898);
nor U2887 (N_2887,N_1950,N_1563);
and U2888 (N_2888,N_1064,N_1070);
xor U2889 (N_2889,N_1919,N_1181);
nand U2890 (N_2890,N_1405,N_1587);
or U2891 (N_2891,N_1474,N_1692);
and U2892 (N_2892,N_1104,N_1050);
or U2893 (N_2893,N_1118,N_1779);
xnor U2894 (N_2894,N_1958,N_1366);
and U2895 (N_2895,N_1338,N_1402);
nor U2896 (N_2896,N_1143,N_1453);
and U2897 (N_2897,N_1023,N_1454);
nand U2898 (N_2898,N_1899,N_1948);
nand U2899 (N_2899,N_1299,N_1358);
or U2900 (N_2900,N_1729,N_1857);
nand U2901 (N_2901,N_1292,N_1160);
or U2902 (N_2902,N_1140,N_1306);
nor U2903 (N_2903,N_1776,N_1462);
xnor U2904 (N_2904,N_1087,N_1997);
and U2905 (N_2905,N_1347,N_1570);
xor U2906 (N_2906,N_1636,N_1114);
nor U2907 (N_2907,N_1071,N_1229);
xnor U2908 (N_2908,N_1341,N_1603);
nor U2909 (N_2909,N_1967,N_1878);
xnor U2910 (N_2910,N_1827,N_1404);
or U2911 (N_2911,N_1656,N_1649);
and U2912 (N_2912,N_1690,N_1732);
or U2913 (N_2913,N_1915,N_1579);
nand U2914 (N_2914,N_1625,N_1707);
nand U2915 (N_2915,N_1114,N_1825);
xor U2916 (N_2916,N_1288,N_1499);
xor U2917 (N_2917,N_1442,N_1068);
and U2918 (N_2918,N_1106,N_1072);
nand U2919 (N_2919,N_1809,N_1408);
xnor U2920 (N_2920,N_1334,N_1532);
nand U2921 (N_2921,N_1041,N_1164);
nor U2922 (N_2922,N_1361,N_1808);
xor U2923 (N_2923,N_1317,N_1013);
and U2924 (N_2924,N_1422,N_1841);
nand U2925 (N_2925,N_1900,N_1190);
xnor U2926 (N_2926,N_1853,N_1824);
nor U2927 (N_2927,N_1914,N_1700);
xnor U2928 (N_2928,N_1627,N_1987);
nor U2929 (N_2929,N_1454,N_1644);
nand U2930 (N_2930,N_1479,N_1645);
xnor U2931 (N_2931,N_1924,N_1893);
nor U2932 (N_2932,N_1732,N_1362);
and U2933 (N_2933,N_1433,N_1034);
or U2934 (N_2934,N_1072,N_1686);
and U2935 (N_2935,N_1481,N_1209);
nand U2936 (N_2936,N_1921,N_1043);
and U2937 (N_2937,N_1898,N_1209);
nor U2938 (N_2938,N_1227,N_1913);
xor U2939 (N_2939,N_1672,N_1492);
nand U2940 (N_2940,N_1696,N_1376);
nand U2941 (N_2941,N_1411,N_1644);
and U2942 (N_2942,N_1010,N_1229);
or U2943 (N_2943,N_1717,N_1034);
xor U2944 (N_2944,N_1074,N_1632);
or U2945 (N_2945,N_1443,N_1147);
nand U2946 (N_2946,N_1217,N_1054);
xor U2947 (N_2947,N_1736,N_1176);
nor U2948 (N_2948,N_1465,N_1339);
nor U2949 (N_2949,N_1813,N_1081);
or U2950 (N_2950,N_1318,N_1319);
xnor U2951 (N_2951,N_1578,N_1699);
or U2952 (N_2952,N_1675,N_1695);
nor U2953 (N_2953,N_1308,N_1304);
xor U2954 (N_2954,N_1144,N_1592);
nand U2955 (N_2955,N_1852,N_1628);
or U2956 (N_2956,N_1501,N_1124);
and U2957 (N_2957,N_1316,N_1780);
xor U2958 (N_2958,N_1387,N_1089);
and U2959 (N_2959,N_1920,N_1917);
or U2960 (N_2960,N_1027,N_1058);
and U2961 (N_2961,N_1157,N_1168);
nor U2962 (N_2962,N_1426,N_1743);
nor U2963 (N_2963,N_1200,N_1347);
and U2964 (N_2964,N_1194,N_1814);
nand U2965 (N_2965,N_1881,N_1202);
nor U2966 (N_2966,N_1135,N_1957);
nor U2967 (N_2967,N_1300,N_1353);
or U2968 (N_2968,N_1160,N_1779);
nor U2969 (N_2969,N_1175,N_1242);
nand U2970 (N_2970,N_1243,N_1357);
nand U2971 (N_2971,N_1336,N_1498);
and U2972 (N_2972,N_1128,N_1487);
and U2973 (N_2973,N_1295,N_1131);
or U2974 (N_2974,N_1597,N_1585);
and U2975 (N_2975,N_1190,N_1723);
nand U2976 (N_2976,N_1492,N_1037);
nand U2977 (N_2977,N_1876,N_1460);
xor U2978 (N_2978,N_1630,N_1819);
nand U2979 (N_2979,N_1363,N_1312);
nand U2980 (N_2980,N_1970,N_1773);
xor U2981 (N_2981,N_1921,N_1436);
xnor U2982 (N_2982,N_1564,N_1658);
nand U2983 (N_2983,N_1213,N_1198);
nand U2984 (N_2984,N_1583,N_1017);
nand U2985 (N_2985,N_1053,N_1483);
nand U2986 (N_2986,N_1922,N_1804);
nand U2987 (N_2987,N_1891,N_1174);
nand U2988 (N_2988,N_1019,N_1524);
and U2989 (N_2989,N_1414,N_1479);
nor U2990 (N_2990,N_1736,N_1952);
or U2991 (N_2991,N_1109,N_1099);
nor U2992 (N_2992,N_1692,N_1110);
or U2993 (N_2993,N_1933,N_1139);
or U2994 (N_2994,N_1363,N_1626);
xnor U2995 (N_2995,N_1609,N_1744);
xnor U2996 (N_2996,N_1733,N_1222);
nor U2997 (N_2997,N_1784,N_1972);
nor U2998 (N_2998,N_1200,N_1359);
nand U2999 (N_2999,N_1085,N_1263);
or U3000 (N_3000,N_2683,N_2527);
or U3001 (N_3001,N_2100,N_2994);
or U3002 (N_3002,N_2656,N_2478);
nor U3003 (N_3003,N_2918,N_2812);
xnor U3004 (N_3004,N_2121,N_2090);
xnor U3005 (N_3005,N_2968,N_2707);
and U3006 (N_3006,N_2752,N_2038);
nor U3007 (N_3007,N_2792,N_2068);
nor U3008 (N_3008,N_2980,N_2229);
xor U3009 (N_3009,N_2426,N_2951);
nor U3010 (N_3010,N_2678,N_2954);
nor U3011 (N_3011,N_2844,N_2541);
nand U3012 (N_3012,N_2282,N_2967);
nand U3013 (N_3013,N_2686,N_2446);
nor U3014 (N_3014,N_2636,N_2771);
xnor U3015 (N_3015,N_2999,N_2970);
xnor U3016 (N_3016,N_2084,N_2919);
nor U3017 (N_3017,N_2785,N_2033);
or U3018 (N_3018,N_2168,N_2095);
nor U3019 (N_3019,N_2809,N_2922);
nor U3020 (N_3020,N_2267,N_2709);
nand U3021 (N_3021,N_2540,N_2330);
xnor U3022 (N_3022,N_2895,N_2059);
nand U3023 (N_3023,N_2646,N_2706);
or U3024 (N_3024,N_2515,N_2816);
or U3025 (N_3025,N_2410,N_2164);
and U3026 (N_3026,N_2620,N_2714);
nand U3027 (N_3027,N_2213,N_2116);
nor U3028 (N_3028,N_2754,N_2030);
and U3029 (N_3029,N_2218,N_2206);
and U3030 (N_3030,N_2740,N_2089);
nand U3031 (N_3031,N_2931,N_2603);
or U3032 (N_3032,N_2634,N_2864);
nor U3033 (N_3033,N_2657,N_2648);
nor U3034 (N_3034,N_2998,N_2817);
or U3035 (N_3035,N_2913,N_2061);
nand U3036 (N_3036,N_2548,N_2534);
and U3037 (N_3037,N_2039,N_2940);
nor U3038 (N_3038,N_2256,N_2764);
xnor U3039 (N_3039,N_2856,N_2141);
or U3040 (N_3040,N_2961,N_2641);
and U3041 (N_3041,N_2893,N_2973);
xnor U3042 (N_3042,N_2367,N_2911);
or U3043 (N_3043,N_2437,N_2494);
or U3044 (N_3044,N_2232,N_2081);
nand U3045 (N_3045,N_2445,N_2741);
nand U3046 (N_3046,N_2926,N_2397);
nor U3047 (N_3047,N_2123,N_2680);
or U3048 (N_3048,N_2717,N_2112);
xnor U3049 (N_3049,N_2079,N_2403);
nor U3050 (N_3050,N_2526,N_2246);
nand U3051 (N_3051,N_2828,N_2052);
nand U3052 (N_3052,N_2904,N_2131);
or U3053 (N_3053,N_2133,N_2547);
or U3054 (N_3054,N_2428,N_2850);
xnor U3055 (N_3055,N_2415,N_2008);
or U3056 (N_3056,N_2983,N_2916);
nor U3057 (N_3057,N_2032,N_2604);
xor U3058 (N_3058,N_2266,N_2640);
and U3059 (N_3059,N_2743,N_2150);
xnor U3060 (N_3060,N_2348,N_2517);
nor U3061 (N_3061,N_2903,N_2487);
and U3062 (N_3062,N_2727,N_2783);
nor U3063 (N_3063,N_2108,N_2750);
xnor U3064 (N_3064,N_2659,N_2921);
nand U3065 (N_3065,N_2808,N_2300);
xnor U3066 (N_3066,N_2549,N_2219);
xnor U3067 (N_3067,N_2531,N_2013);
nor U3068 (N_3068,N_2435,N_2731);
xor U3069 (N_3069,N_2544,N_2937);
and U3070 (N_3070,N_2124,N_2609);
nand U3071 (N_3071,N_2091,N_2860);
or U3072 (N_3072,N_2296,N_2867);
nor U3073 (N_3073,N_2057,N_2868);
xor U3074 (N_3074,N_2382,N_2802);
and U3075 (N_3075,N_2987,N_2886);
nor U3076 (N_3076,N_2730,N_2591);
nand U3077 (N_3077,N_2607,N_2777);
and U3078 (N_3078,N_2333,N_2995);
nor U3079 (N_3079,N_2644,N_2009);
and U3080 (N_3080,N_2765,N_2977);
xnor U3081 (N_3081,N_2067,N_2776);
nand U3082 (N_3082,N_2143,N_2383);
xnor U3083 (N_3083,N_2047,N_2972);
or U3084 (N_3084,N_2255,N_2632);
and U3085 (N_3085,N_2877,N_2307);
xnor U3086 (N_3086,N_2044,N_2703);
xnor U3087 (N_3087,N_2181,N_2885);
and U3088 (N_3088,N_2469,N_2763);
nor U3089 (N_3089,N_2674,N_2474);
xnor U3090 (N_3090,N_2508,N_2948);
nand U3091 (N_3091,N_2370,N_2608);
xor U3092 (N_3092,N_2542,N_2688);
and U3093 (N_3093,N_2324,N_2414);
nor U3094 (N_3094,N_2624,N_2914);
nand U3095 (N_3095,N_2756,N_2863);
xor U3096 (N_3096,N_2304,N_2368);
or U3097 (N_3097,N_2025,N_2144);
nor U3098 (N_3098,N_2965,N_2200);
nand U3099 (N_3099,N_2174,N_2355);
and U3100 (N_3100,N_2119,N_2521);
xnor U3101 (N_3101,N_2601,N_2179);
nand U3102 (N_3102,N_2720,N_2723);
or U3103 (N_3103,N_2822,N_2949);
xor U3104 (N_3104,N_2071,N_2344);
and U3105 (N_3105,N_2165,N_2760);
xor U3106 (N_3106,N_2906,N_2910);
nor U3107 (N_3107,N_2424,N_2125);
xnor U3108 (N_3108,N_2421,N_2749);
nor U3109 (N_3109,N_2907,N_2001);
xor U3110 (N_3110,N_2484,N_2075);
nand U3111 (N_3111,N_2069,N_2630);
nor U3112 (N_3112,N_2837,N_2928);
and U3113 (N_3113,N_2022,N_2292);
xor U3114 (N_3114,N_2372,N_2898);
and U3115 (N_3115,N_2126,N_2520);
xnor U3116 (N_3116,N_2036,N_2114);
xnor U3117 (N_3117,N_2045,N_2243);
and U3118 (N_3118,N_2671,N_2713);
nor U3119 (N_3119,N_2347,N_2331);
or U3120 (N_3120,N_2667,N_2842);
nor U3121 (N_3121,N_2099,N_2668);
or U3122 (N_3122,N_2230,N_2467);
xnor U3123 (N_3123,N_2175,N_2400);
and U3124 (N_3124,N_2645,N_2177);
nand U3125 (N_3125,N_2375,N_2779);
nor U3126 (N_3126,N_2773,N_2923);
xor U3127 (N_3127,N_2927,N_2187);
and U3128 (N_3128,N_2139,N_2617);
nand U3129 (N_3129,N_2649,N_2831);
nor U3130 (N_3130,N_2839,N_2287);
xor U3131 (N_3131,N_2476,N_2402);
xnor U3132 (N_3132,N_2909,N_2171);
or U3133 (N_3133,N_2354,N_2679);
or U3134 (N_3134,N_2352,N_2312);
and U3135 (N_3135,N_2793,N_2590);
or U3136 (N_3136,N_2892,N_2662);
or U3137 (N_3137,N_2291,N_2890);
nor U3138 (N_3138,N_2103,N_2449);
nor U3139 (N_3139,N_2026,N_2129);
nor U3140 (N_3140,N_2732,N_2345);
xnor U3141 (N_3141,N_2513,N_2172);
and U3142 (N_3142,N_2346,N_2209);
or U3143 (N_3143,N_2681,N_2434);
nor U3144 (N_3144,N_2512,N_2452);
xor U3145 (N_3145,N_2149,N_2932);
nand U3146 (N_3146,N_2335,N_2669);
nand U3147 (N_3147,N_2107,N_2273);
or U3148 (N_3148,N_2495,N_2380);
or U3149 (N_3149,N_2029,N_2130);
nand U3150 (N_3150,N_2507,N_2212);
nand U3151 (N_3151,N_2385,N_2959);
xor U3152 (N_3152,N_2825,N_2473);
nand U3153 (N_3153,N_2829,N_2700);
nor U3154 (N_3154,N_2392,N_2726);
and U3155 (N_3155,N_2852,N_2570);
nor U3156 (N_3156,N_2409,N_2979);
xnor U3157 (N_3157,N_2113,N_2479);
and U3158 (N_3158,N_2018,N_2028);
and U3159 (N_3159,N_2427,N_2794);
xnor U3160 (N_3160,N_2748,N_2185);
xor U3161 (N_3161,N_2166,N_2578);
xor U3162 (N_3162,N_2249,N_2772);
nor U3163 (N_3163,N_2682,N_2718);
or U3164 (N_3164,N_2610,N_2422);
nor U3165 (N_3165,N_2463,N_2694);
xor U3166 (N_3166,N_2642,N_2612);
and U3167 (N_3167,N_2373,N_2514);
nand U3168 (N_3168,N_2444,N_2672);
nand U3169 (N_3169,N_2160,N_2552);
nand U3170 (N_3170,N_2236,N_2391);
nand U3171 (N_3171,N_2786,N_2199);
nor U3172 (N_3172,N_2436,N_2941);
and U3173 (N_3173,N_2695,N_2652);
xnor U3174 (N_3174,N_2832,N_2908);
nor U3175 (N_3175,N_2823,N_2716);
nor U3176 (N_3176,N_2896,N_2288);
and U3177 (N_3177,N_2336,N_2311);
nand U3178 (N_3178,N_2419,N_2122);
xnor U3179 (N_3179,N_2614,N_2167);
xnor U3180 (N_3180,N_2861,N_2192);
xor U3181 (N_3181,N_2675,N_2389);
nand U3182 (N_3182,N_2454,N_2359);
nor U3183 (N_3183,N_2945,N_2360);
nand U3184 (N_3184,N_2579,N_2819);
xnor U3185 (N_3185,N_2820,N_2394);
nor U3186 (N_3186,N_2377,N_2618);
or U3187 (N_3187,N_2568,N_2677);
and U3188 (N_3188,N_2086,N_2220);
or U3189 (N_3189,N_2705,N_2269);
and U3190 (N_3190,N_2942,N_2074);
and U3191 (N_3191,N_2471,N_2097);
nand U3192 (N_3192,N_2622,N_2365);
nand U3193 (N_3193,N_2334,N_2465);
and U3194 (N_3194,N_2319,N_2884);
and U3195 (N_3195,N_2020,N_2462);
nand U3196 (N_3196,N_2806,N_2654);
nor U3197 (N_3197,N_2739,N_2472);
nor U3198 (N_3198,N_2715,N_2733);
xnor U3199 (N_3199,N_2077,N_2338);
and U3200 (N_3200,N_2301,N_2633);
xnor U3201 (N_3201,N_2691,N_2722);
nor U3202 (N_3202,N_2509,N_2260);
xnor U3203 (N_3203,N_2073,N_2762);
nand U3204 (N_3204,N_2186,N_2275);
nand U3205 (N_3205,N_2768,N_2553);
nand U3206 (N_3206,N_2519,N_2423);
nor U3207 (N_3207,N_2342,N_2592);
nor U3208 (N_3208,N_2076,N_2194);
or U3209 (N_3209,N_2790,N_2092);
xnor U3210 (N_3210,N_2801,N_2673);
xnor U3211 (N_3211,N_2361,N_2339);
nand U3212 (N_3212,N_2593,N_2933);
xnor U3213 (N_3213,N_2332,N_2237);
or U3214 (N_3214,N_2441,N_2374);
or U3215 (N_3215,N_2915,N_2504);
nor U3216 (N_3216,N_2676,N_2900);
and U3217 (N_3217,N_2432,N_2974);
xnor U3218 (N_3218,N_2946,N_2537);
nand U3219 (N_3219,N_2178,N_2117);
nand U3220 (N_3220,N_2277,N_2497);
nand U3221 (N_3221,N_2329,N_2431);
nor U3222 (N_3222,N_2105,N_2658);
nand U3223 (N_3223,N_2647,N_2146);
nand U3224 (N_3224,N_2796,N_2056);
and U3225 (N_3225,N_2587,N_2872);
xor U3226 (N_3226,N_2048,N_2271);
nor U3227 (N_3227,N_2784,N_2501);
or U3228 (N_3228,N_2874,N_2309);
and U3229 (N_3229,N_2145,N_2851);
xnor U3230 (N_3230,N_2093,N_2881);
xnor U3231 (N_3231,N_2247,N_2065);
xnor U3232 (N_3232,N_2498,N_2957);
xor U3233 (N_3233,N_2745,N_2252);
xor U3234 (N_3234,N_2325,N_2651);
or U3235 (N_3235,N_2262,N_2935);
or U3236 (N_3236,N_2795,N_2986);
and U3237 (N_3237,N_2378,N_2060);
or U3238 (N_3238,N_2381,N_2278);
nor U3239 (N_3239,N_2303,N_2284);
nor U3240 (N_3240,N_2975,N_2480);
nand U3241 (N_3241,N_2201,N_2259);
nand U3242 (N_3242,N_2543,N_2466);
or U3243 (N_3243,N_2196,N_2862);
xnor U3244 (N_3244,N_2746,N_2407);
xnor U3245 (N_3245,N_2859,N_2821);
nand U3246 (N_3246,N_2984,N_2152);
nor U3247 (N_3247,N_2664,N_2556);
and U3248 (N_3248,N_2738,N_2523);
nand U3249 (N_3249,N_2613,N_2217);
xnor U3250 (N_3250,N_2947,N_2148);
xnor U3251 (N_3251,N_2737,N_2775);
or U3252 (N_3252,N_2663,N_2666);
nor U3253 (N_3253,N_2379,N_2460);
nor U3254 (N_3254,N_2351,N_2708);
and U3255 (N_3255,N_2978,N_2701);
xnor U3256 (N_3256,N_2897,N_2021);
and U3257 (N_3257,N_2222,N_2606);
nor U3258 (N_3258,N_2510,N_2468);
and U3259 (N_3259,N_2364,N_2982);
nand U3260 (N_3260,N_2182,N_2969);
xor U3261 (N_3261,N_2328,N_2035);
nor U3262 (N_3262,N_2318,N_2558);
or U3263 (N_3263,N_2596,N_2871);
nor U3264 (N_3264,N_2369,N_2376);
xor U3265 (N_3265,N_2619,N_2482);
nand U3266 (N_3266,N_2005,N_2611);
and U3267 (N_3267,N_2461,N_2582);
and U3268 (N_3268,N_2555,N_2807);
and U3269 (N_3269,N_2653,N_2758);
xnor U3270 (N_3270,N_2398,N_2561);
xnor U3271 (N_3271,N_2063,N_2006);
nand U3272 (N_3272,N_2087,N_2450);
nand U3273 (N_3273,N_2173,N_2757);
and U3274 (N_3274,N_2214,N_2778);
nor U3275 (N_3275,N_2202,N_2964);
and U3276 (N_3276,N_2153,N_2159);
or U3277 (N_3277,N_2934,N_2017);
nand U3278 (N_3278,N_2440,N_2416);
and U3279 (N_3279,N_2953,N_2062);
nor U3280 (N_3280,N_2034,N_2492);
nand U3281 (N_3281,N_2629,N_2003);
nand U3282 (N_3282,N_2310,N_2014);
or U3283 (N_3283,N_2051,N_2283);
or U3284 (N_3284,N_2496,N_2157);
and U3285 (N_3285,N_2628,N_2854);
nor U3286 (N_3286,N_2585,N_2425);
xor U3287 (N_3287,N_2388,N_2976);
nand U3288 (N_3288,N_2207,N_2936);
nor U3289 (N_3289,N_2635,N_2846);
xnor U3290 (N_3290,N_2102,N_2226);
xor U3291 (N_3291,N_2721,N_2992);
nand U3292 (N_3292,N_2314,N_2689);
or U3293 (N_3293,N_2855,N_2563);
xor U3294 (N_3294,N_2805,N_2594);
nor U3295 (N_3295,N_2637,N_2420);
xnor U3296 (N_3296,N_2448,N_2597);
or U3297 (N_3297,N_2258,N_2503);
and U3298 (N_3298,N_2362,N_2742);
and U3299 (N_3299,N_2529,N_2767);
nor U3300 (N_3300,N_2228,N_2843);
and U3301 (N_3301,N_2483,N_2250);
xor U3302 (N_3302,N_2971,N_2188);
or U3303 (N_3303,N_2660,N_2401);
nand U3304 (N_3304,N_2015,N_2299);
and U3305 (N_3305,N_2943,N_2952);
xnor U3306 (N_3306,N_2180,N_2322);
nand U3307 (N_3307,N_2010,N_2525);
nor U3308 (N_3308,N_2151,N_2963);
nand U3309 (N_3309,N_2566,N_2834);
or U3310 (N_3310,N_2110,N_2827);
and U3311 (N_3311,N_2567,N_2811);
and U3312 (N_3312,N_2725,N_2858);
nand U3313 (N_3313,N_2205,N_2245);
xnor U3314 (N_3314,N_2626,N_2791);
or U3315 (N_3315,N_2882,N_2598);
nand U3316 (N_3316,N_2627,N_2193);
or U3317 (N_3317,N_2803,N_2841);
xor U3318 (N_3318,N_2290,N_2412);
and U3319 (N_3319,N_2889,N_2393);
nor U3320 (N_3320,N_2279,N_2078);
nand U3321 (N_3321,N_2043,N_2261);
or U3322 (N_3322,N_2458,N_2623);
and U3323 (N_3323,N_2251,N_2583);
or U3324 (N_3324,N_2443,N_2341);
and U3325 (N_3325,N_2459,N_2902);
xor U3326 (N_3326,N_2233,N_2101);
xnor U3327 (N_3327,N_2294,N_2845);
nor U3328 (N_3328,N_2115,N_2536);
xor U3329 (N_3329,N_2696,N_2924);
nor U3330 (N_3330,N_2049,N_2996);
and U3331 (N_3331,N_2699,N_2183);
nand U3332 (N_3332,N_2836,N_2070);
and U3333 (N_3333,N_2925,N_2163);
or U3334 (N_3334,N_2493,N_2390);
xnor U3335 (N_3335,N_2655,N_2865);
xnor U3336 (N_3336,N_2580,N_2240);
and U3337 (N_3337,N_2176,N_2136);
xor U3338 (N_3338,N_2511,N_2257);
and U3339 (N_3339,N_2413,N_2343);
and U3340 (N_3340,N_2327,N_2216);
or U3341 (N_3341,N_2161,N_2798);
nor U3342 (N_3342,N_2875,N_2697);
nand U3343 (N_3343,N_2888,N_2191);
nor U3344 (N_3344,N_2430,N_2132);
xnor U3345 (N_3345,N_2960,N_2438);
or U3346 (N_3346,N_2643,N_2985);
nand U3347 (N_3347,N_2638,N_2464);
nand U3348 (N_3348,N_2572,N_2395);
and U3349 (N_3349,N_2589,N_2268);
or U3350 (N_3350,N_2270,N_2326);
nand U3351 (N_3351,N_2477,N_2481);
or U3352 (N_3352,N_2349,N_2457);
xor U3353 (N_3353,N_2989,N_2363);
nor U3354 (N_3354,N_2138,N_2535);
nor U3355 (N_3355,N_2281,N_2588);
or U3356 (N_3356,N_2866,N_2447);
xor U3357 (N_3357,N_2242,N_2050);
or U3358 (N_3358,N_2147,N_2891);
nor U3359 (N_3359,N_2221,N_2797);
and U3360 (N_3360,N_2804,N_2096);
or U3361 (N_3361,N_2429,N_2616);
nand U3362 (N_3362,N_2238,N_2340);
nor U3363 (N_3363,N_2912,N_2661);
nor U3364 (N_3364,N_2156,N_2787);
and U3365 (N_3365,N_2231,N_2698);
or U3366 (N_3366,N_2766,N_2789);
nand U3367 (N_3367,N_2848,N_2111);
nand U3368 (N_3368,N_2870,N_2711);
xnor U3369 (N_3369,N_2140,N_2499);
nor U3370 (N_3370,N_2031,N_2002);
nor U3371 (N_3371,N_2781,N_2988);
or U3372 (N_3372,N_2569,N_2939);
or U3373 (N_3373,N_2665,N_2042);
and U3374 (N_3374,N_2605,N_2120);
and U3375 (N_3375,N_2500,N_2755);
xnor U3376 (N_3376,N_2337,N_2690);
nor U3377 (N_3377,N_2104,N_2554);
and U3378 (N_3378,N_2004,N_2007);
nand U3379 (N_3379,N_2272,N_2072);
nor U3380 (N_3380,N_2625,N_2704);
xor U3381 (N_3381,N_2204,N_2810);
xnor U3382 (N_3382,N_2956,N_2455);
nand U3383 (N_3383,N_2053,N_2901);
nor U3384 (N_3384,N_2197,N_2293);
and U3385 (N_3385,N_2532,N_2584);
and U3386 (N_3386,N_2158,N_2248);
and U3387 (N_3387,N_2317,N_2106);
nor U3388 (N_3388,N_2518,N_2019);
or U3389 (N_3389,N_2442,N_2528);
nor U3390 (N_3390,N_2734,N_2162);
nand U3391 (N_3391,N_2263,N_2276);
and U3392 (N_3392,N_2169,N_2724);
and U3393 (N_3393,N_2849,N_2573);
nand U3394 (N_3394,N_2405,N_2470);
nor U3395 (N_3395,N_2195,N_2780);
xor U3396 (N_3396,N_2747,N_2702);
and U3397 (N_3397,N_2505,N_2930);
nand U3398 (N_3398,N_2297,N_2575);
or U3399 (N_3399,N_2189,N_2857);
nor U3400 (N_3400,N_2406,N_2456);
nand U3401 (N_3401,N_2687,N_2264);
nor U3402 (N_3402,N_2550,N_2729);
or U3403 (N_3403,N_2350,N_2289);
or U3404 (N_3404,N_2564,N_2137);
xor U3405 (N_3405,N_2782,N_2085);
or U3406 (N_3406,N_2225,N_2894);
or U3407 (N_3407,N_2280,N_2386);
nor U3408 (N_3408,N_2411,N_2869);
or U3409 (N_3409,N_2599,N_2203);
nor U3410 (N_3410,N_2887,N_2530);
xor U3411 (N_3411,N_2082,N_2058);
nand U3412 (N_3412,N_2155,N_2522);
xor U3413 (N_3413,N_2223,N_2128);
nor U3414 (N_3414,N_2064,N_2899);
or U3415 (N_3415,N_2710,N_2524);
xor U3416 (N_3416,N_2302,N_2315);
or U3417 (N_3417,N_2215,N_2208);
nor U3418 (N_3418,N_2308,N_2538);
xor U3419 (N_3419,N_2595,N_2088);
and U3420 (N_3420,N_2486,N_2118);
and U3421 (N_3421,N_2000,N_2560);
nor U3422 (N_3422,N_2211,N_2824);
nand U3423 (N_3423,N_2094,N_2285);
nand U3424 (N_3424,N_2685,N_2833);
nor U3425 (N_3425,N_2838,N_2184);
or U3426 (N_3426,N_2358,N_2135);
and U3427 (N_3427,N_2305,N_2298);
and U3428 (N_3428,N_2955,N_2433);
nand U3429 (N_3429,N_2418,N_2066);
or U3430 (N_3430,N_2761,N_2210);
and U3431 (N_3431,N_2559,N_2353);
nand U3432 (N_3432,N_2577,N_2586);
or U3433 (N_3433,N_2650,N_2800);
nand U3434 (N_3434,N_2408,N_2054);
nand U3435 (N_3435,N_2046,N_2384);
nand U3436 (N_3436,N_2639,N_2826);
nand U3437 (N_3437,N_2274,N_2876);
xnor U3438 (N_3438,N_2950,N_2371);
or U3439 (N_3439,N_2265,N_2997);
and U3440 (N_3440,N_2670,N_2853);
xor U3441 (N_3441,N_2736,N_2815);
or U3442 (N_3442,N_2873,N_2488);
or U3443 (N_3443,N_2545,N_2788);
or U3444 (N_3444,N_2323,N_2387);
xor U3445 (N_3445,N_2878,N_2813);
nand U3446 (N_3446,N_2993,N_2254);
and U3447 (N_3447,N_2814,N_2631);
and U3448 (N_3448,N_2751,N_2453);
and U3449 (N_3449,N_2744,N_2244);
nor U3450 (N_3450,N_2109,N_2565);
xor U3451 (N_3451,N_2234,N_2684);
nor U3452 (N_3452,N_2011,N_2621);
nand U3453 (N_3453,N_2883,N_2502);
xor U3454 (N_3454,N_2396,N_2574);
xnor U3455 (N_3455,N_2712,N_2966);
or U3456 (N_3456,N_2692,N_2576);
nor U3457 (N_3457,N_2539,N_2581);
and U3458 (N_3458,N_2557,N_2083);
nand U3459 (N_3459,N_2170,N_2027);
nor U3460 (N_3460,N_2224,N_2938);
nand U3461 (N_3461,N_2227,N_2818);
or U3462 (N_3462,N_2142,N_2321);
and U3463 (N_3463,N_2571,N_2239);
nor U3464 (N_3464,N_2417,N_2546);
nand U3465 (N_3465,N_2735,N_2991);
or U3466 (N_3466,N_2451,N_2840);
or U3467 (N_3467,N_2253,N_2719);
or U3468 (N_3468,N_2562,N_2981);
and U3469 (N_3469,N_2190,N_2491);
xnor U3470 (N_3470,N_2198,N_2489);
or U3471 (N_3471,N_2154,N_2016);
nor U3472 (N_3472,N_2080,N_2024);
or U3473 (N_3473,N_2920,N_2830);
nand U3474 (N_3474,N_2320,N_2759);
xor U3475 (N_3475,N_2306,N_2012);
nor U3476 (N_3476,N_2439,N_2127);
nand U3477 (N_3477,N_2506,N_2753);
or U3478 (N_3478,N_2055,N_2799);
and U3479 (N_3479,N_2990,N_2847);
or U3480 (N_3480,N_2693,N_2602);
xnor U3481 (N_3481,N_2880,N_2485);
and U3482 (N_3482,N_2366,N_2098);
nand U3483 (N_3483,N_2316,N_2944);
and U3484 (N_3484,N_2313,N_2769);
nor U3485 (N_3485,N_2356,N_2917);
nand U3486 (N_3486,N_2600,N_2774);
xnor U3487 (N_3487,N_2905,N_2958);
nor U3488 (N_3488,N_2286,N_2475);
or U3489 (N_3489,N_2023,N_2399);
or U3490 (N_3490,N_2770,N_2041);
xor U3491 (N_3491,N_2533,N_2879);
and U3492 (N_3492,N_2404,N_2516);
or U3493 (N_3493,N_2728,N_2929);
or U3494 (N_3494,N_2615,N_2490);
xor U3495 (N_3495,N_2241,N_2235);
or U3496 (N_3496,N_2962,N_2134);
nand U3497 (N_3497,N_2835,N_2040);
xor U3498 (N_3498,N_2295,N_2357);
or U3499 (N_3499,N_2037,N_2551);
xor U3500 (N_3500,N_2889,N_2370);
and U3501 (N_3501,N_2755,N_2463);
xnor U3502 (N_3502,N_2099,N_2896);
nor U3503 (N_3503,N_2887,N_2536);
nor U3504 (N_3504,N_2927,N_2871);
nor U3505 (N_3505,N_2958,N_2770);
nand U3506 (N_3506,N_2534,N_2102);
and U3507 (N_3507,N_2549,N_2143);
and U3508 (N_3508,N_2214,N_2011);
xnor U3509 (N_3509,N_2641,N_2578);
or U3510 (N_3510,N_2863,N_2541);
xor U3511 (N_3511,N_2654,N_2439);
xnor U3512 (N_3512,N_2339,N_2784);
or U3513 (N_3513,N_2029,N_2444);
xnor U3514 (N_3514,N_2656,N_2583);
nand U3515 (N_3515,N_2021,N_2158);
nand U3516 (N_3516,N_2702,N_2749);
nor U3517 (N_3517,N_2635,N_2068);
xor U3518 (N_3518,N_2927,N_2001);
nor U3519 (N_3519,N_2068,N_2608);
or U3520 (N_3520,N_2137,N_2289);
and U3521 (N_3521,N_2346,N_2409);
nand U3522 (N_3522,N_2706,N_2999);
xnor U3523 (N_3523,N_2698,N_2607);
nor U3524 (N_3524,N_2675,N_2139);
nor U3525 (N_3525,N_2297,N_2161);
or U3526 (N_3526,N_2097,N_2532);
and U3527 (N_3527,N_2688,N_2547);
xnor U3528 (N_3528,N_2371,N_2711);
or U3529 (N_3529,N_2535,N_2310);
nand U3530 (N_3530,N_2136,N_2438);
or U3531 (N_3531,N_2270,N_2569);
nor U3532 (N_3532,N_2108,N_2870);
nand U3533 (N_3533,N_2173,N_2065);
nand U3534 (N_3534,N_2412,N_2534);
nor U3535 (N_3535,N_2865,N_2396);
nand U3536 (N_3536,N_2509,N_2198);
nor U3537 (N_3537,N_2082,N_2950);
nand U3538 (N_3538,N_2089,N_2559);
nand U3539 (N_3539,N_2556,N_2991);
nand U3540 (N_3540,N_2408,N_2474);
or U3541 (N_3541,N_2517,N_2539);
nand U3542 (N_3542,N_2471,N_2897);
nor U3543 (N_3543,N_2386,N_2863);
or U3544 (N_3544,N_2069,N_2617);
and U3545 (N_3545,N_2990,N_2204);
xnor U3546 (N_3546,N_2911,N_2112);
nand U3547 (N_3547,N_2500,N_2705);
xnor U3548 (N_3548,N_2070,N_2703);
or U3549 (N_3549,N_2346,N_2321);
nor U3550 (N_3550,N_2706,N_2455);
nand U3551 (N_3551,N_2301,N_2814);
nand U3552 (N_3552,N_2761,N_2156);
and U3553 (N_3553,N_2527,N_2064);
xor U3554 (N_3554,N_2568,N_2579);
and U3555 (N_3555,N_2369,N_2031);
or U3556 (N_3556,N_2508,N_2572);
nand U3557 (N_3557,N_2929,N_2763);
nand U3558 (N_3558,N_2712,N_2137);
xnor U3559 (N_3559,N_2507,N_2820);
nor U3560 (N_3560,N_2124,N_2920);
or U3561 (N_3561,N_2270,N_2970);
nor U3562 (N_3562,N_2476,N_2338);
and U3563 (N_3563,N_2245,N_2582);
nor U3564 (N_3564,N_2119,N_2594);
and U3565 (N_3565,N_2693,N_2361);
or U3566 (N_3566,N_2564,N_2959);
or U3567 (N_3567,N_2212,N_2699);
and U3568 (N_3568,N_2920,N_2136);
nand U3569 (N_3569,N_2643,N_2105);
nand U3570 (N_3570,N_2867,N_2859);
nand U3571 (N_3571,N_2451,N_2331);
nor U3572 (N_3572,N_2506,N_2517);
xor U3573 (N_3573,N_2030,N_2643);
or U3574 (N_3574,N_2947,N_2447);
nor U3575 (N_3575,N_2589,N_2032);
nand U3576 (N_3576,N_2816,N_2724);
nor U3577 (N_3577,N_2887,N_2549);
xor U3578 (N_3578,N_2054,N_2230);
nor U3579 (N_3579,N_2178,N_2514);
nand U3580 (N_3580,N_2087,N_2773);
and U3581 (N_3581,N_2361,N_2861);
and U3582 (N_3582,N_2144,N_2115);
xor U3583 (N_3583,N_2901,N_2526);
xnor U3584 (N_3584,N_2185,N_2174);
nor U3585 (N_3585,N_2873,N_2791);
and U3586 (N_3586,N_2576,N_2187);
xor U3587 (N_3587,N_2199,N_2613);
xnor U3588 (N_3588,N_2846,N_2381);
nor U3589 (N_3589,N_2287,N_2667);
nor U3590 (N_3590,N_2444,N_2809);
nand U3591 (N_3591,N_2300,N_2183);
nand U3592 (N_3592,N_2999,N_2435);
or U3593 (N_3593,N_2816,N_2294);
xor U3594 (N_3594,N_2960,N_2871);
and U3595 (N_3595,N_2021,N_2593);
xnor U3596 (N_3596,N_2072,N_2250);
xnor U3597 (N_3597,N_2830,N_2963);
nand U3598 (N_3598,N_2741,N_2442);
nand U3599 (N_3599,N_2113,N_2235);
nand U3600 (N_3600,N_2483,N_2672);
xor U3601 (N_3601,N_2956,N_2006);
nor U3602 (N_3602,N_2958,N_2467);
nand U3603 (N_3603,N_2608,N_2846);
or U3604 (N_3604,N_2756,N_2263);
nor U3605 (N_3605,N_2111,N_2192);
nand U3606 (N_3606,N_2829,N_2005);
nand U3607 (N_3607,N_2886,N_2423);
xor U3608 (N_3608,N_2648,N_2582);
nand U3609 (N_3609,N_2345,N_2288);
and U3610 (N_3610,N_2937,N_2821);
nor U3611 (N_3611,N_2580,N_2409);
or U3612 (N_3612,N_2352,N_2303);
xnor U3613 (N_3613,N_2772,N_2198);
nand U3614 (N_3614,N_2500,N_2771);
and U3615 (N_3615,N_2204,N_2402);
and U3616 (N_3616,N_2846,N_2856);
or U3617 (N_3617,N_2964,N_2487);
nand U3618 (N_3618,N_2838,N_2001);
or U3619 (N_3619,N_2847,N_2367);
or U3620 (N_3620,N_2873,N_2304);
xor U3621 (N_3621,N_2384,N_2441);
xor U3622 (N_3622,N_2892,N_2293);
xnor U3623 (N_3623,N_2436,N_2981);
nor U3624 (N_3624,N_2041,N_2502);
or U3625 (N_3625,N_2584,N_2835);
nand U3626 (N_3626,N_2365,N_2010);
and U3627 (N_3627,N_2123,N_2886);
nand U3628 (N_3628,N_2587,N_2629);
and U3629 (N_3629,N_2051,N_2344);
and U3630 (N_3630,N_2826,N_2489);
or U3631 (N_3631,N_2392,N_2657);
and U3632 (N_3632,N_2452,N_2177);
xor U3633 (N_3633,N_2128,N_2751);
xor U3634 (N_3634,N_2620,N_2661);
or U3635 (N_3635,N_2648,N_2580);
nor U3636 (N_3636,N_2444,N_2466);
xor U3637 (N_3637,N_2904,N_2402);
nor U3638 (N_3638,N_2200,N_2524);
xnor U3639 (N_3639,N_2648,N_2507);
and U3640 (N_3640,N_2627,N_2401);
or U3641 (N_3641,N_2654,N_2700);
xor U3642 (N_3642,N_2292,N_2369);
or U3643 (N_3643,N_2172,N_2817);
nor U3644 (N_3644,N_2422,N_2441);
nand U3645 (N_3645,N_2349,N_2160);
xor U3646 (N_3646,N_2014,N_2965);
or U3647 (N_3647,N_2144,N_2038);
and U3648 (N_3648,N_2946,N_2931);
nor U3649 (N_3649,N_2865,N_2482);
xor U3650 (N_3650,N_2683,N_2998);
or U3651 (N_3651,N_2806,N_2705);
and U3652 (N_3652,N_2773,N_2647);
nor U3653 (N_3653,N_2625,N_2810);
or U3654 (N_3654,N_2415,N_2588);
and U3655 (N_3655,N_2237,N_2715);
and U3656 (N_3656,N_2652,N_2917);
and U3657 (N_3657,N_2413,N_2651);
nand U3658 (N_3658,N_2943,N_2160);
xnor U3659 (N_3659,N_2799,N_2167);
or U3660 (N_3660,N_2235,N_2957);
nor U3661 (N_3661,N_2106,N_2116);
nand U3662 (N_3662,N_2220,N_2715);
nor U3663 (N_3663,N_2847,N_2956);
and U3664 (N_3664,N_2722,N_2195);
xnor U3665 (N_3665,N_2744,N_2764);
and U3666 (N_3666,N_2168,N_2453);
nand U3667 (N_3667,N_2767,N_2073);
nand U3668 (N_3668,N_2027,N_2298);
nor U3669 (N_3669,N_2730,N_2677);
xnor U3670 (N_3670,N_2913,N_2047);
and U3671 (N_3671,N_2533,N_2357);
xnor U3672 (N_3672,N_2952,N_2193);
or U3673 (N_3673,N_2724,N_2271);
and U3674 (N_3674,N_2793,N_2568);
or U3675 (N_3675,N_2799,N_2878);
and U3676 (N_3676,N_2280,N_2172);
nand U3677 (N_3677,N_2936,N_2082);
nor U3678 (N_3678,N_2009,N_2924);
nand U3679 (N_3679,N_2476,N_2015);
nand U3680 (N_3680,N_2054,N_2578);
xor U3681 (N_3681,N_2813,N_2178);
nand U3682 (N_3682,N_2124,N_2306);
xor U3683 (N_3683,N_2086,N_2548);
and U3684 (N_3684,N_2407,N_2890);
and U3685 (N_3685,N_2665,N_2812);
nor U3686 (N_3686,N_2753,N_2670);
and U3687 (N_3687,N_2374,N_2688);
and U3688 (N_3688,N_2705,N_2171);
nor U3689 (N_3689,N_2738,N_2411);
nor U3690 (N_3690,N_2651,N_2767);
and U3691 (N_3691,N_2243,N_2955);
xnor U3692 (N_3692,N_2682,N_2650);
nor U3693 (N_3693,N_2597,N_2008);
nand U3694 (N_3694,N_2816,N_2685);
or U3695 (N_3695,N_2792,N_2225);
and U3696 (N_3696,N_2504,N_2396);
xor U3697 (N_3697,N_2614,N_2558);
nand U3698 (N_3698,N_2712,N_2883);
xnor U3699 (N_3699,N_2620,N_2845);
xor U3700 (N_3700,N_2731,N_2003);
or U3701 (N_3701,N_2847,N_2290);
xor U3702 (N_3702,N_2452,N_2673);
and U3703 (N_3703,N_2767,N_2734);
or U3704 (N_3704,N_2549,N_2517);
nor U3705 (N_3705,N_2195,N_2294);
and U3706 (N_3706,N_2345,N_2439);
xor U3707 (N_3707,N_2531,N_2233);
or U3708 (N_3708,N_2086,N_2819);
and U3709 (N_3709,N_2229,N_2435);
nand U3710 (N_3710,N_2835,N_2819);
nand U3711 (N_3711,N_2394,N_2454);
xnor U3712 (N_3712,N_2143,N_2932);
or U3713 (N_3713,N_2670,N_2424);
xnor U3714 (N_3714,N_2905,N_2806);
and U3715 (N_3715,N_2588,N_2156);
xnor U3716 (N_3716,N_2056,N_2011);
or U3717 (N_3717,N_2870,N_2890);
nor U3718 (N_3718,N_2957,N_2744);
nor U3719 (N_3719,N_2971,N_2522);
and U3720 (N_3720,N_2541,N_2179);
or U3721 (N_3721,N_2452,N_2317);
nor U3722 (N_3722,N_2291,N_2415);
nor U3723 (N_3723,N_2335,N_2548);
nor U3724 (N_3724,N_2694,N_2906);
nand U3725 (N_3725,N_2170,N_2775);
or U3726 (N_3726,N_2664,N_2200);
xor U3727 (N_3727,N_2929,N_2241);
or U3728 (N_3728,N_2973,N_2523);
xor U3729 (N_3729,N_2643,N_2824);
nand U3730 (N_3730,N_2239,N_2547);
xnor U3731 (N_3731,N_2533,N_2826);
nand U3732 (N_3732,N_2369,N_2247);
xnor U3733 (N_3733,N_2236,N_2093);
xor U3734 (N_3734,N_2799,N_2575);
nor U3735 (N_3735,N_2917,N_2408);
xnor U3736 (N_3736,N_2547,N_2884);
xnor U3737 (N_3737,N_2121,N_2471);
xor U3738 (N_3738,N_2930,N_2520);
or U3739 (N_3739,N_2210,N_2419);
nor U3740 (N_3740,N_2331,N_2870);
xor U3741 (N_3741,N_2174,N_2585);
or U3742 (N_3742,N_2364,N_2946);
and U3743 (N_3743,N_2227,N_2789);
or U3744 (N_3744,N_2674,N_2386);
nand U3745 (N_3745,N_2460,N_2205);
or U3746 (N_3746,N_2491,N_2221);
nor U3747 (N_3747,N_2639,N_2222);
nand U3748 (N_3748,N_2115,N_2292);
xnor U3749 (N_3749,N_2361,N_2100);
and U3750 (N_3750,N_2780,N_2388);
nand U3751 (N_3751,N_2836,N_2723);
xor U3752 (N_3752,N_2225,N_2952);
or U3753 (N_3753,N_2742,N_2293);
nand U3754 (N_3754,N_2133,N_2341);
and U3755 (N_3755,N_2623,N_2498);
or U3756 (N_3756,N_2016,N_2322);
or U3757 (N_3757,N_2298,N_2223);
or U3758 (N_3758,N_2185,N_2639);
nand U3759 (N_3759,N_2723,N_2334);
nand U3760 (N_3760,N_2770,N_2181);
nand U3761 (N_3761,N_2632,N_2746);
xor U3762 (N_3762,N_2514,N_2220);
or U3763 (N_3763,N_2190,N_2950);
nor U3764 (N_3764,N_2438,N_2016);
xor U3765 (N_3765,N_2388,N_2298);
or U3766 (N_3766,N_2486,N_2156);
nand U3767 (N_3767,N_2707,N_2097);
nand U3768 (N_3768,N_2754,N_2234);
nor U3769 (N_3769,N_2991,N_2929);
or U3770 (N_3770,N_2780,N_2149);
nand U3771 (N_3771,N_2944,N_2349);
and U3772 (N_3772,N_2696,N_2166);
nor U3773 (N_3773,N_2677,N_2067);
and U3774 (N_3774,N_2398,N_2173);
nor U3775 (N_3775,N_2165,N_2828);
xor U3776 (N_3776,N_2887,N_2240);
nand U3777 (N_3777,N_2726,N_2277);
nor U3778 (N_3778,N_2986,N_2127);
and U3779 (N_3779,N_2276,N_2237);
and U3780 (N_3780,N_2742,N_2788);
nor U3781 (N_3781,N_2918,N_2623);
nor U3782 (N_3782,N_2608,N_2862);
and U3783 (N_3783,N_2699,N_2227);
nor U3784 (N_3784,N_2586,N_2463);
or U3785 (N_3785,N_2740,N_2163);
and U3786 (N_3786,N_2618,N_2645);
and U3787 (N_3787,N_2974,N_2763);
nor U3788 (N_3788,N_2265,N_2168);
or U3789 (N_3789,N_2828,N_2761);
xor U3790 (N_3790,N_2939,N_2541);
or U3791 (N_3791,N_2133,N_2960);
and U3792 (N_3792,N_2125,N_2150);
xor U3793 (N_3793,N_2522,N_2387);
or U3794 (N_3794,N_2115,N_2954);
xor U3795 (N_3795,N_2651,N_2454);
xnor U3796 (N_3796,N_2674,N_2533);
and U3797 (N_3797,N_2785,N_2438);
nand U3798 (N_3798,N_2339,N_2154);
nand U3799 (N_3799,N_2602,N_2932);
nor U3800 (N_3800,N_2153,N_2784);
and U3801 (N_3801,N_2068,N_2924);
nor U3802 (N_3802,N_2989,N_2663);
nor U3803 (N_3803,N_2519,N_2695);
nor U3804 (N_3804,N_2162,N_2772);
xnor U3805 (N_3805,N_2430,N_2804);
or U3806 (N_3806,N_2085,N_2603);
xnor U3807 (N_3807,N_2680,N_2900);
or U3808 (N_3808,N_2423,N_2600);
nand U3809 (N_3809,N_2205,N_2610);
nand U3810 (N_3810,N_2840,N_2523);
and U3811 (N_3811,N_2969,N_2716);
nor U3812 (N_3812,N_2446,N_2378);
nor U3813 (N_3813,N_2398,N_2238);
nor U3814 (N_3814,N_2938,N_2969);
and U3815 (N_3815,N_2780,N_2686);
and U3816 (N_3816,N_2833,N_2651);
xor U3817 (N_3817,N_2852,N_2562);
and U3818 (N_3818,N_2942,N_2724);
or U3819 (N_3819,N_2707,N_2624);
nand U3820 (N_3820,N_2134,N_2089);
or U3821 (N_3821,N_2024,N_2210);
and U3822 (N_3822,N_2141,N_2393);
xnor U3823 (N_3823,N_2735,N_2579);
xor U3824 (N_3824,N_2802,N_2402);
and U3825 (N_3825,N_2323,N_2242);
xnor U3826 (N_3826,N_2230,N_2936);
nor U3827 (N_3827,N_2064,N_2681);
nor U3828 (N_3828,N_2152,N_2405);
or U3829 (N_3829,N_2791,N_2526);
and U3830 (N_3830,N_2482,N_2053);
or U3831 (N_3831,N_2040,N_2968);
xnor U3832 (N_3832,N_2996,N_2233);
xor U3833 (N_3833,N_2303,N_2312);
nor U3834 (N_3834,N_2629,N_2763);
nor U3835 (N_3835,N_2511,N_2950);
xnor U3836 (N_3836,N_2216,N_2474);
or U3837 (N_3837,N_2084,N_2449);
and U3838 (N_3838,N_2890,N_2159);
nor U3839 (N_3839,N_2344,N_2563);
nand U3840 (N_3840,N_2559,N_2837);
xnor U3841 (N_3841,N_2821,N_2510);
nand U3842 (N_3842,N_2945,N_2737);
or U3843 (N_3843,N_2729,N_2024);
or U3844 (N_3844,N_2644,N_2490);
and U3845 (N_3845,N_2289,N_2872);
nor U3846 (N_3846,N_2196,N_2090);
nor U3847 (N_3847,N_2262,N_2353);
nor U3848 (N_3848,N_2227,N_2243);
nor U3849 (N_3849,N_2044,N_2099);
or U3850 (N_3850,N_2735,N_2355);
or U3851 (N_3851,N_2352,N_2449);
nand U3852 (N_3852,N_2902,N_2567);
nor U3853 (N_3853,N_2509,N_2086);
nor U3854 (N_3854,N_2366,N_2388);
nand U3855 (N_3855,N_2317,N_2104);
nand U3856 (N_3856,N_2810,N_2994);
or U3857 (N_3857,N_2832,N_2650);
nand U3858 (N_3858,N_2260,N_2553);
and U3859 (N_3859,N_2308,N_2821);
xnor U3860 (N_3860,N_2448,N_2985);
nand U3861 (N_3861,N_2758,N_2853);
nand U3862 (N_3862,N_2167,N_2020);
nor U3863 (N_3863,N_2987,N_2916);
nor U3864 (N_3864,N_2004,N_2294);
xnor U3865 (N_3865,N_2604,N_2752);
and U3866 (N_3866,N_2208,N_2118);
and U3867 (N_3867,N_2075,N_2126);
nand U3868 (N_3868,N_2268,N_2413);
xor U3869 (N_3869,N_2500,N_2894);
nand U3870 (N_3870,N_2188,N_2266);
and U3871 (N_3871,N_2423,N_2819);
and U3872 (N_3872,N_2670,N_2384);
nand U3873 (N_3873,N_2496,N_2287);
nand U3874 (N_3874,N_2167,N_2545);
nor U3875 (N_3875,N_2673,N_2146);
xor U3876 (N_3876,N_2660,N_2760);
nand U3877 (N_3877,N_2090,N_2957);
nand U3878 (N_3878,N_2157,N_2796);
nor U3879 (N_3879,N_2192,N_2899);
nand U3880 (N_3880,N_2410,N_2497);
nor U3881 (N_3881,N_2276,N_2682);
nor U3882 (N_3882,N_2871,N_2621);
or U3883 (N_3883,N_2619,N_2412);
and U3884 (N_3884,N_2605,N_2750);
or U3885 (N_3885,N_2094,N_2978);
or U3886 (N_3886,N_2719,N_2860);
and U3887 (N_3887,N_2418,N_2593);
or U3888 (N_3888,N_2213,N_2435);
xnor U3889 (N_3889,N_2889,N_2734);
and U3890 (N_3890,N_2560,N_2584);
nand U3891 (N_3891,N_2954,N_2444);
nand U3892 (N_3892,N_2021,N_2613);
or U3893 (N_3893,N_2034,N_2061);
xor U3894 (N_3894,N_2640,N_2295);
and U3895 (N_3895,N_2725,N_2624);
and U3896 (N_3896,N_2611,N_2878);
or U3897 (N_3897,N_2745,N_2411);
or U3898 (N_3898,N_2492,N_2389);
nand U3899 (N_3899,N_2121,N_2886);
nand U3900 (N_3900,N_2955,N_2847);
nor U3901 (N_3901,N_2549,N_2024);
and U3902 (N_3902,N_2372,N_2996);
or U3903 (N_3903,N_2046,N_2844);
xor U3904 (N_3904,N_2860,N_2806);
or U3905 (N_3905,N_2771,N_2689);
xor U3906 (N_3906,N_2840,N_2333);
xor U3907 (N_3907,N_2558,N_2019);
xor U3908 (N_3908,N_2894,N_2022);
nand U3909 (N_3909,N_2560,N_2708);
xor U3910 (N_3910,N_2149,N_2179);
nand U3911 (N_3911,N_2723,N_2171);
and U3912 (N_3912,N_2061,N_2995);
or U3913 (N_3913,N_2233,N_2869);
and U3914 (N_3914,N_2442,N_2300);
or U3915 (N_3915,N_2059,N_2972);
and U3916 (N_3916,N_2256,N_2519);
and U3917 (N_3917,N_2547,N_2472);
nand U3918 (N_3918,N_2888,N_2272);
nand U3919 (N_3919,N_2420,N_2086);
xor U3920 (N_3920,N_2481,N_2937);
and U3921 (N_3921,N_2644,N_2102);
xnor U3922 (N_3922,N_2289,N_2281);
and U3923 (N_3923,N_2585,N_2675);
xnor U3924 (N_3924,N_2498,N_2251);
xnor U3925 (N_3925,N_2114,N_2728);
or U3926 (N_3926,N_2016,N_2911);
nor U3927 (N_3927,N_2037,N_2768);
xor U3928 (N_3928,N_2589,N_2023);
nor U3929 (N_3929,N_2520,N_2988);
nor U3930 (N_3930,N_2358,N_2111);
and U3931 (N_3931,N_2155,N_2502);
xor U3932 (N_3932,N_2801,N_2819);
and U3933 (N_3933,N_2946,N_2874);
and U3934 (N_3934,N_2708,N_2352);
nand U3935 (N_3935,N_2940,N_2440);
or U3936 (N_3936,N_2612,N_2542);
xnor U3937 (N_3937,N_2865,N_2351);
xor U3938 (N_3938,N_2902,N_2439);
nand U3939 (N_3939,N_2099,N_2612);
nor U3940 (N_3940,N_2264,N_2629);
xor U3941 (N_3941,N_2248,N_2584);
nor U3942 (N_3942,N_2460,N_2696);
xor U3943 (N_3943,N_2605,N_2010);
or U3944 (N_3944,N_2425,N_2290);
nand U3945 (N_3945,N_2649,N_2190);
and U3946 (N_3946,N_2264,N_2845);
and U3947 (N_3947,N_2480,N_2701);
xnor U3948 (N_3948,N_2051,N_2111);
xnor U3949 (N_3949,N_2771,N_2032);
nand U3950 (N_3950,N_2913,N_2117);
nor U3951 (N_3951,N_2596,N_2954);
and U3952 (N_3952,N_2402,N_2390);
nand U3953 (N_3953,N_2012,N_2918);
and U3954 (N_3954,N_2607,N_2831);
and U3955 (N_3955,N_2804,N_2429);
xnor U3956 (N_3956,N_2446,N_2611);
xnor U3957 (N_3957,N_2158,N_2575);
and U3958 (N_3958,N_2720,N_2205);
xor U3959 (N_3959,N_2967,N_2619);
xnor U3960 (N_3960,N_2497,N_2185);
and U3961 (N_3961,N_2552,N_2631);
and U3962 (N_3962,N_2786,N_2035);
nor U3963 (N_3963,N_2294,N_2889);
xor U3964 (N_3964,N_2463,N_2154);
or U3965 (N_3965,N_2986,N_2154);
and U3966 (N_3966,N_2127,N_2470);
and U3967 (N_3967,N_2853,N_2612);
nand U3968 (N_3968,N_2742,N_2854);
nor U3969 (N_3969,N_2384,N_2206);
nor U3970 (N_3970,N_2236,N_2671);
and U3971 (N_3971,N_2197,N_2118);
or U3972 (N_3972,N_2008,N_2899);
nor U3973 (N_3973,N_2090,N_2587);
or U3974 (N_3974,N_2430,N_2920);
xnor U3975 (N_3975,N_2338,N_2850);
xor U3976 (N_3976,N_2080,N_2619);
or U3977 (N_3977,N_2981,N_2203);
nand U3978 (N_3978,N_2570,N_2134);
xnor U3979 (N_3979,N_2583,N_2742);
nor U3980 (N_3980,N_2210,N_2435);
nor U3981 (N_3981,N_2158,N_2691);
nor U3982 (N_3982,N_2740,N_2244);
xor U3983 (N_3983,N_2693,N_2452);
xnor U3984 (N_3984,N_2651,N_2530);
nor U3985 (N_3985,N_2697,N_2241);
nand U3986 (N_3986,N_2041,N_2230);
and U3987 (N_3987,N_2912,N_2531);
nand U3988 (N_3988,N_2621,N_2538);
nand U3989 (N_3989,N_2402,N_2467);
and U3990 (N_3990,N_2941,N_2830);
or U3991 (N_3991,N_2127,N_2756);
xnor U3992 (N_3992,N_2400,N_2708);
or U3993 (N_3993,N_2843,N_2913);
nand U3994 (N_3994,N_2059,N_2461);
nand U3995 (N_3995,N_2819,N_2129);
and U3996 (N_3996,N_2520,N_2361);
xnor U3997 (N_3997,N_2699,N_2449);
nor U3998 (N_3998,N_2060,N_2749);
xor U3999 (N_3999,N_2085,N_2048);
xnor U4000 (N_4000,N_3280,N_3800);
or U4001 (N_4001,N_3552,N_3132);
nor U4002 (N_4002,N_3183,N_3651);
nor U4003 (N_4003,N_3432,N_3283);
nand U4004 (N_4004,N_3475,N_3765);
and U4005 (N_4005,N_3102,N_3399);
xnor U4006 (N_4006,N_3645,N_3181);
or U4007 (N_4007,N_3348,N_3076);
xnor U4008 (N_4008,N_3200,N_3692);
or U4009 (N_4009,N_3070,N_3072);
or U4010 (N_4010,N_3809,N_3203);
nor U4011 (N_4011,N_3665,N_3655);
nand U4012 (N_4012,N_3328,N_3731);
nor U4013 (N_4013,N_3929,N_3184);
nor U4014 (N_4014,N_3504,N_3970);
nor U4015 (N_4015,N_3101,N_3729);
or U4016 (N_4016,N_3855,N_3474);
and U4017 (N_4017,N_3741,N_3327);
and U4018 (N_4018,N_3881,N_3600);
nand U4019 (N_4019,N_3957,N_3247);
nand U4020 (N_4020,N_3927,N_3822);
and U4021 (N_4021,N_3336,N_3361);
or U4022 (N_4022,N_3371,N_3051);
nor U4023 (N_4023,N_3823,N_3798);
and U4024 (N_4024,N_3293,N_3171);
xor U4025 (N_4025,N_3078,N_3392);
nor U4026 (N_4026,N_3398,N_3595);
xor U4027 (N_4027,N_3518,N_3267);
nor U4028 (N_4028,N_3893,N_3004);
and U4029 (N_4029,N_3736,N_3013);
and U4030 (N_4030,N_3923,N_3152);
nor U4031 (N_4031,N_3274,N_3766);
and U4032 (N_4032,N_3945,N_3386);
xnor U4033 (N_4033,N_3786,N_3925);
or U4034 (N_4034,N_3826,N_3614);
or U4035 (N_4035,N_3282,N_3983);
or U4036 (N_4036,N_3611,N_3886);
nand U4037 (N_4037,N_3770,N_3034);
nor U4038 (N_4038,N_3199,N_3060);
nand U4039 (N_4039,N_3795,N_3861);
nand U4040 (N_4040,N_3713,N_3428);
nor U4041 (N_4041,N_3363,N_3951);
xnor U4042 (N_4042,N_3663,N_3458);
and U4043 (N_4043,N_3520,N_3804);
xnor U4044 (N_4044,N_3644,N_3106);
nand U4045 (N_4045,N_3792,N_3757);
or U4046 (N_4046,N_3459,N_3169);
and U4047 (N_4047,N_3571,N_3720);
or U4048 (N_4048,N_3670,N_3472);
nor U4049 (N_4049,N_3216,N_3006);
and U4050 (N_4050,N_3719,N_3674);
and U4051 (N_4051,N_3287,N_3149);
and U4052 (N_4052,N_3960,N_3598);
and U4053 (N_4053,N_3512,N_3576);
nand U4054 (N_4054,N_3605,N_3790);
and U4055 (N_4055,N_3236,N_3637);
or U4056 (N_4056,N_3027,N_3478);
nand U4057 (N_4057,N_3974,N_3862);
nand U4058 (N_4058,N_3867,N_3961);
nand U4059 (N_4059,N_3796,N_3608);
nor U4060 (N_4060,N_3193,N_3639);
nor U4061 (N_4061,N_3439,N_3577);
or U4062 (N_4062,N_3198,N_3094);
nand U4063 (N_4063,N_3710,N_3246);
xor U4064 (N_4064,N_3705,N_3372);
nor U4065 (N_4065,N_3320,N_3926);
nand U4066 (N_4066,N_3108,N_3619);
nor U4067 (N_4067,N_3161,N_3612);
or U4068 (N_4068,N_3462,N_3727);
nor U4069 (N_4069,N_3413,N_3683);
and U4070 (N_4070,N_3388,N_3502);
nor U4071 (N_4071,N_3714,N_3788);
xnor U4072 (N_4072,N_3488,N_3780);
or U4073 (N_4073,N_3671,N_3634);
xnor U4074 (N_4074,N_3163,N_3061);
nor U4075 (N_4075,N_3885,N_3722);
xor U4076 (N_4076,N_3565,N_3699);
xor U4077 (N_4077,N_3105,N_3968);
xnor U4078 (N_4078,N_3418,N_3620);
or U4079 (N_4079,N_3022,N_3650);
nor U4080 (N_4080,N_3299,N_3190);
xor U4081 (N_4081,N_3707,N_3441);
nand U4082 (N_4082,N_3436,N_3421);
and U4083 (N_4083,N_3237,N_3335);
and U4084 (N_4084,N_3584,N_3831);
and U4085 (N_4085,N_3467,N_3024);
and U4086 (N_4086,N_3858,N_3890);
or U4087 (N_4087,N_3684,N_3572);
nor U4088 (N_4088,N_3465,N_3165);
xnor U4089 (N_4089,N_3173,N_3774);
nor U4090 (N_4090,N_3080,N_3219);
nor U4091 (N_4091,N_3025,N_3319);
and U4092 (N_4092,N_3748,N_3365);
nor U4093 (N_4093,N_3658,N_3134);
or U4094 (N_4094,N_3700,N_3450);
nor U4095 (N_4095,N_3672,N_3217);
nand U4096 (N_4096,N_3602,N_3759);
and U4097 (N_4097,N_3207,N_3047);
and U4098 (N_4098,N_3583,N_3669);
or U4099 (N_4099,N_3226,N_3668);
and U4100 (N_4100,N_3001,N_3624);
or U4101 (N_4101,N_3850,N_3121);
and U4102 (N_4102,N_3406,N_3318);
and U4103 (N_4103,N_3784,N_3817);
nand U4104 (N_4104,N_3680,N_3218);
and U4105 (N_4105,N_3677,N_3452);
or U4106 (N_4106,N_3876,N_3843);
nor U4107 (N_4107,N_3625,N_3172);
or U4108 (N_4108,N_3284,N_3836);
xor U4109 (N_4109,N_3701,N_3703);
nand U4110 (N_4110,N_3869,N_3420);
nor U4111 (N_4111,N_3249,N_3980);
xor U4112 (N_4112,N_3995,N_3653);
nand U4113 (N_4113,N_3648,N_3628);
or U4114 (N_4114,N_3411,N_3745);
and U4115 (N_4115,N_3214,N_3863);
and U4116 (N_4116,N_3604,N_3578);
nor U4117 (N_4117,N_3542,N_3548);
and U4118 (N_4118,N_3871,N_3593);
and U4119 (N_4119,N_3021,N_3315);
nand U4120 (N_4120,N_3306,N_3050);
or U4121 (N_4121,N_3894,N_3904);
nor U4122 (N_4122,N_3224,N_3597);
nor U4123 (N_4123,N_3735,N_3239);
nor U4124 (N_4124,N_3381,N_3396);
nand U4125 (N_4125,N_3037,N_3821);
xnor U4126 (N_4126,N_3768,N_3895);
and U4127 (N_4127,N_3730,N_3138);
and U4128 (N_4128,N_3374,N_3939);
nand U4129 (N_4129,N_3148,N_3991);
nand U4130 (N_4130,N_3646,N_3370);
nand U4131 (N_4131,N_3129,N_3401);
and U4132 (N_4132,N_3941,N_3394);
nor U4133 (N_4133,N_3304,N_3607);
or U4134 (N_4134,N_3794,N_3379);
or U4135 (N_4135,N_3908,N_3085);
nor U4136 (N_4136,N_3516,N_3942);
nor U4137 (N_4137,N_3213,N_3801);
and U4138 (N_4138,N_3321,N_3225);
nor U4139 (N_4139,N_3194,N_3263);
and U4140 (N_4140,N_3621,N_3787);
or U4141 (N_4141,N_3545,N_3494);
and U4142 (N_4142,N_3676,N_3296);
or U4143 (N_4143,N_3205,N_3708);
xor U4144 (N_4144,N_3525,N_3055);
or U4145 (N_4145,N_3868,N_3311);
and U4146 (N_4146,N_3258,N_3853);
and U4147 (N_4147,N_3781,N_3573);
xnor U4148 (N_4148,N_3879,N_3551);
xnor U4149 (N_4149,N_3367,N_3984);
xor U4150 (N_4150,N_3709,N_3332);
xnor U4151 (N_4151,N_3938,N_3977);
and U4152 (N_4152,N_3403,N_3301);
nor U4153 (N_4153,N_3291,N_3168);
or U4154 (N_4154,N_3090,N_3039);
nor U4155 (N_4155,N_3081,N_3511);
nor U4156 (N_4156,N_3035,N_3889);
xnor U4157 (N_4157,N_3331,N_3985);
and U4158 (N_4158,N_3206,N_3175);
xor U4159 (N_4159,N_3534,N_3058);
and U4160 (N_4160,N_3350,N_3888);
and U4161 (N_4161,N_3368,N_3726);
nor U4162 (N_4162,N_3967,N_3468);
nand U4163 (N_4163,N_3324,N_3018);
or U4164 (N_4164,N_3240,N_3084);
nor U4165 (N_4165,N_3074,N_3191);
nand U4166 (N_4166,N_3872,N_3587);
nor U4167 (N_4167,N_3753,N_3547);
nand U4168 (N_4168,N_3878,N_3227);
and U4169 (N_4169,N_3498,N_3716);
or U4170 (N_4170,N_3174,N_3965);
or U4171 (N_4171,N_3537,N_3490);
nor U4172 (N_4172,N_3891,N_3979);
and U4173 (N_4173,N_3911,N_3725);
nor U4174 (N_4174,N_3176,N_3414);
nor U4175 (N_4175,N_3717,N_3033);
xnor U4176 (N_4176,N_3223,N_3040);
nand U4177 (N_4177,N_3387,N_3118);
and U4178 (N_4178,N_3443,N_3238);
xnor U4179 (N_4179,N_3845,N_3256);
xnor U4180 (N_4180,N_3844,N_3197);
or U4181 (N_4181,N_3359,N_3896);
xor U4182 (N_4182,N_3752,N_3883);
nand U4183 (N_4183,N_3446,N_3559);
nor U4184 (N_4184,N_3124,N_3662);
and U4185 (N_4185,N_3212,N_3434);
xor U4186 (N_4186,N_3943,N_3640);
and U4187 (N_4187,N_3556,N_3747);
xor U4188 (N_4188,N_3501,N_3698);
nand U4189 (N_4189,N_3603,N_3339);
nand U4190 (N_4190,N_3167,N_3310);
nor U4191 (N_4191,N_3630,N_3999);
xnor U4192 (N_4192,N_3859,N_3931);
or U4193 (N_4193,N_3340,N_3016);
and U4194 (N_4194,N_3917,N_3316);
nand U4195 (N_4195,N_3489,N_3128);
nand U4196 (N_4196,N_3567,N_3048);
nor U4197 (N_4197,N_3570,N_3141);
and U4198 (N_4198,N_3521,N_3812);
xnor U4199 (N_4199,N_3277,N_3629);
xnor U4200 (N_4200,N_3153,N_3417);
and U4201 (N_4201,N_3833,N_3679);
nor U4202 (N_4202,N_3797,N_3987);
and U4203 (N_4203,N_3480,N_3989);
nand U4204 (N_4204,N_3902,N_3425);
nand U4205 (N_4205,N_3632,N_3089);
or U4206 (N_4206,N_3626,N_3453);
nor U4207 (N_4207,N_3649,N_3647);
nand U4208 (N_4208,N_3415,N_3230);
and U4209 (N_4209,N_3011,N_3924);
and U4210 (N_4210,N_3063,N_3535);
nand U4211 (N_4211,N_3043,N_3445);
and U4212 (N_4212,N_3789,N_3131);
and U4213 (N_4213,N_3715,N_3935);
nand U4214 (N_4214,N_3002,N_3373);
and U4215 (N_4215,N_3599,N_3835);
or U4216 (N_4216,N_3816,N_3906);
and U4217 (N_4217,N_3536,N_3248);
nor U4218 (N_4218,N_3732,N_3479);
and U4219 (N_4219,N_3484,N_3507);
xor U4220 (N_4220,N_3322,N_3086);
or U4221 (N_4221,N_3107,N_3229);
nor U4222 (N_4222,N_3111,N_3228);
and U4223 (N_4223,N_3451,N_3146);
nor U4224 (N_4224,N_3666,N_3838);
and U4225 (N_4225,N_3323,N_3366);
nor U4226 (N_4226,N_3519,N_3978);
nand U4227 (N_4227,N_3097,N_3819);
or U4228 (N_4228,N_3738,N_3503);
xor U4229 (N_4229,N_3721,N_3654);
and U4230 (N_4230,N_3342,N_3740);
nor U4231 (N_4231,N_3473,N_3723);
and U4232 (N_4232,N_3338,N_3854);
nor U4233 (N_4233,N_3079,N_3919);
and U4234 (N_4234,N_3245,N_3122);
or U4235 (N_4235,N_3384,N_3075);
xnor U4236 (N_4236,N_3009,N_3652);
or U4237 (N_4237,N_3257,N_3763);
xor U4238 (N_4238,N_3857,N_3279);
or U4239 (N_4239,N_3187,N_3582);
or U4240 (N_4240,N_3591,N_3133);
nor U4241 (N_4241,N_3347,N_3673);
and U4242 (N_4242,N_3864,N_3029);
or U4243 (N_4243,N_3066,N_3986);
xor U4244 (N_4244,N_3325,N_3156);
xnor U4245 (N_4245,N_3966,N_3003);
nor U4246 (N_4246,N_3541,N_3390);
nor U4247 (N_4247,N_3531,N_3581);
nor U4248 (N_4248,N_3073,N_3702);
xnor U4249 (N_4249,N_3364,N_3182);
or U4250 (N_4250,N_3920,N_3631);
nand U4251 (N_4251,N_3356,N_3235);
and U4252 (N_4252,N_3959,N_3114);
nand U4253 (N_4253,N_3463,N_3776);
nand U4254 (N_4254,N_3972,N_3088);
and U4255 (N_4255,N_3346,N_3538);
or U4256 (N_4256,N_3405,N_3271);
and U4257 (N_4257,N_3026,N_3196);
nand U4258 (N_4258,N_3313,N_3554);
nor U4259 (N_4259,N_3592,N_3307);
and U4260 (N_4260,N_3030,N_3259);
nor U4261 (N_4261,N_3476,N_3499);
nand U4262 (N_4262,N_3429,N_3988);
nor U4263 (N_4263,N_3244,N_3496);
or U4264 (N_4264,N_3492,N_3433);
and U4265 (N_4265,N_3527,N_3273);
nor U4266 (N_4266,N_3234,N_3136);
or U4267 (N_4267,N_3686,N_3937);
nand U4268 (N_4268,N_3355,N_3529);
xor U4269 (N_4269,N_3380,N_3793);
nor U4270 (N_4270,N_3201,N_3743);
nand U4271 (N_4271,N_3241,N_3157);
nor U4272 (N_4272,N_3948,N_3145);
nor U4273 (N_4273,N_3290,N_3082);
or U4274 (N_4274,N_3481,N_3918);
or U4275 (N_4275,N_3694,N_3160);
or U4276 (N_4276,N_3815,N_3278);
or U4277 (N_4277,N_3285,N_3155);
nor U4278 (N_4278,N_3456,N_3378);
nand U4279 (N_4279,N_3555,N_3294);
and U4280 (N_4280,N_3358,N_3982);
or U4281 (N_4281,N_3659,N_3762);
and U4282 (N_4282,N_3546,N_3195);
xnor U4283 (N_4283,N_3375,N_3773);
or U4284 (N_4284,N_3882,N_3427);
xor U4285 (N_4285,N_3549,N_3360);
nand U4286 (N_4286,N_3471,N_3772);
nor U4287 (N_4287,N_3964,N_3955);
and U4288 (N_4288,N_3849,N_3408);
or U4289 (N_4289,N_3007,N_3934);
nor U4290 (N_4290,N_3954,N_3297);
nor U4291 (N_4291,N_3588,N_3352);
nor U4292 (N_4292,N_3712,N_3903);
nor U4293 (N_4293,N_3117,N_3949);
nor U4294 (N_4294,N_3750,N_3261);
or U4295 (N_4295,N_3564,N_3901);
or U4296 (N_4296,N_3431,N_3834);
and U4297 (N_4297,N_3276,N_3973);
and U4298 (N_4298,N_3691,N_3761);
nor U4299 (N_4299,N_3343,N_3664);
nor U4300 (N_4300,N_3963,N_3505);
and U4301 (N_4301,N_3349,N_3820);
and U4302 (N_4302,N_3522,N_3020);
xnor U4303 (N_4303,N_3438,N_3211);
or U4304 (N_4304,N_3272,N_3870);
nand U4305 (N_4305,N_3553,N_3326);
and U4306 (N_4306,N_3933,N_3341);
and U4307 (N_4307,N_3144,N_3760);
or U4308 (N_4308,N_3460,N_3469);
nor U4309 (N_4309,N_3435,N_3936);
xor U4310 (N_4310,N_3220,N_3756);
nand U4311 (N_4311,N_3046,N_3667);
and U4312 (N_4312,N_3779,N_3540);
nor U4313 (N_4313,N_3910,N_3569);
nand U4314 (N_4314,N_3265,N_3015);
and U4315 (N_4315,N_3574,N_3830);
nor U4316 (N_4316,N_3251,N_3744);
nand U4317 (N_4317,N_3302,N_3126);
nand U4318 (N_4318,N_3814,N_3231);
nand U4319 (N_4319,N_3579,N_3091);
nor U4320 (N_4320,N_3609,N_3580);
xnor U4321 (N_4321,N_3693,N_3877);
nand U4322 (N_4322,N_3110,N_3533);
or U4323 (N_4323,N_3103,N_3696);
or U4324 (N_4324,N_3104,N_3135);
and U4325 (N_4325,N_3192,N_3281);
nor U4326 (N_4326,N_3866,N_3014);
or U4327 (N_4327,N_3179,N_3049);
or U4328 (N_4328,N_3455,N_3028);
or U4329 (N_4329,N_3695,N_3164);
nand U4330 (N_4330,N_3589,N_3594);
nand U4331 (N_4331,N_3897,N_3054);
nor U4332 (N_4332,N_3706,N_3158);
or U4333 (N_4333,N_3487,N_3068);
or U4334 (N_4334,N_3847,N_3286);
and U4335 (N_4335,N_3586,N_3932);
nand U4336 (N_4336,N_3269,N_3170);
and U4337 (N_4337,N_3791,N_3383);
and U4338 (N_4338,N_3517,N_3288);
nor U4339 (N_4339,N_3099,N_3312);
or U4340 (N_4340,N_3958,N_3407);
or U4341 (N_4341,N_3921,N_3242);
xor U4342 (N_4342,N_3852,N_3333);
xor U4343 (N_4343,N_3530,N_3243);
nand U4344 (N_4344,N_3113,N_3777);
nor U4345 (N_4345,N_3617,N_3746);
nand U4346 (N_4346,N_3975,N_3642);
nand U4347 (N_4347,N_3395,N_3742);
nand U4348 (N_4348,N_3946,N_3430);
nand U4349 (N_4349,N_3444,N_3147);
and U4350 (N_4350,N_3940,N_3539);
xnor U4351 (N_4351,N_3657,N_3806);
nand U4352 (N_4352,N_3127,N_3440);
and U4353 (N_4353,N_3253,N_3514);
nand U4354 (N_4354,N_3874,N_3802);
xor U4355 (N_4355,N_3208,N_3907);
xor U4356 (N_4356,N_3012,N_3532);
or U4357 (N_4357,N_3067,N_3807);
xor U4358 (N_4358,N_3221,N_3887);
nand U4359 (N_4359,N_3391,N_3769);
and U4360 (N_4360,N_3252,N_3329);
nor U4361 (N_4361,N_3064,N_3397);
and U4362 (N_4362,N_3944,N_3485);
nor U4363 (N_4363,N_3947,N_3210);
xor U4364 (N_4364,N_3305,N_3426);
nand U4365 (N_4365,N_3083,N_3660);
and U4366 (N_4366,N_3180,N_3856);
nand U4367 (N_4367,N_3019,N_3005);
and U4368 (N_4368,N_3204,N_3185);
xor U4369 (N_4369,N_3601,N_3828);
xnor U4370 (N_4370,N_3875,N_3803);
or U4371 (N_4371,N_3513,N_3087);
or U4372 (N_4372,N_3615,N_3410);
nand U4373 (N_4373,N_3733,N_3300);
and U4374 (N_4374,N_3448,N_3262);
nor U4375 (N_4375,N_3275,N_3841);
nand U4376 (N_4376,N_3656,N_3354);
nor U4377 (N_4377,N_3913,N_3053);
nor U4378 (N_4378,N_3402,N_3873);
or U4379 (N_4379,N_3357,N_3996);
or U4380 (N_4380,N_3568,N_3317);
xnor U4381 (N_4381,N_3865,N_3848);
or U4382 (N_4382,N_3486,N_3233);
and U4383 (N_4383,N_3728,N_3497);
nand U4384 (N_4384,N_3162,N_3880);
nand U4385 (N_4385,N_3376,N_3767);
xor U4386 (N_4386,N_3557,N_3998);
nor U4387 (N_4387,N_3098,N_3641);
xor U4388 (N_4388,N_3093,N_3524);
xor U4389 (N_4389,N_3618,N_3308);
or U4390 (N_4390,N_3337,N_3523);
nand U4391 (N_4391,N_3116,N_3560);
xnor U4392 (N_4392,N_3851,N_3596);
nand U4393 (N_4393,N_3832,N_3898);
and U4394 (N_4394,N_3412,N_3825);
and U4395 (N_4395,N_3404,N_3045);
nor U4396 (N_4396,N_3369,N_3032);
or U4397 (N_4397,N_3056,N_3751);
and U4398 (N_4398,N_3254,N_3334);
and U4399 (N_4399,N_3997,N_3096);
or U4400 (N_4400,N_3330,N_3457);
and U4401 (N_4401,N_3992,N_3689);
and U4402 (N_4402,N_3295,N_3092);
or U4403 (N_4403,N_3260,N_3697);
nor U4404 (N_4404,N_3508,N_3860);
xor U4405 (N_4405,N_3749,N_3956);
xnor U4406 (N_4406,N_3052,N_3976);
or U4407 (N_4407,N_3962,N_3813);
nor U4408 (N_4408,N_3590,N_3437);
nor U4409 (N_4409,N_3466,N_3805);
nor U4410 (N_4410,N_3351,N_3119);
and U4411 (N_4411,N_3447,N_3755);
nand U4412 (N_4412,N_3041,N_3303);
xnor U4413 (N_4413,N_3635,N_3678);
nor U4414 (N_4414,N_3264,N_3031);
nor U4415 (N_4415,N_3829,N_3345);
or U4416 (N_4416,N_3385,N_3177);
or U4417 (N_4417,N_3069,N_3362);
xor U4418 (N_4418,N_3142,N_3509);
nand U4419 (N_4419,N_3682,N_3950);
nor U4420 (N_4420,N_3528,N_3289);
and U4421 (N_4421,N_3151,N_3685);
nand U4422 (N_4422,N_3166,N_3255);
nand U4423 (N_4423,N_3419,N_3930);
nand U4424 (N_4424,N_3491,N_3400);
or U4425 (N_4425,N_3495,N_3266);
or U4426 (N_4426,N_3842,N_3922);
nor U4427 (N_4427,N_3544,N_3688);
nand U4428 (N_4428,N_3928,N_3482);
or U4429 (N_4429,N_3892,N_3506);
or U4430 (N_4430,N_3000,N_3818);
or U4431 (N_4431,N_3232,N_3899);
xnor U4432 (N_4432,N_3042,N_3675);
and U4433 (N_4433,N_3178,N_3298);
or U4434 (N_4434,N_3140,N_3734);
nand U4435 (N_4435,N_3477,N_3969);
or U4436 (N_4436,N_3077,N_3008);
nor U4437 (N_4437,N_3139,N_3017);
or U4438 (N_4438,N_3981,N_3159);
nand U4439 (N_4439,N_3915,N_3449);
xor U4440 (N_4440,N_3754,N_3309);
xor U4441 (N_4441,N_3704,N_3561);
and U4442 (N_4442,N_3125,N_3764);
nand U4443 (N_4443,N_3799,N_3130);
xor U4444 (N_4444,N_3739,N_3344);
nand U4445 (N_4445,N_3515,N_3643);
nand U4446 (N_4446,N_3423,N_3377);
nor U4447 (N_4447,N_3454,N_3353);
or U4448 (N_4448,N_3095,N_3771);
and U4449 (N_4449,N_3827,N_3994);
nand U4450 (N_4450,N_3038,N_3057);
xnor U4451 (N_4451,N_3464,N_3470);
xnor U4452 (N_4452,N_3036,N_3627);
nand U4453 (N_4453,N_3824,N_3202);
and U4454 (N_4454,N_3785,N_3839);
and U4455 (N_4455,N_3566,N_3737);
nand U4456 (N_4456,N_3416,N_3209);
nor U4457 (N_4457,N_3023,N_3222);
xor U4458 (N_4458,N_3613,N_3846);
xnor U4459 (N_4459,N_3562,N_3188);
and U4460 (N_4460,N_3585,N_3150);
and U4461 (N_4461,N_3952,N_3575);
nand U4462 (N_4462,N_3550,N_3112);
nand U4463 (N_4463,N_3971,N_3993);
nor U4464 (N_4464,N_3758,N_3840);
and U4465 (N_4465,N_3724,N_3914);
nand U4466 (N_4466,N_3912,N_3681);
nand U4467 (N_4467,N_3616,N_3493);
and U4468 (N_4468,N_3044,N_3558);
xnor U4469 (N_4469,N_3783,N_3461);
or U4470 (N_4470,N_3510,N_3143);
or U4471 (N_4471,N_3409,N_3884);
nand U4472 (N_4472,N_3215,N_3382);
or U4473 (N_4473,N_3610,N_3661);
and U4474 (N_4474,N_3109,N_3189);
nand U4475 (N_4475,N_3483,N_3010);
and U4476 (N_4476,N_3442,N_3186);
and U4477 (N_4477,N_3810,N_3718);
and U4478 (N_4478,N_3292,N_3953);
or U4479 (N_4479,N_3622,N_3389);
nor U4480 (N_4480,N_3120,N_3314);
nor U4481 (N_4481,N_3623,N_3990);
nand U4482 (N_4482,N_3268,N_3062);
nor U4483 (N_4483,N_3775,N_3422);
nor U4484 (N_4484,N_3543,N_3778);
xnor U4485 (N_4485,N_3606,N_3123);
nor U4486 (N_4486,N_3100,N_3526);
xnor U4487 (N_4487,N_3638,N_3905);
nand U4488 (N_4488,N_3808,N_3500);
and U4489 (N_4489,N_3687,N_3811);
and U4490 (N_4490,N_3059,N_3633);
nand U4491 (N_4491,N_3270,N_3071);
or U4492 (N_4492,N_3250,N_3900);
and U4493 (N_4493,N_3636,N_3690);
nand U4494 (N_4494,N_3393,N_3711);
xnor U4495 (N_4495,N_3065,N_3424);
and U4496 (N_4496,N_3154,N_3563);
xnor U4497 (N_4497,N_3115,N_3782);
and U4498 (N_4498,N_3909,N_3916);
nor U4499 (N_4499,N_3837,N_3137);
nor U4500 (N_4500,N_3173,N_3302);
or U4501 (N_4501,N_3620,N_3524);
and U4502 (N_4502,N_3811,N_3981);
nor U4503 (N_4503,N_3593,N_3633);
xnor U4504 (N_4504,N_3516,N_3116);
nand U4505 (N_4505,N_3019,N_3764);
xor U4506 (N_4506,N_3193,N_3492);
and U4507 (N_4507,N_3312,N_3866);
and U4508 (N_4508,N_3005,N_3180);
nor U4509 (N_4509,N_3891,N_3963);
nand U4510 (N_4510,N_3215,N_3300);
nand U4511 (N_4511,N_3041,N_3271);
xnor U4512 (N_4512,N_3976,N_3568);
and U4513 (N_4513,N_3108,N_3448);
xor U4514 (N_4514,N_3275,N_3348);
or U4515 (N_4515,N_3227,N_3436);
or U4516 (N_4516,N_3929,N_3506);
and U4517 (N_4517,N_3474,N_3829);
xnor U4518 (N_4518,N_3100,N_3857);
nor U4519 (N_4519,N_3357,N_3289);
nand U4520 (N_4520,N_3507,N_3534);
xor U4521 (N_4521,N_3866,N_3801);
nor U4522 (N_4522,N_3340,N_3993);
nand U4523 (N_4523,N_3402,N_3593);
and U4524 (N_4524,N_3868,N_3316);
nand U4525 (N_4525,N_3657,N_3650);
or U4526 (N_4526,N_3929,N_3084);
nor U4527 (N_4527,N_3578,N_3906);
nand U4528 (N_4528,N_3238,N_3153);
nand U4529 (N_4529,N_3665,N_3009);
nor U4530 (N_4530,N_3843,N_3942);
nand U4531 (N_4531,N_3232,N_3345);
nand U4532 (N_4532,N_3858,N_3072);
nor U4533 (N_4533,N_3501,N_3523);
xor U4534 (N_4534,N_3705,N_3776);
nor U4535 (N_4535,N_3561,N_3466);
nor U4536 (N_4536,N_3015,N_3381);
or U4537 (N_4537,N_3422,N_3739);
nor U4538 (N_4538,N_3568,N_3400);
xnor U4539 (N_4539,N_3518,N_3234);
nand U4540 (N_4540,N_3087,N_3577);
xnor U4541 (N_4541,N_3751,N_3766);
xor U4542 (N_4542,N_3726,N_3837);
or U4543 (N_4543,N_3275,N_3388);
nand U4544 (N_4544,N_3699,N_3611);
nor U4545 (N_4545,N_3719,N_3950);
nand U4546 (N_4546,N_3240,N_3495);
xor U4547 (N_4547,N_3299,N_3538);
and U4548 (N_4548,N_3372,N_3865);
or U4549 (N_4549,N_3383,N_3431);
or U4550 (N_4550,N_3761,N_3768);
nor U4551 (N_4551,N_3619,N_3210);
nor U4552 (N_4552,N_3488,N_3782);
xor U4553 (N_4553,N_3694,N_3747);
or U4554 (N_4554,N_3499,N_3865);
or U4555 (N_4555,N_3532,N_3552);
and U4556 (N_4556,N_3894,N_3858);
nor U4557 (N_4557,N_3338,N_3646);
or U4558 (N_4558,N_3921,N_3410);
nor U4559 (N_4559,N_3917,N_3741);
or U4560 (N_4560,N_3089,N_3742);
xor U4561 (N_4561,N_3307,N_3602);
xnor U4562 (N_4562,N_3196,N_3434);
nand U4563 (N_4563,N_3923,N_3078);
nand U4564 (N_4564,N_3108,N_3396);
nor U4565 (N_4565,N_3493,N_3283);
xor U4566 (N_4566,N_3222,N_3983);
nand U4567 (N_4567,N_3603,N_3287);
nand U4568 (N_4568,N_3792,N_3433);
nand U4569 (N_4569,N_3787,N_3318);
and U4570 (N_4570,N_3068,N_3896);
nor U4571 (N_4571,N_3257,N_3064);
xnor U4572 (N_4572,N_3772,N_3544);
and U4573 (N_4573,N_3102,N_3825);
nor U4574 (N_4574,N_3668,N_3373);
xor U4575 (N_4575,N_3737,N_3246);
nand U4576 (N_4576,N_3085,N_3913);
xor U4577 (N_4577,N_3547,N_3133);
or U4578 (N_4578,N_3057,N_3907);
nor U4579 (N_4579,N_3708,N_3754);
nor U4580 (N_4580,N_3175,N_3517);
and U4581 (N_4581,N_3786,N_3845);
nand U4582 (N_4582,N_3880,N_3293);
nor U4583 (N_4583,N_3634,N_3708);
nor U4584 (N_4584,N_3038,N_3462);
nor U4585 (N_4585,N_3346,N_3789);
xnor U4586 (N_4586,N_3071,N_3311);
or U4587 (N_4587,N_3575,N_3092);
xnor U4588 (N_4588,N_3459,N_3584);
xnor U4589 (N_4589,N_3709,N_3333);
or U4590 (N_4590,N_3728,N_3705);
and U4591 (N_4591,N_3160,N_3409);
xor U4592 (N_4592,N_3842,N_3752);
nand U4593 (N_4593,N_3194,N_3058);
nand U4594 (N_4594,N_3849,N_3547);
and U4595 (N_4595,N_3255,N_3394);
and U4596 (N_4596,N_3854,N_3560);
or U4597 (N_4597,N_3566,N_3271);
and U4598 (N_4598,N_3988,N_3851);
or U4599 (N_4599,N_3170,N_3835);
xnor U4600 (N_4600,N_3042,N_3071);
xnor U4601 (N_4601,N_3967,N_3151);
xnor U4602 (N_4602,N_3468,N_3139);
or U4603 (N_4603,N_3059,N_3227);
nand U4604 (N_4604,N_3957,N_3089);
or U4605 (N_4605,N_3982,N_3059);
and U4606 (N_4606,N_3803,N_3357);
and U4607 (N_4607,N_3537,N_3547);
xor U4608 (N_4608,N_3021,N_3019);
or U4609 (N_4609,N_3924,N_3332);
nor U4610 (N_4610,N_3269,N_3547);
and U4611 (N_4611,N_3476,N_3248);
nand U4612 (N_4612,N_3526,N_3758);
nand U4613 (N_4613,N_3829,N_3940);
and U4614 (N_4614,N_3753,N_3453);
xnor U4615 (N_4615,N_3426,N_3752);
nor U4616 (N_4616,N_3028,N_3467);
nand U4617 (N_4617,N_3826,N_3748);
nand U4618 (N_4618,N_3317,N_3255);
xnor U4619 (N_4619,N_3209,N_3226);
nand U4620 (N_4620,N_3081,N_3876);
and U4621 (N_4621,N_3063,N_3421);
or U4622 (N_4622,N_3378,N_3488);
and U4623 (N_4623,N_3694,N_3994);
nand U4624 (N_4624,N_3308,N_3265);
and U4625 (N_4625,N_3502,N_3773);
nand U4626 (N_4626,N_3231,N_3088);
nand U4627 (N_4627,N_3036,N_3301);
or U4628 (N_4628,N_3258,N_3038);
xnor U4629 (N_4629,N_3916,N_3114);
xnor U4630 (N_4630,N_3531,N_3703);
nor U4631 (N_4631,N_3503,N_3124);
nand U4632 (N_4632,N_3197,N_3640);
nor U4633 (N_4633,N_3804,N_3806);
or U4634 (N_4634,N_3588,N_3259);
nor U4635 (N_4635,N_3431,N_3258);
nor U4636 (N_4636,N_3735,N_3947);
and U4637 (N_4637,N_3250,N_3577);
or U4638 (N_4638,N_3413,N_3881);
or U4639 (N_4639,N_3663,N_3796);
nand U4640 (N_4640,N_3933,N_3514);
nor U4641 (N_4641,N_3020,N_3304);
or U4642 (N_4642,N_3838,N_3607);
and U4643 (N_4643,N_3202,N_3050);
nand U4644 (N_4644,N_3866,N_3526);
and U4645 (N_4645,N_3511,N_3348);
nand U4646 (N_4646,N_3028,N_3910);
xnor U4647 (N_4647,N_3940,N_3484);
xor U4648 (N_4648,N_3724,N_3038);
xor U4649 (N_4649,N_3816,N_3936);
or U4650 (N_4650,N_3443,N_3047);
and U4651 (N_4651,N_3678,N_3248);
and U4652 (N_4652,N_3068,N_3913);
xnor U4653 (N_4653,N_3999,N_3881);
and U4654 (N_4654,N_3820,N_3645);
nand U4655 (N_4655,N_3175,N_3434);
xnor U4656 (N_4656,N_3996,N_3894);
nand U4657 (N_4657,N_3533,N_3521);
or U4658 (N_4658,N_3916,N_3207);
nor U4659 (N_4659,N_3671,N_3165);
nor U4660 (N_4660,N_3322,N_3261);
and U4661 (N_4661,N_3391,N_3091);
or U4662 (N_4662,N_3596,N_3361);
nor U4663 (N_4663,N_3645,N_3499);
or U4664 (N_4664,N_3489,N_3570);
or U4665 (N_4665,N_3995,N_3309);
nand U4666 (N_4666,N_3578,N_3138);
and U4667 (N_4667,N_3771,N_3821);
or U4668 (N_4668,N_3007,N_3386);
nand U4669 (N_4669,N_3462,N_3107);
nand U4670 (N_4670,N_3900,N_3488);
xnor U4671 (N_4671,N_3259,N_3846);
and U4672 (N_4672,N_3716,N_3488);
xnor U4673 (N_4673,N_3472,N_3722);
or U4674 (N_4674,N_3334,N_3290);
nand U4675 (N_4675,N_3725,N_3394);
or U4676 (N_4676,N_3514,N_3426);
nand U4677 (N_4677,N_3342,N_3628);
nand U4678 (N_4678,N_3795,N_3785);
or U4679 (N_4679,N_3937,N_3609);
nor U4680 (N_4680,N_3614,N_3182);
nor U4681 (N_4681,N_3716,N_3516);
xnor U4682 (N_4682,N_3306,N_3108);
nand U4683 (N_4683,N_3834,N_3927);
nor U4684 (N_4684,N_3240,N_3835);
nor U4685 (N_4685,N_3311,N_3554);
nor U4686 (N_4686,N_3656,N_3446);
or U4687 (N_4687,N_3657,N_3161);
and U4688 (N_4688,N_3627,N_3259);
or U4689 (N_4689,N_3557,N_3493);
xnor U4690 (N_4690,N_3234,N_3236);
nand U4691 (N_4691,N_3646,N_3305);
nor U4692 (N_4692,N_3757,N_3728);
and U4693 (N_4693,N_3364,N_3717);
xor U4694 (N_4694,N_3261,N_3053);
nand U4695 (N_4695,N_3011,N_3415);
xor U4696 (N_4696,N_3756,N_3801);
nand U4697 (N_4697,N_3466,N_3727);
and U4698 (N_4698,N_3627,N_3034);
or U4699 (N_4699,N_3182,N_3077);
nor U4700 (N_4700,N_3698,N_3282);
nor U4701 (N_4701,N_3017,N_3941);
xnor U4702 (N_4702,N_3787,N_3643);
xor U4703 (N_4703,N_3260,N_3414);
or U4704 (N_4704,N_3883,N_3763);
or U4705 (N_4705,N_3912,N_3742);
xnor U4706 (N_4706,N_3940,N_3723);
or U4707 (N_4707,N_3533,N_3157);
nor U4708 (N_4708,N_3838,N_3092);
or U4709 (N_4709,N_3315,N_3176);
nand U4710 (N_4710,N_3879,N_3185);
nor U4711 (N_4711,N_3505,N_3436);
or U4712 (N_4712,N_3414,N_3637);
nand U4713 (N_4713,N_3271,N_3236);
xor U4714 (N_4714,N_3136,N_3268);
nor U4715 (N_4715,N_3943,N_3944);
xor U4716 (N_4716,N_3698,N_3362);
xor U4717 (N_4717,N_3148,N_3798);
and U4718 (N_4718,N_3530,N_3534);
and U4719 (N_4719,N_3248,N_3268);
and U4720 (N_4720,N_3669,N_3910);
nor U4721 (N_4721,N_3428,N_3040);
nand U4722 (N_4722,N_3346,N_3855);
xor U4723 (N_4723,N_3875,N_3267);
nand U4724 (N_4724,N_3522,N_3508);
nor U4725 (N_4725,N_3449,N_3001);
and U4726 (N_4726,N_3569,N_3555);
or U4727 (N_4727,N_3565,N_3762);
xnor U4728 (N_4728,N_3667,N_3011);
or U4729 (N_4729,N_3176,N_3756);
or U4730 (N_4730,N_3631,N_3356);
xnor U4731 (N_4731,N_3358,N_3546);
or U4732 (N_4732,N_3154,N_3846);
and U4733 (N_4733,N_3460,N_3230);
nand U4734 (N_4734,N_3782,N_3277);
or U4735 (N_4735,N_3180,N_3332);
nand U4736 (N_4736,N_3229,N_3165);
or U4737 (N_4737,N_3161,N_3805);
and U4738 (N_4738,N_3589,N_3824);
nand U4739 (N_4739,N_3285,N_3400);
nand U4740 (N_4740,N_3649,N_3760);
xnor U4741 (N_4741,N_3957,N_3942);
xor U4742 (N_4742,N_3608,N_3880);
and U4743 (N_4743,N_3690,N_3018);
nor U4744 (N_4744,N_3178,N_3347);
nor U4745 (N_4745,N_3217,N_3389);
nand U4746 (N_4746,N_3613,N_3209);
and U4747 (N_4747,N_3079,N_3548);
or U4748 (N_4748,N_3294,N_3999);
nor U4749 (N_4749,N_3374,N_3305);
or U4750 (N_4750,N_3055,N_3565);
xnor U4751 (N_4751,N_3905,N_3267);
nor U4752 (N_4752,N_3396,N_3101);
xor U4753 (N_4753,N_3421,N_3481);
xnor U4754 (N_4754,N_3896,N_3728);
nand U4755 (N_4755,N_3705,N_3228);
or U4756 (N_4756,N_3492,N_3365);
nand U4757 (N_4757,N_3956,N_3664);
and U4758 (N_4758,N_3351,N_3475);
nor U4759 (N_4759,N_3921,N_3956);
or U4760 (N_4760,N_3971,N_3220);
xor U4761 (N_4761,N_3134,N_3756);
and U4762 (N_4762,N_3324,N_3849);
nand U4763 (N_4763,N_3159,N_3689);
nand U4764 (N_4764,N_3592,N_3928);
or U4765 (N_4765,N_3123,N_3037);
or U4766 (N_4766,N_3544,N_3953);
xnor U4767 (N_4767,N_3638,N_3236);
nand U4768 (N_4768,N_3603,N_3803);
nand U4769 (N_4769,N_3012,N_3392);
nand U4770 (N_4770,N_3208,N_3553);
nand U4771 (N_4771,N_3169,N_3537);
nor U4772 (N_4772,N_3653,N_3374);
or U4773 (N_4773,N_3889,N_3192);
nand U4774 (N_4774,N_3540,N_3134);
xor U4775 (N_4775,N_3772,N_3381);
xor U4776 (N_4776,N_3752,N_3517);
or U4777 (N_4777,N_3089,N_3154);
xnor U4778 (N_4778,N_3307,N_3979);
xor U4779 (N_4779,N_3715,N_3552);
nand U4780 (N_4780,N_3142,N_3924);
nor U4781 (N_4781,N_3354,N_3550);
and U4782 (N_4782,N_3311,N_3728);
xnor U4783 (N_4783,N_3562,N_3918);
nor U4784 (N_4784,N_3952,N_3793);
or U4785 (N_4785,N_3880,N_3177);
xor U4786 (N_4786,N_3151,N_3424);
nor U4787 (N_4787,N_3936,N_3337);
and U4788 (N_4788,N_3398,N_3179);
nor U4789 (N_4789,N_3488,N_3198);
or U4790 (N_4790,N_3282,N_3507);
nand U4791 (N_4791,N_3227,N_3596);
and U4792 (N_4792,N_3774,N_3878);
nor U4793 (N_4793,N_3353,N_3552);
nand U4794 (N_4794,N_3284,N_3998);
or U4795 (N_4795,N_3351,N_3594);
nand U4796 (N_4796,N_3371,N_3030);
xor U4797 (N_4797,N_3460,N_3382);
and U4798 (N_4798,N_3458,N_3763);
xor U4799 (N_4799,N_3515,N_3107);
nand U4800 (N_4800,N_3230,N_3257);
xor U4801 (N_4801,N_3300,N_3798);
and U4802 (N_4802,N_3688,N_3459);
and U4803 (N_4803,N_3522,N_3304);
nand U4804 (N_4804,N_3856,N_3137);
xnor U4805 (N_4805,N_3027,N_3468);
nand U4806 (N_4806,N_3846,N_3871);
and U4807 (N_4807,N_3740,N_3953);
nand U4808 (N_4808,N_3604,N_3159);
and U4809 (N_4809,N_3609,N_3443);
nand U4810 (N_4810,N_3499,N_3697);
or U4811 (N_4811,N_3999,N_3771);
or U4812 (N_4812,N_3807,N_3138);
or U4813 (N_4813,N_3518,N_3537);
xor U4814 (N_4814,N_3680,N_3205);
or U4815 (N_4815,N_3574,N_3710);
nand U4816 (N_4816,N_3996,N_3352);
and U4817 (N_4817,N_3502,N_3360);
or U4818 (N_4818,N_3142,N_3040);
xnor U4819 (N_4819,N_3351,N_3649);
nand U4820 (N_4820,N_3606,N_3598);
or U4821 (N_4821,N_3909,N_3252);
or U4822 (N_4822,N_3354,N_3107);
or U4823 (N_4823,N_3273,N_3885);
xor U4824 (N_4824,N_3169,N_3805);
or U4825 (N_4825,N_3982,N_3917);
xor U4826 (N_4826,N_3146,N_3622);
and U4827 (N_4827,N_3772,N_3248);
nand U4828 (N_4828,N_3493,N_3054);
nand U4829 (N_4829,N_3094,N_3559);
or U4830 (N_4830,N_3844,N_3610);
nor U4831 (N_4831,N_3164,N_3184);
or U4832 (N_4832,N_3115,N_3064);
nor U4833 (N_4833,N_3732,N_3498);
nor U4834 (N_4834,N_3230,N_3430);
or U4835 (N_4835,N_3483,N_3247);
and U4836 (N_4836,N_3402,N_3950);
nor U4837 (N_4837,N_3723,N_3457);
xnor U4838 (N_4838,N_3823,N_3792);
and U4839 (N_4839,N_3145,N_3799);
nand U4840 (N_4840,N_3480,N_3841);
and U4841 (N_4841,N_3805,N_3352);
or U4842 (N_4842,N_3166,N_3178);
nor U4843 (N_4843,N_3096,N_3731);
xor U4844 (N_4844,N_3822,N_3021);
nor U4845 (N_4845,N_3613,N_3506);
or U4846 (N_4846,N_3918,N_3821);
and U4847 (N_4847,N_3828,N_3045);
nand U4848 (N_4848,N_3146,N_3410);
and U4849 (N_4849,N_3005,N_3511);
and U4850 (N_4850,N_3181,N_3580);
xnor U4851 (N_4851,N_3351,N_3310);
xnor U4852 (N_4852,N_3655,N_3188);
and U4853 (N_4853,N_3654,N_3442);
nor U4854 (N_4854,N_3434,N_3405);
nand U4855 (N_4855,N_3850,N_3144);
xnor U4856 (N_4856,N_3080,N_3718);
nor U4857 (N_4857,N_3431,N_3731);
nor U4858 (N_4858,N_3401,N_3585);
or U4859 (N_4859,N_3332,N_3952);
xnor U4860 (N_4860,N_3246,N_3900);
nand U4861 (N_4861,N_3140,N_3122);
nor U4862 (N_4862,N_3894,N_3643);
xnor U4863 (N_4863,N_3854,N_3075);
or U4864 (N_4864,N_3057,N_3720);
nand U4865 (N_4865,N_3624,N_3673);
nor U4866 (N_4866,N_3551,N_3902);
nand U4867 (N_4867,N_3652,N_3314);
and U4868 (N_4868,N_3275,N_3615);
nor U4869 (N_4869,N_3328,N_3019);
nor U4870 (N_4870,N_3104,N_3751);
nor U4871 (N_4871,N_3335,N_3484);
nand U4872 (N_4872,N_3933,N_3531);
and U4873 (N_4873,N_3883,N_3077);
nand U4874 (N_4874,N_3685,N_3215);
nand U4875 (N_4875,N_3702,N_3128);
nor U4876 (N_4876,N_3042,N_3649);
or U4877 (N_4877,N_3835,N_3860);
or U4878 (N_4878,N_3153,N_3918);
and U4879 (N_4879,N_3000,N_3451);
xor U4880 (N_4880,N_3524,N_3247);
nand U4881 (N_4881,N_3787,N_3834);
nand U4882 (N_4882,N_3313,N_3943);
nor U4883 (N_4883,N_3258,N_3333);
nor U4884 (N_4884,N_3137,N_3398);
nor U4885 (N_4885,N_3531,N_3067);
xor U4886 (N_4886,N_3607,N_3652);
xnor U4887 (N_4887,N_3006,N_3065);
and U4888 (N_4888,N_3304,N_3115);
xnor U4889 (N_4889,N_3234,N_3423);
xor U4890 (N_4890,N_3738,N_3768);
nand U4891 (N_4891,N_3894,N_3311);
and U4892 (N_4892,N_3474,N_3934);
nor U4893 (N_4893,N_3087,N_3657);
nand U4894 (N_4894,N_3903,N_3877);
or U4895 (N_4895,N_3522,N_3917);
and U4896 (N_4896,N_3580,N_3836);
and U4897 (N_4897,N_3377,N_3190);
and U4898 (N_4898,N_3884,N_3612);
nor U4899 (N_4899,N_3498,N_3402);
or U4900 (N_4900,N_3402,N_3836);
and U4901 (N_4901,N_3516,N_3677);
and U4902 (N_4902,N_3383,N_3201);
and U4903 (N_4903,N_3886,N_3918);
nor U4904 (N_4904,N_3262,N_3283);
or U4905 (N_4905,N_3742,N_3980);
xnor U4906 (N_4906,N_3065,N_3892);
xnor U4907 (N_4907,N_3061,N_3317);
and U4908 (N_4908,N_3115,N_3399);
xnor U4909 (N_4909,N_3957,N_3749);
and U4910 (N_4910,N_3080,N_3828);
nor U4911 (N_4911,N_3974,N_3216);
nor U4912 (N_4912,N_3478,N_3796);
nand U4913 (N_4913,N_3626,N_3322);
nand U4914 (N_4914,N_3356,N_3937);
nor U4915 (N_4915,N_3756,N_3166);
nor U4916 (N_4916,N_3459,N_3060);
and U4917 (N_4917,N_3122,N_3614);
and U4918 (N_4918,N_3412,N_3491);
nand U4919 (N_4919,N_3458,N_3861);
and U4920 (N_4920,N_3921,N_3543);
and U4921 (N_4921,N_3627,N_3131);
nor U4922 (N_4922,N_3814,N_3315);
xnor U4923 (N_4923,N_3068,N_3225);
nor U4924 (N_4924,N_3909,N_3882);
nor U4925 (N_4925,N_3301,N_3878);
and U4926 (N_4926,N_3072,N_3992);
nor U4927 (N_4927,N_3300,N_3000);
and U4928 (N_4928,N_3674,N_3620);
nand U4929 (N_4929,N_3877,N_3020);
nor U4930 (N_4930,N_3211,N_3922);
or U4931 (N_4931,N_3997,N_3408);
and U4932 (N_4932,N_3387,N_3627);
nor U4933 (N_4933,N_3357,N_3879);
nand U4934 (N_4934,N_3464,N_3584);
xnor U4935 (N_4935,N_3851,N_3694);
nor U4936 (N_4936,N_3757,N_3331);
nand U4937 (N_4937,N_3357,N_3297);
xor U4938 (N_4938,N_3422,N_3255);
and U4939 (N_4939,N_3390,N_3453);
nand U4940 (N_4940,N_3090,N_3336);
or U4941 (N_4941,N_3830,N_3631);
and U4942 (N_4942,N_3539,N_3960);
and U4943 (N_4943,N_3551,N_3504);
nand U4944 (N_4944,N_3621,N_3519);
nand U4945 (N_4945,N_3485,N_3142);
nor U4946 (N_4946,N_3354,N_3514);
nor U4947 (N_4947,N_3217,N_3510);
and U4948 (N_4948,N_3210,N_3995);
nand U4949 (N_4949,N_3086,N_3804);
and U4950 (N_4950,N_3434,N_3939);
xnor U4951 (N_4951,N_3996,N_3651);
or U4952 (N_4952,N_3489,N_3853);
and U4953 (N_4953,N_3073,N_3576);
or U4954 (N_4954,N_3876,N_3304);
or U4955 (N_4955,N_3926,N_3135);
nor U4956 (N_4956,N_3581,N_3378);
and U4957 (N_4957,N_3614,N_3150);
nor U4958 (N_4958,N_3868,N_3196);
or U4959 (N_4959,N_3241,N_3928);
nand U4960 (N_4960,N_3717,N_3564);
xor U4961 (N_4961,N_3285,N_3981);
nor U4962 (N_4962,N_3173,N_3275);
or U4963 (N_4963,N_3284,N_3697);
or U4964 (N_4964,N_3124,N_3543);
and U4965 (N_4965,N_3584,N_3300);
and U4966 (N_4966,N_3904,N_3084);
and U4967 (N_4967,N_3641,N_3736);
nand U4968 (N_4968,N_3263,N_3480);
nor U4969 (N_4969,N_3662,N_3016);
nor U4970 (N_4970,N_3258,N_3148);
nor U4971 (N_4971,N_3082,N_3671);
and U4972 (N_4972,N_3847,N_3787);
nand U4973 (N_4973,N_3129,N_3002);
and U4974 (N_4974,N_3885,N_3619);
xor U4975 (N_4975,N_3586,N_3724);
nor U4976 (N_4976,N_3194,N_3777);
nor U4977 (N_4977,N_3006,N_3525);
nor U4978 (N_4978,N_3508,N_3108);
and U4979 (N_4979,N_3120,N_3726);
and U4980 (N_4980,N_3539,N_3668);
and U4981 (N_4981,N_3239,N_3623);
or U4982 (N_4982,N_3809,N_3790);
or U4983 (N_4983,N_3422,N_3946);
or U4984 (N_4984,N_3749,N_3960);
xor U4985 (N_4985,N_3012,N_3689);
xor U4986 (N_4986,N_3149,N_3526);
and U4987 (N_4987,N_3765,N_3222);
and U4988 (N_4988,N_3075,N_3261);
nor U4989 (N_4989,N_3666,N_3037);
nor U4990 (N_4990,N_3582,N_3722);
nor U4991 (N_4991,N_3213,N_3420);
and U4992 (N_4992,N_3853,N_3539);
and U4993 (N_4993,N_3080,N_3585);
or U4994 (N_4994,N_3063,N_3155);
or U4995 (N_4995,N_3704,N_3487);
xnor U4996 (N_4996,N_3757,N_3136);
or U4997 (N_4997,N_3989,N_3215);
nand U4998 (N_4998,N_3927,N_3004);
or U4999 (N_4999,N_3049,N_3762);
xnor U5000 (N_5000,N_4488,N_4187);
xnor U5001 (N_5001,N_4875,N_4950);
or U5002 (N_5002,N_4991,N_4393);
xor U5003 (N_5003,N_4509,N_4433);
or U5004 (N_5004,N_4873,N_4556);
xnor U5005 (N_5005,N_4767,N_4124);
xnor U5006 (N_5006,N_4659,N_4044);
and U5007 (N_5007,N_4651,N_4982);
xor U5008 (N_5008,N_4614,N_4653);
nand U5009 (N_5009,N_4386,N_4769);
and U5010 (N_5010,N_4588,N_4785);
nand U5011 (N_5011,N_4698,N_4327);
and U5012 (N_5012,N_4405,N_4694);
or U5013 (N_5013,N_4377,N_4086);
or U5014 (N_5014,N_4012,N_4530);
and U5015 (N_5015,N_4236,N_4722);
and U5016 (N_5016,N_4597,N_4103);
xor U5017 (N_5017,N_4691,N_4397);
xor U5018 (N_5018,N_4312,N_4791);
or U5019 (N_5019,N_4316,N_4714);
or U5020 (N_5020,N_4663,N_4543);
and U5021 (N_5021,N_4381,N_4454);
nor U5022 (N_5022,N_4265,N_4972);
xor U5023 (N_5023,N_4775,N_4523);
xor U5024 (N_5024,N_4915,N_4190);
xor U5025 (N_5025,N_4286,N_4737);
nor U5026 (N_5026,N_4962,N_4887);
nand U5027 (N_5027,N_4413,N_4084);
nor U5028 (N_5028,N_4717,N_4021);
and U5029 (N_5029,N_4980,N_4612);
xnor U5030 (N_5030,N_4109,N_4290);
and U5031 (N_5031,N_4102,N_4716);
nor U5032 (N_5032,N_4045,N_4798);
or U5033 (N_5033,N_4673,N_4149);
and U5034 (N_5034,N_4215,N_4827);
nor U5035 (N_5035,N_4213,N_4648);
nor U5036 (N_5036,N_4844,N_4173);
or U5037 (N_5037,N_4028,N_4170);
and U5038 (N_5038,N_4831,N_4943);
or U5039 (N_5039,N_4174,N_4457);
nand U5040 (N_5040,N_4501,N_4819);
and U5041 (N_5041,N_4595,N_4340);
nand U5042 (N_5042,N_4579,N_4230);
nand U5043 (N_5043,N_4184,N_4476);
nor U5044 (N_5044,N_4701,N_4626);
nand U5045 (N_5045,N_4249,N_4994);
or U5046 (N_5046,N_4687,N_4304);
or U5047 (N_5047,N_4814,N_4233);
or U5048 (N_5048,N_4458,N_4771);
nor U5049 (N_5049,N_4997,N_4738);
nor U5050 (N_5050,N_4764,N_4262);
nand U5051 (N_5051,N_4970,N_4404);
nand U5052 (N_5052,N_4058,N_4126);
or U5053 (N_5053,N_4641,N_4605);
and U5054 (N_5054,N_4890,N_4931);
or U5055 (N_5055,N_4212,N_4253);
nand U5056 (N_5056,N_4960,N_4346);
and U5057 (N_5057,N_4546,N_4709);
nand U5058 (N_5058,N_4739,N_4319);
nand U5059 (N_5059,N_4450,N_4995);
or U5060 (N_5060,N_4732,N_4895);
and U5061 (N_5061,N_4809,N_4857);
xor U5062 (N_5062,N_4024,N_4150);
nand U5063 (N_5063,N_4447,N_4942);
or U5064 (N_5064,N_4622,N_4901);
xnor U5065 (N_5065,N_4254,N_4479);
nand U5066 (N_5066,N_4400,N_4919);
nand U5067 (N_5067,N_4348,N_4521);
or U5068 (N_5068,N_4088,N_4842);
or U5069 (N_5069,N_4807,N_4802);
nand U5070 (N_5070,N_4051,N_4421);
nor U5071 (N_5071,N_4604,N_4146);
or U5072 (N_5072,N_4870,N_4792);
xor U5073 (N_5073,N_4006,N_4141);
xor U5074 (N_5074,N_4815,N_4677);
xor U5075 (N_5075,N_4925,N_4990);
xor U5076 (N_5076,N_4520,N_4825);
nand U5077 (N_5077,N_4060,N_4718);
or U5078 (N_5078,N_4214,N_4891);
nor U5079 (N_5079,N_4562,N_4328);
nand U5080 (N_5080,N_4795,N_4255);
nor U5081 (N_5081,N_4531,N_4706);
xnor U5082 (N_5082,N_4625,N_4632);
xnor U5083 (N_5083,N_4369,N_4448);
nor U5084 (N_5084,N_4325,N_4363);
and U5085 (N_5085,N_4042,N_4329);
nor U5086 (N_5086,N_4489,N_4953);
xnor U5087 (N_5087,N_4854,N_4693);
nand U5088 (N_5088,N_4884,N_4968);
and U5089 (N_5089,N_4243,N_4818);
xor U5090 (N_5090,N_4583,N_4205);
or U5091 (N_5091,N_4470,N_4689);
or U5092 (N_5092,N_4049,N_4550);
or U5093 (N_5093,N_4118,N_4617);
nand U5094 (N_5094,N_4406,N_4935);
xnor U5095 (N_5095,N_4005,N_4337);
nor U5096 (N_5096,N_4451,N_4323);
nor U5097 (N_5097,N_4292,N_4181);
or U5098 (N_5098,N_4441,N_4987);
nor U5099 (N_5099,N_4655,N_4993);
or U5100 (N_5100,N_4267,N_4957);
nand U5101 (N_5101,N_4046,N_4453);
nand U5102 (N_5102,N_4565,N_4074);
and U5103 (N_5103,N_4621,N_4749);
nor U5104 (N_5104,N_4429,N_4535);
and U5105 (N_5105,N_4491,N_4756);
nand U5106 (N_5106,N_4395,N_4881);
nor U5107 (N_5107,N_4114,N_4244);
xor U5108 (N_5108,N_4061,N_4786);
or U5109 (N_5109,N_4022,N_4513);
xor U5110 (N_5110,N_4789,N_4507);
and U5111 (N_5111,N_4894,N_4171);
or U5112 (N_5112,N_4198,N_4680);
xor U5113 (N_5113,N_4161,N_4865);
and U5114 (N_5114,N_4311,N_4667);
xor U5115 (N_5115,N_4030,N_4742);
nand U5116 (N_5116,N_4889,N_4226);
or U5117 (N_5117,N_4496,N_4007);
and U5118 (N_5118,N_4428,N_4148);
and U5119 (N_5119,N_4768,N_4934);
nor U5120 (N_5120,N_4868,N_4760);
and U5121 (N_5121,N_4390,N_4182);
xnor U5122 (N_5122,N_4281,N_4425);
or U5123 (N_5123,N_4782,N_4284);
xnor U5124 (N_5124,N_4611,N_4917);
xnor U5125 (N_5125,N_4526,N_4211);
xnor U5126 (N_5126,N_4493,N_4142);
and U5127 (N_5127,N_4926,N_4983);
or U5128 (N_5128,N_4057,N_4553);
nor U5129 (N_5129,N_4362,N_4300);
nand U5130 (N_5130,N_4947,N_4902);
or U5131 (N_5131,N_4452,N_4027);
or U5132 (N_5132,N_4371,N_4330);
and U5133 (N_5133,N_4954,N_4751);
nand U5134 (N_5134,N_4370,N_4838);
and U5135 (N_5135,N_4153,N_4978);
nor U5136 (N_5136,N_4952,N_4757);
or U5137 (N_5137,N_4351,N_4098);
and U5138 (N_5138,N_4018,N_4541);
and U5139 (N_5139,N_4590,N_4237);
xnor U5140 (N_5140,N_4026,N_4420);
nand U5141 (N_5141,N_4229,N_4684);
and U5142 (N_5142,N_4055,N_4582);
nor U5143 (N_5143,N_4218,N_4289);
nand U5144 (N_5144,N_4068,N_4811);
or U5145 (N_5145,N_4678,N_4867);
xor U5146 (N_5146,N_4922,N_4665);
nand U5147 (N_5147,N_4241,N_4201);
xnor U5148 (N_5148,N_4398,N_4710);
nand U5149 (N_5149,N_4038,N_4577);
nor U5150 (N_5150,N_4116,N_4227);
nand U5151 (N_5151,N_4828,N_4469);
nor U5152 (N_5152,N_4610,N_4314);
nor U5153 (N_5153,N_4485,N_4361);
or U5154 (N_5154,N_4216,N_4713);
nor U5155 (N_5155,N_4298,N_4010);
xnor U5156 (N_5156,N_4586,N_4246);
xnor U5157 (N_5157,N_4047,N_4918);
or U5158 (N_5158,N_4293,N_4686);
xnor U5159 (N_5159,N_4778,N_4260);
nand U5160 (N_5160,N_4969,N_4996);
nand U5161 (N_5161,N_4475,N_4193);
nor U5162 (N_5162,N_4637,N_4195);
nor U5163 (N_5163,N_4747,N_4367);
nand U5164 (N_5164,N_4821,N_4856);
nand U5165 (N_5165,N_4859,N_4512);
nand U5166 (N_5166,N_4675,N_4559);
nor U5167 (N_5167,N_4963,N_4017);
nand U5168 (N_5168,N_4067,N_4909);
xor U5169 (N_5169,N_4107,N_4138);
nand U5170 (N_5170,N_4113,N_4248);
or U5171 (N_5171,N_4683,N_4981);
nand U5172 (N_5172,N_4380,N_4221);
and U5173 (N_5173,N_4008,N_4157);
or U5174 (N_5174,N_4692,N_4951);
or U5175 (N_5175,N_4341,N_4851);
xnor U5176 (N_5176,N_4662,N_4128);
nor U5177 (N_5177,N_4412,N_4774);
or U5178 (N_5178,N_4359,N_4204);
nor U5179 (N_5179,N_4777,N_4445);
xor U5180 (N_5180,N_4162,N_4494);
xor U5181 (N_5181,N_4104,N_4900);
nor U5182 (N_5182,N_4191,N_4973);
or U5183 (N_5183,N_4115,N_4711);
and U5184 (N_5184,N_4755,N_4168);
and U5185 (N_5185,N_4269,N_4893);
nand U5186 (N_5186,N_4898,N_4331);
or U5187 (N_5187,N_4139,N_4882);
or U5188 (N_5188,N_4580,N_4636);
or U5189 (N_5189,N_4735,N_4374);
nand U5190 (N_5190,N_4100,N_4869);
or U5191 (N_5191,N_4514,N_4548);
nand U5192 (N_5192,N_4779,N_4944);
and U5193 (N_5193,N_4129,N_4423);
xor U5194 (N_5194,N_4570,N_4242);
nor U5195 (N_5195,N_4091,N_4619);
nor U5196 (N_5196,N_4877,N_4728);
nor U5197 (N_5197,N_4384,N_4599);
nor U5198 (N_5198,N_4321,N_4896);
xor U5199 (N_5199,N_4183,N_4816);
or U5200 (N_5200,N_4752,N_4634);
nand U5201 (N_5201,N_4538,N_4880);
nor U5202 (N_5202,N_4121,N_4671);
xnor U5203 (N_5203,N_4720,N_4180);
nor U5204 (N_5204,N_4130,N_4569);
xnor U5205 (N_5205,N_4812,N_4704);
and U5206 (N_5206,N_4135,N_4471);
nor U5207 (N_5207,N_4210,N_4840);
or U5208 (N_5208,N_4466,N_4350);
xor U5209 (N_5209,N_4552,N_4878);
and U5210 (N_5210,N_4486,N_4324);
and U5211 (N_5211,N_4930,N_4519);
nand U5212 (N_5212,N_4871,N_4432);
nand U5213 (N_5213,N_4207,N_4291);
xnor U5214 (N_5214,N_4202,N_4349);
nand U5215 (N_5215,N_4772,N_4864);
nor U5216 (N_5216,N_4169,N_4905);
nand U5217 (N_5217,N_4417,N_4401);
xor U5218 (N_5218,N_4387,N_4615);
nor U5219 (N_5219,N_4136,N_4696);
xnor U5220 (N_5220,N_4506,N_4295);
and U5221 (N_5221,N_4726,N_4016);
nor U5222 (N_5222,N_4724,N_4499);
nand U5223 (N_5223,N_4702,N_4598);
nor U5224 (N_5224,N_4373,N_4998);
or U5225 (N_5225,N_4770,N_4776);
and U5226 (N_5226,N_4533,N_4504);
and U5227 (N_5227,N_4613,N_4487);
or U5228 (N_5228,N_4426,N_4092);
or U5229 (N_5229,N_4578,N_4761);
xnor U5230 (N_5230,N_4872,N_4585);
nand U5231 (N_5231,N_4906,N_4977);
xnor U5232 (N_5232,N_4054,N_4143);
nand U5233 (N_5233,N_4003,N_4568);
or U5234 (N_5234,N_4836,N_4245);
and U5235 (N_5235,N_4946,N_4522);
xnor U5236 (N_5236,N_4638,N_4172);
and U5237 (N_5237,N_4200,N_4062);
or U5238 (N_5238,N_4594,N_4736);
xor U5239 (N_5239,N_4383,N_4674);
or U5240 (N_5240,N_4431,N_4516);
and U5241 (N_5241,N_4070,N_4083);
nor U5242 (N_5242,N_4366,N_4072);
and U5243 (N_5243,N_4797,N_4343);
or U5244 (N_5244,N_4788,N_4729);
xor U5245 (N_5245,N_4961,N_4924);
and U5246 (N_5246,N_4414,N_4832);
or U5247 (N_5247,N_4988,N_4861);
nand U5248 (N_5248,N_4719,N_4572);
nand U5249 (N_5249,N_4700,N_4823);
xor U5250 (N_5250,N_4059,N_4261);
and U5251 (N_5251,N_4631,N_4784);
xor U5252 (N_5252,N_4551,N_4270);
nand U5253 (N_5253,N_4307,N_4616);
or U5254 (N_5254,N_4656,N_4320);
nand U5255 (N_5255,N_4829,N_4589);
nor U5256 (N_5256,N_4031,N_4940);
nor U5257 (N_5257,N_4892,N_4155);
xor U5258 (N_5258,N_4029,N_4679);
and U5259 (N_5259,N_4463,N_4664);
xnor U5260 (N_5260,N_4257,N_4309);
nor U5261 (N_5261,N_4273,N_4399);
nand U5262 (N_5262,N_4365,N_4294);
or U5263 (N_5263,N_4939,N_4620);
nand U5264 (N_5264,N_4301,N_4633);
or U5265 (N_5265,N_4490,N_4484);
nor U5266 (N_5266,N_4108,N_4862);
nand U5267 (N_5267,N_4534,N_4544);
nand U5268 (N_5268,N_4219,N_4547);
nand U5269 (N_5269,N_4110,N_4075);
and U5270 (N_5270,N_4697,N_4503);
xnor U5271 (N_5271,N_4804,N_4574);
xnor U5272 (N_5272,N_4385,N_4699);
and U5273 (N_5273,N_4502,N_4002);
nand U5274 (N_5274,N_4670,N_4666);
xnor U5275 (N_5275,N_4333,N_4746);
xor U5276 (N_5276,N_4179,N_4833);
or U5277 (N_5277,N_4754,N_4885);
and U5278 (N_5278,N_4646,N_4630);
xnor U5279 (N_5279,N_4907,N_4354);
xnor U5280 (N_5280,N_4936,N_4927);
xor U5281 (N_5281,N_4079,N_4278);
nor U5282 (N_5282,N_4941,N_4635);
or U5283 (N_5283,N_4763,N_4837);
nor U5284 (N_5284,N_4147,N_4629);
and U5285 (N_5285,N_4609,N_4053);
xor U5286 (N_5286,N_4876,N_4056);
xor U5287 (N_5287,N_4932,N_4418);
or U5288 (N_5288,N_4965,N_4288);
xnor U5289 (N_5289,N_4071,N_4658);
or U5290 (N_5290,N_4623,N_4217);
nor U5291 (N_5291,N_4145,N_4753);
nor U5292 (N_5292,N_4481,N_4920);
or U5293 (N_5293,N_4912,N_4654);
or U5294 (N_5294,N_4587,N_4101);
nor U5295 (N_5295,N_4120,N_4593);
nor U5296 (N_5296,N_4571,N_4855);
nor U5297 (N_5297,N_4524,N_4731);
nand U5298 (N_5298,N_4185,N_4140);
and U5299 (N_5299,N_4899,N_4783);
and U5300 (N_5300,N_4251,N_4093);
and U5301 (N_5301,N_4438,N_4596);
nand U5302 (N_5302,N_4967,N_4483);
nor U5303 (N_5303,N_4879,N_4652);
and U5304 (N_5304,N_4618,N_4403);
and U5305 (N_5305,N_4178,N_4705);
xor U5306 (N_5306,N_4497,N_4549);
or U5307 (N_5307,N_4883,N_4188);
and U5308 (N_5308,N_4322,N_4052);
or U5309 (N_5309,N_4601,N_4517);
nand U5310 (N_5310,N_4449,N_4886);
or U5311 (N_5311,N_4745,N_4020);
nor U5312 (N_5312,N_4040,N_4105);
and U5313 (N_5313,N_4703,N_4539);
and U5314 (N_5314,N_4592,N_4511);
and U5315 (N_5315,N_4561,N_4081);
nor U5316 (N_5316,N_4437,N_4986);
nor U5317 (N_5317,N_4069,N_4087);
xor U5318 (N_5318,N_4411,N_4163);
nand U5319 (N_5319,N_4527,N_4858);
nor U5320 (N_5320,N_4681,N_4462);
and U5321 (N_5321,N_4695,N_4310);
nor U5322 (N_5322,N_4813,N_4649);
nor U5323 (N_5323,N_4131,N_4167);
and U5324 (N_5324,N_4106,N_4296);
or U5325 (N_5325,N_4368,N_4308);
and U5326 (N_5326,N_4014,N_4566);
xnor U5327 (N_5327,N_4076,N_4228);
or U5328 (N_5328,N_4099,N_4644);
nor U5329 (N_5329,N_4382,N_4558);
xor U5330 (N_5330,N_4043,N_4657);
or U5331 (N_5331,N_4004,N_4743);
nand U5332 (N_5332,N_4806,N_4165);
nand U5333 (N_5333,N_4971,N_4306);
nand U5334 (N_5334,N_4419,N_4647);
nor U5335 (N_5335,N_4672,N_4639);
or U5336 (N_5336,N_4339,N_4326);
xor U5337 (N_5337,N_4235,N_4035);
xor U5338 (N_5338,N_4525,N_4472);
or U5339 (N_5339,N_4766,N_4555);
xor U5340 (N_5340,N_4468,N_4707);
nand U5341 (N_5341,N_4794,N_4208);
nand U5342 (N_5342,N_4446,N_4958);
nor U5343 (N_5343,N_4643,N_4863);
xnor U5344 (N_5344,N_4209,N_4280);
nand U5345 (N_5345,N_4063,N_4271);
nor U5346 (N_5346,N_4356,N_4335);
xnor U5347 (N_5347,N_4834,N_4465);
nor U5348 (N_5348,N_4025,N_4282);
or U5349 (N_5349,N_4317,N_4408);
and U5350 (N_5350,N_4125,N_4608);
xnor U5351 (N_5351,N_4781,N_4250);
xnor U5352 (N_5352,N_4495,N_4276);
nor U5353 (N_5353,N_4966,N_4758);
and U5354 (N_5354,N_4305,N_4467);
and U5355 (N_5355,N_4564,N_4554);
and U5356 (N_5356,N_4508,N_4256);
nand U5357 (N_5357,N_4800,N_4796);
nand U5358 (N_5358,N_4482,N_4725);
xor U5359 (N_5359,N_4841,N_4232);
xor U5360 (N_5360,N_4492,N_4443);
nor U5361 (N_5361,N_4283,N_4206);
and U5362 (N_5362,N_4773,N_4041);
nand U5363 (N_5363,N_4956,N_4357);
nor U5364 (N_5364,N_4843,N_4921);
or U5365 (N_5365,N_4334,N_4203);
and U5366 (N_5366,N_4336,N_4032);
xor U5367 (N_5367,N_4094,N_4225);
nor U5368 (N_5368,N_4189,N_4734);
and U5369 (N_5369,N_4668,N_4847);
nand U5370 (N_5370,N_4799,N_4455);
nand U5371 (N_5371,N_4231,N_4762);
or U5372 (N_5372,N_4669,N_4741);
nor U5373 (N_5373,N_4015,N_4790);
and U5374 (N_5374,N_4624,N_4793);
and U5375 (N_5375,N_4442,N_4576);
xor U5376 (N_5376,N_4272,N_4019);
and U5377 (N_5377,N_4133,N_4801);
and U5378 (N_5378,N_4388,N_4464);
or U5379 (N_5379,N_4440,N_4478);
and U5380 (N_5380,N_4730,N_4817);
or U5381 (N_5381,N_4345,N_4159);
and U5382 (N_5382,N_4302,N_4975);
and U5383 (N_5383,N_4050,N_4456);
nand U5384 (N_5384,N_4748,N_4913);
nand U5385 (N_5385,N_4410,N_4089);
and U5386 (N_5386,N_4460,N_4222);
nor U5387 (N_5387,N_4480,N_4224);
and U5388 (N_5388,N_4938,N_4712);
xnor U5389 (N_5389,N_4567,N_4259);
and U5390 (N_5390,N_4937,N_4378);
nand U5391 (N_5391,N_4389,N_4536);
and U5392 (N_5392,N_4355,N_4112);
nand U5393 (N_5393,N_4923,N_4929);
and U5394 (N_5394,N_4822,N_4557);
xnor U5395 (N_5395,N_4911,N_4708);
xnor U5396 (N_5396,N_4853,N_4117);
or U5397 (N_5397,N_4846,N_4082);
or U5398 (N_5398,N_4177,N_4948);
xnor U5399 (N_5399,N_4860,N_4258);
nand U5400 (N_5400,N_4036,N_4034);
or U5401 (N_5401,N_4344,N_4949);
and U5402 (N_5402,N_4979,N_4436);
and U5403 (N_5403,N_4164,N_4928);
and U5404 (N_5404,N_4009,N_4315);
nand U5405 (N_5405,N_4394,N_4127);
nor U5406 (N_5406,N_4223,N_4850);
nor U5407 (N_5407,N_4715,N_4744);
and U5408 (N_5408,N_4396,N_4435);
nand U5409 (N_5409,N_4360,N_4154);
xor U5410 (N_5410,N_4676,N_4933);
xnor U5411 (N_5411,N_4826,N_4379);
xor U5412 (N_5412,N_4376,N_4285);
and U5413 (N_5413,N_4064,N_4976);
nor U5414 (N_5414,N_4439,N_4560);
nor U5415 (N_5415,N_4252,N_4808);
nor U5416 (N_5416,N_4097,N_4266);
and U5417 (N_5417,N_4358,N_4810);
nand U5418 (N_5418,N_4196,N_4033);
nor U5419 (N_5419,N_4277,N_4835);
xnor U5420 (N_5420,N_4852,N_4914);
and U5421 (N_5421,N_4537,N_4607);
and U5422 (N_5422,N_4575,N_4156);
nor U5423 (N_5423,N_4830,N_4584);
xnor U5424 (N_5424,N_4364,N_4955);
nor U5425 (N_5425,N_4845,N_4078);
or U5426 (N_5426,N_4721,N_4959);
xnor U5427 (N_5427,N_4085,N_4152);
nor U5428 (N_5428,N_4532,N_4001);
xor U5429 (N_5429,N_4077,N_4650);
and U5430 (N_5430,N_4573,N_4529);
xor U5431 (N_5431,N_4600,N_4240);
or U5432 (N_5432,N_4916,N_4318);
nor U5433 (N_5433,N_4264,N_4848);
nor U5434 (N_5434,N_4194,N_4591);
xor U5435 (N_5435,N_4897,N_4151);
xnor U5436 (N_5436,N_4459,N_4352);
and U5437 (N_5437,N_4945,N_4545);
and U5438 (N_5438,N_4199,N_4908);
nand U5439 (N_5439,N_4080,N_4498);
nor U5440 (N_5440,N_4013,N_4910);
xor U5441 (N_5441,N_4332,N_4175);
and U5442 (N_5442,N_4984,N_4992);
nand U5443 (N_5443,N_4096,N_4186);
and U5444 (N_5444,N_4268,N_4473);
and U5445 (N_5445,N_4904,N_4065);
xnor U5446 (N_5446,N_4299,N_4238);
xnor U5447 (N_5447,N_4528,N_4303);
nor U5448 (N_5448,N_4628,N_4444);
xor U5449 (N_5449,N_4477,N_4690);
nand U5450 (N_5450,N_4424,N_4111);
or U5451 (N_5451,N_4158,N_4903);
xor U5452 (N_5452,N_4999,N_4874);
nand U5453 (N_5453,N_4342,N_4392);
nand U5454 (N_5454,N_4759,N_4176);
xnor U5455 (N_5455,N_4500,N_4780);
xnor U5456 (N_5456,N_4123,N_4606);
xor U5457 (N_5457,N_4740,N_4402);
nand U5458 (N_5458,N_4274,N_4220);
and U5459 (N_5459,N_4372,N_4137);
or U5460 (N_5460,N_4338,N_4765);
nand U5461 (N_5461,N_4542,N_4685);
nor U5462 (N_5462,N_4430,N_4563);
nand U5463 (N_5463,N_4416,N_4640);
nand U5464 (N_5464,N_4688,N_4422);
nor U5465 (N_5465,N_4239,N_4048);
nor U5466 (N_5466,N_4391,N_4824);
nor U5467 (N_5467,N_4134,N_4297);
xnor U5468 (N_5468,N_4166,N_4000);
nor U5469 (N_5469,N_4434,N_4642);
xnor U5470 (N_5470,N_4660,N_4505);
nand U5471 (N_5471,N_4353,N_4011);
nand U5472 (N_5472,N_4275,N_4805);
or U5473 (N_5473,N_4247,N_4461);
and U5474 (N_5474,N_4375,N_4347);
and U5475 (N_5475,N_4515,N_4023);
and U5476 (N_5476,N_4839,N_4985);
xor U5477 (N_5477,N_4095,N_4733);
or U5478 (N_5478,N_4510,N_4723);
and U5479 (N_5479,N_4066,N_4313);
nand U5480 (N_5480,N_4627,N_4581);
or U5481 (N_5481,N_4803,N_4849);
or U5482 (N_5482,N_4866,N_4540);
and U5483 (N_5483,N_4263,N_4727);
nor U5484 (N_5484,N_4192,N_4160);
xor U5485 (N_5485,N_4073,N_4645);
and U5486 (N_5486,N_4132,N_4415);
nor U5487 (N_5487,N_4603,N_4197);
xnor U5488 (N_5488,N_4820,N_4122);
xnor U5489 (N_5489,N_4037,N_4279);
nand U5490 (N_5490,N_4888,N_4750);
xnor U5491 (N_5491,N_4144,N_4682);
xor U5492 (N_5492,N_4602,N_4518);
or U5493 (N_5493,N_4661,N_4989);
or U5494 (N_5494,N_4787,N_4234);
xor U5495 (N_5495,N_4287,N_4090);
nor U5496 (N_5496,N_4119,N_4427);
nand U5497 (N_5497,N_4964,N_4474);
nand U5498 (N_5498,N_4407,N_4409);
xnor U5499 (N_5499,N_4974,N_4039);
xor U5500 (N_5500,N_4279,N_4934);
or U5501 (N_5501,N_4052,N_4885);
or U5502 (N_5502,N_4103,N_4509);
and U5503 (N_5503,N_4683,N_4983);
nand U5504 (N_5504,N_4168,N_4022);
nor U5505 (N_5505,N_4400,N_4527);
and U5506 (N_5506,N_4749,N_4747);
xor U5507 (N_5507,N_4968,N_4457);
and U5508 (N_5508,N_4877,N_4787);
nor U5509 (N_5509,N_4276,N_4552);
and U5510 (N_5510,N_4857,N_4549);
and U5511 (N_5511,N_4562,N_4994);
or U5512 (N_5512,N_4480,N_4261);
nor U5513 (N_5513,N_4803,N_4086);
nor U5514 (N_5514,N_4439,N_4964);
xor U5515 (N_5515,N_4232,N_4696);
and U5516 (N_5516,N_4304,N_4568);
nor U5517 (N_5517,N_4416,N_4556);
or U5518 (N_5518,N_4937,N_4873);
or U5519 (N_5519,N_4153,N_4602);
or U5520 (N_5520,N_4934,N_4840);
xnor U5521 (N_5521,N_4229,N_4040);
xor U5522 (N_5522,N_4272,N_4509);
and U5523 (N_5523,N_4343,N_4556);
and U5524 (N_5524,N_4933,N_4480);
and U5525 (N_5525,N_4354,N_4958);
and U5526 (N_5526,N_4127,N_4980);
nand U5527 (N_5527,N_4562,N_4085);
nor U5528 (N_5528,N_4352,N_4665);
or U5529 (N_5529,N_4577,N_4133);
or U5530 (N_5530,N_4600,N_4862);
nand U5531 (N_5531,N_4223,N_4598);
and U5532 (N_5532,N_4257,N_4505);
and U5533 (N_5533,N_4796,N_4194);
xor U5534 (N_5534,N_4141,N_4926);
or U5535 (N_5535,N_4756,N_4680);
and U5536 (N_5536,N_4677,N_4133);
nor U5537 (N_5537,N_4735,N_4627);
or U5538 (N_5538,N_4239,N_4117);
xor U5539 (N_5539,N_4871,N_4087);
nand U5540 (N_5540,N_4391,N_4791);
and U5541 (N_5541,N_4944,N_4071);
nand U5542 (N_5542,N_4251,N_4162);
or U5543 (N_5543,N_4949,N_4325);
or U5544 (N_5544,N_4166,N_4765);
and U5545 (N_5545,N_4750,N_4765);
nor U5546 (N_5546,N_4165,N_4737);
nand U5547 (N_5547,N_4633,N_4574);
nor U5548 (N_5548,N_4380,N_4461);
or U5549 (N_5549,N_4134,N_4950);
and U5550 (N_5550,N_4569,N_4456);
xor U5551 (N_5551,N_4728,N_4209);
xor U5552 (N_5552,N_4501,N_4944);
and U5553 (N_5553,N_4421,N_4950);
nand U5554 (N_5554,N_4582,N_4353);
nor U5555 (N_5555,N_4465,N_4001);
nor U5556 (N_5556,N_4975,N_4115);
or U5557 (N_5557,N_4950,N_4982);
or U5558 (N_5558,N_4290,N_4258);
nor U5559 (N_5559,N_4115,N_4022);
or U5560 (N_5560,N_4215,N_4423);
nor U5561 (N_5561,N_4724,N_4043);
xnor U5562 (N_5562,N_4102,N_4235);
nor U5563 (N_5563,N_4511,N_4876);
nor U5564 (N_5564,N_4337,N_4388);
nor U5565 (N_5565,N_4315,N_4067);
nor U5566 (N_5566,N_4196,N_4057);
or U5567 (N_5567,N_4966,N_4525);
xor U5568 (N_5568,N_4940,N_4990);
and U5569 (N_5569,N_4695,N_4940);
and U5570 (N_5570,N_4961,N_4043);
xnor U5571 (N_5571,N_4220,N_4880);
nand U5572 (N_5572,N_4650,N_4806);
nor U5573 (N_5573,N_4874,N_4566);
nand U5574 (N_5574,N_4478,N_4776);
xnor U5575 (N_5575,N_4037,N_4677);
nor U5576 (N_5576,N_4589,N_4010);
nand U5577 (N_5577,N_4256,N_4574);
nand U5578 (N_5578,N_4242,N_4351);
nor U5579 (N_5579,N_4581,N_4036);
nand U5580 (N_5580,N_4432,N_4332);
nor U5581 (N_5581,N_4918,N_4113);
nand U5582 (N_5582,N_4945,N_4671);
and U5583 (N_5583,N_4528,N_4339);
or U5584 (N_5584,N_4645,N_4890);
and U5585 (N_5585,N_4892,N_4420);
or U5586 (N_5586,N_4084,N_4365);
and U5587 (N_5587,N_4815,N_4838);
nand U5588 (N_5588,N_4378,N_4992);
nor U5589 (N_5589,N_4950,N_4888);
and U5590 (N_5590,N_4481,N_4317);
nor U5591 (N_5591,N_4111,N_4245);
or U5592 (N_5592,N_4885,N_4372);
xor U5593 (N_5593,N_4141,N_4102);
and U5594 (N_5594,N_4335,N_4498);
nand U5595 (N_5595,N_4305,N_4237);
xor U5596 (N_5596,N_4055,N_4410);
xor U5597 (N_5597,N_4190,N_4410);
or U5598 (N_5598,N_4311,N_4851);
xnor U5599 (N_5599,N_4795,N_4774);
or U5600 (N_5600,N_4565,N_4398);
nor U5601 (N_5601,N_4240,N_4026);
nor U5602 (N_5602,N_4520,N_4104);
nor U5603 (N_5603,N_4966,N_4010);
xor U5604 (N_5604,N_4115,N_4672);
xnor U5605 (N_5605,N_4340,N_4279);
xor U5606 (N_5606,N_4897,N_4636);
nor U5607 (N_5607,N_4261,N_4742);
or U5608 (N_5608,N_4299,N_4697);
nor U5609 (N_5609,N_4286,N_4548);
nor U5610 (N_5610,N_4146,N_4245);
nor U5611 (N_5611,N_4136,N_4734);
xor U5612 (N_5612,N_4087,N_4757);
or U5613 (N_5613,N_4558,N_4295);
nand U5614 (N_5614,N_4596,N_4473);
nand U5615 (N_5615,N_4304,N_4966);
and U5616 (N_5616,N_4915,N_4130);
xor U5617 (N_5617,N_4135,N_4474);
xor U5618 (N_5618,N_4923,N_4297);
nand U5619 (N_5619,N_4347,N_4041);
nor U5620 (N_5620,N_4653,N_4924);
nand U5621 (N_5621,N_4142,N_4538);
or U5622 (N_5622,N_4201,N_4221);
nor U5623 (N_5623,N_4712,N_4526);
nor U5624 (N_5624,N_4696,N_4040);
nor U5625 (N_5625,N_4490,N_4730);
nand U5626 (N_5626,N_4061,N_4060);
or U5627 (N_5627,N_4634,N_4612);
nor U5628 (N_5628,N_4649,N_4907);
and U5629 (N_5629,N_4747,N_4075);
nand U5630 (N_5630,N_4803,N_4606);
nor U5631 (N_5631,N_4551,N_4430);
and U5632 (N_5632,N_4407,N_4196);
nor U5633 (N_5633,N_4953,N_4684);
xor U5634 (N_5634,N_4802,N_4147);
nor U5635 (N_5635,N_4327,N_4192);
or U5636 (N_5636,N_4357,N_4477);
nor U5637 (N_5637,N_4829,N_4297);
nand U5638 (N_5638,N_4758,N_4380);
nor U5639 (N_5639,N_4447,N_4553);
nand U5640 (N_5640,N_4598,N_4372);
and U5641 (N_5641,N_4355,N_4857);
nand U5642 (N_5642,N_4095,N_4673);
or U5643 (N_5643,N_4379,N_4509);
nand U5644 (N_5644,N_4367,N_4329);
or U5645 (N_5645,N_4265,N_4608);
or U5646 (N_5646,N_4142,N_4602);
and U5647 (N_5647,N_4926,N_4561);
nand U5648 (N_5648,N_4608,N_4638);
xor U5649 (N_5649,N_4557,N_4399);
nor U5650 (N_5650,N_4076,N_4621);
nor U5651 (N_5651,N_4671,N_4758);
nor U5652 (N_5652,N_4238,N_4134);
nor U5653 (N_5653,N_4841,N_4541);
or U5654 (N_5654,N_4150,N_4059);
or U5655 (N_5655,N_4067,N_4652);
nor U5656 (N_5656,N_4174,N_4644);
nor U5657 (N_5657,N_4725,N_4865);
nand U5658 (N_5658,N_4630,N_4958);
and U5659 (N_5659,N_4473,N_4076);
or U5660 (N_5660,N_4675,N_4363);
or U5661 (N_5661,N_4262,N_4059);
nand U5662 (N_5662,N_4493,N_4876);
xor U5663 (N_5663,N_4689,N_4063);
and U5664 (N_5664,N_4372,N_4382);
nor U5665 (N_5665,N_4177,N_4945);
nor U5666 (N_5666,N_4548,N_4044);
and U5667 (N_5667,N_4887,N_4704);
or U5668 (N_5668,N_4843,N_4599);
and U5669 (N_5669,N_4222,N_4328);
xor U5670 (N_5670,N_4446,N_4047);
nor U5671 (N_5671,N_4237,N_4713);
nand U5672 (N_5672,N_4355,N_4936);
nand U5673 (N_5673,N_4503,N_4997);
xnor U5674 (N_5674,N_4138,N_4682);
nand U5675 (N_5675,N_4564,N_4288);
and U5676 (N_5676,N_4975,N_4267);
xor U5677 (N_5677,N_4171,N_4127);
or U5678 (N_5678,N_4228,N_4582);
nand U5679 (N_5679,N_4748,N_4389);
nor U5680 (N_5680,N_4397,N_4490);
nor U5681 (N_5681,N_4029,N_4807);
and U5682 (N_5682,N_4615,N_4766);
xor U5683 (N_5683,N_4744,N_4257);
xor U5684 (N_5684,N_4632,N_4909);
xor U5685 (N_5685,N_4085,N_4385);
nor U5686 (N_5686,N_4894,N_4167);
and U5687 (N_5687,N_4179,N_4718);
xor U5688 (N_5688,N_4112,N_4229);
or U5689 (N_5689,N_4288,N_4513);
xor U5690 (N_5690,N_4541,N_4078);
xor U5691 (N_5691,N_4700,N_4736);
and U5692 (N_5692,N_4167,N_4250);
xnor U5693 (N_5693,N_4258,N_4701);
and U5694 (N_5694,N_4317,N_4370);
xnor U5695 (N_5695,N_4102,N_4780);
and U5696 (N_5696,N_4595,N_4591);
nor U5697 (N_5697,N_4049,N_4236);
xor U5698 (N_5698,N_4345,N_4198);
nand U5699 (N_5699,N_4089,N_4366);
xnor U5700 (N_5700,N_4769,N_4316);
nor U5701 (N_5701,N_4794,N_4591);
xnor U5702 (N_5702,N_4936,N_4410);
or U5703 (N_5703,N_4214,N_4667);
and U5704 (N_5704,N_4060,N_4163);
and U5705 (N_5705,N_4681,N_4863);
xor U5706 (N_5706,N_4500,N_4687);
nand U5707 (N_5707,N_4570,N_4275);
nand U5708 (N_5708,N_4595,N_4074);
or U5709 (N_5709,N_4147,N_4761);
and U5710 (N_5710,N_4833,N_4903);
xor U5711 (N_5711,N_4546,N_4272);
nor U5712 (N_5712,N_4716,N_4217);
and U5713 (N_5713,N_4611,N_4653);
nand U5714 (N_5714,N_4678,N_4854);
nand U5715 (N_5715,N_4440,N_4670);
and U5716 (N_5716,N_4423,N_4024);
xnor U5717 (N_5717,N_4134,N_4719);
nand U5718 (N_5718,N_4041,N_4786);
nand U5719 (N_5719,N_4138,N_4398);
xnor U5720 (N_5720,N_4309,N_4992);
nand U5721 (N_5721,N_4553,N_4153);
nand U5722 (N_5722,N_4114,N_4805);
and U5723 (N_5723,N_4534,N_4061);
or U5724 (N_5724,N_4835,N_4042);
nor U5725 (N_5725,N_4673,N_4403);
or U5726 (N_5726,N_4959,N_4088);
or U5727 (N_5727,N_4751,N_4393);
or U5728 (N_5728,N_4645,N_4684);
nor U5729 (N_5729,N_4341,N_4308);
and U5730 (N_5730,N_4117,N_4817);
xor U5731 (N_5731,N_4079,N_4252);
and U5732 (N_5732,N_4415,N_4319);
xor U5733 (N_5733,N_4400,N_4939);
and U5734 (N_5734,N_4358,N_4368);
xnor U5735 (N_5735,N_4593,N_4443);
and U5736 (N_5736,N_4577,N_4480);
xor U5737 (N_5737,N_4176,N_4771);
nor U5738 (N_5738,N_4993,N_4839);
and U5739 (N_5739,N_4285,N_4887);
and U5740 (N_5740,N_4249,N_4047);
and U5741 (N_5741,N_4138,N_4523);
or U5742 (N_5742,N_4462,N_4630);
and U5743 (N_5743,N_4710,N_4559);
or U5744 (N_5744,N_4762,N_4064);
and U5745 (N_5745,N_4877,N_4618);
xor U5746 (N_5746,N_4582,N_4985);
or U5747 (N_5747,N_4615,N_4099);
and U5748 (N_5748,N_4101,N_4713);
and U5749 (N_5749,N_4132,N_4830);
nand U5750 (N_5750,N_4110,N_4509);
and U5751 (N_5751,N_4895,N_4005);
xor U5752 (N_5752,N_4655,N_4458);
nor U5753 (N_5753,N_4150,N_4829);
nand U5754 (N_5754,N_4842,N_4668);
and U5755 (N_5755,N_4812,N_4634);
nand U5756 (N_5756,N_4021,N_4096);
nor U5757 (N_5757,N_4581,N_4058);
xor U5758 (N_5758,N_4304,N_4340);
nor U5759 (N_5759,N_4792,N_4743);
or U5760 (N_5760,N_4398,N_4271);
nor U5761 (N_5761,N_4440,N_4604);
nor U5762 (N_5762,N_4020,N_4724);
or U5763 (N_5763,N_4572,N_4677);
and U5764 (N_5764,N_4608,N_4591);
or U5765 (N_5765,N_4126,N_4842);
or U5766 (N_5766,N_4219,N_4763);
nand U5767 (N_5767,N_4554,N_4470);
nand U5768 (N_5768,N_4299,N_4640);
or U5769 (N_5769,N_4563,N_4772);
nor U5770 (N_5770,N_4746,N_4818);
nor U5771 (N_5771,N_4296,N_4038);
xor U5772 (N_5772,N_4219,N_4730);
nor U5773 (N_5773,N_4208,N_4462);
and U5774 (N_5774,N_4442,N_4675);
nor U5775 (N_5775,N_4814,N_4000);
or U5776 (N_5776,N_4325,N_4068);
or U5777 (N_5777,N_4371,N_4127);
nand U5778 (N_5778,N_4629,N_4456);
xor U5779 (N_5779,N_4287,N_4000);
xnor U5780 (N_5780,N_4605,N_4980);
nand U5781 (N_5781,N_4738,N_4953);
and U5782 (N_5782,N_4509,N_4861);
or U5783 (N_5783,N_4693,N_4998);
nand U5784 (N_5784,N_4610,N_4546);
nor U5785 (N_5785,N_4969,N_4966);
and U5786 (N_5786,N_4263,N_4309);
nand U5787 (N_5787,N_4060,N_4964);
and U5788 (N_5788,N_4243,N_4165);
nand U5789 (N_5789,N_4571,N_4939);
and U5790 (N_5790,N_4998,N_4291);
nand U5791 (N_5791,N_4491,N_4121);
nor U5792 (N_5792,N_4736,N_4297);
or U5793 (N_5793,N_4332,N_4850);
xor U5794 (N_5794,N_4457,N_4721);
xnor U5795 (N_5795,N_4695,N_4746);
nor U5796 (N_5796,N_4010,N_4378);
nand U5797 (N_5797,N_4893,N_4588);
or U5798 (N_5798,N_4826,N_4676);
xnor U5799 (N_5799,N_4580,N_4634);
xor U5800 (N_5800,N_4042,N_4103);
nand U5801 (N_5801,N_4605,N_4559);
or U5802 (N_5802,N_4155,N_4813);
and U5803 (N_5803,N_4339,N_4717);
or U5804 (N_5804,N_4306,N_4942);
nor U5805 (N_5805,N_4381,N_4114);
xor U5806 (N_5806,N_4505,N_4781);
or U5807 (N_5807,N_4492,N_4950);
and U5808 (N_5808,N_4612,N_4334);
and U5809 (N_5809,N_4878,N_4387);
and U5810 (N_5810,N_4436,N_4360);
nor U5811 (N_5811,N_4986,N_4633);
and U5812 (N_5812,N_4062,N_4286);
or U5813 (N_5813,N_4080,N_4759);
and U5814 (N_5814,N_4365,N_4523);
nor U5815 (N_5815,N_4843,N_4157);
nor U5816 (N_5816,N_4401,N_4703);
and U5817 (N_5817,N_4258,N_4099);
or U5818 (N_5818,N_4601,N_4161);
xnor U5819 (N_5819,N_4373,N_4621);
nor U5820 (N_5820,N_4435,N_4903);
nand U5821 (N_5821,N_4527,N_4126);
nand U5822 (N_5822,N_4252,N_4953);
or U5823 (N_5823,N_4778,N_4528);
and U5824 (N_5824,N_4928,N_4683);
nor U5825 (N_5825,N_4048,N_4841);
nor U5826 (N_5826,N_4420,N_4141);
xor U5827 (N_5827,N_4164,N_4448);
and U5828 (N_5828,N_4021,N_4564);
nand U5829 (N_5829,N_4821,N_4992);
nor U5830 (N_5830,N_4820,N_4849);
nand U5831 (N_5831,N_4356,N_4610);
xnor U5832 (N_5832,N_4024,N_4178);
or U5833 (N_5833,N_4993,N_4272);
or U5834 (N_5834,N_4820,N_4271);
nand U5835 (N_5835,N_4309,N_4381);
or U5836 (N_5836,N_4557,N_4917);
and U5837 (N_5837,N_4539,N_4813);
and U5838 (N_5838,N_4927,N_4028);
nand U5839 (N_5839,N_4230,N_4884);
xnor U5840 (N_5840,N_4552,N_4311);
and U5841 (N_5841,N_4680,N_4294);
and U5842 (N_5842,N_4607,N_4347);
and U5843 (N_5843,N_4437,N_4895);
nand U5844 (N_5844,N_4279,N_4729);
nor U5845 (N_5845,N_4976,N_4645);
and U5846 (N_5846,N_4481,N_4419);
or U5847 (N_5847,N_4217,N_4870);
xor U5848 (N_5848,N_4696,N_4851);
nor U5849 (N_5849,N_4391,N_4457);
or U5850 (N_5850,N_4157,N_4808);
xor U5851 (N_5851,N_4388,N_4683);
or U5852 (N_5852,N_4762,N_4239);
nand U5853 (N_5853,N_4278,N_4234);
nand U5854 (N_5854,N_4146,N_4984);
or U5855 (N_5855,N_4404,N_4936);
nor U5856 (N_5856,N_4327,N_4380);
nor U5857 (N_5857,N_4857,N_4345);
nand U5858 (N_5858,N_4870,N_4006);
nor U5859 (N_5859,N_4317,N_4166);
nor U5860 (N_5860,N_4370,N_4081);
xnor U5861 (N_5861,N_4916,N_4826);
and U5862 (N_5862,N_4658,N_4179);
nor U5863 (N_5863,N_4122,N_4464);
xnor U5864 (N_5864,N_4691,N_4322);
or U5865 (N_5865,N_4094,N_4744);
and U5866 (N_5866,N_4496,N_4200);
nand U5867 (N_5867,N_4363,N_4017);
and U5868 (N_5868,N_4483,N_4972);
or U5869 (N_5869,N_4543,N_4697);
nand U5870 (N_5870,N_4506,N_4110);
and U5871 (N_5871,N_4210,N_4889);
nor U5872 (N_5872,N_4631,N_4823);
nand U5873 (N_5873,N_4152,N_4284);
and U5874 (N_5874,N_4128,N_4207);
and U5875 (N_5875,N_4969,N_4742);
or U5876 (N_5876,N_4857,N_4620);
or U5877 (N_5877,N_4696,N_4439);
xor U5878 (N_5878,N_4497,N_4537);
nor U5879 (N_5879,N_4946,N_4620);
nand U5880 (N_5880,N_4331,N_4906);
xnor U5881 (N_5881,N_4495,N_4441);
xor U5882 (N_5882,N_4931,N_4212);
nand U5883 (N_5883,N_4555,N_4267);
and U5884 (N_5884,N_4122,N_4502);
and U5885 (N_5885,N_4693,N_4116);
nor U5886 (N_5886,N_4048,N_4938);
and U5887 (N_5887,N_4509,N_4609);
or U5888 (N_5888,N_4617,N_4165);
nor U5889 (N_5889,N_4139,N_4932);
or U5890 (N_5890,N_4508,N_4044);
nor U5891 (N_5891,N_4010,N_4316);
xnor U5892 (N_5892,N_4086,N_4226);
nand U5893 (N_5893,N_4724,N_4175);
and U5894 (N_5894,N_4665,N_4415);
xnor U5895 (N_5895,N_4814,N_4148);
nand U5896 (N_5896,N_4818,N_4195);
or U5897 (N_5897,N_4279,N_4408);
nand U5898 (N_5898,N_4204,N_4959);
xor U5899 (N_5899,N_4104,N_4439);
xor U5900 (N_5900,N_4462,N_4825);
or U5901 (N_5901,N_4182,N_4243);
nor U5902 (N_5902,N_4716,N_4677);
and U5903 (N_5903,N_4256,N_4697);
and U5904 (N_5904,N_4573,N_4034);
or U5905 (N_5905,N_4207,N_4570);
or U5906 (N_5906,N_4465,N_4650);
and U5907 (N_5907,N_4906,N_4893);
xor U5908 (N_5908,N_4969,N_4339);
and U5909 (N_5909,N_4745,N_4823);
nor U5910 (N_5910,N_4100,N_4910);
nand U5911 (N_5911,N_4461,N_4886);
or U5912 (N_5912,N_4653,N_4525);
nor U5913 (N_5913,N_4631,N_4257);
or U5914 (N_5914,N_4338,N_4670);
nand U5915 (N_5915,N_4544,N_4931);
xnor U5916 (N_5916,N_4713,N_4869);
nand U5917 (N_5917,N_4114,N_4604);
and U5918 (N_5918,N_4542,N_4203);
and U5919 (N_5919,N_4730,N_4179);
and U5920 (N_5920,N_4098,N_4708);
or U5921 (N_5921,N_4405,N_4117);
and U5922 (N_5922,N_4639,N_4293);
xor U5923 (N_5923,N_4061,N_4072);
and U5924 (N_5924,N_4390,N_4642);
nor U5925 (N_5925,N_4227,N_4386);
and U5926 (N_5926,N_4547,N_4149);
and U5927 (N_5927,N_4010,N_4944);
xnor U5928 (N_5928,N_4458,N_4776);
xor U5929 (N_5929,N_4726,N_4025);
nand U5930 (N_5930,N_4836,N_4991);
or U5931 (N_5931,N_4833,N_4657);
and U5932 (N_5932,N_4551,N_4694);
or U5933 (N_5933,N_4539,N_4347);
xnor U5934 (N_5934,N_4206,N_4132);
and U5935 (N_5935,N_4666,N_4949);
nand U5936 (N_5936,N_4547,N_4985);
nand U5937 (N_5937,N_4860,N_4439);
nand U5938 (N_5938,N_4623,N_4119);
and U5939 (N_5939,N_4124,N_4108);
nand U5940 (N_5940,N_4908,N_4738);
and U5941 (N_5941,N_4933,N_4389);
xnor U5942 (N_5942,N_4157,N_4406);
or U5943 (N_5943,N_4700,N_4862);
xor U5944 (N_5944,N_4451,N_4391);
nor U5945 (N_5945,N_4109,N_4232);
or U5946 (N_5946,N_4388,N_4964);
or U5947 (N_5947,N_4130,N_4157);
nor U5948 (N_5948,N_4855,N_4328);
nand U5949 (N_5949,N_4668,N_4824);
or U5950 (N_5950,N_4880,N_4246);
nand U5951 (N_5951,N_4361,N_4759);
nand U5952 (N_5952,N_4681,N_4798);
and U5953 (N_5953,N_4945,N_4704);
or U5954 (N_5954,N_4567,N_4863);
nand U5955 (N_5955,N_4561,N_4973);
xnor U5956 (N_5956,N_4810,N_4528);
nand U5957 (N_5957,N_4228,N_4459);
xor U5958 (N_5958,N_4859,N_4880);
or U5959 (N_5959,N_4875,N_4383);
and U5960 (N_5960,N_4806,N_4154);
and U5961 (N_5961,N_4708,N_4030);
or U5962 (N_5962,N_4431,N_4443);
nand U5963 (N_5963,N_4773,N_4253);
xnor U5964 (N_5964,N_4019,N_4381);
nor U5965 (N_5965,N_4041,N_4171);
xnor U5966 (N_5966,N_4976,N_4490);
and U5967 (N_5967,N_4357,N_4569);
nor U5968 (N_5968,N_4772,N_4902);
or U5969 (N_5969,N_4967,N_4152);
and U5970 (N_5970,N_4831,N_4930);
nand U5971 (N_5971,N_4431,N_4104);
xor U5972 (N_5972,N_4655,N_4252);
or U5973 (N_5973,N_4161,N_4778);
nand U5974 (N_5974,N_4025,N_4795);
or U5975 (N_5975,N_4762,N_4034);
nand U5976 (N_5976,N_4340,N_4213);
nand U5977 (N_5977,N_4526,N_4938);
or U5978 (N_5978,N_4246,N_4132);
nor U5979 (N_5979,N_4786,N_4682);
or U5980 (N_5980,N_4404,N_4859);
or U5981 (N_5981,N_4947,N_4436);
or U5982 (N_5982,N_4375,N_4331);
or U5983 (N_5983,N_4122,N_4050);
xor U5984 (N_5984,N_4803,N_4685);
and U5985 (N_5985,N_4120,N_4580);
and U5986 (N_5986,N_4894,N_4917);
nand U5987 (N_5987,N_4791,N_4365);
xor U5988 (N_5988,N_4785,N_4026);
nand U5989 (N_5989,N_4452,N_4090);
or U5990 (N_5990,N_4556,N_4829);
nand U5991 (N_5991,N_4509,N_4624);
or U5992 (N_5992,N_4927,N_4243);
nor U5993 (N_5993,N_4396,N_4552);
nor U5994 (N_5994,N_4041,N_4589);
xnor U5995 (N_5995,N_4073,N_4279);
and U5996 (N_5996,N_4482,N_4484);
nand U5997 (N_5997,N_4847,N_4059);
and U5998 (N_5998,N_4447,N_4862);
nor U5999 (N_5999,N_4037,N_4602);
or U6000 (N_6000,N_5907,N_5603);
and U6001 (N_6001,N_5678,N_5873);
nand U6002 (N_6002,N_5789,N_5507);
xnor U6003 (N_6003,N_5473,N_5087);
nor U6004 (N_6004,N_5876,N_5656);
nand U6005 (N_6005,N_5301,N_5872);
or U6006 (N_6006,N_5016,N_5319);
nand U6007 (N_6007,N_5897,N_5639);
nand U6008 (N_6008,N_5042,N_5403);
xnor U6009 (N_6009,N_5485,N_5154);
and U6010 (N_6010,N_5327,N_5129);
nand U6011 (N_6011,N_5882,N_5350);
nor U6012 (N_6012,N_5927,N_5256);
nand U6013 (N_6013,N_5930,N_5431);
and U6014 (N_6014,N_5267,N_5901);
xor U6015 (N_6015,N_5516,N_5850);
xnor U6016 (N_6016,N_5264,N_5309);
xor U6017 (N_6017,N_5034,N_5056);
nand U6018 (N_6018,N_5620,N_5320);
nor U6019 (N_6019,N_5462,N_5705);
or U6020 (N_6020,N_5112,N_5941);
or U6021 (N_6021,N_5675,N_5402);
nor U6022 (N_6022,N_5800,N_5008);
and U6023 (N_6023,N_5219,N_5415);
and U6024 (N_6024,N_5761,N_5020);
xnor U6025 (N_6025,N_5381,N_5704);
and U6026 (N_6026,N_5802,N_5839);
or U6027 (N_6027,N_5856,N_5725);
or U6028 (N_6028,N_5973,N_5749);
or U6029 (N_6029,N_5121,N_5125);
nand U6030 (N_6030,N_5660,N_5292);
nor U6031 (N_6031,N_5239,N_5191);
and U6032 (N_6032,N_5146,N_5242);
nand U6033 (N_6033,N_5086,N_5611);
nand U6034 (N_6034,N_5355,N_5065);
xnor U6035 (N_6035,N_5547,N_5263);
nand U6036 (N_6036,N_5073,N_5149);
and U6037 (N_6037,N_5390,N_5985);
nor U6038 (N_6038,N_5898,N_5364);
or U6039 (N_6039,N_5829,N_5550);
or U6040 (N_6040,N_5614,N_5870);
nor U6041 (N_6041,N_5312,N_5588);
and U6042 (N_6042,N_5427,N_5579);
or U6043 (N_6043,N_5464,N_5774);
or U6044 (N_6044,N_5230,N_5047);
or U6045 (N_6045,N_5088,N_5158);
and U6046 (N_6046,N_5541,N_5006);
nand U6047 (N_6047,N_5497,N_5391);
or U6048 (N_6048,N_5680,N_5892);
nand U6049 (N_6049,N_5116,N_5643);
and U6050 (N_6050,N_5176,N_5801);
xor U6051 (N_6051,N_5366,N_5270);
or U6052 (N_6052,N_5583,N_5720);
nor U6053 (N_6053,N_5529,N_5666);
and U6054 (N_6054,N_5947,N_5616);
or U6055 (N_6055,N_5069,N_5100);
and U6056 (N_6056,N_5492,N_5997);
and U6057 (N_6057,N_5508,N_5834);
nand U6058 (N_6058,N_5463,N_5280);
nand U6059 (N_6059,N_5605,N_5661);
xor U6060 (N_6060,N_5282,N_5428);
nand U6061 (N_6061,N_5569,N_5686);
and U6062 (N_6062,N_5886,N_5582);
and U6063 (N_6063,N_5424,N_5671);
or U6064 (N_6064,N_5739,N_5003);
nand U6065 (N_6065,N_5806,N_5394);
and U6066 (N_6066,N_5468,N_5828);
or U6067 (N_6067,N_5912,N_5517);
nor U6068 (N_6068,N_5593,N_5352);
nand U6069 (N_6069,N_5759,N_5970);
xor U6070 (N_6070,N_5524,N_5096);
or U6071 (N_6071,N_5204,N_5826);
xor U6072 (N_6072,N_5181,N_5652);
and U6073 (N_6073,N_5337,N_5330);
or U6074 (N_6074,N_5438,N_5793);
and U6075 (N_6075,N_5360,N_5887);
nand U6076 (N_6076,N_5931,N_5689);
and U6077 (N_6077,N_5226,N_5799);
nor U6078 (N_6078,N_5119,N_5079);
nor U6079 (N_6079,N_5916,N_5142);
or U6080 (N_6080,N_5764,N_5991);
or U6081 (N_6081,N_5027,N_5693);
nor U6082 (N_6082,N_5388,N_5938);
or U6083 (N_6083,N_5198,N_5307);
nor U6084 (N_6084,N_5928,N_5228);
nor U6085 (N_6085,N_5284,N_5180);
and U6086 (N_6086,N_5030,N_5067);
xor U6087 (N_6087,N_5147,N_5920);
nor U6088 (N_6088,N_5383,N_5445);
nand U6089 (N_6089,N_5288,N_5184);
nand U6090 (N_6090,N_5225,N_5878);
nor U6091 (N_6091,N_5542,N_5037);
nand U6092 (N_6092,N_5838,N_5755);
nor U6093 (N_6093,N_5874,N_5268);
nand U6094 (N_6094,N_5854,N_5858);
xnor U6095 (N_6095,N_5363,N_5559);
nand U6096 (N_6096,N_5566,N_5714);
xnor U6097 (N_6097,N_5455,N_5905);
nor U6098 (N_6098,N_5115,N_5948);
or U6099 (N_6099,N_5676,N_5519);
or U6100 (N_6100,N_5279,N_5805);
nor U6101 (N_6101,N_5244,N_5963);
nor U6102 (N_6102,N_5724,N_5640);
xnor U6103 (N_6103,N_5193,N_5471);
and U6104 (N_6104,N_5078,N_5979);
and U6105 (N_6105,N_5695,N_5369);
nand U6106 (N_6106,N_5341,N_5013);
nand U6107 (N_6107,N_5083,N_5536);
and U6108 (N_6108,N_5012,N_5164);
or U6109 (N_6109,N_5744,N_5356);
nand U6110 (N_6110,N_5814,N_5000);
xnor U6111 (N_6111,N_5123,N_5071);
nand U6112 (N_6112,N_5945,N_5135);
and U6113 (N_6113,N_5861,N_5255);
or U6114 (N_6114,N_5532,N_5311);
and U6115 (N_6115,N_5038,N_5103);
and U6116 (N_6116,N_5189,N_5213);
nor U6117 (N_6117,N_5172,N_5097);
nor U6118 (N_6118,N_5241,N_5731);
or U6119 (N_6119,N_5664,N_5389);
xnor U6120 (N_6120,N_5503,N_5537);
and U6121 (N_6121,N_5227,N_5792);
nor U6122 (N_6122,N_5410,N_5325);
or U6123 (N_6123,N_5484,N_5405);
xnor U6124 (N_6124,N_5788,N_5830);
and U6125 (N_6125,N_5419,N_5051);
or U6126 (N_6126,N_5303,N_5106);
nor U6127 (N_6127,N_5883,N_5560);
xnor U6128 (N_6128,N_5223,N_5049);
nand U6129 (N_6129,N_5701,N_5090);
and U6130 (N_6130,N_5375,N_5632);
nor U6131 (N_6131,N_5551,N_5054);
or U6132 (N_6132,N_5203,N_5477);
xnor U6133 (N_6133,N_5766,N_5269);
xnor U6134 (N_6134,N_5214,N_5956);
and U6135 (N_6135,N_5893,N_5565);
or U6136 (N_6136,N_5563,N_5266);
and U6137 (N_6137,N_5348,N_5163);
nor U6138 (N_6138,N_5913,N_5216);
or U6139 (N_6139,N_5601,N_5148);
or U6140 (N_6140,N_5429,N_5253);
nand U6141 (N_6141,N_5776,N_5277);
xnor U6142 (N_6142,N_5846,N_5672);
nand U6143 (N_6143,N_5777,N_5107);
nand U6144 (N_6144,N_5592,N_5160);
or U6145 (N_6145,N_5345,N_5654);
nor U6146 (N_6146,N_5708,N_5716);
or U6147 (N_6147,N_5460,N_5845);
nor U6148 (N_6148,N_5141,N_5298);
xnor U6149 (N_6149,N_5753,N_5526);
nor U6150 (N_6150,N_5339,N_5314);
nor U6151 (N_6151,N_5059,N_5844);
and U6152 (N_6152,N_5732,N_5633);
or U6153 (N_6153,N_5752,N_5333);
and U6154 (N_6154,N_5796,N_5577);
nand U6155 (N_6155,N_5833,N_5265);
nor U6156 (N_6156,N_5118,N_5594);
xor U6157 (N_6157,N_5243,N_5919);
nor U6158 (N_6158,N_5804,N_5781);
nand U6159 (N_6159,N_5040,N_5807);
xnor U6160 (N_6160,N_5698,N_5498);
nor U6161 (N_6161,N_5981,N_5452);
xor U6162 (N_6162,N_5976,N_5412);
or U6163 (N_6163,N_5514,N_5868);
or U6164 (N_6164,N_5835,N_5756);
and U6165 (N_6165,N_5480,N_5548);
or U6166 (N_6166,N_5370,N_5983);
and U6167 (N_6167,N_5543,N_5949);
or U6168 (N_6168,N_5994,N_5426);
xor U6169 (N_6169,N_5523,N_5609);
or U6170 (N_6170,N_5033,N_5398);
and U6171 (N_6171,N_5336,N_5518);
xor U6172 (N_6172,N_5064,N_5943);
xnor U6173 (N_6173,N_5420,N_5124);
nor U6174 (N_6174,N_5585,N_5362);
nor U6175 (N_6175,N_5866,N_5074);
and U6176 (N_6176,N_5762,N_5702);
nor U6177 (N_6177,N_5031,N_5816);
xor U6178 (N_6178,N_5287,N_5760);
nor U6179 (N_6179,N_5200,N_5133);
or U6180 (N_6180,N_5029,N_5902);
or U6181 (N_6181,N_5599,N_5852);
or U6182 (N_6182,N_5053,N_5884);
xor U6183 (N_6183,N_5045,N_5153);
nand U6184 (N_6184,N_5323,N_5914);
xor U6185 (N_6185,N_5177,N_5344);
nand U6186 (N_6186,N_5433,N_5276);
or U6187 (N_6187,N_5556,N_5262);
and U6188 (N_6188,N_5354,N_5975);
and U6189 (N_6189,N_5260,N_5758);
and U6190 (N_6190,N_5466,N_5773);
or U6191 (N_6191,N_5824,N_5329);
or U6192 (N_6192,N_5722,N_5745);
or U6193 (N_6193,N_5554,N_5171);
nor U6194 (N_6194,N_5769,N_5746);
or U6195 (N_6195,N_5933,N_5023);
or U6196 (N_6196,N_5950,N_5767);
xor U6197 (N_6197,N_5990,N_5812);
nor U6198 (N_6198,N_5748,N_5965);
nand U6199 (N_6199,N_5940,N_5952);
and U6200 (N_6200,N_5231,N_5899);
xor U6201 (N_6201,N_5393,N_5969);
or U6202 (N_6202,N_5297,N_5785);
and U6203 (N_6203,N_5971,N_5891);
nor U6204 (N_6204,N_5044,N_5509);
xor U6205 (N_6205,N_5794,N_5063);
xor U6206 (N_6206,N_5808,N_5867);
nor U6207 (N_6207,N_5215,N_5677);
and U6208 (N_6208,N_5502,N_5019);
and U6209 (N_6209,N_5286,N_5659);
xnor U6210 (N_6210,N_5235,N_5010);
or U6211 (N_6211,N_5022,N_5864);
nor U6212 (N_6212,N_5499,N_5707);
xor U6213 (N_6213,N_5840,N_5778);
or U6214 (N_6214,N_5447,N_5351);
xnor U6215 (N_6215,N_5598,N_5472);
xnor U6216 (N_6216,N_5627,N_5888);
xnor U6217 (N_6217,N_5684,N_5076);
nor U6218 (N_6218,N_5557,N_5136);
nor U6219 (N_6219,N_5070,N_5454);
nor U6220 (N_6220,N_5757,N_5972);
xor U6221 (N_6221,N_5449,N_5169);
nand U6222 (N_6222,N_5437,N_5929);
and U6223 (N_6223,N_5951,N_5946);
and U6224 (N_6224,N_5111,N_5910);
or U6225 (N_6225,N_5934,N_5662);
nor U6226 (N_6226,N_5787,N_5205);
nor U6227 (N_6227,N_5634,N_5733);
xor U6228 (N_6228,N_5709,N_5495);
or U6229 (N_6229,N_5152,N_5906);
nor U6230 (N_6230,N_5335,N_5467);
xnor U6231 (N_6231,N_5909,N_5058);
nand U6232 (N_6232,N_5855,N_5150);
xnor U6233 (N_6233,N_5522,N_5966);
or U6234 (N_6234,N_5558,N_5607);
or U6235 (N_6235,N_5233,N_5430);
nor U6236 (N_6236,N_5657,N_5173);
nand U6237 (N_6237,N_5028,N_5823);
or U6238 (N_6238,N_5075,N_5168);
or U6239 (N_6239,N_5104,N_5877);
xnor U6240 (N_6240,N_5663,N_5359);
nor U6241 (N_6241,N_5655,N_5510);
xnor U6242 (N_6242,N_5458,N_5417);
and U6243 (N_6243,N_5977,N_5400);
xnor U6244 (N_6244,N_5290,N_5117);
nor U6245 (N_6245,N_5848,N_5857);
nor U6246 (N_6246,N_5317,N_5372);
and U6247 (N_6247,N_5612,N_5373);
and U6248 (N_6248,N_5957,N_5487);
nor U6249 (N_6249,N_5629,N_5797);
and U6250 (N_6250,N_5817,N_5580);
or U6251 (N_6251,N_5052,N_5863);
nor U6252 (N_6252,N_5576,N_5831);
and U6253 (N_6253,N_5347,N_5668);
or U6254 (N_6254,N_5224,N_5250);
nand U6255 (N_6255,N_5179,N_5122);
xor U6256 (N_6256,N_5025,N_5456);
xnor U6257 (N_6257,N_5474,N_5259);
and U6258 (N_6258,N_5316,N_5229);
or U6259 (N_6259,N_5544,N_5974);
and U6260 (N_6260,N_5005,N_5338);
and U6261 (N_6261,N_5326,N_5036);
and U6262 (N_6262,N_5322,N_5637);
nand U6263 (N_6263,N_5610,N_5289);
and U6264 (N_6264,N_5847,N_5880);
or U6265 (N_6265,N_5521,N_5192);
or U6266 (N_6266,N_5795,N_5525);
or U6267 (N_6267,N_5178,N_5751);
nand U6268 (N_6268,N_5679,N_5597);
xnor U6269 (N_6269,N_5315,N_5836);
nand U6270 (N_6270,N_5257,N_5651);
xor U6271 (N_6271,N_5367,N_5730);
xnor U6272 (N_6272,N_5217,N_5159);
or U6273 (N_6273,N_5143,N_5574);
nor U6274 (N_6274,N_5131,N_5889);
and U6275 (N_6275,N_5481,N_5258);
nand U6276 (N_6276,N_5763,N_5132);
and U6277 (N_6277,N_5349,N_5803);
nand U6278 (N_6278,N_5409,N_5780);
nor U6279 (N_6279,N_5923,N_5674);
and U6280 (N_6280,N_5469,N_5535);
nor U6281 (N_6281,N_5175,N_5182);
or U6282 (N_6282,N_5711,N_5822);
nor U6283 (N_6283,N_5055,N_5187);
xnor U6284 (N_6284,N_5735,N_5331);
xor U6285 (N_6285,N_5162,N_5515);
nand U6286 (N_6286,N_5723,N_5932);
or U6287 (N_6287,N_5306,N_5218);
nor U6288 (N_6288,N_5291,N_5682);
or U6289 (N_6289,N_5604,N_5470);
xor U6290 (N_6290,N_5134,N_5294);
or U6291 (N_6291,N_5128,N_5572);
nand U6292 (N_6292,N_5209,N_5685);
xnor U6293 (N_6293,N_5166,N_5505);
or U6294 (N_6294,N_5827,N_5486);
or U6295 (N_6295,N_5077,N_5591);
nor U6296 (N_6296,N_5493,N_5261);
and U6297 (N_6297,N_5986,N_5964);
nor U6298 (N_6298,N_5479,N_5696);
nor U6299 (N_6299,N_5528,N_5248);
and U6300 (N_6300,N_5500,N_5894);
xnor U6301 (N_6301,N_5924,N_5476);
or U6302 (N_6302,N_5283,N_5821);
nand U6303 (N_6303,N_5018,N_5623);
and U6304 (N_6304,N_5719,N_5407);
nor U6305 (N_6305,N_5304,N_5819);
or U6306 (N_6306,N_5046,N_5959);
or U6307 (N_6307,N_5921,N_5721);
and U6308 (N_6308,N_5491,N_5254);
nand U6309 (N_6309,N_5453,N_5457);
nor U6310 (N_6310,N_5084,N_5099);
and U6311 (N_6311,N_5734,N_5353);
and U6312 (N_6312,N_5137,N_5954);
or U6313 (N_6313,N_5413,N_5120);
nand U6314 (N_6314,N_5645,N_5552);
or U6315 (N_6315,N_5531,N_5108);
or U6316 (N_6316,N_5313,N_5618);
and U6317 (N_6317,N_5813,N_5386);
or U6318 (N_6318,N_5001,N_5207);
nand U6319 (N_6319,N_5841,N_5962);
nor U6320 (N_6320,N_5057,N_5396);
nand U6321 (N_6321,N_5443,N_5195);
or U6322 (N_6322,N_5667,N_5860);
nor U6323 (N_6323,N_5451,N_5770);
nor U6324 (N_6324,N_5904,N_5414);
and U6325 (N_6325,N_5953,N_5436);
xnor U6326 (N_6326,N_5561,N_5376);
and U6327 (N_6327,N_5617,N_5918);
xor U6328 (N_6328,N_5922,N_5527);
nor U6329 (N_6329,N_5729,N_5595);
xor U6330 (N_6330,N_5619,N_5811);
xnor U6331 (N_6331,N_5700,N_5385);
or U6332 (N_6332,N_5300,N_5377);
and U6333 (N_6333,N_5202,N_5533);
xnor U6334 (N_6334,N_5395,N_5201);
and U6335 (N_6335,N_5513,N_5600);
or U6336 (N_6336,N_5140,N_5843);
or U6337 (N_6337,N_5138,N_5996);
and U6338 (N_6338,N_5387,N_5697);
or U6339 (N_6339,N_5423,N_5881);
nand U6340 (N_6340,N_5139,N_5092);
nand U6341 (N_6341,N_5562,N_5435);
nor U6342 (N_6342,N_5450,N_5622);
xor U6343 (N_6343,N_5581,N_5465);
xor U6344 (N_6344,N_5271,N_5397);
xor U6345 (N_6345,N_5890,N_5713);
and U6346 (N_6346,N_5825,N_5853);
nand U6347 (N_6347,N_5903,N_5862);
nor U6348 (N_6348,N_5236,N_5737);
and U6349 (N_6349,N_5982,N_5590);
nor U6350 (N_6350,N_5165,N_5710);
nand U6351 (N_6351,N_5692,N_5081);
nor U6352 (N_6352,N_5130,N_5371);
and U6353 (N_6353,N_5098,N_5538);
xnor U6354 (N_6354,N_5285,N_5900);
and U6355 (N_6355,N_5673,N_5775);
xnor U6356 (N_6356,N_5810,N_5411);
or U6357 (N_6357,N_5448,N_5418);
nor U6358 (N_6358,N_5728,N_5174);
or U6359 (N_6359,N_5095,N_5658);
xor U6360 (N_6360,N_5185,N_5818);
xnor U6361 (N_6361,N_5043,N_5621);
xnor U6362 (N_6362,N_5157,N_5727);
and U6363 (N_6363,N_5343,N_5589);
and U6364 (N_6364,N_5186,N_5534);
xnor U6365 (N_6365,N_5779,N_5101);
xnor U6366 (N_6366,N_5832,N_5444);
or U6367 (N_6367,N_5439,N_5608);
or U6368 (N_6368,N_5014,N_5050);
nor U6369 (N_6369,N_5308,N_5082);
and U6370 (N_6370,N_5293,N_5626);
nor U6371 (N_6371,N_5879,N_5571);
xnor U6372 (N_6372,N_5520,N_5568);
nor U6373 (N_6373,N_5549,N_5489);
xor U6374 (N_6374,N_5332,N_5606);
nor U6375 (N_6375,N_5635,N_5988);
nor U6376 (N_6376,N_5602,N_5295);
xnor U6377 (N_6377,N_5646,N_5578);
and U6378 (N_6378,N_5699,N_5992);
nand U6379 (N_6379,N_5404,N_5302);
or U6380 (N_6380,N_5512,N_5978);
nor U6381 (N_6381,N_5305,N_5066);
or U6382 (N_6382,N_5274,N_5488);
or U6383 (N_6383,N_5741,N_5815);
xor U6384 (N_6384,N_5432,N_5167);
and U6385 (N_6385,N_5401,N_5908);
and U6386 (N_6386,N_5478,N_5380);
nand U6387 (N_6387,N_5220,N_5015);
nand U6388 (N_6388,N_5506,N_5670);
nand U6389 (N_6389,N_5002,N_5384);
nor U6390 (N_6390,N_5007,N_5851);
or U6391 (N_6391,N_5688,N_5272);
xnor U6392 (N_6392,N_5546,N_5939);
xor U6393 (N_6393,N_5772,N_5669);
nor U6394 (N_6394,N_5252,N_5555);
nand U6395 (N_6395,N_5747,N_5368);
or U6396 (N_6396,N_5357,N_5736);
or U6397 (N_6397,N_5809,N_5511);
nand U6398 (N_6398,N_5278,N_5416);
xnor U6399 (N_6399,N_5342,N_5726);
nor U6400 (N_6400,N_5089,N_5026);
nand U6401 (N_6401,N_5379,N_5820);
nor U6402 (N_6402,N_5190,N_5683);
nand U6403 (N_6403,N_5221,N_5211);
nor U6404 (N_6404,N_5238,N_5647);
and U6405 (N_6405,N_5496,N_5573);
nand U6406 (N_6406,N_5786,N_5170);
nor U6407 (N_6407,N_5859,N_5771);
xnor U6408 (N_6408,N_5989,N_5068);
or U6409 (N_6409,N_5584,N_5754);
nor U6410 (N_6410,N_5378,N_5035);
and U6411 (N_6411,N_5461,N_5650);
and U6412 (N_6412,N_5743,N_5105);
or U6413 (N_6413,N_5009,N_5328);
nor U6414 (N_6414,N_5630,N_5374);
xor U6415 (N_6415,N_5738,N_5365);
nor U6416 (N_6416,N_5024,N_5564);
and U6417 (N_6417,N_5649,N_5482);
xnor U6418 (N_6418,N_5937,N_5060);
nand U6419 (N_6419,N_5712,N_5494);
nor U6420 (N_6420,N_5896,N_5798);
nand U6421 (N_6421,N_5980,N_5871);
or U6422 (N_6422,N_5540,N_5628);
and U6423 (N_6423,N_5987,N_5783);
nor U6424 (N_6424,N_5895,N_5665);
nand U6425 (N_6425,N_5340,N_5837);
nor U6426 (N_6426,N_5197,N_5791);
and U6427 (N_6427,N_5275,N_5995);
nand U6428 (N_6428,N_5199,N_5249);
or U6429 (N_6429,N_5425,N_5936);
xnor U6430 (N_6430,N_5039,N_5869);
or U6431 (N_6431,N_5032,N_5631);
nor U6432 (N_6432,N_5358,N_5596);
nand U6433 (N_6433,N_5504,N_5212);
nor U6434 (N_6434,N_5382,N_5094);
and U6435 (N_6435,N_5334,N_5072);
or U6436 (N_6436,N_5145,N_5392);
nor U6437 (N_6437,N_5984,N_5321);
xor U6438 (N_6438,N_5690,N_5232);
nor U6439 (N_6439,N_5422,N_5183);
or U6440 (N_6440,N_5636,N_5080);
nand U6441 (N_6441,N_5641,N_5062);
or U6442 (N_6442,N_5296,N_5750);
xor U6443 (N_6443,N_5110,N_5644);
and U6444 (N_6444,N_5717,N_5126);
nor U6445 (N_6445,N_5586,N_5102);
and U6446 (N_6446,N_5399,N_5742);
nor U6447 (N_6447,N_5648,N_5361);
nand U6448 (N_6448,N_5567,N_5993);
nand U6449 (N_6449,N_5790,N_5251);
nor U6450 (N_6450,N_5206,N_5151);
nand U6451 (N_6451,N_5715,N_5091);
or U6452 (N_6452,N_5475,N_5017);
or U6453 (N_6453,N_5539,N_5247);
or U6454 (N_6454,N_5483,N_5113);
xnor U6455 (N_6455,N_5849,N_5782);
or U6456 (N_6456,N_5246,N_5346);
or U6457 (N_6457,N_5653,N_5545);
and U6458 (N_6458,N_5310,N_5011);
xor U6459 (N_6459,N_5703,N_5196);
xnor U6460 (N_6460,N_5434,N_5638);
nand U6461 (N_6461,N_5915,N_5406);
or U6462 (N_6462,N_5967,N_5061);
nor U6463 (N_6463,N_5625,N_5109);
xor U6464 (N_6464,N_5208,N_5240);
xor U6465 (N_6465,N_5530,N_5441);
or U6466 (N_6466,N_5875,N_5935);
nor U6467 (N_6467,N_5570,N_5188);
or U6468 (N_6468,N_5575,N_5004);
xor U6469 (N_6469,N_5917,N_5885);
and U6470 (N_6470,N_5156,N_5926);
nor U6471 (N_6471,N_5245,N_5865);
nand U6472 (N_6472,N_5968,N_5442);
or U6473 (N_6473,N_5446,N_5842);
nand U6474 (N_6474,N_5960,N_5021);
nor U6475 (N_6475,N_5127,N_5687);
nand U6476 (N_6476,N_5681,N_5273);
nor U6477 (N_6477,N_5161,N_5041);
or U6478 (N_6478,N_5085,N_5955);
or U6479 (N_6479,N_5925,N_5155);
or U6480 (N_6480,N_5318,N_5691);
or U6481 (N_6481,N_5615,N_5144);
xnor U6482 (N_6482,N_5440,N_5421);
xor U6483 (N_6483,N_5237,N_5210);
xnor U6484 (N_6484,N_5587,N_5299);
and U6485 (N_6485,N_5093,N_5706);
nand U6486 (N_6486,N_5768,N_5958);
nor U6487 (N_6487,N_5613,N_5114);
nor U6488 (N_6488,N_5408,N_5765);
xnor U6489 (N_6489,N_5694,N_5942);
xor U6490 (N_6490,N_5501,N_5624);
xor U6491 (N_6491,N_5234,N_5999);
xor U6492 (N_6492,N_5553,N_5961);
nor U6493 (N_6493,N_5718,N_5222);
nand U6494 (N_6494,N_5194,N_5998);
nand U6495 (N_6495,N_5784,N_5048);
xnor U6496 (N_6496,N_5459,N_5490);
nand U6497 (N_6497,N_5740,N_5642);
nand U6498 (N_6498,N_5944,N_5324);
and U6499 (N_6499,N_5911,N_5281);
nor U6500 (N_6500,N_5077,N_5552);
nand U6501 (N_6501,N_5322,N_5927);
nand U6502 (N_6502,N_5621,N_5146);
or U6503 (N_6503,N_5000,N_5110);
or U6504 (N_6504,N_5043,N_5118);
or U6505 (N_6505,N_5906,N_5274);
nor U6506 (N_6506,N_5939,N_5702);
or U6507 (N_6507,N_5789,N_5484);
nand U6508 (N_6508,N_5777,N_5476);
xor U6509 (N_6509,N_5275,N_5106);
and U6510 (N_6510,N_5188,N_5987);
nor U6511 (N_6511,N_5043,N_5653);
xor U6512 (N_6512,N_5628,N_5373);
or U6513 (N_6513,N_5415,N_5463);
or U6514 (N_6514,N_5186,N_5252);
xor U6515 (N_6515,N_5180,N_5915);
nand U6516 (N_6516,N_5761,N_5408);
and U6517 (N_6517,N_5272,N_5529);
and U6518 (N_6518,N_5917,N_5312);
nor U6519 (N_6519,N_5392,N_5991);
nor U6520 (N_6520,N_5245,N_5238);
nand U6521 (N_6521,N_5533,N_5345);
nor U6522 (N_6522,N_5745,N_5121);
xnor U6523 (N_6523,N_5352,N_5736);
and U6524 (N_6524,N_5672,N_5347);
nor U6525 (N_6525,N_5668,N_5842);
nand U6526 (N_6526,N_5426,N_5186);
and U6527 (N_6527,N_5684,N_5516);
nor U6528 (N_6528,N_5338,N_5879);
or U6529 (N_6529,N_5103,N_5767);
and U6530 (N_6530,N_5588,N_5571);
and U6531 (N_6531,N_5086,N_5770);
xor U6532 (N_6532,N_5123,N_5996);
xnor U6533 (N_6533,N_5927,N_5196);
xnor U6534 (N_6534,N_5093,N_5705);
xnor U6535 (N_6535,N_5012,N_5953);
and U6536 (N_6536,N_5699,N_5146);
nor U6537 (N_6537,N_5129,N_5271);
nor U6538 (N_6538,N_5804,N_5081);
nor U6539 (N_6539,N_5918,N_5952);
and U6540 (N_6540,N_5851,N_5787);
and U6541 (N_6541,N_5695,N_5562);
and U6542 (N_6542,N_5318,N_5646);
nor U6543 (N_6543,N_5822,N_5540);
nor U6544 (N_6544,N_5614,N_5611);
nand U6545 (N_6545,N_5571,N_5857);
nor U6546 (N_6546,N_5960,N_5970);
nand U6547 (N_6547,N_5507,N_5071);
xor U6548 (N_6548,N_5026,N_5913);
nand U6549 (N_6549,N_5132,N_5709);
and U6550 (N_6550,N_5739,N_5443);
or U6551 (N_6551,N_5061,N_5150);
nand U6552 (N_6552,N_5913,N_5401);
xnor U6553 (N_6553,N_5570,N_5287);
or U6554 (N_6554,N_5784,N_5097);
nor U6555 (N_6555,N_5891,N_5094);
and U6556 (N_6556,N_5735,N_5508);
or U6557 (N_6557,N_5229,N_5187);
xor U6558 (N_6558,N_5814,N_5774);
and U6559 (N_6559,N_5267,N_5363);
nand U6560 (N_6560,N_5293,N_5337);
nand U6561 (N_6561,N_5526,N_5886);
and U6562 (N_6562,N_5979,N_5943);
xor U6563 (N_6563,N_5884,N_5543);
nor U6564 (N_6564,N_5468,N_5771);
or U6565 (N_6565,N_5664,N_5351);
nand U6566 (N_6566,N_5325,N_5579);
nand U6567 (N_6567,N_5011,N_5292);
nor U6568 (N_6568,N_5761,N_5297);
and U6569 (N_6569,N_5088,N_5863);
nor U6570 (N_6570,N_5698,N_5380);
nor U6571 (N_6571,N_5646,N_5603);
and U6572 (N_6572,N_5475,N_5883);
and U6573 (N_6573,N_5743,N_5010);
or U6574 (N_6574,N_5764,N_5843);
xor U6575 (N_6575,N_5224,N_5078);
and U6576 (N_6576,N_5359,N_5906);
nor U6577 (N_6577,N_5128,N_5038);
or U6578 (N_6578,N_5121,N_5516);
xnor U6579 (N_6579,N_5963,N_5101);
nor U6580 (N_6580,N_5017,N_5305);
xnor U6581 (N_6581,N_5266,N_5373);
nor U6582 (N_6582,N_5237,N_5402);
xor U6583 (N_6583,N_5785,N_5261);
nand U6584 (N_6584,N_5007,N_5811);
and U6585 (N_6585,N_5289,N_5564);
nand U6586 (N_6586,N_5210,N_5230);
nor U6587 (N_6587,N_5228,N_5115);
or U6588 (N_6588,N_5348,N_5054);
nand U6589 (N_6589,N_5146,N_5996);
or U6590 (N_6590,N_5757,N_5328);
and U6591 (N_6591,N_5209,N_5626);
or U6592 (N_6592,N_5970,N_5375);
nand U6593 (N_6593,N_5719,N_5680);
nor U6594 (N_6594,N_5754,N_5626);
nand U6595 (N_6595,N_5474,N_5324);
nand U6596 (N_6596,N_5385,N_5297);
xor U6597 (N_6597,N_5492,N_5738);
nand U6598 (N_6598,N_5725,N_5526);
and U6599 (N_6599,N_5455,N_5980);
or U6600 (N_6600,N_5615,N_5412);
nor U6601 (N_6601,N_5958,N_5883);
and U6602 (N_6602,N_5088,N_5995);
or U6603 (N_6603,N_5349,N_5901);
xor U6604 (N_6604,N_5129,N_5739);
nor U6605 (N_6605,N_5938,N_5603);
nor U6606 (N_6606,N_5597,N_5361);
or U6607 (N_6607,N_5096,N_5383);
nor U6608 (N_6608,N_5925,N_5156);
nand U6609 (N_6609,N_5390,N_5001);
nand U6610 (N_6610,N_5091,N_5170);
nor U6611 (N_6611,N_5707,N_5395);
and U6612 (N_6612,N_5651,N_5056);
nand U6613 (N_6613,N_5184,N_5628);
nor U6614 (N_6614,N_5569,N_5570);
nor U6615 (N_6615,N_5666,N_5659);
or U6616 (N_6616,N_5518,N_5249);
xor U6617 (N_6617,N_5003,N_5542);
and U6618 (N_6618,N_5346,N_5813);
nand U6619 (N_6619,N_5777,N_5367);
and U6620 (N_6620,N_5020,N_5061);
nor U6621 (N_6621,N_5472,N_5916);
or U6622 (N_6622,N_5544,N_5744);
xnor U6623 (N_6623,N_5038,N_5714);
xnor U6624 (N_6624,N_5394,N_5342);
and U6625 (N_6625,N_5539,N_5662);
nor U6626 (N_6626,N_5606,N_5212);
or U6627 (N_6627,N_5121,N_5262);
or U6628 (N_6628,N_5549,N_5394);
nor U6629 (N_6629,N_5793,N_5188);
nand U6630 (N_6630,N_5911,N_5415);
xor U6631 (N_6631,N_5502,N_5242);
nor U6632 (N_6632,N_5679,N_5165);
nand U6633 (N_6633,N_5041,N_5611);
and U6634 (N_6634,N_5774,N_5547);
and U6635 (N_6635,N_5930,N_5567);
or U6636 (N_6636,N_5787,N_5180);
and U6637 (N_6637,N_5030,N_5560);
or U6638 (N_6638,N_5721,N_5927);
nand U6639 (N_6639,N_5842,N_5323);
and U6640 (N_6640,N_5222,N_5846);
xnor U6641 (N_6641,N_5302,N_5628);
and U6642 (N_6642,N_5839,N_5296);
and U6643 (N_6643,N_5965,N_5157);
xnor U6644 (N_6644,N_5367,N_5089);
xor U6645 (N_6645,N_5586,N_5471);
nand U6646 (N_6646,N_5394,N_5684);
and U6647 (N_6647,N_5367,N_5953);
nand U6648 (N_6648,N_5813,N_5364);
xor U6649 (N_6649,N_5009,N_5190);
nor U6650 (N_6650,N_5648,N_5068);
and U6651 (N_6651,N_5033,N_5707);
nor U6652 (N_6652,N_5517,N_5421);
or U6653 (N_6653,N_5336,N_5797);
or U6654 (N_6654,N_5777,N_5885);
or U6655 (N_6655,N_5483,N_5691);
and U6656 (N_6656,N_5543,N_5244);
or U6657 (N_6657,N_5689,N_5548);
and U6658 (N_6658,N_5965,N_5913);
and U6659 (N_6659,N_5763,N_5672);
nand U6660 (N_6660,N_5205,N_5436);
and U6661 (N_6661,N_5491,N_5282);
nand U6662 (N_6662,N_5220,N_5524);
and U6663 (N_6663,N_5978,N_5232);
or U6664 (N_6664,N_5104,N_5770);
nand U6665 (N_6665,N_5136,N_5379);
nor U6666 (N_6666,N_5537,N_5165);
and U6667 (N_6667,N_5346,N_5535);
and U6668 (N_6668,N_5974,N_5367);
or U6669 (N_6669,N_5764,N_5620);
nand U6670 (N_6670,N_5719,N_5606);
nor U6671 (N_6671,N_5024,N_5463);
and U6672 (N_6672,N_5344,N_5175);
and U6673 (N_6673,N_5784,N_5435);
xor U6674 (N_6674,N_5896,N_5074);
xnor U6675 (N_6675,N_5122,N_5324);
xnor U6676 (N_6676,N_5403,N_5691);
and U6677 (N_6677,N_5936,N_5324);
xnor U6678 (N_6678,N_5638,N_5184);
nor U6679 (N_6679,N_5053,N_5099);
nor U6680 (N_6680,N_5218,N_5523);
or U6681 (N_6681,N_5525,N_5601);
or U6682 (N_6682,N_5789,N_5887);
or U6683 (N_6683,N_5879,N_5560);
nor U6684 (N_6684,N_5777,N_5335);
and U6685 (N_6685,N_5179,N_5215);
or U6686 (N_6686,N_5912,N_5128);
and U6687 (N_6687,N_5544,N_5329);
xor U6688 (N_6688,N_5904,N_5755);
xor U6689 (N_6689,N_5628,N_5930);
and U6690 (N_6690,N_5935,N_5723);
and U6691 (N_6691,N_5282,N_5229);
and U6692 (N_6692,N_5696,N_5189);
or U6693 (N_6693,N_5338,N_5258);
or U6694 (N_6694,N_5802,N_5496);
xor U6695 (N_6695,N_5646,N_5087);
nor U6696 (N_6696,N_5718,N_5974);
nand U6697 (N_6697,N_5197,N_5324);
and U6698 (N_6698,N_5250,N_5927);
and U6699 (N_6699,N_5466,N_5715);
and U6700 (N_6700,N_5675,N_5021);
xnor U6701 (N_6701,N_5852,N_5887);
nand U6702 (N_6702,N_5970,N_5091);
and U6703 (N_6703,N_5050,N_5983);
and U6704 (N_6704,N_5338,N_5185);
nand U6705 (N_6705,N_5959,N_5468);
or U6706 (N_6706,N_5948,N_5237);
xnor U6707 (N_6707,N_5538,N_5218);
and U6708 (N_6708,N_5584,N_5779);
nand U6709 (N_6709,N_5910,N_5522);
and U6710 (N_6710,N_5110,N_5423);
and U6711 (N_6711,N_5855,N_5254);
nand U6712 (N_6712,N_5828,N_5330);
or U6713 (N_6713,N_5222,N_5900);
xor U6714 (N_6714,N_5329,N_5011);
nand U6715 (N_6715,N_5289,N_5442);
or U6716 (N_6716,N_5305,N_5948);
xor U6717 (N_6717,N_5925,N_5657);
or U6718 (N_6718,N_5372,N_5535);
or U6719 (N_6719,N_5843,N_5122);
xor U6720 (N_6720,N_5247,N_5770);
or U6721 (N_6721,N_5280,N_5142);
and U6722 (N_6722,N_5691,N_5965);
nand U6723 (N_6723,N_5029,N_5293);
nor U6724 (N_6724,N_5583,N_5136);
or U6725 (N_6725,N_5318,N_5506);
and U6726 (N_6726,N_5417,N_5442);
and U6727 (N_6727,N_5595,N_5139);
xor U6728 (N_6728,N_5473,N_5230);
nor U6729 (N_6729,N_5773,N_5168);
and U6730 (N_6730,N_5614,N_5945);
nor U6731 (N_6731,N_5681,N_5719);
and U6732 (N_6732,N_5693,N_5731);
nand U6733 (N_6733,N_5961,N_5109);
nor U6734 (N_6734,N_5123,N_5630);
nor U6735 (N_6735,N_5582,N_5141);
nor U6736 (N_6736,N_5211,N_5318);
xnor U6737 (N_6737,N_5579,N_5232);
xor U6738 (N_6738,N_5840,N_5794);
or U6739 (N_6739,N_5855,N_5142);
nor U6740 (N_6740,N_5293,N_5486);
xnor U6741 (N_6741,N_5383,N_5619);
nand U6742 (N_6742,N_5976,N_5439);
nand U6743 (N_6743,N_5667,N_5396);
xnor U6744 (N_6744,N_5791,N_5870);
nand U6745 (N_6745,N_5031,N_5472);
nand U6746 (N_6746,N_5873,N_5048);
nor U6747 (N_6747,N_5016,N_5064);
and U6748 (N_6748,N_5962,N_5918);
nand U6749 (N_6749,N_5701,N_5391);
and U6750 (N_6750,N_5648,N_5954);
nor U6751 (N_6751,N_5841,N_5105);
and U6752 (N_6752,N_5154,N_5982);
xor U6753 (N_6753,N_5603,N_5285);
or U6754 (N_6754,N_5229,N_5562);
nand U6755 (N_6755,N_5659,N_5241);
and U6756 (N_6756,N_5535,N_5115);
nand U6757 (N_6757,N_5143,N_5003);
or U6758 (N_6758,N_5275,N_5760);
nor U6759 (N_6759,N_5899,N_5375);
or U6760 (N_6760,N_5054,N_5399);
or U6761 (N_6761,N_5532,N_5608);
and U6762 (N_6762,N_5608,N_5617);
or U6763 (N_6763,N_5086,N_5590);
nor U6764 (N_6764,N_5856,N_5575);
or U6765 (N_6765,N_5521,N_5335);
or U6766 (N_6766,N_5797,N_5012);
nor U6767 (N_6767,N_5207,N_5098);
nor U6768 (N_6768,N_5786,N_5958);
and U6769 (N_6769,N_5603,N_5465);
and U6770 (N_6770,N_5314,N_5383);
xor U6771 (N_6771,N_5847,N_5738);
or U6772 (N_6772,N_5288,N_5576);
nand U6773 (N_6773,N_5346,N_5052);
nor U6774 (N_6774,N_5183,N_5092);
xor U6775 (N_6775,N_5297,N_5172);
nand U6776 (N_6776,N_5862,N_5210);
xnor U6777 (N_6777,N_5238,N_5546);
nand U6778 (N_6778,N_5862,N_5556);
and U6779 (N_6779,N_5769,N_5334);
xnor U6780 (N_6780,N_5472,N_5456);
and U6781 (N_6781,N_5458,N_5626);
nor U6782 (N_6782,N_5235,N_5278);
nor U6783 (N_6783,N_5501,N_5479);
and U6784 (N_6784,N_5376,N_5627);
nand U6785 (N_6785,N_5103,N_5708);
xnor U6786 (N_6786,N_5589,N_5870);
and U6787 (N_6787,N_5265,N_5994);
and U6788 (N_6788,N_5930,N_5968);
nand U6789 (N_6789,N_5304,N_5900);
nor U6790 (N_6790,N_5240,N_5590);
xor U6791 (N_6791,N_5137,N_5707);
and U6792 (N_6792,N_5679,N_5574);
and U6793 (N_6793,N_5470,N_5884);
xor U6794 (N_6794,N_5954,N_5766);
or U6795 (N_6795,N_5411,N_5923);
nor U6796 (N_6796,N_5101,N_5039);
nor U6797 (N_6797,N_5198,N_5258);
xor U6798 (N_6798,N_5588,N_5814);
and U6799 (N_6799,N_5311,N_5417);
and U6800 (N_6800,N_5196,N_5295);
nand U6801 (N_6801,N_5336,N_5448);
nand U6802 (N_6802,N_5113,N_5370);
nor U6803 (N_6803,N_5519,N_5163);
nand U6804 (N_6804,N_5468,N_5505);
and U6805 (N_6805,N_5010,N_5411);
or U6806 (N_6806,N_5575,N_5018);
and U6807 (N_6807,N_5233,N_5084);
and U6808 (N_6808,N_5887,N_5370);
or U6809 (N_6809,N_5532,N_5702);
nand U6810 (N_6810,N_5589,N_5184);
or U6811 (N_6811,N_5717,N_5893);
nand U6812 (N_6812,N_5729,N_5328);
or U6813 (N_6813,N_5850,N_5694);
xor U6814 (N_6814,N_5021,N_5635);
xor U6815 (N_6815,N_5181,N_5187);
nand U6816 (N_6816,N_5267,N_5850);
nor U6817 (N_6817,N_5882,N_5666);
nor U6818 (N_6818,N_5092,N_5782);
nor U6819 (N_6819,N_5768,N_5021);
and U6820 (N_6820,N_5090,N_5575);
or U6821 (N_6821,N_5777,N_5457);
nor U6822 (N_6822,N_5488,N_5449);
or U6823 (N_6823,N_5048,N_5095);
and U6824 (N_6824,N_5929,N_5417);
nor U6825 (N_6825,N_5186,N_5142);
or U6826 (N_6826,N_5642,N_5259);
xor U6827 (N_6827,N_5648,N_5608);
or U6828 (N_6828,N_5391,N_5095);
nor U6829 (N_6829,N_5875,N_5234);
or U6830 (N_6830,N_5576,N_5240);
xnor U6831 (N_6831,N_5204,N_5437);
xnor U6832 (N_6832,N_5433,N_5969);
and U6833 (N_6833,N_5462,N_5587);
xnor U6834 (N_6834,N_5016,N_5030);
nand U6835 (N_6835,N_5247,N_5025);
nand U6836 (N_6836,N_5233,N_5024);
and U6837 (N_6837,N_5061,N_5394);
and U6838 (N_6838,N_5866,N_5539);
or U6839 (N_6839,N_5353,N_5746);
and U6840 (N_6840,N_5075,N_5239);
or U6841 (N_6841,N_5959,N_5124);
nand U6842 (N_6842,N_5129,N_5671);
nor U6843 (N_6843,N_5818,N_5550);
or U6844 (N_6844,N_5419,N_5884);
or U6845 (N_6845,N_5730,N_5894);
xor U6846 (N_6846,N_5499,N_5272);
or U6847 (N_6847,N_5142,N_5951);
nor U6848 (N_6848,N_5664,N_5974);
nor U6849 (N_6849,N_5611,N_5154);
xor U6850 (N_6850,N_5412,N_5765);
and U6851 (N_6851,N_5331,N_5800);
nand U6852 (N_6852,N_5278,N_5831);
and U6853 (N_6853,N_5818,N_5518);
xnor U6854 (N_6854,N_5762,N_5085);
nand U6855 (N_6855,N_5398,N_5371);
nor U6856 (N_6856,N_5342,N_5356);
or U6857 (N_6857,N_5287,N_5559);
and U6858 (N_6858,N_5670,N_5981);
or U6859 (N_6859,N_5143,N_5414);
nor U6860 (N_6860,N_5988,N_5272);
and U6861 (N_6861,N_5731,N_5770);
or U6862 (N_6862,N_5423,N_5221);
nor U6863 (N_6863,N_5778,N_5960);
or U6864 (N_6864,N_5847,N_5913);
xnor U6865 (N_6865,N_5209,N_5570);
xnor U6866 (N_6866,N_5235,N_5705);
nand U6867 (N_6867,N_5810,N_5361);
or U6868 (N_6868,N_5365,N_5285);
nor U6869 (N_6869,N_5996,N_5620);
xor U6870 (N_6870,N_5894,N_5013);
xor U6871 (N_6871,N_5638,N_5302);
xor U6872 (N_6872,N_5155,N_5799);
xnor U6873 (N_6873,N_5617,N_5523);
xor U6874 (N_6874,N_5966,N_5450);
and U6875 (N_6875,N_5968,N_5362);
nor U6876 (N_6876,N_5928,N_5065);
nor U6877 (N_6877,N_5108,N_5383);
nor U6878 (N_6878,N_5342,N_5993);
nor U6879 (N_6879,N_5127,N_5290);
or U6880 (N_6880,N_5285,N_5532);
nor U6881 (N_6881,N_5892,N_5043);
xnor U6882 (N_6882,N_5876,N_5119);
nand U6883 (N_6883,N_5625,N_5676);
xor U6884 (N_6884,N_5582,N_5390);
nand U6885 (N_6885,N_5710,N_5516);
xor U6886 (N_6886,N_5933,N_5807);
or U6887 (N_6887,N_5351,N_5883);
xnor U6888 (N_6888,N_5814,N_5334);
xor U6889 (N_6889,N_5234,N_5548);
or U6890 (N_6890,N_5346,N_5105);
nor U6891 (N_6891,N_5466,N_5780);
or U6892 (N_6892,N_5563,N_5679);
nand U6893 (N_6893,N_5567,N_5929);
nor U6894 (N_6894,N_5904,N_5540);
nand U6895 (N_6895,N_5057,N_5795);
xor U6896 (N_6896,N_5349,N_5062);
or U6897 (N_6897,N_5627,N_5984);
and U6898 (N_6898,N_5220,N_5305);
and U6899 (N_6899,N_5426,N_5442);
or U6900 (N_6900,N_5061,N_5806);
nand U6901 (N_6901,N_5423,N_5367);
nor U6902 (N_6902,N_5115,N_5236);
or U6903 (N_6903,N_5439,N_5420);
or U6904 (N_6904,N_5860,N_5414);
and U6905 (N_6905,N_5219,N_5894);
nand U6906 (N_6906,N_5550,N_5463);
xnor U6907 (N_6907,N_5179,N_5752);
xnor U6908 (N_6908,N_5045,N_5260);
or U6909 (N_6909,N_5057,N_5159);
or U6910 (N_6910,N_5548,N_5237);
or U6911 (N_6911,N_5864,N_5677);
xnor U6912 (N_6912,N_5833,N_5438);
or U6913 (N_6913,N_5841,N_5890);
nor U6914 (N_6914,N_5683,N_5261);
nand U6915 (N_6915,N_5177,N_5269);
xor U6916 (N_6916,N_5299,N_5955);
xnor U6917 (N_6917,N_5705,N_5374);
or U6918 (N_6918,N_5686,N_5422);
nor U6919 (N_6919,N_5030,N_5132);
and U6920 (N_6920,N_5282,N_5107);
and U6921 (N_6921,N_5057,N_5455);
nor U6922 (N_6922,N_5612,N_5326);
nor U6923 (N_6923,N_5849,N_5523);
nor U6924 (N_6924,N_5352,N_5381);
or U6925 (N_6925,N_5792,N_5252);
and U6926 (N_6926,N_5023,N_5307);
and U6927 (N_6927,N_5267,N_5528);
nor U6928 (N_6928,N_5469,N_5244);
xor U6929 (N_6929,N_5554,N_5337);
xnor U6930 (N_6930,N_5686,N_5449);
or U6931 (N_6931,N_5151,N_5522);
xor U6932 (N_6932,N_5764,N_5603);
and U6933 (N_6933,N_5231,N_5255);
and U6934 (N_6934,N_5150,N_5323);
nor U6935 (N_6935,N_5522,N_5377);
or U6936 (N_6936,N_5714,N_5805);
nor U6937 (N_6937,N_5487,N_5416);
xor U6938 (N_6938,N_5878,N_5705);
or U6939 (N_6939,N_5073,N_5417);
nand U6940 (N_6940,N_5910,N_5958);
or U6941 (N_6941,N_5664,N_5763);
xnor U6942 (N_6942,N_5100,N_5743);
and U6943 (N_6943,N_5881,N_5677);
or U6944 (N_6944,N_5171,N_5086);
xor U6945 (N_6945,N_5389,N_5279);
or U6946 (N_6946,N_5163,N_5699);
nand U6947 (N_6947,N_5963,N_5141);
xnor U6948 (N_6948,N_5074,N_5674);
nor U6949 (N_6949,N_5278,N_5425);
nor U6950 (N_6950,N_5437,N_5232);
and U6951 (N_6951,N_5230,N_5506);
xnor U6952 (N_6952,N_5994,N_5831);
and U6953 (N_6953,N_5434,N_5090);
nand U6954 (N_6954,N_5754,N_5333);
xnor U6955 (N_6955,N_5882,N_5260);
nor U6956 (N_6956,N_5043,N_5639);
nor U6957 (N_6957,N_5398,N_5013);
and U6958 (N_6958,N_5367,N_5599);
xnor U6959 (N_6959,N_5650,N_5860);
nor U6960 (N_6960,N_5921,N_5076);
nor U6961 (N_6961,N_5273,N_5539);
nor U6962 (N_6962,N_5421,N_5918);
or U6963 (N_6963,N_5767,N_5663);
nor U6964 (N_6964,N_5382,N_5242);
nor U6965 (N_6965,N_5186,N_5418);
nor U6966 (N_6966,N_5214,N_5604);
or U6967 (N_6967,N_5909,N_5806);
nand U6968 (N_6968,N_5267,N_5654);
nand U6969 (N_6969,N_5731,N_5122);
nand U6970 (N_6970,N_5617,N_5780);
or U6971 (N_6971,N_5290,N_5384);
nand U6972 (N_6972,N_5599,N_5008);
or U6973 (N_6973,N_5137,N_5180);
xnor U6974 (N_6974,N_5206,N_5089);
xor U6975 (N_6975,N_5191,N_5238);
nand U6976 (N_6976,N_5111,N_5742);
and U6977 (N_6977,N_5345,N_5438);
xor U6978 (N_6978,N_5350,N_5576);
or U6979 (N_6979,N_5114,N_5904);
and U6980 (N_6980,N_5787,N_5557);
nand U6981 (N_6981,N_5401,N_5730);
xnor U6982 (N_6982,N_5223,N_5134);
and U6983 (N_6983,N_5351,N_5382);
nand U6984 (N_6984,N_5123,N_5363);
or U6985 (N_6985,N_5638,N_5781);
nand U6986 (N_6986,N_5195,N_5238);
xor U6987 (N_6987,N_5851,N_5168);
nand U6988 (N_6988,N_5854,N_5396);
or U6989 (N_6989,N_5738,N_5376);
xor U6990 (N_6990,N_5916,N_5155);
nor U6991 (N_6991,N_5300,N_5545);
or U6992 (N_6992,N_5728,N_5200);
xnor U6993 (N_6993,N_5403,N_5875);
or U6994 (N_6994,N_5088,N_5516);
nor U6995 (N_6995,N_5674,N_5179);
nand U6996 (N_6996,N_5597,N_5278);
nor U6997 (N_6997,N_5001,N_5571);
nor U6998 (N_6998,N_5587,N_5653);
or U6999 (N_6999,N_5396,N_5993);
nor U7000 (N_7000,N_6925,N_6068);
and U7001 (N_7001,N_6070,N_6502);
or U7002 (N_7002,N_6717,N_6791);
xor U7003 (N_7003,N_6125,N_6247);
or U7004 (N_7004,N_6965,N_6268);
nor U7005 (N_7005,N_6083,N_6968);
xnor U7006 (N_7006,N_6778,N_6138);
nand U7007 (N_7007,N_6693,N_6215);
or U7008 (N_7008,N_6029,N_6359);
nor U7009 (N_7009,N_6167,N_6098);
xnor U7010 (N_7010,N_6905,N_6042);
nand U7011 (N_7011,N_6869,N_6183);
xor U7012 (N_7012,N_6309,N_6976);
or U7013 (N_7013,N_6588,N_6746);
nand U7014 (N_7014,N_6766,N_6940);
and U7015 (N_7015,N_6512,N_6942);
nand U7016 (N_7016,N_6639,N_6995);
or U7017 (N_7017,N_6593,N_6440);
nor U7018 (N_7018,N_6744,N_6326);
or U7019 (N_7019,N_6808,N_6185);
nor U7020 (N_7020,N_6437,N_6462);
or U7021 (N_7021,N_6612,N_6299);
nor U7022 (N_7022,N_6413,N_6292);
nor U7023 (N_7023,N_6434,N_6738);
xnor U7024 (N_7024,N_6811,N_6850);
nand U7025 (N_7025,N_6445,N_6980);
xor U7026 (N_7026,N_6586,N_6684);
nor U7027 (N_7027,N_6862,N_6227);
and U7028 (N_7028,N_6160,N_6891);
nand U7029 (N_7029,N_6102,N_6943);
nor U7030 (N_7030,N_6672,N_6751);
nor U7031 (N_7031,N_6654,N_6323);
nor U7032 (N_7032,N_6762,N_6786);
xor U7033 (N_7033,N_6483,N_6514);
nor U7034 (N_7034,N_6077,N_6590);
and U7035 (N_7035,N_6468,N_6250);
or U7036 (N_7036,N_6967,N_6715);
nand U7037 (N_7037,N_6822,N_6423);
or U7038 (N_7038,N_6561,N_6547);
and U7039 (N_7039,N_6722,N_6801);
or U7040 (N_7040,N_6447,N_6741);
nand U7041 (N_7041,N_6010,N_6071);
xor U7042 (N_7042,N_6284,N_6847);
nand U7043 (N_7043,N_6795,N_6582);
xor U7044 (N_7044,N_6355,N_6490);
nand U7045 (N_7045,N_6998,N_6016);
xor U7046 (N_7046,N_6039,N_6742);
nand U7047 (N_7047,N_6719,N_6599);
nand U7048 (N_7048,N_6855,N_6930);
nor U7049 (N_7049,N_6202,N_6350);
nand U7050 (N_7050,N_6062,N_6537);
nor U7051 (N_7051,N_6119,N_6837);
or U7052 (N_7052,N_6142,N_6319);
or U7053 (N_7053,N_6321,N_6765);
and U7054 (N_7054,N_6712,N_6685);
and U7055 (N_7055,N_6024,N_6784);
nand U7056 (N_7056,N_6034,N_6579);
nand U7057 (N_7057,N_6477,N_6286);
nor U7058 (N_7058,N_6473,N_6902);
nand U7059 (N_7059,N_6376,N_6667);
nor U7060 (N_7060,N_6867,N_6369);
and U7061 (N_7061,N_6030,N_6567);
nor U7062 (N_7062,N_6615,N_6997);
and U7063 (N_7063,N_6379,N_6111);
and U7064 (N_7064,N_6670,N_6175);
xor U7065 (N_7065,N_6994,N_6732);
nand U7066 (N_7066,N_6075,N_6523);
or U7067 (N_7067,N_6475,N_6365);
nand U7068 (N_7068,N_6014,N_6373);
or U7069 (N_7069,N_6418,N_6021);
or U7070 (N_7070,N_6900,N_6086);
nor U7071 (N_7071,N_6508,N_6929);
nand U7072 (N_7072,N_6009,N_6252);
nand U7073 (N_7073,N_6770,N_6129);
or U7074 (N_7074,N_6787,N_6427);
or U7075 (N_7075,N_6398,N_6349);
nand U7076 (N_7076,N_6296,N_6311);
or U7077 (N_7077,N_6581,N_6640);
nand U7078 (N_7078,N_6216,N_6117);
nor U7079 (N_7079,N_6132,N_6450);
and U7080 (N_7080,N_6317,N_6723);
and U7081 (N_7081,N_6658,N_6970);
xnor U7082 (N_7082,N_6458,N_6033);
and U7083 (N_7083,N_6608,N_6318);
or U7084 (N_7084,N_6118,N_6446);
nand U7085 (N_7085,N_6084,N_6331);
nand U7086 (N_7086,N_6152,N_6169);
nor U7087 (N_7087,N_6294,N_6552);
xor U7088 (N_7088,N_6903,N_6168);
and U7089 (N_7089,N_6079,N_6155);
nand U7090 (N_7090,N_6573,N_6006);
and U7091 (N_7091,N_6686,N_6443);
nand U7092 (N_7092,N_6709,N_6878);
nor U7093 (N_7093,N_6148,N_6949);
nor U7094 (N_7094,N_6781,N_6767);
nand U7095 (N_7095,N_6257,N_6491);
xor U7096 (N_7096,N_6624,N_6244);
nor U7097 (N_7097,N_6176,N_6966);
xor U7098 (N_7098,N_6237,N_6826);
xnor U7099 (N_7099,N_6554,N_6282);
or U7100 (N_7100,N_6269,N_6324);
or U7101 (N_7101,N_6828,N_6865);
xor U7102 (N_7102,N_6571,N_6270);
or U7103 (N_7103,N_6213,N_6153);
nand U7104 (N_7104,N_6163,N_6652);
nor U7105 (N_7105,N_6803,N_6402);
nor U7106 (N_7106,N_6421,N_6173);
nand U7107 (N_7107,N_6546,N_6749);
nand U7108 (N_7108,N_6510,N_6184);
and U7109 (N_7109,N_6756,N_6442);
or U7110 (N_7110,N_6708,N_6619);
nand U7111 (N_7111,N_6698,N_6013);
nor U7112 (N_7112,N_6971,N_6472);
nor U7113 (N_7113,N_6578,N_6794);
nand U7114 (N_7114,N_6883,N_6978);
nor U7115 (N_7115,N_6651,N_6879);
xor U7116 (N_7116,N_6726,N_6687);
or U7117 (N_7117,N_6135,N_6604);
nor U7118 (N_7118,N_6671,N_6428);
and U7119 (N_7119,N_6236,N_6898);
xor U7120 (N_7120,N_6541,N_6931);
and U7121 (N_7121,N_6375,N_6842);
and U7122 (N_7122,N_6975,N_6591);
xor U7123 (N_7123,N_6179,N_6191);
nor U7124 (N_7124,N_6069,N_6852);
and U7125 (N_7125,N_6908,N_6342);
nand U7126 (N_7126,N_6165,N_6097);
or U7127 (N_7127,N_6154,N_6983);
and U7128 (N_7128,N_6876,N_6406);
and U7129 (N_7129,N_6381,N_6739);
and U7130 (N_7130,N_6868,N_6653);
or U7131 (N_7131,N_6088,N_6315);
xnor U7132 (N_7132,N_6981,N_6048);
xnor U7133 (N_7133,N_6948,N_6166);
and U7134 (N_7134,N_6002,N_6890);
xnor U7135 (N_7135,N_6404,N_6397);
nand U7136 (N_7136,N_6559,N_6638);
nor U7137 (N_7137,N_6478,N_6779);
nor U7138 (N_7138,N_6461,N_6258);
xnor U7139 (N_7139,N_6424,N_6938);
nand U7140 (N_7140,N_6611,N_6821);
nor U7141 (N_7141,N_6919,N_6377);
or U7142 (N_7142,N_6694,N_6729);
or U7143 (N_7143,N_6889,N_6700);
nand U7144 (N_7144,N_6977,N_6556);
xor U7145 (N_7145,N_6740,N_6587);
or U7146 (N_7146,N_6133,N_6633);
xor U7147 (N_7147,N_6809,N_6989);
xnor U7148 (N_7148,N_6449,N_6810);
nor U7149 (N_7149,N_6730,N_6410);
xor U7150 (N_7150,N_6212,N_6448);
and U7151 (N_7151,N_6368,N_6843);
and U7152 (N_7152,N_6911,N_6705);
xor U7153 (N_7153,N_6469,N_6856);
nand U7154 (N_7154,N_6772,N_6598);
xor U7155 (N_7155,N_6544,N_6594);
or U7156 (N_7156,N_6728,N_6807);
or U7157 (N_7157,N_6208,N_6157);
nor U7158 (N_7158,N_6566,N_6231);
or U7159 (N_7159,N_6841,N_6626);
or U7160 (N_7160,N_6242,N_6361);
or U7161 (N_7161,N_6961,N_6482);
nand U7162 (N_7162,N_6374,N_6226);
nor U7163 (N_7163,N_6939,N_6456);
nand U7164 (N_7164,N_6053,N_6235);
nand U7165 (N_7165,N_6812,N_6436);
nor U7166 (N_7166,N_6771,N_6993);
nor U7167 (N_7167,N_6453,N_6312);
nand U7168 (N_7168,N_6047,N_6804);
xor U7169 (N_7169,N_6695,N_6577);
nand U7170 (N_7170,N_6228,N_6589);
or U7171 (N_7171,N_6113,N_6489);
nand U7172 (N_7172,N_6710,N_6727);
and U7173 (N_7173,N_6407,N_6952);
xnor U7174 (N_7174,N_6289,N_6602);
nor U7175 (N_7175,N_6790,N_6576);
and U7176 (N_7176,N_6348,N_6764);
and U7177 (N_7177,N_6080,N_6507);
and U7178 (N_7178,N_6894,N_6699);
nor U7179 (N_7179,N_6660,N_6303);
nor U7180 (N_7180,N_6945,N_6022);
xnor U7181 (N_7181,N_6836,N_6872);
xor U7182 (N_7182,N_6569,N_6063);
nand U7183 (N_7183,N_6219,N_6390);
xnor U7184 (N_7184,N_6614,N_6799);
or U7185 (N_7185,N_6067,N_6805);
and U7186 (N_7186,N_6007,N_6542);
nor U7187 (N_7187,N_6485,N_6736);
or U7188 (N_7188,N_6217,N_6103);
and U7189 (N_7189,N_6681,N_6255);
and U7190 (N_7190,N_6545,N_6260);
or U7191 (N_7191,N_6180,N_6986);
nor U7192 (N_7192,N_6871,N_6956);
nand U7193 (N_7193,N_6613,N_6372);
and U7194 (N_7194,N_6720,N_6463);
nand U7195 (N_7195,N_6854,N_6848);
nand U7196 (N_7196,N_6702,N_6528);
nor U7197 (N_7197,N_6896,N_6240);
nand U7198 (N_7198,N_6057,N_6832);
or U7199 (N_7199,N_6074,N_6392);
xnor U7200 (N_7200,N_6106,N_6927);
nor U7201 (N_7201,N_6457,N_6099);
and U7202 (N_7202,N_6038,N_6607);
or U7203 (N_7203,N_6011,N_6680);
and U7204 (N_7204,N_6302,N_6387);
xnor U7205 (N_7205,N_6385,N_6108);
nor U7206 (N_7206,N_6470,N_6314);
nor U7207 (N_7207,N_6414,N_6497);
nor U7208 (N_7208,N_6845,N_6425);
nor U7209 (N_7209,N_6144,N_6486);
xor U7210 (N_7210,N_6109,N_6618);
xnor U7211 (N_7211,N_6636,N_6634);
xnor U7212 (N_7212,N_6935,N_6078);
and U7213 (N_7213,N_6574,N_6955);
xor U7214 (N_7214,N_6416,N_6754);
nand U7215 (N_7215,N_6954,N_6417);
nor U7216 (N_7216,N_6487,N_6743);
nor U7217 (N_7217,N_6263,N_6123);
or U7218 (N_7218,N_6422,N_6459);
xnor U7219 (N_7219,N_6584,N_6769);
and U7220 (N_7220,N_6857,N_6830);
or U7221 (N_7221,N_6580,N_6530);
xor U7222 (N_7222,N_6037,N_6277);
xnor U7223 (N_7223,N_6933,N_6238);
or U7224 (N_7224,N_6001,N_6913);
or U7225 (N_7225,N_6846,N_6182);
nand U7226 (N_7226,N_6526,N_6813);
xor U7227 (N_7227,N_6711,N_6840);
and U7228 (N_7228,N_6972,N_6110);
nand U7229 (N_7229,N_6267,N_6454);
xor U7230 (N_7230,N_6072,N_6378);
nor U7231 (N_7231,N_6521,N_6988);
nand U7232 (N_7232,N_6673,N_6924);
nand U7233 (N_7233,N_6085,N_6957);
xor U7234 (N_7234,N_6600,N_6256);
xor U7235 (N_7235,N_6595,N_6538);
or U7236 (N_7236,N_6748,N_6666);
or U7237 (N_7237,N_6172,N_6987);
nor U7238 (N_7238,N_6675,N_6543);
xnor U7239 (N_7239,N_6026,N_6439);
xor U7240 (N_7240,N_6788,N_6320);
xnor U7241 (N_7241,N_6937,N_6982);
or U7242 (N_7242,N_6094,N_6230);
xnor U7243 (N_7243,N_6713,N_6669);
and U7244 (N_7244,N_6283,N_6895);
or U7245 (N_7245,N_6901,N_6120);
nand U7246 (N_7246,N_6245,N_6689);
and U7247 (N_7247,N_6496,N_6853);
nand U7248 (N_7248,N_6800,N_6535);
xor U7249 (N_7249,N_6802,N_6115);
xnor U7250 (N_7250,N_6564,N_6218);
nor U7251 (N_7251,N_6861,N_6550);
xnor U7252 (N_7252,N_6960,N_6885);
nor U7253 (N_7253,N_6753,N_6399);
or U7254 (N_7254,N_6291,N_6341);
or U7255 (N_7255,N_6706,N_6207);
and U7256 (N_7256,N_6782,N_6015);
nor U7257 (N_7257,N_6297,N_6196);
or U7258 (N_7258,N_6540,N_6198);
or U7259 (N_7259,N_6917,N_6904);
and U7260 (N_7260,N_6204,N_6733);
or U7261 (N_7261,N_6281,N_6246);
xnor U7262 (N_7262,N_6334,N_6565);
xnor U7263 (N_7263,N_6785,N_6912);
and U7264 (N_7264,N_6363,N_6195);
xor U7265 (N_7265,N_6276,N_6310);
nand U7266 (N_7266,N_6745,N_6059);
nand U7267 (N_7267,N_6187,N_6023);
xnor U7268 (N_7268,N_6677,N_6190);
or U7269 (N_7269,N_6122,N_6386);
xor U7270 (N_7270,N_6300,N_6092);
nor U7271 (N_7271,N_6629,N_6663);
nor U7272 (N_7272,N_6683,N_6322);
xor U7273 (N_7273,N_6768,N_6553);
and U7274 (N_7274,N_6839,N_6107);
nor U7275 (N_7275,N_6357,N_6650);
and U7276 (N_7276,N_6969,N_6332);
nor U7277 (N_7277,N_6632,N_6731);
nor U7278 (N_7278,N_6337,N_6481);
nor U7279 (N_7279,N_6460,N_6431);
or U7280 (N_7280,N_6877,N_6944);
or U7281 (N_7281,N_6504,N_6290);
or U7282 (N_7282,N_6145,N_6529);
xor U7283 (N_7283,N_6147,N_6503);
nand U7284 (N_7284,N_6928,N_6548);
or U7285 (N_7285,N_6798,N_6055);
or U7286 (N_7286,N_6484,N_6206);
nor U7287 (N_7287,N_6774,N_6233);
and U7288 (N_7288,N_6985,N_6188);
or U7289 (N_7289,N_6366,N_6916);
or U7290 (N_7290,N_6575,N_6162);
nand U7291 (N_7291,N_6494,N_6274);
xor U7292 (N_7292,N_6662,N_6759);
and U7293 (N_7293,N_6882,N_6558);
nor U7294 (N_7294,N_6266,N_6620);
nand U7295 (N_7295,N_6064,N_6696);
and U7296 (N_7296,N_6158,N_6382);
and U7297 (N_7297,N_6307,N_6049);
nor U7298 (N_7298,N_6682,N_6214);
nand U7299 (N_7299,N_6346,N_6004);
nor U7300 (N_7300,N_6052,N_6513);
nand U7301 (N_7301,N_6664,N_6721);
or U7302 (N_7302,N_6171,N_6657);
nor U7303 (N_7303,N_6466,N_6305);
nor U7304 (N_7304,N_6921,N_6285);
nor U7305 (N_7305,N_6763,N_6251);
xor U7306 (N_7306,N_6833,N_6661);
and U7307 (N_7307,N_6134,N_6536);
xnor U7308 (N_7308,N_6498,N_6714);
or U7309 (N_7309,N_6444,N_6313);
nand U7310 (N_7310,N_6095,N_6465);
nand U7311 (N_7311,N_6505,N_6922);
nand U7312 (N_7312,N_6601,N_6495);
nor U7313 (N_7313,N_6716,N_6910);
nand U7314 (N_7314,N_6923,N_6345);
nor U7315 (N_7315,N_6058,N_6892);
and U7316 (N_7316,N_6426,N_6429);
and U7317 (N_7317,N_6555,N_6127);
nor U7318 (N_7318,N_6926,N_6124);
nand U7319 (N_7319,N_6051,N_6492);
or U7320 (N_7320,N_6295,N_6899);
nor U7321 (N_7321,N_6367,N_6036);
nor U7322 (N_7322,N_6958,N_6827);
nor U7323 (N_7323,N_6551,N_6356);
xor U7324 (N_7324,N_6962,N_6091);
or U7325 (N_7325,N_6441,N_6203);
and U7326 (N_7326,N_6941,N_6354);
xnor U7327 (N_7327,N_6126,N_6211);
or U7328 (N_7328,N_6792,N_6951);
nor U7329 (N_7329,N_6197,N_6973);
nand U7330 (N_7330,N_6017,N_6796);
nor U7331 (N_7331,N_6433,N_6881);
nand U7332 (N_7332,N_6806,N_6330);
nand U7333 (N_7333,N_6121,N_6934);
and U7334 (N_7334,N_6776,N_6773);
nand U7335 (N_7335,N_6241,N_6020);
or U7336 (N_7336,N_6012,N_6400);
xor U7337 (N_7337,N_6953,N_6479);
xor U7338 (N_7338,N_6760,N_6560);
xor U7339 (N_7339,N_6511,N_6897);
xor U7340 (N_7340,N_6679,N_6688);
nor U7341 (N_7341,N_6027,N_6617);
xor U7342 (N_7342,N_6524,N_6271);
nand U7343 (N_7343,N_6974,N_6616);
and U7344 (N_7344,N_6293,N_6499);
and U7345 (N_7345,N_6298,N_6050);
nor U7346 (N_7346,N_6471,N_6019);
xor U7347 (N_7347,N_6136,N_6265);
or U7348 (N_7348,N_6819,N_6520);
nor U7349 (N_7349,N_6060,N_6866);
or U7350 (N_7350,N_6534,N_6644);
or U7351 (N_7351,N_6532,N_6384);
nand U7352 (N_7352,N_6875,N_6835);
nor U7353 (N_7353,N_6880,N_6141);
xor U7354 (N_7354,N_6488,N_6452);
and U7355 (N_7355,N_6750,N_6280);
xor U7356 (N_7356,N_6412,N_6140);
or U7357 (N_7357,N_6793,N_6641);
and U7358 (N_7358,N_6333,N_6394);
xnor U7359 (N_7359,N_6339,N_6432);
xnor U7360 (N_7360,N_6186,N_6161);
xor U7361 (N_7361,N_6278,N_6411);
xnor U7362 (N_7362,N_6920,N_6347);
nor U7363 (N_7363,N_6371,N_6557);
xor U7364 (N_7364,N_6340,N_6752);
nand U7365 (N_7365,N_6874,N_6518);
xor U7366 (N_7366,N_6408,N_6419);
and U7367 (N_7367,N_6304,N_6325);
nand U7368 (N_7368,N_6335,N_6817);
nor U7369 (N_7369,N_6625,N_6222);
nor U7370 (N_7370,N_6451,N_6849);
nor U7371 (N_7371,N_6032,N_6480);
and U7372 (N_7372,N_6918,N_6150);
nand U7373 (N_7373,N_6229,N_6596);
or U7374 (N_7374,N_6151,N_6181);
nor U7375 (N_7375,N_6964,N_6914);
nand U7376 (N_7376,N_6789,N_6851);
nand U7377 (N_7377,N_6455,N_6435);
or U7378 (N_7378,N_6225,N_6525);
nor U7379 (N_7379,N_6870,N_6501);
xnor U7380 (N_7380,N_6568,N_6338);
xnor U7381 (N_7381,N_6275,N_6775);
nor U7382 (N_7382,N_6090,N_6301);
nor U7383 (N_7383,N_6081,N_6676);
nand U7384 (N_7384,N_6758,N_6844);
and U7385 (N_7385,N_6128,N_6909);
xnor U7386 (N_7386,N_6815,N_6056);
nor U7387 (N_7387,N_6192,N_6635);
or U7388 (N_7388,N_6193,N_6737);
nor U7389 (N_7389,N_6005,N_6220);
or U7390 (N_7390,N_6649,N_6308);
and U7391 (N_7391,N_6253,N_6279);
or U7392 (N_7392,N_6264,N_6003);
nor U7393 (N_7393,N_6205,N_6621);
or U7394 (N_7394,N_6655,N_6539);
nor U7395 (N_7395,N_6389,N_6288);
or U7396 (N_7396,N_6864,N_6028);
xnor U7397 (N_7397,N_6999,N_6248);
xnor U7398 (N_7398,N_6031,N_6597);
nor U7399 (N_7399,N_6201,N_6984);
xor U7400 (N_7400,N_6224,N_6637);
or U7401 (N_7401,N_6401,N_6018);
xnor U7402 (N_7402,N_6200,N_6522);
nand U7403 (N_7403,N_6096,N_6823);
or U7404 (N_7404,N_6838,N_6045);
and U7405 (N_7405,N_6701,N_6234);
nand U7406 (N_7406,N_6834,N_6221);
nor U7407 (N_7407,N_6627,N_6816);
and U7408 (N_7408,N_6370,N_6065);
xnor U7409 (N_7409,N_6415,N_6570);
and U7410 (N_7410,N_6177,N_6915);
nand U7411 (N_7411,N_6757,N_6076);
xnor U7412 (N_7412,N_6209,N_6131);
or U7413 (N_7413,N_6647,N_6380);
or U7414 (N_7414,N_6592,N_6178);
nand U7415 (N_7415,N_6143,N_6572);
nor U7416 (N_7416,N_6887,N_6362);
xor U7417 (N_7417,N_6360,N_6066);
nor U7418 (N_7418,N_6979,N_6893);
nor U7419 (N_7419,N_6606,N_6189);
and U7420 (N_7420,N_6464,N_6114);
nor U7421 (N_7421,N_6725,N_6697);
nor U7422 (N_7422,N_6438,N_6692);
and U7423 (N_7423,N_6254,N_6395);
or U7424 (N_7424,N_6690,N_6859);
xnor U7425 (N_7425,N_6605,N_6210);
and U7426 (N_7426,N_6932,N_6863);
and U7427 (N_7427,N_6884,N_6306);
nor U7428 (N_7428,N_6531,N_6474);
xnor U7429 (N_7429,N_6156,N_6358);
nor U7430 (N_7430,N_6405,N_6603);
or U7431 (N_7431,N_6035,N_6659);
or U7432 (N_7432,N_6364,N_6691);
nor U7433 (N_7433,N_6643,N_6630);
nand U7434 (N_7434,N_6873,N_6272);
nand U7435 (N_7435,N_6820,N_6139);
nor U7436 (N_7436,N_6383,N_6089);
and U7437 (N_7437,N_6351,N_6223);
or U7438 (N_7438,N_6761,N_6149);
and U7439 (N_7439,N_6533,N_6703);
or U7440 (N_7440,N_6343,N_6388);
and U7441 (N_7441,N_6583,N_6829);
or U7442 (N_7442,N_6164,N_6665);
nand U7443 (N_7443,N_6500,N_6199);
xor U7444 (N_7444,N_6467,N_6420);
or U7445 (N_7445,N_6087,N_6824);
nor U7446 (N_7446,N_6735,N_6232);
or U7447 (N_7447,N_6194,N_6755);
nor U7448 (N_7448,N_6780,N_6777);
and U7449 (N_7449,N_6327,N_6718);
nand U7450 (N_7450,N_6963,N_6734);
or U7451 (N_7451,N_6509,N_6329);
or U7452 (N_7452,N_6054,N_6082);
and U7453 (N_7453,N_6061,N_6947);
and U7454 (N_7454,N_6622,N_6858);
nor U7455 (N_7455,N_6403,N_6249);
or U7456 (N_7456,N_6527,N_6116);
or U7457 (N_7457,N_6112,N_6391);
or U7458 (N_7458,N_6646,N_6261);
nor U7459 (N_7459,N_6724,N_6515);
nand U7460 (N_7460,N_6860,N_6476);
and U7461 (N_7461,N_6287,N_6825);
nor U7462 (N_7462,N_6563,N_6628);
or U7463 (N_7463,N_6674,N_6818);
nor U7464 (N_7464,N_6992,N_6170);
or U7465 (N_7465,N_6043,N_6707);
xnor U7466 (N_7466,N_6631,N_6783);
xor U7467 (N_7467,N_6668,N_6519);
or U7468 (N_7468,N_6000,N_6101);
and U7469 (N_7469,N_6353,N_6328);
nor U7470 (N_7470,N_6093,N_6814);
xnor U7471 (N_7471,N_6409,N_6262);
or U7472 (N_7472,N_6100,N_6610);
nor U7473 (N_7473,N_6831,N_6174);
xor U7474 (N_7474,N_6273,N_6493);
xnor U7475 (N_7475,N_6396,N_6886);
and U7476 (N_7476,N_6623,N_6516);
nand U7477 (N_7477,N_6073,N_6946);
nor U7478 (N_7478,N_6159,N_6316);
or U7479 (N_7479,N_6562,N_6046);
nand U7480 (N_7480,N_6950,N_6044);
and U7481 (N_7481,N_6008,N_6025);
xor U7482 (N_7482,N_6642,N_6907);
nor U7483 (N_7483,N_6959,N_6797);
or U7484 (N_7484,N_6243,N_6906);
nand U7485 (N_7485,N_6105,N_6506);
xnor U7486 (N_7486,N_6104,N_6430);
nand U7487 (N_7487,N_6137,N_6549);
nand U7488 (N_7488,N_6336,N_6609);
nand U7489 (N_7489,N_6585,N_6344);
nor U7490 (N_7490,N_6990,N_6656);
nand U7491 (N_7491,N_6352,N_6991);
and U7492 (N_7492,N_6648,N_6678);
nor U7493 (N_7493,N_6936,N_6239);
and U7494 (N_7494,N_6645,N_6130);
xnor U7495 (N_7495,N_6040,N_6996);
xnor U7496 (N_7496,N_6704,N_6888);
or U7497 (N_7497,N_6146,N_6259);
and U7498 (N_7498,N_6393,N_6747);
xor U7499 (N_7499,N_6041,N_6517);
nor U7500 (N_7500,N_6828,N_6378);
and U7501 (N_7501,N_6402,N_6864);
nor U7502 (N_7502,N_6936,N_6613);
nand U7503 (N_7503,N_6300,N_6760);
nand U7504 (N_7504,N_6197,N_6505);
nand U7505 (N_7505,N_6225,N_6962);
or U7506 (N_7506,N_6803,N_6600);
or U7507 (N_7507,N_6370,N_6703);
nand U7508 (N_7508,N_6222,N_6722);
or U7509 (N_7509,N_6946,N_6810);
and U7510 (N_7510,N_6878,N_6198);
nand U7511 (N_7511,N_6514,N_6093);
xor U7512 (N_7512,N_6829,N_6585);
nor U7513 (N_7513,N_6317,N_6560);
or U7514 (N_7514,N_6781,N_6104);
xor U7515 (N_7515,N_6813,N_6030);
xnor U7516 (N_7516,N_6766,N_6142);
and U7517 (N_7517,N_6991,N_6329);
nor U7518 (N_7518,N_6899,N_6781);
xnor U7519 (N_7519,N_6204,N_6294);
nor U7520 (N_7520,N_6377,N_6230);
xor U7521 (N_7521,N_6149,N_6458);
nand U7522 (N_7522,N_6051,N_6461);
and U7523 (N_7523,N_6406,N_6030);
nor U7524 (N_7524,N_6139,N_6794);
and U7525 (N_7525,N_6268,N_6266);
and U7526 (N_7526,N_6091,N_6860);
nand U7527 (N_7527,N_6661,N_6359);
nor U7528 (N_7528,N_6284,N_6010);
xor U7529 (N_7529,N_6860,N_6102);
xor U7530 (N_7530,N_6817,N_6699);
and U7531 (N_7531,N_6333,N_6641);
nor U7532 (N_7532,N_6483,N_6488);
xnor U7533 (N_7533,N_6305,N_6041);
nor U7534 (N_7534,N_6864,N_6883);
or U7535 (N_7535,N_6801,N_6709);
or U7536 (N_7536,N_6636,N_6523);
nor U7537 (N_7537,N_6776,N_6574);
and U7538 (N_7538,N_6884,N_6574);
and U7539 (N_7539,N_6866,N_6919);
nand U7540 (N_7540,N_6967,N_6835);
xor U7541 (N_7541,N_6115,N_6104);
or U7542 (N_7542,N_6190,N_6104);
nand U7543 (N_7543,N_6187,N_6380);
xnor U7544 (N_7544,N_6943,N_6806);
xor U7545 (N_7545,N_6133,N_6019);
xnor U7546 (N_7546,N_6821,N_6040);
nand U7547 (N_7547,N_6512,N_6389);
xor U7548 (N_7548,N_6571,N_6392);
or U7549 (N_7549,N_6352,N_6068);
or U7550 (N_7550,N_6587,N_6530);
xnor U7551 (N_7551,N_6496,N_6742);
xnor U7552 (N_7552,N_6650,N_6904);
xnor U7553 (N_7553,N_6933,N_6642);
xor U7554 (N_7554,N_6983,N_6210);
xnor U7555 (N_7555,N_6268,N_6844);
nor U7556 (N_7556,N_6873,N_6470);
and U7557 (N_7557,N_6031,N_6281);
and U7558 (N_7558,N_6798,N_6942);
and U7559 (N_7559,N_6634,N_6708);
nor U7560 (N_7560,N_6229,N_6029);
nor U7561 (N_7561,N_6527,N_6294);
or U7562 (N_7562,N_6901,N_6644);
nand U7563 (N_7563,N_6775,N_6501);
nand U7564 (N_7564,N_6685,N_6485);
nor U7565 (N_7565,N_6056,N_6699);
or U7566 (N_7566,N_6560,N_6527);
and U7567 (N_7567,N_6636,N_6625);
xnor U7568 (N_7568,N_6720,N_6242);
xnor U7569 (N_7569,N_6573,N_6066);
nand U7570 (N_7570,N_6246,N_6433);
and U7571 (N_7571,N_6056,N_6484);
xor U7572 (N_7572,N_6548,N_6904);
nand U7573 (N_7573,N_6252,N_6506);
xnor U7574 (N_7574,N_6032,N_6845);
and U7575 (N_7575,N_6892,N_6324);
nand U7576 (N_7576,N_6377,N_6681);
or U7577 (N_7577,N_6342,N_6318);
or U7578 (N_7578,N_6462,N_6819);
nand U7579 (N_7579,N_6704,N_6863);
and U7580 (N_7580,N_6560,N_6907);
and U7581 (N_7581,N_6748,N_6893);
nor U7582 (N_7582,N_6935,N_6644);
xnor U7583 (N_7583,N_6067,N_6503);
xnor U7584 (N_7584,N_6282,N_6387);
nand U7585 (N_7585,N_6584,N_6859);
xor U7586 (N_7586,N_6621,N_6023);
or U7587 (N_7587,N_6192,N_6176);
xnor U7588 (N_7588,N_6610,N_6006);
xor U7589 (N_7589,N_6290,N_6196);
or U7590 (N_7590,N_6037,N_6835);
and U7591 (N_7591,N_6527,N_6911);
or U7592 (N_7592,N_6774,N_6584);
nand U7593 (N_7593,N_6604,N_6446);
and U7594 (N_7594,N_6728,N_6634);
nor U7595 (N_7595,N_6771,N_6905);
nand U7596 (N_7596,N_6576,N_6363);
nor U7597 (N_7597,N_6654,N_6294);
nand U7598 (N_7598,N_6463,N_6244);
nor U7599 (N_7599,N_6939,N_6755);
xor U7600 (N_7600,N_6742,N_6969);
nor U7601 (N_7601,N_6298,N_6702);
xor U7602 (N_7602,N_6471,N_6921);
nor U7603 (N_7603,N_6780,N_6968);
nand U7604 (N_7604,N_6285,N_6497);
and U7605 (N_7605,N_6627,N_6429);
xnor U7606 (N_7606,N_6359,N_6875);
nand U7607 (N_7607,N_6929,N_6423);
nand U7608 (N_7608,N_6587,N_6976);
xnor U7609 (N_7609,N_6097,N_6577);
or U7610 (N_7610,N_6627,N_6618);
and U7611 (N_7611,N_6339,N_6411);
nor U7612 (N_7612,N_6140,N_6193);
xnor U7613 (N_7613,N_6412,N_6215);
and U7614 (N_7614,N_6844,N_6335);
xor U7615 (N_7615,N_6512,N_6695);
xnor U7616 (N_7616,N_6876,N_6243);
xnor U7617 (N_7617,N_6449,N_6368);
xor U7618 (N_7618,N_6403,N_6717);
nand U7619 (N_7619,N_6160,N_6754);
nand U7620 (N_7620,N_6363,N_6517);
or U7621 (N_7621,N_6240,N_6618);
or U7622 (N_7622,N_6480,N_6735);
xor U7623 (N_7623,N_6904,N_6073);
nor U7624 (N_7624,N_6875,N_6758);
xor U7625 (N_7625,N_6181,N_6513);
and U7626 (N_7626,N_6547,N_6962);
xnor U7627 (N_7627,N_6512,N_6470);
and U7628 (N_7628,N_6786,N_6613);
or U7629 (N_7629,N_6534,N_6950);
nor U7630 (N_7630,N_6297,N_6777);
xnor U7631 (N_7631,N_6189,N_6940);
nor U7632 (N_7632,N_6093,N_6288);
or U7633 (N_7633,N_6267,N_6768);
and U7634 (N_7634,N_6341,N_6269);
xnor U7635 (N_7635,N_6335,N_6117);
or U7636 (N_7636,N_6039,N_6864);
or U7637 (N_7637,N_6308,N_6442);
or U7638 (N_7638,N_6580,N_6374);
or U7639 (N_7639,N_6089,N_6219);
and U7640 (N_7640,N_6599,N_6906);
nand U7641 (N_7641,N_6456,N_6231);
and U7642 (N_7642,N_6734,N_6731);
and U7643 (N_7643,N_6539,N_6185);
nand U7644 (N_7644,N_6493,N_6127);
xnor U7645 (N_7645,N_6225,N_6841);
and U7646 (N_7646,N_6013,N_6263);
and U7647 (N_7647,N_6123,N_6935);
or U7648 (N_7648,N_6236,N_6803);
xor U7649 (N_7649,N_6774,N_6968);
xor U7650 (N_7650,N_6266,N_6624);
xor U7651 (N_7651,N_6465,N_6957);
nor U7652 (N_7652,N_6121,N_6562);
xor U7653 (N_7653,N_6621,N_6556);
nand U7654 (N_7654,N_6318,N_6234);
nor U7655 (N_7655,N_6681,N_6776);
and U7656 (N_7656,N_6248,N_6750);
nand U7657 (N_7657,N_6956,N_6066);
and U7658 (N_7658,N_6366,N_6061);
or U7659 (N_7659,N_6043,N_6475);
and U7660 (N_7660,N_6841,N_6665);
or U7661 (N_7661,N_6823,N_6365);
nor U7662 (N_7662,N_6813,N_6017);
or U7663 (N_7663,N_6051,N_6924);
nand U7664 (N_7664,N_6828,N_6056);
nand U7665 (N_7665,N_6782,N_6771);
nor U7666 (N_7666,N_6319,N_6379);
nor U7667 (N_7667,N_6403,N_6645);
or U7668 (N_7668,N_6033,N_6698);
nor U7669 (N_7669,N_6178,N_6295);
and U7670 (N_7670,N_6537,N_6833);
xnor U7671 (N_7671,N_6181,N_6085);
xnor U7672 (N_7672,N_6449,N_6836);
and U7673 (N_7673,N_6179,N_6428);
nor U7674 (N_7674,N_6201,N_6238);
nor U7675 (N_7675,N_6320,N_6994);
xor U7676 (N_7676,N_6846,N_6826);
nand U7677 (N_7677,N_6449,N_6953);
and U7678 (N_7678,N_6963,N_6962);
xor U7679 (N_7679,N_6837,N_6780);
nor U7680 (N_7680,N_6308,N_6101);
xnor U7681 (N_7681,N_6948,N_6764);
xnor U7682 (N_7682,N_6646,N_6004);
nor U7683 (N_7683,N_6492,N_6496);
nor U7684 (N_7684,N_6224,N_6796);
xnor U7685 (N_7685,N_6961,N_6440);
or U7686 (N_7686,N_6871,N_6175);
nor U7687 (N_7687,N_6046,N_6043);
or U7688 (N_7688,N_6050,N_6951);
or U7689 (N_7689,N_6751,N_6989);
or U7690 (N_7690,N_6181,N_6063);
nor U7691 (N_7691,N_6647,N_6264);
or U7692 (N_7692,N_6232,N_6600);
nand U7693 (N_7693,N_6704,N_6322);
xor U7694 (N_7694,N_6674,N_6015);
and U7695 (N_7695,N_6790,N_6286);
nor U7696 (N_7696,N_6644,N_6324);
xor U7697 (N_7697,N_6486,N_6762);
and U7698 (N_7698,N_6885,N_6251);
and U7699 (N_7699,N_6603,N_6203);
nor U7700 (N_7700,N_6809,N_6530);
nand U7701 (N_7701,N_6792,N_6305);
nor U7702 (N_7702,N_6311,N_6039);
and U7703 (N_7703,N_6280,N_6622);
and U7704 (N_7704,N_6398,N_6775);
nand U7705 (N_7705,N_6064,N_6687);
xor U7706 (N_7706,N_6715,N_6983);
nand U7707 (N_7707,N_6467,N_6150);
xnor U7708 (N_7708,N_6195,N_6039);
xor U7709 (N_7709,N_6321,N_6528);
nand U7710 (N_7710,N_6862,N_6624);
nand U7711 (N_7711,N_6436,N_6309);
nor U7712 (N_7712,N_6504,N_6299);
nand U7713 (N_7713,N_6005,N_6343);
nor U7714 (N_7714,N_6963,N_6001);
nand U7715 (N_7715,N_6522,N_6033);
nor U7716 (N_7716,N_6534,N_6788);
nand U7717 (N_7717,N_6928,N_6811);
nor U7718 (N_7718,N_6185,N_6430);
nor U7719 (N_7719,N_6044,N_6552);
xor U7720 (N_7720,N_6372,N_6144);
xnor U7721 (N_7721,N_6869,N_6115);
nand U7722 (N_7722,N_6754,N_6963);
nand U7723 (N_7723,N_6749,N_6751);
nand U7724 (N_7724,N_6986,N_6953);
and U7725 (N_7725,N_6408,N_6997);
nor U7726 (N_7726,N_6113,N_6512);
or U7727 (N_7727,N_6189,N_6241);
and U7728 (N_7728,N_6297,N_6830);
nor U7729 (N_7729,N_6630,N_6648);
nand U7730 (N_7730,N_6671,N_6002);
xnor U7731 (N_7731,N_6206,N_6683);
and U7732 (N_7732,N_6304,N_6822);
xor U7733 (N_7733,N_6106,N_6084);
xor U7734 (N_7734,N_6532,N_6047);
or U7735 (N_7735,N_6965,N_6197);
nand U7736 (N_7736,N_6455,N_6605);
nand U7737 (N_7737,N_6659,N_6924);
nand U7738 (N_7738,N_6865,N_6117);
xnor U7739 (N_7739,N_6881,N_6856);
or U7740 (N_7740,N_6533,N_6523);
xor U7741 (N_7741,N_6779,N_6714);
xnor U7742 (N_7742,N_6538,N_6241);
and U7743 (N_7743,N_6106,N_6048);
xor U7744 (N_7744,N_6201,N_6329);
and U7745 (N_7745,N_6270,N_6442);
nor U7746 (N_7746,N_6121,N_6900);
or U7747 (N_7747,N_6421,N_6032);
or U7748 (N_7748,N_6240,N_6766);
nor U7749 (N_7749,N_6109,N_6541);
xor U7750 (N_7750,N_6229,N_6239);
xor U7751 (N_7751,N_6072,N_6619);
or U7752 (N_7752,N_6862,N_6870);
xnor U7753 (N_7753,N_6398,N_6742);
nor U7754 (N_7754,N_6975,N_6684);
and U7755 (N_7755,N_6390,N_6751);
nor U7756 (N_7756,N_6113,N_6106);
nand U7757 (N_7757,N_6288,N_6596);
xor U7758 (N_7758,N_6670,N_6696);
nor U7759 (N_7759,N_6340,N_6794);
nor U7760 (N_7760,N_6731,N_6170);
or U7761 (N_7761,N_6989,N_6818);
and U7762 (N_7762,N_6809,N_6900);
nor U7763 (N_7763,N_6733,N_6606);
and U7764 (N_7764,N_6372,N_6193);
xor U7765 (N_7765,N_6234,N_6340);
nand U7766 (N_7766,N_6622,N_6398);
nor U7767 (N_7767,N_6009,N_6925);
or U7768 (N_7768,N_6766,N_6023);
xnor U7769 (N_7769,N_6667,N_6069);
nor U7770 (N_7770,N_6507,N_6569);
xnor U7771 (N_7771,N_6323,N_6601);
xor U7772 (N_7772,N_6650,N_6514);
nand U7773 (N_7773,N_6651,N_6769);
and U7774 (N_7774,N_6570,N_6912);
xor U7775 (N_7775,N_6814,N_6770);
xor U7776 (N_7776,N_6933,N_6343);
or U7777 (N_7777,N_6368,N_6539);
xnor U7778 (N_7778,N_6505,N_6119);
and U7779 (N_7779,N_6531,N_6512);
nand U7780 (N_7780,N_6470,N_6025);
xnor U7781 (N_7781,N_6029,N_6806);
nor U7782 (N_7782,N_6657,N_6080);
or U7783 (N_7783,N_6225,N_6952);
nand U7784 (N_7784,N_6691,N_6102);
and U7785 (N_7785,N_6207,N_6469);
or U7786 (N_7786,N_6812,N_6125);
and U7787 (N_7787,N_6381,N_6294);
and U7788 (N_7788,N_6343,N_6265);
and U7789 (N_7789,N_6195,N_6520);
nand U7790 (N_7790,N_6499,N_6990);
or U7791 (N_7791,N_6096,N_6359);
or U7792 (N_7792,N_6272,N_6196);
xnor U7793 (N_7793,N_6934,N_6848);
and U7794 (N_7794,N_6874,N_6909);
and U7795 (N_7795,N_6755,N_6125);
nand U7796 (N_7796,N_6425,N_6860);
xnor U7797 (N_7797,N_6775,N_6808);
nand U7798 (N_7798,N_6048,N_6627);
or U7799 (N_7799,N_6068,N_6821);
xnor U7800 (N_7800,N_6459,N_6482);
xor U7801 (N_7801,N_6418,N_6317);
nand U7802 (N_7802,N_6212,N_6138);
or U7803 (N_7803,N_6040,N_6427);
or U7804 (N_7804,N_6700,N_6691);
and U7805 (N_7805,N_6100,N_6399);
and U7806 (N_7806,N_6581,N_6754);
xnor U7807 (N_7807,N_6834,N_6611);
and U7808 (N_7808,N_6181,N_6923);
nand U7809 (N_7809,N_6558,N_6959);
and U7810 (N_7810,N_6157,N_6756);
nand U7811 (N_7811,N_6614,N_6260);
or U7812 (N_7812,N_6266,N_6586);
xnor U7813 (N_7813,N_6047,N_6498);
and U7814 (N_7814,N_6033,N_6928);
and U7815 (N_7815,N_6393,N_6377);
xnor U7816 (N_7816,N_6666,N_6526);
nand U7817 (N_7817,N_6663,N_6703);
or U7818 (N_7818,N_6546,N_6369);
or U7819 (N_7819,N_6598,N_6634);
nand U7820 (N_7820,N_6303,N_6593);
and U7821 (N_7821,N_6238,N_6532);
or U7822 (N_7822,N_6797,N_6282);
nand U7823 (N_7823,N_6655,N_6186);
nor U7824 (N_7824,N_6290,N_6926);
and U7825 (N_7825,N_6837,N_6659);
xor U7826 (N_7826,N_6315,N_6693);
and U7827 (N_7827,N_6422,N_6792);
or U7828 (N_7828,N_6183,N_6561);
nand U7829 (N_7829,N_6935,N_6224);
and U7830 (N_7830,N_6350,N_6851);
nand U7831 (N_7831,N_6806,N_6363);
nor U7832 (N_7832,N_6286,N_6053);
and U7833 (N_7833,N_6232,N_6058);
and U7834 (N_7834,N_6360,N_6889);
nand U7835 (N_7835,N_6908,N_6562);
and U7836 (N_7836,N_6652,N_6255);
nor U7837 (N_7837,N_6158,N_6786);
nor U7838 (N_7838,N_6279,N_6651);
nand U7839 (N_7839,N_6606,N_6541);
or U7840 (N_7840,N_6056,N_6186);
or U7841 (N_7841,N_6419,N_6611);
nor U7842 (N_7842,N_6128,N_6476);
xnor U7843 (N_7843,N_6459,N_6211);
nand U7844 (N_7844,N_6591,N_6127);
or U7845 (N_7845,N_6711,N_6886);
nand U7846 (N_7846,N_6371,N_6526);
nor U7847 (N_7847,N_6013,N_6966);
or U7848 (N_7848,N_6448,N_6269);
xnor U7849 (N_7849,N_6551,N_6147);
and U7850 (N_7850,N_6854,N_6514);
nor U7851 (N_7851,N_6548,N_6408);
or U7852 (N_7852,N_6391,N_6440);
xor U7853 (N_7853,N_6686,N_6607);
nor U7854 (N_7854,N_6456,N_6177);
and U7855 (N_7855,N_6974,N_6298);
or U7856 (N_7856,N_6774,N_6800);
and U7857 (N_7857,N_6140,N_6877);
nor U7858 (N_7858,N_6748,N_6177);
xor U7859 (N_7859,N_6255,N_6537);
and U7860 (N_7860,N_6673,N_6741);
and U7861 (N_7861,N_6824,N_6914);
and U7862 (N_7862,N_6196,N_6210);
and U7863 (N_7863,N_6549,N_6821);
or U7864 (N_7864,N_6132,N_6193);
xor U7865 (N_7865,N_6029,N_6589);
xnor U7866 (N_7866,N_6211,N_6637);
nor U7867 (N_7867,N_6170,N_6321);
nor U7868 (N_7868,N_6686,N_6659);
xor U7869 (N_7869,N_6978,N_6565);
nor U7870 (N_7870,N_6025,N_6614);
or U7871 (N_7871,N_6313,N_6412);
nand U7872 (N_7872,N_6515,N_6625);
nand U7873 (N_7873,N_6898,N_6764);
nor U7874 (N_7874,N_6168,N_6329);
nor U7875 (N_7875,N_6017,N_6011);
or U7876 (N_7876,N_6779,N_6094);
nor U7877 (N_7877,N_6559,N_6676);
xor U7878 (N_7878,N_6492,N_6843);
nand U7879 (N_7879,N_6299,N_6152);
nor U7880 (N_7880,N_6512,N_6433);
nor U7881 (N_7881,N_6816,N_6776);
nand U7882 (N_7882,N_6078,N_6324);
nand U7883 (N_7883,N_6123,N_6743);
xor U7884 (N_7884,N_6625,N_6423);
nor U7885 (N_7885,N_6831,N_6786);
nand U7886 (N_7886,N_6161,N_6850);
nand U7887 (N_7887,N_6059,N_6853);
xnor U7888 (N_7888,N_6743,N_6710);
and U7889 (N_7889,N_6092,N_6469);
nor U7890 (N_7890,N_6484,N_6086);
xnor U7891 (N_7891,N_6595,N_6988);
xor U7892 (N_7892,N_6532,N_6852);
and U7893 (N_7893,N_6145,N_6296);
nor U7894 (N_7894,N_6149,N_6099);
nand U7895 (N_7895,N_6859,N_6611);
and U7896 (N_7896,N_6376,N_6691);
nand U7897 (N_7897,N_6963,N_6434);
nand U7898 (N_7898,N_6915,N_6030);
nand U7899 (N_7899,N_6843,N_6006);
xnor U7900 (N_7900,N_6927,N_6489);
nor U7901 (N_7901,N_6217,N_6500);
xor U7902 (N_7902,N_6091,N_6582);
nor U7903 (N_7903,N_6521,N_6600);
nand U7904 (N_7904,N_6067,N_6183);
nand U7905 (N_7905,N_6064,N_6029);
nand U7906 (N_7906,N_6489,N_6332);
nor U7907 (N_7907,N_6521,N_6382);
xor U7908 (N_7908,N_6263,N_6265);
nor U7909 (N_7909,N_6231,N_6984);
or U7910 (N_7910,N_6756,N_6193);
xor U7911 (N_7911,N_6932,N_6755);
xor U7912 (N_7912,N_6438,N_6681);
nor U7913 (N_7913,N_6231,N_6911);
xnor U7914 (N_7914,N_6413,N_6416);
xor U7915 (N_7915,N_6549,N_6130);
nand U7916 (N_7916,N_6382,N_6862);
nand U7917 (N_7917,N_6397,N_6527);
nor U7918 (N_7918,N_6316,N_6662);
and U7919 (N_7919,N_6589,N_6778);
or U7920 (N_7920,N_6297,N_6991);
nand U7921 (N_7921,N_6423,N_6116);
xnor U7922 (N_7922,N_6167,N_6306);
nand U7923 (N_7923,N_6207,N_6523);
and U7924 (N_7924,N_6289,N_6803);
or U7925 (N_7925,N_6668,N_6901);
nor U7926 (N_7926,N_6169,N_6704);
xor U7927 (N_7927,N_6491,N_6074);
or U7928 (N_7928,N_6924,N_6126);
or U7929 (N_7929,N_6103,N_6139);
nand U7930 (N_7930,N_6270,N_6880);
nor U7931 (N_7931,N_6359,N_6403);
nor U7932 (N_7932,N_6904,N_6538);
or U7933 (N_7933,N_6912,N_6825);
nand U7934 (N_7934,N_6071,N_6448);
nand U7935 (N_7935,N_6822,N_6454);
and U7936 (N_7936,N_6688,N_6101);
xor U7937 (N_7937,N_6974,N_6776);
nand U7938 (N_7938,N_6353,N_6337);
nor U7939 (N_7939,N_6207,N_6883);
or U7940 (N_7940,N_6244,N_6075);
or U7941 (N_7941,N_6768,N_6192);
and U7942 (N_7942,N_6504,N_6901);
nand U7943 (N_7943,N_6861,N_6925);
or U7944 (N_7944,N_6643,N_6584);
nor U7945 (N_7945,N_6914,N_6101);
nor U7946 (N_7946,N_6874,N_6939);
or U7947 (N_7947,N_6924,N_6716);
xor U7948 (N_7948,N_6347,N_6338);
nor U7949 (N_7949,N_6723,N_6965);
or U7950 (N_7950,N_6278,N_6817);
nand U7951 (N_7951,N_6125,N_6168);
nor U7952 (N_7952,N_6268,N_6807);
nor U7953 (N_7953,N_6996,N_6437);
nor U7954 (N_7954,N_6223,N_6175);
and U7955 (N_7955,N_6336,N_6927);
nor U7956 (N_7956,N_6662,N_6911);
or U7957 (N_7957,N_6016,N_6669);
or U7958 (N_7958,N_6204,N_6050);
and U7959 (N_7959,N_6401,N_6488);
and U7960 (N_7960,N_6985,N_6631);
nor U7961 (N_7961,N_6149,N_6434);
nor U7962 (N_7962,N_6492,N_6331);
xnor U7963 (N_7963,N_6200,N_6774);
and U7964 (N_7964,N_6740,N_6309);
xor U7965 (N_7965,N_6635,N_6691);
or U7966 (N_7966,N_6110,N_6487);
and U7967 (N_7967,N_6748,N_6079);
and U7968 (N_7968,N_6891,N_6134);
or U7969 (N_7969,N_6706,N_6080);
nor U7970 (N_7970,N_6597,N_6180);
xor U7971 (N_7971,N_6155,N_6623);
and U7972 (N_7972,N_6260,N_6169);
nand U7973 (N_7973,N_6924,N_6481);
xor U7974 (N_7974,N_6382,N_6114);
nand U7975 (N_7975,N_6202,N_6544);
xnor U7976 (N_7976,N_6416,N_6408);
nor U7977 (N_7977,N_6282,N_6521);
nand U7978 (N_7978,N_6675,N_6876);
nor U7979 (N_7979,N_6498,N_6392);
or U7980 (N_7980,N_6248,N_6139);
and U7981 (N_7981,N_6585,N_6026);
and U7982 (N_7982,N_6670,N_6949);
nor U7983 (N_7983,N_6767,N_6297);
xnor U7984 (N_7984,N_6440,N_6142);
and U7985 (N_7985,N_6043,N_6184);
and U7986 (N_7986,N_6981,N_6498);
and U7987 (N_7987,N_6199,N_6440);
or U7988 (N_7988,N_6030,N_6699);
xnor U7989 (N_7989,N_6192,N_6366);
xor U7990 (N_7990,N_6730,N_6799);
xor U7991 (N_7991,N_6187,N_6111);
and U7992 (N_7992,N_6858,N_6235);
xor U7993 (N_7993,N_6086,N_6076);
or U7994 (N_7994,N_6131,N_6311);
and U7995 (N_7995,N_6097,N_6698);
and U7996 (N_7996,N_6106,N_6808);
xor U7997 (N_7997,N_6994,N_6568);
and U7998 (N_7998,N_6317,N_6287);
nor U7999 (N_7999,N_6413,N_6032);
or U8000 (N_8000,N_7218,N_7639);
nor U8001 (N_8001,N_7907,N_7585);
nand U8002 (N_8002,N_7875,N_7988);
nand U8003 (N_8003,N_7860,N_7443);
or U8004 (N_8004,N_7305,N_7631);
nor U8005 (N_8005,N_7161,N_7086);
nor U8006 (N_8006,N_7844,N_7427);
and U8007 (N_8007,N_7945,N_7145);
or U8008 (N_8008,N_7455,N_7377);
nor U8009 (N_8009,N_7966,N_7887);
xnor U8010 (N_8010,N_7210,N_7211);
nor U8011 (N_8011,N_7622,N_7714);
or U8012 (N_8012,N_7277,N_7140);
nand U8013 (N_8013,N_7178,N_7496);
nor U8014 (N_8014,N_7510,N_7659);
nor U8015 (N_8015,N_7785,N_7416);
and U8016 (N_8016,N_7334,N_7570);
and U8017 (N_8017,N_7062,N_7414);
nand U8018 (N_8018,N_7101,N_7647);
nor U8019 (N_8019,N_7621,N_7993);
or U8020 (N_8020,N_7963,N_7445);
or U8021 (N_8021,N_7095,N_7671);
xnor U8022 (N_8022,N_7578,N_7012);
nand U8023 (N_8023,N_7971,N_7944);
xnor U8024 (N_8024,N_7475,N_7319);
or U8025 (N_8025,N_7358,N_7855);
nand U8026 (N_8026,N_7282,N_7630);
nor U8027 (N_8027,N_7538,N_7839);
and U8028 (N_8028,N_7782,N_7953);
and U8029 (N_8029,N_7199,N_7330);
xor U8030 (N_8030,N_7060,N_7940);
xnor U8031 (N_8031,N_7991,N_7428);
or U8032 (N_8032,N_7473,N_7852);
or U8033 (N_8033,N_7515,N_7661);
and U8034 (N_8034,N_7776,N_7133);
nor U8035 (N_8035,N_7636,N_7359);
and U8036 (N_8036,N_7504,N_7200);
xnor U8037 (N_8037,N_7118,N_7582);
or U8038 (N_8038,N_7307,N_7077);
nand U8039 (N_8039,N_7000,N_7741);
nor U8040 (N_8040,N_7650,N_7353);
and U8041 (N_8041,N_7460,N_7057);
nor U8042 (N_8042,N_7204,N_7419);
nand U8043 (N_8043,N_7237,N_7586);
or U8044 (N_8044,N_7895,N_7928);
nand U8045 (N_8045,N_7613,N_7084);
or U8046 (N_8046,N_7503,N_7157);
nand U8047 (N_8047,N_7398,N_7828);
or U8048 (N_8048,N_7891,N_7010);
or U8049 (N_8049,N_7616,N_7092);
and U8050 (N_8050,N_7535,N_7313);
xor U8051 (N_8051,N_7122,N_7581);
nand U8052 (N_8052,N_7138,N_7555);
xor U8053 (N_8053,N_7765,N_7451);
xnor U8054 (N_8054,N_7853,N_7790);
nand U8055 (N_8055,N_7041,N_7549);
nand U8056 (N_8056,N_7556,N_7863);
or U8057 (N_8057,N_7242,N_7034);
nor U8058 (N_8058,N_7873,N_7320);
and U8059 (N_8059,N_7097,N_7684);
or U8060 (N_8060,N_7514,N_7896);
and U8061 (N_8061,N_7685,N_7634);
or U8062 (N_8062,N_7625,N_7109);
xnor U8063 (N_8063,N_7415,N_7640);
nor U8064 (N_8064,N_7547,N_7546);
or U8065 (N_8065,N_7395,N_7673);
xor U8066 (N_8066,N_7396,N_7185);
or U8067 (N_8067,N_7656,N_7151);
nor U8068 (N_8068,N_7219,N_7899);
and U8069 (N_8069,N_7332,N_7522);
nand U8070 (N_8070,N_7708,N_7882);
nand U8071 (N_8071,N_7106,N_7879);
or U8072 (N_8072,N_7754,N_7272);
nand U8073 (N_8073,N_7830,N_7652);
xnor U8074 (N_8074,N_7850,N_7354);
nand U8075 (N_8075,N_7175,N_7123);
or U8076 (N_8076,N_7584,N_7566);
and U8077 (N_8077,N_7864,N_7926);
xnor U8078 (N_8078,N_7382,N_7847);
xnor U8079 (N_8079,N_7069,N_7781);
nor U8080 (N_8080,N_7369,N_7375);
nand U8081 (N_8081,N_7087,N_7252);
or U8082 (N_8082,N_7187,N_7543);
xor U8083 (N_8083,N_7311,N_7271);
nor U8084 (N_8084,N_7227,N_7592);
nor U8085 (N_8085,N_7892,N_7615);
xnor U8086 (N_8086,N_7324,N_7935);
nand U8087 (N_8087,N_7308,N_7479);
and U8088 (N_8088,N_7399,N_7737);
and U8089 (N_8089,N_7540,N_7082);
or U8090 (N_8090,N_7653,N_7164);
and U8091 (N_8091,N_7858,N_7348);
or U8092 (N_8092,N_7816,N_7246);
or U8093 (N_8093,N_7572,N_7417);
nand U8094 (N_8094,N_7264,N_7600);
xor U8095 (N_8095,N_7552,N_7391);
and U8096 (N_8096,N_7142,N_7498);
nand U8097 (N_8097,N_7778,N_7179);
nor U8098 (N_8098,N_7598,N_7405);
xor U8099 (N_8099,N_7948,N_7280);
or U8100 (N_8100,N_7511,N_7247);
xor U8101 (N_8101,N_7147,N_7682);
or U8102 (N_8102,N_7126,N_7134);
nor U8103 (N_8103,N_7036,N_7927);
xor U8104 (N_8104,N_7638,N_7571);
or U8105 (N_8105,N_7533,N_7728);
and U8106 (N_8106,N_7904,N_7031);
and U8107 (N_8107,N_7667,N_7901);
xor U8108 (N_8108,N_7569,N_7002);
or U8109 (N_8109,N_7564,N_7772);
or U8110 (N_8110,N_7253,N_7591);
nor U8111 (N_8111,N_7005,N_7422);
and U8112 (N_8112,N_7787,N_7788);
and U8113 (N_8113,N_7693,N_7325);
nand U8114 (N_8114,N_7658,N_7426);
nor U8115 (N_8115,N_7825,N_7418);
and U8116 (N_8116,N_7646,N_7085);
nor U8117 (N_8117,N_7183,N_7703);
or U8118 (N_8118,N_7394,N_7180);
xnor U8119 (N_8119,N_7628,N_7287);
or U8120 (N_8120,N_7799,N_7937);
nor U8121 (N_8121,N_7442,N_7339);
or U8122 (N_8122,N_7822,N_7029);
or U8123 (N_8123,N_7736,N_7516);
and U8124 (N_8124,N_7859,N_7038);
nand U8125 (N_8125,N_7681,N_7470);
nor U8126 (N_8126,N_7297,N_7701);
xnor U8127 (N_8127,N_7824,N_7017);
xnor U8128 (N_8128,N_7477,N_7314);
nand U8129 (N_8129,N_7385,N_7420);
xor U8130 (N_8130,N_7491,N_7662);
xor U8131 (N_8131,N_7088,N_7248);
and U8132 (N_8132,N_7286,N_7517);
xor U8133 (N_8133,N_7360,N_7832);
or U8134 (N_8134,N_7722,N_7367);
or U8135 (N_8135,N_7996,N_7649);
nand U8136 (N_8136,N_7763,N_7411);
or U8137 (N_8137,N_7440,N_7645);
nor U8138 (N_8138,N_7257,N_7866);
xor U8139 (N_8139,N_7119,N_7501);
nand U8140 (N_8140,N_7058,N_7458);
and U8141 (N_8141,N_7072,N_7651);
and U8142 (N_8142,N_7750,N_7743);
nor U8143 (N_8143,N_7273,N_7212);
and U8144 (N_8144,N_7296,N_7934);
and U8145 (N_8145,N_7129,N_7453);
and U8146 (N_8146,N_7090,N_7762);
or U8147 (N_8147,N_7910,N_7141);
xor U8148 (N_8148,N_7430,N_7346);
nor U8149 (N_8149,N_7826,N_7979);
xor U8150 (N_8150,N_7527,N_7465);
nand U8151 (N_8151,N_7006,N_7176);
nor U8152 (N_8152,N_7235,N_7529);
nand U8153 (N_8153,N_7042,N_7435);
xnor U8154 (N_8154,N_7506,N_7654);
or U8155 (N_8155,N_7502,N_7323);
and U8156 (N_8156,N_7663,N_7987);
xnor U8157 (N_8157,N_7223,N_7489);
nor U8158 (N_8158,N_7956,N_7292);
xnor U8159 (N_8159,N_7403,N_7810);
or U8160 (N_8160,N_7102,N_7194);
nand U8161 (N_8161,N_7055,N_7793);
or U8162 (N_8162,N_7507,N_7773);
nand U8163 (N_8163,N_7691,N_7734);
and U8164 (N_8164,N_7168,N_7263);
and U8165 (N_8165,N_7051,N_7486);
xor U8166 (N_8166,N_7366,N_7376);
and U8167 (N_8167,N_7897,N_7717);
nand U8168 (N_8168,N_7744,N_7982);
or U8169 (N_8169,N_7441,N_7021);
xnor U8170 (N_8170,N_7677,N_7689);
nand U8171 (N_8171,N_7694,N_7946);
or U8172 (N_8172,N_7929,N_7295);
nand U8173 (N_8173,N_7597,N_7885);
nand U8174 (N_8174,N_7124,N_7712);
or U8175 (N_8175,N_7814,N_7047);
xor U8176 (N_8176,N_7488,N_7160);
xnor U8177 (N_8177,N_7152,N_7229);
or U8178 (N_8178,N_7939,N_7545);
nand U8179 (N_8179,N_7550,N_7534);
and U8180 (N_8180,N_7997,N_7833);
nand U8181 (N_8181,N_7789,N_7846);
nor U8182 (N_8182,N_7687,N_7742);
or U8183 (N_8183,N_7715,N_7867);
and U8184 (N_8184,N_7672,N_7579);
nand U8185 (N_8185,N_7393,N_7089);
xnor U8186 (N_8186,N_7181,N_7849);
xor U8187 (N_8187,N_7880,N_7177);
nor U8188 (N_8188,N_7955,N_7144);
nand U8189 (N_8189,N_7642,N_7719);
nor U8190 (N_8190,N_7240,N_7462);
xor U8191 (N_8191,N_7232,N_7521);
or U8192 (N_8192,N_7513,N_7356);
or U8193 (N_8193,N_7562,N_7484);
and U8194 (N_8194,N_7196,N_7052);
and U8195 (N_8195,N_7525,N_7698);
or U8196 (N_8196,N_7125,N_7224);
nor U8197 (N_8197,N_7054,N_7463);
nand U8198 (N_8198,N_7329,N_7884);
or U8199 (N_8199,N_7723,N_7143);
nand U8200 (N_8200,N_7070,N_7355);
xnor U8201 (N_8201,N_7753,N_7542);
xor U8202 (N_8202,N_7039,N_7664);
nor U8203 (N_8203,N_7675,N_7401);
and U8204 (N_8204,N_7048,N_7641);
and U8205 (N_8205,N_7374,N_7217);
or U8206 (N_8206,N_7947,N_7795);
and U8207 (N_8207,N_7568,N_7009);
or U8208 (N_8208,N_7267,N_7942);
nor U8209 (N_8209,N_7528,N_7384);
xnor U8210 (N_8210,N_7096,N_7819);
and U8211 (N_8211,N_7265,N_7446);
nor U8212 (N_8212,N_7167,N_7322);
or U8213 (N_8213,N_7372,N_7472);
or U8214 (N_8214,N_7611,N_7811);
xnor U8215 (N_8215,N_7439,N_7027);
or U8216 (N_8216,N_7238,N_7886);
xor U8217 (N_8217,N_7033,N_7025);
and U8218 (N_8218,N_7509,N_7373);
xor U8219 (N_8219,N_7831,N_7107);
xor U8220 (N_8220,N_7081,N_7764);
nand U8221 (N_8221,N_7854,N_7350);
or U8222 (N_8222,N_7409,N_7759);
or U8223 (N_8223,N_7024,N_7362);
xnor U8224 (N_8224,N_7720,N_7718);
and U8225 (N_8225,N_7862,N_7871);
nand U8226 (N_8226,N_7068,N_7397);
xor U8227 (N_8227,N_7075,N_7104);
nand U8228 (N_8228,N_7965,N_7735);
and U8229 (N_8229,N_7908,N_7061);
and U8230 (N_8230,N_7154,N_7679);
xnor U8231 (N_8231,N_7577,N_7222);
xnor U8232 (N_8232,N_7558,N_7207);
nand U8233 (N_8233,N_7467,N_7407);
and U8234 (N_8234,N_7303,N_7284);
or U8235 (N_8235,N_7665,N_7894);
nand U8236 (N_8236,N_7328,N_7318);
or U8237 (N_8237,N_7040,N_7030);
xnor U8238 (N_8238,N_7551,N_7083);
nand U8239 (N_8239,N_7756,N_7471);
nand U8240 (N_8240,N_7537,N_7829);
and U8241 (N_8241,N_7730,N_7733);
and U8242 (N_8242,N_7791,N_7392);
or U8243 (N_8243,N_7575,N_7711);
or U8244 (N_8244,N_7158,N_7783);
and U8245 (N_8245,N_7244,N_7881);
or U8246 (N_8246,N_7189,N_7576);
or U8247 (N_8247,N_7333,N_7293);
nand U8248 (N_8248,N_7281,N_7236);
and U8249 (N_8249,N_7792,N_7842);
nor U8250 (N_8250,N_7950,N_7343);
or U8251 (N_8251,N_7526,N_7697);
xor U8252 (N_8252,N_7580,N_7310);
and U8253 (N_8253,N_7784,N_7163);
xor U8254 (N_8254,N_7105,N_7215);
xor U8255 (N_8255,N_7259,N_7678);
nor U8256 (N_8256,N_7091,N_7856);
xor U8257 (N_8257,N_7802,N_7388);
nor U8258 (N_8258,N_7868,N_7053);
and U8259 (N_8259,N_7958,N_7952);
xor U8260 (N_8260,N_7113,N_7056);
xnor U8261 (N_8261,N_7593,N_7596);
xnor U8262 (N_8262,N_7905,N_7923);
and U8263 (N_8263,N_7174,N_7595);
and U8264 (N_8264,N_7796,N_7890);
nor U8265 (N_8265,N_7028,N_7813);
nand U8266 (N_8266,N_7379,N_7561);
nand U8267 (N_8267,N_7695,N_7476);
and U8268 (N_8268,N_7941,N_7389);
nand U8269 (N_8269,N_7524,N_7120);
and U8270 (N_8270,N_7370,N_7459);
nor U8271 (N_8271,N_7383,N_7618);
xor U8272 (N_8272,N_7794,N_7548);
xor U8273 (N_8273,N_7962,N_7699);
and U8274 (N_8274,N_7452,N_7268);
and U8275 (N_8275,N_7874,N_7380);
nor U8276 (N_8276,N_7003,N_7022);
nand U8277 (N_8277,N_7637,N_7827);
or U8278 (N_8278,N_7780,N_7182);
nor U8279 (N_8279,N_7726,N_7877);
nand U8280 (N_8280,N_7721,N_7933);
nor U8281 (N_8281,N_7239,N_7774);
nand U8282 (N_8282,N_7450,N_7925);
xnor U8283 (N_8283,N_7469,N_7220);
nor U8284 (N_8284,N_7078,N_7171);
xnor U8285 (N_8285,N_7197,N_7706);
or U8286 (N_8286,N_7688,N_7841);
or U8287 (N_8287,N_7869,N_7657);
and U8288 (N_8288,N_7834,N_7992);
and U8289 (N_8289,N_7977,N_7755);
or U8290 (N_8290,N_7709,N_7713);
or U8291 (N_8291,N_7587,N_7387);
nor U8292 (N_8292,N_7285,N_7567);
and U8293 (N_8293,N_7740,N_7690);
nor U8294 (N_8294,N_7225,N_7255);
or U8295 (N_8295,N_7099,N_7902);
and U8296 (N_8296,N_7249,N_7306);
or U8297 (N_8297,N_7400,N_7609);
and U8298 (N_8298,N_7602,N_7302);
nand U8299 (N_8299,N_7076,N_7127);
xnor U8300 (N_8300,N_7512,N_7206);
nor U8301 (N_8301,N_7378,N_7233);
xnor U8302 (N_8302,N_7447,N_7195);
xnor U8303 (N_8303,N_7975,N_7998);
or U8304 (N_8304,N_7132,N_7406);
nor U8305 (N_8305,N_7767,N_7800);
nand U8306 (N_8306,N_7186,N_7606);
nor U8307 (N_8307,N_7505,N_7725);
and U8308 (N_8308,N_7610,N_7063);
or U8309 (N_8309,N_7114,N_7191);
nand U8310 (N_8310,N_7312,N_7234);
and U8311 (N_8311,N_7539,N_7363);
or U8312 (N_8312,N_7492,N_7920);
xor U8313 (N_8313,N_7497,N_7903);
xnor U8314 (N_8314,N_7412,N_7961);
xor U8315 (N_8315,N_7316,N_7974);
and U8316 (N_8316,N_7779,N_7617);
and U8317 (N_8317,N_7130,N_7909);
and U8318 (N_8318,N_7251,N_7648);
xor U8319 (N_8319,N_7423,N_7433);
or U8320 (N_8320,N_7523,N_7071);
nor U8321 (N_8321,N_7770,N_7074);
xnor U8322 (N_8322,N_7331,N_7110);
nor U8323 (N_8323,N_7739,N_7761);
nand U8324 (N_8324,N_7241,N_7337);
xor U8325 (N_8325,N_7007,N_7635);
xor U8326 (N_8326,N_7932,N_7913);
or U8327 (N_8327,N_7976,N_7806);
nand U8328 (N_8328,N_7013,N_7843);
and U8329 (N_8329,N_7632,N_7804);
and U8330 (N_8330,N_7483,N_7493);
nor U8331 (N_8331,N_7301,N_7456);
xor U8332 (N_8332,N_7898,N_7900);
xnor U8333 (N_8333,N_7261,N_7731);
xor U8334 (N_8334,N_7914,N_7468);
and U8335 (N_8335,N_7751,N_7188);
nor U8336 (N_8336,N_7357,N_7845);
or U8337 (N_8337,N_7768,N_7589);
xor U8338 (N_8338,N_7044,N_7565);
and U8339 (N_8339,N_7413,N_7985);
and U8340 (N_8340,N_7590,N_7404);
nand U8341 (N_8341,N_7482,N_7098);
nor U8342 (N_8342,N_7912,N_7727);
or U8343 (N_8343,N_7531,N_7250);
and U8344 (N_8344,N_7274,N_7915);
xnor U8345 (N_8345,N_7760,N_7386);
nand U8346 (N_8346,N_7588,N_7878);
nor U8347 (N_8347,N_7049,N_7438);
and U8348 (N_8348,N_7990,N_7254);
xor U8349 (N_8349,N_7173,N_7969);
and U8350 (N_8350,N_7162,N_7605);
nor U8351 (N_8351,N_7437,N_7115);
nand U8352 (N_8352,N_7193,N_7745);
nand U8353 (N_8353,N_7079,N_7361);
or U8354 (N_8354,N_7532,N_7258);
nand U8355 (N_8355,N_7298,N_7574);
xor U8356 (N_8356,N_7202,N_7820);
nand U8357 (N_8357,N_7166,N_7365);
xnor U8358 (N_8358,N_7559,N_7117);
and U8359 (N_8359,N_7938,N_7669);
nor U8360 (N_8360,N_7836,N_7190);
or U8361 (N_8361,N_7015,N_7153);
nor U8362 (N_8362,N_7111,N_7629);
and U8363 (N_8363,N_7352,N_7700);
and U8364 (N_8364,N_7291,N_7518);
or U8365 (N_8365,N_7931,N_7364);
nor U8366 (N_8366,N_7732,N_7276);
xnor U8367 (N_8367,N_7560,N_7984);
nor U8368 (N_8368,N_7705,N_7876);
and U8369 (N_8369,N_7777,N_7683);
nor U8370 (N_8370,N_7954,N_7627);
nand U8371 (N_8371,N_7801,N_7073);
and U8372 (N_8372,N_7536,N_7968);
or U8373 (N_8373,N_7951,N_7748);
nand U8374 (N_8374,N_7674,N_7349);
nor U8375 (N_8375,N_7208,N_7815);
nor U8376 (N_8376,N_7037,N_7508);
or U8377 (N_8377,N_7917,N_7922);
or U8378 (N_8378,N_7149,N_7563);
xnor U8379 (N_8379,N_7304,N_7410);
xor U8380 (N_8380,N_7279,N_7771);
nand U8381 (N_8381,N_7919,N_7100);
nor U8382 (N_8382,N_7775,N_7883);
nor U8383 (N_8383,N_7214,N_7752);
nor U8384 (N_8384,N_7421,N_7345);
xnor U8385 (N_8385,N_7490,N_7429);
xnor U8386 (N_8386,N_7434,N_7448);
xor U8387 (N_8387,N_7747,N_7494);
and U8388 (N_8388,N_7108,N_7911);
nor U8389 (N_8389,N_7619,N_7710);
or U8390 (N_8390,N_7749,N_7967);
or U8391 (N_8391,N_7766,N_7738);
and U8392 (N_8392,N_7980,N_7924);
nor U8393 (N_8393,N_7485,N_7676);
and U8394 (N_8394,N_7260,N_7872);
and U8395 (N_8395,N_7624,N_7228);
and U8396 (N_8396,N_7457,N_7432);
nand U8397 (N_8397,N_7554,N_7341);
nand U8398 (N_8398,N_7480,N_7461);
and U8399 (N_8399,N_7851,N_7425);
and U8400 (N_8400,N_7146,N_7026);
nor U8401 (N_8401,N_7746,N_7481);
nor U8402 (N_8402,N_7205,N_7798);
nand U8403 (N_8403,N_7557,N_7184);
xnor U8404 (N_8404,N_7916,N_7893);
or U8405 (N_8405,N_7275,N_7262);
or U8406 (N_8406,N_7614,N_7972);
xnor U8407 (N_8407,N_7643,N_7159);
nand U8408 (N_8408,N_7623,N_7011);
xnor U8409 (N_8409,N_7192,N_7466);
nand U8410 (N_8410,N_7612,N_7608);
and U8411 (N_8411,N_7368,N_7336);
xnor U8412 (N_8412,N_7520,N_7066);
nand U8413 (N_8413,N_7213,N_7805);
or U8414 (N_8414,N_7390,N_7995);
and U8415 (N_8415,N_7408,N_7889);
and U8416 (N_8416,N_7155,N_7198);
nor U8417 (N_8417,N_7949,N_7838);
and U8418 (N_8418,N_7112,N_7121);
or U8419 (N_8419,N_7424,N_7921);
nor U8420 (N_8420,N_7032,N_7172);
nand U8421 (N_8421,N_7150,N_7023);
or U8422 (N_8422,N_7103,N_7812);
nand U8423 (N_8423,N_7035,N_7067);
nor U8424 (N_8424,N_7626,N_7474);
or U8425 (N_8425,N_7809,N_7821);
nor U8426 (N_8426,N_7541,N_7583);
or U8427 (N_8427,N_7599,N_7655);
nor U8428 (N_8428,N_7094,N_7573);
nor U8429 (N_8429,N_7553,N_7128);
nor U8430 (N_8430,N_7999,N_7870);
nand U8431 (N_8431,N_7594,N_7837);
and U8432 (N_8432,N_7169,N_7660);
or U8433 (N_8433,N_7808,N_7973);
nor U8434 (N_8434,N_7270,N_7769);
and U8435 (N_8435,N_7131,N_7807);
or U8436 (N_8436,N_7607,N_7707);
and U8437 (N_8437,N_7960,N_7986);
nand U8438 (N_8438,N_7020,N_7116);
and U8439 (N_8439,N_7137,N_7321);
or U8440 (N_8440,N_7139,N_7500);
xor U8441 (N_8441,N_7256,N_7797);
nor U8442 (N_8442,N_7666,N_7729);
or U8443 (N_8443,N_7603,N_7317);
nor U8444 (N_8444,N_7970,N_7817);
nor U8445 (N_8445,N_7680,N_7050);
nor U8446 (N_8446,N_7043,N_7487);
nor U8447 (N_8447,N_7449,N_7283);
nor U8448 (N_8448,N_7957,N_7989);
nand U8449 (N_8449,N_7300,N_7018);
nor U8450 (N_8450,N_7001,N_7704);
xnor U8451 (N_8451,N_7983,N_7045);
nor U8452 (N_8452,N_7315,N_7530);
and U8453 (N_8453,N_7059,N_7309);
nand U8454 (N_8454,N_7266,N_7165);
and U8455 (N_8455,N_7786,N_7080);
nor U8456 (N_8456,N_7170,N_7840);
nand U8457 (N_8457,N_7818,N_7888);
nand U8458 (N_8458,N_7444,N_7544);
or U8459 (N_8459,N_7065,N_7290);
and U8460 (N_8460,N_7964,N_7857);
nand U8461 (N_8461,N_7351,N_7335);
nor U8462 (N_8462,N_7431,N_7633);
and U8463 (N_8463,N_7269,N_7757);
or U8464 (N_8464,N_7014,N_7371);
nand U8465 (N_8465,N_7019,N_7478);
xnor U8466 (N_8466,N_7294,N_7136);
nand U8467 (N_8467,N_7495,N_7436);
nor U8468 (N_8468,N_7221,N_7008);
xor U8469 (N_8469,N_7601,N_7930);
and U8470 (N_8470,N_7716,N_7064);
nor U8471 (N_8471,N_7278,N_7381);
nor U8472 (N_8472,N_7906,N_7046);
and U8473 (N_8473,N_7604,N_7327);
or U8474 (N_8474,N_7245,N_7758);
nand U8475 (N_8475,N_7093,N_7981);
or U8476 (N_8476,N_7203,N_7668);
xnor U8477 (N_8477,N_7288,N_7216);
nor U8478 (N_8478,N_7620,N_7226);
nor U8479 (N_8479,N_7338,N_7135);
and U8480 (N_8480,N_7499,N_7299);
or U8481 (N_8481,N_7289,N_7209);
nand U8482 (N_8482,N_7861,N_7230);
xnor U8483 (N_8483,N_7344,N_7936);
nor U8484 (N_8484,N_7686,N_7959);
and U8485 (N_8485,N_7454,N_7519);
and U8486 (N_8486,N_7803,N_7326);
xnor U8487 (N_8487,N_7692,N_7823);
nand U8488 (N_8488,N_7347,N_7402);
or U8489 (N_8489,N_7016,N_7835);
nor U8490 (N_8490,N_7724,N_7464);
nor U8491 (N_8491,N_7342,N_7231);
nor U8492 (N_8492,N_7848,N_7148);
xor U8493 (N_8493,N_7004,N_7644);
nor U8494 (N_8494,N_7943,N_7696);
or U8495 (N_8495,N_7156,N_7670);
nand U8496 (N_8496,N_7702,N_7340);
or U8497 (N_8497,N_7994,N_7978);
nand U8498 (N_8498,N_7243,N_7201);
or U8499 (N_8499,N_7865,N_7918);
nand U8500 (N_8500,N_7187,N_7668);
xor U8501 (N_8501,N_7276,N_7317);
and U8502 (N_8502,N_7877,N_7236);
and U8503 (N_8503,N_7078,N_7271);
nand U8504 (N_8504,N_7835,N_7374);
nand U8505 (N_8505,N_7031,N_7627);
nor U8506 (N_8506,N_7899,N_7544);
and U8507 (N_8507,N_7951,N_7609);
or U8508 (N_8508,N_7779,N_7932);
xor U8509 (N_8509,N_7494,N_7450);
xor U8510 (N_8510,N_7175,N_7076);
and U8511 (N_8511,N_7256,N_7225);
xor U8512 (N_8512,N_7799,N_7532);
or U8513 (N_8513,N_7618,N_7069);
nor U8514 (N_8514,N_7413,N_7624);
or U8515 (N_8515,N_7954,N_7592);
nand U8516 (N_8516,N_7456,N_7314);
nor U8517 (N_8517,N_7721,N_7826);
xnor U8518 (N_8518,N_7974,N_7997);
xor U8519 (N_8519,N_7218,N_7208);
xor U8520 (N_8520,N_7580,N_7957);
and U8521 (N_8521,N_7186,N_7197);
or U8522 (N_8522,N_7961,N_7748);
nand U8523 (N_8523,N_7950,N_7775);
xor U8524 (N_8524,N_7739,N_7713);
nand U8525 (N_8525,N_7167,N_7847);
nand U8526 (N_8526,N_7980,N_7118);
nor U8527 (N_8527,N_7760,N_7204);
nor U8528 (N_8528,N_7220,N_7658);
nor U8529 (N_8529,N_7729,N_7161);
and U8530 (N_8530,N_7435,N_7592);
nand U8531 (N_8531,N_7419,N_7543);
or U8532 (N_8532,N_7316,N_7983);
or U8533 (N_8533,N_7245,N_7532);
xnor U8534 (N_8534,N_7233,N_7035);
nand U8535 (N_8535,N_7523,N_7787);
or U8536 (N_8536,N_7898,N_7598);
nor U8537 (N_8537,N_7493,N_7136);
and U8538 (N_8538,N_7928,N_7189);
nor U8539 (N_8539,N_7841,N_7628);
nor U8540 (N_8540,N_7465,N_7394);
xnor U8541 (N_8541,N_7077,N_7287);
nor U8542 (N_8542,N_7616,N_7043);
nand U8543 (N_8543,N_7104,N_7238);
nand U8544 (N_8544,N_7869,N_7825);
or U8545 (N_8545,N_7079,N_7321);
xor U8546 (N_8546,N_7993,N_7956);
nand U8547 (N_8547,N_7428,N_7707);
nand U8548 (N_8548,N_7492,N_7885);
or U8549 (N_8549,N_7603,N_7653);
nor U8550 (N_8550,N_7933,N_7561);
and U8551 (N_8551,N_7844,N_7022);
nand U8552 (N_8552,N_7661,N_7327);
and U8553 (N_8553,N_7497,N_7778);
xor U8554 (N_8554,N_7646,N_7818);
xnor U8555 (N_8555,N_7720,N_7143);
xor U8556 (N_8556,N_7380,N_7560);
and U8557 (N_8557,N_7225,N_7048);
nor U8558 (N_8558,N_7275,N_7644);
and U8559 (N_8559,N_7080,N_7270);
nor U8560 (N_8560,N_7428,N_7838);
or U8561 (N_8561,N_7987,N_7613);
nor U8562 (N_8562,N_7576,N_7106);
nand U8563 (N_8563,N_7432,N_7203);
nand U8564 (N_8564,N_7306,N_7711);
nand U8565 (N_8565,N_7198,N_7751);
nor U8566 (N_8566,N_7536,N_7933);
and U8567 (N_8567,N_7283,N_7506);
xor U8568 (N_8568,N_7305,N_7479);
and U8569 (N_8569,N_7741,N_7420);
nor U8570 (N_8570,N_7606,N_7286);
nand U8571 (N_8571,N_7850,N_7755);
xnor U8572 (N_8572,N_7072,N_7563);
or U8573 (N_8573,N_7020,N_7156);
nor U8574 (N_8574,N_7979,N_7040);
and U8575 (N_8575,N_7501,N_7829);
nand U8576 (N_8576,N_7037,N_7817);
xnor U8577 (N_8577,N_7834,N_7787);
xor U8578 (N_8578,N_7344,N_7364);
nor U8579 (N_8579,N_7387,N_7576);
and U8580 (N_8580,N_7534,N_7304);
nand U8581 (N_8581,N_7931,N_7348);
and U8582 (N_8582,N_7657,N_7856);
or U8583 (N_8583,N_7444,N_7763);
and U8584 (N_8584,N_7559,N_7962);
nand U8585 (N_8585,N_7760,N_7714);
nand U8586 (N_8586,N_7854,N_7221);
nor U8587 (N_8587,N_7465,N_7368);
or U8588 (N_8588,N_7884,N_7468);
and U8589 (N_8589,N_7330,N_7379);
nand U8590 (N_8590,N_7350,N_7977);
and U8591 (N_8591,N_7395,N_7037);
and U8592 (N_8592,N_7163,N_7157);
and U8593 (N_8593,N_7348,N_7881);
nand U8594 (N_8594,N_7790,N_7126);
nand U8595 (N_8595,N_7792,N_7256);
nor U8596 (N_8596,N_7796,N_7432);
and U8597 (N_8597,N_7746,N_7675);
nand U8598 (N_8598,N_7659,N_7452);
nor U8599 (N_8599,N_7368,N_7903);
nand U8600 (N_8600,N_7557,N_7349);
and U8601 (N_8601,N_7991,N_7327);
or U8602 (N_8602,N_7108,N_7020);
xor U8603 (N_8603,N_7582,N_7216);
or U8604 (N_8604,N_7679,N_7785);
and U8605 (N_8605,N_7799,N_7170);
nor U8606 (N_8606,N_7960,N_7250);
or U8607 (N_8607,N_7906,N_7412);
and U8608 (N_8608,N_7746,N_7740);
and U8609 (N_8609,N_7272,N_7360);
nor U8610 (N_8610,N_7416,N_7730);
xnor U8611 (N_8611,N_7162,N_7863);
nor U8612 (N_8612,N_7175,N_7782);
and U8613 (N_8613,N_7170,N_7877);
xnor U8614 (N_8614,N_7143,N_7814);
nor U8615 (N_8615,N_7902,N_7167);
nor U8616 (N_8616,N_7878,N_7802);
and U8617 (N_8617,N_7028,N_7194);
xor U8618 (N_8618,N_7006,N_7329);
xnor U8619 (N_8619,N_7576,N_7324);
xor U8620 (N_8620,N_7325,N_7916);
nor U8621 (N_8621,N_7879,N_7316);
nor U8622 (N_8622,N_7281,N_7074);
and U8623 (N_8623,N_7901,N_7120);
nor U8624 (N_8624,N_7577,N_7319);
and U8625 (N_8625,N_7914,N_7402);
xor U8626 (N_8626,N_7150,N_7670);
nor U8627 (N_8627,N_7072,N_7668);
or U8628 (N_8628,N_7152,N_7283);
or U8629 (N_8629,N_7632,N_7001);
nor U8630 (N_8630,N_7149,N_7748);
nor U8631 (N_8631,N_7360,N_7606);
nand U8632 (N_8632,N_7638,N_7714);
and U8633 (N_8633,N_7474,N_7748);
and U8634 (N_8634,N_7542,N_7859);
nor U8635 (N_8635,N_7211,N_7731);
or U8636 (N_8636,N_7142,N_7924);
or U8637 (N_8637,N_7211,N_7925);
nor U8638 (N_8638,N_7991,N_7939);
nand U8639 (N_8639,N_7158,N_7177);
nor U8640 (N_8640,N_7969,N_7763);
nand U8641 (N_8641,N_7444,N_7910);
nor U8642 (N_8642,N_7009,N_7079);
xnor U8643 (N_8643,N_7315,N_7924);
nand U8644 (N_8644,N_7269,N_7437);
and U8645 (N_8645,N_7293,N_7299);
nor U8646 (N_8646,N_7757,N_7099);
and U8647 (N_8647,N_7082,N_7396);
nor U8648 (N_8648,N_7518,N_7722);
nor U8649 (N_8649,N_7567,N_7190);
nor U8650 (N_8650,N_7275,N_7597);
xor U8651 (N_8651,N_7217,N_7306);
and U8652 (N_8652,N_7486,N_7857);
nand U8653 (N_8653,N_7907,N_7114);
and U8654 (N_8654,N_7432,N_7142);
nor U8655 (N_8655,N_7828,N_7708);
xor U8656 (N_8656,N_7867,N_7459);
or U8657 (N_8657,N_7079,N_7163);
and U8658 (N_8658,N_7084,N_7964);
or U8659 (N_8659,N_7624,N_7334);
xnor U8660 (N_8660,N_7743,N_7505);
xor U8661 (N_8661,N_7481,N_7204);
nand U8662 (N_8662,N_7360,N_7265);
nand U8663 (N_8663,N_7477,N_7243);
xnor U8664 (N_8664,N_7866,N_7067);
and U8665 (N_8665,N_7387,N_7847);
or U8666 (N_8666,N_7444,N_7930);
or U8667 (N_8667,N_7466,N_7202);
or U8668 (N_8668,N_7177,N_7485);
or U8669 (N_8669,N_7651,N_7213);
and U8670 (N_8670,N_7943,N_7779);
xnor U8671 (N_8671,N_7372,N_7643);
or U8672 (N_8672,N_7666,N_7252);
xor U8673 (N_8673,N_7152,N_7974);
nand U8674 (N_8674,N_7132,N_7731);
or U8675 (N_8675,N_7325,N_7277);
or U8676 (N_8676,N_7754,N_7495);
and U8677 (N_8677,N_7750,N_7556);
and U8678 (N_8678,N_7769,N_7972);
or U8679 (N_8679,N_7398,N_7489);
nand U8680 (N_8680,N_7052,N_7820);
nor U8681 (N_8681,N_7804,N_7945);
or U8682 (N_8682,N_7770,N_7703);
or U8683 (N_8683,N_7762,N_7395);
nand U8684 (N_8684,N_7216,N_7256);
xor U8685 (N_8685,N_7148,N_7822);
and U8686 (N_8686,N_7878,N_7196);
nor U8687 (N_8687,N_7092,N_7446);
nand U8688 (N_8688,N_7663,N_7246);
xnor U8689 (N_8689,N_7307,N_7105);
nand U8690 (N_8690,N_7914,N_7327);
xor U8691 (N_8691,N_7181,N_7250);
xnor U8692 (N_8692,N_7906,N_7426);
xnor U8693 (N_8693,N_7803,N_7057);
xnor U8694 (N_8694,N_7903,N_7732);
and U8695 (N_8695,N_7465,N_7241);
and U8696 (N_8696,N_7962,N_7680);
and U8697 (N_8697,N_7108,N_7917);
nor U8698 (N_8698,N_7077,N_7769);
or U8699 (N_8699,N_7429,N_7857);
nor U8700 (N_8700,N_7732,N_7610);
nand U8701 (N_8701,N_7885,N_7638);
or U8702 (N_8702,N_7072,N_7257);
or U8703 (N_8703,N_7502,N_7850);
or U8704 (N_8704,N_7362,N_7184);
nand U8705 (N_8705,N_7491,N_7763);
nor U8706 (N_8706,N_7482,N_7910);
nor U8707 (N_8707,N_7735,N_7780);
and U8708 (N_8708,N_7581,N_7332);
nor U8709 (N_8709,N_7975,N_7884);
and U8710 (N_8710,N_7073,N_7481);
nor U8711 (N_8711,N_7211,N_7026);
or U8712 (N_8712,N_7561,N_7045);
or U8713 (N_8713,N_7638,N_7141);
nor U8714 (N_8714,N_7847,N_7605);
or U8715 (N_8715,N_7779,N_7118);
nor U8716 (N_8716,N_7806,N_7758);
nor U8717 (N_8717,N_7407,N_7092);
nor U8718 (N_8718,N_7630,N_7026);
or U8719 (N_8719,N_7127,N_7608);
nor U8720 (N_8720,N_7108,N_7122);
xor U8721 (N_8721,N_7203,N_7436);
or U8722 (N_8722,N_7806,N_7093);
nor U8723 (N_8723,N_7130,N_7085);
nor U8724 (N_8724,N_7548,N_7087);
and U8725 (N_8725,N_7444,N_7103);
nor U8726 (N_8726,N_7715,N_7879);
nand U8727 (N_8727,N_7932,N_7048);
or U8728 (N_8728,N_7830,N_7899);
and U8729 (N_8729,N_7545,N_7449);
and U8730 (N_8730,N_7605,N_7809);
nand U8731 (N_8731,N_7707,N_7201);
nand U8732 (N_8732,N_7882,N_7858);
and U8733 (N_8733,N_7062,N_7045);
nand U8734 (N_8734,N_7919,N_7578);
nor U8735 (N_8735,N_7161,N_7360);
and U8736 (N_8736,N_7878,N_7902);
nand U8737 (N_8737,N_7120,N_7073);
xor U8738 (N_8738,N_7071,N_7959);
and U8739 (N_8739,N_7595,N_7671);
and U8740 (N_8740,N_7208,N_7402);
and U8741 (N_8741,N_7181,N_7028);
and U8742 (N_8742,N_7600,N_7307);
or U8743 (N_8743,N_7427,N_7164);
or U8744 (N_8744,N_7520,N_7983);
nor U8745 (N_8745,N_7525,N_7415);
xor U8746 (N_8746,N_7698,N_7092);
or U8747 (N_8747,N_7845,N_7014);
or U8748 (N_8748,N_7121,N_7758);
nand U8749 (N_8749,N_7088,N_7949);
xor U8750 (N_8750,N_7672,N_7629);
and U8751 (N_8751,N_7568,N_7929);
and U8752 (N_8752,N_7525,N_7207);
nor U8753 (N_8753,N_7493,N_7870);
and U8754 (N_8754,N_7828,N_7492);
nand U8755 (N_8755,N_7999,N_7568);
or U8756 (N_8756,N_7603,N_7138);
and U8757 (N_8757,N_7085,N_7847);
or U8758 (N_8758,N_7615,N_7337);
xnor U8759 (N_8759,N_7447,N_7813);
xor U8760 (N_8760,N_7021,N_7988);
or U8761 (N_8761,N_7466,N_7213);
nor U8762 (N_8762,N_7452,N_7789);
nor U8763 (N_8763,N_7118,N_7371);
or U8764 (N_8764,N_7324,N_7922);
or U8765 (N_8765,N_7252,N_7647);
and U8766 (N_8766,N_7847,N_7661);
nand U8767 (N_8767,N_7287,N_7010);
xnor U8768 (N_8768,N_7021,N_7087);
and U8769 (N_8769,N_7321,N_7522);
nor U8770 (N_8770,N_7640,N_7099);
xnor U8771 (N_8771,N_7055,N_7378);
nor U8772 (N_8772,N_7118,N_7175);
xor U8773 (N_8773,N_7088,N_7875);
xor U8774 (N_8774,N_7772,N_7313);
nand U8775 (N_8775,N_7711,N_7347);
nand U8776 (N_8776,N_7104,N_7014);
nor U8777 (N_8777,N_7305,N_7626);
nand U8778 (N_8778,N_7744,N_7090);
or U8779 (N_8779,N_7262,N_7209);
xnor U8780 (N_8780,N_7531,N_7338);
or U8781 (N_8781,N_7374,N_7589);
and U8782 (N_8782,N_7285,N_7124);
or U8783 (N_8783,N_7492,N_7471);
or U8784 (N_8784,N_7273,N_7474);
xor U8785 (N_8785,N_7867,N_7687);
nor U8786 (N_8786,N_7561,N_7740);
and U8787 (N_8787,N_7797,N_7200);
nor U8788 (N_8788,N_7216,N_7186);
nor U8789 (N_8789,N_7242,N_7788);
or U8790 (N_8790,N_7604,N_7664);
xnor U8791 (N_8791,N_7906,N_7696);
nor U8792 (N_8792,N_7895,N_7283);
and U8793 (N_8793,N_7103,N_7614);
xor U8794 (N_8794,N_7015,N_7736);
or U8795 (N_8795,N_7020,N_7511);
nand U8796 (N_8796,N_7661,N_7222);
xor U8797 (N_8797,N_7010,N_7333);
xnor U8798 (N_8798,N_7265,N_7918);
xor U8799 (N_8799,N_7135,N_7421);
or U8800 (N_8800,N_7560,N_7814);
nand U8801 (N_8801,N_7254,N_7766);
nand U8802 (N_8802,N_7611,N_7582);
xnor U8803 (N_8803,N_7835,N_7265);
nand U8804 (N_8804,N_7309,N_7241);
or U8805 (N_8805,N_7842,N_7522);
nor U8806 (N_8806,N_7602,N_7471);
xor U8807 (N_8807,N_7866,N_7685);
xnor U8808 (N_8808,N_7557,N_7767);
nand U8809 (N_8809,N_7702,N_7534);
or U8810 (N_8810,N_7822,N_7103);
xnor U8811 (N_8811,N_7382,N_7834);
and U8812 (N_8812,N_7550,N_7209);
nor U8813 (N_8813,N_7678,N_7093);
xnor U8814 (N_8814,N_7015,N_7816);
or U8815 (N_8815,N_7949,N_7033);
and U8816 (N_8816,N_7249,N_7887);
or U8817 (N_8817,N_7630,N_7878);
nand U8818 (N_8818,N_7105,N_7627);
nand U8819 (N_8819,N_7019,N_7085);
nand U8820 (N_8820,N_7041,N_7351);
nor U8821 (N_8821,N_7997,N_7579);
xnor U8822 (N_8822,N_7967,N_7589);
or U8823 (N_8823,N_7746,N_7509);
and U8824 (N_8824,N_7709,N_7972);
or U8825 (N_8825,N_7130,N_7335);
xnor U8826 (N_8826,N_7005,N_7247);
and U8827 (N_8827,N_7270,N_7989);
or U8828 (N_8828,N_7203,N_7053);
and U8829 (N_8829,N_7543,N_7002);
xnor U8830 (N_8830,N_7951,N_7138);
xnor U8831 (N_8831,N_7989,N_7574);
nor U8832 (N_8832,N_7664,N_7960);
nand U8833 (N_8833,N_7294,N_7853);
nand U8834 (N_8834,N_7376,N_7883);
or U8835 (N_8835,N_7149,N_7761);
or U8836 (N_8836,N_7241,N_7649);
xnor U8837 (N_8837,N_7995,N_7085);
and U8838 (N_8838,N_7001,N_7231);
nor U8839 (N_8839,N_7124,N_7738);
nand U8840 (N_8840,N_7352,N_7106);
xor U8841 (N_8841,N_7153,N_7624);
xor U8842 (N_8842,N_7019,N_7733);
nor U8843 (N_8843,N_7095,N_7699);
nand U8844 (N_8844,N_7501,N_7856);
nor U8845 (N_8845,N_7405,N_7076);
or U8846 (N_8846,N_7664,N_7748);
and U8847 (N_8847,N_7564,N_7747);
xnor U8848 (N_8848,N_7883,N_7071);
and U8849 (N_8849,N_7850,N_7589);
nor U8850 (N_8850,N_7466,N_7876);
nor U8851 (N_8851,N_7245,N_7655);
nor U8852 (N_8852,N_7332,N_7338);
nand U8853 (N_8853,N_7105,N_7011);
xnor U8854 (N_8854,N_7674,N_7248);
xnor U8855 (N_8855,N_7153,N_7835);
xor U8856 (N_8856,N_7526,N_7166);
nand U8857 (N_8857,N_7658,N_7941);
nand U8858 (N_8858,N_7694,N_7877);
and U8859 (N_8859,N_7848,N_7545);
nor U8860 (N_8860,N_7913,N_7640);
xnor U8861 (N_8861,N_7683,N_7194);
xor U8862 (N_8862,N_7686,N_7141);
and U8863 (N_8863,N_7613,N_7302);
xnor U8864 (N_8864,N_7466,N_7498);
nor U8865 (N_8865,N_7762,N_7039);
or U8866 (N_8866,N_7400,N_7504);
xor U8867 (N_8867,N_7138,N_7009);
and U8868 (N_8868,N_7678,N_7118);
or U8869 (N_8869,N_7787,N_7073);
xnor U8870 (N_8870,N_7476,N_7075);
xnor U8871 (N_8871,N_7800,N_7655);
nor U8872 (N_8872,N_7689,N_7848);
nand U8873 (N_8873,N_7640,N_7841);
nand U8874 (N_8874,N_7958,N_7634);
nor U8875 (N_8875,N_7381,N_7592);
or U8876 (N_8876,N_7313,N_7056);
xor U8877 (N_8877,N_7450,N_7139);
nand U8878 (N_8878,N_7233,N_7120);
nand U8879 (N_8879,N_7767,N_7490);
and U8880 (N_8880,N_7621,N_7704);
nand U8881 (N_8881,N_7594,N_7097);
and U8882 (N_8882,N_7562,N_7541);
xnor U8883 (N_8883,N_7434,N_7386);
nand U8884 (N_8884,N_7045,N_7886);
or U8885 (N_8885,N_7073,N_7610);
nand U8886 (N_8886,N_7723,N_7651);
or U8887 (N_8887,N_7857,N_7091);
nor U8888 (N_8888,N_7011,N_7256);
xnor U8889 (N_8889,N_7921,N_7506);
nand U8890 (N_8890,N_7161,N_7361);
nand U8891 (N_8891,N_7533,N_7582);
nand U8892 (N_8892,N_7695,N_7262);
nor U8893 (N_8893,N_7257,N_7059);
xor U8894 (N_8894,N_7404,N_7796);
and U8895 (N_8895,N_7220,N_7215);
or U8896 (N_8896,N_7927,N_7905);
nor U8897 (N_8897,N_7519,N_7924);
and U8898 (N_8898,N_7017,N_7771);
xor U8899 (N_8899,N_7975,N_7091);
and U8900 (N_8900,N_7600,N_7948);
or U8901 (N_8901,N_7368,N_7460);
nor U8902 (N_8902,N_7931,N_7209);
nor U8903 (N_8903,N_7752,N_7067);
nor U8904 (N_8904,N_7262,N_7383);
or U8905 (N_8905,N_7200,N_7566);
and U8906 (N_8906,N_7113,N_7616);
nor U8907 (N_8907,N_7815,N_7836);
xor U8908 (N_8908,N_7829,N_7993);
xnor U8909 (N_8909,N_7045,N_7924);
xor U8910 (N_8910,N_7185,N_7412);
or U8911 (N_8911,N_7759,N_7046);
or U8912 (N_8912,N_7990,N_7886);
xnor U8913 (N_8913,N_7698,N_7032);
nand U8914 (N_8914,N_7257,N_7354);
nor U8915 (N_8915,N_7591,N_7738);
nand U8916 (N_8916,N_7046,N_7908);
and U8917 (N_8917,N_7970,N_7457);
xor U8918 (N_8918,N_7860,N_7407);
or U8919 (N_8919,N_7493,N_7538);
and U8920 (N_8920,N_7029,N_7962);
and U8921 (N_8921,N_7164,N_7673);
or U8922 (N_8922,N_7160,N_7715);
or U8923 (N_8923,N_7104,N_7974);
or U8924 (N_8924,N_7573,N_7624);
xnor U8925 (N_8925,N_7163,N_7562);
xnor U8926 (N_8926,N_7247,N_7117);
xor U8927 (N_8927,N_7886,N_7846);
nor U8928 (N_8928,N_7060,N_7077);
nor U8929 (N_8929,N_7515,N_7301);
and U8930 (N_8930,N_7461,N_7122);
xor U8931 (N_8931,N_7397,N_7795);
or U8932 (N_8932,N_7909,N_7812);
nor U8933 (N_8933,N_7536,N_7744);
and U8934 (N_8934,N_7981,N_7364);
xor U8935 (N_8935,N_7042,N_7978);
nor U8936 (N_8936,N_7670,N_7755);
and U8937 (N_8937,N_7472,N_7827);
nor U8938 (N_8938,N_7707,N_7649);
and U8939 (N_8939,N_7229,N_7263);
nor U8940 (N_8940,N_7078,N_7410);
nor U8941 (N_8941,N_7410,N_7620);
or U8942 (N_8942,N_7134,N_7215);
xor U8943 (N_8943,N_7432,N_7552);
nor U8944 (N_8944,N_7960,N_7545);
or U8945 (N_8945,N_7353,N_7519);
xor U8946 (N_8946,N_7821,N_7030);
nand U8947 (N_8947,N_7311,N_7561);
and U8948 (N_8948,N_7295,N_7787);
nor U8949 (N_8949,N_7381,N_7262);
and U8950 (N_8950,N_7615,N_7903);
and U8951 (N_8951,N_7575,N_7163);
nand U8952 (N_8952,N_7167,N_7389);
xor U8953 (N_8953,N_7368,N_7608);
or U8954 (N_8954,N_7869,N_7177);
nor U8955 (N_8955,N_7066,N_7461);
nand U8956 (N_8956,N_7536,N_7466);
and U8957 (N_8957,N_7463,N_7023);
and U8958 (N_8958,N_7931,N_7339);
xnor U8959 (N_8959,N_7221,N_7191);
and U8960 (N_8960,N_7569,N_7304);
xnor U8961 (N_8961,N_7230,N_7635);
and U8962 (N_8962,N_7841,N_7856);
nand U8963 (N_8963,N_7970,N_7954);
and U8964 (N_8964,N_7674,N_7772);
or U8965 (N_8965,N_7753,N_7392);
nand U8966 (N_8966,N_7635,N_7288);
and U8967 (N_8967,N_7679,N_7885);
or U8968 (N_8968,N_7228,N_7112);
and U8969 (N_8969,N_7478,N_7898);
nor U8970 (N_8970,N_7463,N_7812);
xnor U8971 (N_8971,N_7566,N_7465);
xor U8972 (N_8972,N_7159,N_7064);
or U8973 (N_8973,N_7984,N_7115);
xor U8974 (N_8974,N_7866,N_7391);
and U8975 (N_8975,N_7184,N_7301);
nor U8976 (N_8976,N_7154,N_7612);
nand U8977 (N_8977,N_7680,N_7043);
nand U8978 (N_8978,N_7725,N_7207);
or U8979 (N_8979,N_7911,N_7561);
xnor U8980 (N_8980,N_7816,N_7043);
nor U8981 (N_8981,N_7334,N_7054);
or U8982 (N_8982,N_7726,N_7138);
xor U8983 (N_8983,N_7086,N_7514);
xor U8984 (N_8984,N_7375,N_7250);
xor U8985 (N_8985,N_7262,N_7950);
xor U8986 (N_8986,N_7867,N_7232);
xor U8987 (N_8987,N_7378,N_7652);
and U8988 (N_8988,N_7965,N_7159);
nand U8989 (N_8989,N_7128,N_7182);
and U8990 (N_8990,N_7649,N_7806);
nand U8991 (N_8991,N_7952,N_7564);
and U8992 (N_8992,N_7483,N_7594);
or U8993 (N_8993,N_7356,N_7804);
and U8994 (N_8994,N_7154,N_7856);
and U8995 (N_8995,N_7932,N_7256);
nor U8996 (N_8996,N_7946,N_7528);
nand U8997 (N_8997,N_7847,N_7750);
xor U8998 (N_8998,N_7073,N_7847);
or U8999 (N_8999,N_7550,N_7335);
nand U9000 (N_9000,N_8124,N_8429);
or U9001 (N_9001,N_8994,N_8688);
and U9002 (N_9002,N_8712,N_8562);
and U9003 (N_9003,N_8921,N_8896);
and U9004 (N_9004,N_8052,N_8526);
nand U9005 (N_9005,N_8380,N_8414);
nor U9006 (N_9006,N_8598,N_8021);
or U9007 (N_9007,N_8156,N_8684);
nor U9008 (N_9008,N_8547,N_8845);
nand U9009 (N_9009,N_8357,N_8633);
xor U9010 (N_9010,N_8116,N_8563);
and U9011 (N_9011,N_8827,N_8410);
nand U9012 (N_9012,N_8325,N_8850);
nand U9013 (N_9013,N_8370,N_8589);
xnor U9014 (N_9014,N_8530,N_8915);
xnor U9015 (N_9015,N_8159,N_8846);
nand U9016 (N_9016,N_8222,N_8946);
nand U9017 (N_9017,N_8791,N_8165);
or U9018 (N_9018,N_8236,N_8487);
or U9019 (N_9019,N_8465,N_8076);
xor U9020 (N_9020,N_8592,N_8331);
xor U9021 (N_9021,N_8498,N_8652);
and U9022 (N_9022,N_8777,N_8211);
nand U9023 (N_9023,N_8054,N_8287);
xnor U9024 (N_9024,N_8018,N_8205);
nand U9025 (N_9025,N_8286,N_8735);
nand U9026 (N_9026,N_8233,N_8208);
or U9027 (N_9027,N_8333,N_8740);
nand U9028 (N_9028,N_8085,N_8677);
nor U9029 (N_9029,N_8985,N_8982);
and U9030 (N_9030,N_8489,N_8171);
nor U9031 (N_9031,N_8948,N_8014);
and U9032 (N_9032,N_8394,N_8893);
nor U9033 (N_9033,N_8901,N_8306);
nor U9034 (N_9034,N_8464,N_8163);
nor U9035 (N_9035,N_8518,N_8265);
nor U9036 (N_9036,N_8651,N_8919);
nand U9037 (N_9037,N_8935,N_8483);
and U9038 (N_9038,N_8904,N_8412);
nand U9039 (N_9039,N_8296,N_8593);
xnor U9040 (N_9040,N_8198,N_8486);
or U9041 (N_9041,N_8046,N_8324);
xnor U9042 (N_9042,N_8476,N_8223);
xor U9043 (N_9043,N_8319,N_8241);
or U9044 (N_9044,N_8199,N_8491);
or U9045 (N_9045,N_8421,N_8685);
or U9046 (N_9046,N_8601,N_8271);
or U9047 (N_9047,N_8079,N_8709);
nor U9048 (N_9048,N_8642,N_8504);
and U9049 (N_9049,N_8187,N_8767);
or U9050 (N_9050,N_8965,N_8871);
and U9051 (N_9051,N_8248,N_8913);
and U9052 (N_9052,N_8023,N_8981);
xnor U9053 (N_9053,N_8978,N_8797);
xor U9054 (N_9054,N_8989,N_8837);
or U9055 (N_9055,N_8903,N_8335);
nand U9056 (N_9056,N_8449,N_8392);
or U9057 (N_9057,N_8471,N_8283);
nand U9058 (N_9058,N_8717,N_8454);
or U9059 (N_9059,N_8969,N_8127);
and U9060 (N_9060,N_8799,N_8524);
or U9061 (N_9061,N_8334,N_8502);
xor U9062 (N_9062,N_8275,N_8117);
nor U9063 (N_9063,N_8875,N_8359);
xor U9064 (N_9064,N_8765,N_8890);
nor U9065 (N_9065,N_8231,N_8868);
or U9066 (N_9066,N_8129,N_8702);
xor U9067 (N_9067,N_8847,N_8250);
and U9068 (N_9068,N_8861,N_8910);
xnor U9069 (N_9069,N_8361,N_8182);
nor U9070 (N_9070,N_8907,N_8457);
xnor U9071 (N_9071,N_8103,N_8654);
nor U9072 (N_9072,N_8555,N_8713);
and U9073 (N_9073,N_8751,N_8836);
or U9074 (N_9074,N_8295,N_8379);
nor U9075 (N_9075,N_8191,N_8297);
and U9076 (N_9076,N_8584,N_8136);
xnor U9077 (N_9077,N_8812,N_8973);
xnor U9078 (N_9078,N_8667,N_8822);
nor U9079 (N_9079,N_8309,N_8459);
nor U9080 (N_9080,N_8927,N_8849);
nor U9081 (N_9081,N_8075,N_8147);
nand U9082 (N_9082,N_8118,N_8824);
nor U9083 (N_9083,N_8255,N_8062);
or U9084 (N_9084,N_8436,N_8643);
nor U9085 (N_9085,N_8467,N_8523);
nand U9086 (N_9086,N_8603,N_8407);
nor U9087 (N_9087,N_8839,N_8285);
and U9088 (N_9088,N_8902,N_8786);
or U9089 (N_9089,N_8121,N_8444);
and U9090 (N_9090,N_8605,N_8888);
xor U9091 (N_9091,N_8550,N_8556);
nand U9092 (N_9092,N_8269,N_8762);
nor U9093 (N_9093,N_8142,N_8932);
xor U9094 (N_9094,N_8829,N_8646);
xor U9095 (N_9095,N_8573,N_8472);
and U9096 (N_9096,N_8814,N_8192);
or U9097 (N_9097,N_8945,N_8671);
nand U9098 (N_9098,N_8899,N_8680);
and U9099 (N_9099,N_8425,N_8608);
and U9100 (N_9100,N_8235,N_8461);
or U9101 (N_9101,N_8662,N_8660);
or U9102 (N_9102,N_8322,N_8544);
or U9103 (N_9103,N_8466,N_8928);
or U9104 (N_9104,N_8534,N_8403);
nand U9105 (N_9105,N_8013,N_8715);
nor U9106 (N_9106,N_8417,N_8186);
xor U9107 (N_9107,N_8724,N_8962);
xnor U9108 (N_9108,N_8941,N_8298);
or U9109 (N_9109,N_8661,N_8863);
nor U9110 (N_9110,N_8923,N_8036);
or U9111 (N_9111,N_8882,N_8282);
and U9112 (N_9112,N_8115,N_8207);
xnor U9113 (N_9113,N_8374,N_8914);
and U9114 (N_9114,N_8826,N_8637);
nor U9115 (N_9115,N_8060,N_8760);
and U9116 (N_9116,N_8545,N_8126);
nor U9117 (N_9117,N_8011,N_8521);
nor U9118 (N_9118,N_8405,N_8996);
nand U9119 (N_9119,N_8745,N_8656);
and U9120 (N_9120,N_8574,N_8632);
nor U9121 (N_9121,N_8299,N_8068);
nor U9122 (N_9122,N_8369,N_8067);
nor U9123 (N_9123,N_8423,N_8691);
nor U9124 (N_9124,N_8422,N_8936);
or U9125 (N_9125,N_8727,N_8259);
or U9126 (N_9126,N_8307,N_8585);
nor U9127 (N_9127,N_8440,N_8830);
xor U9128 (N_9128,N_8352,N_8986);
and U9129 (N_9129,N_8097,N_8228);
or U9130 (N_9130,N_8100,N_8516);
nand U9131 (N_9131,N_8772,N_8610);
nand U9132 (N_9132,N_8279,N_8818);
xnor U9133 (N_9133,N_8693,N_8704);
and U9134 (N_9134,N_8729,N_8096);
and U9135 (N_9135,N_8859,N_8758);
and U9136 (N_9136,N_8597,N_8153);
xnor U9137 (N_9137,N_8569,N_8719);
or U9138 (N_9138,N_8088,N_8943);
and U9139 (N_9139,N_8220,N_8918);
nor U9140 (N_9140,N_8794,N_8533);
or U9141 (N_9141,N_8615,N_8017);
nor U9142 (N_9142,N_8674,N_8304);
xnor U9143 (N_9143,N_8694,N_8764);
or U9144 (N_9144,N_8061,N_8215);
and U9145 (N_9145,N_8441,N_8672);
nand U9146 (N_9146,N_8462,N_8320);
or U9147 (N_9147,N_8711,N_8290);
nand U9148 (N_9148,N_8512,N_8501);
nor U9149 (N_9149,N_8788,N_8810);
nand U9150 (N_9150,N_8108,N_8963);
and U9151 (N_9151,N_8773,N_8225);
nor U9152 (N_9152,N_8184,N_8120);
nor U9153 (N_9153,N_8503,N_8431);
nor U9154 (N_9154,N_8926,N_8594);
or U9155 (N_9155,N_8623,N_8009);
nor U9156 (N_9156,N_8987,N_8832);
or U9157 (N_9157,N_8876,N_8289);
nand U9158 (N_9158,N_8496,N_8621);
or U9159 (N_9159,N_8453,N_8995);
nand U9160 (N_9160,N_8212,N_8189);
or U9161 (N_9161,N_8313,N_8239);
or U9162 (N_9162,N_8291,N_8133);
or U9163 (N_9163,N_8485,N_8976);
xnor U9164 (N_9164,N_8625,N_8778);
or U9165 (N_9165,N_8527,N_8174);
xor U9166 (N_9166,N_8734,N_8540);
nor U9167 (N_9167,N_8575,N_8151);
xnor U9168 (N_9168,N_8455,N_8531);
nand U9169 (N_9169,N_8595,N_8041);
and U9170 (N_9170,N_8302,N_8537);
xnor U9171 (N_9171,N_8865,N_8368);
nand U9172 (N_9172,N_8099,N_8549);
xnor U9173 (N_9173,N_8439,N_8327);
nand U9174 (N_9174,N_8841,N_8007);
or U9175 (N_9175,N_8647,N_8609);
and U9176 (N_9176,N_8803,N_8084);
nor U9177 (N_9177,N_8842,N_8063);
nand U9178 (N_9178,N_8348,N_8000);
nand U9179 (N_9179,N_8853,N_8072);
nor U9180 (N_9180,N_8687,N_8997);
xnor U9181 (N_9181,N_8966,N_8696);
nor U9182 (N_9182,N_8137,N_8624);
nor U9183 (N_9183,N_8578,N_8329);
xnor U9184 (N_9184,N_8897,N_8627);
or U9185 (N_9185,N_8351,N_8409);
xnor U9186 (N_9186,N_8415,N_8917);
or U9187 (N_9187,N_8456,N_8170);
nand U9188 (N_9188,N_8194,N_8513);
nor U9189 (N_9189,N_8251,N_8006);
nand U9190 (N_9190,N_8190,N_8834);
nand U9191 (N_9191,N_8668,N_8769);
or U9192 (N_9192,N_8635,N_8056);
or U9193 (N_9193,N_8355,N_8484);
or U9194 (N_9194,N_8612,N_8536);
nand U9195 (N_9195,N_8344,N_8507);
xnor U9196 (N_9196,N_8905,N_8860);
nor U9197 (N_9197,N_8071,N_8892);
xor U9198 (N_9198,N_8188,N_8253);
nor U9199 (N_9199,N_8038,N_8149);
nor U9200 (N_9200,N_8529,N_8360);
xnor U9201 (N_9201,N_8820,N_8977);
or U9202 (N_9202,N_8775,N_8238);
or U9203 (N_9203,N_8553,N_8796);
xnor U9204 (N_9204,N_8774,N_8397);
or U9205 (N_9205,N_8998,N_8446);
and U9206 (N_9206,N_8636,N_8130);
nor U9207 (N_9207,N_8474,N_8604);
nor U9208 (N_9208,N_8204,N_8364);
or U9209 (N_9209,N_8787,N_8073);
or U9210 (N_9210,N_8864,N_8931);
or U9211 (N_9211,N_8318,N_8132);
or U9212 (N_9212,N_8771,N_8937);
nand U9213 (N_9213,N_8398,N_8268);
nand U9214 (N_9214,N_8200,N_8469);
xnor U9215 (N_9215,N_8183,N_8858);
and U9216 (N_9216,N_8128,N_8588);
or U9217 (N_9217,N_8798,N_8257);
nor U9218 (N_9218,N_8037,N_8866);
xor U9219 (N_9219,N_8664,N_8064);
and U9220 (N_9220,N_8505,N_8019);
and U9221 (N_9221,N_8254,N_8424);
nand U9222 (N_9222,N_8669,N_8363);
and U9223 (N_9223,N_8066,N_8003);
nor U9224 (N_9224,N_8305,N_8784);
or U9225 (N_9225,N_8975,N_8070);
nand U9226 (N_9226,N_8280,N_8756);
or U9227 (N_9227,N_8059,N_8809);
nor U9228 (N_9228,N_8166,N_8748);
or U9229 (N_9229,N_8157,N_8728);
xnor U9230 (N_9230,N_8087,N_8972);
xor U9231 (N_9231,N_8494,N_8206);
nor U9232 (N_9232,N_8707,N_8232);
nand U9233 (N_9233,N_8558,N_8631);
or U9234 (N_9234,N_8263,N_8947);
xnor U9235 (N_9235,N_8452,N_8924);
or U9236 (N_9236,N_8091,N_8045);
nor U9237 (N_9237,N_8856,N_8463);
nor U9238 (N_9238,N_8336,N_8991);
xnor U9239 (N_9239,N_8451,N_8539);
or U9240 (N_9240,N_8141,N_8144);
or U9241 (N_9241,N_8763,N_8990);
nand U9242 (N_9242,N_8710,N_8221);
xnor U9243 (N_9243,N_8833,N_8004);
nor U9244 (N_9244,N_8210,N_8025);
and U9245 (N_9245,N_8152,N_8964);
xor U9246 (N_9246,N_8532,N_8113);
nor U9247 (N_9247,N_8673,N_8051);
and U9248 (N_9248,N_8139,N_8074);
and U9249 (N_9249,N_8470,N_8872);
xor U9250 (N_9250,N_8567,N_8332);
xor U9251 (N_9251,N_8804,N_8001);
and U9252 (N_9252,N_8857,N_8506);
nand U9253 (N_9253,N_8042,N_8385);
and U9254 (N_9254,N_8802,N_8922);
or U9255 (N_9255,N_8743,N_8260);
nand U9256 (N_9256,N_8303,N_8277);
or U9257 (N_9257,N_8988,N_8581);
or U9258 (N_9258,N_8010,N_8244);
and U9259 (N_9259,N_8107,N_8600);
xnor U9260 (N_9260,N_8723,N_8911);
and U9261 (N_9261,N_8399,N_8522);
nor U9262 (N_9262,N_8146,N_8193);
or U9263 (N_9263,N_8081,N_8196);
xnor U9264 (N_9264,N_8362,N_8906);
nor U9265 (N_9265,N_8273,N_8747);
and U9266 (N_9266,N_8663,N_8721);
nor U9267 (N_9267,N_8779,N_8511);
nor U9268 (N_9268,N_8434,N_8202);
nand U9269 (N_9269,N_8095,N_8252);
and U9270 (N_9270,N_8817,N_8613);
and U9271 (N_9271,N_8216,N_8381);
nand U9272 (N_9272,N_8920,N_8877);
nor U9273 (N_9273,N_8759,N_8404);
nor U9274 (N_9274,N_8458,N_8909);
xnor U9275 (N_9275,N_8326,N_8638);
nor U9276 (N_9276,N_8201,N_8065);
nor U9277 (N_9277,N_8420,N_8816);
nand U9278 (N_9278,N_8616,N_8925);
and U9279 (N_9279,N_8722,N_8580);
nand U9280 (N_9280,N_8475,N_8078);
and U9281 (N_9281,N_8958,N_8838);
and U9282 (N_9282,N_8950,N_8565);
nand U9283 (N_9283,N_8135,N_8173);
nor U9284 (N_9284,N_8916,N_8180);
and U9285 (N_9285,N_8002,N_8338);
xor U9286 (N_9286,N_8703,N_8618);
nand U9287 (N_9287,N_8757,N_8898);
nand U9288 (N_9288,N_8264,N_8795);
nor U9289 (N_9289,N_8886,N_8161);
nor U9290 (N_9290,N_8761,N_8739);
or U9291 (N_9291,N_8267,N_8870);
xnor U9292 (N_9292,N_8406,N_8102);
xnor U9293 (N_9293,N_8376,N_8214);
or U9294 (N_9294,N_8175,N_8396);
nand U9295 (N_9295,N_8961,N_8270);
nor U9296 (N_9296,N_8587,N_8256);
and U9297 (N_9297,N_8577,N_8579);
and U9298 (N_9298,N_8626,N_8878);
nor U9299 (N_9299,N_8840,N_8249);
and U9300 (N_9300,N_8162,N_8828);
nor U9301 (N_9301,N_8552,N_8288);
xor U9302 (N_9302,N_8445,N_8675);
and U9303 (N_9303,N_8234,N_8330);
nand U9304 (N_9304,N_8611,N_8971);
xor U9305 (N_9305,N_8123,N_8387);
or U9306 (N_9306,N_8509,N_8730);
and U9307 (N_9307,N_8993,N_8705);
nand U9308 (N_9308,N_8493,N_8477);
nor U9309 (N_9309,N_8317,N_8093);
or U9310 (N_9310,N_8177,N_8891);
and U9311 (N_9311,N_8641,N_8430);
xnor U9312 (N_9312,N_8560,N_8571);
and U9313 (N_9313,N_8815,N_8008);
nand U9314 (N_9314,N_8110,N_8698);
xnor U9315 (N_9315,N_8155,N_8040);
nand U9316 (N_9316,N_8960,N_8793);
xor U9317 (N_9317,N_8980,N_8879);
or U9318 (N_9318,N_8999,N_8776);
or U9319 (N_9319,N_8077,N_8554);
or U9320 (N_9320,N_8586,N_8293);
and U9321 (N_9321,N_8572,N_8057);
nand U9322 (N_9322,N_8938,N_8154);
nand U9323 (N_9323,N_8310,N_8510);
and U9324 (N_9324,N_8167,N_8261);
and U9325 (N_9325,N_8679,N_8683);
or U9326 (N_9326,N_8855,N_8419);
and U9327 (N_9327,N_8754,N_8366);
and U9328 (N_9328,N_8746,N_8590);
nand U9329 (N_9329,N_8676,N_8557);
xnor U9330 (N_9330,N_8105,N_8490);
xor U9331 (N_9331,N_8356,N_8854);
xnor U9332 (N_9332,N_8435,N_8949);
nor U9333 (N_9333,N_8346,N_8653);
xnor U9334 (N_9334,N_8753,N_8178);
and U9335 (N_9335,N_8805,N_8952);
xnor U9336 (N_9336,N_8525,N_8350);
or U9337 (N_9337,N_8389,N_8808);
nor U9338 (N_9338,N_8104,N_8650);
and U9339 (N_9339,N_8957,N_8657);
xor U9340 (N_9340,N_8024,N_8033);
or U9341 (N_9341,N_8339,N_8617);
and U9342 (N_9342,N_8145,N_8031);
xnor U9343 (N_9343,N_8227,N_8515);
and U9344 (N_9344,N_8378,N_8602);
or U9345 (N_9345,N_8258,N_8959);
nand U9346 (N_9346,N_8224,N_8542);
xnor U9347 (N_9347,N_8328,N_8681);
and U9348 (N_9348,N_8082,N_8718);
nor U9349 (N_9349,N_8951,N_8874);
nand U9350 (N_9350,N_8852,N_8242);
and U9351 (N_9351,N_8825,N_8873);
xor U9352 (N_9352,N_8245,N_8488);
xnor U9353 (N_9353,N_8596,N_8195);
nand U9354 (N_9354,N_8372,N_8185);
or U9355 (N_9355,N_8321,N_8591);
and U9356 (N_9356,N_8744,N_8164);
xor U9357 (N_9357,N_8114,N_8634);
nand U9358 (N_9358,N_8974,N_8884);
and U9359 (N_9359,N_8934,N_8301);
nand U9360 (N_9360,N_8246,N_8276);
nand U9361 (N_9361,N_8628,N_8714);
or U9362 (N_9362,N_8416,N_8112);
and U9363 (N_9363,N_8738,N_8094);
or U9364 (N_9364,N_8029,N_8811);
or U9365 (N_9365,N_8499,N_8433);
or U9366 (N_9366,N_8150,N_8438);
xor U9367 (N_9367,N_8016,N_8384);
nor U9368 (N_9368,N_8785,N_8312);
nand U9369 (N_9369,N_8039,N_8851);
or U9370 (N_9370,N_8473,N_8284);
and U9371 (N_9371,N_8551,N_8823);
and U9372 (N_9372,N_8408,N_8342);
xor U9373 (N_9373,N_8732,N_8092);
nand U9374 (N_9374,N_8766,N_8880);
or U9375 (N_9375,N_8226,N_8749);
xnor U9376 (N_9376,N_8930,N_8413);
nand U9377 (N_9377,N_8391,N_8752);
and U9378 (N_9378,N_8442,N_8418);
nand U9379 (N_9379,N_8300,N_8701);
nor U9380 (N_9380,N_8055,N_8665);
and U9381 (N_9381,N_8427,N_8122);
nand U9382 (N_9382,N_8022,N_8725);
nand U9383 (N_9383,N_8692,N_8005);
or U9384 (N_9384,N_8807,N_8316);
nand U9385 (N_9385,N_8026,N_8939);
and U9386 (N_9386,N_8292,N_8620);
nor U9387 (N_9387,N_8349,N_8619);
nand U9388 (N_9388,N_8240,N_8800);
or U9389 (N_9389,N_8143,N_8365);
and U9390 (N_9390,N_8311,N_8341);
nor U9391 (N_9391,N_8862,N_8889);
or U9392 (N_9392,N_8479,N_8848);
or U9393 (N_9393,N_8655,N_8308);
nand U9394 (N_9394,N_8520,N_8670);
nand U9395 (N_9395,N_8209,N_8426);
and U9396 (N_9396,N_8373,N_8895);
nor U9397 (N_9397,N_8607,N_8028);
and U9398 (N_9398,N_8648,N_8835);
nand U9399 (N_9399,N_8219,N_8630);
nor U9400 (N_9400,N_8908,N_8168);
xnor U9401 (N_9401,N_8032,N_8885);
xor U9402 (N_9402,N_8682,N_8383);
and U9403 (N_9403,N_8929,N_8755);
nand U9404 (N_9404,N_8700,N_8218);
nand U9405 (N_9405,N_8266,N_8559);
and U9406 (N_9406,N_8375,N_8131);
or U9407 (N_9407,N_8992,N_8367);
xnor U9408 (N_9408,N_8478,N_8111);
xnor U9409 (N_9409,N_8649,N_8247);
nor U9410 (N_9410,N_8371,N_8109);
xnor U9411 (N_9411,N_8514,N_8789);
xnor U9412 (N_9412,N_8720,N_8148);
nor U9413 (N_9413,N_8314,N_8272);
or U9414 (N_9414,N_8582,N_8020);
or U9415 (N_9415,N_8347,N_8213);
nor U9416 (N_9416,N_8048,N_8699);
nand U9417 (N_9417,N_8294,N_8782);
nor U9418 (N_9418,N_8015,N_8912);
xnor U9419 (N_9419,N_8497,N_8736);
nor U9420 (N_9420,N_8706,N_8535);
xnor U9421 (N_9421,N_8731,N_8315);
or U9422 (N_9422,N_8933,N_8716);
nor U9423 (N_9423,N_8733,N_8134);
and U9424 (N_9424,N_8495,N_8690);
nor U9425 (N_9425,N_8393,N_8750);
or U9426 (N_9426,N_8337,N_8323);
nor U9427 (N_9427,N_8158,N_8781);
nor U9428 (N_9428,N_8844,N_8447);
or U9429 (N_9429,N_8086,N_8203);
and U9430 (N_9430,N_8353,N_8027);
nand U9431 (N_9431,N_8528,N_8644);
or U9432 (N_9432,N_8401,N_8639);
nor U9433 (N_9433,N_8894,N_8069);
or U9434 (N_9434,N_8181,N_8443);
nand U9435 (N_9435,N_8695,N_8354);
nand U9436 (N_9436,N_8138,N_8737);
or U9437 (N_9437,N_8140,N_8278);
or U9438 (N_9438,N_8450,N_8678);
nand U9439 (N_9439,N_8570,N_8564);
nor U9440 (N_9440,N_8281,N_8448);
or U9441 (N_9441,N_8172,N_8437);
or U9442 (N_9442,N_8770,N_8119);
nand U9443 (N_9443,N_8358,N_8400);
nand U9444 (N_9444,N_8566,N_8090);
xnor U9445 (N_9445,N_8508,N_8519);
xnor U9446 (N_9446,N_8819,N_8954);
nor U9447 (N_9447,N_8274,N_8377);
and U9448 (N_9448,N_8053,N_8217);
nor U9449 (N_9449,N_8382,N_8390);
nand U9450 (N_9450,N_8098,N_8806);
nand U9451 (N_9451,N_8243,N_8869);
xor U9452 (N_9452,N_8500,N_8125);
xor U9453 (N_9453,N_8395,N_8726);
xnor U9454 (N_9454,N_8237,N_8900);
nand U9455 (N_9455,N_8768,N_8742);
xor U9456 (N_9456,N_8813,N_8229);
and U9457 (N_9457,N_8546,N_8080);
xnor U9458 (N_9458,N_8881,N_8083);
xnor U9459 (N_9459,N_8049,N_8942);
and U9460 (N_9460,N_8801,N_8583);
or U9461 (N_9461,N_8780,N_8340);
xor U9462 (N_9462,N_8940,N_8050);
xor U9463 (N_9463,N_8968,N_8468);
nor U9464 (N_9464,N_8388,N_8599);
and U9465 (N_9465,N_8179,N_8689);
nand U9466 (N_9466,N_8030,N_8058);
and U9467 (N_9467,N_8944,N_8169);
xor U9468 (N_9468,N_8614,N_8983);
nor U9469 (N_9469,N_8659,N_8831);
or U9470 (N_9470,N_8012,N_8043);
and U9471 (N_9471,N_8492,N_8955);
nand U9472 (N_9472,N_8568,N_8541);
and U9473 (N_9473,N_8034,N_8480);
nand U9474 (N_9474,N_8606,N_8460);
and U9475 (N_9475,N_8979,N_8956);
and U9476 (N_9476,N_8345,N_8686);
or U9477 (N_9477,N_8790,N_8481);
nand U9478 (N_9478,N_8658,N_8622);
nor U9479 (N_9479,N_8843,N_8047);
and U9480 (N_9480,N_8402,N_8561);
nand U9481 (N_9481,N_8432,N_8343);
and U9482 (N_9482,N_8101,N_8645);
or U9483 (N_9483,N_8953,N_8089);
or U9484 (N_9484,N_8482,N_8821);
nor U9485 (N_9485,N_8708,N_8640);
and U9486 (N_9486,N_8883,N_8697);
and U9487 (N_9487,N_8197,N_8783);
xnor U9488 (N_9488,N_8666,N_8984);
nor U9489 (N_9489,N_8967,N_8428);
nor U9490 (N_9490,N_8887,N_8262);
nor U9491 (N_9491,N_8176,N_8792);
or U9492 (N_9492,N_8970,N_8867);
or U9493 (N_9493,N_8517,N_8538);
and U9494 (N_9494,N_8548,N_8629);
xnor U9495 (N_9495,N_8230,N_8160);
and U9496 (N_9496,N_8741,N_8035);
xnor U9497 (N_9497,N_8044,N_8386);
or U9498 (N_9498,N_8576,N_8411);
xnor U9499 (N_9499,N_8543,N_8106);
nand U9500 (N_9500,N_8326,N_8892);
and U9501 (N_9501,N_8661,N_8551);
and U9502 (N_9502,N_8014,N_8327);
nor U9503 (N_9503,N_8790,N_8951);
nand U9504 (N_9504,N_8275,N_8309);
xnor U9505 (N_9505,N_8080,N_8763);
and U9506 (N_9506,N_8949,N_8295);
nand U9507 (N_9507,N_8601,N_8886);
nor U9508 (N_9508,N_8297,N_8636);
nand U9509 (N_9509,N_8503,N_8355);
or U9510 (N_9510,N_8510,N_8795);
nor U9511 (N_9511,N_8598,N_8398);
or U9512 (N_9512,N_8880,N_8519);
xor U9513 (N_9513,N_8275,N_8815);
nor U9514 (N_9514,N_8107,N_8710);
nand U9515 (N_9515,N_8830,N_8595);
xor U9516 (N_9516,N_8964,N_8652);
nand U9517 (N_9517,N_8727,N_8961);
and U9518 (N_9518,N_8581,N_8406);
nor U9519 (N_9519,N_8601,N_8439);
and U9520 (N_9520,N_8298,N_8446);
xor U9521 (N_9521,N_8797,N_8867);
or U9522 (N_9522,N_8080,N_8924);
xor U9523 (N_9523,N_8726,N_8014);
xnor U9524 (N_9524,N_8509,N_8258);
nor U9525 (N_9525,N_8638,N_8290);
xnor U9526 (N_9526,N_8170,N_8590);
xor U9527 (N_9527,N_8374,N_8820);
and U9528 (N_9528,N_8123,N_8385);
and U9529 (N_9529,N_8805,N_8353);
or U9530 (N_9530,N_8405,N_8756);
and U9531 (N_9531,N_8332,N_8744);
nand U9532 (N_9532,N_8338,N_8285);
xor U9533 (N_9533,N_8892,N_8799);
nor U9534 (N_9534,N_8055,N_8699);
nor U9535 (N_9535,N_8960,N_8840);
nand U9536 (N_9536,N_8297,N_8902);
xnor U9537 (N_9537,N_8743,N_8367);
and U9538 (N_9538,N_8221,N_8368);
nor U9539 (N_9539,N_8709,N_8786);
xnor U9540 (N_9540,N_8642,N_8084);
xor U9541 (N_9541,N_8513,N_8028);
nand U9542 (N_9542,N_8844,N_8467);
nor U9543 (N_9543,N_8083,N_8193);
nand U9544 (N_9544,N_8042,N_8194);
and U9545 (N_9545,N_8440,N_8427);
or U9546 (N_9546,N_8173,N_8393);
or U9547 (N_9547,N_8899,N_8228);
or U9548 (N_9548,N_8636,N_8493);
nand U9549 (N_9549,N_8065,N_8009);
nand U9550 (N_9550,N_8143,N_8838);
or U9551 (N_9551,N_8104,N_8836);
and U9552 (N_9552,N_8134,N_8124);
nand U9553 (N_9553,N_8406,N_8687);
xor U9554 (N_9554,N_8733,N_8711);
nor U9555 (N_9555,N_8244,N_8466);
and U9556 (N_9556,N_8737,N_8773);
and U9557 (N_9557,N_8442,N_8760);
or U9558 (N_9558,N_8758,N_8650);
and U9559 (N_9559,N_8905,N_8230);
nor U9560 (N_9560,N_8415,N_8647);
xnor U9561 (N_9561,N_8613,N_8157);
or U9562 (N_9562,N_8762,N_8524);
nor U9563 (N_9563,N_8478,N_8816);
nand U9564 (N_9564,N_8979,N_8863);
nand U9565 (N_9565,N_8007,N_8708);
and U9566 (N_9566,N_8507,N_8459);
nor U9567 (N_9567,N_8710,N_8123);
nor U9568 (N_9568,N_8571,N_8976);
nor U9569 (N_9569,N_8896,N_8048);
nand U9570 (N_9570,N_8171,N_8347);
nor U9571 (N_9571,N_8921,N_8040);
and U9572 (N_9572,N_8467,N_8862);
nand U9573 (N_9573,N_8476,N_8866);
nor U9574 (N_9574,N_8059,N_8347);
or U9575 (N_9575,N_8270,N_8928);
xnor U9576 (N_9576,N_8654,N_8381);
and U9577 (N_9577,N_8451,N_8392);
or U9578 (N_9578,N_8457,N_8641);
nand U9579 (N_9579,N_8627,N_8952);
xnor U9580 (N_9580,N_8715,N_8707);
nor U9581 (N_9581,N_8304,N_8563);
or U9582 (N_9582,N_8178,N_8708);
nor U9583 (N_9583,N_8999,N_8920);
or U9584 (N_9584,N_8173,N_8026);
and U9585 (N_9585,N_8650,N_8076);
and U9586 (N_9586,N_8206,N_8400);
and U9587 (N_9587,N_8501,N_8786);
or U9588 (N_9588,N_8932,N_8758);
or U9589 (N_9589,N_8428,N_8437);
and U9590 (N_9590,N_8575,N_8663);
and U9591 (N_9591,N_8654,N_8616);
nor U9592 (N_9592,N_8572,N_8657);
or U9593 (N_9593,N_8224,N_8631);
xor U9594 (N_9594,N_8953,N_8381);
or U9595 (N_9595,N_8394,N_8761);
xor U9596 (N_9596,N_8872,N_8273);
or U9597 (N_9597,N_8422,N_8781);
nand U9598 (N_9598,N_8405,N_8204);
nand U9599 (N_9599,N_8639,N_8379);
or U9600 (N_9600,N_8468,N_8357);
xor U9601 (N_9601,N_8736,N_8961);
xor U9602 (N_9602,N_8005,N_8032);
nand U9603 (N_9603,N_8098,N_8318);
and U9604 (N_9604,N_8215,N_8563);
nand U9605 (N_9605,N_8406,N_8768);
nor U9606 (N_9606,N_8772,N_8165);
nor U9607 (N_9607,N_8538,N_8151);
xor U9608 (N_9608,N_8155,N_8448);
nand U9609 (N_9609,N_8180,N_8104);
nand U9610 (N_9610,N_8072,N_8704);
nand U9611 (N_9611,N_8078,N_8455);
or U9612 (N_9612,N_8529,N_8547);
xnor U9613 (N_9613,N_8802,N_8215);
or U9614 (N_9614,N_8838,N_8754);
nor U9615 (N_9615,N_8172,N_8867);
nor U9616 (N_9616,N_8320,N_8456);
or U9617 (N_9617,N_8773,N_8035);
nand U9618 (N_9618,N_8695,N_8788);
xnor U9619 (N_9619,N_8911,N_8325);
nand U9620 (N_9620,N_8917,N_8667);
or U9621 (N_9621,N_8321,N_8947);
nor U9622 (N_9622,N_8940,N_8258);
nand U9623 (N_9623,N_8507,N_8602);
nor U9624 (N_9624,N_8896,N_8181);
nand U9625 (N_9625,N_8825,N_8492);
nor U9626 (N_9626,N_8669,N_8812);
or U9627 (N_9627,N_8832,N_8353);
xor U9628 (N_9628,N_8996,N_8888);
nor U9629 (N_9629,N_8419,N_8236);
or U9630 (N_9630,N_8240,N_8797);
xor U9631 (N_9631,N_8210,N_8178);
xnor U9632 (N_9632,N_8407,N_8052);
xor U9633 (N_9633,N_8700,N_8342);
nand U9634 (N_9634,N_8198,N_8923);
and U9635 (N_9635,N_8790,N_8722);
nor U9636 (N_9636,N_8378,N_8294);
xnor U9637 (N_9637,N_8659,N_8291);
nand U9638 (N_9638,N_8925,N_8097);
or U9639 (N_9639,N_8195,N_8192);
xnor U9640 (N_9640,N_8969,N_8630);
nand U9641 (N_9641,N_8806,N_8047);
or U9642 (N_9642,N_8221,N_8951);
or U9643 (N_9643,N_8971,N_8454);
or U9644 (N_9644,N_8886,N_8570);
or U9645 (N_9645,N_8519,N_8401);
nor U9646 (N_9646,N_8542,N_8278);
or U9647 (N_9647,N_8722,N_8013);
nor U9648 (N_9648,N_8065,N_8545);
or U9649 (N_9649,N_8428,N_8678);
or U9650 (N_9650,N_8157,N_8383);
nor U9651 (N_9651,N_8189,N_8891);
and U9652 (N_9652,N_8666,N_8491);
nand U9653 (N_9653,N_8641,N_8644);
nor U9654 (N_9654,N_8864,N_8183);
nand U9655 (N_9655,N_8440,N_8408);
nor U9656 (N_9656,N_8818,N_8920);
nand U9657 (N_9657,N_8484,N_8683);
xor U9658 (N_9658,N_8927,N_8963);
and U9659 (N_9659,N_8554,N_8492);
nand U9660 (N_9660,N_8642,N_8759);
and U9661 (N_9661,N_8169,N_8813);
nor U9662 (N_9662,N_8493,N_8633);
xor U9663 (N_9663,N_8476,N_8204);
nand U9664 (N_9664,N_8841,N_8583);
and U9665 (N_9665,N_8323,N_8146);
xnor U9666 (N_9666,N_8186,N_8327);
xor U9667 (N_9667,N_8820,N_8059);
and U9668 (N_9668,N_8123,N_8729);
nor U9669 (N_9669,N_8668,N_8807);
xor U9670 (N_9670,N_8581,N_8045);
nor U9671 (N_9671,N_8296,N_8249);
nand U9672 (N_9672,N_8884,N_8204);
xor U9673 (N_9673,N_8575,N_8589);
nor U9674 (N_9674,N_8976,N_8359);
xor U9675 (N_9675,N_8809,N_8214);
xnor U9676 (N_9676,N_8702,N_8077);
nor U9677 (N_9677,N_8406,N_8032);
nand U9678 (N_9678,N_8758,N_8519);
nand U9679 (N_9679,N_8276,N_8552);
xor U9680 (N_9680,N_8586,N_8369);
or U9681 (N_9681,N_8126,N_8572);
xor U9682 (N_9682,N_8717,N_8615);
nand U9683 (N_9683,N_8634,N_8495);
nor U9684 (N_9684,N_8283,N_8034);
nand U9685 (N_9685,N_8003,N_8167);
and U9686 (N_9686,N_8776,N_8772);
nor U9687 (N_9687,N_8049,N_8582);
nor U9688 (N_9688,N_8435,N_8210);
nand U9689 (N_9689,N_8521,N_8806);
nand U9690 (N_9690,N_8546,N_8831);
xnor U9691 (N_9691,N_8638,N_8135);
and U9692 (N_9692,N_8544,N_8010);
and U9693 (N_9693,N_8687,N_8681);
xor U9694 (N_9694,N_8993,N_8444);
and U9695 (N_9695,N_8395,N_8611);
nand U9696 (N_9696,N_8768,N_8036);
nor U9697 (N_9697,N_8311,N_8184);
nand U9698 (N_9698,N_8315,N_8685);
and U9699 (N_9699,N_8665,N_8654);
nor U9700 (N_9700,N_8799,N_8752);
xnor U9701 (N_9701,N_8999,N_8626);
and U9702 (N_9702,N_8292,N_8503);
nand U9703 (N_9703,N_8838,N_8658);
or U9704 (N_9704,N_8170,N_8937);
xnor U9705 (N_9705,N_8747,N_8185);
or U9706 (N_9706,N_8038,N_8079);
and U9707 (N_9707,N_8891,N_8047);
xnor U9708 (N_9708,N_8620,N_8052);
xnor U9709 (N_9709,N_8880,N_8078);
nor U9710 (N_9710,N_8335,N_8933);
nand U9711 (N_9711,N_8341,N_8742);
nor U9712 (N_9712,N_8548,N_8471);
nand U9713 (N_9713,N_8012,N_8304);
nand U9714 (N_9714,N_8520,N_8142);
nand U9715 (N_9715,N_8945,N_8507);
nor U9716 (N_9716,N_8584,N_8278);
or U9717 (N_9717,N_8390,N_8697);
nor U9718 (N_9718,N_8733,N_8087);
nand U9719 (N_9719,N_8678,N_8623);
or U9720 (N_9720,N_8373,N_8989);
and U9721 (N_9721,N_8506,N_8339);
xnor U9722 (N_9722,N_8089,N_8231);
nand U9723 (N_9723,N_8002,N_8352);
and U9724 (N_9724,N_8687,N_8822);
nand U9725 (N_9725,N_8880,N_8064);
nand U9726 (N_9726,N_8525,N_8026);
nor U9727 (N_9727,N_8684,N_8903);
xor U9728 (N_9728,N_8656,N_8267);
and U9729 (N_9729,N_8019,N_8014);
nand U9730 (N_9730,N_8688,N_8014);
nor U9731 (N_9731,N_8356,N_8977);
xnor U9732 (N_9732,N_8755,N_8650);
or U9733 (N_9733,N_8941,N_8869);
and U9734 (N_9734,N_8890,N_8649);
xor U9735 (N_9735,N_8610,N_8540);
nand U9736 (N_9736,N_8072,N_8712);
xor U9737 (N_9737,N_8315,N_8301);
nor U9738 (N_9738,N_8908,N_8961);
nor U9739 (N_9739,N_8759,N_8400);
nand U9740 (N_9740,N_8899,N_8096);
nor U9741 (N_9741,N_8556,N_8212);
and U9742 (N_9742,N_8366,N_8762);
nor U9743 (N_9743,N_8012,N_8289);
nor U9744 (N_9744,N_8383,N_8410);
nand U9745 (N_9745,N_8805,N_8266);
xnor U9746 (N_9746,N_8368,N_8148);
nor U9747 (N_9747,N_8153,N_8752);
and U9748 (N_9748,N_8659,N_8267);
or U9749 (N_9749,N_8816,N_8223);
xor U9750 (N_9750,N_8132,N_8088);
xnor U9751 (N_9751,N_8717,N_8909);
and U9752 (N_9752,N_8069,N_8994);
and U9753 (N_9753,N_8750,N_8256);
and U9754 (N_9754,N_8881,N_8573);
and U9755 (N_9755,N_8245,N_8843);
nor U9756 (N_9756,N_8318,N_8140);
nor U9757 (N_9757,N_8632,N_8273);
nand U9758 (N_9758,N_8884,N_8015);
xor U9759 (N_9759,N_8776,N_8919);
or U9760 (N_9760,N_8931,N_8332);
and U9761 (N_9761,N_8819,N_8332);
xnor U9762 (N_9762,N_8910,N_8692);
xnor U9763 (N_9763,N_8219,N_8350);
nand U9764 (N_9764,N_8543,N_8104);
and U9765 (N_9765,N_8567,N_8328);
or U9766 (N_9766,N_8509,N_8449);
nor U9767 (N_9767,N_8192,N_8476);
xnor U9768 (N_9768,N_8172,N_8372);
nand U9769 (N_9769,N_8923,N_8988);
or U9770 (N_9770,N_8191,N_8760);
xnor U9771 (N_9771,N_8022,N_8419);
xor U9772 (N_9772,N_8947,N_8175);
and U9773 (N_9773,N_8743,N_8459);
nor U9774 (N_9774,N_8195,N_8393);
or U9775 (N_9775,N_8614,N_8432);
and U9776 (N_9776,N_8595,N_8300);
and U9777 (N_9777,N_8817,N_8234);
nor U9778 (N_9778,N_8425,N_8729);
nand U9779 (N_9779,N_8837,N_8595);
nor U9780 (N_9780,N_8282,N_8440);
nor U9781 (N_9781,N_8128,N_8291);
and U9782 (N_9782,N_8467,N_8875);
nand U9783 (N_9783,N_8903,N_8119);
and U9784 (N_9784,N_8213,N_8385);
and U9785 (N_9785,N_8275,N_8164);
and U9786 (N_9786,N_8331,N_8246);
or U9787 (N_9787,N_8382,N_8151);
nand U9788 (N_9788,N_8836,N_8221);
xor U9789 (N_9789,N_8902,N_8241);
and U9790 (N_9790,N_8588,N_8903);
and U9791 (N_9791,N_8433,N_8582);
nor U9792 (N_9792,N_8310,N_8777);
nand U9793 (N_9793,N_8889,N_8799);
nor U9794 (N_9794,N_8142,N_8412);
or U9795 (N_9795,N_8848,N_8354);
or U9796 (N_9796,N_8008,N_8038);
xnor U9797 (N_9797,N_8971,N_8974);
and U9798 (N_9798,N_8145,N_8698);
or U9799 (N_9799,N_8901,N_8268);
and U9800 (N_9800,N_8437,N_8813);
xor U9801 (N_9801,N_8597,N_8686);
or U9802 (N_9802,N_8146,N_8682);
and U9803 (N_9803,N_8140,N_8369);
or U9804 (N_9804,N_8541,N_8561);
nor U9805 (N_9805,N_8228,N_8624);
nand U9806 (N_9806,N_8928,N_8206);
and U9807 (N_9807,N_8851,N_8091);
xor U9808 (N_9808,N_8231,N_8327);
nor U9809 (N_9809,N_8675,N_8820);
or U9810 (N_9810,N_8294,N_8357);
xnor U9811 (N_9811,N_8932,N_8735);
or U9812 (N_9812,N_8724,N_8812);
nand U9813 (N_9813,N_8434,N_8719);
and U9814 (N_9814,N_8867,N_8468);
xor U9815 (N_9815,N_8283,N_8953);
and U9816 (N_9816,N_8798,N_8996);
nand U9817 (N_9817,N_8716,N_8330);
xnor U9818 (N_9818,N_8167,N_8967);
or U9819 (N_9819,N_8182,N_8039);
nor U9820 (N_9820,N_8370,N_8867);
and U9821 (N_9821,N_8835,N_8072);
nand U9822 (N_9822,N_8809,N_8496);
or U9823 (N_9823,N_8904,N_8010);
xor U9824 (N_9824,N_8413,N_8286);
or U9825 (N_9825,N_8821,N_8940);
xor U9826 (N_9826,N_8472,N_8083);
nor U9827 (N_9827,N_8974,N_8816);
nor U9828 (N_9828,N_8655,N_8871);
or U9829 (N_9829,N_8260,N_8213);
and U9830 (N_9830,N_8958,N_8955);
nand U9831 (N_9831,N_8637,N_8491);
xor U9832 (N_9832,N_8888,N_8297);
nand U9833 (N_9833,N_8851,N_8733);
and U9834 (N_9834,N_8635,N_8407);
xnor U9835 (N_9835,N_8307,N_8276);
xor U9836 (N_9836,N_8321,N_8916);
and U9837 (N_9837,N_8250,N_8706);
and U9838 (N_9838,N_8865,N_8458);
and U9839 (N_9839,N_8179,N_8693);
nor U9840 (N_9840,N_8024,N_8940);
nand U9841 (N_9841,N_8666,N_8022);
xnor U9842 (N_9842,N_8828,N_8296);
or U9843 (N_9843,N_8052,N_8223);
nor U9844 (N_9844,N_8059,N_8702);
or U9845 (N_9845,N_8528,N_8142);
and U9846 (N_9846,N_8042,N_8689);
nand U9847 (N_9847,N_8317,N_8498);
nor U9848 (N_9848,N_8304,N_8167);
or U9849 (N_9849,N_8372,N_8858);
or U9850 (N_9850,N_8800,N_8545);
nor U9851 (N_9851,N_8773,N_8637);
or U9852 (N_9852,N_8694,N_8156);
xor U9853 (N_9853,N_8805,N_8290);
and U9854 (N_9854,N_8408,N_8260);
nor U9855 (N_9855,N_8619,N_8106);
and U9856 (N_9856,N_8561,N_8474);
or U9857 (N_9857,N_8632,N_8787);
nor U9858 (N_9858,N_8719,N_8340);
nand U9859 (N_9859,N_8270,N_8585);
nand U9860 (N_9860,N_8938,N_8699);
and U9861 (N_9861,N_8019,N_8824);
nand U9862 (N_9862,N_8651,N_8572);
xnor U9863 (N_9863,N_8087,N_8266);
nand U9864 (N_9864,N_8946,N_8390);
nand U9865 (N_9865,N_8704,N_8520);
and U9866 (N_9866,N_8453,N_8011);
or U9867 (N_9867,N_8491,N_8433);
nand U9868 (N_9868,N_8968,N_8875);
nand U9869 (N_9869,N_8051,N_8713);
and U9870 (N_9870,N_8954,N_8763);
xnor U9871 (N_9871,N_8885,N_8868);
nand U9872 (N_9872,N_8322,N_8372);
or U9873 (N_9873,N_8255,N_8919);
xnor U9874 (N_9874,N_8387,N_8085);
and U9875 (N_9875,N_8943,N_8203);
and U9876 (N_9876,N_8210,N_8699);
nor U9877 (N_9877,N_8321,N_8205);
nand U9878 (N_9878,N_8716,N_8108);
xnor U9879 (N_9879,N_8424,N_8761);
and U9880 (N_9880,N_8993,N_8031);
and U9881 (N_9881,N_8344,N_8408);
nor U9882 (N_9882,N_8453,N_8603);
nor U9883 (N_9883,N_8055,N_8979);
and U9884 (N_9884,N_8042,N_8381);
nand U9885 (N_9885,N_8863,N_8223);
xor U9886 (N_9886,N_8814,N_8762);
and U9887 (N_9887,N_8578,N_8271);
nor U9888 (N_9888,N_8586,N_8287);
and U9889 (N_9889,N_8292,N_8347);
or U9890 (N_9890,N_8129,N_8267);
and U9891 (N_9891,N_8508,N_8678);
xor U9892 (N_9892,N_8455,N_8672);
xnor U9893 (N_9893,N_8962,N_8931);
xnor U9894 (N_9894,N_8807,N_8601);
nand U9895 (N_9895,N_8460,N_8495);
xor U9896 (N_9896,N_8351,N_8485);
nor U9897 (N_9897,N_8289,N_8090);
xnor U9898 (N_9898,N_8429,N_8560);
and U9899 (N_9899,N_8411,N_8033);
xor U9900 (N_9900,N_8772,N_8574);
or U9901 (N_9901,N_8879,N_8948);
xnor U9902 (N_9902,N_8625,N_8326);
or U9903 (N_9903,N_8244,N_8214);
xor U9904 (N_9904,N_8286,N_8318);
or U9905 (N_9905,N_8754,N_8375);
nor U9906 (N_9906,N_8857,N_8914);
nand U9907 (N_9907,N_8277,N_8198);
nand U9908 (N_9908,N_8842,N_8596);
or U9909 (N_9909,N_8339,N_8641);
and U9910 (N_9910,N_8775,N_8101);
nor U9911 (N_9911,N_8810,N_8961);
xnor U9912 (N_9912,N_8051,N_8293);
xor U9913 (N_9913,N_8484,N_8377);
or U9914 (N_9914,N_8736,N_8302);
nor U9915 (N_9915,N_8109,N_8372);
nor U9916 (N_9916,N_8437,N_8518);
nand U9917 (N_9917,N_8296,N_8747);
and U9918 (N_9918,N_8311,N_8260);
or U9919 (N_9919,N_8476,N_8498);
or U9920 (N_9920,N_8591,N_8239);
and U9921 (N_9921,N_8913,N_8656);
xnor U9922 (N_9922,N_8299,N_8193);
nor U9923 (N_9923,N_8845,N_8403);
nand U9924 (N_9924,N_8343,N_8037);
nor U9925 (N_9925,N_8381,N_8629);
xnor U9926 (N_9926,N_8037,N_8170);
nand U9927 (N_9927,N_8852,N_8321);
or U9928 (N_9928,N_8415,N_8911);
nand U9929 (N_9929,N_8388,N_8103);
xor U9930 (N_9930,N_8847,N_8168);
xnor U9931 (N_9931,N_8037,N_8429);
xnor U9932 (N_9932,N_8985,N_8822);
xor U9933 (N_9933,N_8142,N_8107);
or U9934 (N_9934,N_8055,N_8282);
or U9935 (N_9935,N_8919,N_8288);
and U9936 (N_9936,N_8509,N_8065);
nand U9937 (N_9937,N_8146,N_8988);
and U9938 (N_9938,N_8698,N_8026);
and U9939 (N_9939,N_8329,N_8361);
xor U9940 (N_9940,N_8162,N_8696);
xnor U9941 (N_9941,N_8689,N_8382);
nand U9942 (N_9942,N_8615,N_8141);
and U9943 (N_9943,N_8520,N_8058);
nand U9944 (N_9944,N_8205,N_8700);
or U9945 (N_9945,N_8831,N_8620);
nor U9946 (N_9946,N_8794,N_8179);
nor U9947 (N_9947,N_8015,N_8062);
xor U9948 (N_9948,N_8722,N_8227);
nand U9949 (N_9949,N_8733,N_8659);
nor U9950 (N_9950,N_8178,N_8086);
xor U9951 (N_9951,N_8361,N_8189);
and U9952 (N_9952,N_8622,N_8227);
nand U9953 (N_9953,N_8910,N_8778);
and U9954 (N_9954,N_8232,N_8408);
xnor U9955 (N_9955,N_8526,N_8323);
nor U9956 (N_9956,N_8758,N_8380);
xnor U9957 (N_9957,N_8531,N_8553);
and U9958 (N_9958,N_8146,N_8319);
and U9959 (N_9959,N_8716,N_8553);
or U9960 (N_9960,N_8710,N_8850);
nand U9961 (N_9961,N_8126,N_8151);
and U9962 (N_9962,N_8793,N_8324);
nand U9963 (N_9963,N_8291,N_8300);
nor U9964 (N_9964,N_8158,N_8726);
and U9965 (N_9965,N_8745,N_8560);
xor U9966 (N_9966,N_8290,N_8844);
or U9967 (N_9967,N_8217,N_8870);
and U9968 (N_9968,N_8336,N_8480);
nand U9969 (N_9969,N_8437,N_8805);
nor U9970 (N_9970,N_8737,N_8955);
xnor U9971 (N_9971,N_8676,N_8156);
or U9972 (N_9972,N_8119,N_8398);
nand U9973 (N_9973,N_8346,N_8844);
nand U9974 (N_9974,N_8544,N_8707);
and U9975 (N_9975,N_8666,N_8068);
xor U9976 (N_9976,N_8673,N_8332);
nor U9977 (N_9977,N_8685,N_8364);
or U9978 (N_9978,N_8247,N_8965);
nor U9979 (N_9979,N_8703,N_8366);
nand U9980 (N_9980,N_8127,N_8667);
nor U9981 (N_9981,N_8619,N_8309);
nand U9982 (N_9982,N_8105,N_8489);
xnor U9983 (N_9983,N_8899,N_8382);
and U9984 (N_9984,N_8337,N_8567);
or U9985 (N_9985,N_8607,N_8474);
or U9986 (N_9986,N_8630,N_8417);
nand U9987 (N_9987,N_8904,N_8398);
nand U9988 (N_9988,N_8291,N_8378);
xnor U9989 (N_9989,N_8154,N_8901);
or U9990 (N_9990,N_8246,N_8343);
and U9991 (N_9991,N_8199,N_8531);
xor U9992 (N_9992,N_8718,N_8690);
nor U9993 (N_9993,N_8924,N_8670);
and U9994 (N_9994,N_8572,N_8711);
nand U9995 (N_9995,N_8318,N_8387);
nor U9996 (N_9996,N_8562,N_8084);
nand U9997 (N_9997,N_8768,N_8225);
nand U9998 (N_9998,N_8593,N_8521);
xor U9999 (N_9999,N_8251,N_8324);
and U10000 (N_10000,N_9971,N_9270);
nor U10001 (N_10001,N_9635,N_9380);
xnor U10002 (N_10002,N_9662,N_9758);
xnor U10003 (N_10003,N_9455,N_9894);
or U10004 (N_10004,N_9610,N_9931);
or U10005 (N_10005,N_9210,N_9226);
and U10006 (N_10006,N_9535,N_9554);
and U10007 (N_10007,N_9784,N_9128);
xor U10008 (N_10008,N_9550,N_9006);
nor U10009 (N_10009,N_9812,N_9413);
nor U10010 (N_10010,N_9332,N_9645);
nor U10011 (N_10011,N_9384,N_9239);
or U10012 (N_10012,N_9630,N_9161);
nand U10013 (N_10013,N_9860,N_9268);
and U10014 (N_10014,N_9866,N_9633);
nor U10015 (N_10015,N_9488,N_9793);
xor U10016 (N_10016,N_9598,N_9427);
and U10017 (N_10017,N_9158,N_9277);
xnor U10018 (N_10018,N_9521,N_9743);
and U10019 (N_10019,N_9478,N_9673);
xnor U10020 (N_10020,N_9134,N_9719);
or U10021 (N_10021,N_9555,N_9731);
or U10022 (N_10022,N_9829,N_9467);
xor U10023 (N_10023,N_9573,N_9257);
nor U10024 (N_10024,N_9604,N_9497);
or U10025 (N_10025,N_9648,N_9443);
or U10026 (N_10026,N_9343,N_9863);
nor U10027 (N_10027,N_9964,N_9386);
nor U10028 (N_10028,N_9086,N_9375);
and U10029 (N_10029,N_9755,N_9068);
or U10030 (N_10030,N_9798,N_9563);
nor U10031 (N_10031,N_9523,N_9369);
or U10032 (N_10032,N_9641,N_9877);
or U10033 (N_10033,N_9895,N_9440);
or U10034 (N_10034,N_9490,N_9962);
and U10035 (N_10035,N_9355,N_9241);
xnor U10036 (N_10036,N_9568,N_9791);
and U10037 (N_10037,N_9307,N_9830);
nor U10038 (N_10038,N_9026,N_9833);
xor U10039 (N_10039,N_9152,N_9916);
nor U10040 (N_10040,N_9489,N_9339);
and U10041 (N_10041,N_9388,N_9527);
and U10042 (N_10042,N_9311,N_9501);
or U10043 (N_10043,N_9400,N_9244);
and U10044 (N_10044,N_9363,N_9783);
and U10045 (N_10045,N_9294,N_9750);
xnor U10046 (N_10046,N_9200,N_9148);
and U10047 (N_10047,N_9033,N_9799);
nor U10048 (N_10048,N_9510,N_9898);
nand U10049 (N_10049,N_9892,N_9016);
nor U10050 (N_10050,N_9336,N_9276);
nand U10051 (N_10051,N_9986,N_9441);
xnor U10052 (N_10052,N_9978,N_9144);
and U10053 (N_10053,N_9117,N_9020);
or U10054 (N_10054,N_9350,N_9483);
nand U10055 (N_10055,N_9620,N_9553);
or U10056 (N_10056,N_9428,N_9461);
or U10057 (N_10057,N_9126,N_9147);
and U10058 (N_10058,N_9714,N_9937);
and U10059 (N_10059,N_9544,N_9379);
nor U10060 (N_10060,N_9253,N_9954);
nor U10061 (N_10061,N_9410,N_9782);
and U10062 (N_10062,N_9721,N_9306);
nand U10063 (N_10063,N_9031,N_9372);
xor U10064 (N_10064,N_9974,N_9811);
nand U10065 (N_10065,N_9653,N_9424);
xnor U10066 (N_10066,N_9464,N_9412);
or U10067 (N_10067,N_9319,N_9491);
and U10068 (N_10068,N_9248,N_9957);
and U10069 (N_10069,N_9520,N_9206);
nor U10070 (N_10070,N_9906,N_9001);
nand U10071 (N_10071,N_9768,N_9655);
and U10072 (N_10072,N_9463,N_9110);
xnor U10073 (N_10073,N_9999,N_9063);
nor U10074 (N_10074,N_9274,N_9669);
or U10075 (N_10075,N_9171,N_9847);
nor U10076 (N_10076,N_9718,N_9871);
and U10077 (N_10077,N_9280,N_9909);
or U10078 (N_10078,N_9361,N_9802);
or U10079 (N_10079,N_9968,N_9912);
or U10080 (N_10080,N_9725,N_9227);
nor U10081 (N_10081,N_9426,N_9235);
nor U10082 (N_10082,N_9600,N_9080);
and U10083 (N_10083,N_9220,N_9506);
or U10084 (N_10084,N_9810,N_9159);
nand U10085 (N_10085,N_9449,N_9670);
and U10086 (N_10086,N_9612,N_9228);
nand U10087 (N_10087,N_9136,N_9543);
nand U10088 (N_10088,N_9146,N_9901);
nand U10089 (N_10089,N_9345,N_9558);
or U10090 (N_10090,N_9943,N_9175);
nor U10091 (N_10091,N_9019,N_9591);
nor U10092 (N_10092,N_9278,N_9298);
and U10093 (N_10093,N_9292,N_9177);
nor U10094 (N_10094,N_9611,N_9037);
xnor U10095 (N_10095,N_9756,N_9308);
nand U10096 (N_10096,N_9930,N_9764);
xnor U10097 (N_10097,N_9973,N_9772);
or U10098 (N_10098,N_9524,N_9084);
nand U10099 (N_10099,N_9367,N_9212);
nand U10100 (N_10100,N_9780,N_9649);
or U10101 (N_10101,N_9886,N_9509);
nor U10102 (N_10102,N_9104,N_9472);
or U10103 (N_10103,N_9786,N_9835);
or U10104 (N_10104,N_9823,N_9849);
and U10105 (N_10105,N_9000,N_9541);
or U10106 (N_10106,N_9328,N_9088);
nor U10107 (N_10107,N_9947,N_9806);
and U10108 (N_10108,N_9745,N_9700);
and U10109 (N_10109,N_9221,N_9419);
or U10110 (N_10110,N_9804,N_9879);
xor U10111 (N_10111,N_9751,N_9279);
xor U10112 (N_10112,N_9627,N_9789);
nor U10113 (N_10113,N_9211,N_9317);
and U10114 (N_10114,N_9165,N_9956);
or U10115 (N_10115,N_9862,N_9242);
and U10116 (N_10116,N_9511,N_9095);
xnor U10117 (N_10117,N_9773,N_9851);
or U10118 (N_10118,N_9250,N_9093);
nand U10119 (N_10119,N_9352,N_9138);
and U10120 (N_10120,N_9448,N_9053);
xnor U10121 (N_10121,N_9561,N_9920);
nor U10122 (N_10122,N_9639,N_9284);
nand U10123 (N_10123,N_9264,N_9644);
and U10124 (N_10124,N_9418,N_9011);
xor U10125 (N_10125,N_9106,N_9681);
or U10126 (N_10126,N_9818,N_9403);
nand U10127 (N_10127,N_9321,N_9192);
xnor U10128 (N_10128,N_9251,N_9007);
and U10129 (N_10129,N_9252,N_9907);
nor U10130 (N_10130,N_9888,N_9765);
nor U10131 (N_10131,N_9752,N_9853);
or U10132 (N_10132,N_9097,N_9471);
or U10133 (N_10133,N_9632,N_9434);
xnor U10134 (N_10134,N_9269,N_9980);
nor U10135 (N_10135,N_9243,N_9733);
nor U10136 (N_10136,N_9487,N_9874);
xnor U10137 (N_10137,N_9499,N_9728);
xor U10138 (N_10138,N_9723,N_9651);
and U10139 (N_10139,N_9997,N_9951);
nand U10140 (N_10140,N_9302,N_9364);
xor U10141 (N_10141,N_9392,N_9626);
nand U10142 (N_10142,N_9452,N_9289);
and U10143 (N_10143,N_9163,N_9314);
nor U10144 (N_10144,N_9817,N_9762);
nor U10145 (N_10145,N_9290,N_9625);
nor U10146 (N_10146,N_9405,N_9697);
or U10147 (N_10147,N_9530,N_9111);
or U10148 (N_10148,N_9178,N_9918);
xnor U10149 (N_10149,N_9952,N_9065);
nand U10150 (N_10150,N_9042,N_9771);
nand U10151 (N_10151,N_9942,N_9459);
or U10152 (N_10152,N_9526,N_9120);
nor U10153 (N_10153,N_9323,N_9166);
nor U10154 (N_10154,N_9052,N_9127);
nand U10155 (N_10155,N_9690,N_9621);
and U10156 (N_10156,N_9024,N_9828);
or U10157 (N_10157,N_9469,N_9194);
or U10158 (N_10158,N_9846,N_9987);
and U10159 (N_10159,N_9542,N_9734);
and U10160 (N_10160,N_9593,N_9844);
xnor U10161 (N_10161,N_9606,N_9891);
and U10162 (N_10162,N_9225,N_9688);
or U10163 (N_10163,N_9946,N_9036);
xnor U10164 (N_10164,N_9822,N_9255);
nor U10165 (N_10165,N_9421,N_9528);
nor U10166 (N_10166,N_9614,N_9536);
or U10167 (N_10167,N_9376,N_9503);
xor U10168 (N_10168,N_9186,N_9445);
and U10169 (N_10169,N_9301,N_9949);
or U10170 (N_10170,N_9699,N_9660);
xor U10171 (N_10171,N_9650,N_9291);
xor U10172 (N_10172,N_9601,N_9518);
and U10173 (N_10173,N_9562,N_9236);
xnor U10174 (N_10174,N_9885,N_9961);
or U10175 (N_10175,N_9899,N_9204);
nand U10176 (N_10176,N_9125,N_9083);
and U10177 (N_10177,N_9958,N_9263);
xor U10178 (N_10178,N_9522,N_9816);
nand U10179 (N_10179,N_9131,N_9423);
xor U10180 (N_10180,N_9890,N_9049);
or U10181 (N_10181,N_9840,N_9484);
xor U10182 (N_10182,N_9356,N_9399);
nand U10183 (N_10183,N_9638,N_9800);
xor U10184 (N_10184,N_9139,N_9203);
or U10185 (N_10185,N_9834,N_9201);
and U10186 (N_10186,N_9123,N_9389);
nand U10187 (N_10187,N_9230,N_9991);
and U10188 (N_10188,N_9454,N_9896);
xnor U10189 (N_10189,N_9337,N_9508);
nand U10190 (N_10190,N_9713,N_9826);
xor U10191 (N_10191,N_9303,N_9013);
nand U10192 (N_10192,N_9564,N_9071);
and U10193 (N_10193,N_9922,N_9790);
nand U10194 (N_10194,N_9855,N_9746);
and U10195 (N_10195,N_9893,N_9282);
and U10196 (N_10196,N_9453,N_9470);
or U10197 (N_10197,N_9041,N_9824);
xnor U10198 (N_10198,N_9473,N_9054);
nor U10199 (N_10199,N_9691,N_9658);
xor U10200 (N_10200,N_9034,N_9722);
or U10201 (N_10201,N_9119,N_9371);
nand U10202 (N_10202,N_9950,N_9038);
xor U10203 (N_10203,N_9383,N_9393);
nand U10204 (N_10204,N_9333,N_9229);
xnor U10205 (N_10205,N_9545,N_9602);
nand U10206 (N_10206,N_9836,N_9805);
and U10207 (N_10207,N_9841,N_9603);
nor U10208 (N_10208,N_9061,N_9926);
nor U10209 (N_10209,N_9567,N_9636);
and U10210 (N_10210,N_9348,N_9778);
or U10211 (N_10211,N_9995,N_9374);
or U10212 (N_10212,N_9969,N_9300);
xnor U10213 (N_10213,N_9525,N_9358);
and U10214 (N_10214,N_9397,N_9727);
nand U10215 (N_10215,N_9047,N_9537);
and U10216 (N_10216,N_9223,N_9359);
or U10217 (N_10217,N_9077,N_9992);
nor U10218 (N_10218,N_9797,N_9704);
nand U10219 (N_10219,N_9720,N_9249);
and U10220 (N_10220,N_9378,N_9928);
and U10221 (N_10221,N_9616,N_9776);
nor U10222 (N_10222,N_9096,N_9854);
or U10223 (N_10223,N_9039,N_9316);
or U10224 (N_10224,N_9875,N_9173);
nand U10225 (N_10225,N_9664,N_9135);
nand U10226 (N_10226,N_9759,N_9905);
nor U10227 (N_10227,N_9025,N_9747);
nand U10228 (N_10228,N_9092,N_9945);
nand U10229 (N_10229,N_9266,N_9130);
and U10230 (N_10230,N_9184,N_9654);
nor U10231 (N_10231,N_9507,N_9187);
nand U10232 (N_10232,N_9067,N_9794);
nand U10233 (N_10233,N_9676,N_9100);
xnor U10234 (N_10234,N_9193,N_9787);
nand U10235 (N_10235,N_9792,N_9628);
or U10236 (N_10236,N_9739,N_9556);
nand U10237 (N_10237,N_9565,N_9970);
nor U10238 (N_10238,N_9597,N_9133);
xnor U10239 (N_10239,N_9433,N_9017);
and U10240 (N_10240,N_9740,N_9199);
or U10241 (N_10241,N_9154,N_9517);
or U10242 (N_10242,N_9108,N_9259);
nand U10243 (N_10243,N_9861,N_9996);
nand U10244 (N_10244,N_9458,N_9344);
and U10245 (N_10245,N_9208,N_9760);
xnor U10246 (N_10246,N_9432,N_9021);
and U10247 (N_10247,N_9659,N_9238);
or U10248 (N_10248,N_9195,N_9493);
nor U10249 (N_10249,N_9366,N_9176);
nor U10250 (N_10250,N_9082,N_9105);
and U10251 (N_10251,N_9275,N_9640);
or U10252 (N_10252,N_9587,N_9261);
or U10253 (N_10253,N_9709,N_9420);
and U10254 (N_10254,N_9923,N_9219);
nor U10255 (N_10255,N_9058,N_9647);
and U10256 (N_10256,N_9185,N_9076);
nand U10257 (N_10257,N_9737,N_9028);
or U10258 (N_10258,N_9415,N_9579);
and U10259 (N_10259,N_9103,N_9538);
xnor U10260 (N_10260,N_9354,N_9075);
nor U10261 (N_10261,N_9921,N_9757);
and U10262 (N_10262,N_9619,N_9607);
xnor U10263 (N_10263,N_9113,N_9247);
nor U10264 (N_10264,N_9993,N_9679);
xor U10265 (N_10265,N_9583,N_9581);
or U10266 (N_10266,N_9533,N_9904);
nor U10267 (N_10267,N_9883,N_9590);
nor U10268 (N_10268,N_9532,N_9692);
and U10269 (N_10269,N_9548,N_9057);
or U10270 (N_10270,N_9191,N_9297);
and U10271 (N_10271,N_9258,N_9569);
and U10272 (N_10272,N_9008,N_9570);
and U10273 (N_10273,N_9837,N_9143);
xor U10274 (N_10274,N_9989,N_9205);
xor U10275 (N_10275,N_9324,N_9329);
or U10276 (N_10276,N_9476,N_9051);
and U10277 (N_10277,N_9132,N_9151);
or U10278 (N_10278,N_9761,N_9631);
nor U10279 (N_10279,N_9801,N_9707);
xnor U10280 (N_10280,N_9189,N_9213);
nor U10281 (N_10281,N_9687,N_9234);
and U10282 (N_10282,N_9730,N_9012);
or U10283 (N_10283,N_9486,N_9529);
nand U10284 (N_10284,N_9557,N_9429);
xnor U10285 (N_10285,N_9813,N_9512);
xor U10286 (N_10286,N_9629,N_9450);
nor U10287 (N_10287,N_9754,N_9584);
xnor U10288 (N_10288,N_9142,N_9982);
xnor U10289 (N_10289,N_9078,N_9819);
xor U10290 (N_10290,N_9272,N_9156);
or U10291 (N_10291,N_9140,N_9414);
nor U10292 (N_10292,N_9401,N_9385);
xor U10293 (N_10293,N_9098,N_9781);
nand U10294 (N_10294,N_9137,N_9362);
nand U10295 (N_10295,N_9514,N_9373);
nand U10296 (N_10296,N_9406,N_9404);
nor U10297 (N_10297,N_9665,N_9766);
nand U10298 (N_10298,N_9066,N_9683);
nor U10299 (N_10299,N_9852,N_9929);
nor U10300 (N_10300,N_9674,N_9360);
xnor U10301 (N_10301,N_9122,N_9657);
xor U10302 (N_10302,N_9365,N_9468);
nand U10303 (N_10303,N_9821,N_9677);
and U10304 (N_10304,N_9069,N_9685);
and U10305 (N_10305,N_9305,N_9285);
nand U10306 (N_10306,N_9839,N_9145);
nand U10307 (N_10307,N_9150,N_9504);
or U10308 (N_10308,N_9121,N_9091);
or U10309 (N_10309,N_9157,N_9004);
nor U10310 (N_10310,N_9395,N_9495);
or U10311 (N_10311,N_9288,N_9981);
and U10312 (N_10312,N_9889,N_9900);
and U10313 (N_10313,N_9571,N_9845);
and U10314 (N_10314,N_9182,N_9742);
nor U10315 (N_10315,N_9357,N_9155);
or U10316 (N_10316,N_9966,N_9983);
or U10317 (N_10317,N_9293,N_9589);
nand U10318 (N_10318,N_9202,N_9732);
nand U10319 (N_10319,N_9310,N_9582);
nor U10320 (N_10320,N_9050,N_9624);
nand U10321 (N_10321,N_9064,N_9546);
and U10322 (N_10322,N_9959,N_9387);
nand U10323 (N_10323,N_9796,N_9753);
nor U10324 (N_10324,N_9417,N_9479);
or U10325 (N_10325,N_9035,N_9960);
or U10326 (N_10326,N_9975,N_9435);
nand U10327 (N_10327,N_9169,N_9617);
or U10328 (N_10328,N_9112,N_9578);
and U10329 (N_10329,N_9708,N_9576);
nand U10330 (N_10330,N_9838,N_9595);
nand U10331 (N_10331,N_9903,N_9908);
nor U10332 (N_10332,N_9872,N_9585);
nand U10333 (N_10333,N_9736,N_9304);
and U10334 (N_10334,N_9271,N_9882);
xnor U10335 (N_10335,N_9586,N_9124);
nand U10336 (N_10336,N_9370,N_9513);
xor U10337 (N_10337,N_9820,N_9442);
xnor U10338 (N_10338,N_9869,N_9170);
xnor U10339 (N_10339,N_9174,N_9390);
and U10340 (N_10340,N_9180,N_9197);
xnor U10341 (N_10341,N_9914,N_9808);
nor U10342 (N_10342,N_9646,N_9018);
xor U10343 (N_10343,N_9179,N_9254);
nand U10344 (N_10344,N_9940,N_9976);
and U10345 (N_10345,N_9710,N_9162);
xor U10346 (N_10346,N_9368,N_9726);
nor U10347 (N_10347,N_9224,N_9701);
nor U10348 (N_10348,N_9596,N_9283);
or U10349 (N_10349,N_9560,N_9515);
xor U10350 (N_10350,N_9775,N_9711);
nand U10351 (N_10351,N_9087,N_9850);
xor U10352 (N_10352,N_9325,N_9438);
nand U10353 (N_10353,N_9919,N_9456);
or U10354 (N_10354,N_9539,N_9911);
or U10355 (N_10355,N_9594,N_9643);
nor U10356 (N_10356,N_9897,N_9233);
or U10357 (N_10357,N_9749,N_9474);
nor U10358 (N_10358,N_9827,N_9216);
xor U10359 (N_10359,N_9446,N_9099);
xor U10360 (N_10360,N_9377,N_9972);
xnor U10361 (N_10361,N_9608,N_9618);
nand U10362 (N_10362,N_9313,N_9465);
and U10363 (N_10363,N_9857,N_9622);
or U10364 (N_10364,N_9715,N_9482);
nor U10365 (N_10365,N_9073,N_9196);
or U10366 (N_10366,N_9712,N_9663);
xnor U10367 (N_10367,N_9864,N_9217);
nand U10368 (N_10368,N_9994,N_9580);
xor U10369 (N_10369,N_9101,N_9114);
and U10370 (N_10370,N_9613,N_9656);
nor U10371 (N_10371,N_9689,N_9237);
xnor U10372 (N_10372,N_9858,N_9915);
xor U10373 (N_10373,N_9164,N_9167);
nor U10374 (N_10374,N_9967,N_9118);
nand U10375 (N_10375,N_9927,N_9988);
nand U10376 (N_10376,N_9948,N_9868);
nand U10377 (N_10377,N_9085,N_9215);
or U10378 (N_10378,N_9934,N_9984);
and U10379 (N_10379,N_9190,N_9060);
or U10380 (N_10380,N_9703,N_9462);
xor U10381 (N_10381,N_9494,N_9735);
and U10382 (N_10382,N_9675,N_9309);
and U10383 (N_10383,N_9788,N_9496);
nor U10384 (N_10384,N_9029,N_9777);
or U10385 (N_10385,N_9944,N_9460);
or U10386 (N_10386,N_9925,N_9540);
or U10387 (N_10387,N_9667,N_9843);
or U10388 (N_10388,N_9245,N_9807);
xor U10389 (N_10389,N_9457,N_9141);
xor U10390 (N_10390,N_9661,N_9267);
xor U10391 (N_10391,N_9327,N_9043);
nor U10392 (N_10392,N_9716,N_9382);
nor U10393 (N_10393,N_9634,N_9998);
or U10394 (N_10394,N_9492,N_9881);
nand U10395 (N_10395,N_9695,N_9214);
xor U10396 (N_10396,N_9682,N_9615);
nand U10397 (N_10397,N_9684,N_9402);
and U10398 (N_10398,N_9349,N_9686);
nor U10399 (N_10399,N_9338,N_9265);
xor U10400 (N_10400,N_9048,N_9046);
xnor U10401 (N_10401,N_9519,N_9599);
xnor U10402 (N_10402,N_9027,N_9032);
and U10403 (N_10403,N_9865,N_9502);
and U10404 (N_10404,N_9312,N_9717);
nand U10405 (N_10405,N_9411,N_9870);
xnor U10406 (N_10406,N_9500,N_9209);
nand U10407 (N_10407,N_9430,N_9588);
or U10408 (N_10408,N_9181,N_9936);
xnor U10409 (N_10409,N_9832,N_9040);
or U10410 (N_10410,N_9577,N_9287);
nor U10411 (N_10411,N_9341,N_9022);
or U10412 (N_10412,N_9516,N_9566);
nand U10413 (N_10413,N_9985,N_9741);
xor U10414 (N_10414,N_9055,N_9431);
or U10415 (N_10415,N_9070,N_9391);
nand U10416 (N_10416,N_9637,N_9436);
nand U10417 (N_10417,N_9262,N_9910);
and U10418 (N_10418,N_9416,N_9090);
xor U10419 (N_10419,N_9256,N_9437);
nand U10420 (N_10420,N_9115,N_9842);
nor U10421 (N_10421,N_9102,N_9081);
xnor U10422 (N_10422,N_9814,N_9678);
nor U10423 (N_10423,N_9172,N_9706);
or U10424 (N_10424,N_9698,N_9693);
or U10425 (N_10425,N_9045,N_9398);
nor U10426 (N_10426,N_9666,N_9299);
or U10427 (N_10427,N_9394,N_9009);
nor U10428 (N_10428,N_9409,N_9353);
and U10429 (N_10429,N_9059,N_9062);
or U10430 (N_10430,N_9880,N_9407);
xnor U10431 (N_10431,N_9605,N_9671);
or U10432 (N_10432,N_9825,N_9198);
nand U10433 (N_10433,N_9779,N_9422);
nor U10434 (N_10434,N_9938,N_9340);
xor U10435 (N_10435,N_9246,N_9856);
nand U10436 (N_10436,N_9444,N_9876);
and U10437 (N_10437,N_9466,N_9505);
or U10438 (N_10438,N_9551,N_9315);
nand U10439 (N_10439,N_9342,N_9592);
xnor U10440 (N_10440,N_9873,N_9232);
xnor U10441 (N_10441,N_9222,N_9023);
or U10442 (N_10442,N_9168,N_9335);
nand U10443 (N_10443,N_9439,N_9447);
nor U10444 (N_10444,N_9785,N_9729);
or U10445 (N_10445,N_9748,N_9218);
nand U10446 (N_10446,N_9149,N_9296);
and U10447 (N_10447,N_9153,N_9116);
nor U10448 (N_10448,N_9705,N_9694);
or U10449 (N_10449,N_9326,N_9887);
or U10450 (N_10450,N_9738,N_9953);
nor U10451 (N_10451,N_9322,N_9867);
and U10452 (N_10452,N_9831,N_9260);
nand U10453 (N_10453,N_9079,N_9129);
and U10454 (N_10454,N_9668,N_9498);
and U10455 (N_10455,N_9795,N_9549);
and U10456 (N_10456,N_9330,N_9913);
and U10457 (N_10457,N_9094,N_9044);
and U10458 (N_10458,N_9231,N_9652);
xnor U10459 (N_10459,N_9320,N_9072);
xnor U10460 (N_10460,N_9559,N_9188);
xor U10461 (N_10461,N_9933,N_9769);
nor U10462 (N_10462,N_9425,N_9030);
and U10463 (N_10463,N_9696,N_9346);
nor U10464 (N_10464,N_9941,N_9240);
and U10465 (N_10465,N_9902,N_9878);
nand U10466 (N_10466,N_9408,N_9977);
xor U10467 (N_10467,N_9273,N_9744);
nand U10468 (N_10468,N_9334,N_9109);
or U10469 (N_10469,N_9318,N_9859);
and U10470 (N_10470,N_9680,N_9295);
nand U10471 (N_10471,N_9965,N_9623);
nand U10472 (N_10472,N_9774,N_9574);
xnor U10473 (N_10473,N_9010,N_9534);
nor U10474 (N_10474,N_9160,N_9935);
nor U10475 (N_10475,N_9056,N_9815);
and U10476 (N_10476,N_9107,N_9396);
xnor U10477 (N_10477,N_9979,N_9917);
or U10478 (N_10478,N_9963,N_9074);
or U10479 (N_10479,N_9481,N_9477);
xor U10480 (N_10480,N_9672,N_9331);
or U10481 (N_10481,N_9702,N_9552);
nand U10482 (N_10482,N_9480,N_9015);
or U10483 (N_10483,N_9848,N_9451);
xnor U10484 (N_10484,N_9572,N_9531);
and U10485 (N_10485,N_9351,N_9281);
and U10486 (N_10486,N_9767,N_9183);
xnor U10487 (N_10487,N_9003,N_9575);
or U10488 (N_10488,N_9990,N_9809);
nor U10489 (N_10489,N_9609,N_9955);
xor U10490 (N_10490,N_9286,N_9089);
xor U10491 (N_10491,N_9475,N_9381);
and U10492 (N_10492,N_9002,N_9939);
and U10493 (N_10493,N_9724,N_9924);
nor U10494 (N_10494,N_9642,N_9207);
or U10495 (N_10495,N_9763,N_9770);
nor U10496 (N_10496,N_9005,N_9932);
and U10497 (N_10497,N_9547,N_9803);
xnor U10498 (N_10498,N_9884,N_9014);
xor U10499 (N_10499,N_9485,N_9347);
nor U10500 (N_10500,N_9036,N_9615);
and U10501 (N_10501,N_9717,N_9601);
or U10502 (N_10502,N_9650,N_9488);
and U10503 (N_10503,N_9404,N_9345);
or U10504 (N_10504,N_9889,N_9105);
or U10505 (N_10505,N_9193,N_9200);
or U10506 (N_10506,N_9064,N_9595);
or U10507 (N_10507,N_9834,N_9589);
and U10508 (N_10508,N_9576,N_9401);
nand U10509 (N_10509,N_9886,N_9220);
or U10510 (N_10510,N_9932,N_9575);
or U10511 (N_10511,N_9257,N_9092);
nand U10512 (N_10512,N_9006,N_9470);
nor U10513 (N_10513,N_9344,N_9413);
or U10514 (N_10514,N_9374,N_9828);
xor U10515 (N_10515,N_9695,N_9813);
xor U10516 (N_10516,N_9962,N_9767);
and U10517 (N_10517,N_9113,N_9435);
or U10518 (N_10518,N_9269,N_9662);
nand U10519 (N_10519,N_9661,N_9696);
xnor U10520 (N_10520,N_9126,N_9574);
or U10521 (N_10521,N_9443,N_9707);
nand U10522 (N_10522,N_9488,N_9720);
nand U10523 (N_10523,N_9425,N_9288);
xnor U10524 (N_10524,N_9988,N_9870);
and U10525 (N_10525,N_9127,N_9005);
nor U10526 (N_10526,N_9234,N_9704);
nor U10527 (N_10527,N_9035,N_9469);
or U10528 (N_10528,N_9817,N_9610);
and U10529 (N_10529,N_9830,N_9449);
and U10530 (N_10530,N_9257,N_9582);
xnor U10531 (N_10531,N_9322,N_9433);
xnor U10532 (N_10532,N_9437,N_9929);
nand U10533 (N_10533,N_9643,N_9460);
xor U10534 (N_10534,N_9732,N_9543);
xnor U10535 (N_10535,N_9620,N_9441);
xor U10536 (N_10536,N_9859,N_9282);
nand U10537 (N_10537,N_9570,N_9892);
xnor U10538 (N_10538,N_9475,N_9175);
xor U10539 (N_10539,N_9278,N_9402);
nand U10540 (N_10540,N_9366,N_9941);
xnor U10541 (N_10541,N_9996,N_9634);
xnor U10542 (N_10542,N_9660,N_9760);
nand U10543 (N_10543,N_9378,N_9859);
xor U10544 (N_10544,N_9124,N_9029);
nand U10545 (N_10545,N_9009,N_9384);
xor U10546 (N_10546,N_9424,N_9361);
xnor U10547 (N_10547,N_9740,N_9188);
or U10548 (N_10548,N_9011,N_9008);
nor U10549 (N_10549,N_9468,N_9323);
xnor U10550 (N_10550,N_9741,N_9260);
nor U10551 (N_10551,N_9650,N_9941);
xnor U10552 (N_10552,N_9774,N_9758);
xnor U10553 (N_10553,N_9097,N_9721);
xnor U10554 (N_10554,N_9269,N_9509);
nor U10555 (N_10555,N_9144,N_9142);
xnor U10556 (N_10556,N_9812,N_9794);
and U10557 (N_10557,N_9442,N_9679);
or U10558 (N_10558,N_9787,N_9418);
or U10559 (N_10559,N_9799,N_9039);
nor U10560 (N_10560,N_9035,N_9836);
and U10561 (N_10561,N_9457,N_9369);
or U10562 (N_10562,N_9340,N_9636);
nand U10563 (N_10563,N_9434,N_9246);
xnor U10564 (N_10564,N_9401,N_9134);
xor U10565 (N_10565,N_9468,N_9630);
xnor U10566 (N_10566,N_9135,N_9256);
nor U10567 (N_10567,N_9113,N_9654);
nand U10568 (N_10568,N_9049,N_9530);
and U10569 (N_10569,N_9824,N_9284);
or U10570 (N_10570,N_9453,N_9076);
nand U10571 (N_10571,N_9100,N_9752);
or U10572 (N_10572,N_9604,N_9338);
or U10573 (N_10573,N_9453,N_9239);
nor U10574 (N_10574,N_9327,N_9234);
or U10575 (N_10575,N_9561,N_9221);
or U10576 (N_10576,N_9816,N_9883);
xnor U10577 (N_10577,N_9595,N_9732);
and U10578 (N_10578,N_9257,N_9634);
xnor U10579 (N_10579,N_9277,N_9220);
xor U10580 (N_10580,N_9865,N_9587);
nor U10581 (N_10581,N_9266,N_9850);
nor U10582 (N_10582,N_9135,N_9909);
nand U10583 (N_10583,N_9258,N_9380);
nand U10584 (N_10584,N_9582,N_9468);
nand U10585 (N_10585,N_9101,N_9505);
or U10586 (N_10586,N_9397,N_9723);
nand U10587 (N_10587,N_9899,N_9234);
nand U10588 (N_10588,N_9573,N_9698);
nor U10589 (N_10589,N_9303,N_9518);
and U10590 (N_10590,N_9477,N_9919);
xnor U10591 (N_10591,N_9495,N_9362);
or U10592 (N_10592,N_9042,N_9854);
xor U10593 (N_10593,N_9377,N_9562);
or U10594 (N_10594,N_9545,N_9786);
and U10595 (N_10595,N_9795,N_9264);
xnor U10596 (N_10596,N_9768,N_9805);
nor U10597 (N_10597,N_9211,N_9132);
or U10598 (N_10598,N_9061,N_9100);
nand U10599 (N_10599,N_9750,N_9846);
or U10600 (N_10600,N_9687,N_9302);
nand U10601 (N_10601,N_9775,N_9209);
or U10602 (N_10602,N_9851,N_9324);
and U10603 (N_10603,N_9737,N_9072);
and U10604 (N_10604,N_9360,N_9167);
xor U10605 (N_10605,N_9197,N_9490);
nand U10606 (N_10606,N_9058,N_9587);
nor U10607 (N_10607,N_9550,N_9451);
nand U10608 (N_10608,N_9255,N_9680);
or U10609 (N_10609,N_9417,N_9989);
nand U10610 (N_10610,N_9556,N_9708);
xor U10611 (N_10611,N_9588,N_9916);
nor U10612 (N_10612,N_9515,N_9571);
or U10613 (N_10613,N_9049,N_9714);
and U10614 (N_10614,N_9346,N_9769);
xnor U10615 (N_10615,N_9055,N_9461);
and U10616 (N_10616,N_9000,N_9184);
xnor U10617 (N_10617,N_9778,N_9558);
or U10618 (N_10618,N_9345,N_9909);
or U10619 (N_10619,N_9547,N_9680);
or U10620 (N_10620,N_9506,N_9726);
xnor U10621 (N_10621,N_9595,N_9361);
nand U10622 (N_10622,N_9952,N_9867);
xnor U10623 (N_10623,N_9296,N_9151);
or U10624 (N_10624,N_9217,N_9691);
and U10625 (N_10625,N_9723,N_9852);
nor U10626 (N_10626,N_9613,N_9376);
or U10627 (N_10627,N_9430,N_9745);
nor U10628 (N_10628,N_9760,N_9056);
and U10629 (N_10629,N_9198,N_9386);
nand U10630 (N_10630,N_9519,N_9455);
nand U10631 (N_10631,N_9002,N_9178);
nor U10632 (N_10632,N_9169,N_9145);
xor U10633 (N_10633,N_9069,N_9825);
and U10634 (N_10634,N_9990,N_9249);
nand U10635 (N_10635,N_9471,N_9617);
xor U10636 (N_10636,N_9576,N_9507);
or U10637 (N_10637,N_9179,N_9143);
or U10638 (N_10638,N_9257,N_9985);
or U10639 (N_10639,N_9533,N_9228);
or U10640 (N_10640,N_9002,N_9225);
and U10641 (N_10641,N_9421,N_9125);
nand U10642 (N_10642,N_9609,N_9155);
or U10643 (N_10643,N_9021,N_9445);
and U10644 (N_10644,N_9693,N_9315);
nor U10645 (N_10645,N_9690,N_9984);
nand U10646 (N_10646,N_9759,N_9610);
nor U10647 (N_10647,N_9232,N_9063);
nand U10648 (N_10648,N_9215,N_9782);
or U10649 (N_10649,N_9163,N_9011);
nor U10650 (N_10650,N_9564,N_9690);
nor U10651 (N_10651,N_9131,N_9998);
or U10652 (N_10652,N_9473,N_9116);
nor U10653 (N_10653,N_9069,N_9496);
nand U10654 (N_10654,N_9168,N_9552);
or U10655 (N_10655,N_9511,N_9163);
and U10656 (N_10656,N_9571,N_9337);
nand U10657 (N_10657,N_9534,N_9061);
and U10658 (N_10658,N_9008,N_9064);
or U10659 (N_10659,N_9915,N_9537);
or U10660 (N_10660,N_9231,N_9528);
and U10661 (N_10661,N_9664,N_9405);
and U10662 (N_10662,N_9502,N_9668);
xor U10663 (N_10663,N_9964,N_9137);
and U10664 (N_10664,N_9115,N_9368);
and U10665 (N_10665,N_9633,N_9290);
or U10666 (N_10666,N_9066,N_9875);
nand U10667 (N_10667,N_9370,N_9393);
or U10668 (N_10668,N_9768,N_9750);
nor U10669 (N_10669,N_9562,N_9456);
nand U10670 (N_10670,N_9821,N_9793);
nor U10671 (N_10671,N_9684,N_9718);
and U10672 (N_10672,N_9915,N_9003);
or U10673 (N_10673,N_9060,N_9216);
nand U10674 (N_10674,N_9237,N_9907);
nand U10675 (N_10675,N_9767,N_9656);
xor U10676 (N_10676,N_9024,N_9366);
xnor U10677 (N_10677,N_9661,N_9063);
or U10678 (N_10678,N_9092,N_9808);
nand U10679 (N_10679,N_9371,N_9128);
xnor U10680 (N_10680,N_9367,N_9900);
xor U10681 (N_10681,N_9195,N_9459);
nor U10682 (N_10682,N_9637,N_9739);
nand U10683 (N_10683,N_9317,N_9993);
and U10684 (N_10684,N_9126,N_9367);
or U10685 (N_10685,N_9102,N_9612);
nand U10686 (N_10686,N_9760,N_9848);
and U10687 (N_10687,N_9398,N_9844);
or U10688 (N_10688,N_9972,N_9948);
nor U10689 (N_10689,N_9373,N_9045);
or U10690 (N_10690,N_9427,N_9786);
nor U10691 (N_10691,N_9559,N_9071);
nor U10692 (N_10692,N_9401,N_9273);
nor U10693 (N_10693,N_9771,N_9776);
nor U10694 (N_10694,N_9733,N_9810);
and U10695 (N_10695,N_9487,N_9737);
or U10696 (N_10696,N_9407,N_9402);
and U10697 (N_10697,N_9022,N_9534);
nand U10698 (N_10698,N_9274,N_9949);
nor U10699 (N_10699,N_9787,N_9241);
xor U10700 (N_10700,N_9774,N_9276);
nand U10701 (N_10701,N_9091,N_9142);
and U10702 (N_10702,N_9241,N_9818);
xor U10703 (N_10703,N_9534,N_9851);
nor U10704 (N_10704,N_9975,N_9385);
or U10705 (N_10705,N_9678,N_9006);
xnor U10706 (N_10706,N_9032,N_9373);
xor U10707 (N_10707,N_9680,N_9309);
and U10708 (N_10708,N_9333,N_9701);
or U10709 (N_10709,N_9647,N_9808);
nor U10710 (N_10710,N_9245,N_9586);
nor U10711 (N_10711,N_9678,N_9285);
xnor U10712 (N_10712,N_9105,N_9917);
nand U10713 (N_10713,N_9262,N_9522);
nand U10714 (N_10714,N_9160,N_9622);
and U10715 (N_10715,N_9070,N_9035);
nor U10716 (N_10716,N_9096,N_9486);
xor U10717 (N_10717,N_9404,N_9303);
or U10718 (N_10718,N_9102,N_9588);
nor U10719 (N_10719,N_9302,N_9690);
nor U10720 (N_10720,N_9513,N_9589);
nor U10721 (N_10721,N_9646,N_9641);
xor U10722 (N_10722,N_9948,N_9896);
xor U10723 (N_10723,N_9857,N_9704);
nor U10724 (N_10724,N_9069,N_9608);
or U10725 (N_10725,N_9992,N_9481);
xor U10726 (N_10726,N_9202,N_9354);
or U10727 (N_10727,N_9023,N_9638);
and U10728 (N_10728,N_9038,N_9216);
or U10729 (N_10729,N_9446,N_9359);
nor U10730 (N_10730,N_9229,N_9902);
and U10731 (N_10731,N_9447,N_9284);
or U10732 (N_10732,N_9486,N_9548);
nand U10733 (N_10733,N_9567,N_9452);
nand U10734 (N_10734,N_9491,N_9853);
xor U10735 (N_10735,N_9880,N_9508);
nor U10736 (N_10736,N_9095,N_9984);
and U10737 (N_10737,N_9560,N_9448);
or U10738 (N_10738,N_9352,N_9802);
nor U10739 (N_10739,N_9855,N_9766);
xor U10740 (N_10740,N_9281,N_9543);
nor U10741 (N_10741,N_9049,N_9210);
nor U10742 (N_10742,N_9353,N_9577);
xor U10743 (N_10743,N_9053,N_9682);
nand U10744 (N_10744,N_9092,N_9911);
and U10745 (N_10745,N_9934,N_9504);
xnor U10746 (N_10746,N_9374,N_9839);
or U10747 (N_10747,N_9737,N_9272);
nor U10748 (N_10748,N_9534,N_9295);
and U10749 (N_10749,N_9911,N_9892);
xnor U10750 (N_10750,N_9824,N_9858);
and U10751 (N_10751,N_9659,N_9143);
xor U10752 (N_10752,N_9862,N_9145);
xor U10753 (N_10753,N_9794,N_9420);
or U10754 (N_10754,N_9832,N_9696);
nor U10755 (N_10755,N_9562,N_9398);
xnor U10756 (N_10756,N_9690,N_9805);
nor U10757 (N_10757,N_9181,N_9177);
and U10758 (N_10758,N_9106,N_9552);
or U10759 (N_10759,N_9899,N_9146);
xor U10760 (N_10760,N_9627,N_9309);
nor U10761 (N_10761,N_9178,N_9731);
nand U10762 (N_10762,N_9040,N_9263);
xnor U10763 (N_10763,N_9253,N_9471);
nand U10764 (N_10764,N_9980,N_9590);
and U10765 (N_10765,N_9871,N_9687);
nor U10766 (N_10766,N_9350,N_9781);
and U10767 (N_10767,N_9926,N_9281);
nor U10768 (N_10768,N_9647,N_9406);
nand U10769 (N_10769,N_9789,N_9329);
or U10770 (N_10770,N_9273,N_9823);
nor U10771 (N_10771,N_9969,N_9410);
and U10772 (N_10772,N_9377,N_9293);
and U10773 (N_10773,N_9491,N_9958);
xnor U10774 (N_10774,N_9852,N_9194);
and U10775 (N_10775,N_9145,N_9683);
nand U10776 (N_10776,N_9292,N_9588);
and U10777 (N_10777,N_9546,N_9537);
or U10778 (N_10778,N_9178,N_9754);
xor U10779 (N_10779,N_9215,N_9339);
and U10780 (N_10780,N_9801,N_9053);
nor U10781 (N_10781,N_9575,N_9796);
nor U10782 (N_10782,N_9267,N_9046);
nand U10783 (N_10783,N_9562,N_9828);
nand U10784 (N_10784,N_9103,N_9416);
and U10785 (N_10785,N_9072,N_9123);
nand U10786 (N_10786,N_9847,N_9831);
or U10787 (N_10787,N_9968,N_9377);
nand U10788 (N_10788,N_9508,N_9910);
xnor U10789 (N_10789,N_9555,N_9051);
or U10790 (N_10790,N_9742,N_9940);
and U10791 (N_10791,N_9707,N_9397);
or U10792 (N_10792,N_9068,N_9815);
and U10793 (N_10793,N_9672,N_9690);
nand U10794 (N_10794,N_9717,N_9880);
nand U10795 (N_10795,N_9753,N_9333);
nand U10796 (N_10796,N_9423,N_9816);
nand U10797 (N_10797,N_9139,N_9644);
nand U10798 (N_10798,N_9622,N_9421);
xor U10799 (N_10799,N_9755,N_9678);
or U10800 (N_10800,N_9294,N_9797);
and U10801 (N_10801,N_9684,N_9846);
nand U10802 (N_10802,N_9017,N_9315);
or U10803 (N_10803,N_9247,N_9606);
and U10804 (N_10804,N_9943,N_9488);
and U10805 (N_10805,N_9874,N_9866);
or U10806 (N_10806,N_9907,N_9712);
or U10807 (N_10807,N_9376,N_9184);
and U10808 (N_10808,N_9455,N_9591);
nand U10809 (N_10809,N_9992,N_9741);
and U10810 (N_10810,N_9378,N_9553);
nor U10811 (N_10811,N_9557,N_9508);
or U10812 (N_10812,N_9987,N_9091);
and U10813 (N_10813,N_9940,N_9082);
or U10814 (N_10814,N_9112,N_9062);
nor U10815 (N_10815,N_9335,N_9477);
and U10816 (N_10816,N_9603,N_9586);
or U10817 (N_10817,N_9803,N_9634);
and U10818 (N_10818,N_9212,N_9479);
xor U10819 (N_10819,N_9474,N_9104);
nand U10820 (N_10820,N_9088,N_9205);
and U10821 (N_10821,N_9185,N_9653);
or U10822 (N_10822,N_9963,N_9621);
nand U10823 (N_10823,N_9212,N_9577);
xnor U10824 (N_10824,N_9787,N_9653);
nand U10825 (N_10825,N_9220,N_9463);
xor U10826 (N_10826,N_9148,N_9797);
xnor U10827 (N_10827,N_9790,N_9454);
and U10828 (N_10828,N_9923,N_9085);
nand U10829 (N_10829,N_9979,N_9683);
xor U10830 (N_10830,N_9021,N_9429);
and U10831 (N_10831,N_9449,N_9861);
or U10832 (N_10832,N_9166,N_9321);
and U10833 (N_10833,N_9280,N_9629);
nor U10834 (N_10834,N_9957,N_9125);
xor U10835 (N_10835,N_9211,N_9270);
or U10836 (N_10836,N_9169,N_9146);
xor U10837 (N_10837,N_9788,N_9143);
nand U10838 (N_10838,N_9924,N_9228);
nor U10839 (N_10839,N_9823,N_9298);
nand U10840 (N_10840,N_9870,N_9684);
and U10841 (N_10841,N_9058,N_9989);
or U10842 (N_10842,N_9655,N_9384);
or U10843 (N_10843,N_9124,N_9882);
nor U10844 (N_10844,N_9383,N_9258);
xor U10845 (N_10845,N_9153,N_9648);
and U10846 (N_10846,N_9088,N_9661);
and U10847 (N_10847,N_9916,N_9339);
and U10848 (N_10848,N_9391,N_9130);
xnor U10849 (N_10849,N_9328,N_9080);
nor U10850 (N_10850,N_9783,N_9447);
nand U10851 (N_10851,N_9153,N_9666);
nor U10852 (N_10852,N_9222,N_9425);
xor U10853 (N_10853,N_9844,N_9599);
nand U10854 (N_10854,N_9239,N_9805);
xor U10855 (N_10855,N_9778,N_9005);
nor U10856 (N_10856,N_9435,N_9045);
nand U10857 (N_10857,N_9689,N_9710);
nand U10858 (N_10858,N_9404,N_9619);
and U10859 (N_10859,N_9120,N_9255);
nor U10860 (N_10860,N_9096,N_9880);
nor U10861 (N_10861,N_9063,N_9773);
xnor U10862 (N_10862,N_9866,N_9776);
nand U10863 (N_10863,N_9850,N_9250);
and U10864 (N_10864,N_9731,N_9067);
nor U10865 (N_10865,N_9011,N_9704);
or U10866 (N_10866,N_9158,N_9297);
nor U10867 (N_10867,N_9611,N_9570);
nor U10868 (N_10868,N_9838,N_9550);
or U10869 (N_10869,N_9602,N_9057);
xnor U10870 (N_10870,N_9912,N_9369);
or U10871 (N_10871,N_9210,N_9983);
nor U10872 (N_10872,N_9794,N_9593);
and U10873 (N_10873,N_9069,N_9543);
nor U10874 (N_10874,N_9332,N_9658);
nor U10875 (N_10875,N_9962,N_9470);
xnor U10876 (N_10876,N_9184,N_9232);
nand U10877 (N_10877,N_9331,N_9682);
nand U10878 (N_10878,N_9329,N_9166);
or U10879 (N_10879,N_9265,N_9411);
nand U10880 (N_10880,N_9163,N_9130);
xor U10881 (N_10881,N_9808,N_9530);
or U10882 (N_10882,N_9138,N_9914);
and U10883 (N_10883,N_9891,N_9875);
xor U10884 (N_10884,N_9854,N_9822);
and U10885 (N_10885,N_9729,N_9689);
nor U10886 (N_10886,N_9427,N_9711);
nor U10887 (N_10887,N_9442,N_9374);
and U10888 (N_10888,N_9017,N_9910);
nor U10889 (N_10889,N_9078,N_9884);
or U10890 (N_10890,N_9660,N_9261);
nor U10891 (N_10891,N_9042,N_9359);
nor U10892 (N_10892,N_9800,N_9030);
xor U10893 (N_10893,N_9280,N_9648);
or U10894 (N_10894,N_9330,N_9487);
nor U10895 (N_10895,N_9395,N_9854);
nor U10896 (N_10896,N_9120,N_9681);
nand U10897 (N_10897,N_9496,N_9981);
nand U10898 (N_10898,N_9004,N_9020);
xnor U10899 (N_10899,N_9243,N_9277);
and U10900 (N_10900,N_9317,N_9729);
or U10901 (N_10901,N_9090,N_9657);
or U10902 (N_10902,N_9159,N_9007);
xor U10903 (N_10903,N_9871,N_9549);
or U10904 (N_10904,N_9174,N_9070);
or U10905 (N_10905,N_9253,N_9249);
or U10906 (N_10906,N_9729,N_9046);
or U10907 (N_10907,N_9871,N_9700);
xor U10908 (N_10908,N_9052,N_9712);
or U10909 (N_10909,N_9356,N_9059);
xor U10910 (N_10910,N_9894,N_9246);
and U10911 (N_10911,N_9764,N_9741);
nand U10912 (N_10912,N_9125,N_9742);
nor U10913 (N_10913,N_9714,N_9828);
xor U10914 (N_10914,N_9713,N_9012);
nand U10915 (N_10915,N_9889,N_9295);
nand U10916 (N_10916,N_9948,N_9370);
nand U10917 (N_10917,N_9656,N_9020);
nand U10918 (N_10918,N_9477,N_9406);
or U10919 (N_10919,N_9280,N_9994);
nor U10920 (N_10920,N_9362,N_9903);
or U10921 (N_10921,N_9368,N_9875);
nand U10922 (N_10922,N_9292,N_9199);
nand U10923 (N_10923,N_9414,N_9840);
or U10924 (N_10924,N_9293,N_9998);
xnor U10925 (N_10925,N_9496,N_9470);
nand U10926 (N_10926,N_9220,N_9608);
nand U10927 (N_10927,N_9062,N_9218);
and U10928 (N_10928,N_9904,N_9057);
or U10929 (N_10929,N_9376,N_9285);
or U10930 (N_10930,N_9920,N_9600);
or U10931 (N_10931,N_9702,N_9591);
nand U10932 (N_10932,N_9873,N_9205);
and U10933 (N_10933,N_9332,N_9088);
and U10934 (N_10934,N_9005,N_9444);
or U10935 (N_10935,N_9494,N_9882);
or U10936 (N_10936,N_9476,N_9340);
and U10937 (N_10937,N_9835,N_9452);
nand U10938 (N_10938,N_9143,N_9797);
xnor U10939 (N_10939,N_9159,N_9125);
or U10940 (N_10940,N_9385,N_9314);
xor U10941 (N_10941,N_9740,N_9253);
or U10942 (N_10942,N_9617,N_9812);
nor U10943 (N_10943,N_9016,N_9941);
or U10944 (N_10944,N_9916,N_9633);
xor U10945 (N_10945,N_9227,N_9072);
nor U10946 (N_10946,N_9106,N_9095);
nand U10947 (N_10947,N_9901,N_9301);
nor U10948 (N_10948,N_9117,N_9517);
nor U10949 (N_10949,N_9622,N_9765);
nand U10950 (N_10950,N_9874,N_9031);
and U10951 (N_10951,N_9794,N_9129);
xnor U10952 (N_10952,N_9750,N_9979);
or U10953 (N_10953,N_9427,N_9189);
xor U10954 (N_10954,N_9347,N_9968);
or U10955 (N_10955,N_9530,N_9776);
or U10956 (N_10956,N_9829,N_9658);
and U10957 (N_10957,N_9877,N_9866);
nand U10958 (N_10958,N_9678,N_9073);
or U10959 (N_10959,N_9136,N_9187);
xnor U10960 (N_10960,N_9729,N_9191);
xnor U10961 (N_10961,N_9236,N_9099);
nor U10962 (N_10962,N_9442,N_9756);
nand U10963 (N_10963,N_9912,N_9220);
or U10964 (N_10964,N_9593,N_9789);
and U10965 (N_10965,N_9707,N_9008);
nor U10966 (N_10966,N_9362,N_9780);
xor U10967 (N_10967,N_9690,N_9375);
and U10968 (N_10968,N_9011,N_9259);
or U10969 (N_10969,N_9776,N_9568);
and U10970 (N_10970,N_9881,N_9675);
or U10971 (N_10971,N_9212,N_9415);
xor U10972 (N_10972,N_9132,N_9470);
or U10973 (N_10973,N_9431,N_9075);
and U10974 (N_10974,N_9666,N_9983);
or U10975 (N_10975,N_9830,N_9340);
nand U10976 (N_10976,N_9645,N_9613);
and U10977 (N_10977,N_9043,N_9417);
nor U10978 (N_10978,N_9074,N_9458);
nand U10979 (N_10979,N_9355,N_9296);
xor U10980 (N_10980,N_9363,N_9472);
nor U10981 (N_10981,N_9925,N_9839);
nor U10982 (N_10982,N_9474,N_9456);
and U10983 (N_10983,N_9415,N_9408);
xnor U10984 (N_10984,N_9415,N_9351);
or U10985 (N_10985,N_9162,N_9241);
and U10986 (N_10986,N_9026,N_9106);
xnor U10987 (N_10987,N_9470,N_9187);
xor U10988 (N_10988,N_9759,N_9039);
or U10989 (N_10989,N_9255,N_9665);
nand U10990 (N_10990,N_9717,N_9120);
nand U10991 (N_10991,N_9361,N_9661);
nand U10992 (N_10992,N_9649,N_9549);
nor U10993 (N_10993,N_9642,N_9578);
xnor U10994 (N_10994,N_9082,N_9123);
xor U10995 (N_10995,N_9879,N_9333);
and U10996 (N_10996,N_9859,N_9498);
nor U10997 (N_10997,N_9755,N_9603);
xor U10998 (N_10998,N_9510,N_9388);
xor U10999 (N_10999,N_9980,N_9387);
and U11000 (N_11000,N_10785,N_10157);
and U11001 (N_11001,N_10675,N_10091);
xnor U11002 (N_11002,N_10196,N_10579);
nor U11003 (N_11003,N_10549,N_10138);
nand U11004 (N_11004,N_10683,N_10954);
nor U11005 (N_11005,N_10655,N_10871);
and U11006 (N_11006,N_10458,N_10709);
nor U11007 (N_11007,N_10797,N_10321);
and U11008 (N_11008,N_10914,N_10996);
or U11009 (N_11009,N_10092,N_10127);
xnor U11010 (N_11010,N_10231,N_10448);
nand U11011 (N_11011,N_10897,N_10434);
nor U11012 (N_11012,N_10457,N_10776);
nand U11013 (N_11013,N_10386,N_10372);
xnor U11014 (N_11014,N_10242,N_10309);
xor U11015 (N_11015,N_10789,N_10481);
xnor U11016 (N_11016,N_10719,N_10819);
nor U11017 (N_11017,N_10426,N_10322);
nor U11018 (N_11018,N_10454,N_10652);
and U11019 (N_11019,N_10404,N_10112);
nor U11020 (N_11020,N_10220,N_10204);
and U11021 (N_11021,N_10915,N_10432);
nor U11022 (N_11022,N_10031,N_10739);
or U11023 (N_11023,N_10574,N_10088);
xnor U11024 (N_11024,N_10859,N_10937);
or U11025 (N_11025,N_10317,N_10491);
or U11026 (N_11026,N_10810,N_10995);
and U11027 (N_11027,N_10017,N_10000);
nor U11028 (N_11028,N_10382,N_10496);
xor U11029 (N_11029,N_10557,N_10755);
and U11030 (N_11030,N_10668,N_10944);
and U11031 (N_11031,N_10994,N_10538);
and U11032 (N_11032,N_10534,N_10703);
xnor U11033 (N_11033,N_10613,N_10854);
xnor U11034 (N_11034,N_10406,N_10616);
nand U11035 (N_11035,N_10069,N_10330);
nand U11036 (N_11036,N_10985,N_10723);
or U11037 (N_11037,N_10378,N_10158);
nand U11038 (N_11038,N_10941,N_10990);
xor U11039 (N_11039,N_10485,N_10249);
nor U11040 (N_11040,N_10548,N_10680);
xnor U11041 (N_11041,N_10277,N_10794);
and U11042 (N_11042,N_10521,N_10877);
and U11043 (N_11043,N_10296,N_10353);
xnor U11044 (N_11044,N_10949,N_10495);
or U11045 (N_11045,N_10352,N_10388);
xnor U11046 (N_11046,N_10621,N_10326);
or U11047 (N_11047,N_10649,N_10377);
and U11048 (N_11048,N_10608,N_10441);
xor U11049 (N_11049,N_10141,N_10498);
and U11050 (N_11050,N_10051,N_10181);
nand U11051 (N_11051,N_10007,N_10325);
nand U11052 (N_11052,N_10427,N_10639);
nand U11053 (N_11053,N_10962,N_10023);
xnor U11054 (N_11054,N_10612,N_10173);
or U11055 (N_11055,N_10053,N_10615);
nor U11056 (N_11056,N_10700,N_10757);
nor U11057 (N_11057,N_10407,N_10845);
nor U11058 (N_11058,N_10115,N_10487);
nand U11059 (N_11059,N_10447,N_10518);
nand U11060 (N_11060,N_10836,N_10967);
nand U11061 (N_11061,N_10024,N_10264);
and U11062 (N_11062,N_10738,N_10812);
and U11063 (N_11063,N_10437,N_10917);
and U11064 (N_11064,N_10807,N_10759);
nor U11065 (N_11065,N_10626,N_10133);
xnor U11066 (N_11066,N_10813,N_10455);
or U11067 (N_11067,N_10188,N_10278);
nor U11068 (N_11068,N_10423,N_10113);
and U11069 (N_11069,N_10106,N_10525);
and U11070 (N_11070,N_10623,N_10085);
nor U11071 (N_11071,N_10934,N_10908);
xor U11072 (N_11072,N_10957,N_10839);
xnor U11073 (N_11073,N_10241,N_10906);
xnor U11074 (N_11074,N_10150,N_10499);
nor U11075 (N_11075,N_10004,N_10850);
xnor U11076 (N_11076,N_10578,N_10860);
or U11077 (N_11077,N_10068,N_10136);
nand U11078 (N_11078,N_10603,N_10258);
or U11079 (N_11079,N_10771,N_10054);
or U11080 (N_11080,N_10885,N_10919);
xor U11081 (N_11081,N_10236,N_10778);
nor U11082 (N_11082,N_10893,N_10540);
nor U11083 (N_11083,N_10275,N_10791);
nor U11084 (N_11084,N_10357,N_10572);
nor U11085 (N_11085,N_10311,N_10001);
nand U11086 (N_11086,N_10130,N_10698);
and U11087 (N_11087,N_10730,N_10878);
or U11088 (N_11088,N_10966,N_10095);
and U11089 (N_11089,N_10899,N_10562);
or U11090 (N_11090,N_10126,N_10254);
xnor U11091 (N_11091,N_10537,N_10221);
or U11092 (N_11092,N_10561,N_10560);
nor U11093 (N_11093,N_10660,N_10940);
and U11094 (N_11094,N_10167,N_10370);
xor U11095 (N_11095,N_10600,N_10299);
or U11096 (N_11096,N_10033,N_10667);
nand U11097 (N_11097,N_10255,N_10857);
or U11098 (N_11098,N_10619,N_10520);
xnor U11099 (N_11099,N_10070,N_10291);
or U11100 (N_11100,N_10341,N_10036);
nand U11101 (N_11101,N_10425,N_10882);
nand U11102 (N_11102,N_10705,N_10013);
xor U11103 (N_11103,N_10643,N_10171);
xor U11104 (N_11104,N_10656,N_10592);
nor U11105 (N_11105,N_10333,N_10380);
or U11106 (N_11106,N_10864,N_10714);
nor U11107 (N_11107,N_10782,N_10064);
or U11108 (N_11108,N_10488,N_10856);
and U11109 (N_11109,N_10222,N_10773);
or U11110 (N_11110,N_10156,N_10065);
xor U11111 (N_11111,N_10722,N_10933);
xor U11112 (N_11112,N_10516,N_10635);
nand U11113 (N_11113,N_10246,N_10411);
nand U11114 (N_11114,N_10227,N_10984);
or U11115 (N_11115,N_10076,N_10170);
nand U11116 (N_11116,N_10169,N_10465);
nand U11117 (N_11117,N_10048,N_10559);
nor U11118 (N_11118,N_10852,N_10148);
and U11119 (N_11119,N_10315,N_10712);
and U11120 (N_11120,N_10783,N_10294);
and U11121 (N_11121,N_10997,N_10664);
or U11122 (N_11122,N_10651,N_10345);
or U11123 (N_11123,N_10861,N_10636);
or U11124 (N_11124,N_10690,N_10213);
and U11125 (N_11125,N_10030,N_10617);
or U11126 (N_11126,N_10653,N_10466);
nand U11127 (N_11127,N_10252,N_10981);
nand U11128 (N_11128,N_10260,N_10887);
and U11129 (N_11129,N_10346,N_10201);
or U11130 (N_11130,N_10618,N_10329);
and U11131 (N_11131,N_10901,N_10266);
xnor U11132 (N_11132,N_10314,N_10038);
or U11133 (N_11133,N_10970,N_10866);
nand U11134 (N_11134,N_10039,N_10144);
and U11135 (N_11135,N_10025,N_10847);
or U11136 (N_11136,N_10890,N_10788);
nand U11137 (N_11137,N_10977,N_10134);
nor U11138 (N_11138,N_10119,N_10565);
or U11139 (N_11139,N_10253,N_10508);
or U11140 (N_11140,N_10176,N_10584);
xor U11141 (N_11141,N_10986,N_10486);
and U11142 (N_11142,N_10028,N_10591);
xor U11143 (N_11143,N_10539,N_10910);
nand U11144 (N_11144,N_10318,N_10765);
and U11145 (N_11145,N_10973,N_10998);
or U11146 (N_11146,N_10100,N_10964);
and U11147 (N_11147,N_10456,N_10146);
or U11148 (N_11148,N_10390,N_10762);
or U11149 (N_11149,N_10745,N_10638);
and U11150 (N_11150,N_10531,N_10831);
or U11151 (N_11151,N_10165,N_10989);
or U11152 (N_11152,N_10582,N_10809);
or U11153 (N_11153,N_10546,N_10245);
nor U11154 (N_11154,N_10558,N_10452);
and U11155 (N_11155,N_10935,N_10728);
and U11156 (N_11156,N_10524,N_10737);
and U11157 (N_11157,N_10770,N_10784);
or U11158 (N_11158,N_10029,N_10371);
xor U11159 (N_11159,N_10210,N_10014);
nand U11160 (N_11160,N_10681,N_10725);
xor U11161 (N_11161,N_10803,N_10695);
or U11162 (N_11162,N_10373,N_10056);
or U11163 (N_11163,N_10567,N_10350);
or U11164 (N_11164,N_10946,N_10354);
and U11165 (N_11165,N_10568,N_10889);
xor U11166 (N_11166,N_10153,N_10238);
nor U11167 (N_11167,N_10356,N_10472);
or U11168 (N_11168,N_10470,N_10290);
nand U11169 (N_11169,N_10775,N_10987);
nand U11170 (N_11170,N_10936,N_10827);
or U11171 (N_11171,N_10921,N_10976);
nand U11172 (N_11172,N_10177,N_10876);
xor U11173 (N_11173,N_10162,N_10554);
nor U11174 (N_11174,N_10159,N_10147);
nand U11175 (N_11175,N_10049,N_10713);
nor U11176 (N_11176,N_10547,N_10331);
nand U11177 (N_11177,N_10172,N_10405);
nand U11178 (N_11178,N_10428,N_10895);
nor U11179 (N_11179,N_10978,N_10818);
nor U11180 (N_11180,N_10610,N_10927);
or U11181 (N_11181,N_10523,N_10923);
nor U11182 (N_11182,N_10402,N_10756);
and U11183 (N_11183,N_10323,N_10109);
nor U11184 (N_11184,N_10896,N_10080);
or U11185 (N_11185,N_10689,N_10436);
nor U11186 (N_11186,N_10090,N_10197);
nand U11187 (N_11187,N_10573,N_10760);
nand U11188 (N_11188,N_10273,N_10606);
and U11189 (N_11189,N_10032,N_10505);
nor U11190 (N_11190,N_10155,N_10805);
or U11191 (N_11191,N_10189,N_10431);
nor U11192 (N_11192,N_10504,N_10947);
xor U11193 (N_11193,N_10293,N_10974);
nor U11194 (N_11194,N_10796,N_10037);
nand U11195 (N_11195,N_10175,N_10217);
or U11196 (N_11196,N_10682,N_10830);
xnor U11197 (N_11197,N_10289,N_10611);
xor U11198 (N_11198,N_10424,N_10892);
xor U11199 (N_11199,N_10648,N_10858);
nand U11200 (N_11200,N_10443,N_10336);
xnor U11201 (N_11201,N_10281,N_10646);
nor U11202 (N_11202,N_10467,N_10747);
xnor U11203 (N_11203,N_10368,N_10512);
or U11204 (N_11204,N_10823,N_10792);
or U11205 (N_11205,N_10409,N_10550);
and U11206 (N_11206,N_10918,N_10510);
and U11207 (N_11207,N_10707,N_10035);
xnor U11208 (N_11208,N_10863,N_10192);
nor U11209 (N_11209,N_10686,N_10663);
nor U11210 (N_11210,N_10596,N_10556);
nor U11211 (N_11211,N_10338,N_10781);
and U11212 (N_11212,N_10825,N_10907);
xnor U11213 (N_11213,N_10151,N_10515);
nand U11214 (N_11214,N_10628,N_10101);
xor U11215 (N_11215,N_10078,N_10284);
nor U11216 (N_11216,N_10125,N_10308);
nor U11217 (N_11217,N_10121,N_10195);
nor U11218 (N_11218,N_10276,N_10103);
xnor U11219 (N_11219,N_10442,N_10459);
and U11220 (N_11220,N_10694,N_10108);
nor U11221 (N_11221,N_10302,N_10593);
or U11222 (N_11222,N_10569,N_10489);
nor U11223 (N_11223,N_10059,N_10022);
nand U11224 (N_11224,N_10640,N_10718);
and U11225 (N_11225,N_10376,N_10193);
or U11226 (N_11226,N_10219,N_10780);
nand U11227 (N_11227,N_10072,N_10421);
and U11228 (N_11228,N_10605,N_10307);
xor U11229 (N_11229,N_10360,N_10837);
and U11230 (N_11230,N_10571,N_10375);
xnor U11231 (N_11231,N_10198,N_10477);
nand U11232 (N_11232,N_10226,N_10900);
and U11233 (N_11233,N_10461,N_10961);
or U11234 (N_11234,N_10821,N_10597);
nor U11235 (N_11235,N_10586,N_10451);
nand U11236 (N_11236,N_10060,N_10642);
nand U11237 (N_11237,N_10229,N_10840);
and U11238 (N_11238,N_10043,N_10116);
nand U11239 (N_11239,N_10764,N_10687);
nand U11240 (N_11240,N_10793,N_10342);
xor U11241 (N_11241,N_10418,N_10834);
nand U11242 (N_11242,N_10006,N_10203);
and U11243 (N_11243,N_10874,N_10234);
and U11244 (N_11244,N_10692,N_10925);
xnor U11245 (N_11245,N_10798,N_10471);
and U11246 (N_11246,N_10816,N_10483);
or U11247 (N_11247,N_10851,N_10979);
and U11248 (N_11248,N_10494,N_10502);
nor U11249 (N_11249,N_10743,N_10880);
or U11250 (N_11250,N_10003,N_10244);
and U11251 (N_11251,N_10800,N_10185);
or U11252 (N_11252,N_10052,N_10853);
or U11253 (N_11253,N_10160,N_10482);
nand U11254 (N_11254,N_10393,N_10152);
nand U11255 (N_11255,N_10678,N_10742);
or U11256 (N_11256,N_10473,N_10806);
nor U11257 (N_11257,N_10609,N_10835);
nand U11258 (N_11258,N_10697,N_10963);
and U11259 (N_11259,N_10826,N_10300);
and U11260 (N_11260,N_10676,N_10020);
xor U11261 (N_11261,N_10319,N_10349);
nand U11262 (N_11262,N_10084,N_10932);
nor U11263 (N_11263,N_10905,N_10625);
or U11264 (N_11264,N_10218,N_10433);
xor U11265 (N_11265,N_10063,N_10268);
nor U11266 (N_11266,N_10911,N_10449);
xnor U11267 (N_11267,N_10122,N_10753);
or U11268 (N_11268,N_10754,N_10057);
and U11269 (N_11269,N_10758,N_10497);
or U11270 (N_11270,N_10945,N_10363);
xnor U11271 (N_11271,N_10161,N_10298);
xor U11272 (N_11272,N_10828,N_10601);
xor U11273 (N_11273,N_10873,N_10143);
nand U11274 (N_11274,N_10468,N_10132);
nand U11275 (N_11275,N_10259,N_10027);
and U11276 (N_11276,N_10243,N_10012);
xor U11277 (N_11277,N_10061,N_10413);
nor U11278 (N_11278,N_10183,N_10726);
nand U11279 (N_11279,N_10991,N_10484);
nor U11280 (N_11280,N_10087,N_10267);
xor U11281 (N_11281,N_10924,N_10952);
nor U11282 (N_11282,N_10566,N_10956);
xnor U11283 (N_11283,N_10083,N_10634);
and U11284 (N_11284,N_10715,N_10779);
nand U11285 (N_11285,N_10948,N_10139);
xor U11286 (N_11286,N_10135,N_10369);
and U11287 (N_11287,N_10479,N_10931);
and U11288 (N_11288,N_10446,N_10492);
nand U11289 (N_11289,N_10644,N_10844);
xnor U11290 (N_11290,N_10862,N_10316);
xnor U11291 (N_11291,N_10891,N_10942);
or U11292 (N_11292,N_10740,N_10665);
nor U11293 (N_11293,N_10872,N_10886);
or U11294 (N_11294,N_10506,N_10503);
or U11295 (N_11295,N_10385,N_10581);
and U11296 (N_11296,N_10699,N_10811);
xor U11297 (N_11297,N_10128,N_10355);
and U11298 (N_11298,N_10677,N_10303);
nor U11299 (N_11299,N_10209,N_10801);
nand U11300 (N_11300,N_10364,N_10768);
nor U11301 (N_11301,N_10731,N_10551);
xnor U11302 (N_11302,N_10833,N_10272);
or U11303 (N_11303,N_10180,N_10968);
and U11304 (N_11304,N_10888,N_10016);
and U11305 (N_11305,N_10055,N_10670);
nor U11306 (N_11306,N_10993,N_10211);
or U11307 (N_11307,N_10062,N_10926);
or U11308 (N_11308,N_10587,N_10046);
and U11309 (N_11309,N_10786,N_10102);
nand U11310 (N_11310,N_10410,N_10366);
nand U11311 (N_11311,N_10645,N_10123);
or U11312 (N_11312,N_10536,N_10313);
nand U11313 (N_11313,N_10445,N_10702);
xor U11314 (N_11314,N_10110,N_10708);
or U11315 (N_11315,N_10178,N_10214);
nor U11316 (N_11316,N_10902,N_10041);
or U11317 (N_11317,N_10654,N_10868);
nor U11318 (N_11318,N_10913,N_10094);
nor U11319 (N_11319,N_10564,N_10588);
xnor U11320 (N_11320,N_10416,N_10002);
xnor U11321 (N_11321,N_10824,N_10478);
nor U11322 (N_11322,N_10474,N_10199);
nand U11323 (N_11323,N_10401,N_10751);
nand U11324 (N_11324,N_10287,N_10684);
nor U11325 (N_11325,N_10832,N_10129);
or U11326 (N_11326,N_10802,N_10589);
and U11327 (N_11327,N_10671,N_10191);
nor U11328 (N_11328,N_10875,N_10735);
nor U11329 (N_11329,N_10408,N_10950);
nor U11330 (N_11330,N_10958,N_10894);
or U11331 (N_11331,N_10790,N_10960);
nand U11332 (N_11332,N_10075,N_10522);
xor U11333 (N_11333,N_10514,N_10335);
xnor U11334 (N_11334,N_10124,N_10955);
nand U11335 (N_11335,N_10939,N_10999);
nor U11336 (N_11336,N_10463,N_10476);
nor U11337 (N_11337,N_10120,N_10187);
or U11338 (N_11338,N_10235,N_10881);
xnor U11339 (N_11339,N_10391,N_10629);
xor U11340 (N_11340,N_10843,N_10420);
and U11341 (N_11341,N_10086,N_10912);
nor U11342 (N_11342,N_10761,N_10280);
and U11343 (N_11343,N_10666,N_10795);
and U11344 (N_11344,N_10412,N_10384);
nand U11345 (N_11345,N_10164,N_10077);
nor U11346 (N_11346,N_10493,N_10674);
nor U11347 (N_11347,N_10182,N_10021);
or U11348 (N_11348,N_10184,N_10711);
and U11349 (N_11349,N_10720,N_10532);
nor U11350 (N_11350,N_10389,N_10282);
xnor U11351 (N_11351,N_10005,N_10724);
nor U11352 (N_11352,N_10168,N_10205);
nor U11353 (N_11353,N_10200,N_10777);
nand U11354 (N_11354,N_10098,N_10396);
nand U11355 (N_11355,N_10570,N_10631);
xnor U11356 (N_11356,N_10849,N_10701);
and U11357 (N_11357,N_10230,N_10240);
nor U11358 (N_11358,N_10019,N_10269);
or U11359 (N_11359,N_10312,N_10542);
nor U11360 (N_11360,N_10543,N_10067);
or U11361 (N_11361,N_10225,N_10206);
or U11362 (N_11362,N_10855,N_10018);
xnor U11363 (N_11363,N_10752,N_10673);
nand U11364 (N_11364,N_10306,N_10305);
and U11365 (N_11365,N_10374,N_10047);
and U11366 (N_11366,N_10535,N_10074);
and U11367 (N_11367,N_10283,N_10553);
xor U11368 (N_11368,N_10544,N_10641);
and U11369 (N_11369,N_10706,N_10362);
nor U11370 (N_11370,N_10526,N_10383);
and U11371 (N_11371,N_10774,N_10620);
or U11372 (N_11372,N_10429,N_10334);
nand U11373 (N_11373,N_10527,N_10089);
xnor U11374 (N_11374,N_10846,N_10105);
nor U11375 (N_11375,N_10594,N_10256);
xor U11376 (N_11376,N_10223,N_10310);
and U11377 (N_11377,N_10361,N_10026);
nor U11378 (N_11378,N_10870,N_10685);
nand U11379 (N_11379,N_10327,N_10261);
or U11380 (N_11380,N_10422,N_10732);
nor U11381 (N_11381,N_10044,N_10118);
or U11382 (N_11382,N_10943,N_10787);
nor U11383 (N_11383,N_10679,N_10270);
and U11384 (N_11384,N_10983,N_10916);
and U11385 (N_11385,N_10010,N_10394);
and U11386 (N_11386,N_10727,N_10224);
xnor U11387 (N_11387,N_10250,N_10716);
and U11388 (N_11388,N_10464,N_10519);
and U11389 (N_11389,N_10545,N_10696);
nor U11390 (N_11390,N_10595,N_10733);
or U11391 (N_11391,N_10721,N_10607);
and U11392 (N_11392,N_10922,N_10343);
nand U11393 (N_11393,N_10734,N_10462);
or U11394 (N_11394,N_10359,N_10079);
or U11395 (N_11395,N_10174,N_10622);
xnor U11396 (N_11396,N_10969,N_10050);
nand U11397 (N_11397,N_10430,N_10590);
or U11398 (N_11398,N_10637,N_10040);
or U11399 (N_11399,N_10627,N_10015);
nand U11400 (N_11400,N_10301,N_10114);
nand U11401 (N_11401,N_10808,N_10507);
xnor U11402 (N_11402,N_10248,N_10884);
and U11403 (N_11403,N_10658,N_10137);
xnor U11404 (N_11404,N_10082,N_10929);
xor U11405 (N_11405,N_10563,N_10661);
or U11406 (N_11406,N_10011,N_10517);
and U11407 (N_11407,N_10710,N_10814);
nor U11408 (N_11408,N_10930,N_10415);
nand U11409 (N_11409,N_10583,N_10140);
nor U11410 (N_11410,N_10951,N_10533);
xnor U11411 (N_11411,N_10980,N_10744);
xnor U11412 (N_11412,N_10513,N_10453);
xnor U11413 (N_11413,N_10107,N_10142);
xnor U11414 (N_11414,N_10228,N_10688);
or U11415 (N_11415,N_10632,N_10304);
nand U11416 (N_11416,N_10480,N_10397);
xnor U11417 (N_11417,N_10216,N_10149);
nor U11418 (N_11418,N_10166,N_10647);
nor U11419 (N_11419,N_10071,N_10920);
or U11420 (N_11420,N_10215,N_10501);
and U11421 (N_11421,N_10659,N_10822);
nor U11422 (N_11422,N_10347,N_10511);
xnor U11423 (N_11423,N_10838,N_10444);
xnor U11424 (N_11424,N_10399,N_10938);
nand U11425 (N_11425,N_10096,N_10469);
nand U11426 (N_11426,N_10403,N_10602);
and U11427 (N_11427,N_10233,N_10576);
or U11428 (N_11428,N_10509,N_10320);
and U11429 (N_11429,N_10392,N_10982);
nor U11430 (N_11430,N_10869,N_10237);
and U11431 (N_11431,N_10528,N_10440);
nand U11432 (N_11432,N_10073,N_10804);
and U11433 (N_11433,N_10657,N_10953);
nor U11434 (N_11434,N_10279,N_10251);
xor U11435 (N_11435,N_10247,N_10763);
xnor U11436 (N_11436,N_10577,N_10598);
nand U11437 (N_11437,N_10207,N_10093);
or U11438 (N_11438,N_10772,N_10820);
or U11439 (N_11439,N_10575,N_10438);
or U11440 (N_11440,N_10332,N_10633);
and U11441 (N_11441,N_10766,N_10604);
nor U11442 (N_11442,N_10741,N_10799);
xnor U11443 (N_11443,N_10693,N_10704);
xor U11444 (N_11444,N_10111,N_10848);
and U11445 (N_11445,N_10624,N_10008);
nor U11446 (N_11446,N_10460,N_10398);
xor U11447 (N_11447,N_10500,N_10351);
or U11448 (N_11448,N_10381,N_10490);
and U11449 (N_11449,N_10965,N_10435);
nor U11450 (N_11450,N_10904,N_10580);
or U11451 (N_11451,N_10841,N_10530);
nor U11452 (N_11452,N_10163,N_10748);
and U11453 (N_11453,N_10271,N_10190);
and U11454 (N_11454,N_10817,N_10552);
nand U11455 (N_11455,N_10417,N_10815);
xnor U11456 (N_11456,N_10630,N_10585);
or U11457 (N_11457,N_10042,N_10292);
nand U11458 (N_11458,N_10344,N_10337);
nor U11459 (N_11459,N_10395,N_10672);
or U11460 (N_11460,N_10104,N_10650);
xnor U11461 (N_11461,N_10614,N_10295);
and U11462 (N_11462,N_10232,N_10265);
nand U11463 (N_11463,N_10339,N_10599);
or U11464 (N_11464,N_10365,N_10274);
or U11465 (N_11465,N_10202,N_10767);
nand U11466 (N_11466,N_10099,N_10058);
nor U11467 (N_11467,N_10898,N_10419);
or U11468 (N_11468,N_10988,N_10879);
nand U11469 (N_11469,N_10529,N_10288);
or U11470 (N_11470,N_10286,N_10297);
or U11471 (N_11471,N_10097,N_10179);
and U11472 (N_11472,N_10414,N_10450);
nand U11473 (N_11473,N_10909,N_10387);
nor U11474 (N_11474,N_10867,N_10358);
nand U11475 (N_11475,N_10928,N_10186);
nor U11476 (N_11476,N_10263,N_10208);
nor U11477 (N_11477,N_10194,N_10400);
xor U11478 (N_11478,N_10009,N_10475);
and U11479 (N_11479,N_10145,N_10662);
xor U11480 (N_11480,N_10975,N_10285);
nor U11481 (N_11481,N_10829,N_10883);
or U11482 (N_11482,N_10239,N_10045);
nand U11483 (N_11483,N_10903,N_10746);
xor U11484 (N_11484,N_10959,N_10555);
or U11485 (N_11485,N_10769,N_10842);
or U11486 (N_11486,N_10865,N_10066);
nor U11487 (N_11487,N_10034,N_10992);
xnor U11488 (N_11488,N_10750,N_10691);
xnor U11489 (N_11489,N_10971,N_10212);
nand U11490 (N_11490,N_10154,N_10328);
and U11491 (N_11491,N_10749,N_10729);
xnor U11492 (N_11492,N_10081,N_10541);
xor U11493 (N_11493,N_10348,N_10379);
and U11494 (N_11494,N_10117,N_10972);
or U11495 (N_11495,N_10717,N_10367);
nor U11496 (N_11496,N_10262,N_10257);
xnor U11497 (N_11497,N_10131,N_10669);
and U11498 (N_11498,N_10439,N_10736);
nand U11499 (N_11499,N_10324,N_10340);
xnor U11500 (N_11500,N_10539,N_10803);
nand U11501 (N_11501,N_10951,N_10936);
nand U11502 (N_11502,N_10210,N_10228);
or U11503 (N_11503,N_10801,N_10905);
or U11504 (N_11504,N_10494,N_10830);
nor U11505 (N_11505,N_10466,N_10365);
nand U11506 (N_11506,N_10968,N_10125);
nand U11507 (N_11507,N_10679,N_10906);
or U11508 (N_11508,N_10761,N_10977);
nand U11509 (N_11509,N_10795,N_10764);
nor U11510 (N_11510,N_10156,N_10851);
nand U11511 (N_11511,N_10338,N_10494);
nor U11512 (N_11512,N_10908,N_10947);
nor U11513 (N_11513,N_10862,N_10199);
nand U11514 (N_11514,N_10915,N_10609);
and U11515 (N_11515,N_10687,N_10386);
nor U11516 (N_11516,N_10878,N_10865);
and U11517 (N_11517,N_10671,N_10064);
and U11518 (N_11518,N_10239,N_10907);
xnor U11519 (N_11519,N_10690,N_10617);
or U11520 (N_11520,N_10344,N_10735);
nor U11521 (N_11521,N_10450,N_10400);
and U11522 (N_11522,N_10349,N_10882);
nor U11523 (N_11523,N_10356,N_10033);
or U11524 (N_11524,N_10804,N_10839);
or U11525 (N_11525,N_10787,N_10984);
nand U11526 (N_11526,N_10538,N_10646);
nand U11527 (N_11527,N_10574,N_10042);
nand U11528 (N_11528,N_10126,N_10243);
and U11529 (N_11529,N_10046,N_10803);
xnor U11530 (N_11530,N_10544,N_10409);
or U11531 (N_11531,N_10416,N_10218);
nor U11532 (N_11532,N_10896,N_10275);
nand U11533 (N_11533,N_10716,N_10436);
nor U11534 (N_11534,N_10847,N_10625);
and U11535 (N_11535,N_10892,N_10937);
nor U11536 (N_11536,N_10661,N_10560);
nand U11537 (N_11537,N_10127,N_10377);
and U11538 (N_11538,N_10095,N_10008);
nor U11539 (N_11539,N_10990,N_10942);
xnor U11540 (N_11540,N_10908,N_10724);
xor U11541 (N_11541,N_10975,N_10503);
and U11542 (N_11542,N_10296,N_10740);
or U11543 (N_11543,N_10848,N_10059);
nand U11544 (N_11544,N_10539,N_10241);
nand U11545 (N_11545,N_10359,N_10712);
nand U11546 (N_11546,N_10125,N_10318);
and U11547 (N_11547,N_10055,N_10535);
or U11548 (N_11548,N_10767,N_10581);
nor U11549 (N_11549,N_10699,N_10646);
nor U11550 (N_11550,N_10692,N_10603);
xnor U11551 (N_11551,N_10013,N_10822);
and U11552 (N_11552,N_10732,N_10117);
nor U11553 (N_11553,N_10688,N_10728);
and U11554 (N_11554,N_10261,N_10064);
xnor U11555 (N_11555,N_10817,N_10942);
or U11556 (N_11556,N_10667,N_10724);
nand U11557 (N_11557,N_10233,N_10789);
and U11558 (N_11558,N_10263,N_10384);
nor U11559 (N_11559,N_10610,N_10727);
nor U11560 (N_11560,N_10508,N_10514);
or U11561 (N_11561,N_10036,N_10323);
xor U11562 (N_11562,N_10557,N_10255);
nor U11563 (N_11563,N_10171,N_10794);
nand U11564 (N_11564,N_10597,N_10164);
nand U11565 (N_11565,N_10748,N_10253);
and U11566 (N_11566,N_10741,N_10549);
nand U11567 (N_11567,N_10463,N_10028);
xor U11568 (N_11568,N_10302,N_10285);
nand U11569 (N_11569,N_10359,N_10450);
xor U11570 (N_11570,N_10686,N_10721);
nor U11571 (N_11571,N_10931,N_10808);
nand U11572 (N_11572,N_10675,N_10646);
and U11573 (N_11573,N_10126,N_10739);
nand U11574 (N_11574,N_10021,N_10924);
nor U11575 (N_11575,N_10322,N_10029);
nor U11576 (N_11576,N_10664,N_10780);
and U11577 (N_11577,N_10113,N_10166);
nor U11578 (N_11578,N_10501,N_10016);
nor U11579 (N_11579,N_10161,N_10952);
or U11580 (N_11580,N_10407,N_10446);
and U11581 (N_11581,N_10797,N_10070);
and U11582 (N_11582,N_10774,N_10017);
xor U11583 (N_11583,N_10480,N_10728);
nor U11584 (N_11584,N_10903,N_10428);
nand U11585 (N_11585,N_10776,N_10544);
nand U11586 (N_11586,N_10441,N_10770);
and U11587 (N_11587,N_10862,N_10847);
nor U11588 (N_11588,N_10212,N_10568);
nor U11589 (N_11589,N_10148,N_10285);
and U11590 (N_11590,N_10613,N_10431);
and U11591 (N_11591,N_10112,N_10296);
nand U11592 (N_11592,N_10266,N_10044);
and U11593 (N_11593,N_10163,N_10671);
nand U11594 (N_11594,N_10905,N_10274);
and U11595 (N_11595,N_10655,N_10839);
xor U11596 (N_11596,N_10189,N_10365);
xor U11597 (N_11597,N_10628,N_10313);
xnor U11598 (N_11598,N_10913,N_10484);
and U11599 (N_11599,N_10397,N_10796);
or U11600 (N_11600,N_10203,N_10642);
nand U11601 (N_11601,N_10890,N_10916);
nor U11602 (N_11602,N_10018,N_10886);
nor U11603 (N_11603,N_10170,N_10954);
xor U11604 (N_11604,N_10721,N_10968);
nand U11605 (N_11605,N_10096,N_10163);
nor U11606 (N_11606,N_10729,N_10325);
and U11607 (N_11607,N_10488,N_10141);
or U11608 (N_11608,N_10324,N_10890);
or U11609 (N_11609,N_10744,N_10145);
xnor U11610 (N_11610,N_10843,N_10102);
or U11611 (N_11611,N_10347,N_10604);
nor U11612 (N_11612,N_10474,N_10947);
xnor U11613 (N_11613,N_10771,N_10640);
xor U11614 (N_11614,N_10550,N_10284);
nand U11615 (N_11615,N_10165,N_10875);
xor U11616 (N_11616,N_10068,N_10080);
nor U11617 (N_11617,N_10723,N_10466);
and U11618 (N_11618,N_10004,N_10783);
xor U11619 (N_11619,N_10936,N_10855);
and U11620 (N_11620,N_10278,N_10802);
nand U11621 (N_11621,N_10630,N_10918);
xor U11622 (N_11622,N_10721,N_10590);
and U11623 (N_11623,N_10758,N_10442);
nor U11624 (N_11624,N_10763,N_10405);
nor U11625 (N_11625,N_10780,N_10915);
xnor U11626 (N_11626,N_10524,N_10622);
or U11627 (N_11627,N_10012,N_10712);
nand U11628 (N_11628,N_10810,N_10287);
nand U11629 (N_11629,N_10010,N_10866);
and U11630 (N_11630,N_10646,N_10702);
nor U11631 (N_11631,N_10567,N_10073);
or U11632 (N_11632,N_10350,N_10272);
xor U11633 (N_11633,N_10069,N_10094);
nor U11634 (N_11634,N_10326,N_10063);
xor U11635 (N_11635,N_10135,N_10317);
xnor U11636 (N_11636,N_10795,N_10441);
nor U11637 (N_11637,N_10709,N_10693);
nand U11638 (N_11638,N_10292,N_10413);
or U11639 (N_11639,N_10710,N_10494);
nand U11640 (N_11640,N_10484,N_10007);
nor U11641 (N_11641,N_10578,N_10632);
nor U11642 (N_11642,N_10625,N_10590);
nor U11643 (N_11643,N_10028,N_10063);
nand U11644 (N_11644,N_10374,N_10053);
nand U11645 (N_11645,N_10561,N_10044);
or U11646 (N_11646,N_10610,N_10124);
or U11647 (N_11647,N_10788,N_10217);
nand U11648 (N_11648,N_10432,N_10158);
xor U11649 (N_11649,N_10408,N_10933);
and U11650 (N_11650,N_10493,N_10333);
and U11651 (N_11651,N_10945,N_10850);
and U11652 (N_11652,N_10044,N_10825);
xor U11653 (N_11653,N_10354,N_10928);
and U11654 (N_11654,N_10990,N_10220);
nor U11655 (N_11655,N_10916,N_10713);
nor U11656 (N_11656,N_10438,N_10357);
or U11657 (N_11657,N_10448,N_10334);
and U11658 (N_11658,N_10092,N_10602);
nand U11659 (N_11659,N_10363,N_10575);
or U11660 (N_11660,N_10200,N_10031);
or U11661 (N_11661,N_10428,N_10976);
and U11662 (N_11662,N_10570,N_10182);
nor U11663 (N_11663,N_10396,N_10807);
nor U11664 (N_11664,N_10700,N_10708);
nand U11665 (N_11665,N_10402,N_10729);
nand U11666 (N_11666,N_10187,N_10900);
or U11667 (N_11667,N_10149,N_10491);
and U11668 (N_11668,N_10054,N_10219);
nand U11669 (N_11669,N_10064,N_10339);
nor U11670 (N_11670,N_10436,N_10395);
xor U11671 (N_11671,N_10155,N_10186);
nand U11672 (N_11672,N_10433,N_10309);
nand U11673 (N_11673,N_10733,N_10762);
nand U11674 (N_11674,N_10854,N_10592);
nand U11675 (N_11675,N_10680,N_10711);
and U11676 (N_11676,N_10452,N_10356);
xor U11677 (N_11677,N_10034,N_10394);
nor U11678 (N_11678,N_10167,N_10909);
xor U11679 (N_11679,N_10995,N_10431);
nand U11680 (N_11680,N_10422,N_10724);
and U11681 (N_11681,N_10235,N_10453);
or U11682 (N_11682,N_10468,N_10614);
nand U11683 (N_11683,N_10561,N_10967);
and U11684 (N_11684,N_10365,N_10664);
nand U11685 (N_11685,N_10694,N_10912);
xor U11686 (N_11686,N_10838,N_10016);
or U11687 (N_11687,N_10014,N_10730);
nand U11688 (N_11688,N_10590,N_10059);
and U11689 (N_11689,N_10662,N_10350);
nor U11690 (N_11690,N_10818,N_10088);
nor U11691 (N_11691,N_10058,N_10221);
nand U11692 (N_11692,N_10866,N_10134);
nor U11693 (N_11693,N_10408,N_10439);
and U11694 (N_11694,N_10298,N_10750);
nor U11695 (N_11695,N_10200,N_10998);
nor U11696 (N_11696,N_10303,N_10118);
or U11697 (N_11697,N_10896,N_10826);
or U11698 (N_11698,N_10666,N_10392);
nor U11699 (N_11699,N_10160,N_10772);
nor U11700 (N_11700,N_10654,N_10276);
or U11701 (N_11701,N_10200,N_10195);
nand U11702 (N_11702,N_10787,N_10853);
nand U11703 (N_11703,N_10729,N_10101);
and U11704 (N_11704,N_10039,N_10312);
xnor U11705 (N_11705,N_10614,N_10826);
nor U11706 (N_11706,N_10548,N_10757);
or U11707 (N_11707,N_10399,N_10957);
or U11708 (N_11708,N_10561,N_10484);
and U11709 (N_11709,N_10102,N_10467);
nand U11710 (N_11710,N_10549,N_10438);
nor U11711 (N_11711,N_10910,N_10865);
and U11712 (N_11712,N_10551,N_10271);
nand U11713 (N_11713,N_10883,N_10332);
or U11714 (N_11714,N_10908,N_10467);
or U11715 (N_11715,N_10222,N_10791);
or U11716 (N_11716,N_10926,N_10791);
and U11717 (N_11717,N_10078,N_10297);
nor U11718 (N_11718,N_10385,N_10127);
or U11719 (N_11719,N_10211,N_10908);
or U11720 (N_11720,N_10226,N_10494);
xor U11721 (N_11721,N_10836,N_10312);
xor U11722 (N_11722,N_10219,N_10314);
xnor U11723 (N_11723,N_10176,N_10488);
nand U11724 (N_11724,N_10542,N_10385);
xor U11725 (N_11725,N_10135,N_10462);
nor U11726 (N_11726,N_10859,N_10383);
and U11727 (N_11727,N_10481,N_10078);
and U11728 (N_11728,N_10165,N_10150);
or U11729 (N_11729,N_10401,N_10105);
and U11730 (N_11730,N_10118,N_10096);
and U11731 (N_11731,N_10715,N_10393);
nor U11732 (N_11732,N_10183,N_10869);
xor U11733 (N_11733,N_10219,N_10809);
xnor U11734 (N_11734,N_10311,N_10604);
or U11735 (N_11735,N_10751,N_10022);
or U11736 (N_11736,N_10914,N_10081);
nor U11737 (N_11737,N_10479,N_10675);
xnor U11738 (N_11738,N_10613,N_10155);
nand U11739 (N_11739,N_10570,N_10914);
or U11740 (N_11740,N_10881,N_10403);
or U11741 (N_11741,N_10905,N_10755);
and U11742 (N_11742,N_10554,N_10618);
xnor U11743 (N_11743,N_10794,N_10644);
xor U11744 (N_11744,N_10084,N_10343);
nand U11745 (N_11745,N_10384,N_10699);
nand U11746 (N_11746,N_10478,N_10400);
or U11747 (N_11747,N_10110,N_10325);
xnor U11748 (N_11748,N_10238,N_10279);
xor U11749 (N_11749,N_10822,N_10012);
xnor U11750 (N_11750,N_10682,N_10242);
or U11751 (N_11751,N_10869,N_10969);
nand U11752 (N_11752,N_10192,N_10392);
and U11753 (N_11753,N_10628,N_10753);
and U11754 (N_11754,N_10367,N_10410);
nor U11755 (N_11755,N_10299,N_10885);
xor U11756 (N_11756,N_10142,N_10238);
and U11757 (N_11757,N_10966,N_10383);
xnor U11758 (N_11758,N_10548,N_10657);
xnor U11759 (N_11759,N_10356,N_10545);
or U11760 (N_11760,N_10074,N_10212);
or U11761 (N_11761,N_10085,N_10965);
nand U11762 (N_11762,N_10495,N_10746);
or U11763 (N_11763,N_10473,N_10618);
or U11764 (N_11764,N_10339,N_10785);
or U11765 (N_11765,N_10657,N_10649);
or U11766 (N_11766,N_10432,N_10289);
nor U11767 (N_11767,N_10476,N_10444);
nor U11768 (N_11768,N_10003,N_10007);
and U11769 (N_11769,N_10056,N_10799);
or U11770 (N_11770,N_10112,N_10704);
nand U11771 (N_11771,N_10069,N_10836);
xor U11772 (N_11772,N_10768,N_10130);
and U11773 (N_11773,N_10137,N_10882);
nand U11774 (N_11774,N_10777,N_10202);
and U11775 (N_11775,N_10167,N_10495);
xnor U11776 (N_11776,N_10076,N_10293);
xor U11777 (N_11777,N_10988,N_10566);
or U11778 (N_11778,N_10891,N_10022);
nor U11779 (N_11779,N_10567,N_10913);
xnor U11780 (N_11780,N_10666,N_10309);
and U11781 (N_11781,N_10796,N_10528);
or U11782 (N_11782,N_10719,N_10135);
or U11783 (N_11783,N_10347,N_10541);
xnor U11784 (N_11784,N_10043,N_10744);
or U11785 (N_11785,N_10859,N_10963);
or U11786 (N_11786,N_10493,N_10944);
and U11787 (N_11787,N_10799,N_10135);
xor U11788 (N_11788,N_10912,N_10227);
and U11789 (N_11789,N_10190,N_10639);
and U11790 (N_11790,N_10253,N_10980);
nand U11791 (N_11791,N_10383,N_10331);
nand U11792 (N_11792,N_10323,N_10387);
xnor U11793 (N_11793,N_10155,N_10261);
nor U11794 (N_11794,N_10842,N_10422);
nor U11795 (N_11795,N_10700,N_10938);
or U11796 (N_11796,N_10452,N_10867);
xnor U11797 (N_11797,N_10277,N_10863);
xnor U11798 (N_11798,N_10989,N_10142);
and U11799 (N_11799,N_10058,N_10077);
nand U11800 (N_11800,N_10497,N_10218);
or U11801 (N_11801,N_10489,N_10546);
nor U11802 (N_11802,N_10610,N_10207);
or U11803 (N_11803,N_10873,N_10920);
xnor U11804 (N_11804,N_10259,N_10192);
or U11805 (N_11805,N_10508,N_10703);
and U11806 (N_11806,N_10141,N_10109);
and U11807 (N_11807,N_10257,N_10394);
xor U11808 (N_11808,N_10461,N_10238);
nand U11809 (N_11809,N_10542,N_10181);
nand U11810 (N_11810,N_10672,N_10283);
and U11811 (N_11811,N_10397,N_10410);
xor U11812 (N_11812,N_10304,N_10546);
or U11813 (N_11813,N_10446,N_10412);
nand U11814 (N_11814,N_10443,N_10681);
or U11815 (N_11815,N_10598,N_10099);
nand U11816 (N_11816,N_10713,N_10931);
nor U11817 (N_11817,N_10922,N_10618);
nor U11818 (N_11818,N_10183,N_10458);
nor U11819 (N_11819,N_10244,N_10635);
nor U11820 (N_11820,N_10060,N_10286);
and U11821 (N_11821,N_10898,N_10075);
nand U11822 (N_11822,N_10509,N_10954);
xor U11823 (N_11823,N_10246,N_10935);
nand U11824 (N_11824,N_10666,N_10011);
xor U11825 (N_11825,N_10632,N_10356);
nor U11826 (N_11826,N_10158,N_10248);
nand U11827 (N_11827,N_10853,N_10847);
or U11828 (N_11828,N_10666,N_10355);
nor U11829 (N_11829,N_10991,N_10135);
or U11830 (N_11830,N_10002,N_10911);
nor U11831 (N_11831,N_10260,N_10647);
and U11832 (N_11832,N_10036,N_10002);
and U11833 (N_11833,N_10210,N_10916);
or U11834 (N_11834,N_10751,N_10635);
nor U11835 (N_11835,N_10505,N_10764);
and U11836 (N_11836,N_10056,N_10261);
nor U11837 (N_11837,N_10819,N_10512);
and U11838 (N_11838,N_10918,N_10967);
and U11839 (N_11839,N_10424,N_10799);
or U11840 (N_11840,N_10112,N_10643);
and U11841 (N_11841,N_10483,N_10595);
nor U11842 (N_11842,N_10830,N_10739);
nand U11843 (N_11843,N_10644,N_10040);
and U11844 (N_11844,N_10033,N_10514);
and U11845 (N_11845,N_10583,N_10354);
nor U11846 (N_11846,N_10207,N_10452);
and U11847 (N_11847,N_10116,N_10010);
nor U11848 (N_11848,N_10034,N_10930);
or U11849 (N_11849,N_10876,N_10651);
nand U11850 (N_11850,N_10014,N_10316);
nand U11851 (N_11851,N_10825,N_10045);
xor U11852 (N_11852,N_10990,N_10567);
xnor U11853 (N_11853,N_10996,N_10397);
or U11854 (N_11854,N_10120,N_10222);
nand U11855 (N_11855,N_10733,N_10428);
xnor U11856 (N_11856,N_10929,N_10984);
or U11857 (N_11857,N_10643,N_10135);
nor U11858 (N_11858,N_10420,N_10269);
nand U11859 (N_11859,N_10684,N_10280);
nand U11860 (N_11860,N_10283,N_10180);
nor U11861 (N_11861,N_10270,N_10500);
or U11862 (N_11862,N_10758,N_10674);
and U11863 (N_11863,N_10066,N_10456);
and U11864 (N_11864,N_10118,N_10789);
or U11865 (N_11865,N_10940,N_10437);
and U11866 (N_11866,N_10626,N_10771);
nand U11867 (N_11867,N_10993,N_10736);
nor U11868 (N_11868,N_10001,N_10266);
nand U11869 (N_11869,N_10717,N_10948);
nand U11870 (N_11870,N_10422,N_10061);
xnor U11871 (N_11871,N_10433,N_10325);
nor U11872 (N_11872,N_10331,N_10967);
or U11873 (N_11873,N_10386,N_10345);
and U11874 (N_11874,N_10663,N_10655);
nand U11875 (N_11875,N_10073,N_10580);
xnor U11876 (N_11876,N_10216,N_10837);
xnor U11877 (N_11877,N_10923,N_10215);
or U11878 (N_11878,N_10498,N_10179);
nor U11879 (N_11879,N_10036,N_10441);
or U11880 (N_11880,N_10530,N_10770);
xor U11881 (N_11881,N_10826,N_10879);
nand U11882 (N_11882,N_10810,N_10065);
xor U11883 (N_11883,N_10291,N_10179);
or U11884 (N_11884,N_10559,N_10980);
or U11885 (N_11885,N_10512,N_10580);
xor U11886 (N_11886,N_10404,N_10632);
nor U11887 (N_11887,N_10748,N_10421);
xor U11888 (N_11888,N_10050,N_10136);
nor U11889 (N_11889,N_10619,N_10208);
xor U11890 (N_11890,N_10471,N_10397);
and U11891 (N_11891,N_10818,N_10163);
and U11892 (N_11892,N_10152,N_10602);
xnor U11893 (N_11893,N_10694,N_10909);
and U11894 (N_11894,N_10990,N_10552);
nor U11895 (N_11895,N_10264,N_10382);
and U11896 (N_11896,N_10826,N_10392);
nand U11897 (N_11897,N_10756,N_10403);
nor U11898 (N_11898,N_10789,N_10762);
and U11899 (N_11899,N_10168,N_10377);
nor U11900 (N_11900,N_10299,N_10241);
xor U11901 (N_11901,N_10542,N_10111);
xor U11902 (N_11902,N_10606,N_10443);
nand U11903 (N_11903,N_10956,N_10173);
nand U11904 (N_11904,N_10945,N_10091);
or U11905 (N_11905,N_10468,N_10693);
nor U11906 (N_11906,N_10783,N_10803);
nand U11907 (N_11907,N_10089,N_10224);
xor U11908 (N_11908,N_10769,N_10525);
nand U11909 (N_11909,N_10060,N_10331);
or U11910 (N_11910,N_10766,N_10351);
nand U11911 (N_11911,N_10179,N_10143);
xor U11912 (N_11912,N_10035,N_10795);
nor U11913 (N_11913,N_10958,N_10136);
nand U11914 (N_11914,N_10624,N_10666);
nor U11915 (N_11915,N_10420,N_10544);
nor U11916 (N_11916,N_10306,N_10874);
nor U11917 (N_11917,N_10619,N_10444);
xor U11918 (N_11918,N_10988,N_10583);
nor U11919 (N_11919,N_10435,N_10455);
xnor U11920 (N_11920,N_10762,N_10679);
nand U11921 (N_11921,N_10477,N_10519);
and U11922 (N_11922,N_10191,N_10271);
or U11923 (N_11923,N_10676,N_10076);
nor U11924 (N_11924,N_10204,N_10074);
nor U11925 (N_11925,N_10024,N_10584);
nand U11926 (N_11926,N_10918,N_10128);
and U11927 (N_11927,N_10163,N_10646);
and U11928 (N_11928,N_10866,N_10905);
nor U11929 (N_11929,N_10626,N_10778);
nand U11930 (N_11930,N_10883,N_10460);
xnor U11931 (N_11931,N_10631,N_10904);
nor U11932 (N_11932,N_10509,N_10435);
nor U11933 (N_11933,N_10589,N_10886);
or U11934 (N_11934,N_10196,N_10896);
or U11935 (N_11935,N_10516,N_10204);
and U11936 (N_11936,N_10880,N_10685);
nor U11937 (N_11937,N_10763,N_10919);
and U11938 (N_11938,N_10936,N_10175);
nand U11939 (N_11939,N_10144,N_10254);
nor U11940 (N_11940,N_10290,N_10585);
xnor U11941 (N_11941,N_10113,N_10469);
xnor U11942 (N_11942,N_10858,N_10239);
nand U11943 (N_11943,N_10287,N_10228);
nand U11944 (N_11944,N_10206,N_10873);
nand U11945 (N_11945,N_10667,N_10588);
or U11946 (N_11946,N_10834,N_10061);
xnor U11947 (N_11947,N_10951,N_10194);
or U11948 (N_11948,N_10560,N_10078);
and U11949 (N_11949,N_10330,N_10993);
nand U11950 (N_11950,N_10104,N_10570);
nor U11951 (N_11951,N_10736,N_10323);
and U11952 (N_11952,N_10521,N_10910);
or U11953 (N_11953,N_10360,N_10505);
nand U11954 (N_11954,N_10586,N_10589);
or U11955 (N_11955,N_10230,N_10079);
xor U11956 (N_11956,N_10790,N_10453);
nor U11957 (N_11957,N_10623,N_10596);
and U11958 (N_11958,N_10378,N_10866);
nor U11959 (N_11959,N_10677,N_10191);
or U11960 (N_11960,N_10826,N_10460);
xnor U11961 (N_11961,N_10954,N_10874);
nand U11962 (N_11962,N_10252,N_10312);
or U11963 (N_11963,N_10643,N_10806);
or U11964 (N_11964,N_10478,N_10903);
nand U11965 (N_11965,N_10225,N_10319);
nand U11966 (N_11966,N_10246,N_10287);
nor U11967 (N_11967,N_10260,N_10225);
or U11968 (N_11968,N_10645,N_10330);
or U11969 (N_11969,N_10529,N_10654);
nand U11970 (N_11970,N_10820,N_10423);
xor U11971 (N_11971,N_10929,N_10530);
nand U11972 (N_11972,N_10064,N_10969);
nor U11973 (N_11973,N_10302,N_10090);
nor U11974 (N_11974,N_10260,N_10556);
xnor U11975 (N_11975,N_10676,N_10673);
and U11976 (N_11976,N_10035,N_10622);
nand U11977 (N_11977,N_10027,N_10805);
nor U11978 (N_11978,N_10936,N_10114);
nand U11979 (N_11979,N_10828,N_10514);
and U11980 (N_11980,N_10905,N_10758);
nand U11981 (N_11981,N_10127,N_10926);
or U11982 (N_11982,N_10147,N_10393);
nand U11983 (N_11983,N_10276,N_10932);
and U11984 (N_11984,N_10809,N_10828);
or U11985 (N_11985,N_10038,N_10253);
and U11986 (N_11986,N_10723,N_10647);
nand U11987 (N_11987,N_10711,N_10329);
xor U11988 (N_11988,N_10893,N_10411);
xnor U11989 (N_11989,N_10032,N_10289);
and U11990 (N_11990,N_10462,N_10589);
and U11991 (N_11991,N_10626,N_10933);
or U11992 (N_11992,N_10188,N_10478);
and U11993 (N_11993,N_10214,N_10807);
and U11994 (N_11994,N_10050,N_10894);
nor U11995 (N_11995,N_10315,N_10827);
nand U11996 (N_11996,N_10652,N_10737);
and U11997 (N_11997,N_10319,N_10329);
nand U11998 (N_11998,N_10252,N_10065);
nor U11999 (N_11999,N_10350,N_10964);
or U12000 (N_12000,N_11629,N_11408);
nor U12001 (N_12001,N_11511,N_11569);
or U12002 (N_12002,N_11519,N_11219);
xnor U12003 (N_12003,N_11248,N_11421);
and U12004 (N_12004,N_11839,N_11991);
and U12005 (N_12005,N_11385,N_11636);
or U12006 (N_12006,N_11759,N_11512);
and U12007 (N_12007,N_11800,N_11309);
or U12008 (N_12008,N_11955,N_11576);
or U12009 (N_12009,N_11648,N_11657);
or U12010 (N_12010,N_11726,N_11483);
and U12011 (N_12011,N_11567,N_11665);
nor U12012 (N_12012,N_11148,N_11589);
or U12013 (N_12013,N_11910,N_11639);
xor U12014 (N_12014,N_11741,N_11689);
xor U12015 (N_12015,N_11238,N_11306);
xnor U12016 (N_12016,N_11480,N_11265);
nor U12017 (N_12017,N_11184,N_11801);
or U12018 (N_12018,N_11938,N_11833);
nor U12019 (N_12019,N_11485,N_11745);
nor U12020 (N_12020,N_11178,N_11062);
or U12021 (N_12021,N_11083,N_11711);
nor U12022 (N_12022,N_11846,N_11431);
nand U12023 (N_12023,N_11021,N_11907);
or U12024 (N_12024,N_11517,N_11273);
nor U12025 (N_12025,N_11840,N_11379);
xor U12026 (N_12026,N_11091,N_11363);
and U12027 (N_12027,N_11961,N_11520);
nor U12028 (N_12028,N_11298,N_11610);
nor U12029 (N_12029,N_11784,N_11289);
xnor U12030 (N_12030,N_11429,N_11165);
or U12031 (N_12031,N_11685,N_11370);
nand U12032 (N_12032,N_11108,N_11218);
xnor U12033 (N_12033,N_11369,N_11339);
nor U12034 (N_12034,N_11879,N_11322);
or U12035 (N_12035,N_11920,N_11865);
nand U12036 (N_12036,N_11070,N_11876);
nand U12037 (N_12037,N_11034,N_11543);
or U12038 (N_12038,N_11964,N_11231);
and U12039 (N_12039,N_11584,N_11783);
nand U12040 (N_12040,N_11175,N_11510);
nand U12041 (N_12041,N_11951,N_11449);
nor U12042 (N_12042,N_11434,N_11808);
and U12043 (N_12043,N_11670,N_11387);
nand U12044 (N_12044,N_11285,N_11487);
and U12045 (N_12045,N_11612,N_11412);
and U12046 (N_12046,N_11287,N_11500);
or U12047 (N_12047,N_11877,N_11710);
nor U12048 (N_12048,N_11697,N_11382);
nor U12049 (N_12049,N_11019,N_11946);
and U12050 (N_12050,N_11630,N_11756);
xor U12051 (N_12051,N_11950,N_11341);
nand U12052 (N_12052,N_11416,N_11459);
nor U12053 (N_12053,N_11651,N_11551);
or U12054 (N_12054,N_11542,N_11059);
and U12055 (N_12055,N_11035,N_11181);
nand U12056 (N_12056,N_11658,N_11654);
xnor U12057 (N_12057,N_11171,N_11229);
nor U12058 (N_12058,N_11197,N_11672);
nand U12059 (N_12059,N_11465,N_11493);
xor U12060 (N_12060,N_11447,N_11696);
xnor U12061 (N_12061,N_11947,N_11509);
nand U12062 (N_12062,N_11361,N_11945);
and U12063 (N_12063,N_11110,N_11869);
nor U12064 (N_12064,N_11242,N_11693);
or U12065 (N_12065,N_11702,N_11668);
xnor U12066 (N_12066,N_11160,N_11841);
nand U12067 (N_12067,N_11297,N_11691);
nand U12068 (N_12068,N_11758,N_11475);
nor U12069 (N_12069,N_11448,N_11226);
or U12070 (N_12070,N_11031,N_11953);
nor U12071 (N_12071,N_11462,N_11954);
and U12072 (N_12072,N_11142,N_11003);
and U12073 (N_12073,N_11191,N_11221);
nand U12074 (N_12074,N_11202,N_11135);
or U12075 (N_12075,N_11056,N_11731);
or U12076 (N_12076,N_11319,N_11497);
nor U12077 (N_12077,N_11366,N_11707);
xnor U12078 (N_12078,N_11729,N_11652);
nand U12079 (N_12079,N_11504,N_11295);
and U12080 (N_12080,N_11327,N_11771);
nand U12081 (N_12081,N_11738,N_11944);
nor U12082 (N_12082,N_11757,N_11897);
or U12083 (N_12083,N_11036,N_11904);
xnor U12084 (N_12084,N_11296,N_11095);
or U12085 (N_12085,N_11455,N_11980);
nor U12086 (N_12086,N_11237,N_11214);
nor U12087 (N_12087,N_11208,N_11958);
nand U12088 (N_12088,N_11858,N_11787);
nor U12089 (N_12089,N_11167,N_11746);
xnor U12090 (N_12090,N_11762,N_11970);
nor U12091 (N_12091,N_11681,N_11033);
nor U12092 (N_12092,N_11502,N_11470);
xnor U12093 (N_12093,N_11852,N_11130);
nor U12094 (N_12094,N_11106,N_11818);
nand U12095 (N_12095,N_11179,N_11097);
or U12096 (N_12096,N_11843,N_11123);
or U12097 (N_12097,N_11701,N_11669);
nand U12098 (N_12098,N_11061,N_11280);
xnor U12099 (N_12099,N_11324,N_11122);
or U12100 (N_12100,N_11541,N_11022);
nor U12101 (N_12101,N_11495,N_11917);
nor U12102 (N_12102,N_11330,N_11891);
xor U12103 (N_12103,N_11402,N_11074);
nor U12104 (N_12104,N_11125,N_11870);
or U12105 (N_12105,N_11640,N_11973);
xnor U12106 (N_12106,N_11825,N_11454);
or U12107 (N_12107,N_11407,N_11260);
or U12108 (N_12108,N_11538,N_11760);
nor U12109 (N_12109,N_11988,N_11461);
or U12110 (N_12110,N_11507,N_11774);
xnor U12111 (N_12111,N_11545,N_11441);
and U12112 (N_12112,N_11633,N_11561);
xnor U12113 (N_12113,N_11992,N_11778);
xnor U12114 (N_12114,N_11092,N_11067);
xor U12115 (N_12115,N_11637,N_11578);
or U12116 (N_12116,N_11401,N_11650);
nor U12117 (N_12117,N_11850,N_11336);
and U12118 (N_12118,N_11041,N_11956);
and U12119 (N_12119,N_11820,N_11788);
xor U12120 (N_12120,N_11749,N_11017);
xnor U12121 (N_12121,N_11356,N_11537);
and U12122 (N_12122,N_11981,N_11423);
nand U12123 (N_12123,N_11700,N_11203);
xnor U12124 (N_12124,N_11884,N_11514);
or U12125 (N_12125,N_11395,N_11124);
nor U12126 (N_12126,N_11527,N_11805);
xnor U12127 (N_12127,N_11393,N_11299);
and U12128 (N_12128,N_11536,N_11655);
nand U12129 (N_12129,N_11119,N_11215);
nand U12130 (N_12130,N_11016,N_11570);
and U12131 (N_12131,N_11239,N_11780);
nand U12132 (N_12132,N_11752,N_11071);
or U12133 (N_12133,N_11560,N_11772);
or U12134 (N_12134,N_11329,N_11427);
or U12135 (N_12135,N_11666,N_11767);
nor U12136 (N_12136,N_11539,N_11557);
nand U12137 (N_12137,N_11066,N_11817);
and U12138 (N_12138,N_11253,N_11283);
or U12139 (N_12139,N_11107,N_11882);
nand U12140 (N_12140,N_11486,N_11896);
or U12141 (N_12141,N_11127,N_11883);
xor U12142 (N_12142,N_11862,N_11140);
and U12143 (N_12143,N_11667,N_11355);
or U12144 (N_12144,N_11813,N_11555);
nor U12145 (N_12145,N_11250,N_11360);
nand U12146 (N_12146,N_11321,N_11837);
nand U12147 (N_12147,N_11653,N_11247);
and U12148 (N_12148,N_11842,N_11574);
or U12149 (N_12149,N_11874,N_11799);
nand U12150 (N_12150,N_11469,N_11679);
nand U12151 (N_12151,N_11604,N_11501);
and U12152 (N_12152,N_11534,N_11976);
nor U12153 (N_12153,N_11742,N_11939);
nand U12154 (N_12154,N_11286,N_11608);
or U12155 (N_12155,N_11886,N_11080);
xnor U12156 (N_12156,N_11764,N_11887);
xor U12157 (N_12157,N_11635,N_11881);
or U12158 (N_12158,N_11332,N_11325);
nand U12159 (N_12159,N_11971,N_11582);
nand U12160 (N_12160,N_11444,N_11414);
nand U12161 (N_12161,N_11709,N_11525);
and U12162 (N_12162,N_11969,N_11819);
or U12163 (N_12163,N_11195,N_11391);
nand U12164 (N_12164,N_11528,N_11078);
and U12165 (N_12165,N_11479,N_11374);
nand U12166 (N_12166,N_11550,N_11262);
nor U12167 (N_12167,N_11699,N_11791);
or U12168 (N_12168,N_11999,N_11645);
or U12169 (N_12169,N_11058,N_11863);
xnor U12170 (N_12170,N_11312,N_11244);
or U12171 (N_12171,N_11935,N_11662);
nand U12172 (N_12172,N_11794,N_11400);
xor U12173 (N_12173,N_11418,N_11169);
xor U12174 (N_12174,N_11198,N_11173);
nand U12175 (N_12175,N_11713,N_11804);
nor U12176 (N_12176,N_11893,N_11723);
nor U12177 (N_12177,N_11753,N_11192);
and U12178 (N_12178,N_11878,N_11556);
and U12179 (N_12179,N_11340,N_11213);
xnor U12180 (N_12180,N_11795,N_11364);
nor U12181 (N_12181,N_11617,N_11380);
and U12182 (N_12182,N_11786,N_11420);
or U12183 (N_12183,N_11090,N_11088);
xor U12184 (N_12184,N_11585,N_11675);
xnor U12185 (N_12185,N_11187,N_11281);
and U12186 (N_12186,N_11763,N_11488);
or U12187 (N_12187,N_11089,N_11424);
xnor U12188 (N_12188,N_11075,N_11730);
xnor U12189 (N_12189,N_11288,N_11264);
nor U12190 (N_12190,N_11252,N_11628);
nand U12191 (N_12191,N_11845,N_11596);
nand U12192 (N_12192,N_11728,N_11766);
and U12193 (N_12193,N_11796,N_11245);
xnor U12194 (N_12194,N_11458,N_11233);
and U12195 (N_12195,N_11673,N_11368);
and U12196 (N_12196,N_11081,N_11750);
and U12197 (N_12197,N_11007,N_11718);
and U12198 (N_12198,N_11932,N_11188);
and U12199 (N_12199,N_11690,N_11384);
and U12200 (N_12200,N_11854,N_11346);
or U12201 (N_12201,N_11099,N_11905);
nand U12202 (N_12202,N_11962,N_11337);
xor U12203 (N_12203,N_11403,N_11398);
nand U12204 (N_12204,N_11712,N_11952);
xnor U12205 (N_12205,N_11616,N_11732);
and U12206 (N_12206,N_11595,N_11937);
or U12207 (N_12207,N_11816,N_11499);
nand U12208 (N_12208,N_11986,N_11522);
or U12209 (N_12209,N_11157,N_11292);
xor U12210 (N_12210,N_11269,N_11810);
xnor U12211 (N_12211,N_11782,N_11474);
nor U12212 (N_12212,N_11143,N_11761);
and U12213 (N_12213,N_11057,N_11684);
or U12214 (N_12214,N_11018,N_11743);
and U12215 (N_12215,N_11934,N_11831);
and U12216 (N_12216,N_11183,N_11591);
nand U12217 (N_12217,N_11204,N_11769);
or U12218 (N_12218,N_11072,N_11377);
nand U12219 (N_12219,N_11998,N_11776);
xor U12220 (N_12220,N_11120,N_11978);
or U12221 (N_12221,N_11503,N_11959);
nand U12222 (N_12222,N_11308,N_11186);
nand U12223 (N_12223,N_11172,N_11674);
nor U12224 (N_12224,N_11413,N_11572);
or U12225 (N_12225,N_11708,N_11030);
and U12226 (N_12226,N_11139,N_11466);
or U12227 (N_12227,N_11524,N_11464);
nand U12228 (N_12228,N_11008,N_11315);
and U12229 (N_12229,N_11193,N_11282);
nor U12230 (N_12230,N_11146,N_11311);
xnor U12231 (N_12231,N_11873,N_11686);
and U12232 (N_12232,N_11386,N_11331);
nor U12233 (N_12233,N_11740,N_11446);
or U12234 (N_12234,N_11261,N_11967);
nor U12235 (N_12235,N_11996,N_11232);
nor U12236 (N_12236,N_11276,N_11602);
nor U12237 (N_12237,N_11043,N_11457);
nand U12238 (N_12238,N_11415,N_11695);
and U12239 (N_12239,N_11358,N_11029);
xor U12240 (N_12240,N_11611,N_11736);
and U12241 (N_12241,N_11812,N_11147);
or U12242 (N_12242,N_11940,N_11647);
nor U12243 (N_12243,N_11848,N_11598);
and U12244 (N_12244,N_11579,N_11544);
or U12245 (N_12245,N_11344,N_11903);
nor U12246 (N_12246,N_11875,N_11859);
nand U12247 (N_12247,N_11348,N_11564);
nor U12248 (N_12248,N_11829,N_11836);
nor U12249 (N_12249,N_11046,N_11987);
and U12250 (N_12250,N_11832,N_11982);
nand U12251 (N_12251,N_11851,N_11154);
xor U12252 (N_12252,N_11605,N_11649);
or U12253 (N_12253,N_11523,N_11453);
or U12254 (N_12254,N_11236,N_11781);
and U12255 (N_12255,N_11467,N_11388);
nor U12256 (N_12256,N_11118,N_11580);
xnor U12257 (N_12257,N_11529,N_11622);
nor U12258 (N_12258,N_11634,N_11271);
xor U12259 (N_12259,N_11554,N_11835);
nor U12260 (N_12260,N_11592,N_11045);
nor U12261 (N_12261,N_11929,N_11293);
nor U12262 (N_12262,N_11603,N_11251);
and U12263 (N_12263,N_11040,N_11806);
xor U12264 (N_12264,N_11692,N_11015);
nor U12265 (N_12265,N_11532,N_11001);
nand U12266 (N_12266,N_11085,N_11716);
or U12267 (N_12267,N_11077,N_11822);
and U12268 (N_12268,N_11456,N_11627);
xnor U12269 (N_12269,N_11985,N_11924);
nor U12270 (N_12270,N_11737,N_11117);
nand U12271 (N_12271,N_11515,N_11868);
and U12272 (N_12272,N_11294,N_11472);
nand U12273 (N_12273,N_11463,N_11396);
nand U12274 (N_12274,N_11350,N_11722);
or U12275 (N_12275,N_11573,N_11301);
xor U12276 (N_12276,N_11618,N_11209);
or U12277 (N_12277,N_11249,N_11302);
xor U12278 (N_12278,N_11642,N_11826);
and U12279 (N_12279,N_11768,N_11751);
nor U12280 (N_12280,N_11367,N_11548);
nor U12281 (N_12281,N_11136,N_11126);
xor U12282 (N_12282,N_11880,N_11688);
nand U12283 (N_12283,N_11609,N_11005);
or U12284 (N_12284,N_11177,N_11552);
nor U12285 (N_12285,N_11397,N_11660);
nor U12286 (N_12286,N_11406,N_11216);
nor U12287 (N_12287,N_11727,N_11682);
and U12288 (N_12288,N_11145,N_11028);
and U12289 (N_12289,N_11275,N_11246);
or U12290 (N_12290,N_11342,N_11676);
nand U12291 (N_12291,N_11733,N_11912);
and U12292 (N_12292,N_11606,N_11254);
nor U12293 (N_12293,N_11051,N_11508);
or U12294 (N_12294,N_11871,N_11200);
xor U12295 (N_12295,N_11452,N_11316);
xor U12296 (N_12296,N_11044,N_11583);
nor U12297 (N_12297,N_11211,N_11168);
nand U12298 (N_12298,N_11274,N_11365);
or U12299 (N_12299,N_11671,N_11053);
nor U12300 (N_12300,N_11563,N_11482);
and U12301 (N_12301,N_11349,N_11565);
or U12302 (N_12302,N_11586,N_11161);
nor U12303 (N_12303,N_11185,N_11176);
xnor U12304 (N_12304,N_11011,N_11323);
xnor U12305 (N_12305,N_11137,N_11558);
xor U12306 (N_12306,N_11755,N_11291);
nor U12307 (N_12307,N_11278,N_11914);
xor U12308 (N_12308,N_11677,N_11720);
xor U12309 (N_12309,N_11948,N_11491);
and U12310 (N_12310,N_11855,N_11659);
xnor U12311 (N_12311,N_11159,N_11392);
nand U12312 (N_12312,N_11490,N_11039);
nand U12313 (N_12313,N_11646,N_11966);
or U12314 (N_12314,N_11343,N_11590);
nor U12315 (N_12315,N_11984,N_11255);
or U12316 (N_12316,N_11000,N_11553);
nand U12317 (N_12317,N_11257,N_11521);
and U12318 (N_12318,N_11477,N_11864);
or U12319 (N_12319,N_11644,N_11112);
nand U12320 (N_12320,N_11121,N_11305);
and U12321 (N_12321,N_11705,N_11638);
and U12322 (N_12322,N_11827,N_11404);
nor U12323 (N_12323,N_11290,N_11259);
and U12324 (N_12324,N_11613,N_11450);
xor U12325 (N_12325,N_11084,N_11484);
nand U12326 (N_12326,N_11196,N_11547);
nand U12327 (N_12327,N_11389,N_11351);
xnor U12328 (N_12328,N_11777,N_11133);
nand U12329 (N_12329,N_11114,N_11908);
or U12330 (N_12330,N_11714,N_11993);
xor U12331 (N_12331,N_11928,N_11531);
nor U12332 (N_12332,N_11180,N_11152);
xor U12333 (N_12333,N_11132,N_11607);
nor U12334 (N_12334,N_11974,N_11698);
and U12335 (N_12335,N_11026,N_11381);
nor U12336 (N_12336,N_11923,N_11076);
nor U12337 (N_12337,N_11437,N_11949);
and U12338 (N_12338,N_11093,N_11199);
or U12339 (N_12339,N_11931,N_11086);
nand U12340 (N_12340,N_11012,N_11773);
xnor U12341 (N_12341,N_11440,N_11048);
or U12342 (N_12342,N_11207,N_11892);
nand U12343 (N_12343,N_11936,N_11739);
or U12344 (N_12344,N_11494,N_11020);
nor U12345 (N_12345,N_11240,N_11919);
nand U12346 (N_12346,N_11797,N_11115);
nand U12347 (N_12347,N_11513,N_11798);
xnor U12348 (N_12348,N_11526,N_11433);
and U12349 (N_12349,N_11861,N_11535);
nand U12350 (N_12350,N_11439,N_11182);
xnor U12351 (N_12351,N_11128,N_11065);
xor U12352 (N_12352,N_11568,N_11037);
or U12353 (N_12353,N_11098,N_11587);
nor U12354 (N_12354,N_11313,N_11930);
nand U12355 (N_12355,N_11793,N_11505);
xor U12356 (N_12356,N_11915,N_11432);
nor U12357 (N_12357,N_11156,N_11303);
and U12358 (N_12358,N_11747,N_11963);
xor U12359 (N_12359,N_11941,N_11201);
nor U12360 (N_12360,N_11038,N_11476);
or U12361 (N_12361,N_11857,N_11588);
and U12362 (N_12362,N_11228,N_11814);
nand U12363 (N_12363,N_11158,N_11506);
nor U12364 (N_12364,N_11821,N_11965);
xor U12365 (N_12365,N_11990,N_11995);
nand U12366 (N_12366,N_11900,N_11489);
and U12367 (N_12367,N_11885,N_11230);
xnor U12368 (N_12368,N_11025,N_11643);
nor U12369 (N_12369,N_11405,N_11663);
nor U12370 (N_12370,N_11721,N_11770);
or U12371 (N_12371,N_11047,N_11748);
nor U12372 (N_12372,N_11134,N_11661);
nor U12373 (N_12373,N_11997,N_11409);
nor U12374 (N_12374,N_11131,N_11419);
nand U12375 (N_12375,N_11268,N_11096);
or U12376 (N_12376,N_11866,N_11889);
or U12377 (N_12377,N_11577,N_11425);
and U12378 (N_12378,N_11581,N_11518);
xnor U12379 (N_12379,N_11050,N_11068);
or U12380 (N_12380,N_11631,N_11478);
and U12381 (N_12381,N_11779,N_11004);
and U12382 (N_12382,N_11378,N_11073);
xnor U12383 (N_12383,N_11849,N_11334);
xor U12384 (N_12384,N_11105,N_11599);
and U12385 (N_12385,N_11223,N_11922);
xnor U12386 (N_12386,N_11422,N_11438);
or U12387 (N_12387,N_11354,N_11023);
and U12388 (N_12388,N_11263,N_11894);
nor U12389 (N_12389,N_11600,N_11704);
or U12390 (N_12390,N_11064,N_11623);
nor U12391 (N_12391,N_11847,N_11943);
nor U12392 (N_12392,N_11918,N_11435);
or U12393 (N_12393,N_11765,N_11373);
nand U12394 (N_12394,N_11149,N_11803);
or U12395 (N_12395,N_11706,N_11362);
nand U12396 (N_12396,N_11925,N_11909);
nand U12397 (N_12397,N_11807,N_11724);
or U12398 (N_12398,N_11898,N_11460);
xnor U12399 (N_12399,N_11678,N_11069);
xnor U12400 (N_12400,N_11926,N_11266);
xor U12401 (N_12401,N_11619,N_11625);
or U12402 (N_12402,N_11615,N_11853);
and U12403 (N_12403,N_11626,N_11789);
or U12404 (N_12404,N_11735,N_11258);
xnor U12405 (N_12405,N_11436,N_11815);
xor U12406 (N_12406,N_11530,N_11277);
nand U12407 (N_12407,N_11844,N_11972);
nor U12408 (N_12408,N_11656,N_11593);
or U12409 (N_12409,N_11913,N_11775);
nor U12410 (N_12410,N_11683,N_11594);
xor U12411 (N_12411,N_11426,N_11575);
nor U12412 (N_12412,N_11024,N_11307);
xnor U12413 (N_12413,N_11310,N_11353);
nor U12414 (N_12414,N_11540,N_11217);
nor U12415 (N_12415,N_11256,N_11333);
xor U12416 (N_12416,N_11009,N_11687);
nor U12417 (N_12417,N_11335,N_11206);
or U12418 (N_12418,N_11189,N_11357);
nand U12419 (N_12419,N_11823,N_11241);
or U12420 (N_12420,N_11054,N_11468);
and U12421 (N_12421,N_11856,N_11006);
or U12422 (N_12422,N_11895,N_11442);
xnor U12423 (N_12423,N_11279,N_11571);
nand U12424 (N_12424,N_11546,N_11496);
and U12425 (N_12425,N_11138,N_11411);
nand U12426 (N_12426,N_11100,N_11566);
and U12427 (N_12427,N_11079,N_11838);
xnor U12428 (N_12428,N_11624,N_11430);
xor U12429 (N_12429,N_11010,N_11481);
nand U12430 (N_12430,N_11272,N_11960);
and U12431 (N_12431,N_11155,N_11060);
or U12432 (N_12432,N_11144,N_11087);
nand U12433 (N_12433,N_11284,N_11890);
nand U12434 (N_12434,N_11399,N_11921);
nor U12435 (N_12435,N_11790,N_11314);
xnor U12436 (N_12436,N_11394,N_11680);
and U12437 (N_12437,N_11927,N_11328);
xor U12438 (N_12438,N_11428,N_11957);
and U12439 (N_12439,N_11225,N_11498);
or U12440 (N_12440,N_11014,N_11170);
nand U12441 (N_12441,N_11163,N_11318);
nor U12442 (N_12442,N_11326,N_11212);
xnor U12443 (N_12443,N_11153,N_11052);
xor U12444 (N_12444,N_11220,N_11664);
or U12445 (N_12445,N_11375,N_11785);
and U12446 (N_12446,N_11443,N_11243);
or U12447 (N_12447,N_11445,N_11151);
and U12448 (N_12448,N_11549,N_11632);
nor U12449 (N_12449,N_11383,N_11562);
nor U12450 (N_12450,N_11224,N_11473);
nand U12451 (N_12451,N_11533,N_11104);
or U12452 (N_12452,N_11744,N_11809);
and U12453 (N_12453,N_11597,N_11270);
and U12454 (N_12454,N_11002,N_11719);
and U12455 (N_12455,N_11162,N_11109);
xnor U12456 (N_12456,N_11032,N_11227);
or U12457 (N_12457,N_11304,N_11975);
or U12458 (N_12458,N_11063,N_11703);
nand U12459 (N_12459,N_11300,N_11129);
or U12460 (N_12460,N_11267,N_11235);
nor U12461 (N_12461,N_11150,N_11103);
xor U12462 (N_12462,N_11390,N_11867);
xnor U12463 (N_12463,N_11614,N_11968);
nand U12464 (N_12464,N_11994,N_11977);
and U12465 (N_12465,N_11013,N_11111);
xor U12466 (N_12466,N_11899,N_11694);
nor U12467 (N_12467,N_11116,N_11164);
and U12468 (N_12468,N_11371,N_11210);
or U12469 (N_12469,N_11824,N_11027);
nor U12470 (N_12470,N_11906,N_11317);
nor U12471 (N_12471,N_11802,N_11205);
or U12472 (N_12472,N_11911,N_11641);
nand U12473 (N_12473,N_11410,N_11338);
and U12474 (N_12474,N_11601,N_11174);
and U12475 (N_12475,N_11376,N_11141);
nor U12476 (N_12476,N_11811,N_11942);
nand U12477 (N_12477,N_11901,N_11754);
or U12478 (N_12478,N_11872,N_11102);
nand U12479 (N_12479,N_11042,N_11516);
or U12480 (N_12480,N_11792,N_11347);
nor U12481 (N_12481,N_11860,N_11979);
xor U12482 (N_12482,N_11715,N_11621);
or U12483 (N_12483,N_11359,N_11725);
nor U12484 (N_12484,N_11989,N_11094);
nor U12485 (N_12485,N_11902,N_11055);
xnor U12486 (N_12486,N_11830,N_11492);
and U12487 (N_12487,N_11933,N_11049);
nand U12488 (N_12488,N_11888,N_11717);
and U12489 (N_12489,N_11559,N_11834);
xnor U12490 (N_12490,N_11620,N_11101);
nand U12491 (N_12491,N_11113,N_11345);
xnor U12492 (N_12492,N_11983,N_11417);
nor U12493 (N_12493,N_11166,N_11352);
nor U12494 (N_12494,N_11194,N_11471);
nand U12495 (N_12495,N_11320,N_11734);
or U12496 (N_12496,N_11222,N_11828);
or U12497 (N_12497,N_11190,N_11916);
or U12498 (N_12498,N_11082,N_11234);
and U12499 (N_12499,N_11372,N_11451);
or U12500 (N_12500,N_11898,N_11650);
xor U12501 (N_12501,N_11836,N_11999);
and U12502 (N_12502,N_11037,N_11839);
nor U12503 (N_12503,N_11728,N_11544);
nor U12504 (N_12504,N_11695,N_11370);
or U12505 (N_12505,N_11406,N_11674);
and U12506 (N_12506,N_11512,N_11288);
nor U12507 (N_12507,N_11754,N_11575);
or U12508 (N_12508,N_11805,N_11187);
or U12509 (N_12509,N_11484,N_11097);
and U12510 (N_12510,N_11510,N_11849);
nand U12511 (N_12511,N_11802,N_11157);
or U12512 (N_12512,N_11562,N_11674);
xor U12513 (N_12513,N_11496,N_11832);
or U12514 (N_12514,N_11307,N_11805);
or U12515 (N_12515,N_11906,N_11560);
nor U12516 (N_12516,N_11230,N_11270);
xnor U12517 (N_12517,N_11207,N_11346);
nand U12518 (N_12518,N_11869,N_11928);
or U12519 (N_12519,N_11776,N_11165);
nor U12520 (N_12520,N_11054,N_11107);
xor U12521 (N_12521,N_11427,N_11753);
nor U12522 (N_12522,N_11440,N_11819);
xor U12523 (N_12523,N_11183,N_11633);
or U12524 (N_12524,N_11029,N_11047);
xnor U12525 (N_12525,N_11198,N_11081);
or U12526 (N_12526,N_11316,N_11511);
xnor U12527 (N_12527,N_11439,N_11925);
nor U12528 (N_12528,N_11992,N_11473);
nand U12529 (N_12529,N_11875,N_11824);
xor U12530 (N_12530,N_11476,N_11567);
or U12531 (N_12531,N_11956,N_11812);
and U12532 (N_12532,N_11396,N_11066);
nand U12533 (N_12533,N_11633,N_11497);
and U12534 (N_12534,N_11114,N_11143);
nor U12535 (N_12535,N_11052,N_11519);
and U12536 (N_12536,N_11765,N_11135);
nand U12537 (N_12537,N_11775,N_11879);
nand U12538 (N_12538,N_11773,N_11147);
nand U12539 (N_12539,N_11307,N_11723);
and U12540 (N_12540,N_11679,N_11842);
nor U12541 (N_12541,N_11019,N_11593);
xnor U12542 (N_12542,N_11145,N_11931);
xnor U12543 (N_12543,N_11399,N_11511);
and U12544 (N_12544,N_11841,N_11278);
and U12545 (N_12545,N_11657,N_11235);
nand U12546 (N_12546,N_11277,N_11765);
xor U12547 (N_12547,N_11062,N_11342);
and U12548 (N_12548,N_11742,N_11242);
and U12549 (N_12549,N_11024,N_11810);
nor U12550 (N_12550,N_11913,N_11258);
xor U12551 (N_12551,N_11950,N_11276);
nor U12552 (N_12552,N_11461,N_11387);
nor U12553 (N_12553,N_11192,N_11046);
and U12554 (N_12554,N_11738,N_11465);
xnor U12555 (N_12555,N_11102,N_11038);
nor U12556 (N_12556,N_11054,N_11425);
xor U12557 (N_12557,N_11105,N_11848);
and U12558 (N_12558,N_11572,N_11218);
nor U12559 (N_12559,N_11697,N_11518);
or U12560 (N_12560,N_11283,N_11128);
and U12561 (N_12561,N_11024,N_11111);
nor U12562 (N_12562,N_11445,N_11145);
nand U12563 (N_12563,N_11603,N_11169);
and U12564 (N_12564,N_11885,N_11315);
or U12565 (N_12565,N_11384,N_11446);
nor U12566 (N_12566,N_11887,N_11347);
xnor U12567 (N_12567,N_11685,N_11932);
or U12568 (N_12568,N_11081,N_11899);
nor U12569 (N_12569,N_11857,N_11289);
nand U12570 (N_12570,N_11271,N_11182);
or U12571 (N_12571,N_11912,N_11139);
and U12572 (N_12572,N_11507,N_11416);
xor U12573 (N_12573,N_11347,N_11046);
nor U12574 (N_12574,N_11270,N_11682);
xnor U12575 (N_12575,N_11715,N_11665);
or U12576 (N_12576,N_11912,N_11089);
and U12577 (N_12577,N_11009,N_11135);
or U12578 (N_12578,N_11201,N_11205);
and U12579 (N_12579,N_11818,N_11710);
nor U12580 (N_12580,N_11762,N_11660);
or U12581 (N_12581,N_11815,N_11218);
and U12582 (N_12582,N_11272,N_11320);
xnor U12583 (N_12583,N_11594,N_11222);
and U12584 (N_12584,N_11338,N_11152);
and U12585 (N_12585,N_11293,N_11875);
nor U12586 (N_12586,N_11278,N_11020);
xnor U12587 (N_12587,N_11417,N_11499);
or U12588 (N_12588,N_11060,N_11192);
or U12589 (N_12589,N_11192,N_11708);
and U12590 (N_12590,N_11867,N_11073);
nand U12591 (N_12591,N_11866,N_11227);
or U12592 (N_12592,N_11940,N_11324);
and U12593 (N_12593,N_11402,N_11419);
xor U12594 (N_12594,N_11375,N_11319);
and U12595 (N_12595,N_11980,N_11128);
nand U12596 (N_12596,N_11153,N_11227);
and U12597 (N_12597,N_11625,N_11401);
or U12598 (N_12598,N_11298,N_11408);
and U12599 (N_12599,N_11206,N_11579);
and U12600 (N_12600,N_11531,N_11919);
or U12601 (N_12601,N_11909,N_11974);
or U12602 (N_12602,N_11164,N_11717);
nand U12603 (N_12603,N_11273,N_11740);
xnor U12604 (N_12604,N_11846,N_11352);
or U12605 (N_12605,N_11540,N_11655);
and U12606 (N_12606,N_11790,N_11692);
or U12607 (N_12607,N_11410,N_11513);
or U12608 (N_12608,N_11439,N_11808);
and U12609 (N_12609,N_11786,N_11983);
nand U12610 (N_12610,N_11789,N_11774);
and U12611 (N_12611,N_11226,N_11845);
nor U12612 (N_12612,N_11605,N_11816);
and U12613 (N_12613,N_11572,N_11277);
nor U12614 (N_12614,N_11071,N_11212);
nand U12615 (N_12615,N_11198,N_11725);
xor U12616 (N_12616,N_11192,N_11463);
nand U12617 (N_12617,N_11197,N_11420);
nor U12618 (N_12618,N_11106,N_11821);
or U12619 (N_12619,N_11319,N_11002);
nor U12620 (N_12620,N_11673,N_11292);
or U12621 (N_12621,N_11646,N_11423);
and U12622 (N_12622,N_11893,N_11878);
nand U12623 (N_12623,N_11406,N_11100);
or U12624 (N_12624,N_11298,N_11062);
xor U12625 (N_12625,N_11862,N_11660);
xnor U12626 (N_12626,N_11658,N_11326);
nor U12627 (N_12627,N_11872,N_11396);
xnor U12628 (N_12628,N_11589,N_11849);
nor U12629 (N_12629,N_11189,N_11443);
nor U12630 (N_12630,N_11222,N_11352);
nand U12631 (N_12631,N_11730,N_11922);
nor U12632 (N_12632,N_11780,N_11205);
or U12633 (N_12633,N_11267,N_11825);
nand U12634 (N_12634,N_11017,N_11097);
and U12635 (N_12635,N_11767,N_11993);
xor U12636 (N_12636,N_11258,N_11255);
or U12637 (N_12637,N_11347,N_11277);
nor U12638 (N_12638,N_11528,N_11531);
and U12639 (N_12639,N_11622,N_11048);
nand U12640 (N_12640,N_11597,N_11509);
and U12641 (N_12641,N_11531,N_11367);
nor U12642 (N_12642,N_11439,N_11869);
nand U12643 (N_12643,N_11339,N_11435);
xnor U12644 (N_12644,N_11428,N_11191);
xor U12645 (N_12645,N_11059,N_11528);
and U12646 (N_12646,N_11403,N_11580);
xnor U12647 (N_12647,N_11286,N_11542);
and U12648 (N_12648,N_11224,N_11105);
nor U12649 (N_12649,N_11639,N_11736);
or U12650 (N_12650,N_11021,N_11018);
and U12651 (N_12651,N_11956,N_11584);
xnor U12652 (N_12652,N_11265,N_11207);
nor U12653 (N_12653,N_11740,N_11774);
xnor U12654 (N_12654,N_11033,N_11661);
xnor U12655 (N_12655,N_11210,N_11369);
and U12656 (N_12656,N_11500,N_11471);
nand U12657 (N_12657,N_11382,N_11506);
nand U12658 (N_12658,N_11844,N_11185);
nor U12659 (N_12659,N_11784,N_11595);
and U12660 (N_12660,N_11659,N_11296);
xnor U12661 (N_12661,N_11024,N_11878);
xnor U12662 (N_12662,N_11868,N_11687);
xor U12663 (N_12663,N_11266,N_11294);
xnor U12664 (N_12664,N_11402,N_11009);
and U12665 (N_12665,N_11110,N_11685);
or U12666 (N_12666,N_11038,N_11330);
nand U12667 (N_12667,N_11787,N_11326);
xor U12668 (N_12668,N_11342,N_11450);
nand U12669 (N_12669,N_11200,N_11128);
xnor U12670 (N_12670,N_11648,N_11836);
or U12671 (N_12671,N_11965,N_11725);
nor U12672 (N_12672,N_11647,N_11600);
xor U12673 (N_12673,N_11400,N_11993);
nor U12674 (N_12674,N_11832,N_11764);
xnor U12675 (N_12675,N_11146,N_11809);
or U12676 (N_12676,N_11203,N_11814);
nand U12677 (N_12677,N_11794,N_11152);
xnor U12678 (N_12678,N_11830,N_11128);
or U12679 (N_12679,N_11382,N_11680);
xnor U12680 (N_12680,N_11049,N_11354);
or U12681 (N_12681,N_11585,N_11905);
nor U12682 (N_12682,N_11506,N_11352);
nand U12683 (N_12683,N_11919,N_11347);
and U12684 (N_12684,N_11127,N_11500);
nor U12685 (N_12685,N_11168,N_11605);
nand U12686 (N_12686,N_11981,N_11454);
nand U12687 (N_12687,N_11582,N_11399);
nand U12688 (N_12688,N_11496,N_11021);
nor U12689 (N_12689,N_11619,N_11802);
xor U12690 (N_12690,N_11900,N_11540);
xor U12691 (N_12691,N_11772,N_11013);
or U12692 (N_12692,N_11821,N_11767);
nor U12693 (N_12693,N_11274,N_11399);
xor U12694 (N_12694,N_11065,N_11166);
nand U12695 (N_12695,N_11593,N_11410);
nand U12696 (N_12696,N_11278,N_11645);
nor U12697 (N_12697,N_11906,N_11484);
and U12698 (N_12698,N_11417,N_11695);
nor U12699 (N_12699,N_11730,N_11602);
and U12700 (N_12700,N_11220,N_11313);
nor U12701 (N_12701,N_11507,N_11934);
nand U12702 (N_12702,N_11166,N_11553);
or U12703 (N_12703,N_11618,N_11935);
and U12704 (N_12704,N_11039,N_11627);
or U12705 (N_12705,N_11357,N_11790);
or U12706 (N_12706,N_11338,N_11129);
or U12707 (N_12707,N_11615,N_11788);
xnor U12708 (N_12708,N_11727,N_11678);
and U12709 (N_12709,N_11215,N_11795);
or U12710 (N_12710,N_11945,N_11013);
xor U12711 (N_12711,N_11912,N_11747);
nor U12712 (N_12712,N_11930,N_11987);
nand U12713 (N_12713,N_11267,N_11184);
nor U12714 (N_12714,N_11034,N_11724);
and U12715 (N_12715,N_11974,N_11164);
or U12716 (N_12716,N_11832,N_11224);
nand U12717 (N_12717,N_11296,N_11609);
or U12718 (N_12718,N_11870,N_11311);
nand U12719 (N_12719,N_11454,N_11897);
nand U12720 (N_12720,N_11405,N_11006);
xnor U12721 (N_12721,N_11964,N_11764);
and U12722 (N_12722,N_11983,N_11129);
xor U12723 (N_12723,N_11516,N_11045);
nor U12724 (N_12724,N_11191,N_11420);
nor U12725 (N_12725,N_11045,N_11141);
nand U12726 (N_12726,N_11529,N_11260);
or U12727 (N_12727,N_11387,N_11421);
nor U12728 (N_12728,N_11822,N_11747);
nor U12729 (N_12729,N_11068,N_11755);
nor U12730 (N_12730,N_11948,N_11165);
nand U12731 (N_12731,N_11703,N_11548);
nand U12732 (N_12732,N_11725,N_11702);
nand U12733 (N_12733,N_11657,N_11553);
and U12734 (N_12734,N_11281,N_11443);
or U12735 (N_12735,N_11405,N_11590);
xor U12736 (N_12736,N_11658,N_11378);
and U12737 (N_12737,N_11947,N_11055);
xnor U12738 (N_12738,N_11337,N_11154);
nor U12739 (N_12739,N_11213,N_11210);
and U12740 (N_12740,N_11101,N_11980);
xor U12741 (N_12741,N_11586,N_11084);
or U12742 (N_12742,N_11190,N_11325);
nor U12743 (N_12743,N_11554,N_11920);
nor U12744 (N_12744,N_11070,N_11449);
nor U12745 (N_12745,N_11779,N_11175);
or U12746 (N_12746,N_11186,N_11367);
nand U12747 (N_12747,N_11356,N_11708);
or U12748 (N_12748,N_11264,N_11882);
nor U12749 (N_12749,N_11649,N_11002);
nor U12750 (N_12750,N_11009,N_11474);
and U12751 (N_12751,N_11524,N_11385);
xor U12752 (N_12752,N_11073,N_11741);
xnor U12753 (N_12753,N_11689,N_11494);
xor U12754 (N_12754,N_11400,N_11840);
nor U12755 (N_12755,N_11837,N_11023);
or U12756 (N_12756,N_11409,N_11120);
xor U12757 (N_12757,N_11590,N_11861);
and U12758 (N_12758,N_11669,N_11974);
nand U12759 (N_12759,N_11536,N_11819);
or U12760 (N_12760,N_11906,N_11210);
or U12761 (N_12761,N_11173,N_11863);
xor U12762 (N_12762,N_11126,N_11400);
nand U12763 (N_12763,N_11305,N_11448);
nand U12764 (N_12764,N_11844,N_11298);
xor U12765 (N_12765,N_11476,N_11674);
nor U12766 (N_12766,N_11103,N_11700);
or U12767 (N_12767,N_11035,N_11989);
xor U12768 (N_12768,N_11884,N_11008);
nor U12769 (N_12769,N_11989,N_11241);
xor U12770 (N_12770,N_11474,N_11043);
nor U12771 (N_12771,N_11300,N_11687);
and U12772 (N_12772,N_11383,N_11016);
or U12773 (N_12773,N_11224,N_11528);
and U12774 (N_12774,N_11651,N_11178);
and U12775 (N_12775,N_11977,N_11197);
nor U12776 (N_12776,N_11463,N_11921);
nor U12777 (N_12777,N_11096,N_11449);
nor U12778 (N_12778,N_11621,N_11736);
nand U12779 (N_12779,N_11655,N_11973);
nor U12780 (N_12780,N_11448,N_11975);
xnor U12781 (N_12781,N_11689,N_11634);
or U12782 (N_12782,N_11186,N_11615);
and U12783 (N_12783,N_11753,N_11777);
xnor U12784 (N_12784,N_11387,N_11033);
xor U12785 (N_12785,N_11662,N_11375);
or U12786 (N_12786,N_11002,N_11908);
or U12787 (N_12787,N_11898,N_11567);
and U12788 (N_12788,N_11248,N_11826);
nor U12789 (N_12789,N_11949,N_11569);
or U12790 (N_12790,N_11716,N_11293);
and U12791 (N_12791,N_11482,N_11069);
nand U12792 (N_12792,N_11998,N_11690);
or U12793 (N_12793,N_11531,N_11584);
nor U12794 (N_12794,N_11305,N_11642);
nor U12795 (N_12795,N_11051,N_11725);
xnor U12796 (N_12796,N_11412,N_11537);
or U12797 (N_12797,N_11579,N_11415);
nand U12798 (N_12798,N_11120,N_11670);
xnor U12799 (N_12799,N_11805,N_11145);
nor U12800 (N_12800,N_11546,N_11164);
nand U12801 (N_12801,N_11015,N_11576);
nor U12802 (N_12802,N_11941,N_11659);
nand U12803 (N_12803,N_11851,N_11846);
or U12804 (N_12804,N_11016,N_11140);
nand U12805 (N_12805,N_11954,N_11428);
xor U12806 (N_12806,N_11663,N_11641);
nand U12807 (N_12807,N_11037,N_11277);
or U12808 (N_12808,N_11340,N_11023);
nand U12809 (N_12809,N_11560,N_11002);
nor U12810 (N_12810,N_11296,N_11103);
xor U12811 (N_12811,N_11098,N_11176);
xor U12812 (N_12812,N_11775,N_11572);
xnor U12813 (N_12813,N_11285,N_11024);
and U12814 (N_12814,N_11027,N_11051);
and U12815 (N_12815,N_11253,N_11585);
or U12816 (N_12816,N_11498,N_11902);
or U12817 (N_12817,N_11399,N_11533);
or U12818 (N_12818,N_11968,N_11619);
nor U12819 (N_12819,N_11865,N_11078);
xor U12820 (N_12820,N_11780,N_11630);
and U12821 (N_12821,N_11731,N_11144);
and U12822 (N_12822,N_11926,N_11368);
nor U12823 (N_12823,N_11517,N_11101);
xor U12824 (N_12824,N_11350,N_11767);
xnor U12825 (N_12825,N_11008,N_11774);
xnor U12826 (N_12826,N_11180,N_11867);
or U12827 (N_12827,N_11816,N_11486);
and U12828 (N_12828,N_11481,N_11191);
nor U12829 (N_12829,N_11284,N_11794);
and U12830 (N_12830,N_11338,N_11892);
xnor U12831 (N_12831,N_11361,N_11102);
nor U12832 (N_12832,N_11195,N_11318);
and U12833 (N_12833,N_11041,N_11007);
xor U12834 (N_12834,N_11449,N_11028);
xor U12835 (N_12835,N_11007,N_11777);
or U12836 (N_12836,N_11938,N_11140);
or U12837 (N_12837,N_11051,N_11542);
or U12838 (N_12838,N_11269,N_11938);
nor U12839 (N_12839,N_11502,N_11003);
nor U12840 (N_12840,N_11080,N_11065);
nand U12841 (N_12841,N_11076,N_11536);
nand U12842 (N_12842,N_11341,N_11375);
or U12843 (N_12843,N_11419,N_11518);
xor U12844 (N_12844,N_11404,N_11601);
nand U12845 (N_12845,N_11400,N_11644);
or U12846 (N_12846,N_11564,N_11954);
nand U12847 (N_12847,N_11179,N_11815);
nand U12848 (N_12848,N_11494,N_11382);
and U12849 (N_12849,N_11251,N_11241);
nand U12850 (N_12850,N_11054,N_11843);
or U12851 (N_12851,N_11507,N_11506);
xor U12852 (N_12852,N_11446,N_11959);
nor U12853 (N_12853,N_11201,N_11946);
nand U12854 (N_12854,N_11349,N_11634);
nor U12855 (N_12855,N_11872,N_11640);
or U12856 (N_12856,N_11950,N_11408);
or U12857 (N_12857,N_11917,N_11301);
and U12858 (N_12858,N_11126,N_11666);
xnor U12859 (N_12859,N_11672,N_11662);
and U12860 (N_12860,N_11018,N_11274);
and U12861 (N_12861,N_11512,N_11982);
or U12862 (N_12862,N_11981,N_11185);
xnor U12863 (N_12863,N_11481,N_11214);
or U12864 (N_12864,N_11742,N_11645);
xnor U12865 (N_12865,N_11572,N_11222);
nor U12866 (N_12866,N_11482,N_11798);
or U12867 (N_12867,N_11072,N_11355);
nor U12868 (N_12868,N_11128,N_11326);
xor U12869 (N_12869,N_11806,N_11082);
nor U12870 (N_12870,N_11518,N_11407);
xnor U12871 (N_12871,N_11726,N_11915);
or U12872 (N_12872,N_11218,N_11216);
nand U12873 (N_12873,N_11499,N_11354);
nand U12874 (N_12874,N_11793,N_11490);
nand U12875 (N_12875,N_11714,N_11185);
and U12876 (N_12876,N_11929,N_11787);
or U12877 (N_12877,N_11086,N_11040);
and U12878 (N_12878,N_11953,N_11049);
nor U12879 (N_12879,N_11546,N_11186);
xnor U12880 (N_12880,N_11998,N_11367);
nand U12881 (N_12881,N_11059,N_11420);
nand U12882 (N_12882,N_11584,N_11012);
xor U12883 (N_12883,N_11367,N_11775);
and U12884 (N_12884,N_11372,N_11171);
nor U12885 (N_12885,N_11647,N_11137);
xor U12886 (N_12886,N_11189,N_11140);
or U12887 (N_12887,N_11991,N_11675);
xnor U12888 (N_12888,N_11319,N_11861);
or U12889 (N_12889,N_11970,N_11412);
xnor U12890 (N_12890,N_11276,N_11037);
and U12891 (N_12891,N_11939,N_11596);
nor U12892 (N_12892,N_11940,N_11093);
and U12893 (N_12893,N_11395,N_11059);
or U12894 (N_12894,N_11447,N_11248);
or U12895 (N_12895,N_11388,N_11828);
nand U12896 (N_12896,N_11486,N_11501);
nand U12897 (N_12897,N_11205,N_11733);
nand U12898 (N_12898,N_11646,N_11014);
or U12899 (N_12899,N_11680,N_11831);
nor U12900 (N_12900,N_11272,N_11734);
and U12901 (N_12901,N_11851,N_11929);
nor U12902 (N_12902,N_11706,N_11216);
nand U12903 (N_12903,N_11025,N_11400);
or U12904 (N_12904,N_11542,N_11925);
nor U12905 (N_12905,N_11414,N_11340);
nor U12906 (N_12906,N_11414,N_11286);
nor U12907 (N_12907,N_11800,N_11036);
or U12908 (N_12908,N_11379,N_11662);
nand U12909 (N_12909,N_11235,N_11647);
and U12910 (N_12910,N_11189,N_11067);
nand U12911 (N_12911,N_11450,N_11384);
xor U12912 (N_12912,N_11639,N_11521);
nand U12913 (N_12913,N_11008,N_11090);
xnor U12914 (N_12914,N_11103,N_11091);
and U12915 (N_12915,N_11336,N_11299);
nor U12916 (N_12916,N_11352,N_11625);
nor U12917 (N_12917,N_11569,N_11726);
xor U12918 (N_12918,N_11575,N_11077);
nand U12919 (N_12919,N_11412,N_11303);
and U12920 (N_12920,N_11934,N_11266);
xnor U12921 (N_12921,N_11288,N_11797);
or U12922 (N_12922,N_11272,N_11217);
nor U12923 (N_12923,N_11710,N_11692);
nor U12924 (N_12924,N_11387,N_11616);
nor U12925 (N_12925,N_11001,N_11315);
xnor U12926 (N_12926,N_11660,N_11226);
xor U12927 (N_12927,N_11681,N_11353);
xnor U12928 (N_12928,N_11367,N_11216);
nand U12929 (N_12929,N_11263,N_11656);
or U12930 (N_12930,N_11025,N_11967);
nor U12931 (N_12931,N_11412,N_11801);
and U12932 (N_12932,N_11477,N_11023);
xnor U12933 (N_12933,N_11495,N_11373);
and U12934 (N_12934,N_11128,N_11076);
or U12935 (N_12935,N_11678,N_11545);
or U12936 (N_12936,N_11396,N_11960);
and U12937 (N_12937,N_11585,N_11940);
nor U12938 (N_12938,N_11158,N_11447);
nor U12939 (N_12939,N_11648,N_11839);
nor U12940 (N_12940,N_11507,N_11564);
nor U12941 (N_12941,N_11674,N_11947);
nor U12942 (N_12942,N_11391,N_11193);
nor U12943 (N_12943,N_11884,N_11557);
or U12944 (N_12944,N_11144,N_11720);
and U12945 (N_12945,N_11656,N_11925);
and U12946 (N_12946,N_11476,N_11745);
nor U12947 (N_12947,N_11442,N_11195);
or U12948 (N_12948,N_11173,N_11020);
nand U12949 (N_12949,N_11678,N_11707);
xnor U12950 (N_12950,N_11984,N_11630);
xnor U12951 (N_12951,N_11375,N_11431);
nor U12952 (N_12952,N_11635,N_11563);
or U12953 (N_12953,N_11780,N_11419);
xor U12954 (N_12954,N_11049,N_11492);
or U12955 (N_12955,N_11600,N_11155);
nor U12956 (N_12956,N_11101,N_11719);
xor U12957 (N_12957,N_11897,N_11516);
xnor U12958 (N_12958,N_11118,N_11099);
nand U12959 (N_12959,N_11245,N_11143);
nand U12960 (N_12960,N_11064,N_11947);
and U12961 (N_12961,N_11499,N_11581);
nor U12962 (N_12962,N_11635,N_11480);
or U12963 (N_12963,N_11634,N_11240);
or U12964 (N_12964,N_11740,N_11336);
xnor U12965 (N_12965,N_11597,N_11136);
or U12966 (N_12966,N_11197,N_11300);
and U12967 (N_12967,N_11267,N_11997);
xnor U12968 (N_12968,N_11527,N_11299);
or U12969 (N_12969,N_11062,N_11935);
nand U12970 (N_12970,N_11035,N_11651);
nand U12971 (N_12971,N_11775,N_11243);
and U12972 (N_12972,N_11016,N_11422);
xor U12973 (N_12973,N_11986,N_11726);
nor U12974 (N_12974,N_11312,N_11670);
nor U12975 (N_12975,N_11422,N_11407);
xnor U12976 (N_12976,N_11647,N_11577);
nand U12977 (N_12977,N_11057,N_11191);
nor U12978 (N_12978,N_11297,N_11254);
nor U12979 (N_12979,N_11914,N_11986);
xnor U12980 (N_12980,N_11853,N_11813);
nand U12981 (N_12981,N_11136,N_11609);
xnor U12982 (N_12982,N_11935,N_11394);
or U12983 (N_12983,N_11476,N_11929);
xor U12984 (N_12984,N_11919,N_11860);
nor U12985 (N_12985,N_11624,N_11033);
and U12986 (N_12986,N_11404,N_11748);
nand U12987 (N_12987,N_11426,N_11905);
xor U12988 (N_12988,N_11175,N_11633);
or U12989 (N_12989,N_11745,N_11969);
nand U12990 (N_12990,N_11732,N_11771);
nor U12991 (N_12991,N_11437,N_11531);
nor U12992 (N_12992,N_11191,N_11246);
xnor U12993 (N_12993,N_11466,N_11574);
xor U12994 (N_12994,N_11942,N_11459);
nand U12995 (N_12995,N_11010,N_11587);
or U12996 (N_12996,N_11815,N_11428);
nand U12997 (N_12997,N_11310,N_11745);
nand U12998 (N_12998,N_11056,N_11543);
nand U12999 (N_12999,N_11883,N_11937);
xor U13000 (N_13000,N_12838,N_12313);
or U13001 (N_13001,N_12680,N_12956);
and U13002 (N_13002,N_12473,N_12162);
or U13003 (N_13003,N_12489,N_12028);
nand U13004 (N_13004,N_12662,N_12106);
nand U13005 (N_13005,N_12309,N_12136);
xnor U13006 (N_13006,N_12395,N_12556);
and U13007 (N_13007,N_12352,N_12580);
or U13008 (N_13008,N_12042,N_12446);
xor U13009 (N_13009,N_12943,N_12876);
and U13010 (N_13010,N_12514,N_12099);
and U13011 (N_13011,N_12942,N_12161);
and U13012 (N_13012,N_12860,N_12209);
and U13013 (N_13013,N_12965,N_12359);
and U13014 (N_13014,N_12432,N_12635);
xnor U13015 (N_13015,N_12597,N_12755);
or U13016 (N_13016,N_12436,N_12717);
and U13017 (N_13017,N_12888,N_12706);
or U13018 (N_13018,N_12955,N_12534);
xor U13019 (N_13019,N_12132,N_12759);
nor U13020 (N_13020,N_12340,N_12734);
nand U13021 (N_13021,N_12894,N_12302);
nand U13022 (N_13022,N_12025,N_12324);
nand U13023 (N_13023,N_12661,N_12409);
nand U13024 (N_13024,N_12601,N_12345);
nor U13025 (N_13025,N_12204,N_12291);
and U13026 (N_13026,N_12554,N_12587);
xor U13027 (N_13027,N_12805,N_12711);
and U13028 (N_13028,N_12913,N_12286);
xnor U13029 (N_13029,N_12865,N_12967);
xor U13030 (N_13030,N_12539,N_12163);
nor U13031 (N_13031,N_12763,N_12142);
and U13032 (N_13032,N_12837,N_12337);
nand U13033 (N_13033,N_12841,N_12590);
or U13034 (N_13034,N_12069,N_12344);
nand U13035 (N_13035,N_12836,N_12783);
and U13036 (N_13036,N_12816,N_12460);
xor U13037 (N_13037,N_12517,N_12884);
and U13038 (N_13038,N_12715,N_12953);
or U13039 (N_13039,N_12819,N_12159);
xor U13040 (N_13040,N_12511,N_12929);
nand U13041 (N_13041,N_12623,N_12001);
and U13042 (N_13042,N_12368,N_12297);
or U13043 (N_13043,N_12505,N_12125);
or U13044 (N_13044,N_12215,N_12533);
xnor U13045 (N_13045,N_12626,N_12552);
nand U13046 (N_13046,N_12806,N_12279);
and U13047 (N_13047,N_12650,N_12979);
xnor U13048 (N_13048,N_12791,N_12969);
and U13049 (N_13049,N_12718,N_12926);
or U13050 (N_13050,N_12604,N_12524);
or U13051 (N_13051,N_12859,N_12295);
or U13052 (N_13052,N_12660,N_12752);
nand U13053 (N_13053,N_12912,N_12919);
nand U13054 (N_13054,N_12729,N_12245);
nor U13055 (N_13055,N_12433,N_12656);
nand U13056 (N_13056,N_12241,N_12257);
nand U13057 (N_13057,N_12108,N_12972);
xor U13058 (N_13058,N_12723,N_12267);
or U13059 (N_13059,N_12992,N_12703);
xor U13060 (N_13060,N_12088,N_12905);
and U13061 (N_13061,N_12644,N_12205);
or U13062 (N_13062,N_12549,N_12252);
and U13063 (N_13063,N_12331,N_12914);
nor U13064 (N_13064,N_12663,N_12450);
nand U13065 (N_13065,N_12802,N_12726);
nor U13066 (N_13066,N_12173,N_12426);
and U13067 (N_13067,N_12684,N_12148);
xnor U13068 (N_13068,N_12011,N_12307);
nor U13069 (N_13069,N_12115,N_12579);
xnor U13070 (N_13070,N_12284,N_12606);
xor U13071 (N_13071,N_12881,N_12230);
nor U13072 (N_13072,N_12641,N_12037);
or U13073 (N_13073,N_12174,N_12855);
nor U13074 (N_13074,N_12476,N_12184);
and U13075 (N_13075,N_12510,N_12893);
and U13076 (N_13076,N_12506,N_12405);
and U13077 (N_13077,N_12039,N_12364);
and U13078 (N_13078,N_12081,N_12885);
or U13079 (N_13079,N_12922,N_12586);
nor U13080 (N_13080,N_12664,N_12281);
or U13081 (N_13081,N_12092,N_12361);
xor U13082 (N_13082,N_12048,N_12997);
and U13083 (N_13083,N_12458,N_12652);
nor U13084 (N_13084,N_12647,N_12558);
nor U13085 (N_13085,N_12852,N_12135);
or U13086 (N_13086,N_12987,N_12072);
nand U13087 (N_13087,N_12126,N_12379);
nand U13088 (N_13088,N_12722,N_12129);
or U13089 (N_13089,N_12444,N_12197);
and U13090 (N_13090,N_12397,N_12832);
or U13091 (N_13091,N_12076,N_12090);
or U13092 (N_13092,N_12293,N_12124);
nor U13093 (N_13093,N_12323,N_12014);
xnor U13094 (N_13094,N_12634,N_12594);
or U13095 (N_13095,N_12431,N_12240);
nand U13096 (N_13096,N_12183,N_12870);
nor U13097 (N_13097,N_12848,N_12598);
or U13098 (N_13098,N_12311,N_12733);
nor U13099 (N_13099,N_12954,N_12145);
nor U13100 (N_13100,N_12053,N_12698);
nand U13101 (N_13101,N_12082,N_12328);
nand U13102 (N_13102,N_12730,N_12677);
or U13103 (N_13103,N_12268,N_12502);
or U13104 (N_13104,N_12471,N_12178);
nor U13105 (N_13105,N_12044,N_12996);
and U13106 (N_13106,N_12957,N_12440);
or U13107 (N_13107,N_12827,N_12310);
nor U13108 (N_13108,N_12550,N_12646);
or U13109 (N_13109,N_12185,N_12574);
or U13110 (N_13110,N_12788,N_12710);
nor U13111 (N_13111,N_12632,N_12420);
nand U13112 (N_13112,N_12330,N_12067);
and U13113 (N_13113,N_12638,N_12765);
nand U13114 (N_13114,N_12847,N_12786);
or U13115 (N_13115,N_12224,N_12864);
nand U13116 (N_13116,N_12984,N_12160);
xor U13117 (N_13117,N_12867,N_12525);
nand U13118 (N_13118,N_12437,N_12519);
or U13119 (N_13119,N_12256,N_12430);
or U13120 (N_13120,N_12298,N_12674);
or U13121 (N_13121,N_12176,N_12180);
nand U13122 (N_13122,N_12269,N_12889);
xnor U13123 (N_13123,N_12949,N_12461);
nor U13124 (N_13124,N_12451,N_12386);
or U13125 (N_13125,N_12610,N_12583);
or U13126 (N_13126,N_12393,N_12109);
and U13127 (N_13127,N_12441,N_12410);
or U13128 (N_13128,N_12625,N_12317);
nor U13129 (N_13129,N_12536,N_12991);
xor U13130 (N_13130,N_12459,N_12333);
nand U13131 (N_13131,N_12339,N_12486);
xor U13132 (N_13132,N_12631,N_12654);
nand U13133 (N_13133,N_12777,N_12123);
or U13134 (N_13134,N_12024,N_12611);
and U13135 (N_13135,N_12974,N_12879);
xor U13136 (N_13136,N_12246,N_12447);
nor U13137 (N_13137,N_12003,N_12941);
and U13138 (N_13138,N_12512,N_12551);
xnor U13139 (N_13139,N_12719,N_12113);
xnor U13140 (N_13140,N_12043,N_12636);
and U13141 (N_13141,N_12541,N_12857);
and U13142 (N_13142,N_12897,N_12272);
nand U13143 (N_13143,N_12232,N_12341);
nor U13144 (N_13144,N_12607,N_12559);
or U13145 (N_13145,N_12998,N_12052);
xnor U13146 (N_13146,N_12553,N_12872);
nand U13147 (N_13147,N_12303,N_12970);
and U13148 (N_13148,N_12620,N_12384);
or U13149 (N_13149,N_12807,N_12016);
xnor U13150 (N_13150,N_12946,N_12417);
nand U13151 (N_13151,N_12983,N_12036);
and U13152 (N_13152,N_12973,N_12285);
nand U13153 (N_13153,N_12371,N_12761);
and U13154 (N_13154,N_12538,N_12801);
nand U13155 (N_13155,N_12002,N_12675);
nor U13156 (N_13156,N_12147,N_12038);
and U13157 (N_13157,N_12040,N_12628);
nand U13158 (N_13158,N_12760,N_12762);
and U13159 (N_13159,N_12784,N_12637);
or U13160 (N_13160,N_12004,N_12182);
nor U13161 (N_13161,N_12753,N_12924);
nor U13162 (N_13162,N_12271,N_12501);
nand U13163 (N_13163,N_12006,N_12110);
nand U13164 (N_13164,N_12214,N_12187);
and U13165 (N_13165,N_12787,N_12665);
xor U13166 (N_13166,N_12336,N_12380);
nor U13167 (N_13167,N_12172,N_12809);
xnor U13168 (N_13168,N_12732,N_12366);
nor U13169 (N_13169,N_12047,N_12105);
nor U13170 (N_13170,N_12362,N_12290);
nor U13171 (N_13171,N_12265,N_12374);
nor U13172 (N_13172,N_12227,N_12455);
nand U13173 (N_13173,N_12804,N_12485);
and U13174 (N_13174,N_12299,N_12645);
nor U13175 (N_13175,N_12225,N_12866);
and U13176 (N_13176,N_12496,N_12790);
nor U13177 (N_13177,N_12414,N_12153);
nor U13178 (N_13178,N_12022,N_12627);
or U13179 (N_13179,N_12679,N_12454);
nand U13180 (N_13180,N_12195,N_12289);
nor U13181 (N_13181,N_12350,N_12475);
nand U13182 (N_13182,N_12915,N_12509);
or U13183 (N_13183,N_12692,N_12716);
or U13184 (N_13184,N_12695,N_12971);
and U13185 (N_13185,N_12070,N_12399);
and U13186 (N_13186,N_12582,N_12988);
xnor U13187 (N_13187,N_12931,N_12743);
xnor U13188 (N_13188,N_12216,N_12798);
and U13189 (N_13189,N_12179,N_12000);
xor U13190 (N_13190,N_12482,N_12168);
or U13191 (N_13191,N_12812,N_12990);
xor U13192 (N_13192,N_12057,N_12027);
nand U13193 (N_13193,N_12061,N_12633);
and U13194 (N_13194,N_12463,N_12466);
nor U13195 (N_13195,N_12744,N_12089);
nor U13196 (N_13196,N_12354,N_12348);
xor U13197 (N_13197,N_12064,N_12966);
nor U13198 (N_13198,N_12562,N_12300);
and U13199 (N_13199,N_12236,N_12308);
nor U13200 (N_13200,N_12681,N_12210);
or U13201 (N_13201,N_12856,N_12874);
nor U13202 (N_13202,N_12797,N_12900);
and U13203 (N_13203,N_12746,N_12372);
nor U13204 (N_13204,N_12342,N_12375);
or U13205 (N_13205,N_12032,N_12814);
or U13206 (N_13206,N_12098,N_12369);
nand U13207 (N_13207,N_12065,N_12139);
or U13208 (N_13208,N_12520,N_12657);
nand U13209 (N_13209,N_12276,N_12731);
nor U13210 (N_13210,N_12425,N_12535);
nand U13211 (N_13211,N_12878,N_12821);
nand U13212 (N_13212,N_12465,N_12909);
and U13213 (N_13213,N_12618,N_12748);
and U13214 (N_13214,N_12521,N_12621);
xnor U13215 (N_13215,N_12690,N_12095);
and U13216 (N_13216,N_12813,N_12356);
and U13217 (N_13217,N_12470,N_12497);
nor U13218 (N_13218,N_12253,N_12051);
or U13219 (N_13219,N_12989,N_12803);
or U13220 (N_13220,N_12778,N_12021);
nor U13221 (N_13221,N_12795,N_12563);
nor U13222 (N_13222,N_12068,N_12704);
and U13223 (N_13223,N_12221,N_12434);
nand U13224 (N_13224,N_12403,N_12448);
xnor U13225 (N_13225,N_12149,N_12902);
xor U13226 (N_13226,N_12443,N_12208);
nor U13227 (N_13227,N_12713,N_12818);
nand U13228 (N_13228,N_12009,N_12054);
nor U13229 (N_13229,N_12916,N_12944);
nand U13230 (N_13230,N_12117,N_12060);
nor U13231 (N_13231,N_12388,N_12899);
xnor U13232 (N_13232,N_12775,N_12391);
or U13233 (N_13233,N_12191,N_12781);
or U13234 (N_13234,N_12581,N_12747);
or U13235 (N_13235,N_12238,N_12008);
nand U13236 (N_13236,N_12602,N_12111);
or U13237 (N_13237,N_12277,N_12616);
xnor U13238 (N_13238,N_12565,N_12377);
nand U13239 (N_13239,N_12322,N_12599);
and U13240 (N_13240,N_12767,N_12937);
and U13241 (N_13241,N_12050,N_12705);
xnor U13242 (N_13242,N_12234,N_12213);
nor U13243 (N_13243,N_12764,N_12921);
xnor U13244 (N_13244,N_12758,N_12958);
nor U13245 (N_13245,N_12190,N_12326);
nor U13246 (N_13246,N_12408,N_12873);
nor U13247 (N_13247,N_12720,N_12868);
nand U13248 (N_13248,N_12688,N_12035);
or U13249 (N_13249,N_12305,N_12155);
and U13250 (N_13250,N_12087,N_12239);
nand U13251 (N_13251,N_12614,N_12167);
or U13252 (N_13252,N_12146,N_12030);
nor U13253 (N_13253,N_12096,N_12651);
or U13254 (N_13254,N_12591,N_12248);
or U13255 (N_13255,N_12062,N_12605);
or U13256 (N_13256,N_12985,N_12367);
nand U13257 (N_13257,N_12423,N_12171);
nor U13258 (N_13258,N_12642,N_12121);
or U13259 (N_13259,N_12382,N_12355);
xnor U13260 (N_13260,N_12796,N_12325);
and U13261 (N_13261,N_12522,N_12863);
xor U13262 (N_13262,N_12250,N_12218);
nand U13263 (N_13263,N_12396,N_12166);
nand U13264 (N_13264,N_12708,N_12570);
nand U13265 (N_13265,N_12964,N_12976);
xor U13266 (N_13266,N_12370,N_12673);
xor U13267 (N_13267,N_12118,N_12274);
nand U13268 (N_13268,N_12363,N_12059);
xnor U13269 (N_13269,N_12378,N_12910);
nand U13270 (N_13270,N_12243,N_12999);
xnor U13271 (N_13271,N_12055,N_12073);
or U13272 (N_13272,N_12066,N_12346);
nand U13273 (N_13273,N_12537,N_12170);
nand U13274 (N_13274,N_12242,N_12456);
and U13275 (N_13275,N_12353,N_12488);
xnor U13276 (N_13276,N_12138,N_12484);
nor U13277 (N_13277,N_12516,N_12398);
nand U13278 (N_13278,N_12228,N_12200);
nor U13279 (N_13279,N_12347,N_12231);
xor U13280 (N_13280,N_12544,N_12993);
and U13281 (N_13281,N_12419,N_12084);
xnor U13282 (N_13282,N_12843,N_12564);
and U13283 (N_13283,N_12810,N_12572);
or U13284 (N_13284,N_12828,N_12203);
xnor U13285 (N_13285,N_12315,N_12503);
xor U13286 (N_13286,N_12593,N_12156);
or U13287 (N_13287,N_12130,N_12280);
nand U13288 (N_13288,N_12817,N_12151);
or U13289 (N_13289,N_12406,N_12928);
nor U13290 (N_13290,N_12413,N_12714);
and U13291 (N_13291,N_12102,N_12515);
and U13292 (N_13292,N_12120,N_12849);
or U13293 (N_13293,N_12617,N_12217);
xor U13294 (N_13294,N_12206,N_12329);
and U13295 (N_13295,N_12199,N_12114);
or U13296 (N_13296,N_12986,N_12415);
and U13297 (N_13297,N_12869,N_12877);
and U13298 (N_13298,N_12493,N_12696);
xor U13299 (N_13299,N_12494,N_12595);
nor U13300 (N_13300,N_12685,N_12567);
nor U13301 (N_13301,N_12980,N_12947);
nor U13302 (N_13302,N_12530,N_12982);
nor U13303 (N_13303,N_12622,N_12404);
xor U13304 (N_13304,N_12697,N_12890);
nor U13305 (N_13305,N_12882,N_12930);
and U13306 (N_13306,N_12938,N_12569);
or U13307 (N_13307,N_12830,N_12133);
xnor U13308 (N_13308,N_12196,N_12422);
or U13309 (N_13309,N_12691,N_12917);
nand U13310 (N_13310,N_12193,N_12799);
nor U13311 (N_13311,N_12895,N_12411);
nor U13312 (N_13312,N_12766,N_12960);
xnor U13313 (N_13313,N_12649,N_12903);
or U13314 (N_13314,N_12825,N_12015);
xor U13315 (N_13315,N_12693,N_12518);
or U13316 (N_13316,N_12737,N_12771);
nand U13317 (N_13317,N_12792,N_12435);
xnor U13318 (N_13318,N_12029,N_12756);
nor U13319 (N_13319,N_12896,N_12270);
or U13320 (N_13320,N_12198,N_12659);
or U13321 (N_13321,N_12507,N_12296);
nand U13322 (N_13322,N_12385,N_12278);
nor U13323 (N_13323,N_12939,N_12316);
nand U13324 (N_13324,N_12392,N_12287);
nand U13325 (N_13325,N_12351,N_12546);
nand U13326 (N_13326,N_12721,N_12480);
nand U13327 (N_13327,N_12951,N_12612);
and U13328 (N_13328,N_12749,N_12835);
or U13329 (N_13329,N_12034,N_12738);
nand U13330 (N_13330,N_12119,N_12429);
nand U13331 (N_13331,N_12334,N_12648);
and U13332 (N_13332,N_12007,N_12264);
or U13333 (N_13333,N_12682,N_12923);
xor U13334 (N_13334,N_12131,N_12258);
xnor U13335 (N_13335,N_12181,N_12741);
or U13336 (N_13336,N_12150,N_12304);
nand U13337 (N_13337,N_12154,N_12306);
nor U13338 (N_13338,N_12247,N_12251);
xor U13339 (N_13339,N_12822,N_12100);
nand U13340 (N_13340,N_12780,N_12031);
and U13341 (N_13341,N_12086,N_12948);
and U13342 (N_13342,N_12143,N_12212);
and U13343 (N_13343,N_12026,N_12573);
nand U13344 (N_13344,N_12672,N_12049);
xnor U13345 (N_13345,N_12523,N_12376);
or U13346 (N_13346,N_12400,N_12940);
xnor U13347 (N_13347,N_12157,N_12144);
and U13348 (N_13348,N_12768,N_12492);
nor U13349 (N_13349,N_12887,N_12933);
and U13350 (N_13350,N_12815,N_12596);
or U13351 (N_13351,N_12401,N_12824);
nor U13352 (N_13352,N_12891,N_12192);
xnor U13353 (N_13353,N_12686,N_12603);
and U13354 (N_13354,N_12235,N_12335);
or U13355 (N_13355,N_12700,N_12770);
nand U13356 (N_13356,N_12935,N_12439);
xor U13357 (N_13357,N_12745,N_12226);
xor U13358 (N_13358,N_12557,N_12629);
and U13359 (N_13359,N_12013,N_12906);
nor U13360 (N_13360,N_12262,N_12023);
nor U13361 (N_13361,N_12462,N_12707);
nand U13362 (N_13362,N_12079,N_12018);
and U13363 (N_13363,N_12107,N_12811);
or U13364 (N_13364,N_12576,N_12671);
or U13365 (N_13365,N_12464,N_12349);
xnor U13366 (N_13366,N_12474,N_12981);
or U13367 (N_13367,N_12689,N_12080);
xnor U13368 (N_13368,N_12880,N_12794);
nor U13369 (N_13369,N_12041,N_12504);
xnor U13370 (N_13370,N_12078,N_12094);
nor U13371 (N_13371,N_12845,N_12585);
and U13372 (N_13372,N_12736,N_12075);
nor U13373 (N_13373,N_12724,N_12609);
xor U13374 (N_13374,N_12207,N_12438);
or U13375 (N_13375,N_12727,N_12140);
and U13376 (N_13376,N_12116,N_12010);
nor U13377 (N_13377,N_12085,N_12853);
nor U13378 (N_13378,N_12449,N_12739);
and U13379 (N_13379,N_12481,N_12694);
or U13380 (N_13380,N_12548,N_12428);
nor U13381 (N_13381,N_12653,N_12421);
and U13382 (N_13382,N_12568,N_12904);
nand U13383 (N_13383,N_12312,N_12012);
and U13384 (N_13384,N_12365,N_12769);
nand U13385 (N_13385,N_12709,N_12319);
or U13386 (N_13386,N_12407,N_12712);
nand U13387 (N_13387,N_12292,N_12020);
nand U13388 (N_13388,N_12219,N_12959);
or U13389 (N_13389,N_12058,N_12263);
or U13390 (N_13390,N_12725,N_12789);
and U13391 (N_13391,N_12445,N_12532);
and U13392 (N_13392,N_12774,N_12630);
nor U13393 (N_13393,N_12266,N_12547);
xor U13394 (N_13394,N_12619,N_12776);
nor U13395 (N_13395,N_12188,N_12963);
or U13396 (N_13396,N_12063,N_12255);
nor U13397 (N_13397,N_12495,N_12531);
or U13398 (N_13398,N_12643,N_12261);
and U13399 (N_13399,N_12165,N_12543);
nand U13400 (N_13400,N_12091,N_12994);
nand U13401 (N_13401,N_12945,N_12927);
and U13402 (N_13402,N_12871,N_12418);
xor U13403 (N_13403,N_12046,N_12540);
nand U13404 (N_13404,N_12137,N_12840);
or U13405 (N_13405,N_12901,N_12045);
nor U13406 (N_13406,N_12338,N_12702);
xnor U13407 (N_13407,N_12735,N_12469);
nor U13408 (N_13408,N_12995,N_12453);
nor U13409 (N_13409,N_12477,N_12678);
nor U13410 (N_13410,N_12152,N_12952);
xor U13411 (N_13411,N_12757,N_12829);
or U13412 (N_13412,N_12483,N_12390);
xor U13413 (N_13413,N_12831,N_12975);
nor U13414 (N_13414,N_12920,N_12833);
and U13415 (N_13415,N_12584,N_12658);
nor U13416 (N_13416,N_12808,N_12850);
xnor U13417 (N_13417,N_12201,N_12093);
or U13418 (N_13418,N_12854,N_12083);
xnor U13419 (N_13419,N_12452,N_12128);
nor U13420 (N_13420,N_12468,N_12779);
nand U13421 (N_13421,N_12592,N_12750);
or U13422 (N_13422,N_12555,N_12898);
nor U13423 (N_13423,N_12186,N_12472);
nand U13424 (N_13424,N_12402,N_12577);
nor U13425 (N_13425,N_12103,N_12498);
or U13426 (N_13426,N_12782,N_12314);
xnor U13427 (N_13427,N_12751,N_12259);
and U13428 (N_13428,N_12785,N_12244);
xnor U13429 (N_13429,N_12608,N_12886);
or U13430 (N_13430,N_12529,N_12071);
and U13431 (N_13431,N_12019,N_12358);
xor U13432 (N_13432,N_12233,N_12260);
and U13433 (N_13433,N_12332,N_12962);
nand U13434 (N_13434,N_12427,N_12578);
or U13435 (N_13435,N_12793,N_12127);
nor U13436 (N_13436,N_12412,N_12177);
nor U13437 (N_13437,N_12613,N_12683);
or U13438 (N_13438,N_12624,N_12542);
nand U13439 (N_13439,N_12842,N_12122);
nand U13440 (N_13440,N_12666,N_12911);
xnor U13441 (N_13441,N_12918,N_12479);
nor U13442 (N_13442,N_12211,N_12588);
or U13443 (N_13443,N_12851,N_12104);
or U13444 (N_13444,N_12288,N_12571);
nor U13445 (N_13445,N_12134,N_12861);
and U13446 (N_13446,N_12978,N_12932);
or U13447 (N_13447,N_12249,N_12934);
nor U13448 (N_13448,N_12977,N_12321);
and U13449 (N_13449,N_12640,N_12820);
xnor U13450 (N_13450,N_12194,N_12318);
and U13451 (N_13451,N_12017,N_12936);
xor U13452 (N_13452,N_12875,N_12033);
xnor U13453 (N_13453,N_12858,N_12357);
xor U13454 (N_13454,N_12005,N_12834);
and U13455 (N_13455,N_12499,N_12600);
nand U13456 (N_13456,N_12175,N_12846);
xor U13457 (N_13457,N_12491,N_12327);
and U13458 (N_13458,N_12381,N_12699);
or U13459 (N_13459,N_12528,N_12908);
or U13460 (N_13460,N_12467,N_12826);
xnor U13461 (N_13461,N_12639,N_12282);
nand U13462 (N_13462,N_12701,N_12373);
nand U13463 (N_13463,N_12112,N_12077);
or U13464 (N_13464,N_12478,N_12237);
or U13465 (N_13465,N_12589,N_12294);
and U13466 (N_13466,N_12545,N_12961);
or U13467 (N_13467,N_12487,N_12925);
or U13468 (N_13468,N_12566,N_12387);
xnor U13469 (N_13469,N_12500,N_12669);
nor U13470 (N_13470,N_12457,N_12220);
xor U13471 (N_13471,N_12742,N_12101);
and U13472 (N_13472,N_12273,N_12074);
or U13473 (N_13473,N_12527,N_12907);
nor U13474 (N_13474,N_12275,N_12950);
nand U13475 (N_13475,N_12169,N_12773);
xnor U13476 (N_13476,N_12508,N_12823);
and U13477 (N_13477,N_12513,N_12687);
nor U13478 (N_13478,N_12561,N_12968);
nand U13479 (N_13479,N_12416,N_12254);
xnor U13480 (N_13480,N_12883,N_12839);
and U13481 (N_13481,N_12800,N_12158);
or U13482 (N_13482,N_12164,N_12383);
xnor U13483 (N_13483,N_12490,N_12320);
and U13484 (N_13484,N_12097,N_12360);
nand U13485 (N_13485,N_12283,N_12667);
nand U13486 (N_13486,N_12676,N_12754);
and U13487 (N_13487,N_12424,N_12301);
and U13488 (N_13488,N_12668,N_12394);
nor U13489 (N_13489,N_12442,N_12862);
xor U13490 (N_13490,N_12655,N_12389);
nor U13491 (N_13491,N_12056,N_12728);
and U13492 (N_13492,N_12526,N_12772);
nor U13493 (N_13493,N_12892,N_12575);
nor U13494 (N_13494,N_12615,N_12202);
xor U13495 (N_13495,N_12223,N_12670);
and U13496 (N_13496,N_12222,N_12189);
nand U13497 (N_13497,N_12229,N_12141);
or U13498 (N_13498,N_12343,N_12844);
or U13499 (N_13499,N_12740,N_12560);
and U13500 (N_13500,N_12267,N_12669);
nor U13501 (N_13501,N_12966,N_12220);
nand U13502 (N_13502,N_12714,N_12111);
nand U13503 (N_13503,N_12719,N_12471);
and U13504 (N_13504,N_12011,N_12309);
or U13505 (N_13505,N_12647,N_12347);
nand U13506 (N_13506,N_12610,N_12185);
xor U13507 (N_13507,N_12867,N_12627);
nor U13508 (N_13508,N_12869,N_12855);
xor U13509 (N_13509,N_12762,N_12225);
xor U13510 (N_13510,N_12290,N_12172);
xor U13511 (N_13511,N_12719,N_12586);
nand U13512 (N_13512,N_12622,N_12437);
and U13513 (N_13513,N_12483,N_12429);
and U13514 (N_13514,N_12095,N_12733);
nor U13515 (N_13515,N_12125,N_12458);
nand U13516 (N_13516,N_12967,N_12818);
nand U13517 (N_13517,N_12449,N_12464);
or U13518 (N_13518,N_12908,N_12060);
nor U13519 (N_13519,N_12180,N_12053);
xnor U13520 (N_13520,N_12988,N_12558);
nor U13521 (N_13521,N_12570,N_12817);
xor U13522 (N_13522,N_12108,N_12005);
nor U13523 (N_13523,N_12829,N_12800);
nand U13524 (N_13524,N_12352,N_12363);
nor U13525 (N_13525,N_12766,N_12709);
and U13526 (N_13526,N_12084,N_12120);
and U13527 (N_13527,N_12678,N_12046);
xor U13528 (N_13528,N_12289,N_12868);
xnor U13529 (N_13529,N_12863,N_12697);
nor U13530 (N_13530,N_12539,N_12896);
xor U13531 (N_13531,N_12109,N_12714);
nand U13532 (N_13532,N_12858,N_12894);
xor U13533 (N_13533,N_12661,N_12214);
xnor U13534 (N_13534,N_12716,N_12647);
or U13535 (N_13535,N_12788,N_12718);
nand U13536 (N_13536,N_12487,N_12974);
and U13537 (N_13537,N_12404,N_12874);
and U13538 (N_13538,N_12314,N_12535);
or U13539 (N_13539,N_12576,N_12364);
xor U13540 (N_13540,N_12309,N_12154);
xnor U13541 (N_13541,N_12085,N_12599);
nor U13542 (N_13542,N_12577,N_12935);
or U13543 (N_13543,N_12055,N_12008);
or U13544 (N_13544,N_12762,N_12179);
nand U13545 (N_13545,N_12146,N_12631);
or U13546 (N_13546,N_12884,N_12298);
or U13547 (N_13547,N_12292,N_12113);
xnor U13548 (N_13548,N_12893,N_12579);
or U13549 (N_13549,N_12869,N_12969);
or U13550 (N_13550,N_12691,N_12299);
and U13551 (N_13551,N_12519,N_12661);
nor U13552 (N_13552,N_12116,N_12072);
xor U13553 (N_13553,N_12283,N_12807);
nor U13554 (N_13554,N_12891,N_12921);
or U13555 (N_13555,N_12520,N_12481);
nand U13556 (N_13556,N_12487,N_12793);
nand U13557 (N_13557,N_12742,N_12091);
or U13558 (N_13558,N_12443,N_12628);
or U13559 (N_13559,N_12227,N_12148);
nand U13560 (N_13560,N_12756,N_12544);
or U13561 (N_13561,N_12506,N_12888);
and U13562 (N_13562,N_12884,N_12190);
nand U13563 (N_13563,N_12692,N_12931);
or U13564 (N_13564,N_12811,N_12466);
nand U13565 (N_13565,N_12966,N_12628);
nand U13566 (N_13566,N_12960,N_12923);
and U13567 (N_13567,N_12462,N_12926);
and U13568 (N_13568,N_12604,N_12059);
and U13569 (N_13569,N_12133,N_12931);
and U13570 (N_13570,N_12353,N_12573);
or U13571 (N_13571,N_12252,N_12954);
and U13572 (N_13572,N_12020,N_12249);
xor U13573 (N_13573,N_12333,N_12254);
nand U13574 (N_13574,N_12060,N_12925);
nand U13575 (N_13575,N_12652,N_12708);
and U13576 (N_13576,N_12819,N_12766);
and U13577 (N_13577,N_12250,N_12071);
nand U13578 (N_13578,N_12099,N_12019);
nor U13579 (N_13579,N_12235,N_12196);
xnor U13580 (N_13580,N_12443,N_12100);
nand U13581 (N_13581,N_12261,N_12677);
nor U13582 (N_13582,N_12949,N_12800);
nor U13583 (N_13583,N_12577,N_12722);
nor U13584 (N_13584,N_12299,N_12951);
nand U13585 (N_13585,N_12739,N_12238);
nor U13586 (N_13586,N_12645,N_12131);
nor U13587 (N_13587,N_12310,N_12449);
nor U13588 (N_13588,N_12627,N_12343);
or U13589 (N_13589,N_12706,N_12914);
xnor U13590 (N_13590,N_12258,N_12722);
and U13591 (N_13591,N_12442,N_12347);
nor U13592 (N_13592,N_12113,N_12224);
nand U13593 (N_13593,N_12124,N_12461);
xnor U13594 (N_13594,N_12405,N_12159);
or U13595 (N_13595,N_12652,N_12315);
nor U13596 (N_13596,N_12209,N_12065);
and U13597 (N_13597,N_12923,N_12461);
nand U13598 (N_13598,N_12545,N_12700);
or U13599 (N_13599,N_12324,N_12685);
nand U13600 (N_13600,N_12393,N_12512);
xor U13601 (N_13601,N_12112,N_12052);
or U13602 (N_13602,N_12979,N_12931);
and U13603 (N_13603,N_12154,N_12993);
or U13604 (N_13604,N_12568,N_12925);
or U13605 (N_13605,N_12722,N_12560);
xor U13606 (N_13606,N_12123,N_12970);
nand U13607 (N_13607,N_12329,N_12350);
nor U13608 (N_13608,N_12369,N_12074);
or U13609 (N_13609,N_12885,N_12048);
or U13610 (N_13610,N_12544,N_12004);
and U13611 (N_13611,N_12049,N_12613);
nand U13612 (N_13612,N_12032,N_12688);
and U13613 (N_13613,N_12526,N_12667);
nand U13614 (N_13614,N_12136,N_12844);
xor U13615 (N_13615,N_12689,N_12136);
and U13616 (N_13616,N_12210,N_12844);
nand U13617 (N_13617,N_12737,N_12556);
and U13618 (N_13618,N_12389,N_12253);
or U13619 (N_13619,N_12193,N_12631);
and U13620 (N_13620,N_12527,N_12072);
nand U13621 (N_13621,N_12184,N_12710);
xor U13622 (N_13622,N_12077,N_12828);
xnor U13623 (N_13623,N_12173,N_12961);
or U13624 (N_13624,N_12671,N_12795);
and U13625 (N_13625,N_12164,N_12444);
xnor U13626 (N_13626,N_12514,N_12210);
and U13627 (N_13627,N_12971,N_12743);
xor U13628 (N_13628,N_12857,N_12932);
nor U13629 (N_13629,N_12325,N_12419);
and U13630 (N_13630,N_12282,N_12321);
nand U13631 (N_13631,N_12548,N_12120);
xor U13632 (N_13632,N_12160,N_12140);
xor U13633 (N_13633,N_12338,N_12019);
xor U13634 (N_13634,N_12843,N_12734);
and U13635 (N_13635,N_12362,N_12504);
and U13636 (N_13636,N_12964,N_12196);
xnor U13637 (N_13637,N_12783,N_12855);
xnor U13638 (N_13638,N_12956,N_12678);
xor U13639 (N_13639,N_12982,N_12448);
xnor U13640 (N_13640,N_12281,N_12853);
and U13641 (N_13641,N_12683,N_12903);
nand U13642 (N_13642,N_12209,N_12898);
or U13643 (N_13643,N_12843,N_12481);
and U13644 (N_13644,N_12567,N_12467);
or U13645 (N_13645,N_12617,N_12976);
nor U13646 (N_13646,N_12717,N_12887);
and U13647 (N_13647,N_12480,N_12145);
nor U13648 (N_13648,N_12979,N_12633);
and U13649 (N_13649,N_12677,N_12869);
or U13650 (N_13650,N_12989,N_12168);
or U13651 (N_13651,N_12813,N_12602);
or U13652 (N_13652,N_12103,N_12475);
or U13653 (N_13653,N_12174,N_12420);
and U13654 (N_13654,N_12108,N_12270);
nand U13655 (N_13655,N_12622,N_12827);
xnor U13656 (N_13656,N_12648,N_12564);
and U13657 (N_13657,N_12508,N_12602);
nand U13658 (N_13658,N_12761,N_12981);
xor U13659 (N_13659,N_12501,N_12403);
xor U13660 (N_13660,N_12133,N_12340);
or U13661 (N_13661,N_12751,N_12442);
xnor U13662 (N_13662,N_12618,N_12932);
and U13663 (N_13663,N_12827,N_12138);
nand U13664 (N_13664,N_12517,N_12271);
nor U13665 (N_13665,N_12214,N_12096);
nor U13666 (N_13666,N_12495,N_12168);
and U13667 (N_13667,N_12570,N_12595);
nand U13668 (N_13668,N_12328,N_12303);
xor U13669 (N_13669,N_12246,N_12036);
and U13670 (N_13670,N_12894,N_12363);
xor U13671 (N_13671,N_12197,N_12817);
and U13672 (N_13672,N_12928,N_12502);
or U13673 (N_13673,N_12366,N_12023);
nand U13674 (N_13674,N_12552,N_12229);
nor U13675 (N_13675,N_12013,N_12399);
nor U13676 (N_13676,N_12711,N_12513);
and U13677 (N_13677,N_12830,N_12998);
nand U13678 (N_13678,N_12171,N_12737);
xor U13679 (N_13679,N_12430,N_12425);
and U13680 (N_13680,N_12725,N_12578);
xor U13681 (N_13681,N_12270,N_12484);
xor U13682 (N_13682,N_12656,N_12636);
nand U13683 (N_13683,N_12250,N_12233);
xnor U13684 (N_13684,N_12543,N_12170);
or U13685 (N_13685,N_12997,N_12469);
nand U13686 (N_13686,N_12947,N_12163);
xnor U13687 (N_13687,N_12137,N_12594);
and U13688 (N_13688,N_12110,N_12232);
or U13689 (N_13689,N_12990,N_12283);
nand U13690 (N_13690,N_12122,N_12423);
nand U13691 (N_13691,N_12867,N_12283);
and U13692 (N_13692,N_12720,N_12903);
nand U13693 (N_13693,N_12711,N_12933);
and U13694 (N_13694,N_12666,N_12266);
nor U13695 (N_13695,N_12432,N_12012);
and U13696 (N_13696,N_12131,N_12610);
nand U13697 (N_13697,N_12238,N_12231);
xor U13698 (N_13698,N_12624,N_12342);
nor U13699 (N_13699,N_12550,N_12803);
nor U13700 (N_13700,N_12423,N_12747);
and U13701 (N_13701,N_12323,N_12888);
or U13702 (N_13702,N_12187,N_12713);
xor U13703 (N_13703,N_12647,N_12914);
nor U13704 (N_13704,N_12067,N_12847);
or U13705 (N_13705,N_12243,N_12199);
nor U13706 (N_13706,N_12817,N_12227);
and U13707 (N_13707,N_12001,N_12104);
nand U13708 (N_13708,N_12846,N_12592);
nor U13709 (N_13709,N_12683,N_12359);
and U13710 (N_13710,N_12452,N_12094);
or U13711 (N_13711,N_12658,N_12285);
nand U13712 (N_13712,N_12932,N_12323);
xor U13713 (N_13713,N_12296,N_12242);
xnor U13714 (N_13714,N_12190,N_12990);
and U13715 (N_13715,N_12340,N_12348);
or U13716 (N_13716,N_12136,N_12462);
nor U13717 (N_13717,N_12978,N_12625);
and U13718 (N_13718,N_12534,N_12840);
and U13719 (N_13719,N_12691,N_12159);
nor U13720 (N_13720,N_12194,N_12163);
xnor U13721 (N_13721,N_12074,N_12903);
nor U13722 (N_13722,N_12032,N_12666);
and U13723 (N_13723,N_12666,N_12596);
and U13724 (N_13724,N_12326,N_12105);
xor U13725 (N_13725,N_12990,N_12669);
or U13726 (N_13726,N_12570,N_12805);
nand U13727 (N_13727,N_12902,N_12658);
and U13728 (N_13728,N_12685,N_12319);
and U13729 (N_13729,N_12593,N_12438);
xor U13730 (N_13730,N_12447,N_12666);
nand U13731 (N_13731,N_12310,N_12171);
nand U13732 (N_13732,N_12383,N_12196);
xor U13733 (N_13733,N_12544,N_12743);
and U13734 (N_13734,N_12546,N_12459);
or U13735 (N_13735,N_12402,N_12890);
nor U13736 (N_13736,N_12312,N_12228);
and U13737 (N_13737,N_12614,N_12152);
xor U13738 (N_13738,N_12305,N_12663);
nor U13739 (N_13739,N_12518,N_12555);
xor U13740 (N_13740,N_12367,N_12080);
and U13741 (N_13741,N_12650,N_12106);
and U13742 (N_13742,N_12461,N_12920);
xor U13743 (N_13743,N_12609,N_12813);
xor U13744 (N_13744,N_12698,N_12302);
xnor U13745 (N_13745,N_12903,N_12209);
or U13746 (N_13746,N_12886,N_12065);
nand U13747 (N_13747,N_12895,N_12494);
nor U13748 (N_13748,N_12133,N_12012);
xor U13749 (N_13749,N_12160,N_12011);
and U13750 (N_13750,N_12638,N_12730);
nand U13751 (N_13751,N_12331,N_12159);
and U13752 (N_13752,N_12216,N_12190);
xnor U13753 (N_13753,N_12269,N_12102);
nand U13754 (N_13754,N_12371,N_12835);
nand U13755 (N_13755,N_12924,N_12242);
nor U13756 (N_13756,N_12505,N_12353);
nand U13757 (N_13757,N_12043,N_12980);
nand U13758 (N_13758,N_12943,N_12364);
xnor U13759 (N_13759,N_12715,N_12085);
and U13760 (N_13760,N_12151,N_12016);
nand U13761 (N_13761,N_12202,N_12680);
nand U13762 (N_13762,N_12927,N_12628);
xor U13763 (N_13763,N_12142,N_12692);
and U13764 (N_13764,N_12998,N_12869);
nand U13765 (N_13765,N_12676,N_12686);
xor U13766 (N_13766,N_12534,N_12078);
and U13767 (N_13767,N_12637,N_12336);
nor U13768 (N_13768,N_12270,N_12124);
and U13769 (N_13769,N_12189,N_12460);
nor U13770 (N_13770,N_12787,N_12713);
nand U13771 (N_13771,N_12631,N_12928);
nand U13772 (N_13772,N_12500,N_12827);
or U13773 (N_13773,N_12593,N_12925);
and U13774 (N_13774,N_12046,N_12376);
nand U13775 (N_13775,N_12658,N_12605);
or U13776 (N_13776,N_12855,N_12143);
nand U13777 (N_13777,N_12701,N_12430);
or U13778 (N_13778,N_12711,N_12152);
nand U13779 (N_13779,N_12391,N_12941);
and U13780 (N_13780,N_12398,N_12323);
or U13781 (N_13781,N_12775,N_12257);
and U13782 (N_13782,N_12142,N_12418);
nor U13783 (N_13783,N_12956,N_12110);
xor U13784 (N_13784,N_12139,N_12792);
xnor U13785 (N_13785,N_12667,N_12163);
or U13786 (N_13786,N_12456,N_12897);
or U13787 (N_13787,N_12559,N_12203);
xor U13788 (N_13788,N_12401,N_12563);
nor U13789 (N_13789,N_12874,N_12036);
nand U13790 (N_13790,N_12927,N_12910);
and U13791 (N_13791,N_12186,N_12044);
or U13792 (N_13792,N_12410,N_12472);
and U13793 (N_13793,N_12080,N_12384);
or U13794 (N_13794,N_12498,N_12212);
nor U13795 (N_13795,N_12345,N_12381);
or U13796 (N_13796,N_12761,N_12781);
nor U13797 (N_13797,N_12494,N_12383);
nor U13798 (N_13798,N_12090,N_12248);
nor U13799 (N_13799,N_12994,N_12789);
xor U13800 (N_13800,N_12225,N_12141);
nor U13801 (N_13801,N_12414,N_12949);
or U13802 (N_13802,N_12139,N_12660);
xor U13803 (N_13803,N_12986,N_12188);
or U13804 (N_13804,N_12711,N_12769);
or U13805 (N_13805,N_12287,N_12603);
nand U13806 (N_13806,N_12205,N_12935);
xnor U13807 (N_13807,N_12298,N_12399);
nor U13808 (N_13808,N_12216,N_12052);
or U13809 (N_13809,N_12012,N_12052);
xnor U13810 (N_13810,N_12199,N_12038);
and U13811 (N_13811,N_12275,N_12476);
or U13812 (N_13812,N_12686,N_12223);
or U13813 (N_13813,N_12128,N_12858);
nor U13814 (N_13814,N_12452,N_12123);
xor U13815 (N_13815,N_12604,N_12518);
nor U13816 (N_13816,N_12538,N_12012);
or U13817 (N_13817,N_12213,N_12088);
xnor U13818 (N_13818,N_12983,N_12546);
and U13819 (N_13819,N_12210,N_12921);
nand U13820 (N_13820,N_12919,N_12794);
nor U13821 (N_13821,N_12855,N_12961);
and U13822 (N_13822,N_12322,N_12089);
and U13823 (N_13823,N_12532,N_12786);
nand U13824 (N_13824,N_12156,N_12074);
nor U13825 (N_13825,N_12700,N_12007);
or U13826 (N_13826,N_12915,N_12889);
and U13827 (N_13827,N_12791,N_12262);
nand U13828 (N_13828,N_12598,N_12738);
nor U13829 (N_13829,N_12595,N_12122);
nand U13830 (N_13830,N_12006,N_12525);
and U13831 (N_13831,N_12935,N_12629);
nor U13832 (N_13832,N_12929,N_12122);
and U13833 (N_13833,N_12793,N_12870);
or U13834 (N_13834,N_12385,N_12094);
or U13835 (N_13835,N_12004,N_12010);
nor U13836 (N_13836,N_12288,N_12613);
xnor U13837 (N_13837,N_12046,N_12988);
xor U13838 (N_13838,N_12383,N_12125);
or U13839 (N_13839,N_12373,N_12353);
nor U13840 (N_13840,N_12908,N_12783);
xor U13841 (N_13841,N_12727,N_12476);
or U13842 (N_13842,N_12936,N_12916);
or U13843 (N_13843,N_12154,N_12493);
or U13844 (N_13844,N_12280,N_12294);
and U13845 (N_13845,N_12452,N_12685);
xor U13846 (N_13846,N_12386,N_12050);
and U13847 (N_13847,N_12507,N_12922);
xnor U13848 (N_13848,N_12170,N_12590);
or U13849 (N_13849,N_12926,N_12785);
and U13850 (N_13850,N_12529,N_12738);
and U13851 (N_13851,N_12286,N_12786);
or U13852 (N_13852,N_12936,N_12763);
xor U13853 (N_13853,N_12002,N_12993);
xor U13854 (N_13854,N_12040,N_12789);
or U13855 (N_13855,N_12584,N_12134);
nor U13856 (N_13856,N_12221,N_12187);
xnor U13857 (N_13857,N_12480,N_12194);
nand U13858 (N_13858,N_12998,N_12789);
nand U13859 (N_13859,N_12873,N_12368);
or U13860 (N_13860,N_12858,N_12422);
nor U13861 (N_13861,N_12761,N_12743);
nor U13862 (N_13862,N_12694,N_12242);
xnor U13863 (N_13863,N_12722,N_12031);
or U13864 (N_13864,N_12552,N_12106);
xor U13865 (N_13865,N_12971,N_12288);
nand U13866 (N_13866,N_12429,N_12454);
and U13867 (N_13867,N_12679,N_12918);
nand U13868 (N_13868,N_12131,N_12137);
nand U13869 (N_13869,N_12103,N_12830);
nor U13870 (N_13870,N_12370,N_12575);
nand U13871 (N_13871,N_12516,N_12417);
xnor U13872 (N_13872,N_12484,N_12734);
or U13873 (N_13873,N_12185,N_12745);
nand U13874 (N_13874,N_12525,N_12543);
nor U13875 (N_13875,N_12373,N_12913);
xnor U13876 (N_13876,N_12258,N_12825);
or U13877 (N_13877,N_12906,N_12086);
or U13878 (N_13878,N_12853,N_12594);
or U13879 (N_13879,N_12878,N_12851);
or U13880 (N_13880,N_12043,N_12656);
xnor U13881 (N_13881,N_12150,N_12158);
xnor U13882 (N_13882,N_12489,N_12790);
xnor U13883 (N_13883,N_12042,N_12577);
nand U13884 (N_13884,N_12126,N_12441);
nor U13885 (N_13885,N_12119,N_12176);
xor U13886 (N_13886,N_12449,N_12674);
xor U13887 (N_13887,N_12610,N_12122);
and U13888 (N_13888,N_12593,N_12412);
nand U13889 (N_13889,N_12972,N_12624);
xor U13890 (N_13890,N_12562,N_12844);
nor U13891 (N_13891,N_12378,N_12099);
nor U13892 (N_13892,N_12197,N_12504);
or U13893 (N_13893,N_12180,N_12148);
xnor U13894 (N_13894,N_12635,N_12190);
or U13895 (N_13895,N_12141,N_12496);
nor U13896 (N_13896,N_12549,N_12292);
and U13897 (N_13897,N_12609,N_12271);
and U13898 (N_13898,N_12660,N_12715);
or U13899 (N_13899,N_12647,N_12064);
or U13900 (N_13900,N_12638,N_12884);
xor U13901 (N_13901,N_12696,N_12450);
or U13902 (N_13902,N_12016,N_12932);
nand U13903 (N_13903,N_12125,N_12691);
or U13904 (N_13904,N_12669,N_12548);
xor U13905 (N_13905,N_12148,N_12897);
or U13906 (N_13906,N_12643,N_12533);
or U13907 (N_13907,N_12719,N_12799);
nor U13908 (N_13908,N_12100,N_12951);
or U13909 (N_13909,N_12994,N_12837);
xnor U13910 (N_13910,N_12919,N_12357);
and U13911 (N_13911,N_12296,N_12728);
nand U13912 (N_13912,N_12153,N_12004);
or U13913 (N_13913,N_12598,N_12156);
or U13914 (N_13914,N_12513,N_12050);
or U13915 (N_13915,N_12991,N_12309);
nand U13916 (N_13916,N_12526,N_12242);
nand U13917 (N_13917,N_12663,N_12715);
nor U13918 (N_13918,N_12005,N_12655);
or U13919 (N_13919,N_12922,N_12346);
nor U13920 (N_13920,N_12395,N_12583);
nand U13921 (N_13921,N_12175,N_12819);
xor U13922 (N_13922,N_12182,N_12268);
or U13923 (N_13923,N_12234,N_12498);
nor U13924 (N_13924,N_12580,N_12547);
nor U13925 (N_13925,N_12535,N_12473);
xor U13926 (N_13926,N_12845,N_12102);
and U13927 (N_13927,N_12166,N_12951);
or U13928 (N_13928,N_12609,N_12051);
xnor U13929 (N_13929,N_12433,N_12738);
and U13930 (N_13930,N_12251,N_12408);
xor U13931 (N_13931,N_12562,N_12820);
nand U13932 (N_13932,N_12961,N_12656);
nor U13933 (N_13933,N_12111,N_12440);
nand U13934 (N_13934,N_12101,N_12711);
and U13935 (N_13935,N_12606,N_12164);
or U13936 (N_13936,N_12444,N_12261);
and U13937 (N_13937,N_12222,N_12056);
nor U13938 (N_13938,N_12328,N_12465);
nand U13939 (N_13939,N_12714,N_12461);
or U13940 (N_13940,N_12204,N_12115);
nand U13941 (N_13941,N_12063,N_12250);
and U13942 (N_13942,N_12677,N_12988);
or U13943 (N_13943,N_12688,N_12482);
nand U13944 (N_13944,N_12631,N_12183);
or U13945 (N_13945,N_12423,N_12330);
nand U13946 (N_13946,N_12843,N_12861);
nor U13947 (N_13947,N_12576,N_12136);
nand U13948 (N_13948,N_12126,N_12202);
xor U13949 (N_13949,N_12808,N_12032);
xnor U13950 (N_13950,N_12776,N_12831);
nand U13951 (N_13951,N_12812,N_12977);
and U13952 (N_13952,N_12704,N_12419);
nor U13953 (N_13953,N_12799,N_12235);
or U13954 (N_13954,N_12971,N_12332);
nand U13955 (N_13955,N_12852,N_12668);
and U13956 (N_13956,N_12356,N_12183);
xnor U13957 (N_13957,N_12349,N_12725);
nand U13958 (N_13958,N_12213,N_12180);
and U13959 (N_13959,N_12272,N_12894);
or U13960 (N_13960,N_12980,N_12977);
xnor U13961 (N_13961,N_12816,N_12403);
nand U13962 (N_13962,N_12041,N_12080);
xor U13963 (N_13963,N_12303,N_12190);
and U13964 (N_13964,N_12037,N_12749);
nor U13965 (N_13965,N_12330,N_12741);
or U13966 (N_13966,N_12904,N_12758);
nor U13967 (N_13967,N_12344,N_12706);
nor U13968 (N_13968,N_12543,N_12778);
and U13969 (N_13969,N_12440,N_12600);
xor U13970 (N_13970,N_12495,N_12826);
or U13971 (N_13971,N_12999,N_12648);
xor U13972 (N_13972,N_12391,N_12821);
nand U13973 (N_13973,N_12820,N_12408);
or U13974 (N_13974,N_12703,N_12518);
and U13975 (N_13975,N_12469,N_12271);
and U13976 (N_13976,N_12447,N_12664);
and U13977 (N_13977,N_12600,N_12243);
xor U13978 (N_13978,N_12718,N_12759);
or U13979 (N_13979,N_12780,N_12648);
and U13980 (N_13980,N_12465,N_12057);
nand U13981 (N_13981,N_12036,N_12317);
nand U13982 (N_13982,N_12675,N_12284);
and U13983 (N_13983,N_12200,N_12480);
nor U13984 (N_13984,N_12482,N_12000);
nor U13985 (N_13985,N_12146,N_12662);
nor U13986 (N_13986,N_12076,N_12662);
nand U13987 (N_13987,N_12447,N_12406);
xor U13988 (N_13988,N_12973,N_12101);
or U13989 (N_13989,N_12973,N_12478);
and U13990 (N_13990,N_12542,N_12193);
or U13991 (N_13991,N_12795,N_12380);
nor U13992 (N_13992,N_12281,N_12145);
nor U13993 (N_13993,N_12812,N_12130);
nor U13994 (N_13994,N_12124,N_12943);
nand U13995 (N_13995,N_12147,N_12526);
xor U13996 (N_13996,N_12156,N_12173);
or U13997 (N_13997,N_12542,N_12320);
nor U13998 (N_13998,N_12917,N_12527);
and U13999 (N_13999,N_12491,N_12275);
nand U14000 (N_14000,N_13693,N_13296);
or U14001 (N_14001,N_13179,N_13147);
nor U14002 (N_14002,N_13608,N_13029);
nand U14003 (N_14003,N_13956,N_13631);
xnor U14004 (N_14004,N_13444,N_13416);
and U14005 (N_14005,N_13541,N_13396);
nand U14006 (N_14006,N_13536,N_13820);
nor U14007 (N_14007,N_13790,N_13648);
xnor U14008 (N_14008,N_13874,N_13867);
nor U14009 (N_14009,N_13316,N_13824);
nand U14010 (N_14010,N_13393,N_13748);
xor U14011 (N_14011,N_13586,N_13896);
or U14012 (N_14012,N_13294,N_13499);
and U14013 (N_14013,N_13616,N_13273);
or U14014 (N_14014,N_13638,N_13921);
xor U14015 (N_14015,N_13251,N_13598);
and U14016 (N_14016,N_13597,N_13665);
nand U14017 (N_14017,N_13359,N_13442);
nand U14018 (N_14018,N_13569,N_13252);
nor U14019 (N_14019,N_13836,N_13568);
nor U14020 (N_14020,N_13967,N_13657);
nor U14021 (N_14021,N_13300,N_13002);
or U14022 (N_14022,N_13533,N_13011);
nand U14023 (N_14023,N_13732,N_13329);
xor U14024 (N_14024,N_13429,N_13534);
and U14025 (N_14025,N_13045,N_13198);
and U14026 (N_14026,N_13245,N_13105);
and U14027 (N_14027,N_13588,N_13057);
nand U14028 (N_14028,N_13843,N_13879);
or U14029 (N_14029,N_13126,N_13152);
or U14030 (N_14030,N_13766,N_13233);
or U14031 (N_14031,N_13942,N_13003);
xnor U14032 (N_14032,N_13215,N_13783);
nor U14033 (N_14033,N_13621,N_13523);
nand U14034 (N_14034,N_13338,N_13256);
nand U14035 (N_14035,N_13821,N_13791);
or U14036 (N_14036,N_13788,N_13682);
xnor U14037 (N_14037,N_13734,N_13760);
nand U14038 (N_14038,N_13862,N_13059);
or U14039 (N_14039,N_13165,N_13009);
nand U14040 (N_14040,N_13004,N_13283);
or U14041 (N_14041,N_13873,N_13288);
or U14042 (N_14042,N_13096,N_13040);
or U14043 (N_14043,N_13809,N_13100);
xnor U14044 (N_14044,N_13992,N_13812);
and U14045 (N_14045,N_13117,N_13542);
nor U14046 (N_14046,N_13438,N_13019);
xor U14047 (N_14047,N_13595,N_13979);
xnor U14048 (N_14048,N_13630,N_13472);
nor U14049 (N_14049,N_13346,N_13448);
nor U14050 (N_14050,N_13954,N_13973);
nor U14051 (N_14051,N_13938,N_13155);
nand U14052 (N_14052,N_13394,N_13168);
and U14053 (N_14053,N_13557,N_13082);
nor U14054 (N_14054,N_13209,N_13030);
or U14055 (N_14055,N_13320,N_13015);
and U14056 (N_14056,N_13347,N_13871);
xnor U14057 (N_14057,N_13414,N_13471);
nor U14058 (N_14058,N_13982,N_13644);
or U14059 (N_14059,N_13380,N_13697);
and U14060 (N_14060,N_13343,N_13340);
or U14061 (N_14061,N_13699,N_13102);
nor U14062 (N_14062,N_13049,N_13708);
nand U14063 (N_14063,N_13959,N_13620);
xnor U14064 (N_14064,N_13845,N_13513);
nand U14065 (N_14065,N_13714,N_13650);
nand U14066 (N_14066,N_13033,N_13039);
nand U14067 (N_14067,N_13728,N_13287);
or U14068 (N_14068,N_13835,N_13086);
and U14069 (N_14069,N_13014,N_13281);
xor U14070 (N_14070,N_13231,N_13461);
nand U14071 (N_14071,N_13143,N_13888);
nor U14072 (N_14072,N_13998,N_13626);
xnor U14073 (N_14073,N_13684,N_13724);
nor U14074 (N_14074,N_13409,N_13988);
or U14075 (N_14075,N_13312,N_13418);
xor U14076 (N_14076,N_13280,N_13218);
and U14077 (N_14077,N_13885,N_13151);
or U14078 (N_14078,N_13801,N_13431);
nand U14079 (N_14079,N_13107,N_13585);
nor U14080 (N_14080,N_13913,N_13512);
or U14081 (N_14081,N_13763,N_13356);
nor U14082 (N_14082,N_13206,N_13920);
nand U14083 (N_14083,N_13103,N_13480);
nor U14084 (N_14084,N_13926,N_13455);
or U14085 (N_14085,N_13309,N_13929);
nor U14086 (N_14086,N_13439,N_13705);
and U14087 (N_14087,N_13656,N_13263);
nand U14088 (N_14088,N_13232,N_13997);
or U14089 (N_14089,N_13796,N_13468);
nand U14090 (N_14090,N_13158,N_13073);
and U14091 (N_14091,N_13905,N_13560);
nor U14092 (N_14092,N_13718,N_13055);
nor U14093 (N_14093,N_13555,N_13420);
nand U14094 (N_14094,N_13036,N_13698);
nand U14095 (N_14095,N_13433,N_13332);
and U14096 (N_14096,N_13031,N_13138);
nand U14097 (N_14097,N_13304,N_13028);
nand U14098 (N_14098,N_13654,N_13012);
nor U14099 (N_14099,N_13743,N_13917);
nor U14100 (N_14100,N_13322,N_13407);
and U14101 (N_14101,N_13238,N_13310);
or U14102 (N_14102,N_13771,N_13141);
nand U14103 (N_14103,N_13047,N_13326);
xor U14104 (N_14104,N_13694,N_13087);
and U14105 (N_14105,N_13001,N_13328);
and U14106 (N_14106,N_13813,N_13331);
nor U14107 (N_14107,N_13951,N_13254);
nand U14108 (N_14108,N_13689,N_13991);
and U14109 (N_14109,N_13008,N_13205);
or U14110 (N_14110,N_13805,N_13878);
or U14111 (N_14111,N_13483,N_13357);
or U14112 (N_14112,N_13118,N_13576);
or U14113 (N_14113,N_13750,N_13278);
and U14114 (N_14114,N_13731,N_13563);
xnor U14115 (N_14115,N_13176,N_13677);
and U14116 (N_14116,N_13594,N_13277);
xor U14117 (N_14117,N_13735,N_13700);
nor U14118 (N_14118,N_13432,N_13434);
nand U14119 (N_14119,N_13108,N_13174);
xor U14120 (N_14120,N_13860,N_13244);
nand U14121 (N_14121,N_13514,N_13520);
nand U14122 (N_14122,N_13833,N_13119);
and U14123 (N_14123,N_13149,N_13032);
xnor U14124 (N_14124,N_13787,N_13160);
and U14125 (N_14125,N_13747,N_13506);
nand U14126 (N_14126,N_13419,N_13491);
xnor U14127 (N_14127,N_13501,N_13016);
and U14128 (N_14128,N_13260,N_13071);
and U14129 (N_14129,N_13671,N_13792);
nor U14130 (N_14130,N_13901,N_13239);
or U14131 (N_14131,N_13084,N_13266);
nand U14132 (N_14132,N_13659,N_13828);
nand U14133 (N_14133,N_13977,N_13891);
and U14134 (N_14134,N_13305,N_13646);
nand U14135 (N_14135,N_13981,N_13823);
xnor U14136 (N_14136,N_13655,N_13890);
nand U14137 (N_14137,N_13240,N_13208);
and U14138 (N_14138,N_13567,N_13246);
nor U14139 (N_14139,N_13410,N_13148);
nor U14140 (N_14140,N_13530,N_13027);
or U14141 (N_14141,N_13966,N_13164);
or U14142 (N_14142,N_13894,N_13302);
or U14143 (N_14143,N_13866,N_13053);
nand U14144 (N_14144,N_13781,N_13863);
or U14145 (N_14145,N_13056,N_13274);
and U14146 (N_14146,N_13802,N_13180);
nor U14147 (N_14147,N_13345,N_13270);
and U14148 (N_14148,N_13996,N_13315);
or U14149 (N_14149,N_13962,N_13319);
and U14150 (N_14150,N_13167,N_13856);
nand U14151 (N_14151,N_13234,N_13295);
xor U14152 (N_14152,N_13465,N_13456);
or U14153 (N_14153,N_13607,N_13189);
or U14154 (N_14154,N_13341,N_13949);
or U14155 (N_14155,N_13947,N_13733);
and U14156 (N_14156,N_13974,N_13615);
nor U14157 (N_14157,N_13127,N_13848);
and U14158 (N_14158,N_13545,N_13154);
nand U14159 (N_14159,N_13637,N_13844);
nand U14160 (N_14160,N_13464,N_13371);
and U14161 (N_14161,N_13069,N_13399);
xor U14162 (N_14162,N_13388,N_13253);
and U14163 (N_14163,N_13619,N_13195);
and U14164 (N_14164,N_13235,N_13043);
or U14165 (N_14165,N_13837,N_13457);
xnor U14166 (N_14166,N_13772,N_13293);
nor U14167 (N_14167,N_13928,N_13144);
and U14168 (N_14168,N_13384,N_13518);
nand U14169 (N_14169,N_13784,N_13739);
and U14170 (N_14170,N_13649,N_13112);
or U14171 (N_14171,N_13354,N_13330);
or U14172 (N_14172,N_13193,N_13869);
and U14173 (N_14173,N_13060,N_13083);
or U14174 (N_14174,N_13614,N_13681);
or U14175 (N_14175,N_13793,N_13628);
nor U14176 (N_14176,N_13258,N_13970);
nand U14177 (N_14177,N_13818,N_13265);
nor U14178 (N_14178,N_13687,N_13170);
nor U14179 (N_14179,N_13192,N_13044);
nand U14180 (N_14180,N_13562,N_13908);
xor U14181 (N_14181,N_13271,N_13853);
nand U14182 (N_14182,N_13255,N_13488);
xor U14183 (N_14183,N_13831,N_13291);
or U14184 (N_14184,N_13889,N_13334);
nand U14185 (N_14185,N_13722,N_13589);
and U14186 (N_14186,N_13596,N_13768);
nor U14187 (N_14187,N_13720,N_13387);
xnor U14188 (N_14188,N_13382,N_13635);
nand U14189 (N_14189,N_13933,N_13919);
and U14190 (N_14190,N_13183,N_13441);
nor U14191 (N_14191,N_13276,N_13572);
nor U14192 (N_14192,N_13157,N_13660);
nor U14193 (N_14193,N_13551,N_13203);
or U14194 (N_14194,N_13746,N_13701);
or U14195 (N_14195,N_13489,N_13453);
or U14196 (N_14196,N_13507,N_13759);
xor U14197 (N_14197,N_13963,N_13153);
nand U14198 (N_14198,N_13115,N_13492);
nor U14199 (N_14199,N_13840,N_13777);
xnor U14200 (N_14200,N_13936,N_13090);
or U14201 (N_14201,N_13636,N_13599);
nor U14202 (N_14202,N_13079,N_13881);
nand U14203 (N_14203,N_13450,N_13046);
nor U14204 (N_14204,N_13696,N_13691);
nand U14205 (N_14205,N_13579,N_13524);
nor U14206 (N_14206,N_13368,N_13940);
xor U14207 (N_14207,N_13757,N_13526);
and U14208 (N_14208,N_13372,N_13738);
nand U14209 (N_14209,N_13651,N_13427);
and U14210 (N_14210,N_13093,N_13237);
xnor U14211 (N_14211,N_13261,N_13826);
nor U14212 (N_14212,N_13110,N_13565);
or U14213 (N_14213,N_13564,N_13900);
or U14214 (N_14214,N_13175,N_13712);
and U14215 (N_14215,N_13887,N_13652);
or U14216 (N_14216,N_13336,N_13484);
xnor U14217 (N_14217,N_13223,N_13404);
or U14218 (N_14218,N_13034,N_13425);
nand U14219 (N_14219,N_13504,N_13999);
and U14220 (N_14220,N_13751,N_13200);
or U14221 (N_14221,N_13552,N_13362);
nor U14222 (N_14222,N_13716,N_13130);
nor U14223 (N_14223,N_13375,N_13762);
nand U14224 (N_14224,N_13789,N_13634);
nand U14225 (N_14225,N_13476,N_13422);
and U14226 (N_14226,N_13965,N_13590);
or U14227 (N_14227,N_13451,N_13411);
nor U14228 (N_14228,N_13937,N_13642);
and U14229 (N_14229,N_13994,N_13035);
nand U14230 (N_14230,N_13201,N_13074);
or U14231 (N_14231,N_13612,N_13509);
nand U14232 (N_14232,N_13647,N_13306);
or U14233 (N_14233,N_13262,N_13786);
xor U14234 (N_14234,N_13876,N_13364);
nor U14235 (N_14235,N_13051,N_13606);
or U14236 (N_14236,N_13064,N_13898);
nor U14237 (N_14237,N_13953,N_13307);
xor U14238 (N_14238,N_13292,N_13097);
xnor U14239 (N_14239,N_13024,N_13975);
xnor U14240 (N_14240,N_13080,N_13686);
nand U14241 (N_14241,N_13186,N_13529);
nor U14242 (N_14242,N_13496,N_13946);
and U14243 (N_14243,N_13139,N_13544);
or U14244 (N_14244,N_13125,N_13600);
xnor U14245 (N_14245,N_13286,N_13111);
and U14246 (N_14246,N_13284,N_13782);
xor U14247 (N_14247,N_13910,N_13886);
nor U14248 (N_14248,N_13842,N_13669);
nand U14249 (N_14249,N_13213,N_13948);
or U14250 (N_14250,N_13473,N_13249);
nand U14251 (N_14251,N_13680,N_13452);
and U14252 (N_14252,N_13062,N_13383);
nor U14253 (N_14253,N_13632,N_13214);
and U14254 (N_14254,N_13884,N_13490);
xnor U14255 (N_14255,N_13521,N_13190);
nand U14256 (N_14256,N_13169,N_13171);
xnor U14257 (N_14257,N_13808,N_13785);
nor U14258 (N_14258,N_13197,N_13449);
xnor U14259 (N_14259,N_13725,N_13817);
nand U14260 (N_14260,N_13868,N_13538);
nor U14261 (N_14261,N_13230,N_13577);
and U14262 (N_14262,N_13578,N_13104);
or U14263 (N_14263,N_13798,N_13548);
and U14264 (N_14264,N_13976,N_13402);
or U14265 (N_14265,N_13516,N_13156);
or U14266 (N_14266,N_13350,N_13892);
xnor U14267 (N_14267,N_13764,N_13730);
xor U14268 (N_14268,N_13077,N_13945);
xor U14269 (N_14269,N_13709,N_13986);
nor U14270 (N_14270,N_13389,N_13072);
nor U14271 (N_14271,N_13711,N_13406);
nand U14272 (N_14272,N_13961,N_13778);
nor U14273 (N_14273,N_13641,N_13374);
or U14274 (N_14274,N_13454,N_13314);
and U14275 (N_14275,N_13395,N_13146);
xor U14276 (N_14276,N_13591,N_13150);
and U14277 (N_14277,N_13930,N_13690);
nor U14278 (N_14278,N_13290,N_13376);
nor U14279 (N_14279,N_13318,N_13078);
nand U14280 (N_14280,N_13745,N_13816);
nor U14281 (N_14281,N_13386,N_13931);
xor U14282 (N_14282,N_13692,N_13510);
or U14283 (N_14283,N_13458,N_13494);
or U14284 (N_14284,N_13497,N_13587);
and U14285 (N_14285,N_13365,N_13918);
and U14286 (N_14286,N_13715,N_13822);
nand U14287 (N_14287,N_13048,N_13352);
nor U14288 (N_14288,N_13633,N_13969);
or U14289 (N_14289,N_13242,N_13247);
xor U14290 (N_14290,N_13091,N_13737);
nor U14291 (N_14291,N_13505,N_13342);
nand U14292 (N_14292,N_13161,N_13726);
and U14293 (N_14293,N_13861,N_13566);
and U14294 (N_14294,N_13575,N_13241);
nand U14295 (N_14295,N_13194,N_13924);
nand U14296 (N_14296,N_13191,N_13116);
or U14297 (N_14297,N_13670,N_13559);
nor U14298 (N_14298,N_13617,N_13547);
nor U14299 (N_14299,N_13089,N_13369);
and U14300 (N_14300,N_13508,N_13775);
nor U14301 (N_14301,N_13553,N_13421);
and U14302 (N_14302,N_13610,N_13515);
and U14303 (N_14303,N_13417,N_13532);
nand U14304 (N_14304,N_13335,N_13006);
and U14305 (N_14305,N_13603,N_13990);
and U14306 (N_14306,N_13475,N_13582);
nand U14307 (N_14307,N_13611,N_13377);
or U14308 (N_14308,N_13339,N_13944);
nand U14309 (N_14309,N_13925,N_13436);
nand U14310 (N_14310,N_13769,N_13477);
xor U14311 (N_14311,N_13435,N_13248);
or U14312 (N_14312,N_13137,N_13640);
or U14313 (N_14313,N_13723,N_13695);
nor U14314 (N_14314,N_13971,N_13960);
nand U14315 (N_14315,N_13989,N_13806);
or U14316 (N_14316,N_13859,N_13478);
nor U14317 (N_14317,N_13841,N_13995);
xnor U14318 (N_14318,N_13145,N_13474);
and U14319 (N_14319,N_13756,N_13065);
xnor U14320 (N_14320,N_13795,N_13957);
and U14321 (N_14321,N_13907,N_13702);
and U14322 (N_14322,N_13401,N_13609);
and U14323 (N_14323,N_13543,N_13729);
nand U14324 (N_14324,N_13939,N_13212);
nor U14325 (N_14325,N_13527,N_13814);
nand U14326 (N_14326,N_13727,N_13958);
xor U14327 (N_14327,N_13366,N_13216);
or U14328 (N_14328,N_13173,N_13272);
nand U14329 (N_14329,N_13187,N_13199);
nand U14330 (N_14330,N_13672,N_13744);
and U14331 (N_14331,N_13094,N_13624);
or U14332 (N_14332,N_13184,N_13397);
and U14333 (N_14333,N_13487,N_13850);
nor U14334 (N_14334,N_13602,N_13865);
xnor U14335 (N_14335,N_13658,N_13437);
nand U14336 (N_14336,N_13182,N_13188);
and U14337 (N_14337,N_13353,N_13210);
nand U14338 (N_14338,N_13964,N_13202);
nand U14339 (N_14339,N_13275,N_13952);
xor U14340 (N_14340,N_13470,N_13704);
xnor U14341 (N_14341,N_13101,N_13325);
or U14342 (N_14342,N_13228,N_13282);
nand U14343 (N_14343,N_13317,N_13131);
nand U14344 (N_14344,N_13993,N_13005);
nor U14345 (N_14345,N_13462,N_13525);
nor U14346 (N_14346,N_13794,N_13554);
nand U14347 (N_14347,N_13870,N_13018);
or U14348 (N_14348,N_13679,N_13303);
or U14349 (N_14349,N_13941,N_13159);
nand U14350 (N_14350,N_13023,N_13259);
nand U14351 (N_14351,N_13909,N_13770);
xor U14352 (N_14352,N_13140,N_13075);
or U14353 (N_14353,N_13227,N_13172);
xnor U14354 (N_14354,N_13528,N_13927);
nand U14355 (N_14355,N_13392,N_13412);
xnor U14356 (N_14356,N_13629,N_13978);
and U14357 (N_14357,N_13264,N_13780);
nand U14358 (N_14358,N_13755,N_13911);
or U14359 (N_14359,N_13706,N_13875);
xnor U14360 (N_14360,N_13721,N_13400);
or U14361 (N_14361,N_13807,N_13899);
and U14362 (N_14362,N_13134,N_13710);
and U14363 (N_14363,N_13135,N_13181);
or U14364 (N_14364,N_13236,N_13855);
and U14365 (N_14365,N_13070,N_13313);
nor U14366 (N_14366,N_13639,N_13185);
or U14367 (N_14367,N_13593,N_13133);
xnor U14368 (N_14368,N_13267,N_13849);
xnor U14369 (N_14369,N_13351,N_13459);
or U14370 (N_14370,N_13381,N_13323);
nor U14371 (N_14371,N_13370,N_13297);
nand U14372 (N_14372,N_13765,N_13985);
xor U14373 (N_14373,N_13872,N_13021);
nor U14374 (N_14374,N_13955,N_13717);
or U14375 (N_14375,N_13675,N_13495);
or U14376 (N_14376,N_13136,N_13479);
xor U14377 (N_14377,N_13950,N_13613);
or U14378 (N_14378,N_13166,N_13882);
or U14379 (N_14379,N_13893,N_13022);
and U14380 (N_14380,N_13038,N_13854);
nor U14381 (N_14381,N_13486,N_13883);
or U14382 (N_14382,N_13664,N_13592);
nor U14383 (N_14383,N_13754,N_13207);
nor U14384 (N_14384,N_13570,N_13423);
nor U14385 (N_14385,N_13688,N_13851);
and U14386 (N_14386,N_13662,N_13561);
nor U14387 (N_14387,N_13467,N_13067);
xnor U14388 (N_14388,N_13289,N_13719);
nand U14389 (N_14389,N_13279,N_13776);
xnor U14390 (N_14390,N_13299,N_13061);
and U14391 (N_14391,N_13408,N_13324);
nand U14392 (N_14392,N_13758,N_13405);
xnor U14393 (N_14393,N_13810,N_13983);
nand U14394 (N_14394,N_13311,N_13819);
nand U14395 (N_14395,N_13852,N_13500);
nor U14396 (N_14396,N_13902,N_13349);
nand U14397 (N_14397,N_13604,N_13880);
nand U14398 (N_14398,N_13858,N_13229);
nor U14399 (N_14399,N_13968,N_13363);
xnor U14400 (N_14400,N_13385,N_13106);
nand U14401 (N_14401,N_13799,N_13839);
or U14402 (N_14402,N_13428,N_13466);
nand U14403 (N_14403,N_13058,N_13327);
nor U14404 (N_14404,N_13774,N_13934);
nand U14405 (N_14405,N_13752,N_13398);
nand U14406 (N_14406,N_13123,N_13460);
xnor U14407 (N_14407,N_13558,N_13426);
nand U14408 (N_14408,N_13622,N_13736);
nor U14409 (N_14409,N_13413,N_13605);
xor U14410 (N_14410,N_13415,N_13224);
nand U14411 (N_14411,N_13403,N_13378);
xnor U14412 (N_14412,N_13076,N_13673);
nand U14413 (N_14413,N_13088,N_13980);
or U14414 (N_14414,N_13574,N_13095);
xor U14415 (N_14415,N_13742,N_13779);
xor U14416 (N_14416,N_13114,N_13447);
nor U14417 (N_14417,N_13661,N_13674);
or U14418 (N_14418,N_13469,N_13485);
and U14419 (N_14419,N_13667,N_13142);
nand U14420 (N_14420,N_13052,N_13539);
or U14421 (N_14421,N_13972,N_13222);
and U14422 (N_14422,N_13333,N_13128);
nor U14423 (N_14423,N_13132,N_13430);
nand U14424 (N_14424,N_13301,N_13618);
nand U14425 (N_14425,N_13099,N_13226);
nor U14426 (N_14426,N_13498,N_13804);
nor U14427 (N_14427,N_13519,N_13463);
nand U14428 (N_14428,N_13916,N_13803);
xor U14429 (N_14429,N_13540,N_13864);
nand U14430 (N_14430,N_13163,N_13571);
xnor U14431 (N_14431,N_13829,N_13042);
and U14432 (N_14432,N_13037,N_13827);
nand U14433 (N_14433,N_13493,N_13098);
xor U14434 (N_14434,N_13666,N_13129);
and U14435 (N_14435,N_13531,N_13741);
and U14436 (N_14436,N_13068,N_13627);
or U14437 (N_14437,N_13124,N_13749);
nor U14438 (N_14438,N_13683,N_13549);
and U14439 (N_14439,N_13020,N_13800);
xnor U14440 (N_14440,N_13285,N_13122);
nand U14441 (N_14441,N_13026,N_13811);
and U14442 (N_14442,N_13573,N_13987);
or U14443 (N_14443,N_13121,N_13391);
or U14444 (N_14444,N_13815,N_13580);
and U14445 (N_14445,N_13676,N_13767);
xor U14446 (N_14446,N_13857,N_13217);
and U14447 (N_14447,N_13601,N_13321);
or U14448 (N_14448,N_13025,N_13066);
nand U14449 (N_14449,N_13196,N_13269);
and U14450 (N_14450,N_13838,N_13984);
nand U14451 (N_14451,N_13424,N_13922);
xor U14452 (N_14452,N_13482,N_13740);
nand U14453 (N_14453,N_13085,N_13643);
and U14454 (N_14454,N_13050,N_13550);
nand U14455 (N_14455,N_13503,N_13897);
and U14456 (N_14456,N_13109,N_13063);
and U14457 (N_14457,N_13379,N_13443);
xor U14458 (N_14458,N_13943,N_13007);
xnor U14459 (N_14459,N_13625,N_13308);
or U14460 (N_14460,N_13663,N_13162);
nand U14461 (N_14461,N_13903,N_13847);
xnor U14462 (N_14462,N_13846,N_13517);
xor U14463 (N_14463,N_13348,N_13010);
and U14464 (N_14464,N_13906,N_13113);
or U14465 (N_14465,N_13932,N_13713);
xor U14466 (N_14466,N_13877,N_13703);
or U14467 (N_14467,N_13583,N_13935);
nor U14468 (N_14468,N_13546,N_13355);
or U14469 (N_14469,N_13390,N_13753);
nor U14470 (N_14470,N_13537,N_13225);
xnor U14471 (N_14471,N_13645,N_13219);
nand U14472 (N_14472,N_13337,N_13707);
nand U14473 (N_14473,N_13367,N_13511);
nand U14474 (N_14474,N_13268,N_13211);
and U14475 (N_14475,N_13502,N_13668);
nor U14476 (N_14476,N_13535,N_13360);
or U14477 (N_14477,N_13678,N_13204);
and U14478 (N_14478,N_13834,N_13481);
nor U14479 (N_14479,N_13221,N_13081);
and U14480 (N_14480,N_13446,N_13177);
xnor U14481 (N_14481,N_13653,N_13120);
nand U14482 (N_14482,N_13923,N_13220);
or U14483 (N_14483,N_13797,N_13623);
and U14484 (N_14484,N_13257,N_13915);
and U14485 (N_14485,N_13440,N_13522);
xnor U14486 (N_14486,N_13358,N_13825);
nand U14487 (N_14487,N_13361,N_13773);
xor U14488 (N_14488,N_13914,N_13373);
nor U14489 (N_14489,N_13243,N_13445);
nor U14490 (N_14490,N_13904,N_13685);
nor U14491 (N_14491,N_13832,N_13761);
nor U14492 (N_14492,N_13000,N_13912);
and U14493 (N_14493,N_13344,N_13092);
nand U14494 (N_14494,N_13041,N_13584);
xor U14495 (N_14495,N_13250,N_13017);
nand U14496 (N_14496,N_13895,N_13013);
nor U14497 (N_14497,N_13830,N_13298);
nor U14498 (N_14498,N_13556,N_13054);
or U14499 (N_14499,N_13178,N_13581);
nor U14500 (N_14500,N_13001,N_13093);
and U14501 (N_14501,N_13542,N_13529);
and U14502 (N_14502,N_13291,N_13451);
or U14503 (N_14503,N_13446,N_13558);
nor U14504 (N_14504,N_13648,N_13441);
or U14505 (N_14505,N_13211,N_13504);
nor U14506 (N_14506,N_13468,N_13433);
or U14507 (N_14507,N_13878,N_13443);
or U14508 (N_14508,N_13256,N_13366);
nand U14509 (N_14509,N_13166,N_13849);
nor U14510 (N_14510,N_13037,N_13508);
or U14511 (N_14511,N_13738,N_13481);
and U14512 (N_14512,N_13844,N_13054);
nor U14513 (N_14513,N_13312,N_13862);
nor U14514 (N_14514,N_13028,N_13038);
xor U14515 (N_14515,N_13635,N_13919);
or U14516 (N_14516,N_13422,N_13602);
and U14517 (N_14517,N_13034,N_13423);
xnor U14518 (N_14518,N_13929,N_13103);
xor U14519 (N_14519,N_13250,N_13075);
nand U14520 (N_14520,N_13015,N_13007);
and U14521 (N_14521,N_13036,N_13392);
and U14522 (N_14522,N_13209,N_13184);
nand U14523 (N_14523,N_13704,N_13285);
nor U14524 (N_14524,N_13441,N_13101);
or U14525 (N_14525,N_13540,N_13000);
or U14526 (N_14526,N_13115,N_13409);
nand U14527 (N_14527,N_13578,N_13354);
xor U14528 (N_14528,N_13911,N_13604);
nor U14529 (N_14529,N_13032,N_13577);
xnor U14530 (N_14530,N_13059,N_13227);
xor U14531 (N_14531,N_13258,N_13877);
nor U14532 (N_14532,N_13732,N_13838);
nor U14533 (N_14533,N_13258,N_13322);
and U14534 (N_14534,N_13462,N_13681);
nor U14535 (N_14535,N_13385,N_13989);
or U14536 (N_14536,N_13622,N_13050);
xor U14537 (N_14537,N_13423,N_13931);
nand U14538 (N_14538,N_13169,N_13476);
xnor U14539 (N_14539,N_13468,N_13356);
nor U14540 (N_14540,N_13808,N_13751);
and U14541 (N_14541,N_13025,N_13414);
nand U14542 (N_14542,N_13724,N_13068);
or U14543 (N_14543,N_13114,N_13738);
xor U14544 (N_14544,N_13022,N_13590);
nor U14545 (N_14545,N_13540,N_13384);
and U14546 (N_14546,N_13641,N_13620);
or U14547 (N_14547,N_13458,N_13008);
and U14548 (N_14548,N_13965,N_13849);
xor U14549 (N_14549,N_13900,N_13764);
or U14550 (N_14550,N_13003,N_13476);
xnor U14551 (N_14551,N_13325,N_13110);
xor U14552 (N_14552,N_13023,N_13124);
or U14553 (N_14553,N_13694,N_13616);
and U14554 (N_14554,N_13297,N_13789);
or U14555 (N_14555,N_13362,N_13004);
xnor U14556 (N_14556,N_13559,N_13741);
or U14557 (N_14557,N_13776,N_13862);
nand U14558 (N_14558,N_13312,N_13186);
or U14559 (N_14559,N_13625,N_13966);
nor U14560 (N_14560,N_13100,N_13830);
or U14561 (N_14561,N_13555,N_13144);
xor U14562 (N_14562,N_13928,N_13751);
and U14563 (N_14563,N_13756,N_13985);
xor U14564 (N_14564,N_13073,N_13962);
nand U14565 (N_14565,N_13645,N_13080);
and U14566 (N_14566,N_13969,N_13616);
and U14567 (N_14567,N_13352,N_13713);
nand U14568 (N_14568,N_13288,N_13222);
nand U14569 (N_14569,N_13262,N_13505);
xnor U14570 (N_14570,N_13500,N_13034);
or U14571 (N_14571,N_13411,N_13050);
and U14572 (N_14572,N_13399,N_13329);
nor U14573 (N_14573,N_13032,N_13692);
or U14574 (N_14574,N_13699,N_13742);
xor U14575 (N_14575,N_13980,N_13922);
xor U14576 (N_14576,N_13052,N_13278);
and U14577 (N_14577,N_13031,N_13847);
nor U14578 (N_14578,N_13508,N_13443);
xnor U14579 (N_14579,N_13539,N_13250);
nand U14580 (N_14580,N_13841,N_13261);
and U14581 (N_14581,N_13033,N_13895);
xor U14582 (N_14582,N_13591,N_13059);
nor U14583 (N_14583,N_13426,N_13640);
nand U14584 (N_14584,N_13056,N_13821);
or U14585 (N_14585,N_13477,N_13267);
or U14586 (N_14586,N_13754,N_13919);
nand U14587 (N_14587,N_13681,N_13386);
and U14588 (N_14588,N_13580,N_13471);
nor U14589 (N_14589,N_13631,N_13578);
nand U14590 (N_14590,N_13020,N_13426);
nor U14591 (N_14591,N_13362,N_13900);
or U14592 (N_14592,N_13301,N_13907);
nor U14593 (N_14593,N_13482,N_13616);
and U14594 (N_14594,N_13241,N_13431);
and U14595 (N_14595,N_13241,N_13593);
nand U14596 (N_14596,N_13986,N_13675);
xnor U14597 (N_14597,N_13623,N_13390);
and U14598 (N_14598,N_13743,N_13452);
or U14599 (N_14599,N_13036,N_13569);
xor U14600 (N_14600,N_13080,N_13020);
and U14601 (N_14601,N_13549,N_13661);
nand U14602 (N_14602,N_13993,N_13294);
and U14603 (N_14603,N_13554,N_13225);
nand U14604 (N_14604,N_13699,N_13938);
and U14605 (N_14605,N_13712,N_13918);
xor U14606 (N_14606,N_13023,N_13676);
nand U14607 (N_14607,N_13607,N_13447);
and U14608 (N_14608,N_13115,N_13825);
nor U14609 (N_14609,N_13278,N_13131);
or U14610 (N_14610,N_13958,N_13205);
xnor U14611 (N_14611,N_13608,N_13516);
or U14612 (N_14612,N_13711,N_13673);
nor U14613 (N_14613,N_13119,N_13889);
nand U14614 (N_14614,N_13473,N_13001);
nand U14615 (N_14615,N_13149,N_13921);
xnor U14616 (N_14616,N_13743,N_13978);
nor U14617 (N_14617,N_13970,N_13082);
nor U14618 (N_14618,N_13691,N_13311);
xor U14619 (N_14619,N_13085,N_13909);
nor U14620 (N_14620,N_13596,N_13923);
and U14621 (N_14621,N_13315,N_13701);
nor U14622 (N_14622,N_13968,N_13136);
nand U14623 (N_14623,N_13616,N_13007);
xnor U14624 (N_14624,N_13216,N_13858);
and U14625 (N_14625,N_13677,N_13595);
nand U14626 (N_14626,N_13168,N_13806);
nand U14627 (N_14627,N_13196,N_13838);
and U14628 (N_14628,N_13847,N_13712);
and U14629 (N_14629,N_13491,N_13231);
and U14630 (N_14630,N_13614,N_13703);
xor U14631 (N_14631,N_13149,N_13774);
nand U14632 (N_14632,N_13998,N_13622);
or U14633 (N_14633,N_13330,N_13841);
nor U14634 (N_14634,N_13162,N_13433);
and U14635 (N_14635,N_13432,N_13630);
or U14636 (N_14636,N_13288,N_13537);
xnor U14637 (N_14637,N_13668,N_13986);
or U14638 (N_14638,N_13362,N_13039);
or U14639 (N_14639,N_13931,N_13570);
nand U14640 (N_14640,N_13625,N_13926);
nor U14641 (N_14641,N_13735,N_13985);
nor U14642 (N_14642,N_13490,N_13736);
and U14643 (N_14643,N_13102,N_13467);
nand U14644 (N_14644,N_13656,N_13507);
or U14645 (N_14645,N_13133,N_13586);
nand U14646 (N_14646,N_13327,N_13127);
nor U14647 (N_14647,N_13006,N_13247);
xnor U14648 (N_14648,N_13415,N_13030);
nand U14649 (N_14649,N_13515,N_13316);
xnor U14650 (N_14650,N_13617,N_13512);
and U14651 (N_14651,N_13218,N_13252);
xnor U14652 (N_14652,N_13221,N_13662);
nand U14653 (N_14653,N_13067,N_13684);
nor U14654 (N_14654,N_13941,N_13759);
nor U14655 (N_14655,N_13655,N_13937);
nand U14656 (N_14656,N_13733,N_13949);
nor U14657 (N_14657,N_13058,N_13560);
nor U14658 (N_14658,N_13146,N_13568);
nand U14659 (N_14659,N_13556,N_13793);
nor U14660 (N_14660,N_13261,N_13452);
or U14661 (N_14661,N_13569,N_13805);
and U14662 (N_14662,N_13105,N_13441);
or U14663 (N_14663,N_13470,N_13265);
and U14664 (N_14664,N_13043,N_13643);
and U14665 (N_14665,N_13729,N_13850);
nand U14666 (N_14666,N_13265,N_13808);
and U14667 (N_14667,N_13643,N_13410);
xnor U14668 (N_14668,N_13187,N_13313);
or U14669 (N_14669,N_13036,N_13235);
and U14670 (N_14670,N_13678,N_13694);
or U14671 (N_14671,N_13977,N_13381);
nand U14672 (N_14672,N_13837,N_13162);
or U14673 (N_14673,N_13263,N_13122);
xnor U14674 (N_14674,N_13039,N_13851);
nand U14675 (N_14675,N_13744,N_13846);
xor U14676 (N_14676,N_13228,N_13932);
nor U14677 (N_14677,N_13715,N_13744);
nor U14678 (N_14678,N_13836,N_13749);
nand U14679 (N_14679,N_13845,N_13618);
xor U14680 (N_14680,N_13121,N_13418);
nor U14681 (N_14681,N_13880,N_13707);
xor U14682 (N_14682,N_13300,N_13363);
nand U14683 (N_14683,N_13708,N_13179);
and U14684 (N_14684,N_13043,N_13069);
or U14685 (N_14685,N_13985,N_13205);
nor U14686 (N_14686,N_13790,N_13722);
xnor U14687 (N_14687,N_13379,N_13297);
nand U14688 (N_14688,N_13983,N_13125);
xor U14689 (N_14689,N_13397,N_13546);
nand U14690 (N_14690,N_13917,N_13018);
xor U14691 (N_14691,N_13938,N_13266);
and U14692 (N_14692,N_13018,N_13899);
or U14693 (N_14693,N_13919,N_13380);
nor U14694 (N_14694,N_13103,N_13922);
or U14695 (N_14695,N_13896,N_13002);
xnor U14696 (N_14696,N_13053,N_13401);
and U14697 (N_14697,N_13799,N_13390);
nor U14698 (N_14698,N_13331,N_13738);
xor U14699 (N_14699,N_13923,N_13940);
xnor U14700 (N_14700,N_13688,N_13554);
and U14701 (N_14701,N_13387,N_13075);
nand U14702 (N_14702,N_13358,N_13956);
and U14703 (N_14703,N_13113,N_13015);
nand U14704 (N_14704,N_13720,N_13593);
nand U14705 (N_14705,N_13695,N_13915);
xor U14706 (N_14706,N_13110,N_13907);
and U14707 (N_14707,N_13773,N_13208);
nor U14708 (N_14708,N_13789,N_13150);
and U14709 (N_14709,N_13238,N_13046);
nor U14710 (N_14710,N_13520,N_13697);
xor U14711 (N_14711,N_13791,N_13505);
xnor U14712 (N_14712,N_13583,N_13721);
and U14713 (N_14713,N_13939,N_13653);
xnor U14714 (N_14714,N_13206,N_13627);
nand U14715 (N_14715,N_13302,N_13001);
xnor U14716 (N_14716,N_13366,N_13547);
and U14717 (N_14717,N_13164,N_13852);
and U14718 (N_14718,N_13805,N_13734);
or U14719 (N_14719,N_13036,N_13748);
nand U14720 (N_14720,N_13014,N_13066);
xnor U14721 (N_14721,N_13805,N_13385);
xor U14722 (N_14722,N_13410,N_13651);
nor U14723 (N_14723,N_13179,N_13989);
nor U14724 (N_14724,N_13474,N_13774);
xor U14725 (N_14725,N_13422,N_13824);
xnor U14726 (N_14726,N_13940,N_13591);
and U14727 (N_14727,N_13769,N_13525);
nor U14728 (N_14728,N_13586,N_13997);
or U14729 (N_14729,N_13143,N_13383);
and U14730 (N_14730,N_13469,N_13243);
nand U14731 (N_14731,N_13507,N_13480);
or U14732 (N_14732,N_13018,N_13053);
nor U14733 (N_14733,N_13673,N_13834);
and U14734 (N_14734,N_13662,N_13927);
nor U14735 (N_14735,N_13701,N_13599);
or U14736 (N_14736,N_13119,N_13982);
xor U14737 (N_14737,N_13191,N_13267);
and U14738 (N_14738,N_13797,N_13847);
nor U14739 (N_14739,N_13759,N_13778);
nand U14740 (N_14740,N_13318,N_13996);
xor U14741 (N_14741,N_13979,N_13967);
and U14742 (N_14742,N_13906,N_13538);
or U14743 (N_14743,N_13293,N_13831);
or U14744 (N_14744,N_13022,N_13677);
or U14745 (N_14745,N_13957,N_13301);
and U14746 (N_14746,N_13081,N_13603);
xnor U14747 (N_14747,N_13295,N_13628);
or U14748 (N_14748,N_13568,N_13355);
nand U14749 (N_14749,N_13961,N_13532);
or U14750 (N_14750,N_13359,N_13157);
nor U14751 (N_14751,N_13687,N_13990);
nand U14752 (N_14752,N_13356,N_13954);
or U14753 (N_14753,N_13432,N_13168);
xnor U14754 (N_14754,N_13960,N_13689);
or U14755 (N_14755,N_13747,N_13751);
xnor U14756 (N_14756,N_13683,N_13979);
and U14757 (N_14757,N_13437,N_13537);
nor U14758 (N_14758,N_13354,N_13373);
nor U14759 (N_14759,N_13945,N_13986);
xor U14760 (N_14760,N_13881,N_13696);
nor U14761 (N_14761,N_13014,N_13155);
or U14762 (N_14762,N_13320,N_13248);
xor U14763 (N_14763,N_13232,N_13908);
and U14764 (N_14764,N_13925,N_13500);
nand U14765 (N_14765,N_13179,N_13866);
or U14766 (N_14766,N_13615,N_13883);
or U14767 (N_14767,N_13808,N_13497);
nor U14768 (N_14768,N_13594,N_13207);
and U14769 (N_14769,N_13852,N_13912);
or U14770 (N_14770,N_13655,N_13710);
nor U14771 (N_14771,N_13871,N_13494);
nand U14772 (N_14772,N_13937,N_13788);
and U14773 (N_14773,N_13713,N_13339);
nand U14774 (N_14774,N_13702,N_13352);
and U14775 (N_14775,N_13372,N_13786);
or U14776 (N_14776,N_13903,N_13122);
and U14777 (N_14777,N_13928,N_13475);
nand U14778 (N_14778,N_13597,N_13028);
nand U14779 (N_14779,N_13827,N_13956);
nand U14780 (N_14780,N_13854,N_13912);
and U14781 (N_14781,N_13272,N_13665);
xor U14782 (N_14782,N_13377,N_13591);
and U14783 (N_14783,N_13840,N_13992);
or U14784 (N_14784,N_13117,N_13808);
and U14785 (N_14785,N_13589,N_13710);
or U14786 (N_14786,N_13199,N_13203);
or U14787 (N_14787,N_13327,N_13968);
xnor U14788 (N_14788,N_13448,N_13084);
or U14789 (N_14789,N_13333,N_13311);
nand U14790 (N_14790,N_13231,N_13044);
and U14791 (N_14791,N_13702,N_13450);
xor U14792 (N_14792,N_13480,N_13367);
xor U14793 (N_14793,N_13580,N_13054);
nor U14794 (N_14794,N_13831,N_13642);
and U14795 (N_14795,N_13598,N_13499);
or U14796 (N_14796,N_13392,N_13550);
nor U14797 (N_14797,N_13938,N_13413);
or U14798 (N_14798,N_13480,N_13487);
nand U14799 (N_14799,N_13387,N_13136);
and U14800 (N_14800,N_13649,N_13398);
and U14801 (N_14801,N_13977,N_13039);
nor U14802 (N_14802,N_13787,N_13521);
and U14803 (N_14803,N_13110,N_13321);
nor U14804 (N_14804,N_13987,N_13910);
nand U14805 (N_14805,N_13663,N_13690);
and U14806 (N_14806,N_13791,N_13929);
and U14807 (N_14807,N_13442,N_13681);
nand U14808 (N_14808,N_13493,N_13927);
or U14809 (N_14809,N_13501,N_13447);
or U14810 (N_14810,N_13904,N_13388);
and U14811 (N_14811,N_13996,N_13466);
nand U14812 (N_14812,N_13497,N_13081);
and U14813 (N_14813,N_13085,N_13539);
nand U14814 (N_14814,N_13295,N_13958);
and U14815 (N_14815,N_13415,N_13497);
nand U14816 (N_14816,N_13488,N_13084);
nand U14817 (N_14817,N_13533,N_13057);
xor U14818 (N_14818,N_13233,N_13013);
nand U14819 (N_14819,N_13027,N_13454);
xor U14820 (N_14820,N_13697,N_13907);
nor U14821 (N_14821,N_13255,N_13542);
xnor U14822 (N_14822,N_13568,N_13783);
and U14823 (N_14823,N_13727,N_13953);
nor U14824 (N_14824,N_13463,N_13385);
or U14825 (N_14825,N_13752,N_13544);
nand U14826 (N_14826,N_13505,N_13873);
nand U14827 (N_14827,N_13360,N_13380);
and U14828 (N_14828,N_13291,N_13292);
and U14829 (N_14829,N_13978,N_13888);
and U14830 (N_14830,N_13425,N_13119);
nor U14831 (N_14831,N_13788,N_13070);
and U14832 (N_14832,N_13080,N_13755);
and U14833 (N_14833,N_13431,N_13595);
xor U14834 (N_14834,N_13161,N_13789);
and U14835 (N_14835,N_13910,N_13120);
nand U14836 (N_14836,N_13594,N_13834);
xor U14837 (N_14837,N_13087,N_13926);
nor U14838 (N_14838,N_13908,N_13524);
or U14839 (N_14839,N_13329,N_13633);
or U14840 (N_14840,N_13247,N_13996);
or U14841 (N_14841,N_13184,N_13009);
or U14842 (N_14842,N_13113,N_13312);
and U14843 (N_14843,N_13816,N_13799);
or U14844 (N_14844,N_13192,N_13199);
or U14845 (N_14845,N_13706,N_13674);
xor U14846 (N_14846,N_13861,N_13880);
nor U14847 (N_14847,N_13673,N_13836);
xnor U14848 (N_14848,N_13847,N_13806);
and U14849 (N_14849,N_13156,N_13997);
xnor U14850 (N_14850,N_13206,N_13610);
or U14851 (N_14851,N_13041,N_13251);
nor U14852 (N_14852,N_13077,N_13747);
nor U14853 (N_14853,N_13829,N_13068);
or U14854 (N_14854,N_13507,N_13318);
xor U14855 (N_14855,N_13233,N_13855);
xnor U14856 (N_14856,N_13206,N_13163);
or U14857 (N_14857,N_13644,N_13529);
or U14858 (N_14858,N_13658,N_13527);
or U14859 (N_14859,N_13752,N_13181);
and U14860 (N_14860,N_13871,N_13358);
and U14861 (N_14861,N_13097,N_13140);
nand U14862 (N_14862,N_13863,N_13631);
nor U14863 (N_14863,N_13979,N_13441);
xnor U14864 (N_14864,N_13852,N_13233);
and U14865 (N_14865,N_13073,N_13150);
nand U14866 (N_14866,N_13402,N_13063);
nand U14867 (N_14867,N_13971,N_13672);
xor U14868 (N_14868,N_13875,N_13663);
xor U14869 (N_14869,N_13254,N_13495);
and U14870 (N_14870,N_13085,N_13176);
nor U14871 (N_14871,N_13392,N_13434);
and U14872 (N_14872,N_13633,N_13698);
xor U14873 (N_14873,N_13724,N_13245);
xnor U14874 (N_14874,N_13364,N_13242);
nor U14875 (N_14875,N_13893,N_13543);
nor U14876 (N_14876,N_13015,N_13767);
nand U14877 (N_14877,N_13337,N_13031);
or U14878 (N_14878,N_13034,N_13522);
nand U14879 (N_14879,N_13545,N_13664);
nand U14880 (N_14880,N_13233,N_13422);
nand U14881 (N_14881,N_13906,N_13850);
nand U14882 (N_14882,N_13103,N_13824);
nor U14883 (N_14883,N_13524,N_13354);
nor U14884 (N_14884,N_13844,N_13192);
xnor U14885 (N_14885,N_13329,N_13488);
nand U14886 (N_14886,N_13475,N_13469);
xnor U14887 (N_14887,N_13184,N_13499);
or U14888 (N_14888,N_13203,N_13336);
xor U14889 (N_14889,N_13903,N_13340);
or U14890 (N_14890,N_13478,N_13253);
xnor U14891 (N_14891,N_13371,N_13028);
nand U14892 (N_14892,N_13202,N_13835);
xnor U14893 (N_14893,N_13694,N_13008);
nor U14894 (N_14894,N_13829,N_13529);
and U14895 (N_14895,N_13102,N_13616);
or U14896 (N_14896,N_13626,N_13507);
nand U14897 (N_14897,N_13324,N_13400);
and U14898 (N_14898,N_13141,N_13811);
and U14899 (N_14899,N_13120,N_13666);
nor U14900 (N_14900,N_13794,N_13904);
nor U14901 (N_14901,N_13486,N_13297);
nand U14902 (N_14902,N_13140,N_13070);
nor U14903 (N_14903,N_13257,N_13011);
or U14904 (N_14904,N_13989,N_13452);
or U14905 (N_14905,N_13641,N_13945);
and U14906 (N_14906,N_13832,N_13820);
and U14907 (N_14907,N_13906,N_13863);
xnor U14908 (N_14908,N_13979,N_13293);
and U14909 (N_14909,N_13318,N_13806);
xnor U14910 (N_14910,N_13977,N_13358);
xnor U14911 (N_14911,N_13368,N_13731);
nand U14912 (N_14912,N_13278,N_13314);
nand U14913 (N_14913,N_13644,N_13654);
or U14914 (N_14914,N_13256,N_13418);
and U14915 (N_14915,N_13672,N_13507);
nand U14916 (N_14916,N_13315,N_13017);
and U14917 (N_14917,N_13064,N_13576);
and U14918 (N_14918,N_13364,N_13237);
nand U14919 (N_14919,N_13348,N_13017);
and U14920 (N_14920,N_13863,N_13636);
xor U14921 (N_14921,N_13014,N_13490);
or U14922 (N_14922,N_13301,N_13392);
xnor U14923 (N_14923,N_13518,N_13463);
nor U14924 (N_14924,N_13019,N_13616);
or U14925 (N_14925,N_13055,N_13128);
and U14926 (N_14926,N_13426,N_13922);
and U14927 (N_14927,N_13326,N_13895);
xor U14928 (N_14928,N_13123,N_13410);
or U14929 (N_14929,N_13020,N_13699);
nor U14930 (N_14930,N_13132,N_13275);
nand U14931 (N_14931,N_13253,N_13892);
nand U14932 (N_14932,N_13849,N_13365);
nor U14933 (N_14933,N_13000,N_13119);
xor U14934 (N_14934,N_13615,N_13368);
or U14935 (N_14935,N_13440,N_13257);
nand U14936 (N_14936,N_13097,N_13492);
nor U14937 (N_14937,N_13835,N_13549);
nand U14938 (N_14938,N_13125,N_13568);
and U14939 (N_14939,N_13491,N_13366);
xor U14940 (N_14940,N_13652,N_13540);
and U14941 (N_14941,N_13531,N_13309);
and U14942 (N_14942,N_13031,N_13482);
nand U14943 (N_14943,N_13522,N_13101);
nor U14944 (N_14944,N_13422,N_13731);
or U14945 (N_14945,N_13463,N_13914);
nand U14946 (N_14946,N_13166,N_13367);
nor U14947 (N_14947,N_13742,N_13535);
xnor U14948 (N_14948,N_13845,N_13592);
or U14949 (N_14949,N_13485,N_13689);
nand U14950 (N_14950,N_13212,N_13806);
nand U14951 (N_14951,N_13481,N_13628);
nor U14952 (N_14952,N_13971,N_13193);
nor U14953 (N_14953,N_13287,N_13431);
and U14954 (N_14954,N_13724,N_13201);
xor U14955 (N_14955,N_13667,N_13827);
nand U14956 (N_14956,N_13378,N_13806);
nand U14957 (N_14957,N_13477,N_13179);
nand U14958 (N_14958,N_13330,N_13680);
nand U14959 (N_14959,N_13310,N_13902);
and U14960 (N_14960,N_13629,N_13919);
xor U14961 (N_14961,N_13463,N_13974);
or U14962 (N_14962,N_13694,N_13273);
nand U14963 (N_14963,N_13756,N_13867);
and U14964 (N_14964,N_13124,N_13557);
xnor U14965 (N_14965,N_13844,N_13449);
or U14966 (N_14966,N_13796,N_13675);
and U14967 (N_14967,N_13163,N_13389);
xnor U14968 (N_14968,N_13017,N_13629);
xor U14969 (N_14969,N_13850,N_13798);
xnor U14970 (N_14970,N_13750,N_13226);
xnor U14971 (N_14971,N_13241,N_13709);
nand U14972 (N_14972,N_13163,N_13626);
xnor U14973 (N_14973,N_13451,N_13393);
nor U14974 (N_14974,N_13791,N_13924);
and U14975 (N_14975,N_13669,N_13733);
and U14976 (N_14976,N_13410,N_13934);
nor U14977 (N_14977,N_13667,N_13892);
xor U14978 (N_14978,N_13632,N_13119);
or U14979 (N_14979,N_13155,N_13907);
xnor U14980 (N_14980,N_13443,N_13860);
or U14981 (N_14981,N_13386,N_13796);
xnor U14982 (N_14982,N_13271,N_13443);
nand U14983 (N_14983,N_13839,N_13143);
or U14984 (N_14984,N_13488,N_13340);
xor U14985 (N_14985,N_13789,N_13030);
nand U14986 (N_14986,N_13258,N_13947);
or U14987 (N_14987,N_13917,N_13269);
and U14988 (N_14988,N_13820,N_13070);
xnor U14989 (N_14989,N_13228,N_13862);
nor U14990 (N_14990,N_13664,N_13309);
xnor U14991 (N_14991,N_13947,N_13840);
xor U14992 (N_14992,N_13726,N_13703);
or U14993 (N_14993,N_13033,N_13653);
nand U14994 (N_14994,N_13701,N_13318);
or U14995 (N_14995,N_13923,N_13085);
or U14996 (N_14996,N_13938,N_13610);
nor U14997 (N_14997,N_13590,N_13956);
or U14998 (N_14998,N_13977,N_13320);
xor U14999 (N_14999,N_13377,N_13492);
or U15000 (N_15000,N_14120,N_14236);
nor U15001 (N_15001,N_14444,N_14544);
or U15002 (N_15002,N_14077,N_14469);
nand U15003 (N_15003,N_14428,N_14816);
nand U15004 (N_15004,N_14184,N_14643);
nand U15005 (N_15005,N_14953,N_14356);
xnor U15006 (N_15006,N_14827,N_14148);
or U15007 (N_15007,N_14114,N_14186);
or U15008 (N_15008,N_14113,N_14871);
or U15009 (N_15009,N_14758,N_14717);
and U15010 (N_15010,N_14795,N_14454);
xor U15011 (N_15011,N_14136,N_14368);
nand U15012 (N_15012,N_14941,N_14505);
or U15013 (N_15013,N_14354,N_14274);
nor U15014 (N_15014,N_14825,N_14894);
nor U15015 (N_15015,N_14310,N_14111);
nand U15016 (N_15016,N_14088,N_14338);
nor U15017 (N_15017,N_14439,N_14848);
or U15018 (N_15018,N_14786,N_14202);
and U15019 (N_15019,N_14245,N_14143);
or U15020 (N_15020,N_14597,N_14616);
and U15021 (N_15021,N_14079,N_14278);
and U15022 (N_15022,N_14966,N_14584);
xor U15023 (N_15023,N_14458,N_14563);
xnor U15024 (N_15024,N_14963,N_14060);
or U15025 (N_15025,N_14456,N_14002);
xor U15026 (N_15026,N_14714,N_14090);
or U15027 (N_15027,N_14750,N_14367);
or U15028 (N_15028,N_14414,N_14059);
nor U15029 (N_15029,N_14776,N_14523);
or U15030 (N_15030,N_14965,N_14728);
and U15031 (N_15031,N_14067,N_14460);
or U15032 (N_15032,N_14653,N_14430);
nor U15033 (N_15033,N_14527,N_14341);
nor U15034 (N_15034,N_14760,N_14247);
and U15035 (N_15035,N_14064,N_14753);
nand U15036 (N_15036,N_14238,N_14323);
and U15037 (N_15037,N_14945,N_14520);
nor U15038 (N_15038,N_14560,N_14076);
or U15039 (N_15039,N_14392,N_14098);
nor U15040 (N_15040,N_14438,N_14072);
and U15041 (N_15041,N_14618,N_14665);
xor U15042 (N_15042,N_14801,N_14054);
nand U15043 (N_15043,N_14057,N_14065);
and U15044 (N_15044,N_14969,N_14422);
xor U15045 (N_15045,N_14693,N_14904);
nor U15046 (N_15046,N_14929,N_14283);
or U15047 (N_15047,N_14780,N_14106);
and U15048 (N_15048,N_14187,N_14704);
nor U15049 (N_15049,N_14551,N_14348);
nor U15050 (N_15050,N_14897,N_14755);
or U15051 (N_15051,N_14126,N_14366);
or U15052 (N_15052,N_14003,N_14547);
xor U15053 (N_15053,N_14195,N_14974);
nand U15054 (N_15054,N_14888,N_14865);
and U15055 (N_15055,N_14504,N_14211);
and U15056 (N_15056,N_14706,N_14206);
nor U15057 (N_15057,N_14849,N_14992);
xor U15058 (N_15058,N_14474,N_14715);
xnor U15059 (N_15059,N_14982,N_14612);
or U15060 (N_15060,N_14398,N_14462);
nand U15061 (N_15061,N_14221,N_14068);
nand U15062 (N_15062,N_14431,N_14832);
nand U15063 (N_15063,N_14224,N_14287);
nor U15064 (N_15064,N_14978,N_14713);
xor U15065 (N_15065,N_14290,N_14554);
or U15066 (N_15066,N_14732,N_14699);
xnor U15067 (N_15067,N_14011,N_14025);
and U15068 (N_15068,N_14300,N_14617);
nand U15069 (N_15069,N_14977,N_14768);
and U15070 (N_15070,N_14410,N_14638);
or U15071 (N_15071,N_14402,N_14796);
or U15072 (N_15072,N_14679,N_14272);
xor U15073 (N_15073,N_14494,N_14053);
nand U15074 (N_15074,N_14731,N_14646);
and U15075 (N_15075,N_14898,N_14600);
and U15076 (N_15076,N_14027,N_14336);
or U15077 (N_15077,N_14937,N_14662);
nor U15078 (N_15078,N_14286,N_14263);
nand U15079 (N_15079,N_14455,N_14418);
nor U15080 (N_15080,N_14532,N_14809);
and U15081 (N_15081,N_14916,N_14540);
nor U15082 (N_15082,N_14075,N_14204);
and U15083 (N_15083,N_14491,N_14484);
xor U15084 (N_15084,N_14389,N_14103);
nand U15085 (N_15085,N_14362,N_14387);
or U15086 (N_15086,N_14522,N_14445);
and U15087 (N_15087,N_14810,N_14403);
xnor U15088 (N_15088,N_14483,N_14789);
or U15089 (N_15089,N_14481,N_14841);
nand U15090 (N_15090,N_14729,N_14426);
nor U15091 (N_15091,N_14819,N_14920);
xnor U15092 (N_15092,N_14457,N_14569);
or U15093 (N_15093,N_14196,N_14490);
and U15094 (N_15094,N_14495,N_14010);
nand U15095 (N_15095,N_14991,N_14337);
nor U15096 (N_15096,N_14382,N_14837);
and U15097 (N_15097,N_14641,N_14252);
nor U15098 (N_15098,N_14839,N_14411);
xor U15099 (N_15099,N_14331,N_14466);
nor U15100 (N_15100,N_14999,N_14413);
xnor U15101 (N_15101,N_14696,N_14149);
and U15102 (N_15102,N_14026,N_14710);
xor U15103 (N_15103,N_14749,N_14820);
nand U15104 (N_15104,N_14237,N_14774);
xor U15105 (N_15105,N_14767,N_14409);
xor U15106 (N_15106,N_14742,N_14799);
nor U15107 (N_15107,N_14762,N_14657);
xnor U15108 (N_15108,N_14826,N_14235);
nand U15109 (N_15109,N_14378,N_14595);
xnor U15110 (N_15110,N_14633,N_14655);
or U15111 (N_15111,N_14771,N_14640);
nand U15112 (N_15112,N_14203,N_14960);
and U15113 (N_15113,N_14461,N_14571);
xnor U15114 (N_15114,N_14950,N_14669);
xnor U15115 (N_15115,N_14927,N_14073);
and U15116 (N_15116,N_14770,N_14887);
and U15117 (N_15117,N_14257,N_14480);
or U15118 (N_15118,N_14117,N_14174);
and U15119 (N_15119,N_14216,N_14085);
and U15120 (N_15120,N_14123,N_14329);
and U15121 (N_15121,N_14754,N_14074);
nor U15122 (N_15122,N_14070,N_14385);
or U15123 (N_15123,N_14901,N_14166);
and U15124 (N_15124,N_14273,N_14509);
xnor U15125 (N_15125,N_14147,N_14488);
xnor U15126 (N_15126,N_14745,N_14516);
nand U15127 (N_15127,N_14427,N_14702);
and U15128 (N_15128,N_14535,N_14193);
xnor U15129 (N_15129,N_14759,N_14306);
nor U15130 (N_15130,N_14448,N_14518);
nand U15131 (N_15131,N_14205,N_14465);
xor U15132 (N_15132,N_14299,N_14349);
nand U15133 (N_15133,N_14215,N_14269);
nor U15134 (N_15134,N_14705,N_14515);
nor U15135 (N_15135,N_14160,N_14377);
nand U15136 (N_15136,N_14346,N_14083);
and U15137 (N_15137,N_14109,N_14823);
or U15138 (N_15138,N_14261,N_14862);
nor U15139 (N_15139,N_14364,N_14949);
and U15140 (N_15140,N_14021,N_14973);
nand U15141 (N_15141,N_14671,N_14814);
nor U15142 (N_15142,N_14987,N_14581);
or U15143 (N_15143,N_14536,N_14716);
xnor U15144 (N_15144,N_14676,N_14185);
or U15145 (N_15145,N_14276,N_14128);
and U15146 (N_15146,N_14830,N_14051);
or U15147 (N_15147,N_14319,N_14321);
nor U15148 (N_15148,N_14513,N_14824);
nand U15149 (N_15149,N_14621,N_14883);
or U15150 (N_15150,N_14947,N_14453);
nand U15151 (N_15151,N_14808,N_14089);
nand U15152 (N_15152,N_14675,N_14230);
xor U15153 (N_15153,N_14242,N_14399);
xnor U15154 (N_15154,N_14279,N_14962);
nor U15155 (N_15155,N_14511,N_14574);
and U15156 (N_15156,N_14589,N_14464);
xnor U15157 (N_15157,N_14983,N_14416);
nor U15158 (N_15158,N_14586,N_14254);
and U15159 (N_15159,N_14847,N_14163);
or U15160 (N_15160,N_14334,N_14086);
and U15161 (N_15161,N_14419,N_14328);
and U15162 (N_15162,N_14400,N_14219);
xor U15163 (N_15163,N_14437,N_14727);
nor U15164 (N_15164,N_14790,N_14878);
xor U15165 (N_15165,N_14256,N_14007);
and U15166 (N_15166,N_14548,N_14181);
nor U15167 (N_15167,N_14266,N_14441);
nand U15168 (N_15168,N_14353,N_14645);
nand U15169 (N_15169,N_14886,N_14118);
nand U15170 (N_15170,N_14900,N_14095);
nor U15171 (N_15171,N_14942,N_14957);
nand U15172 (N_15172,N_14986,N_14691);
nor U15173 (N_15173,N_14001,N_14097);
or U15174 (N_15174,N_14330,N_14327);
and U15175 (N_15175,N_14874,N_14844);
and U15176 (N_15176,N_14133,N_14890);
or U15177 (N_15177,N_14726,N_14531);
or U15178 (N_15178,N_14173,N_14688);
or U15179 (N_15179,N_14468,N_14802);
nor U15180 (N_15180,N_14333,N_14212);
nor U15181 (N_15181,N_14537,N_14159);
nand U15182 (N_15182,N_14647,N_14231);
nor U15183 (N_15183,N_14719,N_14023);
nor U15184 (N_15184,N_14765,N_14896);
nand U15185 (N_15185,N_14189,N_14043);
xnor U15186 (N_15186,N_14580,N_14359);
or U15187 (N_15187,N_14629,N_14100);
xor U15188 (N_15188,N_14127,N_14940);
nand U15189 (N_15189,N_14931,N_14734);
or U15190 (N_15190,N_14559,N_14066);
nand U15191 (N_15191,N_14994,N_14570);
xnor U15192 (N_15192,N_14194,N_14094);
and U15193 (N_15193,N_14250,N_14956);
and U15194 (N_15194,N_14158,N_14345);
xnor U15195 (N_15195,N_14698,N_14636);
xnor U15196 (N_15196,N_14358,N_14534);
and U15197 (N_15197,N_14817,N_14508);
xor U15198 (N_15198,N_14500,N_14093);
xor U15199 (N_15199,N_14778,N_14425);
and U15200 (N_15200,N_14583,N_14151);
nor U15201 (N_15201,N_14800,N_14502);
and U15202 (N_15202,N_14096,N_14663);
or U15203 (N_15203,N_14388,N_14512);
nand U15204 (N_15204,N_14039,N_14038);
xnor U15205 (N_15205,N_14294,N_14976);
nor U15206 (N_15206,N_14493,N_14668);
and U15207 (N_15207,N_14140,N_14078);
xnor U15208 (N_15208,N_14324,N_14615);
or U15209 (N_15209,N_14303,N_14867);
nand U15210 (N_15210,N_14694,N_14519);
nand U15211 (N_15211,N_14587,N_14594);
or U15212 (N_15212,N_14980,N_14239);
xnor U15213 (N_15213,N_14292,N_14452);
and U15214 (N_15214,N_14144,N_14712);
xor U15215 (N_15215,N_14546,N_14692);
nor U15216 (N_15216,N_14794,N_14008);
nand U15217 (N_15217,N_14320,N_14124);
nand U15218 (N_15218,N_14298,N_14666);
and U15219 (N_15219,N_14834,N_14661);
and U15220 (N_15220,N_14135,N_14415);
nor U15221 (N_15221,N_14659,N_14391);
or U15222 (N_15222,N_14838,N_14592);
and U15223 (N_15223,N_14751,N_14482);
nor U15224 (N_15224,N_14152,N_14225);
xnor U15225 (N_15225,N_14380,N_14280);
nor U15226 (N_15226,N_14525,N_14275);
xor U15227 (N_15227,N_14568,N_14339);
nand U15228 (N_15228,N_14132,N_14930);
nand U15229 (N_15229,N_14872,N_14222);
nand U15230 (N_15230,N_14471,N_14860);
nor U15231 (N_15231,N_14833,N_14463);
and U15232 (N_15232,N_14130,N_14855);
xnor U15233 (N_15233,N_14854,N_14701);
and U15234 (N_15234,N_14394,N_14139);
nor U15235 (N_15235,N_14177,N_14922);
xor U15236 (N_15236,N_14384,N_14308);
or U15237 (N_15237,N_14879,N_14861);
xnor U15238 (N_15238,N_14169,N_14030);
or U15239 (N_15239,N_14155,N_14209);
xnor U15240 (N_15240,N_14249,N_14335);
xor U15241 (N_15241,N_14302,N_14386);
xor U15242 (N_15242,N_14365,N_14542);
nor U15243 (N_15243,N_14869,N_14288);
xor U15244 (N_15244,N_14405,N_14539);
nand U15245 (N_15245,N_14793,N_14029);
nor U15246 (N_15246,N_14434,N_14932);
nand U15247 (N_15247,N_14910,N_14707);
or U15248 (N_15248,N_14325,N_14782);
nand U15249 (N_15249,N_14764,N_14440);
and U15250 (N_15250,N_14936,N_14036);
or U15251 (N_15251,N_14803,N_14424);
nand U15252 (N_15252,N_14406,N_14777);
xnor U15253 (N_15253,N_14876,N_14903);
nor U15254 (N_15254,N_14958,N_14926);
nor U15255 (N_15255,N_14603,N_14735);
nand U15256 (N_15256,N_14304,N_14743);
xor U15257 (N_15257,N_14044,N_14244);
nand U15258 (N_15258,N_14091,N_14375);
xnor U15259 (N_15259,N_14081,N_14214);
or U15260 (N_15260,N_14915,N_14138);
or U15261 (N_15261,N_14955,N_14253);
or U15262 (N_15262,N_14889,N_14572);
xnor U15263 (N_15263,N_14305,N_14747);
xor U15264 (N_15264,N_14575,N_14228);
and U15265 (N_15265,N_14626,N_14315);
nor U15266 (N_15266,N_14260,N_14251);
xor U15267 (N_15267,N_14582,N_14884);
and U15268 (N_15268,N_14052,N_14737);
nand U15269 (N_15269,N_14708,N_14881);
or U15270 (N_15270,N_14013,N_14034);
and U15271 (N_15271,N_14087,N_14614);
nor U15272 (N_15272,N_14567,N_14040);
and U15273 (N_15273,N_14161,N_14773);
or U15274 (N_15274,N_14557,N_14379);
or U15275 (N_15275,N_14864,N_14902);
or U15276 (N_15276,N_14198,N_14170);
nor U15277 (N_15277,N_14492,N_14047);
xnor U15278 (N_15278,N_14141,N_14099);
nor U15279 (N_15279,N_14284,N_14340);
and U15280 (N_15280,N_14909,N_14374);
and U15281 (N_15281,N_14813,N_14168);
or U15282 (N_15282,N_14805,N_14316);
xor U15283 (N_15283,N_14401,N_14882);
nor U15284 (N_15284,N_14162,N_14101);
nor U15285 (N_15285,N_14720,N_14852);
nand U15286 (N_15286,N_14550,N_14217);
nand U15287 (N_15287,N_14301,N_14923);
and U15288 (N_15288,N_14297,N_14895);
or U15289 (N_15289,N_14613,N_14993);
xnor U15290 (N_15290,N_14677,N_14733);
nor U15291 (N_15291,N_14223,N_14517);
and U15292 (N_15292,N_14703,N_14296);
and U15293 (N_15293,N_14639,N_14019);
xnor U15294 (N_15294,N_14906,N_14579);
nor U15295 (N_15295,N_14390,N_14718);
xnor U15296 (N_15296,N_14804,N_14351);
nand U15297 (N_15297,N_14110,N_14724);
and U15298 (N_15298,N_14635,N_14108);
nor U15299 (N_15299,N_14233,N_14851);
nor U15300 (N_15300,N_14119,N_14487);
or U15301 (N_15301,N_14009,N_14084);
nand U15302 (N_15302,N_14609,N_14450);
xnor U15303 (N_15303,N_14741,N_14192);
xnor U15304 (N_15304,N_14656,N_14016);
or U15305 (N_15305,N_14218,N_14309);
and U15306 (N_15306,N_14006,N_14711);
or U15307 (N_15307,N_14658,N_14918);
and U15308 (N_15308,N_14056,N_14420);
or U15309 (N_15309,N_14725,N_14408);
xor U15310 (N_15310,N_14673,N_14899);
nor U15311 (N_15311,N_14165,N_14970);
nor U15312 (N_15312,N_14107,N_14467);
nor U15313 (N_15313,N_14129,N_14530);
xor U15314 (N_15314,N_14180,N_14154);
xor U15315 (N_15315,N_14285,N_14892);
nand U15316 (N_15316,N_14921,N_14372);
and U15317 (N_15317,N_14840,N_14772);
nand U15318 (N_15318,N_14012,N_14479);
and U15319 (N_15319,N_14134,N_14623);
nor U15320 (N_15320,N_14499,N_14082);
or U15321 (N_15321,N_14566,N_14606);
and U15322 (N_15322,N_14905,N_14681);
and U15323 (N_15323,N_14891,N_14050);
nand U15324 (N_15324,N_14510,N_14024);
nor U15325 (N_15325,N_14037,N_14806);
and U15326 (N_15326,N_14829,N_14317);
or U15327 (N_15327,N_14648,N_14137);
and U15328 (N_15328,N_14478,N_14102);
xor U15329 (N_15329,N_14311,N_14031);
nand U15330 (N_15330,N_14875,N_14873);
or U15331 (N_15331,N_14763,N_14289);
nor U15332 (N_15332,N_14270,N_14553);
xor U15333 (N_15333,N_14689,N_14943);
xnor U15334 (N_15334,N_14291,N_14501);
and U15335 (N_15335,N_14684,N_14062);
nor U15336 (N_15336,N_14259,N_14475);
xor U15337 (N_15337,N_14045,N_14514);
nand U15338 (N_15338,N_14486,N_14925);
and U15339 (N_15339,N_14061,N_14775);
and U15340 (N_15340,N_14678,N_14226);
nand U15341 (N_15341,N_14815,N_14634);
and U15342 (N_15342,N_14271,N_14295);
xnor U15343 (N_15343,N_14447,N_14914);
xor U15344 (N_15344,N_14981,N_14080);
xnor U15345 (N_15345,N_14756,N_14821);
nand U15346 (N_15346,N_14831,N_14828);
or U15347 (N_15347,N_14856,N_14967);
xnor U15348 (N_15348,N_14652,N_14343);
nand U15349 (N_15349,N_14866,N_14241);
or U15350 (N_15350,N_14984,N_14243);
nand U15351 (N_15351,N_14210,N_14680);
nand U15352 (N_15352,N_14318,N_14361);
and U15353 (N_15353,N_14369,N_14761);
nor U15354 (N_15354,N_14432,N_14435);
nor U15355 (N_15355,N_14229,N_14443);
nand U15356 (N_15356,N_14277,N_14845);
xor U15357 (N_15357,N_14035,N_14220);
and U15358 (N_15358,N_14055,N_14893);
or U15359 (N_15359,N_14146,N_14370);
or U15360 (N_15360,N_14442,N_14541);
xnor U15361 (N_15361,N_14267,N_14588);
xor U15362 (N_15362,N_14783,N_14971);
nand U15363 (N_15363,N_14314,N_14015);
nor U15364 (N_15364,N_14934,N_14150);
xnor U15365 (N_15365,N_14545,N_14213);
and U15366 (N_15366,N_14654,N_14651);
nor U15367 (N_15367,N_14240,N_14561);
nor U15368 (N_15368,N_14470,N_14812);
xor U15369 (N_15369,N_14730,N_14262);
nor U15370 (N_15370,N_14017,N_14995);
nor U15371 (N_15371,N_14352,N_14000);
xor U15372 (N_15372,N_14004,N_14556);
or U15373 (N_15373,N_14171,N_14573);
nor U15374 (N_15374,N_14042,N_14631);
nand U15375 (N_15375,N_14281,N_14757);
xnor U15376 (N_15376,N_14020,N_14996);
xnor U15377 (N_15377,N_14779,N_14695);
xor U15378 (N_15378,N_14682,N_14627);
and U15379 (N_15379,N_14473,N_14429);
or U15380 (N_15380,N_14611,N_14234);
nor U15381 (N_15381,N_14131,N_14048);
nand U15382 (N_15382,N_14178,N_14912);
or U15383 (N_15383,N_14121,N_14690);
nor U15384 (N_15384,N_14459,N_14046);
nand U15385 (N_15385,N_14917,N_14997);
nand U15386 (N_15386,N_14938,N_14911);
nor U15387 (N_15387,N_14664,N_14208);
xor U15388 (N_15388,N_14877,N_14395);
and U15389 (N_15389,N_14928,N_14248);
nor U15390 (N_15390,N_14787,N_14788);
or U15391 (N_15391,N_14312,N_14990);
and U15392 (N_15392,N_14687,N_14863);
xor U15393 (N_15393,N_14069,N_14342);
nand U15394 (N_15394,N_14959,N_14552);
xor U15395 (N_15395,N_14122,N_14521);
xnor U15396 (N_15396,N_14625,N_14005);
xnor U15397 (N_15397,N_14620,N_14497);
xor U15398 (N_15398,N_14393,N_14766);
or U15399 (N_15399,N_14596,N_14125);
nor U15400 (N_15400,N_14989,N_14092);
or U15401 (N_15401,N_14964,N_14985);
nor U15402 (N_15402,N_14948,N_14642);
xor U15403 (N_15403,N_14028,N_14538);
nand U15404 (N_15404,N_14175,N_14112);
nand U15405 (N_15405,N_14397,N_14979);
or U15406 (N_15406,N_14752,N_14818);
or U15407 (N_15407,N_14565,N_14421);
and U15408 (N_15408,N_14578,N_14417);
nand U15409 (N_15409,N_14506,N_14373);
nand U15410 (N_15410,N_14954,N_14781);
xor U15411 (N_15411,N_14451,N_14396);
nand U15412 (N_15412,N_14179,N_14357);
xor U15413 (N_15413,N_14628,N_14748);
nand U15414 (N_15414,N_14630,N_14722);
nand U15415 (N_15415,N_14105,N_14907);
nand U15416 (N_15416,N_14489,N_14913);
nand U15417 (N_15417,N_14258,N_14857);
or U15418 (N_15418,N_14842,N_14822);
xnor U15419 (N_15419,N_14784,N_14649);
nor U15420 (N_15420,N_14674,N_14507);
and U15421 (N_15421,N_14182,N_14104);
nand U15422 (N_15422,N_14191,N_14407);
or U15423 (N_15423,N_14721,N_14988);
xnor U15424 (N_15424,N_14700,N_14610);
and U15425 (N_15425,N_14807,N_14293);
nand U15426 (N_15426,N_14738,N_14200);
nand U15427 (N_15427,N_14683,N_14939);
or U15428 (N_15428,N_14476,N_14919);
nand U15429 (N_15429,N_14371,N_14014);
or U15430 (N_15430,N_14326,N_14142);
or U15431 (N_15431,N_14885,N_14870);
nor U15432 (N_15432,N_14836,N_14798);
nand U15433 (N_15433,N_14951,N_14585);
nand U15434 (N_15434,N_14601,N_14412);
and U15435 (N_15435,N_14071,N_14032);
and U15436 (N_15436,N_14190,N_14858);
and U15437 (N_15437,N_14608,N_14156);
nor U15438 (N_15438,N_14853,N_14347);
xnor U15439 (N_15439,N_14167,N_14791);
or U15440 (N_15440,N_14153,N_14041);
and U15441 (N_15441,N_14360,N_14593);
and U15442 (N_15442,N_14558,N_14543);
xnor U15443 (N_15443,N_14496,N_14018);
or U15444 (N_15444,N_14355,N_14322);
nor U15445 (N_15445,N_14176,N_14622);
nand U15446 (N_15446,N_14785,N_14116);
xnor U15447 (N_15447,N_14199,N_14183);
or U15448 (N_15448,N_14590,N_14644);
nor U15449 (N_15449,N_14063,N_14404);
or U15450 (N_15450,N_14350,N_14528);
nand U15451 (N_15451,N_14723,N_14232);
xnor U15452 (N_15452,N_14555,N_14811);
and U15453 (N_15453,N_14255,N_14188);
and U15454 (N_15454,N_14598,N_14946);
xor U15455 (N_15455,N_14022,N_14564);
nand U15456 (N_15456,N_14498,N_14526);
nor U15457 (N_15457,N_14503,N_14058);
and U15458 (N_15458,N_14672,N_14268);
nand U15459 (N_15459,N_14933,N_14952);
xnor U15460 (N_15460,N_14577,N_14769);
nand U15461 (N_15461,N_14944,N_14332);
nand U15462 (N_15462,N_14792,N_14744);
and U15463 (N_15463,N_14591,N_14549);
xor U15464 (N_15464,N_14604,N_14605);
or U15465 (N_15465,N_14529,N_14576);
xnor U15466 (N_15466,N_14164,N_14197);
nor U15467 (N_15467,N_14201,N_14650);
nor U15468 (N_15468,N_14049,N_14961);
and U15469 (N_15469,N_14697,N_14172);
nor U15470 (N_15470,N_14797,N_14533);
and U15471 (N_15471,N_14908,N_14624);
or U15472 (N_15472,N_14868,N_14619);
and U15473 (N_15473,N_14363,N_14739);
or U15474 (N_15474,N_14307,N_14670);
nand U15475 (N_15475,N_14846,N_14383);
or U15476 (N_15476,N_14446,N_14033);
or U15477 (N_15477,N_14686,N_14968);
xor U15478 (N_15478,N_14850,N_14660);
nand U15479 (N_15479,N_14859,N_14265);
or U15480 (N_15480,N_14423,N_14313);
and U15481 (N_15481,N_14433,N_14472);
nor U15482 (N_15482,N_14436,N_14115);
nor U15483 (N_15483,N_14998,N_14449);
and U15484 (N_15484,N_14972,N_14975);
or U15485 (N_15485,N_14880,N_14736);
and U15486 (N_15486,N_14282,N_14835);
nand U15487 (N_15487,N_14602,N_14740);
or U15488 (N_15488,N_14485,N_14709);
nand U15489 (N_15489,N_14746,N_14344);
xor U15490 (N_15490,N_14843,N_14145);
nor U15491 (N_15491,N_14599,N_14524);
or U15492 (N_15492,N_14264,N_14207);
nand U15493 (N_15493,N_14562,N_14935);
nand U15494 (N_15494,N_14667,N_14637);
or U15495 (N_15495,N_14924,N_14157);
xor U15496 (N_15496,N_14227,N_14376);
nand U15497 (N_15497,N_14632,N_14477);
nand U15498 (N_15498,N_14685,N_14381);
nor U15499 (N_15499,N_14607,N_14246);
nor U15500 (N_15500,N_14048,N_14851);
nor U15501 (N_15501,N_14072,N_14387);
or U15502 (N_15502,N_14264,N_14647);
and U15503 (N_15503,N_14886,N_14360);
xor U15504 (N_15504,N_14254,N_14747);
nand U15505 (N_15505,N_14815,N_14761);
or U15506 (N_15506,N_14668,N_14443);
or U15507 (N_15507,N_14568,N_14305);
and U15508 (N_15508,N_14036,N_14388);
and U15509 (N_15509,N_14362,N_14975);
and U15510 (N_15510,N_14061,N_14503);
and U15511 (N_15511,N_14816,N_14161);
nor U15512 (N_15512,N_14764,N_14187);
and U15513 (N_15513,N_14641,N_14188);
xnor U15514 (N_15514,N_14775,N_14047);
xnor U15515 (N_15515,N_14372,N_14816);
and U15516 (N_15516,N_14881,N_14484);
nor U15517 (N_15517,N_14764,N_14977);
and U15518 (N_15518,N_14927,N_14492);
nor U15519 (N_15519,N_14093,N_14707);
nor U15520 (N_15520,N_14483,N_14707);
nand U15521 (N_15521,N_14030,N_14100);
nor U15522 (N_15522,N_14763,N_14320);
nand U15523 (N_15523,N_14759,N_14834);
or U15524 (N_15524,N_14088,N_14124);
and U15525 (N_15525,N_14737,N_14913);
nor U15526 (N_15526,N_14595,N_14467);
and U15527 (N_15527,N_14011,N_14451);
nor U15528 (N_15528,N_14523,N_14994);
or U15529 (N_15529,N_14029,N_14071);
nor U15530 (N_15530,N_14648,N_14338);
and U15531 (N_15531,N_14866,N_14611);
nor U15532 (N_15532,N_14663,N_14632);
and U15533 (N_15533,N_14426,N_14400);
xor U15534 (N_15534,N_14930,N_14337);
or U15535 (N_15535,N_14331,N_14049);
nor U15536 (N_15536,N_14657,N_14492);
nand U15537 (N_15537,N_14922,N_14596);
nor U15538 (N_15538,N_14737,N_14480);
nand U15539 (N_15539,N_14602,N_14592);
xnor U15540 (N_15540,N_14733,N_14233);
or U15541 (N_15541,N_14241,N_14978);
or U15542 (N_15542,N_14345,N_14957);
and U15543 (N_15543,N_14627,N_14797);
nor U15544 (N_15544,N_14557,N_14804);
nand U15545 (N_15545,N_14808,N_14437);
or U15546 (N_15546,N_14840,N_14064);
and U15547 (N_15547,N_14199,N_14738);
nor U15548 (N_15548,N_14397,N_14944);
xor U15549 (N_15549,N_14197,N_14029);
or U15550 (N_15550,N_14515,N_14806);
nand U15551 (N_15551,N_14406,N_14364);
xnor U15552 (N_15552,N_14209,N_14586);
xor U15553 (N_15553,N_14458,N_14033);
nor U15554 (N_15554,N_14770,N_14006);
or U15555 (N_15555,N_14814,N_14558);
or U15556 (N_15556,N_14848,N_14365);
and U15557 (N_15557,N_14879,N_14289);
and U15558 (N_15558,N_14270,N_14708);
and U15559 (N_15559,N_14432,N_14332);
nand U15560 (N_15560,N_14497,N_14759);
and U15561 (N_15561,N_14160,N_14460);
nor U15562 (N_15562,N_14641,N_14479);
nor U15563 (N_15563,N_14064,N_14546);
xnor U15564 (N_15564,N_14832,N_14134);
or U15565 (N_15565,N_14459,N_14135);
xnor U15566 (N_15566,N_14614,N_14719);
xnor U15567 (N_15567,N_14279,N_14421);
or U15568 (N_15568,N_14119,N_14413);
or U15569 (N_15569,N_14393,N_14450);
and U15570 (N_15570,N_14966,N_14562);
and U15571 (N_15571,N_14925,N_14383);
nor U15572 (N_15572,N_14356,N_14137);
xnor U15573 (N_15573,N_14237,N_14332);
xnor U15574 (N_15574,N_14165,N_14271);
nand U15575 (N_15575,N_14824,N_14430);
nand U15576 (N_15576,N_14172,N_14302);
and U15577 (N_15577,N_14416,N_14944);
and U15578 (N_15578,N_14971,N_14081);
and U15579 (N_15579,N_14465,N_14831);
nand U15580 (N_15580,N_14468,N_14657);
or U15581 (N_15581,N_14290,N_14423);
or U15582 (N_15582,N_14975,N_14009);
and U15583 (N_15583,N_14750,N_14097);
nand U15584 (N_15584,N_14629,N_14734);
nand U15585 (N_15585,N_14367,N_14003);
and U15586 (N_15586,N_14499,N_14653);
nand U15587 (N_15587,N_14838,N_14996);
nand U15588 (N_15588,N_14719,N_14546);
nand U15589 (N_15589,N_14122,N_14382);
xnor U15590 (N_15590,N_14223,N_14360);
nor U15591 (N_15591,N_14574,N_14549);
and U15592 (N_15592,N_14575,N_14184);
nand U15593 (N_15593,N_14460,N_14129);
and U15594 (N_15594,N_14728,N_14819);
and U15595 (N_15595,N_14808,N_14560);
nand U15596 (N_15596,N_14965,N_14318);
nor U15597 (N_15597,N_14315,N_14471);
or U15598 (N_15598,N_14646,N_14803);
or U15599 (N_15599,N_14826,N_14509);
and U15600 (N_15600,N_14428,N_14358);
and U15601 (N_15601,N_14630,N_14868);
nor U15602 (N_15602,N_14317,N_14764);
nor U15603 (N_15603,N_14100,N_14567);
nor U15604 (N_15604,N_14807,N_14459);
or U15605 (N_15605,N_14716,N_14848);
or U15606 (N_15606,N_14902,N_14845);
nand U15607 (N_15607,N_14879,N_14748);
nor U15608 (N_15608,N_14933,N_14371);
and U15609 (N_15609,N_14491,N_14257);
or U15610 (N_15610,N_14620,N_14108);
xor U15611 (N_15611,N_14966,N_14190);
nand U15612 (N_15612,N_14113,N_14070);
nand U15613 (N_15613,N_14368,N_14936);
or U15614 (N_15614,N_14367,N_14105);
and U15615 (N_15615,N_14658,N_14992);
nand U15616 (N_15616,N_14610,N_14693);
and U15617 (N_15617,N_14113,N_14625);
or U15618 (N_15618,N_14656,N_14663);
nand U15619 (N_15619,N_14705,N_14343);
nor U15620 (N_15620,N_14241,N_14459);
xnor U15621 (N_15621,N_14101,N_14284);
or U15622 (N_15622,N_14026,N_14591);
and U15623 (N_15623,N_14005,N_14137);
nand U15624 (N_15624,N_14966,N_14843);
xor U15625 (N_15625,N_14011,N_14449);
xnor U15626 (N_15626,N_14015,N_14732);
nand U15627 (N_15627,N_14372,N_14016);
xor U15628 (N_15628,N_14658,N_14810);
or U15629 (N_15629,N_14144,N_14325);
nor U15630 (N_15630,N_14041,N_14151);
nor U15631 (N_15631,N_14107,N_14237);
nor U15632 (N_15632,N_14732,N_14976);
nand U15633 (N_15633,N_14236,N_14143);
xnor U15634 (N_15634,N_14009,N_14355);
or U15635 (N_15635,N_14322,N_14202);
or U15636 (N_15636,N_14360,N_14858);
and U15637 (N_15637,N_14751,N_14371);
and U15638 (N_15638,N_14474,N_14570);
nand U15639 (N_15639,N_14872,N_14885);
nand U15640 (N_15640,N_14832,N_14396);
nor U15641 (N_15641,N_14593,N_14084);
nor U15642 (N_15642,N_14014,N_14657);
nand U15643 (N_15643,N_14479,N_14149);
and U15644 (N_15644,N_14882,N_14171);
and U15645 (N_15645,N_14741,N_14255);
xnor U15646 (N_15646,N_14692,N_14903);
nor U15647 (N_15647,N_14093,N_14686);
nand U15648 (N_15648,N_14003,N_14094);
nor U15649 (N_15649,N_14767,N_14689);
nor U15650 (N_15650,N_14376,N_14955);
xor U15651 (N_15651,N_14709,N_14511);
and U15652 (N_15652,N_14639,N_14053);
nand U15653 (N_15653,N_14022,N_14115);
nor U15654 (N_15654,N_14010,N_14206);
or U15655 (N_15655,N_14817,N_14561);
and U15656 (N_15656,N_14845,N_14658);
or U15657 (N_15657,N_14290,N_14396);
or U15658 (N_15658,N_14656,N_14611);
and U15659 (N_15659,N_14383,N_14138);
or U15660 (N_15660,N_14665,N_14493);
nand U15661 (N_15661,N_14992,N_14511);
xor U15662 (N_15662,N_14248,N_14745);
and U15663 (N_15663,N_14949,N_14550);
and U15664 (N_15664,N_14892,N_14491);
xor U15665 (N_15665,N_14797,N_14532);
or U15666 (N_15666,N_14324,N_14892);
and U15667 (N_15667,N_14863,N_14300);
nor U15668 (N_15668,N_14134,N_14667);
xnor U15669 (N_15669,N_14199,N_14813);
or U15670 (N_15670,N_14735,N_14253);
nor U15671 (N_15671,N_14140,N_14819);
nor U15672 (N_15672,N_14157,N_14908);
nor U15673 (N_15673,N_14785,N_14576);
nand U15674 (N_15674,N_14254,N_14231);
xor U15675 (N_15675,N_14401,N_14495);
or U15676 (N_15676,N_14909,N_14411);
nand U15677 (N_15677,N_14415,N_14275);
or U15678 (N_15678,N_14765,N_14328);
nor U15679 (N_15679,N_14939,N_14006);
and U15680 (N_15680,N_14755,N_14924);
and U15681 (N_15681,N_14891,N_14523);
nand U15682 (N_15682,N_14489,N_14634);
nor U15683 (N_15683,N_14552,N_14744);
nor U15684 (N_15684,N_14888,N_14861);
or U15685 (N_15685,N_14550,N_14972);
nand U15686 (N_15686,N_14283,N_14757);
xor U15687 (N_15687,N_14054,N_14080);
nand U15688 (N_15688,N_14765,N_14947);
nand U15689 (N_15689,N_14012,N_14995);
nor U15690 (N_15690,N_14815,N_14159);
nand U15691 (N_15691,N_14553,N_14499);
or U15692 (N_15692,N_14358,N_14505);
nand U15693 (N_15693,N_14293,N_14962);
nor U15694 (N_15694,N_14304,N_14264);
and U15695 (N_15695,N_14155,N_14435);
or U15696 (N_15696,N_14107,N_14804);
xnor U15697 (N_15697,N_14030,N_14754);
and U15698 (N_15698,N_14287,N_14380);
xnor U15699 (N_15699,N_14510,N_14853);
xor U15700 (N_15700,N_14932,N_14016);
or U15701 (N_15701,N_14793,N_14761);
xor U15702 (N_15702,N_14274,N_14911);
and U15703 (N_15703,N_14641,N_14574);
xor U15704 (N_15704,N_14018,N_14140);
nand U15705 (N_15705,N_14353,N_14891);
nand U15706 (N_15706,N_14336,N_14801);
and U15707 (N_15707,N_14928,N_14491);
and U15708 (N_15708,N_14394,N_14579);
nor U15709 (N_15709,N_14942,N_14469);
nor U15710 (N_15710,N_14041,N_14548);
and U15711 (N_15711,N_14517,N_14368);
nor U15712 (N_15712,N_14190,N_14537);
nor U15713 (N_15713,N_14013,N_14736);
or U15714 (N_15714,N_14467,N_14724);
or U15715 (N_15715,N_14606,N_14154);
nor U15716 (N_15716,N_14839,N_14241);
nand U15717 (N_15717,N_14698,N_14980);
nand U15718 (N_15718,N_14870,N_14417);
or U15719 (N_15719,N_14236,N_14383);
nor U15720 (N_15720,N_14637,N_14410);
nand U15721 (N_15721,N_14277,N_14282);
xor U15722 (N_15722,N_14669,N_14261);
nand U15723 (N_15723,N_14330,N_14055);
nor U15724 (N_15724,N_14100,N_14084);
nand U15725 (N_15725,N_14312,N_14366);
nand U15726 (N_15726,N_14587,N_14743);
nor U15727 (N_15727,N_14232,N_14359);
or U15728 (N_15728,N_14122,N_14316);
and U15729 (N_15729,N_14413,N_14387);
and U15730 (N_15730,N_14519,N_14658);
xnor U15731 (N_15731,N_14630,N_14534);
xor U15732 (N_15732,N_14044,N_14772);
xor U15733 (N_15733,N_14538,N_14217);
or U15734 (N_15734,N_14482,N_14912);
xnor U15735 (N_15735,N_14706,N_14857);
nand U15736 (N_15736,N_14102,N_14010);
nand U15737 (N_15737,N_14698,N_14828);
nand U15738 (N_15738,N_14886,N_14890);
nand U15739 (N_15739,N_14269,N_14875);
xnor U15740 (N_15740,N_14387,N_14388);
xor U15741 (N_15741,N_14109,N_14273);
nor U15742 (N_15742,N_14490,N_14438);
xor U15743 (N_15743,N_14317,N_14681);
nor U15744 (N_15744,N_14924,N_14717);
xnor U15745 (N_15745,N_14135,N_14937);
and U15746 (N_15746,N_14305,N_14457);
nand U15747 (N_15747,N_14370,N_14173);
and U15748 (N_15748,N_14175,N_14043);
nor U15749 (N_15749,N_14793,N_14827);
or U15750 (N_15750,N_14320,N_14402);
nor U15751 (N_15751,N_14822,N_14479);
xnor U15752 (N_15752,N_14307,N_14393);
and U15753 (N_15753,N_14069,N_14905);
xor U15754 (N_15754,N_14004,N_14546);
nand U15755 (N_15755,N_14451,N_14101);
and U15756 (N_15756,N_14976,N_14653);
or U15757 (N_15757,N_14706,N_14488);
or U15758 (N_15758,N_14248,N_14038);
nor U15759 (N_15759,N_14900,N_14918);
and U15760 (N_15760,N_14665,N_14903);
xnor U15761 (N_15761,N_14901,N_14672);
or U15762 (N_15762,N_14937,N_14088);
or U15763 (N_15763,N_14141,N_14107);
nor U15764 (N_15764,N_14788,N_14896);
nand U15765 (N_15765,N_14515,N_14813);
xnor U15766 (N_15766,N_14521,N_14235);
and U15767 (N_15767,N_14686,N_14667);
or U15768 (N_15768,N_14942,N_14007);
and U15769 (N_15769,N_14862,N_14665);
or U15770 (N_15770,N_14088,N_14198);
and U15771 (N_15771,N_14261,N_14676);
and U15772 (N_15772,N_14496,N_14263);
nor U15773 (N_15773,N_14068,N_14032);
nand U15774 (N_15774,N_14714,N_14473);
nand U15775 (N_15775,N_14094,N_14425);
xnor U15776 (N_15776,N_14192,N_14800);
or U15777 (N_15777,N_14743,N_14907);
xnor U15778 (N_15778,N_14258,N_14863);
and U15779 (N_15779,N_14570,N_14839);
nor U15780 (N_15780,N_14081,N_14768);
nor U15781 (N_15781,N_14579,N_14764);
nand U15782 (N_15782,N_14501,N_14485);
xor U15783 (N_15783,N_14750,N_14024);
xnor U15784 (N_15784,N_14107,N_14821);
nor U15785 (N_15785,N_14713,N_14099);
or U15786 (N_15786,N_14236,N_14345);
nand U15787 (N_15787,N_14710,N_14687);
and U15788 (N_15788,N_14057,N_14086);
xor U15789 (N_15789,N_14531,N_14999);
nor U15790 (N_15790,N_14681,N_14530);
nor U15791 (N_15791,N_14032,N_14791);
and U15792 (N_15792,N_14251,N_14681);
nor U15793 (N_15793,N_14238,N_14188);
nand U15794 (N_15794,N_14064,N_14080);
or U15795 (N_15795,N_14239,N_14950);
nor U15796 (N_15796,N_14482,N_14410);
xor U15797 (N_15797,N_14783,N_14590);
nand U15798 (N_15798,N_14292,N_14977);
xor U15799 (N_15799,N_14823,N_14597);
and U15800 (N_15800,N_14398,N_14433);
nor U15801 (N_15801,N_14248,N_14473);
or U15802 (N_15802,N_14673,N_14999);
xnor U15803 (N_15803,N_14271,N_14235);
xnor U15804 (N_15804,N_14221,N_14237);
xor U15805 (N_15805,N_14513,N_14496);
xor U15806 (N_15806,N_14415,N_14241);
or U15807 (N_15807,N_14727,N_14109);
nor U15808 (N_15808,N_14705,N_14534);
or U15809 (N_15809,N_14048,N_14110);
or U15810 (N_15810,N_14264,N_14749);
and U15811 (N_15811,N_14048,N_14116);
xor U15812 (N_15812,N_14858,N_14221);
and U15813 (N_15813,N_14588,N_14116);
or U15814 (N_15814,N_14097,N_14306);
nor U15815 (N_15815,N_14502,N_14378);
or U15816 (N_15816,N_14486,N_14321);
or U15817 (N_15817,N_14019,N_14419);
or U15818 (N_15818,N_14260,N_14708);
and U15819 (N_15819,N_14093,N_14299);
nand U15820 (N_15820,N_14482,N_14190);
xnor U15821 (N_15821,N_14795,N_14107);
nand U15822 (N_15822,N_14166,N_14276);
and U15823 (N_15823,N_14571,N_14049);
xor U15824 (N_15824,N_14981,N_14817);
and U15825 (N_15825,N_14866,N_14788);
and U15826 (N_15826,N_14294,N_14877);
xnor U15827 (N_15827,N_14708,N_14421);
or U15828 (N_15828,N_14212,N_14296);
and U15829 (N_15829,N_14532,N_14023);
nor U15830 (N_15830,N_14720,N_14657);
and U15831 (N_15831,N_14426,N_14229);
nand U15832 (N_15832,N_14810,N_14716);
nand U15833 (N_15833,N_14591,N_14480);
and U15834 (N_15834,N_14739,N_14889);
or U15835 (N_15835,N_14243,N_14508);
xnor U15836 (N_15836,N_14419,N_14580);
or U15837 (N_15837,N_14919,N_14809);
or U15838 (N_15838,N_14764,N_14521);
and U15839 (N_15839,N_14532,N_14389);
xnor U15840 (N_15840,N_14784,N_14584);
xor U15841 (N_15841,N_14027,N_14283);
nor U15842 (N_15842,N_14560,N_14189);
nand U15843 (N_15843,N_14731,N_14328);
nand U15844 (N_15844,N_14951,N_14196);
and U15845 (N_15845,N_14351,N_14411);
nor U15846 (N_15846,N_14621,N_14605);
nand U15847 (N_15847,N_14511,N_14861);
nand U15848 (N_15848,N_14750,N_14022);
nor U15849 (N_15849,N_14052,N_14094);
nor U15850 (N_15850,N_14176,N_14401);
nand U15851 (N_15851,N_14837,N_14637);
nand U15852 (N_15852,N_14009,N_14465);
nor U15853 (N_15853,N_14885,N_14123);
and U15854 (N_15854,N_14472,N_14695);
nor U15855 (N_15855,N_14032,N_14161);
nand U15856 (N_15856,N_14471,N_14596);
nand U15857 (N_15857,N_14273,N_14798);
or U15858 (N_15858,N_14463,N_14887);
nor U15859 (N_15859,N_14748,N_14865);
xnor U15860 (N_15860,N_14488,N_14662);
or U15861 (N_15861,N_14677,N_14775);
nand U15862 (N_15862,N_14318,N_14159);
xnor U15863 (N_15863,N_14841,N_14212);
nand U15864 (N_15864,N_14150,N_14961);
nand U15865 (N_15865,N_14528,N_14836);
and U15866 (N_15866,N_14863,N_14636);
or U15867 (N_15867,N_14725,N_14793);
and U15868 (N_15868,N_14466,N_14097);
and U15869 (N_15869,N_14299,N_14562);
nand U15870 (N_15870,N_14187,N_14175);
and U15871 (N_15871,N_14814,N_14440);
nor U15872 (N_15872,N_14543,N_14793);
or U15873 (N_15873,N_14926,N_14854);
and U15874 (N_15874,N_14093,N_14507);
nor U15875 (N_15875,N_14183,N_14924);
nand U15876 (N_15876,N_14107,N_14289);
and U15877 (N_15877,N_14126,N_14945);
or U15878 (N_15878,N_14114,N_14547);
xor U15879 (N_15879,N_14205,N_14333);
and U15880 (N_15880,N_14826,N_14665);
or U15881 (N_15881,N_14727,N_14151);
or U15882 (N_15882,N_14184,N_14858);
nand U15883 (N_15883,N_14899,N_14221);
and U15884 (N_15884,N_14969,N_14170);
or U15885 (N_15885,N_14348,N_14043);
nand U15886 (N_15886,N_14781,N_14902);
and U15887 (N_15887,N_14050,N_14151);
nand U15888 (N_15888,N_14468,N_14143);
or U15889 (N_15889,N_14794,N_14698);
or U15890 (N_15890,N_14628,N_14106);
xnor U15891 (N_15891,N_14085,N_14672);
xor U15892 (N_15892,N_14866,N_14318);
nand U15893 (N_15893,N_14515,N_14410);
xor U15894 (N_15894,N_14327,N_14446);
nor U15895 (N_15895,N_14695,N_14942);
nand U15896 (N_15896,N_14182,N_14885);
nand U15897 (N_15897,N_14470,N_14447);
nand U15898 (N_15898,N_14641,N_14113);
nor U15899 (N_15899,N_14709,N_14500);
or U15900 (N_15900,N_14821,N_14894);
or U15901 (N_15901,N_14065,N_14178);
nor U15902 (N_15902,N_14447,N_14546);
or U15903 (N_15903,N_14429,N_14750);
and U15904 (N_15904,N_14084,N_14709);
and U15905 (N_15905,N_14130,N_14666);
nand U15906 (N_15906,N_14907,N_14077);
or U15907 (N_15907,N_14823,N_14275);
nor U15908 (N_15908,N_14422,N_14578);
and U15909 (N_15909,N_14622,N_14294);
nand U15910 (N_15910,N_14369,N_14263);
xor U15911 (N_15911,N_14806,N_14429);
and U15912 (N_15912,N_14637,N_14840);
and U15913 (N_15913,N_14461,N_14106);
nor U15914 (N_15914,N_14529,N_14994);
and U15915 (N_15915,N_14849,N_14261);
nor U15916 (N_15916,N_14487,N_14399);
nor U15917 (N_15917,N_14799,N_14203);
or U15918 (N_15918,N_14162,N_14513);
nor U15919 (N_15919,N_14953,N_14290);
xnor U15920 (N_15920,N_14525,N_14302);
or U15921 (N_15921,N_14594,N_14068);
or U15922 (N_15922,N_14517,N_14641);
nor U15923 (N_15923,N_14425,N_14284);
xnor U15924 (N_15924,N_14011,N_14946);
and U15925 (N_15925,N_14954,N_14575);
and U15926 (N_15926,N_14004,N_14164);
nor U15927 (N_15927,N_14554,N_14151);
and U15928 (N_15928,N_14028,N_14782);
xnor U15929 (N_15929,N_14666,N_14132);
or U15930 (N_15930,N_14956,N_14925);
nor U15931 (N_15931,N_14475,N_14817);
nor U15932 (N_15932,N_14684,N_14219);
nand U15933 (N_15933,N_14719,N_14705);
nor U15934 (N_15934,N_14874,N_14949);
or U15935 (N_15935,N_14567,N_14200);
and U15936 (N_15936,N_14382,N_14786);
xor U15937 (N_15937,N_14942,N_14334);
nor U15938 (N_15938,N_14386,N_14083);
and U15939 (N_15939,N_14815,N_14458);
or U15940 (N_15940,N_14916,N_14077);
or U15941 (N_15941,N_14517,N_14196);
and U15942 (N_15942,N_14439,N_14062);
xnor U15943 (N_15943,N_14713,N_14843);
xnor U15944 (N_15944,N_14119,N_14591);
nand U15945 (N_15945,N_14481,N_14324);
and U15946 (N_15946,N_14455,N_14733);
nor U15947 (N_15947,N_14283,N_14025);
or U15948 (N_15948,N_14817,N_14824);
and U15949 (N_15949,N_14237,N_14040);
and U15950 (N_15950,N_14645,N_14011);
nor U15951 (N_15951,N_14122,N_14793);
xor U15952 (N_15952,N_14376,N_14685);
xnor U15953 (N_15953,N_14034,N_14808);
nor U15954 (N_15954,N_14735,N_14167);
nand U15955 (N_15955,N_14259,N_14159);
or U15956 (N_15956,N_14804,N_14899);
and U15957 (N_15957,N_14418,N_14723);
nor U15958 (N_15958,N_14377,N_14118);
xnor U15959 (N_15959,N_14615,N_14513);
nand U15960 (N_15960,N_14764,N_14255);
and U15961 (N_15961,N_14540,N_14841);
nand U15962 (N_15962,N_14416,N_14912);
xnor U15963 (N_15963,N_14478,N_14132);
and U15964 (N_15964,N_14045,N_14608);
or U15965 (N_15965,N_14560,N_14995);
xor U15966 (N_15966,N_14895,N_14842);
xor U15967 (N_15967,N_14135,N_14979);
xnor U15968 (N_15968,N_14036,N_14830);
or U15969 (N_15969,N_14444,N_14552);
nand U15970 (N_15970,N_14596,N_14609);
xnor U15971 (N_15971,N_14530,N_14841);
nand U15972 (N_15972,N_14410,N_14371);
and U15973 (N_15973,N_14737,N_14732);
nand U15974 (N_15974,N_14794,N_14714);
nand U15975 (N_15975,N_14493,N_14894);
nand U15976 (N_15976,N_14834,N_14966);
nand U15977 (N_15977,N_14194,N_14789);
xnor U15978 (N_15978,N_14978,N_14348);
nand U15979 (N_15979,N_14452,N_14281);
and U15980 (N_15980,N_14952,N_14075);
nor U15981 (N_15981,N_14519,N_14345);
or U15982 (N_15982,N_14761,N_14388);
or U15983 (N_15983,N_14239,N_14223);
or U15984 (N_15984,N_14612,N_14546);
xor U15985 (N_15985,N_14272,N_14344);
or U15986 (N_15986,N_14254,N_14886);
or U15987 (N_15987,N_14453,N_14321);
or U15988 (N_15988,N_14019,N_14499);
nor U15989 (N_15989,N_14986,N_14497);
nand U15990 (N_15990,N_14755,N_14616);
nand U15991 (N_15991,N_14872,N_14384);
xnor U15992 (N_15992,N_14895,N_14965);
nor U15993 (N_15993,N_14690,N_14339);
or U15994 (N_15994,N_14579,N_14176);
or U15995 (N_15995,N_14754,N_14063);
and U15996 (N_15996,N_14802,N_14427);
or U15997 (N_15997,N_14440,N_14462);
nand U15998 (N_15998,N_14723,N_14023);
xor U15999 (N_15999,N_14324,N_14485);
or U16000 (N_16000,N_15378,N_15639);
nor U16001 (N_16001,N_15573,N_15039);
nor U16002 (N_16002,N_15389,N_15477);
nor U16003 (N_16003,N_15607,N_15559);
nand U16004 (N_16004,N_15671,N_15269);
and U16005 (N_16005,N_15251,N_15244);
nor U16006 (N_16006,N_15513,N_15261);
and U16007 (N_16007,N_15098,N_15268);
xor U16008 (N_16008,N_15318,N_15439);
nor U16009 (N_16009,N_15015,N_15434);
nor U16010 (N_16010,N_15081,N_15887);
nand U16011 (N_16011,N_15515,N_15694);
and U16012 (N_16012,N_15067,N_15606);
xnor U16013 (N_16013,N_15262,N_15721);
nor U16014 (N_16014,N_15171,N_15294);
or U16015 (N_16015,N_15023,N_15846);
xnor U16016 (N_16016,N_15528,N_15463);
xor U16017 (N_16017,N_15824,N_15665);
nand U16018 (N_16018,N_15502,N_15973);
or U16019 (N_16019,N_15919,N_15172);
and U16020 (N_16020,N_15494,N_15614);
or U16021 (N_16021,N_15759,N_15806);
nand U16022 (N_16022,N_15041,N_15022);
xnor U16023 (N_16023,N_15282,N_15427);
nand U16024 (N_16024,N_15977,N_15140);
and U16025 (N_16025,N_15619,N_15769);
and U16026 (N_16026,N_15801,N_15475);
nor U16027 (N_16027,N_15110,N_15873);
nand U16028 (N_16028,N_15672,N_15828);
nand U16029 (N_16029,N_15643,N_15382);
nand U16030 (N_16030,N_15926,N_15401);
and U16031 (N_16031,N_15895,N_15629);
xnor U16032 (N_16032,N_15101,N_15001);
or U16033 (N_16033,N_15615,N_15490);
or U16034 (N_16034,N_15877,N_15960);
or U16035 (N_16035,N_15538,N_15812);
nor U16036 (N_16036,N_15542,N_15498);
xnor U16037 (N_16037,N_15603,N_15831);
xnor U16038 (N_16038,N_15307,N_15979);
nor U16039 (N_16039,N_15184,N_15805);
nand U16040 (N_16040,N_15596,N_15419);
or U16041 (N_16041,N_15600,N_15178);
and U16042 (N_16042,N_15305,N_15563);
or U16043 (N_16043,N_15435,N_15106);
nor U16044 (N_16044,N_15837,N_15962);
and U16045 (N_16045,N_15117,N_15774);
nor U16046 (N_16046,N_15526,N_15739);
xor U16047 (N_16047,N_15154,N_15925);
xnor U16048 (N_16048,N_15815,N_15552);
xor U16049 (N_16049,N_15814,N_15767);
nand U16050 (N_16050,N_15851,N_15618);
nand U16051 (N_16051,N_15511,N_15737);
and U16052 (N_16052,N_15093,N_15544);
and U16053 (N_16053,N_15817,N_15776);
nand U16054 (N_16054,N_15113,N_15756);
xnor U16055 (N_16055,N_15062,N_15592);
or U16056 (N_16056,N_15821,N_15488);
or U16057 (N_16057,N_15397,N_15912);
and U16058 (N_16058,N_15866,N_15219);
xor U16059 (N_16059,N_15902,N_15599);
nand U16060 (N_16060,N_15228,N_15561);
xnor U16061 (N_16061,N_15601,N_15345);
nor U16062 (N_16062,N_15868,N_15373);
nand U16063 (N_16063,N_15211,N_15365);
xnor U16064 (N_16064,N_15743,N_15313);
or U16065 (N_16065,N_15857,N_15679);
nor U16066 (N_16066,N_15414,N_15223);
or U16067 (N_16067,N_15638,N_15928);
nor U16068 (N_16068,N_15405,N_15809);
nand U16069 (N_16069,N_15421,N_15204);
nor U16070 (N_16070,N_15578,N_15650);
nor U16071 (N_16071,N_15316,N_15705);
or U16072 (N_16072,N_15451,N_15342);
or U16073 (N_16073,N_15509,N_15764);
nand U16074 (N_16074,N_15186,N_15945);
nor U16075 (N_16075,N_15403,N_15630);
nor U16076 (N_16076,N_15433,N_15715);
nand U16077 (N_16077,N_15042,N_15727);
nor U16078 (N_16078,N_15275,N_15392);
nor U16079 (N_16079,N_15400,N_15384);
nor U16080 (N_16080,N_15602,N_15330);
nand U16081 (N_16081,N_15850,N_15840);
xor U16082 (N_16082,N_15280,N_15930);
nor U16083 (N_16083,N_15843,N_15900);
xnor U16084 (N_16084,N_15044,N_15982);
nor U16085 (N_16085,N_15816,N_15899);
or U16086 (N_16086,N_15700,N_15993);
nand U16087 (N_16087,N_15966,N_15872);
and U16088 (N_16088,N_15339,N_15864);
or U16089 (N_16089,N_15888,N_15369);
nand U16090 (N_16090,N_15297,N_15447);
xor U16091 (N_16091,N_15683,N_15792);
nand U16092 (N_16092,N_15119,N_15548);
or U16093 (N_16093,N_15018,N_15445);
or U16094 (N_16094,N_15108,N_15353);
nand U16095 (N_16095,N_15356,N_15380);
and U16096 (N_16096,N_15901,N_15331);
nor U16097 (N_16097,N_15111,N_15628);
nand U16098 (N_16098,N_15319,N_15835);
or U16099 (N_16099,N_15968,N_15415);
nor U16100 (N_16100,N_15860,N_15971);
nand U16101 (N_16101,N_15489,N_15613);
nand U16102 (N_16102,N_15781,N_15728);
xnor U16103 (N_16103,N_15685,N_15554);
nand U16104 (N_16104,N_15799,N_15916);
or U16105 (N_16105,N_15123,N_15917);
nand U16106 (N_16106,N_15684,N_15051);
nand U16107 (N_16107,N_15571,N_15078);
and U16108 (N_16108,N_15758,N_15121);
and U16109 (N_16109,N_15362,N_15163);
nand U16110 (N_16110,N_15190,N_15141);
and U16111 (N_16111,N_15351,N_15139);
and U16112 (N_16112,N_15243,N_15393);
nand U16113 (N_16113,N_15045,N_15161);
nand U16114 (N_16114,N_15304,N_15744);
and U16115 (N_16115,N_15506,N_15149);
or U16116 (N_16116,N_15826,N_15545);
nand U16117 (N_16117,N_15976,N_15355);
and U16118 (N_16118,N_15696,N_15398);
or U16119 (N_16119,N_15852,N_15048);
nor U16120 (N_16120,N_15151,N_15867);
or U16121 (N_16121,N_15882,N_15595);
nor U16122 (N_16122,N_15795,N_15199);
nand U16123 (N_16123,N_15220,N_15550);
nor U16124 (N_16124,N_15751,N_15712);
or U16125 (N_16125,N_15274,N_15802);
nor U16126 (N_16126,N_15742,N_15390);
and U16127 (N_16127,N_15474,N_15660);
and U16128 (N_16128,N_15593,N_15453);
xnor U16129 (N_16129,N_15138,N_15749);
nand U16130 (N_16130,N_15049,N_15931);
nand U16131 (N_16131,N_15730,N_15693);
or U16132 (N_16132,N_15541,N_15181);
nor U16133 (N_16133,N_15366,N_15647);
and U16134 (N_16134,N_15168,N_15670);
and U16135 (N_16135,N_15485,N_15621);
xnor U16136 (N_16136,N_15567,N_15127);
and U16137 (N_16137,N_15818,N_15037);
xnor U16138 (N_16138,N_15009,N_15587);
nor U16139 (N_16139,N_15033,N_15285);
or U16140 (N_16140,N_15103,N_15478);
xor U16141 (N_16141,N_15950,N_15272);
or U16142 (N_16142,N_15320,N_15296);
nor U16143 (N_16143,N_15247,N_15310);
nand U16144 (N_16144,N_15649,N_15423);
nor U16145 (N_16145,N_15317,N_15132);
nand U16146 (N_16146,N_15420,N_15745);
nor U16147 (N_16147,N_15777,N_15845);
nand U16148 (N_16148,N_15890,N_15590);
and U16149 (N_16149,N_15214,N_15855);
xnor U16150 (N_16150,N_15825,N_15978);
xnor U16151 (N_16151,N_15589,N_15061);
xnor U16152 (N_16152,N_15703,N_15609);
nand U16153 (N_16153,N_15079,N_15134);
xor U16154 (N_16154,N_15175,N_15077);
and U16155 (N_16155,N_15543,N_15284);
nor U16156 (N_16156,N_15517,N_15129);
and U16157 (N_16157,N_15784,N_15412);
nand U16158 (N_16158,N_15765,N_15233);
nand U16159 (N_16159,N_15681,N_15100);
and U16160 (N_16160,N_15271,N_15135);
nand U16161 (N_16161,N_15063,N_15834);
and U16162 (N_16162,N_15669,N_15344);
nand U16163 (N_16163,N_15236,N_15540);
nor U16164 (N_16164,N_15519,N_15143);
nor U16165 (N_16165,N_15066,N_15258);
nand U16166 (N_16166,N_15510,N_15725);
nand U16167 (N_16167,N_15856,N_15499);
and U16168 (N_16168,N_15859,N_15588);
nand U16169 (N_16169,N_15952,N_15634);
nor U16170 (N_16170,N_15794,N_15698);
or U16171 (N_16171,N_15457,N_15796);
nor U16172 (N_16172,N_15381,N_15597);
or U16173 (N_16173,N_15975,N_15229);
or U16174 (N_16174,N_15025,N_15476);
xor U16175 (N_16175,N_15640,N_15083);
and U16176 (N_16176,N_15341,N_15565);
nor U16177 (N_16177,N_15723,N_15898);
nand U16178 (N_16178,N_15455,N_15118);
xor U16179 (N_16179,N_15833,N_15354);
and U16180 (N_16180,N_15883,N_15273);
and U16181 (N_16181,N_15438,N_15880);
xnor U16182 (N_16182,N_15653,N_15052);
nand U16183 (N_16183,N_15946,N_15906);
or U16184 (N_16184,N_15689,N_15753);
xor U16185 (N_16185,N_15686,N_15459);
nor U16186 (N_16186,N_15065,N_15594);
or U16187 (N_16187,N_15343,N_15377);
and U16188 (N_16188,N_15636,N_15935);
and U16189 (N_16189,N_15335,N_15006);
nand U16190 (N_16190,N_15820,N_15875);
nor U16191 (N_16191,N_15329,N_15804);
or U16192 (N_16192,N_15185,N_15326);
xnor U16193 (N_16193,N_15626,N_15667);
or U16194 (N_16194,N_15608,N_15980);
and U16195 (N_16195,N_15688,N_15003);
or U16196 (N_16196,N_15525,N_15292);
nor U16197 (N_16197,N_15965,N_15800);
nor U16198 (N_16198,N_15413,N_15738);
or U16199 (N_16199,N_15183,N_15162);
or U16200 (N_16200,N_15361,N_15673);
and U16201 (N_16201,N_15974,N_15286);
nor U16202 (N_16202,N_15075,N_15446);
and U16203 (N_16203,N_15972,N_15215);
or U16204 (N_16204,N_15735,N_15270);
nand U16205 (N_16205,N_15617,N_15921);
xnor U16206 (N_16206,N_15652,N_15203);
or U16207 (N_16207,N_15658,N_15238);
or U16208 (N_16208,N_15907,N_15002);
nor U16209 (N_16209,N_15610,N_15512);
or U16210 (N_16210,N_15748,N_15473);
or U16211 (N_16211,N_15555,N_15762);
or U16212 (N_16212,N_15924,N_15763);
nor U16213 (N_16213,N_15131,N_15216);
nor U16214 (N_16214,N_15625,N_15704);
or U16215 (N_16215,N_15169,N_15778);
xnor U16216 (N_16216,N_15417,N_15126);
and U16217 (N_16217,N_15089,N_15922);
or U16218 (N_16218,N_15470,N_15249);
or U16219 (N_16219,N_15456,N_15325);
xnor U16220 (N_16220,N_15699,N_15441);
nor U16221 (N_16221,N_15583,N_15133);
or U16222 (N_16222,N_15201,N_15056);
xnor U16223 (N_16223,N_15182,N_15224);
nor U16224 (N_16224,N_15449,N_15871);
or U16225 (N_16225,N_15808,N_15388);
and U16226 (N_16226,N_15232,N_15291);
nand U16227 (N_16227,N_15616,N_15073);
or U16228 (N_16228,N_15213,N_15797);
nor U16229 (N_16229,N_15987,N_15469);
nand U16230 (N_16230,N_15349,N_15150);
or U16231 (N_16231,N_15556,N_15740);
nand U16232 (N_16232,N_15532,N_15363);
nand U16233 (N_16233,N_15411,N_15237);
and U16234 (N_16234,N_15787,N_15088);
nand U16235 (N_16235,N_15722,N_15920);
nand U16236 (N_16236,N_15299,N_15208);
nand U16237 (N_16237,N_15357,N_15605);
or U16238 (N_16238,N_15893,N_15881);
or U16239 (N_16239,N_15364,N_15265);
nand U16240 (N_16240,N_15306,N_15430);
nor U16241 (N_16241,N_15841,N_15690);
xnor U16242 (N_16242,N_15995,N_15482);
xor U16243 (N_16243,N_15053,N_15050);
or U16244 (N_16244,N_15012,N_15496);
nor U16245 (N_16245,N_15137,N_15927);
nor U16246 (N_16246,N_15210,N_15255);
and U16247 (N_16247,N_15340,N_15192);
nand U16248 (N_16248,N_15557,N_15783);
and U16249 (N_16249,N_15788,N_15252);
nand U16250 (N_16250,N_15963,N_15848);
nand U16251 (N_16251,N_15295,N_15189);
xor U16252 (N_16252,N_15507,N_15897);
or U16253 (N_16253,N_15454,N_15155);
or U16254 (N_16254,N_15315,N_15218);
and U16255 (N_16255,N_15716,N_15779);
and U16256 (N_16256,N_15004,N_15071);
nand U16257 (N_16257,N_15207,N_15682);
and U16258 (N_16258,N_15308,N_15662);
or U16259 (N_16259,N_15558,N_15998);
xor U16260 (N_16260,N_15472,N_15539);
nor U16261 (N_16261,N_15082,N_15575);
nor U16262 (N_16262,N_15124,N_15905);
xor U16263 (N_16263,N_15598,N_15337);
and U16264 (N_16264,N_15780,N_15941);
or U16265 (N_16265,N_15947,N_15157);
nor U16266 (N_16266,N_15409,N_15577);
or U16267 (N_16267,N_15957,N_15152);
nor U16268 (N_16268,N_15448,N_15109);
xnor U16269 (N_16269,N_15142,N_15572);
and U16270 (N_16270,N_15064,N_15120);
nand U16271 (N_16271,N_15144,N_15352);
nand U16272 (N_16272,N_15279,N_15560);
or U16273 (N_16273,N_15300,N_15462);
and U16274 (N_16274,N_15766,N_15505);
nand U16275 (N_16275,N_15115,N_15706);
xnor U16276 (N_16276,N_15654,N_15503);
or U16277 (N_16277,N_15146,N_15633);
nand U16278 (N_16278,N_15964,N_15536);
nor U16279 (N_16279,N_15466,N_15032);
or U16280 (N_16280,N_15399,N_15914);
nor U16281 (N_16281,N_15695,N_15309);
nand U16282 (N_16282,N_15027,N_15677);
xor U16283 (N_16283,N_15368,N_15458);
and U16284 (N_16284,N_15508,N_15180);
nor U16285 (N_16285,N_15070,N_15711);
and U16286 (N_16286,N_15933,N_15076);
or U16287 (N_16287,N_15226,N_15798);
and U16288 (N_16288,N_15311,N_15239);
and U16289 (N_16289,N_15253,N_15293);
nand U16290 (N_16290,N_15394,N_15426);
nor U16291 (N_16291,N_15418,N_15813);
nand U16292 (N_16292,N_15580,N_15334);
or U16293 (N_16293,N_15198,N_15655);
or U16294 (N_16294,N_15884,N_15529);
nand U16295 (N_16295,N_15495,N_15819);
or U16296 (N_16296,N_15358,N_15122);
xnor U16297 (N_16297,N_15534,N_15301);
xnor U16298 (N_16298,N_15896,N_15581);
xnor U16299 (N_16299,N_15011,N_15627);
xnor U16300 (N_16300,N_15114,N_15624);
nor U16301 (N_16301,N_15659,N_15954);
and U16302 (N_16302,N_15811,N_15046);
and U16303 (N_16303,N_15775,N_15836);
xnor U16304 (N_16304,N_15990,N_15460);
nand U16305 (N_16305,N_15604,N_15350);
or U16306 (N_16306,N_15153,N_15793);
or U16307 (N_16307,N_15328,N_15029);
and U16308 (N_16308,N_15112,N_15170);
and U16309 (N_16309,N_15464,N_15520);
xor U16310 (N_16310,N_15323,N_15225);
and U16311 (N_16311,N_15096,N_15918);
and U16312 (N_16312,N_15188,N_15648);
or U16313 (N_16313,N_15631,N_15091);
or U16314 (N_16314,N_15092,N_15217);
xnor U16315 (N_16315,N_15424,N_15068);
nand U16316 (N_16316,N_15549,N_15790);
nor U16317 (N_16317,N_15371,N_15010);
xnor U16318 (N_16318,N_15407,N_15314);
or U16319 (N_16319,N_15611,N_15383);
and U16320 (N_16320,N_15518,N_15145);
and U16321 (N_16321,N_15522,N_15984);
or U16322 (N_16322,N_15017,N_15030);
xor U16323 (N_16323,N_15467,N_15870);
nor U16324 (N_16324,N_15264,N_15200);
xor U16325 (N_16325,N_15854,N_15564);
xor U16326 (N_16326,N_15641,N_15047);
and U16327 (N_16327,N_15791,N_15431);
xnor U16328 (N_16328,N_15360,N_15886);
xor U16329 (N_16329,N_15632,N_15692);
and U16330 (N_16330,N_15989,N_15359);
or U16331 (N_16331,N_15988,N_15026);
or U16332 (N_16332,N_15375,N_15234);
and U16333 (N_16333,N_15007,N_15322);
nor U16334 (N_16334,N_15165,N_15736);
or U16335 (N_16335,N_15090,N_15332);
nor U16336 (N_16336,N_15250,N_15347);
nand U16337 (N_16337,N_15194,N_15789);
nor U16338 (N_16338,N_15701,N_15934);
nor U16339 (N_16339,N_15746,N_15158);
xnor U16340 (N_16340,N_15391,N_15955);
and U16341 (N_16341,N_15102,N_15830);
or U16342 (N_16342,N_15923,N_15497);
nand U16343 (N_16343,N_15635,N_15034);
xor U16344 (N_16344,N_15038,N_15105);
or U16345 (N_16345,N_15031,N_15387);
or U16346 (N_16346,N_15060,N_15442);
and U16347 (N_16347,N_15773,N_15094);
nand U16348 (N_16348,N_15084,N_15014);
nor U16349 (N_16349,N_15338,N_15174);
nor U16350 (N_16350,N_15085,N_15942);
nand U16351 (N_16351,N_15099,N_15013);
and U16352 (N_16352,N_15770,N_15125);
or U16353 (N_16353,N_15847,N_15346);
or U16354 (N_16354,N_15348,N_15479);
or U16355 (N_16355,N_15107,N_15491);
nor U16356 (N_16356,N_15678,N_15983);
xor U16357 (N_16357,N_15932,N_15087);
nor U16358 (N_16358,N_15404,N_15254);
and U16359 (N_16359,N_15147,N_15747);
nor U16360 (N_16360,N_15668,N_15493);
nand U16361 (N_16361,N_15680,N_15288);
xor U16362 (N_16362,N_15687,N_15876);
and U16363 (N_16363,N_15863,N_15374);
xor U16364 (N_16364,N_15651,N_15862);
nand U16365 (N_16365,N_15710,N_15786);
nor U16366 (N_16366,N_15771,N_15005);
xor U16367 (N_16367,N_15524,N_15043);
nand U16368 (N_16368,N_15324,N_15527);
xor U16369 (N_16369,N_15750,N_15177);
or U16370 (N_16370,N_15757,N_15533);
xnor U16371 (N_16371,N_15230,N_15241);
xnor U16372 (N_16372,N_15246,N_15436);
nor U16373 (N_16373,N_15879,N_15953);
nand U16374 (N_16374,N_15958,N_15656);
nand U16375 (N_16375,N_15996,N_15336);
xnor U16376 (N_16376,N_15432,N_15376);
and U16377 (N_16377,N_15810,N_15481);
and U16378 (N_16378,N_15967,N_15657);
xnor U16379 (N_16379,N_15637,N_15839);
or U16380 (N_16380,N_15385,N_15807);
or U16381 (N_16381,N_15231,N_15205);
or U16382 (N_16382,N_15874,N_15903);
or U16383 (N_16383,N_15553,N_15136);
nand U16384 (N_16384,N_15734,N_15281);
nor U16385 (N_16385,N_15256,N_15167);
xor U16386 (N_16386,N_15991,N_15531);
xor U16387 (N_16387,N_15909,N_15842);
or U16388 (N_16388,N_15622,N_15944);
nand U16389 (N_16389,N_15720,N_15303);
or U16390 (N_16390,N_15772,N_15222);
or U16391 (N_16391,N_15838,N_15724);
nand U16392 (N_16392,N_15915,N_15731);
nand U16393 (N_16393,N_15913,N_15530);
nor U16394 (N_16394,N_15019,N_15410);
or U16395 (N_16395,N_15719,N_15097);
xor U16396 (N_16396,N_15970,N_15452);
nor U16397 (N_16397,N_15104,N_15212);
nand U16398 (N_16398,N_15242,N_15487);
xnor U16399 (N_16399,N_15267,N_15869);
nand U16400 (N_16400,N_15058,N_15196);
or U16401 (N_16401,N_15501,N_15537);
or U16402 (N_16402,N_15861,N_15500);
and U16403 (N_16403,N_15729,N_15904);
and U16404 (N_16404,N_15666,N_15803);
nor U16405 (N_16405,N_15733,N_15760);
and U16406 (N_16406,N_15853,N_15259);
nor U16407 (N_16407,N_15504,N_15785);
nor U16408 (N_16408,N_15202,N_15367);
and U16409 (N_16409,N_15889,N_15663);
or U16410 (N_16410,N_15761,N_15021);
and U16411 (N_16411,N_15028,N_15483);
nor U16412 (N_16412,N_15675,N_15072);
nand U16413 (N_16413,N_15159,N_15823);
nand U16414 (N_16414,N_15197,N_15276);
nor U16415 (N_16415,N_15492,N_15484);
and U16416 (N_16416,N_15885,N_15570);
and U16417 (N_16417,N_15298,N_15969);
and U16418 (N_16418,N_15372,N_15891);
nand U16419 (N_16419,N_15849,N_15406);
nand U16420 (N_16420,N_15908,N_15176);
xnor U16421 (N_16421,N_15148,N_15844);
or U16422 (N_16422,N_15546,N_15386);
xor U16423 (N_16423,N_15095,N_15471);
nor U16424 (N_16424,N_15646,N_15961);
nand U16425 (N_16425,N_15156,N_15187);
and U16426 (N_16426,N_15959,N_15951);
xnor U16427 (N_16427,N_15260,N_15582);
or U16428 (N_16428,N_15985,N_15894);
nor U16429 (N_16429,N_15266,N_15576);
nand U16430 (N_16430,N_15086,N_15016);
nand U16431 (N_16431,N_15302,N_15257);
nand U16432 (N_16432,N_15832,N_15206);
and U16433 (N_16433,N_15160,N_15221);
xnor U16434 (N_16434,N_15547,N_15055);
or U16435 (N_16435,N_15691,N_15911);
nor U16436 (N_16436,N_15523,N_15128);
nand U16437 (N_16437,N_15248,N_15191);
or U16438 (N_16438,N_15562,N_15069);
nor U16439 (N_16439,N_15535,N_15579);
and U16440 (N_16440,N_15752,N_15948);
nor U16441 (N_16441,N_15910,N_15321);
nor U16442 (N_16442,N_15878,N_15986);
or U16443 (N_16443,N_15584,N_15283);
nor U16444 (N_16444,N_15591,N_15620);
xnor U16445 (N_16445,N_15024,N_15726);
xor U16446 (N_16446,N_15713,N_15179);
or U16447 (N_16447,N_15702,N_15707);
and U16448 (N_16448,N_15644,N_15929);
xnor U16449 (N_16449,N_15057,N_15054);
nand U16450 (N_16450,N_15661,N_15676);
or U16451 (N_16451,N_15568,N_15674);
xor U16452 (N_16452,N_15195,N_15829);
xnor U16453 (N_16453,N_15235,N_15664);
nand U16454 (N_16454,N_15949,N_15566);
nand U16455 (N_16455,N_15858,N_15333);
nand U16456 (N_16456,N_15395,N_15645);
and U16457 (N_16457,N_15612,N_15465);
or U16458 (N_16458,N_15379,N_15697);
nand U16459 (N_16459,N_15516,N_15939);
xnor U16460 (N_16460,N_15059,N_15289);
or U16461 (N_16461,N_15440,N_15396);
nor U16462 (N_16462,N_15402,N_15754);
nor U16463 (N_16463,N_15623,N_15450);
or U16464 (N_16464,N_15585,N_15938);
xnor U16465 (N_16465,N_15994,N_15782);
or U16466 (N_16466,N_15461,N_15040);
nand U16467 (N_16467,N_15822,N_15768);
or U16468 (N_16468,N_15408,N_15997);
xor U16469 (N_16469,N_15290,N_15444);
and U16470 (N_16470,N_15940,N_15551);
nor U16471 (N_16471,N_15327,N_15443);
or U16472 (N_16472,N_15020,N_15209);
or U16473 (N_16473,N_15429,N_15569);
or U16474 (N_16474,N_15263,N_15116);
nand U16475 (N_16475,N_15865,N_15416);
xor U16476 (N_16476,N_15036,N_15008);
nor U16477 (N_16477,N_15717,N_15173);
nor U16478 (N_16478,N_15370,N_15936);
or U16479 (N_16479,N_15827,N_15287);
and U16480 (N_16480,N_15240,N_15278);
nor U16481 (N_16481,N_15193,N_15166);
nand U16482 (N_16482,N_15732,N_15718);
or U16483 (N_16483,N_15468,N_15708);
nor U16484 (N_16484,N_15164,N_15755);
nand U16485 (N_16485,N_15312,N_15574);
xnor U16486 (N_16486,N_15514,N_15709);
nand U16487 (N_16487,N_15130,N_15943);
nand U16488 (N_16488,N_15245,N_15480);
or U16489 (N_16489,N_15642,N_15956);
nand U16490 (N_16490,N_15422,N_15937);
and U16491 (N_16491,N_15277,N_15074);
and U16492 (N_16492,N_15521,N_15486);
xor U16493 (N_16493,N_15437,N_15035);
and U16494 (N_16494,N_15428,N_15892);
and U16495 (N_16495,N_15586,N_15080);
nand U16496 (N_16496,N_15425,N_15981);
xnor U16497 (N_16497,N_15992,N_15227);
or U16498 (N_16498,N_15741,N_15714);
nand U16499 (N_16499,N_15999,N_15000);
and U16500 (N_16500,N_15370,N_15192);
or U16501 (N_16501,N_15738,N_15417);
or U16502 (N_16502,N_15619,N_15268);
or U16503 (N_16503,N_15943,N_15568);
nor U16504 (N_16504,N_15884,N_15994);
nand U16505 (N_16505,N_15210,N_15291);
or U16506 (N_16506,N_15780,N_15440);
and U16507 (N_16507,N_15258,N_15182);
or U16508 (N_16508,N_15877,N_15130);
nand U16509 (N_16509,N_15787,N_15210);
or U16510 (N_16510,N_15164,N_15050);
xor U16511 (N_16511,N_15911,N_15192);
and U16512 (N_16512,N_15740,N_15944);
nand U16513 (N_16513,N_15342,N_15575);
nor U16514 (N_16514,N_15399,N_15977);
xnor U16515 (N_16515,N_15234,N_15330);
xnor U16516 (N_16516,N_15070,N_15725);
nor U16517 (N_16517,N_15059,N_15106);
nand U16518 (N_16518,N_15198,N_15741);
nand U16519 (N_16519,N_15417,N_15708);
and U16520 (N_16520,N_15178,N_15425);
or U16521 (N_16521,N_15521,N_15100);
nand U16522 (N_16522,N_15295,N_15966);
nor U16523 (N_16523,N_15609,N_15905);
and U16524 (N_16524,N_15580,N_15458);
and U16525 (N_16525,N_15884,N_15499);
and U16526 (N_16526,N_15697,N_15571);
nor U16527 (N_16527,N_15500,N_15444);
and U16528 (N_16528,N_15393,N_15861);
or U16529 (N_16529,N_15031,N_15894);
nor U16530 (N_16530,N_15676,N_15862);
or U16531 (N_16531,N_15507,N_15711);
and U16532 (N_16532,N_15761,N_15784);
and U16533 (N_16533,N_15651,N_15083);
nor U16534 (N_16534,N_15958,N_15942);
and U16535 (N_16535,N_15597,N_15549);
nor U16536 (N_16536,N_15226,N_15428);
nand U16537 (N_16537,N_15661,N_15002);
and U16538 (N_16538,N_15855,N_15832);
nor U16539 (N_16539,N_15446,N_15077);
nor U16540 (N_16540,N_15066,N_15723);
and U16541 (N_16541,N_15331,N_15557);
nor U16542 (N_16542,N_15999,N_15985);
xnor U16543 (N_16543,N_15311,N_15833);
nand U16544 (N_16544,N_15266,N_15320);
nand U16545 (N_16545,N_15929,N_15080);
nand U16546 (N_16546,N_15197,N_15199);
or U16547 (N_16547,N_15459,N_15906);
nor U16548 (N_16548,N_15129,N_15617);
nand U16549 (N_16549,N_15545,N_15862);
xor U16550 (N_16550,N_15305,N_15050);
xor U16551 (N_16551,N_15795,N_15892);
xor U16552 (N_16552,N_15552,N_15565);
and U16553 (N_16553,N_15835,N_15817);
nor U16554 (N_16554,N_15889,N_15787);
xnor U16555 (N_16555,N_15224,N_15143);
nor U16556 (N_16556,N_15380,N_15886);
and U16557 (N_16557,N_15399,N_15687);
nand U16558 (N_16558,N_15051,N_15757);
or U16559 (N_16559,N_15223,N_15623);
nand U16560 (N_16560,N_15571,N_15111);
xor U16561 (N_16561,N_15165,N_15077);
nand U16562 (N_16562,N_15383,N_15350);
xor U16563 (N_16563,N_15076,N_15181);
nand U16564 (N_16564,N_15950,N_15081);
and U16565 (N_16565,N_15871,N_15867);
xor U16566 (N_16566,N_15575,N_15497);
nand U16567 (N_16567,N_15328,N_15379);
or U16568 (N_16568,N_15701,N_15896);
nor U16569 (N_16569,N_15527,N_15432);
nand U16570 (N_16570,N_15816,N_15831);
nor U16571 (N_16571,N_15171,N_15740);
xor U16572 (N_16572,N_15039,N_15964);
or U16573 (N_16573,N_15733,N_15962);
xor U16574 (N_16574,N_15190,N_15248);
and U16575 (N_16575,N_15957,N_15549);
and U16576 (N_16576,N_15597,N_15264);
nor U16577 (N_16577,N_15823,N_15275);
or U16578 (N_16578,N_15241,N_15380);
or U16579 (N_16579,N_15022,N_15584);
or U16580 (N_16580,N_15925,N_15729);
nand U16581 (N_16581,N_15966,N_15864);
or U16582 (N_16582,N_15279,N_15436);
nand U16583 (N_16583,N_15067,N_15906);
xnor U16584 (N_16584,N_15266,N_15406);
nand U16585 (N_16585,N_15029,N_15567);
xnor U16586 (N_16586,N_15970,N_15445);
xnor U16587 (N_16587,N_15190,N_15247);
nand U16588 (N_16588,N_15111,N_15383);
or U16589 (N_16589,N_15321,N_15632);
or U16590 (N_16590,N_15215,N_15848);
xor U16591 (N_16591,N_15387,N_15053);
nand U16592 (N_16592,N_15369,N_15049);
or U16593 (N_16593,N_15813,N_15428);
or U16594 (N_16594,N_15749,N_15772);
nand U16595 (N_16595,N_15415,N_15010);
nor U16596 (N_16596,N_15652,N_15181);
nand U16597 (N_16597,N_15737,N_15256);
nor U16598 (N_16598,N_15743,N_15231);
or U16599 (N_16599,N_15722,N_15148);
or U16600 (N_16600,N_15938,N_15110);
nor U16601 (N_16601,N_15931,N_15668);
nor U16602 (N_16602,N_15467,N_15323);
nand U16603 (N_16603,N_15483,N_15584);
or U16604 (N_16604,N_15023,N_15485);
or U16605 (N_16605,N_15723,N_15984);
and U16606 (N_16606,N_15520,N_15359);
nand U16607 (N_16607,N_15996,N_15573);
and U16608 (N_16608,N_15481,N_15663);
nand U16609 (N_16609,N_15238,N_15096);
and U16610 (N_16610,N_15236,N_15467);
xor U16611 (N_16611,N_15280,N_15981);
xor U16612 (N_16612,N_15384,N_15589);
nor U16613 (N_16613,N_15560,N_15031);
xor U16614 (N_16614,N_15448,N_15278);
xnor U16615 (N_16615,N_15553,N_15429);
or U16616 (N_16616,N_15784,N_15896);
nand U16617 (N_16617,N_15053,N_15463);
or U16618 (N_16618,N_15469,N_15786);
nand U16619 (N_16619,N_15170,N_15818);
and U16620 (N_16620,N_15881,N_15741);
and U16621 (N_16621,N_15145,N_15665);
nand U16622 (N_16622,N_15140,N_15863);
or U16623 (N_16623,N_15521,N_15877);
and U16624 (N_16624,N_15664,N_15519);
nor U16625 (N_16625,N_15919,N_15388);
xnor U16626 (N_16626,N_15786,N_15729);
and U16627 (N_16627,N_15707,N_15544);
xor U16628 (N_16628,N_15844,N_15710);
and U16629 (N_16629,N_15804,N_15201);
nand U16630 (N_16630,N_15599,N_15355);
nor U16631 (N_16631,N_15827,N_15672);
or U16632 (N_16632,N_15021,N_15802);
nor U16633 (N_16633,N_15231,N_15650);
or U16634 (N_16634,N_15953,N_15775);
and U16635 (N_16635,N_15863,N_15174);
or U16636 (N_16636,N_15873,N_15802);
nor U16637 (N_16637,N_15435,N_15256);
or U16638 (N_16638,N_15769,N_15629);
xnor U16639 (N_16639,N_15973,N_15926);
nor U16640 (N_16640,N_15720,N_15277);
nor U16641 (N_16641,N_15632,N_15235);
nor U16642 (N_16642,N_15086,N_15174);
xor U16643 (N_16643,N_15018,N_15325);
or U16644 (N_16644,N_15874,N_15364);
and U16645 (N_16645,N_15961,N_15699);
or U16646 (N_16646,N_15816,N_15448);
nor U16647 (N_16647,N_15304,N_15345);
and U16648 (N_16648,N_15282,N_15701);
nand U16649 (N_16649,N_15629,N_15121);
and U16650 (N_16650,N_15465,N_15301);
nor U16651 (N_16651,N_15248,N_15717);
or U16652 (N_16652,N_15070,N_15937);
nor U16653 (N_16653,N_15614,N_15377);
or U16654 (N_16654,N_15031,N_15377);
xor U16655 (N_16655,N_15633,N_15183);
nand U16656 (N_16656,N_15516,N_15208);
or U16657 (N_16657,N_15633,N_15729);
or U16658 (N_16658,N_15106,N_15489);
nand U16659 (N_16659,N_15039,N_15220);
xor U16660 (N_16660,N_15231,N_15005);
xnor U16661 (N_16661,N_15425,N_15855);
or U16662 (N_16662,N_15327,N_15204);
and U16663 (N_16663,N_15192,N_15094);
xor U16664 (N_16664,N_15980,N_15318);
xor U16665 (N_16665,N_15597,N_15295);
or U16666 (N_16666,N_15770,N_15761);
nor U16667 (N_16667,N_15839,N_15301);
and U16668 (N_16668,N_15330,N_15815);
xor U16669 (N_16669,N_15734,N_15386);
nand U16670 (N_16670,N_15318,N_15153);
nand U16671 (N_16671,N_15243,N_15056);
nand U16672 (N_16672,N_15171,N_15004);
and U16673 (N_16673,N_15092,N_15045);
and U16674 (N_16674,N_15724,N_15082);
and U16675 (N_16675,N_15499,N_15983);
nor U16676 (N_16676,N_15015,N_15356);
nand U16677 (N_16677,N_15495,N_15933);
xor U16678 (N_16678,N_15944,N_15336);
xnor U16679 (N_16679,N_15355,N_15600);
nor U16680 (N_16680,N_15277,N_15003);
nor U16681 (N_16681,N_15277,N_15182);
xor U16682 (N_16682,N_15252,N_15874);
xor U16683 (N_16683,N_15785,N_15253);
nor U16684 (N_16684,N_15524,N_15338);
and U16685 (N_16685,N_15721,N_15813);
and U16686 (N_16686,N_15873,N_15500);
and U16687 (N_16687,N_15839,N_15377);
nor U16688 (N_16688,N_15953,N_15473);
and U16689 (N_16689,N_15411,N_15195);
or U16690 (N_16690,N_15844,N_15838);
and U16691 (N_16691,N_15884,N_15124);
nor U16692 (N_16692,N_15869,N_15799);
nand U16693 (N_16693,N_15030,N_15656);
xnor U16694 (N_16694,N_15916,N_15913);
xnor U16695 (N_16695,N_15556,N_15276);
nor U16696 (N_16696,N_15096,N_15376);
or U16697 (N_16697,N_15559,N_15736);
or U16698 (N_16698,N_15964,N_15556);
nor U16699 (N_16699,N_15010,N_15149);
or U16700 (N_16700,N_15803,N_15962);
or U16701 (N_16701,N_15425,N_15865);
and U16702 (N_16702,N_15532,N_15595);
and U16703 (N_16703,N_15738,N_15586);
nor U16704 (N_16704,N_15679,N_15305);
or U16705 (N_16705,N_15829,N_15594);
or U16706 (N_16706,N_15358,N_15031);
xor U16707 (N_16707,N_15947,N_15720);
nand U16708 (N_16708,N_15862,N_15236);
and U16709 (N_16709,N_15022,N_15580);
or U16710 (N_16710,N_15223,N_15301);
or U16711 (N_16711,N_15780,N_15679);
nand U16712 (N_16712,N_15984,N_15552);
or U16713 (N_16713,N_15432,N_15054);
xnor U16714 (N_16714,N_15995,N_15583);
nand U16715 (N_16715,N_15813,N_15329);
xnor U16716 (N_16716,N_15222,N_15976);
nor U16717 (N_16717,N_15781,N_15908);
or U16718 (N_16718,N_15375,N_15211);
and U16719 (N_16719,N_15543,N_15495);
nand U16720 (N_16720,N_15058,N_15441);
nor U16721 (N_16721,N_15509,N_15280);
and U16722 (N_16722,N_15935,N_15503);
and U16723 (N_16723,N_15129,N_15986);
and U16724 (N_16724,N_15137,N_15834);
nand U16725 (N_16725,N_15649,N_15856);
xor U16726 (N_16726,N_15923,N_15698);
xnor U16727 (N_16727,N_15687,N_15388);
nor U16728 (N_16728,N_15507,N_15964);
and U16729 (N_16729,N_15864,N_15274);
nand U16730 (N_16730,N_15411,N_15397);
and U16731 (N_16731,N_15704,N_15231);
xnor U16732 (N_16732,N_15973,N_15033);
nand U16733 (N_16733,N_15694,N_15180);
or U16734 (N_16734,N_15800,N_15761);
and U16735 (N_16735,N_15741,N_15634);
xor U16736 (N_16736,N_15191,N_15561);
xor U16737 (N_16737,N_15405,N_15042);
and U16738 (N_16738,N_15358,N_15716);
nor U16739 (N_16739,N_15895,N_15213);
or U16740 (N_16740,N_15578,N_15815);
or U16741 (N_16741,N_15674,N_15273);
and U16742 (N_16742,N_15927,N_15598);
or U16743 (N_16743,N_15041,N_15769);
xnor U16744 (N_16744,N_15948,N_15786);
xor U16745 (N_16745,N_15517,N_15217);
and U16746 (N_16746,N_15894,N_15313);
and U16747 (N_16747,N_15251,N_15114);
and U16748 (N_16748,N_15406,N_15658);
or U16749 (N_16749,N_15899,N_15911);
or U16750 (N_16750,N_15870,N_15545);
nor U16751 (N_16751,N_15079,N_15551);
xnor U16752 (N_16752,N_15853,N_15245);
nand U16753 (N_16753,N_15672,N_15169);
nor U16754 (N_16754,N_15442,N_15491);
xnor U16755 (N_16755,N_15276,N_15653);
nor U16756 (N_16756,N_15074,N_15565);
or U16757 (N_16757,N_15201,N_15289);
nand U16758 (N_16758,N_15428,N_15534);
xnor U16759 (N_16759,N_15159,N_15185);
or U16760 (N_16760,N_15207,N_15553);
xor U16761 (N_16761,N_15345,N_15480);
xnor U16762 (N_16762,N_15840,N_15071);
or U16763 (N_16763,N_15914,N_15180);
and U16764 (N_16764,N_15822,N_15101);
and U16765 (N_16765,N_15373,N_15396);
or U16766 (N_16766,N_15747,N_15813);
nor U16767 (N_16767,N_15933,N_15396);
xnor U16768 (N_16768,N_15238,N_15794);
nor U16769 (N_16769,N_15147,N_15499);
or U16770 (N_16770,N_15533,N_15506);
xor U16771 (N_16771,N_15365,N_15794);
nand U16772 (N_16772,N_15980,N_15956);
nand U16773 (N_16773,N_15495,N_15969);
xor U16774 (N_16774,N_15949,N_15722);
and U16775 (N_16775,N_15195,N_15660);
nand U16776 (N_16776,N_15787,N_15783);
nand U16777 (N_16777,N_15880,N_15216);
nand U16778 (N_16778,N_15203,N_15325);
nand U16779 (N_16779,N_15969,N_15370);
nor U16780 (N_16780,N_15988,N_15548);
xnor U16781 (N_16781,N_15979,N_15901);
or U16782 (N_16782,N_15418,N_15557);
and U16783 (N_16783,N_15253,N_15936);
nor U16784 (N_16784,N_15236,N_15680);
nand U16785 (N_16785,N_15072,N_15570);
and U16786 (N_16786,N_15376,N_15416);
and U16787 (N_16787,N_15044,N_15829);
nor U16788 (N_16788,N_15064,N_15058);
or U16789 (N_16789,N_15503,N_15406);
nand U16790 (N_16790,N_15655,N_15712);
or U16791 (N_16791,N_15727,N_15625);
nand U16792 (N_16792,N_15914,N_15796);
and U16793 (N_16793,N_15863,N_15625);
nor U16794 (N_16794,N_15928,N_15809);
or U16795 (N_16795,N_15445,N_15249);
xnor U16796 (N_16796,N_15832,N_15817);
nor U16797 (N_16797,N_15342,N_15113);
and U16798 (N_16798,N_15378,N_15714);
nor U16799 (N_16799,N_15714,N_15291);
xnor U16800 (N_16800,N_15299,N_15762);
nor U16801 (N_16801,N_15648,N_15393);
and U16802 (N_16802,N_15255,N_15376);
or U16803 (N_16803,N_15201,N_15951);
nand U16804 (N_16804,N_15316,N_15396);
xor U16805 (N_16805,N_15509,N_15143);
nor U16806 (N_16806,N_15604,N_15524);
and U16807 (N_16807,N_15984,N_15086);
nand U16808 (N_16808,N_15681,N_15090);
xnor U16809 (N_16809,N_15134,N_15255);
and U16810 (N_16810,N_15893,N_15286);
nand U16811 (N_16811,N_15872,N_15422);
nor U16812 (N_16812,N_15876,N_15642);
xor U16813 (N_16813,N_15039,N_15185);
or U16814 (N_16814,N_15135,N_15267);
and U16815 (N_16815,N_15645,N_15345);
nand U16816 (N_16816,N_15924,N_15625);
or U16817 (N_16817,N_15190,N_15590);
or U16818 (N_16818,N_15954,N_15056);
nor U16819 (N_16819,N_15852,N_15186);
or U16820 (N_16820,N_15233,N_15592);
and U16821 (N_16821,N_15055,N_15449);
nand U16822 (N_16822,N_15386,N_15934);
or U16823 (N_16823,N_15399,N_15226);
and U16824 (N_16824,N_15153,N_15477);
or U16825 (N_16825,N_15066,N_15030);
and U16826 (N_16826,N_15555,N_15898);
xnor U16827 (N_16827,N_15721,N_15991);
or U16828 (N_16828,N_15989,N_15828);
or U16829 (N_16829,N_15066,N_15827);
or U16830 (N_16830,N_15069,N_15290);
and U16831 (N_16831,N_15926,N_15459);
or U16832 (N_16832,N_15221,N_15848);
or U16833 (N_16833,N_15530,N_15467);
nor U16834 (N_16834,N_15997,N_15085);
and U16835 (N_16835,N_15508,N_15296);
nand U16836 (N_16836,N_15924,N_15792);
nand U16837 (N_16837,N_15278,N_15202);
and U16838 (N_16838,N_15621,N_15240);
nand U16839 (N_16839,N_15647,N_15437);
or U16840 (N_16840,N_15926,N_15080);
nand U16841 (N_16841,N_15848,N_15001);
and U16842 (N_16842,N_15694,N_15658);
nor U16843 (N_16843,N_15436,N_15646);
or U16844 (N_16844,N_15952,N_15731);
xnor U16845 (N_16845,N_15930,N_15734);
and U16846 (N_16846,N_15551,N_15775);
or U16847 (N_16847,N_15274,N_15095);
or U16848 (N_16848,N_15813,N_15621);
nor U16849 (N_16849,N_15928,N_15454);
or U16850 (N_16850,N_15979,N_15990);
nor U16851 (N_16851,N_15951,N_15523);
nor U16852 (N_16852,N_15140,N_15425);
nor U16853 (N_16853,N_15969,N_15583);
nor U16854 (N_16854,N_15230,N_15424);
nor U16855 (N_16855,N_15655,N_15558);
and U16856 (N_16856,N_15901,N_15074);
or U16857 (N_16857,N_15003,N_15495);
or U16858 (N_16858,N_15191,N_15173);
nor U16859 (N_16859,N_15824,N_15691);
or U16860 (N_16860,N_15784,N_15778);
nand U16861 (N_16861,N_15717,N_15918);
xor U16862 (N_16862,N_15044,N_15998);
or U16863 (N_16863,N_15013,N_15284);
or U16864 (N_16864,N_15252,N_15822);
nor U16865 (N_16865,N_15657,N_15843);
nand U16866 (N_16866,N_15945,N_15122);
or U16867 (N_16867,N_15603,N_15274);
or U16868 (N_16868,N_15139,N_15557);
or U16869 (N_16869,N_15414,N_15251);
or U16870 (N_16870,N_15268,N_15120);
nand U16871 (N_16871,N_15512,N_15442);
xnor U16872 (N_16872,N_15570,N_15010);
or U16873 (N_16873,N_15749,N_15819);
and U16874 (N_16874,N_15840,N_15524);
or U16875 (N_16875,N_15333,N_15689);
nor U16876 (N_16876,N_15830,N_15704);
nand U16877 (N_16877,N_15639,N_15279);
and U16878 (N_16878,N_15877,N_15777);
xnor U16879 (N_16879,N_15712,N_15123);
nor U16880 (N_16880,N_15006,N_15821);
and U16881 (N_16881,N_15555,N_15838);
or U16882 (N_16882,N_15452,N_15049);
nand U16883 (N_16883,N_15844,N_15614);
nor U16884 (N_16884,N_15348,N_15809);
or U16885 (N_16885,N_15908,N_15657);
and U16886 (N_16886,N_15693,N_15155);
or U16887 (N_16887,N_15905,N_15161);
nor U16888 (N_16888,N_15165,N_15404);
and U16889 (N_16889,N_15376,N_15789);
or U16890 (N_16890,N_15755,N_15956);
and U16891 (N_16891,N_15064,N_15385);
nor U16892 (N_16892,N_15342,N_15525);
or U16893 (N_16893,N_15576,N_15587);
and U16894 (N_16894,N_15904,N_15992);
or U16895 (N_16895,N_15611,N_15530);
or U16896 (N_16896,N_15997,N_15999);
xnor U16897 (N_16897,N_15020,N_15019);
xor U16898 (N_16898,N_15606,N_15937);
nor U16899 (N_16899,N_15184,N_15339);
nor U16900 (N_16900,N_15091,N_15057);
xor U16901 (N_16901,N_15325,N_15811);
or U16902 (N_16902,N_15317,N_15277);
nor U16903 (N_16903,N_15816,N_15863);
and U16904 (N_16904,N_15400,N_15893);
xnor U16905 (N_16905,N_15453,N_15677);
nor U16906 (N_16906,N_15001,N_15473);
xnor U16907 (N_16907,N_15230,N_15659);
or U16908 (N_16908,N_15510,N_15465);
nand U16909 (N_16909,N_15653,N_15277);
or U16910 (N_16910,N_15624,N_15815);
nor U16911 (N_16911,N_15643,N_15972);
xor U16912 (N_16912,N_15181,N_15614);
xor U16913 (N_16913,N_15341,N_15181);
or U16914 (N_16914,N_15831,N_15303);
nand U16915 (N_16915,N_15956,N_15341);
xnor U16916 (N_16916,N_15690,N_15695);
and U16917 (N_16917,N_15016,N_15004);
or U16918 (N_16918,N_15998,N_15560);
nor U16919 (N_16919,N_15105,N_15426);
and U16920 (N_16920,N_15795,N_15497);
nand U16921 (N_16921,N_15098,N_15835);
or U16922 (N_16922,N_15451,N_15665);
or U16923 (N_16923,N_15202,N_15564);
or U16924 (N_16924,N_15065,N_15354);
xor U16925 (N_16925,N_15706,N_15770);
nand U16926 (N_16926,N_15994,N_15267);
and U16927 (N_16927,N_15658,N_15787);
and U16928 (N_16928,N_15016,N_15014);
nor U16929 (N_16929,N_15166,N_15040);
or U16930 (N_16930,N_15342,N_15884);
and U16931 (N_16931,N_15683,N_15250);
or U16932 (N_16932,N_15641,N_15982);
and U16933 (N_16933,N_15047,N_15878);
and U16934 (N_16934,N_15991,N_15273);
or U16935 (N_16935,N_15679,N_15510);
nand U16936 (N_16936,N_15620,N_15734);
or U16937 (N_16937,N_15157,N_15767);
and U16938 (N_16938,N_15470,N_15507);
nand U16939 (N_16939,N_15364,N_15904);
and U16940 (N_16940,N_15677,N_15282);
xnor U16941 (N_16941,N_15843,N_15169);
and U16942 (N_16942,N_15282,N_15940);
or U16943 (N_16943,N_15011,N_15015);
nor U16944 (N_16944,N_15732,N_15079);
or U16945 (N_16945,N_15052,N_15010);
nand U16946 (N_16946,N_15281,N_15705);
nor U16947 (N_16947,N_15450,N_15432);
and U16948 (N_16948,N_15917,N_15663);
and U16949 (N_16949,N_15241,N_15362);
or U16950 (N_16950,N_15828,N_15165);
or U16951 (N_16951,N_15311,N_15406);
nand U16952 (N_16952,N_15719,N_15328);
xnor U16953 (N_16953,N_15821,N_15301);
nor U16954 (N_16954,N_15634,N_15201);
nor U16955 (N_16955,N_15066,N_15715);
xnor U16956 (N_16956,N_15940,N_15125);
xor U16957 (N_16957,N_15938,N_15365);
xnor U16958 (N_16958,N_15811,N_15419);
or U16959 (N_16959,N_15248,N_15783);
nor U16960 (N_16960,N_15448,N_15884);
nor U16961 (N_16961,N_15592,N_15611);
or U16962 (N_16962,N_15159,N_15226);
and U16963 (N_16963,N_15114,N_15985);
xor U16964 (N_16964,N_15050,N_15444);
and U16965 (N_16965,N_15902,N_15042);
nor U16966 (N_16966,N_15888,N_15233);
nand U16967 (N_16967,N_15065,N_15753);
and U16968 (N_16968,N_15464,N_15273);
or U16969 (N_16969,N_15706,N_15935);
nand U16970 (N_16970,N_15189,N_15441);
or U16971 (N_16971,N_15486,N_15314);
or U16972 (N_16972,N_15322,N_15512);
nand U16973 (N_16973,N_15526,N_15798);
and U16974 (N_16974,N_15089,N_15693);
and U16975 (N_16975,N_15725,N_15752);
nor U16976 (N_16976,N_15582,N_15442);
and U16977 (N_16977,N_15072,N_15950);
xor U16978 (N_16978,N_15326,N_15759);
and U16979 (N_16979,N_15553,N_15899);
or U16980 (N_16980,N_15065,N_15905);
or U16981 (N_16981,N_15108,N_15426);
nor U16982 (N_16982,N_15867,N_15550);
and U16983 (N_16983,N_15916,N_15080);
or U16984 (N_16984,N_15960,N_15390);
nand U16985 (N_16985,N_15705,N_15074);
or U16986 (N_16986,N_15704,N_15542);
or U16987 (N_16987,N_15089,N_15864);
nand U16988 (N_16988,N_15989,N_15011);
xor U16989 (N_16989,N_15097,N_15024);
or U16990 (N_16990,N_15774,N_15951);
nor U16991 (N_16991,N_15410,N_15530);
nand U16992 (N_16992,N_15572,N_15960);
xnor U16993 (N_16993,N_15892,N_15380);
or U16994 (N_16994,N_15532,N_15995);
and U16995 (N_16995,N_15131,N_15929);
and U16996 (N_16996,N_15955,N_15192);
or U16997 (N_16997,N_15434,N_15911);
nor U16998 (N_16998,N_15395,N_15406);
xnor U16999 (N_16999,N_15855,N_15321);
or U17000 (N_17000,N_16173,N_16796);
xnor U17001 (N_17001,N_16007,N_16309);
nand U17002 (N_17002,N_16122,N_16810);
nor U17003 (N_17003,N_16944,N_16166);
and U17004 (N_17004,N_16013,N_16237);
nor U17005 (N_17005,N_16652,N_16439);
or U17006 (N_17006,N_16224,N_16413);
and U17007 (N_17007,N_16400,N_16664);
or U17008 (N_17008,N_16424,N_16996);
xnor U17009 (N_17009,N_16759,N_16615);
and U17010 (N_17010,N_16164,N_16351);
and U17011 (N_17011,N_16849,N_16573);
or U17012 (N_17012,N_16828,N_16109);
xor U17013 (N_17013,N_16307,N_16291);
xnor U17014 (N_17014,N_16199,N_16375);
nand U17015 (N_17015,N_16865,N_16541);
nor U17016 (N_17016,N_16232,N_16257);
xnor U17017 (N_17017,N_16586,N_16948);
nand U17018 (N_17018,N_16911,N_16967);
xnor U17019 (N_17019,N_16775,N_16107);
nand U17020 (N_17020,N_16547,N_16298);
nor U17021 (N_17021,N_16635,N_16834);
nand U17022 (N_17022,N_16373,N_16151);
nand U17023 (N_17023,N_16879,N_16843);
nor U17024 (N_17024,N_16123,N_16467);
and U17025 (N_17025,N_16859,N_16786);
and U17026 (N_17026,N_16031,N_16874);
or U17027 (N_17027,N_16645,N_16126);
or U17028 (N_17028,N_16771,N_16281);
nor U17029 (N_17029,N_16113,N_16130);
or U17030 (N_17030,N_16358,N_16557);
and U17031 (N_17031,N_16788,N_16612);
xnor U17032 (N_17032,N_16082,N_16215);
nand U17033 (N_17033,N_16114,N_16914);
nor U17034 (N_17034,N_16794,N_16324);
and U17035 (N_17035,N_16686,N_16345);
or U17036 (N_17036,N_16198,N_16561);
nand U17037 (N_17037,N_16760,N_16527);
xnor U17038 (N_17038,N_16384,N_16691);
nand U17039 (N_17039,N_16427,N_16341);
and U17040 (N_17040,N_16722,N_16010);
or U17041 (N_17041,N_16390,N_16473);
or U17042 (N_17042,N_16693,N_16779);
or U17043 (N_17043,N_16105,N_16209);
nor U17044 (N_17044,N_16054,N_16617);
nand U17045 (N_17045,N_16753,N_16295);
nor U17046 (N_17046,N_16012,N_16918);
xor U17047 (N_17047,N_16866,N_16804);
xnor U17048 (N_17048,N_16334,N_16930);
and U17049 (N_17049,N_16726,N_16651);
xor U17050 (N_17050,N_16285,N_16666);
nand U17051 (N_17051,N_16220,N_16023);
nor U17052 (N_17052,N_16658,N_16250);
or U17053 (N_17053,N_16063,N_16368);
xnor U17054 (N_17054,N_16174,N_16141);
or U17055 (N_17055,N_16803,N_16370);
xnor U17056 (N_17056,N_16349,N_16070);
nor U17057 (N_17057,N_16221,N_16036);
nand U17058 (N_17058,N_16171,N_16044);
nand U17059 (N_17059,N_16102,N_16144);
or U17060 (N_17060,N_16569,N_16361);
xnor U17061 (N_17061,N_16040,N_16764);
nor U17062 (N_17062,N_16533,N_16405);
nand U17063 (N_17063,N_16793,N_16266);
nor U17064 (N_17064,N_16742,N_16327);
or U17065 (N_17065,N_16820,N_16520);
xor U17066 (N_17066,N_16156,N_16618);
nor U17067 (N_17067,N_16850,N_16430);
and U17068 (N_17068,N_16366,N_16041);
nor U17069 (N_17069,N_16657,N_16555);
xor U17070 (N_17070,N_16584,N_16603);
and U17071 (N_17071,N_16488,N_16087);
nand U17072 (N_17072,N_16184,N_16821);
or U17073 (N_17073,N_16489,N_16714);
xor U17074 (N_17074,N_16409,N_16931);
nor U17075 (N_17075,N_16238,N_16043);
xnor U17076 (N_17076,N_16441,N_16449);
and U17077 (N_17077,N_16412,N_16721);
xor U17078 (N_17078,N_16460,N_16050);
nor U17079 (N_17079,N_16301,N_16127);
and U17080 (N_17080,N_16668,N_16862);
and U17081 (N_17081,N_16567,N_16538);
xor U17082 (N_17082,N_16505,N_16328);
or U17083 (N_17083,N_16983,N_16492);
xor U17084 (N_17084,N_16592,N_16813);
nand U17085 (N_17085,N_16957,N_16097);
xnor U17086 (N_17086,N_16723,N_16801);
or U17087 (N_17087,N_16827,N_16112);
nor U17088 (N_17088,N_16515,N_16069);
nand U17089 (N_17089,N_16032,N_16320);
nand U17090 (N_17090,N_16682,N_16522);
nand U17091 (N_17091,N_16696,N_16818);
or U17092 (N_17092,N_16797,N_16213);
nor U17093 (N_17093,N_16971,N_16554);
nand U17094 (N_17094,N_16734,N_16244);
nor U17095 (N_17095,N_16442,N_16056);
nand U17096 (N_17096,N_16816,N_16643);
and U17097 (N_17097,N_16511,N_16832);
nor U17098 (N_17098,N_16240,N_16030);
nor U17099 (N_17099,N_16392,N_16282);
or U17100 (N_17100,N_16839,N_16762);
nor U17101 (N_17101,N_16672,N_16229);
nor U17102 (N_17102,N_16096,N_16429);
xnor U17103 (N_17103,N_16684,N_16275);
nand U17104 (N_17104,N_16873,N_16108);
nor U17105 (N_17105,N_16508,N_16419);
nand U17106 (N_17106,N_16552,N_16894);
nor U17107 (N_17107,N_16751,N_16490);
nor U17108 (N_17108,N_16665,N_16809);
or U17109 (N_17109,N_16770,N_16758);
nand U17110 (N_17110,N_16381,N_16134);
and U17111 (N_17111,N_16808,N_16984);
nor U17112 (N_17112,N_16332,N_16104);
nor U17113 (N_17113,N_16811,N_16098);
nor U17114 (N_17114,N_16423,N_16812);
nand U17115 (N_17115,N_16523,N_16744);
and U17116 (N_17116,N_16896,N_16646);
and U17117 (N_17117,N_16431,N_16579);
nand U17118 (N_17118,N_16611,N_16667);
or U17119 (N_17119,N_16656,N_16973);
xor U17120 (N_17120,N_16989,N_16288);
or U17121 (N_17121,N_16057,N_16754);
nand U17122 (N_17122,N_16729,N_16622);
nand U17123 (N_17123,N_16374,N_16993);
xnor U17124 (N_17124,N_16219,N_16319);
or U17125 (N_17125,N_16922,N_16575);
and U17126 (N_17126,N_16673,N_16662);
and U17127 (N_17127,N_16895,N_16225);
xnor U17128 (N_17128,N_16958,N_16011);
and U17129 (N_17129,N_16230,N_16774);
nand U17130 (N_17130,N_16443,N_16417);
or U17131 (N_17131,N_16582,N_16871);
xor U17132 (N_17132,N_16580,N_16551);
or U17133 (N_17133,N_16572,N_16035);
xnor U17134 (N_17134,N_16343,N_16318);
or U17135 (N_17135,N_16780,N_16197);
nor U17136 (N_17136,N_16607,N_16929);
or U17137 (N_17137,N_16073,N_16461);
nand U17138 (N_17138,N_16325,N_16946);
and U17139 (N_17139,N_16840,N_16806);
and U17140 (N_17140,N_16891,N_16317);
xnor U17141 (N_17141,N_16453,N_16350);
and U17142 (N_17142,N_16120,N_16480);
and U17143 (N_17143,N_16704,N_16718);
xnor U17144 (N_17144,N_16943,N_16814);
xnor U17145 (N_17145,N_16649,N_16919);
and U17146 (N_17146,N_16934,N_16258);
and U17147 (N_17147,N_16176,N_16581);
nor U17148 (N_17148,N_16792,N_16578);
or U17149 (N_17149,N_16360,N_16132);
nand U17150 (N_17150,N_16017,N_16819);
xor U17151 (N_17151,N_16302,N_16817);
and U17152 (N_17152,N_16773,N_16708);
and U17153 (N_17153,N_16585,N_16624);
nand U17154 (N_17154,N_16293,N_16273);
and U17155 (N_17155,N_16836,N_16529);
or U17156 (N_17156,N_16600,N_16954);
nand U17157 (N_17157,N_16484,N_16616);
nand U17158 (N_17158,N_16383,N_16245);
nor U17159 (N_17159,N_16394,N_16550);
nand U17160 (N_17160,N_16937,N_16464);
or U17161 (N_17161,N_16660,N_16732);
and U17162 (N_17162,N_16494,N_16239);
xnor U17163 (N_17163,N_16716,N_16641);
or U17164 (N_17164,N_16982,N_16211);
and U17165 (N_17165,N_16287,N_16458);
xor U17166 (N_17166,N_16678,N_16393);
and U17167 (N_17167,N_16588,N_16795);
or U17168 (N_17168,N_16083,N_16103);
or U17169 (N_17169,N_16844,N_16933);
or U17170 (N_17170,N_16669,N_16433);
xnor U17171 (N_17171,N_16680,N_16995);
or U17172 (N_17172,N_16998,N_16500);
xnor U17173 (N_17173,N_16084,N_16081);
and U17174 (N_17174,N_16162,N_16885);
nor U17175 (N_17175,N_16904,N_16997);
nor U17176 (N_17176,N_16064,N_16822);
or U17177 (N_17177,N_16408,N_16829);
xnor U17178 (N_17178,N_16340,N_16479);
nand U17179 (N_17179,N_16605,N_16259);
xor U17180 (N_17180,N_16227,N_16493);
nor U17181 (N_17181,N_16614,N_16707);
and U17182 (N_17182,N_16299,N_16181);
or U17183 (N_17183,N_16938,N_16459);
nand U17184 (N_17184,N_16071,N_16025);
nor U17185 (N_17185,N_16719,N_16205);
nand U17186 (N_17186,N_16304,N_16698);
xnor U17187 (N_17187,N_16015,N_16175);
nor U17188 (N_17188,N_16642,N_16941);
nand U17189 (N_17189,N_16034,N_16677);
nor U17190 (N_17190,N_16711,N_16457);
and U17191 (N_17191,N_16422,N_16653);
and U17192 (N_17192,N_16481,N_16100);
nor U17193 (N_17193,N_16524,N_16969);
nand U17194 (N_17194,N_16870,N_16671);
nor U17195 (N_17195,N_16783,N_16356);
or U17196 (N_17196,N_16777,N_16236);
nand U17197 (N_17197,N_16060,N_16474);
or U17198 (N_17198,N_16532,N_16210);
xnor U17199 (N_17199,N_16344,N_16853);
nand U17200 (N_17200,N_16029,N_16633);
xor U17201 (N_17201,N_16387,N_16968);
or U17202 (N_17202,N_16976,N_16496);
or U17203 (N_17203,N_16226,N_16475);
nand U17204 (N_17204,N_16644,N_16663);
xnor U17205 (N_17205,N_16906,N_16313);
or U17206 (N_17206,N_16516,N_16689);
nand U17207 (N_17207,N_16949,N_16487);
xor U17208 (N_17208,N_16452,N_16763);
or U17209 (N_17209,N_16602,N_16994);
nor U17210 (N_17210,N_16051,N_16207);
and U17211 (N_17211,N_16129,N_16274);
xor U17212 (N_17212,N_16756,N_16899);
nand U17213 (N_17213,N_16978,N_16518);
nor U17214 (N_17214,N_16599,N_16267);
nor U17215 (N_17215,N_16333,N_16628);
xnor U17216 (N_17216,N_16425,N_16868);
nor U17217 (N_17217,N_16090,N_16901);
nand U17218 (N_17218,N_16420,N_16396);
nor U17219 (N_17219,N_16039,N_16253);
xnor U17220 (N_17220,N_16388,N_16000);
xor U17221 (N_17221,N_16296,N_16284);
and U17222 (N_17222,N_16619,N_16887);
nand U17223 (N_17223,N_16466,N_16234);
nor U17224 (N_17224,N_16765,N_16093);
nor U17225 (N_17225,N_16709,N_16512);
or U17226 (N_17226,N_16790,N_16322);
nor U17227 (N_17227,N_16451,N_16848);
nor U17228 (N_17228,N_16428,N_16263);
or U17229 (N_17229,N_16372,N_16182);
nor U17230 (N_17230,N_16143,N_16079);
or U17231 (N_17231,N_16179,N_16336);
and U17232 (N_17232,N_16647,N_16142);
xnor U17233 (N_17233,N_16787,N_16359);
nand U17234 (N_17234,N_16153,N_16300);
and U17235 (N_17235,N_16228,N_16426);
nand U17236 (N_17236,N_16528,N_16674);
nand U17237 (N_17237,N_16727,N_16942);
and U17238 (N_17238,N_16486,N_16566);
nor U17239 (N_17239,N_16331,N_16315);
nand U17240 (N_17240,N_16119,N_16864);
or U17241 (N_17241,N_16625,N_16927);
nand U17242 (N_17242,N_16498,N_16217);
and U17243 (N_17243,N_16246,N_16306);
nand U17244 (N_17244,N_16634,N_16154);
nor U17245 (N_17245,N_16363,N_16297);
or U17246 (N_17246,N_16837,N_16308);
nand U17247 (N_17247,N_16735,N_16769);
nor U17248 (N_17248,N_16111,N_16415);
xnor U17249 (N_17249,N_16124,N_16601);
xnor U17250 (N_17250,N_16563,N_16776);
or U17251 (N_17251,N_16590,N_16469);
xnor U17252 (N_17252,N_16110,N_16168);
xor U17253 (N_17253,N_16835,N_16861);
nor U17254 (N_17254,N_16909,N_16330);
nor U17255 (N_17255,N_16831,N_16212);
or U17256 (N_17256,N_16986,N_16101);
nor U17257 (N_17257,N_16398,N_16546);
nor U17258 (N_17258,N_16980,N_16021);
xnor U17259 (N_17259,N_16401,N_16167);
or U17260 (N_17260,N_16379,N_16977);
xnor U17261 (N_17261,N_16339,N_16465);
nand U17262 (N_17262,N_16889,N_16826);
nor U17263 (N_17263,N_16755,N_16235);
nor U17264 (N_17264,N_16856,N_16289);
nor U17265 (N_17265,N_16730,N_16655);
nand U17266 (N_17266,N_16278,N_16935);
nor U17267 (N_17267,N_16781,N_16362);
xnor U17268 (N_17268,N_16138,N_16845);
or U17269 (N_17269,N_16076,N_16193);
xor U17270 (N_17270,N_16369,N_16888);
xor U17271 (N_17271,N_16145,N_16847);
xnor U17272 (N_17272,N_16782,N_16728);
xor U17273 (N_17273,N_16846,N_16531);
nand U17274 (N_17274,N_16536,N_16432);
xnor U17275 (N_17275,N_16312,N_16936);
or U17276 (N_17276,N_16118,N_16875);
and U17277 (N_17277,N_16654,N_16157);
xnor U17278 (N_17278,N_16066,N_16947);
nor U17279 (N_17279,N_16049,N_16446);
nor U17280 (N_17280,N_16725,N_16715);
or U17281 (N_17281,N_16881,N_16807);
xnor U17282 (N_17282,N_16216,N_16706);
and U17283 (N_17283,N_16337,N_16276);
or U17284 (N_17284,N_16953,N_16610);
nand U17285 (N_17285,N_16506,N_16009);
nand U17286 (N_17286,N_16410,N_16397);
or U17287 (N_17287,N_16477,N_16152);
or U17288 (N_17288,N_16893,N_16921);
xnor U17289 (N_17289,N_16833,N_16208);
and U17290 (N_17290,N_16086,N_16277);
nor U17291 (N_17291,N_16194,N_16077);
and U17292 (N_17292,N_16137,N_16188);
nand U17293 (N_17293,N_16172,N_16192);
or U17294 (N_17294,N_16890,N_16435);
xor U17295 (N_17295,N_16418,N_16699);
xnor U17296 (N_17296,N_16731,N_16106);
nor U17297 (N_17297,N_16380,N_16648);
nand U17298 (N_17298,N_16596,N_16627);
or U17299 (N_17299,N_16437,N_16553);
xnor U17300 (N_17300,N_16860,N_16200);
and U17301 (N_17301,N_16008,N_16975);
nor U17302 (N_17302,N_16987,N_16979);
xor U17303 (N_17303,N_16187,N_16434);
nand U17304 (N_17304,N_16687,N_16824);
nand U17305 (N_17305,N_16591,N_16231);
xor U17306 (N_17306,N_16038,N_16544);
xor U17307 (N_17307,N_16741,N_16037);
nor U17308 (N_17308,N_16447,N_16990);
nor U17309 (N_17309,N_16757,N_16951);
and U17310 (N_17310,N_16170,N_16745);
or U17311 (N_17311,N_16637,N_16700);
nand U17312 (N_17312,N_16499,N_16883);
or U17313 (N_17313,N_16202,N_16046);
nor U17314 (N_17314,N_16863,N_16004);
and U17315 (N_17315,N_16365,N_16915);
or U17316 (N_17316,N_16342,N_16454);
and U17317 (N_17317,N_16815,N_16355);
nor U17318 (N_17318,N_16713,N_16024);
and U17319 (N_17319,N_16404,N_16444);
and U17320 (N_17320,N_16950,N_16399);
nor U17321 (N_17321,N_16115,N_16631);
nand U17322 (N_17322,N_16683,N_16504);
nor U17323 (N_17323,N_16346,N_16970);
nor U17324 (N_17324,N_16088,N_16436);
and U17325 (N_17325,N_16543,N_16456);
nand U17326 (N_17326,N_16352,N_16403);
and U17327 (N_17327,N_16857,N_16353);
nand U17328 (N_17328,N_16406,N_16639);
xnor U17329 (N_17329,N_16303,N_16147);
nor U17330 (N_17330,N_16802,N_16574);
nand U17331 (N_17331,N_16882,N_16905);
xnor U17332 (N_17332,N_16926,N_16099);
nor U17333 (N_17333,N_16048,N_16752);
xnor U17334 (N_17334,N_16470,N_16535);
nor U17335 (N_17335,N_16165,N_16135);
and U17336 (N_17336,N_16169,N_16521);
xnor U17337 (N_17337,N_16485,N_16163);
xnor U17338 (N_17338,N_16981,N_16326);
nand U17339 (N_17339,N_16471,N_16468);
nor U17340 (N_17340,N_16005,N_16548);
xor U17341 (N_17341,N_16694,N_16695);
and U17342 (N_17342,N_16159,N_16242);
or U17343 (N_17343,N_16146,N_16247);
and U17344 (N_17344,N_16478,N_16907);
and U17345 (N_17345,N_16438,N_16903);
nor U17346 (N_17346,N_16377,N_16960);
and U17347 (N_17347,N_16670,N_16502);
nand U17348 (N_17348,N_16006,N_16201);
xor U17349 (N_17349,N_16183,N_16150);
xor U17350 (N_17350,N_16558,N_16280);
nand U17351 (N_17351,N_16851,N_16988);
xnor U17352 (N_17352,N_16290,N_16196);
nor U17353 (N_17353,N_16078,N_16450);
or U17354 (N_17354,N_16898,N_16630);
nor U17355 (N_17355,N_16329,N_16241);
and U17356 (N_17356,N_16710,N_16052);
nor U17357 (N_17357,N_16910,N_16869);
or U17358 (N_17358,N_16877,N_16391);
or U17359 (N_17359,N_16286,N_16402);
nand U17360 (N_17360,N_16260,N_16149);
xor U17361 (N_17361,N_16772,N_16133);
or U17362 (N_17362,N_16992,N_16854);
xor U17363 (N_17363,N_16606,N_16002);
xor U17364 (N_17364,N_16206,N_16676);
or U17365 (N_17365,N_16269,N_16026);
or U17366 (N_17366,N_16621,N_16852);
or U17367 (N_17367,N_16195,N_16019);
and U17368 (N_17368,N_16513,N_16095);
xnor U17369 (N_17369,N_16092,N_16091);
nand U17370 (N_17370,N_16738,N_16872);
nand U17371 (N_17371,N_16491,N_16638);
xnor U17372 (N_17372,N_16233,N_16749);
nor U17373 (N_17373,N_16629,N_16924);
nand U17374 (N_17374,N_16094,N_16913);
nand U17375 (N_17375,N_16072,N_16576);
nor U17376 (N_17376,N_16061,N_16784);
or U17377 (N_17377,N_16311,N_16371);
xor U17378 (N_17378,N_16161,N_16539);
nand U17379 (N_17379,N_16577,N_16027);
xor U17380 (N_17380,N_16594,N_16128);
or U17381 (N_17381,N_16675,N_16445);
nor U17382 (N_17382,N_16746,N_16799);
or U17383 (N_17383,N_16568,N_16160);
nand U17384 (N_17384,N_16136,N_16705);
and U17385 (N_17385,N_16902,N_16085);
nand U17386 (N_17386,N_16892,N_16766);
nand U17387 (N_17387,N_16067,N_16357);
and U17388 (N_17388,N_16559,N_16495);
and U17389 (N_17389,N_16254,N_16823);
xnor U17390 (N_17390,N_16501,N_16310);
or U17391 (N_17391,N_16867,N_16932);
xor U17392 (N_17392,N_16016,N_16940);
nand U17393 (N_17393,N_16305,N_16956);
or U17394 (N_17394,N_16283,N_16761);
nand U17395 (N_17395,N_16570,N_16701);
nor U17396 (N_17396,N_16203,N_16962);
xor U17397 (N_17397,N_16540,N_16367);
or U17398 (N_17398,N_16798,N_16650);
xor U17399 (N_17399,N_16855,N_16014);
nor U17400 (N_17400,N_16791,N_16908);
or U17401 (N_17401,N_16321,N_16121);
or U17402 (N_17402,N_16800,N_16571);
xnor U17403 (N_17403,N_16830,N_16661);
nand U17404 (N_17404,N_16264,N_16117);
or U17405 (N_17405,N_16858,N_16131);
nor U17406 (N_17406,N_16251,N_16916);
and U17407 (N_17407,N_16534,N_16679);
and U17408 (N_17408,N_16003,N_16743);
nor U17409 (N_17409,N_16062,N_16271);
nor U17410 (N_17410,N_16537,N_16560);
nor U17411 (N_17411,N_16598,N_16985);
nor U17412 (N_17412,N_16878,N_16065);
nor U17413 (N_17413,N_16116,N_16632);
nand U17414 (N_17414,N_16385,N_16270);
nor U17415 (N_17415,N_16335,N_16692);
and U17416 (N_17416,N_16733,N_16750);
nand U17417 (N_17417,N_16900,N_16497);
nand U17418 (N_17418,N_16389,N_16747);
xor U17419 (N_17419,N_16549,N_16059);
and U17420 (N_17420,N_16964,N_16055);
nand U17421 (N_17421,N_16255,N_16767);
nor U17422 (N_17422,N_16825,N_16125);
and U17423 (N_17423,N_16256,N_16685);
nand U17424 (N_17424,N_16440,N_16525);
and U17425 (N_17425,N_16636,N_16503);
and U17426 (N_17426,N_16681,N_16785);
and U17427 (N_17427,N_16354,N_16789);
xor U17428 (N_17428,N_16688,N_16020);
nor U17429 (N_17429,N_16414,N_16884);
and U17430 (N_17430,N_16186,N_16880);
nor U17431 (N_17431,N_16876,N_16462);
or U17432 (N_17432,N_16952,N_16659);
and U17433 (N_17433,N_16028,N_16542);
or U17434 (N_17434,N_16348,N_16920);
nand U17435 (N_17435,N_16620,N_16075);
and U17436 (N_17436,N_16925,N_16139);
nor U17437 (N_17437,N_16294,N_16421);
or U17438 (N_17438,N_16378,N_16448);
or U17439 (N_17439,N_16190,N_16045);
nor U17440 (N_17440,N_16955,N_16185);
nor U17441 (N_17441,N_16476,N_16080);
xnor U17442 (N_17442,N_16712,N_16047);
xnor U17443 (N_17443,N_16292,N_16376);
and U17444 (N_17444,N_16974,N_16140);
or U17445 (N_17445,N_16805,N_16223);
xor U17446 (N_17446,N_16177,N_16609);
nand U17447 (N_17447,N_16702,N_16963);
or U17448 (N_17448,N_16626,N_16737);
nor U17449 (N_17449,N_16961,N_16033);
and U17450 (N_17450,N_16268,N_16608);
xnor U17451 (N_17451,N_16068,N_16178);
and U17452 (N_17452,N_16514,N_16519);
xnor U17453 (N_17453,N_16966,N_16697);
xnor U17454 (N_17454,N_16768,N_16214);
and U17455 (N_17455,N_16597,N_16917);
xnor U17456 (N_17456,N_16739,N_16623);
nand U17457 (N_17457,N_16042,N_16510);
nand U17458 (N_17458,N_16841,N_16928);
nand U17459 (N_17459,N_16564,N_16074);
xor U17460 (N_17460,N_16483,N_16472);
nand U17461 (N_17461,N_16395,N_16222);
or U17462 (N_17462,N_16022,N_16886);
nor U17463 (N_17463,N_16939,N_16556);
xor U17464 (N_17464,N_16243,N_16338);
xnor U17465 (N_17465,N_16314,N_16261);
nor U17466 (N_17466,N_16316,N_16604);
nand U17467 (N_17467,N_16583,N_16416);
nand U17468 (N_17468,N_16640,N_16740);
xnor U17469 (N_17469,N_16509,N_16058);
and U17470 (N_17470,N_16279,N_16018);
xor U17471 (N_17471,N_16897,N_16972);
or U17472 (N_17472,N_16191,N_16180);
nand U17473 (N_17473,N_16703,N_16545);
nor U17474 (N_17474,N_16158,N_16736);
nand U17475 (N_17475,N_16562,N_16089);
nor U17476 (N_17476,N_16463,N_16218);
nand U17477 (N_17477,N_16249,N_16526);
and U17478 (N_17478,N_16364,N_16595);
nor U17479 (N_17479,N_16999,N_16517);
xor U17480 (N_17480,N_16189,N_16262);
or U17481 (N_17481,N_16838,N_16455);
or U17482 (N_17482,N_16347,N_16690);
and U17483 (N_17483,N_16482,N_16748);
nor U17484 (N_17484,N_16204,N_16001);
nor U17485 (N_17485,N_16842,N_16382);
nor U17486 (N_17486,N_16386,N_16411);
or U17487 (N_17487,N_16252,N_16565);
nand U17488 (N_17488,N_16923,N_16272);
nor U17489 (N_17489,N_16148,N_16265);
xor U17490 (N_17490,N_16530,N_16613);
xor U17491 (N_17491,N_16155,N_16912);
or U17492 (N_17492,N_16053,N_16323);
or U17493 (N_17493,N_16724,N_16778);
nand U17494 (N_17494,N_16959,N_16587);
and U17495 (N_17495,N_16991,N_16248);
xnor U17496 (N_17496,N_16945,N_16717);
and U17497 (N_17497,N_16965,N_16407);
or U17498 (N_17498,N_16720,N_16593);
xnor U17499 (N_17499,N_16507,N_16589);
or U17500 (N_17500,N_16692,N_16471);
nor U17501 (N_17501,N_16508,N_16477);
or U17502 (N_17502,N_16736,N_16840);
or U17503 (N_17503,N_16833,N_16715);
nand U17504 (N_17504,N_16302,N_16172);
or U17505 (N_17505,N_16045,N_16757);
nand U17506 (N_17506,N_16516,N_16125);
nor U17507 (N_17507,N_16928,N_16872);
nor U17508 (N_17508,N_16204,N_16056);
nand U17509 (N_17509,N_16911,N_16282);
xor U17510 (N_17510,N_16631,N_16442);
and U17511 (N_17511,N_16163,N_16956);
and U17512 (N_17512,N_16252,N_16996);
xor U17513 (N_17513,N_16333,N_16433);
nand U17514 (N_17514,N_16453,N_16837);
and U17515 (N_17515,N_16215,N_16258);
and U17516 (N_17516,N_16936,N_16849);
nand U17517 (N_17517,N_16574,N_16534);
nand U17518 (N_17518,N_16782,N_16036);
or U17519 (N_17519,N_16344,N_16065);
nand U17520 (N_17520,N_16907,N_16876);
nor U17521 (N_17521,N_16280,N_16763);
xnor U17522 (N_17522,N_16608,N_16762);
nand U17523 (N_17523,N_16785,N_16720);
nor U17524 (N_17524,N_16204,N_16036);
and U17525 (N_17525,N_16841,N_16597);
or U17526 (N_17526,N_16025,N_16385);
nand U17527 (N_17527,N_16588,N_16689);
nand U17528 (N_17528,N_16529,N_16554);
and U17529 (N_17529,N_16569,N_16811);
or U17530 (N_17530,N_16303,N_16162);
and U17531 (N_17531,N_16630,N_16172);
xor U17532 (N_17532,N_16104,N_16440);
xor U17533 (N_17533,N_16007,N_16336);
xor U17534 (N_17534,N_16299,N_16348);
nand U17535 (N_17535,N_16238,N_16956);
nand U17536 (N_17536,N_16317,N_16263);
nand U17537 (N_17537,N_16573,N_16025);
and U17538 (N_17538,N_16877,N_16220);
xnor U17539 (N_17539,N_16093,N_16152);
and U17540 (N_17540,N_16618,N_16694);
xor U17541 (N_17541,N_16690,N_16084);
xor U17542 (N_17542,N_16898,N_16616);
nand U17543 (N_17543,N_16246,N_16455);
nor U17544 (N_17544,N_16918,N_16196);
nand U17545 (N_17545,N_16212,N_16146);
xnor U17546 (N_17546,N_16815,N_16978);
or U17547 (N_17547,N_16632,N_16230);
nor U17548 (N_17548,N_16234,N_16812);
or U17549 (N_17549,N_16496,N_16123);
nor U17550 (N_17550,N_16691,N_16057);
nand U17551 (N_17551,N_16038,N_16473);
and U17552 (N_17552,N_16651,N_16919);
nor U17553 (N_17553,N_16692,N_16807);
nand U17554 (N_17554,N_16565,N_16085);
and U17555 (N_17555,N_16524,N_16134);
nand U17556 (N_17556,N_16380,N_16026);
or U17557 (N_17557,N_16435,N_16245);
xor U17558 (N_17558,N_16346,N_16435);
xnor U17559 (N_17559,N_16128,N_16740);
or U17560 (N_17560,N_16090,N_16741);
or U17561 (N_17561,N_16169,N_16147);
xor U17562 (N_17562,N_16278,N_16001);
or U17563 (N_17563,N_16116,N_16570);
xnor U17564 (N_17564,N_16380,N_16943);
nand U17565 (N_17565,N_16496,N_16242);
nor U17566 (N_17566,N_16328,N_16240);
or U17567 (N_17567,N_16970,N_16746);
nand U17568 (N_17568,N_16613,N_16840);
nand U17569 (N_17569,N_16266,N_16231);
nand U17570 (N_17570,N_16242,N_16531);
nor U17571 (N_17571,N_16529,N_16776);
and U17572 (N_17572,N_16164,N_16992);
or U17573 (N_17573,N_16300,N_16773);
xor U17574 (N_17574,N_16016,N_16391);
nand U17575 (N_17575,N_16784,N_16131);
nand U17576 (N_17576,N_16704,N_16449);
nand U17577 (N_17577,N_16552,N_16519);
and U17578 (N_17578,N_16522,N_16832);
and U17579 (N_17579,N_16189,N_16823);
and U17580 (N_17580,N_16698,N_16651);
nand U17581 (N_17581,N_16581,N_16121);
or U17582 (N_17582,N_16243,N_16778);
nor U17583 (N_17583,N_16093,N_16467);
xnor U17584 (N_17584,N_16470,N_16769);
and U17585 (N_17585,N_16537,N_16758);
or U17586 (N_17586,N_16210,N_16585);
and U17587 (N_17587,N_16671,N_16262);
nor U17588 (N_17588,N_16068,N_16171);
nor U17589 (N_17589,N_16691,N_16302);
and U17590 (N_17590,N_16921,N_16907);
xor U17591 (N_17591,N_16765,N_16272);
and U17592 (N_17592,N_16184,N_16221);
xnor U17593 (N_17593,N_16472,N_16639);
nor U17594 (N_17594,N_16192,N_16517);
and U17595 (N_17595,N_16231,N_16836);
and U17596 (N_17596,N_16343,N_16726);
nor U17597 (N_17597,N_16173,N_16843);
or U17598 (N_17598,N_16533,N_16429);
xnor U17599 (N_17599,N_16295,N_16106);
or U17600 (N_17600,N_16363,N_16459);
nand U17601 (N_17601,N_16550,N_16112);
and U17602 (N_17602,N_16308,N_16890);
nor U17603 (N_17603,N_16312,N_16125);
xor U17604 (N_17604,N_16830,N_16816);
nand U17605 (N_17605,N_16861,N_16687);
nand U17606 (N_17606,N_16038,N_16760);
nand U17607 (N_17607,N_16631,N_16855);
and U17608 (N_17608,N_16310,N_16902);
nor U17609 (N_17609,N_16390,N_16695);
nor U17610 (N_17610,N_16027,N_16003);
xor U17611 (N_17611,N_16239,N_16923);
nand U17612 (N_17612,N_16340,N_16979);
nand U17613 (N_17613,N_16569,N_16182);
nand U17614 (N_17614,N_16733,N_16319);
nor U17615 (N_17615,N_16017,N_16835);
or U17616 (N_17616,N_16310,N_16247);
xor U17617 (N_17617,N_16274,N_16316);
and U17618 (N_17618,N_16921,N_16732);
nor U17619 (N_17619,N_16543,N_16377);
xnor U17620 (N_17620,N_16757,N_16679);
and U17621 (N_17621,N_16400,N_16857);
xnor U17622 (N_17622,N_16784,N_16291);
nor U17623 (N_17623,N_16705,N_16987);
or U17624 (N_17624,N_16541,N_16811);
nor U17625 (N_17625,N_16240,N_16531);
and U17626 (N_17626,N_16674,N_16141);
or U17627 (N_17627,N_16326,N_16797);
xnor U17628 (N_17628,N_16613,N_16713);
xor U17629 (N_17629,N_16163,N_16685);
or U17630 (N_17630,N_16107,N_16913);
xor U17631 (N_17631,N_16380,N_16882);
xor U17632 (N_17632,N_16012,N_16975);
and U17633 (N_17633,N_16846,N_16225);
and U17634 (N_17634,N_16054,N_16371);
nor U17635 (N_17635,N_16959,N_16539);
nor U17636 (N_17636,N_16098,N_16477);
or U17637 (N_17637,N_16440,N_16395);
xor U17638 (N_17638,N_16697,N_16865);
xor U17639 (N_17639,N_16421,N_16525);
or U17640 (N_17640,N_16058,N_16700);
and U17641 (N_17641,N_16898,N_16276);
and U17642 (N_17642,N_16780,N_16517);
xor U17643 (N_17643,N_16867,N_16831);
nor U17644 (N_17644,N_16078,N_16961);
or U17645 (N_17645,N_16802,N_16669);
nor U17646 (N_17646,N_16406,N_16190);
and U17647 (N_17647,N_16710,N_16665);
xnor U17648 (N_17648,N_16107,N_16528);
or U17649 (N_17649,N_16872,N_16400);
xor U17650 (N_17650,N_16367,N_16076);
xor U17651 (N_17651,N_16802,N_16321);
or U17652 (N_17652,N_16673,N_16062);
nor U17653 (N_17653,N_16091,N_16858);
and U17654 (N_17654,N_16489,N_16367);
nor U17655 (N_17655,N_16148,N_16683);
nor U17656 (N_17656,N_16280,N_16303);
and U17657 (N_17657,N_16240,N_16144);
and U17658 (N_17658,N_16526,N_16373);
xor U17659 (N_17659,N_16813,N_16797);
xor U17660 (N_17660,N_16733,N_16798);
and U17661 (N_17661,N_16361,N_16866);
nor U17662 (N_17662,N_16917,N_16452);
xor U17663 (N_17663,N_16508,N_16980);
xor U17664 (N_17664,N_16210,N_16709);
nor U17665 (N_17665,N_16760,N_16457);
or U17666 (N_17666,N_16691,N_16121);
nand U17667 (N_17667,N_16187,N_16961);
xor U17668 (N_17668,N_16941,N_16236);
nor U17669 (N_17669,N_16715,N_16947);
xor U17670 (N_17670,N_16294,N_16754);
and U17671 (N_17671,N_16957,N_16875);
nor U17672 (N_17672,N_16126,N_16983);
xor U17673 (N_17673,N_16544,N_16485);
nor U17674 (N_17674,N_16946,N_16492);
or U17675 (N_17675,N_16806,N_16009);
or U17676 (N_17676,N_16395,N_16993);
or U17677 (N_17677,N_16653,N_16885);
nand U17678 (N_17678,N_16431,N_16360);
nor U17679 (N_17679,N_16064,N_16913);
nor U17680 (N_17680,N_16350,N_16015);
nor U17681 (N_17681,N_16286,N_16823);
xnor U17682 (N_17682,N_16288,N_16235);
nand U17683 (N_17683,N_16766,N_16153);
or U17684 (N_17684,N_16887,N_16106);
nand U17685 (N_17685,N_16210,N_16775);
and U17686 (N_17686,N_16346,N_16188);
and U17687 (N_17687,N_16785,N_16176);
and U17688 (N_17688,N_16867,N_16302);
nor U17689 (N_17689,N_16740,N_16686);
nand U17690 (N_17690,N_16241,N_16597);
nand U17691 (N_17691,N_16130,N_16492);
or U17692 (N_17692,N_16480,N_16932);
xnor U17693 (N_17693,N_16156,N_16304);
nor U17694 (N_17694,N_16161,N_16824);
and U17695 (N_17695,N_16678,N_16585);
nor U17696 (N_17696,N_16217,N_16956);
nor U17697 (N_17697,N_16642,N_16254);
nor U17698 (N_17698,N_16444,N_16717);
or U17699 (N_17699,N_16386,N_16726);
nand U17700 (N_17700,N_16898,N_16158);
nand U17701 (N_17701,N_16713,N_16844);
or U17702 (N_17702,N_16589,N_16176);
nor U17703 (N_17703,N_16539,N_16560);
or U17704 (N_17704,N_16451,N_16020);
and U17705 (N_17705,N_16362,N_16949);
and U17706 (N_17706,N_16625,N_16270);
and U17707 (N_17707,N_16456,N_16648);
xor U17708 (N_17708,N_16199,N_16784);
xor U17709 (N_17709,N_16981,N_16742);
or U17710 (N_17710,N_16968,N_16638);
nor U17711 (N_17711,N_16860,N_16984);
xor U17712 (N_17712,N_16121,N_16231);
nand U17713 (N_17713,N_16779,N_16379);
and U17714 (N_17714,N_16654,N_16124);
or U17715 (N_17715,N_16213,N_16193);
nand U17716 (N_17716,N_16377,N_16915);
nor U17717 (N_17717,N_16703,N_16695);
xor U17718 (N_17718,N_16499,N_16594);
nand U17719 (N_17719,N_16218,N_16890);
and U17720 (N_17720,N_16284,N_16747);
xor U17721 (N_17721,N_16492,N_16368);
and U17722 (N_17722,N_16228,N_16814);
nor U17723 (N_17723,N_16353,N_16920);
and U17724 (N_17724,N_16835,N_16155);
and U17725 (N_17725,N_16205,N_16049);
xnor U17726 (N_17726,N_16615,N_16811);
and U17727 (N_17727,N_16080,N_16913);
nor U17728 (N_17728,N_16205,N_16328);
nor U17729 (N_17729,N_16950,N_16635);
xnor U17730 (N_17730,N_16751,N_16859);
and U17731 (N_17731,N_16663,N_16924);
and U17732 (N_17732,N_16072,N_16775);
and U17733 (N_17733,N_16113,N_16059);
nand U17734 (N_17734,N_16795,N_16676);
and U17735 (N_17735,N_16213,N_16677);
xnor U17736 (N_17736,N_16491,N_16395);
nand U17737 (N_17737,N_16672,N_16490);
and U17738 (N_17738,N_16655,N_16004);
or U17739 (N_17739,N_16339,N_16035);
or U17740 (N_17740,N_16046,N_16366);
xnor U17741 (N_17741,N_16162,N_16079);
xor U17742 (N_17742,N_16466,N_16344);
nor U17743 (N_17743,N_16269,N_16330);
and U17744 (N_17744,N_16326,N_16606);
and U17745 (N_17745,N_16731,N_16349);
and U17746 (N_17746,N_16300,N_16403);
nand U17747 (N_17747,N_16338,N_16777);
and U17748 (N_17748,N_16053,N_16709);
or U17749 (N_17749,N_16644,N_16530);
nor U17750 (N_17750,N_16573,N_16169);
and U17751 (N_17751,N_16190,N_16814);
or U17752 (N_17752,N_16488,N_16003);
nand U17753 (N_17753,N_16085,N_16240);
nor U17754 (N_17754,N_16113,N_16532);
and U17755 (N_17755,N_16029,N_16840);
and U17756 (N_17756,N_16944,N_16998);
xnor U17757 (N_17757,N_16317,N_16840);
xor U17758 (N_17758,N_16162,N_16749);
nand U17759 (N_17759,N_16436,N_16077);
nor U17760 (N_17760,N_16810,N_16585);
or U17761 (N_17761,N_16609,N_16824);
and U17762 (N_17762,N_16600,N_16675);
nand U17763 (N_17763,N_16073,N_16516);
xnor U17764 (N_17764,N_16171,N_16322);
nor U17765 (N_17765,N_16204,N_16707);
nand U17766 (N_17766,N_16492,N_16772);
nand U17767 (N_17767,N_16430,N_16265);
nand U17768 (N_17768,N_16632,N_16200);
and U17769 (N_17769,N_16253,N_16609);
nor U17770 (N_17770,N_16120,N_16181);
xor U17771 (N_17771,N_16836,N_16165);
or U17772 (N_17772,N_16963,N_16722);
nand U17773 (N_17773,N_16795,N_16013);
nor U17774 (N_17774,N_16125,N_16137);
or U17775 (N_17775,N_16273,N_16196);
and U17776 (N_17776,N_16954,N_16544);
or U17777 (N_17777,N_16843,N_16352);
xnor U17778 (N_17778,N_16665,N_16045);
nand U17779 (N_17779,N_16498,N_16643);
or U17780 (N_17780,N_16223,N_16885);
nand U17781 (N_17781,N_16529,N_16626);
nor U17782 (N_17782,N_16605,N_16123);
or U17783 (N_17783,N_16139,N_16057);
xnor U17784 (N_17784,N_16160,N_16893);
nand U17785 (N_17785,N_16326,N_16580);
or U17786 (N_17786,N_16288,N_16930);
nor U17787 (N_17787,N_16750,N_16744);
or U17788 (N_17788,N_16532,N_16902);
nor U17789 (N_17789,N_16920,N_16405);
and U17790 (N_17790,N_16728,N_16848);
or U17791 (N_17791,N_16474,N_16626);
nor U17792 (N_17792,N_16515,N_16747);
xnor U17793 (N_17793,N_16167,N_16032);
or U17794 (N_17794,N_16313,N_16066);
or U17795 (N_17795,N_16756,N_16291);
nand U17796 (N_17796,N_16273,N_16500);
and U17797 (N_17797,N_16133,N_16245);
nor U17798 (N_17798,N_16084,N_16154);
xor U17799 (N_17799,N_16897,N_16630);
nor U17800 (N_17800,N_16581,N_16062);
nor U17801 (N_17801,N_16246,N_16024);
or U17802 (N_17802,N_16659,N_16693);
or U17803 (N_17803,N_16421,N_16176);
or U17804 (N_17804,N_16339,N_16259);
xnor U17805 (N_17805,N_16628,N_16673);
or U17806 (N_17806,N_16630,N_16386);
and U17807 (N_17807,N_16702,N_16677);
and U17808 (N_17808,N_16975,N_16567);
and U17809 (N_17809,N_16273,N_16334);
xnor U17810 (N_17810,N_16404,N_16350);
nor U17811 (N_17811,N_16065,N_16360);
xnor U17812 (N_17812,N_16044,N_16642);
or U17813 (N_17813,N_16224,N_16209);
xnor U17814 (N_17814,N_16978,N_16895);
nand U17815 (N_17815,N_16807,N_16277);
xnor U17816 (N_17816,N_16494,N_16388);
xnor U17817 (N_17817,N_16145,N_16082);
nand U17818 (N_17818,N_16764,N_16916);
nor U17819 (N_17819,N_16920,N_16518);
xor U17820 (N_17820,N_16852,N_16423);
or U17821 (N_17821,N_16669,N_16147);
or U17822 (N_17822,N_16151,N_16300);
xnor U17823 (N_17823,N_16827,N_16394);
and U17824 (N_17824,N_16529,N_16216);
or U17825 (N_17825,N_16692,N_16040);
nand U17826 (N_17826,N_16863,N_16445);
nand U17827 (N_17827,N_16807,N_16232);
and U17828 (N_17828,N_16841,N_16542);
or U17829 (N_17829,N_16326,N_16871);
xor U17830 (N_17830,N_16393,N_16333);
nand U17831 (N_17831,N_16968,N_16311);
nand U17832 (N_17832,N_16964,N_16644);
nor U17833 (N_17833,N_16872,N_16810);
xor U17834 (N_17834,N_16237,N_16483);
and U17835 (N_17835,N_16447,N_16443);
nor U17836 (N_17836,N_16663,N_16094);
nor U17837 (N_17837,N_16715,N_16604);
or U17838 (N_17838,N_16478,N_16876);
nor U17839 (N_17839,N_16069,N_16362);
and U17840 (N_17840,N_16432,N_16201);
xor U17841 (N_17841,N_16206,N_16231);
xnor U17842 (N_17842,N_16938,N_16668);
nand U17843 (N_17843,N_16055,N_16915);
xor U17844 (N_17844,N_16421,N_16511);
nand U17845 (N_17845,N_16028,N_16845);
or U17846 (N_17846,N_16783,N_16344);
and U17847 (N_17847,N_16574,N_16587);
or U17848 (N_17848,N_16002,N_16036);
xor U17849 (N_17849,N_16608,N_16830);
nor U17850 (N_17850,N_16142,N_16902);
nand U17851 (N_17851,N_16603,N_16482);
nor U17852 (N_17852,N_16646,N_16759);
and U17853 (N_17853,N_16626,N_16262);
nor U17854 (N_17854,N_16737,N_16942);
and U17855 (N_17855,N_16241,N_16455);
and U17856 (N_17856,N_16110,N_16229);
and U17857 (N_17857,N_16690,N_16479);
nor U17858 (N_17858,N_16863,N_16666);
xnor U17859 (N_17859,N_16530,N_16251);
and U17860 (N_17860,N_16687,N_16877);
nor U17861 (N_17861,N_16687,N_16980);
nand U17862 (N_17862,N_16337,N_16414);
xnor U17863 (N_17863,N_16816,N_16834);
nor U17864 (N_17864,N_16611,N_16312);
xor U17865 (N_17865,N_16116,N_16193);
nand U17866 (N_17866,N_16360,N_16335);
and U17867 (N_17867,N_16045,N_16933);
xor U17868 (N_17868,N_16617,N_16212);
xor U17869 (N_17869,N_16167,N_16139);
nand U17870 (N_17870,N_16133,N_16539);
nor U17871 (N_17871,N_16715,N_16143);
and U17872 (N_17872,N_16499,N_16469);
nand U17873 (N_17873,N_16902,N_16908);
nor U17874 (N_17874,N_16776,N_16351);
nand U17875 (N_17875,N_16782,N_16409);
and U17876 (N_17876,N_16850,N_16217);
nor U17877 (N_17877,N_16732,N_16930);
nor U17878 (N_17878,N_16784,N_16975);
or U17879 (N_17879,N_16809,N_16570);
nand U17880 (N_17880,N_16753,N_16320);
and U17881 (N_17881,N_16466,N_16513);
nand U17882 (N_17882,N_16626,N_16402);
nand U17883 (N_17883,N_16562,N_16451);
or U17884 (N_17884,N_16784,N_16404);
nand U17885 (N_17885,N_16665,N_16043);
xor U17886 (N_17886,N_16613,N_16909);
and U17887 (N_17887,N_16096,N_16354);
nor U17888 (N_17888,N_16424,N_16408);
nand U17889 (N_17889,N_16836,N_16882);
nor U17890 (N_17890,N_16461,N_16052);
xnor U17891 (N_17891,N_16629,N_16697);
or U17892 (N_17892,N_16480,N_16703);
nor U17893 (N_17893,N_16176,N_16932);
nor U17894 (N_17894,N_16302,N_16426);
xnor U17895 (N_17895,N_16327,N_16094);
nor U17896 (N_17896,N_16085,N_16942);
xnor U17897 (N_17897,N_16030,N_16870);
xnor U17898 (N_17898,N_16585,N_16380);
nand U17899 (N_17899,N_16930,N_16681);
or U17900 (N_17900,N_16643,N_16663);
nor U17901 (N_17901,N_16348,N_16651);
xor U17902 (N_17902,N_16809,N_16178);
xnor U17903 (N_17903,N_16367,N_16788);
nand U17904 (N_17904,N_16270,N_16124);
xnor U17905 (N_17905,N_16630,N_16593);
nor U17906 (N_17906,N_16606,N_16697);
nor U17907 (N_17907,N_16994,N_16520);
xnor U17908 (N_17908,N_16172,N_16698);
nand U17909 (N_17909,N_16282,N_16264);
nand U17910 (N_17910,N_16883,N_16823);
nor U17911 (N_17911,N_16921,N_16556);
and U17912 (N_17912,N_16374,N_16527);
nand U17913 (N_17913,N_16148,N_16969);
nor U17914 (N_17914,N_16469,N_16707);
nor U17915 (N_17915,N_16704,N_16787);
xor U17916 (N_17916,N_16730,N_16310);
nand U17917 (N_17917,N_16783,N_16739);
nor U17918 (N_17918,N_16343,N_16455);
or U17919 (N_17919,N_16131,N_16912);
nand U17920 (N_17920,N_16535,N_16844);
nand U17921 (N_17921,N_16037,N_16221);
and U17922 (N_17922,N_16874,N_16013);
nand U17923 (N_17923,N_16876,N_16403);
nor U17924 (N_17924,N_16280,N_16688);
or U17925 (N_17925,N_16882,N_16581);
and U17926 (N_17926,N_16683,N_16338);
nand U17927 (N_17927,N_16938,N_16660);
nor U17928 (N_17928,N_16951,N_16189);
xnor U17929 (N_17929,N_16563,N_16962);
xnor U17930 (N_17930,N_16911,N_16595);
xnor U17931 (N_17931,N_16528,N_16658);
or U17932 (N_17932,N_16336,N_16164);
and U17933 (N_17933,N_16307,N_16900);
and U17934 (N_17934,N_16294,N_16271);
xnor U17935 (N_17935,N_16927,N_16566);
and U17936 (N_17936,N_16231,N_16323);
nand U17937 (N_17937,N_16138,N_16285);
or U17938 (N_17938,N_16568,N_16557);
nand U17939 (N_17939,N_16953,N_16338);
nand U17940 (N_17940,N_16054,N_16441);
nor U17941 (N_17941,N_16453,N_16438);
or U17942 (N_17942,N_16196,N_16589);
nor U17943 (N_17943,N_16459,N_16314);
xor U17944 (N_17944,N_16012,N_16426);
xor U17945 (N_17945,N_16778,N_16798);
or U17946 (N_17946,N_16206,N_16092);
and U17947 (N_17947,N_16620,N_16501);
or U17948 (N_17948,N_16469,N_16928);
or U17949 (N_17949,N_16651,N_16429);
xor U17950 (N_17950,N_16222,N_16434);
xor U17951 (N_17951,N_16441,N_16517);
xor U17952 (N_17952,N_16689,N_16573);
and U17953 (N_17953,N_16705,N_16506);
and U17954 (N_17954,N_16047,N_16984);
and U17955 (N_17955,N_16093,N_16761);
and U17956 (N_17956,N_16159,N_16823);
or U17957 (N_17957,N_16069,N_16008);
nor U17958 (N_17958,N_16124,N_16572);
and U17959 (N_17959,N_16940,N_16920);
xnor U17960 (N_17960,N_16765,N_16219);
xor U17961 (N_17961,N_16927,N_16485);
nor U17962 (N_17962,N_16477,N_16069);
xnor U17963 (N_17963,N_16231,N_16957);
nor U17964 (N_17964,N_16547,N_16529);
or U17965 (N_17965,N_16321,N_16366);
xnor U17966 (N_17966,N_16001,N_16250);
xnor U17967 (N_17967,N_16657,N_16243);
nor U17968 (N_17968,N_16872,N_16133);
nand U17969 (N_17969,N_16516,N_16666);
nor U17970 (N_17970,N_16151,N_16552);
and U17971 (N_17971,N_16150,N_16407);
nand U17972 (N_17972,N_16540,N_16240);
and U17973 (N_17973,N_16888,N_16197);
nand U17974 (N_17974,N_16975,N_16484);
or U17975 (N_17975,N_16815,N_16692);
or U17976 (N_17976,N_16002,N_16184);
and U17977 (N_17977,N_16169,N_16641);
nor U17978 (N_17978,N_16938,N_16708);
xnor U17979 (N_17979,N_16494,N_16330);
nand U17980 (N_17980,N_16095,N_16720);
and U17981 (N_17981,N_16917,N_16417);
xor U17982 (N_17982,N_16888,N_16758);
nor U17983 (N_17983,N_16209,N_16167);
or U17984 (N_17984,N_16626,N_16013);
nand U17985 (N_17985,N_16428,N_16213);
xor U17986 (N_17986,N_16819,N_16991);
or U17987 (N_17987,N_16047,N_16746);
nand U17988 (N_17988,N_16961,N_16100);
nand U17989 (N_17989,N_16695,N_16528);
nand U17990 (N_17990,N_16223,N_16363);
and U17991 (N_17991,N_16310,N_16723);
nor U17992 (N_17992,N_16387,N_16640);
and U17993 (N_17993,N_16879,N_16285);
nor U17994 (N_17994,N_16347,N_16329);
nor U17995 (N_17995,N_16380,N_16017);
nand U17996 (N_17996,N_16859,N_16829);
or U17997 (N_17997,N_16842,N_16747);
nand U17998 (N_17998,N_16702,N_16471);
and U17999 (N_17999,N_16586,N_16650);
nor U18000 (N_18000,N_17954,N_17540);
nor U18001 (N_18001,N_17375,N_17413);
nor U18002 (N_18002,N_17192,N_17275);
and U18003 (N_18003,N_17218,N_17877);
xnor U18004 (N_18004,N_17497,N_17755);
and U18005 (N_18005,N_17743,N_17258);
or U18006 (N_18006,N_17080,N_17582);
and U18007 (N_18007,N_17622,N_17821);
and U18008 (N_18008,N_17443,N_17051);
nand U18009 (N_18009,N_17974,N_17912);
xnor U18010 (N_18010,N_17179,N_17641);
nand U18011 (N_18011,N_17826,N_17099);
nor U18012 (N_18012,N_17868,N_17549);
and U18013 (N_18013,N_17160,N_17469);
nor U18014 (N_18014,N_17955,N_17085);
and U18015 (N_18015,N_17007,N_17617);
xor U18016 (N_18016,N_17405,N_17283);
and U18017 (N_18017,N_17168,N_17410);
xnor U18018 (N_18018,N_17020,N_17752);
nand U18019 (N_18019,N_17625,N_17013);
or U18020 (N_18020,N_17914,N_17562);
xor U18021 (N_18021,N_17980,N_17344);
and U18022 (N_18022,N_17543,N_17606);
nand U18023 (N_18023,N_17418,N_17044);
nand U18024 (N_18024,N_17873,N_17399);
and U18025 (N_18025,N_17411,N_17573);
nor U18026 (N_18026,N_17175,N_17639);
nor U18027 (N_18027,N_17255,N_17857);
nor U18028 (N_18028,N_17629,N_17789);
nor U18029 (N_18029,N_17198,N_17377);
nor U18030 (N_18030,N_17651,N_17815);
and U18031 (N_18031,N_17546,N_17057);
nand U18032 (N_18032,N_17662,N_17668);
nor U18033 (N_18033,N_17503,N_17822);
nor U18034 (N_18034,N_17227,N_17016);
or U18035 (N_18035,N_17456,N_17769);
and U18036 (N_18036,N_17680,N_17450);
nor U18037 (N_18037,N_17539,N_17446);
nor U18038 (N_18038,N_17706,N_17626);
or U18039 (N_18039,N_17087,N_17196);
nand U18040 (N_18040,N_17913,N_17674);
and U18041 (N_18041,N_17833,N_17048);
xnor U18042 (N_18042,N_17829,N_17421);
or U18043 (N_18043,N_17766,N_17261);
or U18044 (N_18044,N_17654,N_17378);
nand U18045 (N_18045,N_17118,N_17270);
and U18046 (N_18046,N_17817,N_17334);
nand U18047 (N_18047,N_17983,N_17849);
and U18048 (N_18048,N_17730,N_17447);
or U18049 (N_18049,N_17145,N_17478);
or U18050 (N_18050,N_17844,N_17104);
or U18051 (N_18051,N_17870,N_17733);
nand U18052 (N_18052,N_17551,N_17116);
and U18053 (N_18053,N_17262,N_17157);
and U18054 (N_18054,N_17343,N_17757);
nor U18055 (N_18055,N_17468,N_17357);
nand U18056 (N_18056,N_17881,N_17216);
xor U18057 (N_18057,N_17796,N_17664);
and U18058 (N_18058,N_17265,N_17222);
xnor U18059 (N_18059,N_17150,N_17990);
and U18060 (N_18060,N_17441,N_17217);
nand U18061 (N_18061,N_17461,N_17337);
nand U18062 (N_18062,N_17518,N_17591);
xor U18063 (N_18063,N_17322,N_17548);
and U18064 (N_18064,N_17074,N_17507);
and U18065 (N_18065,N_17071,N_17864);
nor U18066 (N_18066,N_17713,N_17311);
nor U18067 (N_18067,N_17612,N_17678);
nand U18068 (N_18068,N_17891,N_17184);
xnor U18069 (N_18069,N_17679,N_17351);
or U18070 (N_18070,N_17519,N_17962);
and U18071 (N_18071,N_17723,N_17021);
or U18072 (N_18072,N_17401,N_17472);
xnor U18073 (N_18073,N_17950,N_17008);
nor U18074 (N_18074,N_17001,N_17092);
or U18075 (N_18075,N_17395,N_17896);
xor U18076 (N_18076,N_17906,N_17177);
nor U18077 (N_18077,N_17560,N_17717);
nor U18078 (N_18078,N_17928,N_17598);
or U18079 (N_18079,N_17874,N_17783);
nor U18080 (N_18080,N_17956,N_17957);
and U18081 (N_18081,N_17508,N_17657);
or U18082 (N_18082,N_17326,N_17088);
and U18083 (N_18083,N_17075,N_17635);
or U18084 (N_18084,N_17512,N_17267);
and U18085 (N_18085,N_17424,N_17510);
xnor U18086 (N_18086,N_17702,N_17155);
nor U18087 (N_18087,N_17046,N_17439);
xnor U18088 (N_18088,N_17566,N_17091);
or U18089 (N_18089,N_17537,N_17797);
nor U18090 (N_18090,N_17333,N_17368);
xor U18091 (N_18091,N_17644,N_17941);
or U18092 (N_18092,N_17047,N_17762);
or U18093 (N_18093,N_17340,N_17787);
nand U18094 (N_18094,N_17727,N_17388);
nor U18095 (N_18095,N_17522,N_17908);
nor U18096 (N_18096,N_17670,N_17187);
nand U18097 (N_18097,N_17367,N_17393);
or U18098 (N_18098,N_17581,N_17299);
and U18099 (N_18099,N_17785,N_17136);
nand U18100 (N_18100,N_17305,N_17526);
and U18101 (N_18101,N_17922,N_17176);
xnor U18102 (N_18102,N_17200,N_17193);
xnor U18103 (N_18103,N_17223,N_17294);
and U18104 (N_18104,N_17704,N_17675);
and U18105 (N_18105,N_17023,N_17824);
nor U18106 (N_18106,N_17746,N_17452);
xnor U18107 (N_18107,N_17930,N_17404);
nand U18108 (N_18108,N_17454,N_17570);
and U18109 (N_18109,N_17676,N_17542);
nor U18110 (N_18110,N_17127,N_17940);
and U18111 (N_18111,N_17319,N_17105);
nand U18112 (N_18112,N_17620,N_17342);
xnor U18113 (N_18113,N_17332,N_17135);
xor U18114 (N_18114,N_17805,N_17103);
nor U18115 (N_18115,N_17114,N_17987);
and U18116 (N_18116,N_17627,N_17649);
or U18117 (N_18117,N_17521,N_17171);
xnor U18118 (N_18118,N_17500,N_17655);
or U18119 (N_18119,N_17030,N_17807);
xor U18120 (N_18120,N_17100,N_17451);
and U18121 (N_18121,N_17005,N_17281);
nor U18122 (N_18122,N_17673,N_17584);
nor U18123 (N_18123,N_17455,N_17055);
xor U18124 (N_18124,N_17580,N_17861);
nor U18125 (N_18125,N_17967,N_17583);
xnor U18126 (N_18126,N_17169,N_17414);
nor U18127 (N_18127,N_17671,N_17130);
xor U18128 (N_18128,N_17939,N_17489);
xnor U18129 (N_18129,N_17603,N_17384);
xnor U18130 (N_18130,N_17541,N_17473);
nand U18131 (N_18131,N_17068,N_17613);
nand U18132 (N_18132,N_17856,N_17318);
nor U18133 (N_18133,N_17205,N_17736);
and U18134 (N_18134,N_17061,N_17231);
nand U18135 (N_18135,N_17009,N_17398);
xnor U18136 (N_18136,N_17709,N_17277);
xnor U18137 (N_18137,N_17475,N_17308);
and U18138 (N_18138,N_17089,N_17616);
nand U18139 (N_18139,N_17741,N_17827);
xor U18140 (N_18140,N_17098,N_17365);
xnor U18141 (N_18141,N_17535,N_17210);
nor U18142 (N_18142,N_17499,N_17372);
or U18143 (N_18143,N_17937,N_17031);
xnor U18144 (N_18144,N_17213,N_17250);
and U18145 (N_18145,N_17683,N_17381);
or U18146 (N_18146,N_17120,N_17350);
xor U18147 (N_18147,N_17872,N_17689);
or U18148 (N_18148,N_17772,N_17840);
and U18149 (N_18149,N_17828,N_17324);
xor U18150 (N_18150,N_17920,N_17970);
xor U18151 (N_18151,N_17911,N_17793);
and U18152 (N_18152,N_17645,N_17558);
and U18153 (N_18153,N_17385,N_17776);
nor U18154 (N_18154,N_17491,N_17533);
xor U18155 (N_18155,N_17137,N_17093);
nor U18156 (N_18156,N_17747,N_17686);
nor U18157 (N_18157,N_17909,N_17492);
xnor U18158 (N_18158,N_17076,N_17520);
xor U18159 (N_18159,N_17180,N_17285);
nand U18160 (N_18160,N_17585,N_17147);
xnor U18161 (N_18161,N_17479,N_17630);
nand U18162 (N_18162,N_17524,N_17208);
and U18163 (N_18163,N_17316,N_17938);
and U18164 (N_18164,N_17079,N_17434);
and U18165 (N_18165,N_17910,N_17437);
nand U18166 (N_18166,N_17483,N_17391);
or U18167 (N_18167,N_17774,N_17237);
nand U18168 (N_18168,N_17315,N_17495);
and U18169 (N_18169,N_17597,N_17442);
nor U18170 (N_18170,N_17360,N_17345);
xor U18171 (N_18171,N_17715,N_17049);
nor U18172 (N_18172,N_17677,N_17515);
and U18173 (N_18173,N_17219,N_17808);
nor U18174 (N_18174,N_17988,N_17975);
xor U18175 (N_18175,N_17790,N_17428);
nor U18176 (N_18176,N_17719,N_17595);
nor U18177 (N_18177,N_17292,N_17830);
xor U18178 (N_18178,N_17392,N_17396);
or U18179 (N_18179,N_17040,N_17062);
or U18180 (N_18180,N_17601,N_17588);
and U18181 (N_18181,N_17382,N_17471);
and U18182 (N_18182,N_17027,N_17904);
nor U18183 (N_18183,N_17720,N_17667);
and U18184 (N_18184,N_17209,N_17780);
or U18185 (N_18185,N_17138,N_17972);
nor U18186 (N_18186,N_17467,N_17331);
and U18187 (N_18187,N_17965,N_17813);
nand U18188 (N_18188,N_17577,N_17660);
nor U18189 (N_18189,N_17435,N_17036);
xor U18190 (N_18190,N_17317,N_17514);
nand U18191 (N_18191,N_17681,N_17876);
or U18192 (N_18192,N_17905,N_17899);
nand U18193 (N_18193,N_17221,N_17786);
nand U18194 (N_18194,N_17893,N_17614);
or U18195 (N_18195,N_17672,N_17353);
and U18196 (N_18196,N_17430,N_17665);
xnor U18197 (N_18197,N_17571,N_17059);
xnor U18198 (N_18198,N_17724,N_17482);
nor U18199 (N_18199,N_17569,N_17148);
and U18200 (N_18200,N_17532,N_17274);
or U18201 (N_18201,N_17761,N_17457);
or U18202 (N_18202,N_17341,N_17273);
or U18203 (N_18203,N_17778,N_17431);
nor U18204 (N_18204,N_17504,N_17712);
nor U18205 (N_18205,N_17971,N_17167);
nor U18206 (N_18206,N_17470,N_17642);
or U18207 (N_18207,N_17403,N_17096);
or U18208 (N_18208,N_17149,N_17948);
and U18209 (N_18209,N_17860,N_17942);
xor U18210 (N_18210,N_17271,N_17146);
or U18211 (N_18211,N_17758,N_17996);
and U18212 (N_18212,N_17890,N_17550);
nand U18213 (N_18213,N_17698,N_17234);
or U18214 (N_18214,N_17090,N_17015);
or U18215 (N_18215,N_17511,N_17125);
nand U18216 (N_18216,N_17944,N_17043);
and U18217 (N_18217,N_17767,N_17081);
nor U18218 (N_18218,N_17230,N_17918);
or U18219 (N_18219,N_17014,N_17831);
or U18220 (N_18220,N_17916,N_17599);
or U18221 (N_18221,N_17352,N_17835);
nand U18222 (N_18222,N_17108,N_17017);
or U18223 (N_18223,N_17244,N_17211);
nand U18224 (N_18224,N_17576,N_17336);
nand U18225 (N_18225,N_17379,N_17634);
xor U18226 (N_18226,N_17459,N_17658);
nor U18227 (N_18227,N_17369,N_17509);
nand U18228 (N_18228,N_17530,N_17409);
xnor U18229 (N_18229,N_17124,N_17764);
nor U18230 (N_18230,N_17083,N_17838);
xor U18231 (N_18231,N_17084,N_17968);
xnor U18232 (N_18232,N_17628,N_17233);
and U18233 (N_18233,N_17820,N_17993);
or U18234 (N_18234,N_17842,N_17513);
and U18235 (N_18235,N_17763,N_17587);
nand U18236 (N_18236,N_17701,N_17376);
nor U18237 (N_18237,N_17552,N_17173);
and U18238 (N_18238,N_17812,N_17257);
and U18239 (N_18239,N_17888,N_17960);
xor U18240 (N_18240,N_17865,N_17185);
xor U18241 (N_18241,N_17033,N_17609);
nand U18242 (N_18242,N_17523,N_17128);
or U18243 (N_18243,N_17158,N_17374);
and U18244 (N_18244,N_17371,N_17024);
or U18245 (N_18245,N_17839,N_17029);
and U18246 (N_18246,N_17695,N_17416);
xnor U18247 (N_18247,N_17768,N_17314);
or U18248 (N_18248,N_17659,N_17339);
and U18249 (N_18249,N_17338,N_17982);
nand U18250 (N_18250,N_17915,N_17460);
and U18251 (N_18251,N_17973,N_17653);
nand U18252 (N_18252,N_17536,N_17754);
and U18253 (N_18253,N_17243,N_17879);
nand U18254 (N_18254,N_17791,N_17253);
and U18255 (N_18255,N_17624,N_17348);
nand U18256 (N_18256,N_17094,N_17117);
nand U18257 (N_18257,N_17992,N_17553);
or U18258 (N_18258,N_17214,N_17966);
or U18259 (N_18259,N_17517,N_17053);
nor U18260 (N_18260,N_17765,N_17189);
nand U18261 (N_18261,N_17528,N_17394);
nand U18262 (N_18262,N_17464,N_17263);
nand U18263 (N_18263,N_17364,N_17195);
nor U18264 (N_18264,N_17759,N_17887);
nand U18265 (N_18265,N_17929,N_17494);
nor U18266 (N_18266,N_17781,N_17837);
xnor U18267 (N_18267,N_17563,N_17480);
nor U18268 (N_18268,N_17919,N_17863);
or U18269 (N_18269,N_17711,N_17298);
and U18270 (N_18270,N_17567,N_17615);
or U18271 (N_18271,N_17306,N_17534);
xnor U18272 (N_18272,N_17788,N_17531);
nor U18273 (N_18273,N_17745,N_17538);
xnor U18274 (N_18274,N_17852,N_17354);
nand U18275 (N_18275,N_17438,N_17107);
xnor U18276 (N_18276,N_17985,N_17693);
or U18277 (N_18277,N_17356,N_17643);
or U18278 (N_18278,N_17449,N_17238);
or U18279 (N_18279,N_17433,N_17771);
xor U18280 (N_18280,N_17440,N_17203);
xnor U18281 (N_18281,N_17018,N_17153);
and U18282 (N_18282,N_17592,N_17760);
xnor U18283 (N_18283,N_17383,N_17363);
or U18284 (N_18284,N_17229,N_17697);
or U18285 (N_18285,N_17462,N_17402);
nor U18286 (N_18286,N_17307,N_17832);
xor U18287 (N_18287,N_17045,N_17802);
and U18288 (N_18288,N_17871,N_17026);
or U18289 (N_18289,N_17154,N_17917);
and U18290 (N_18290,N_17109,N_17481);
or U18291 (N_18291,N_17932,N_17429);
nand U18292 (N_18292,N_17002,N_17579);
nand U18293 (N_18293,N_17151,N_17739);
nand U18294 (N_18294,N_17818,N_17313);
nor U18295 (N_18295,N_17290,N_17346);
and U18296 (N_18296,N_17869,N_17907);
or U18297 (N_18297,N_17052,N_17798);
and U18298 (N_18298,N_17732,N_17997);
nand U18299 (N_18299,N_17728,N_17204);
xnor U18300 (N_18300,N_17115,N_17019);
and U18301 (N_18301,N_17705,N_17854);
nor U18302 (N_18302,N_17823,N_17964);
nor U18303 (N_18303,N_17923,N_17101);
nand U18304 (N_18304,N_17490,N_17846);
nand U18305 (N_18305,N_17493,N_17902);
nand U18306 (N_18306,N_17113,N_17848);
xnor U18307 (N_18307,N_17042,N_17162);
or U18308 (N_18308,N_17866,N_17183);
nand U18309 (N_18309,N_17465,N_17773);
nor U18310 (N_18310,N_17803,N_17633);
or U18311 (N_18311,N_17172,N_17436);
or U18312 (N_18312,N_17804,N_17792);
nand U18313 (N_18313,N_17359,N_17496);
nor U18314 (N_18314,N_17082,N_17097);
or U18315 (N_18315,N_17894,N_17845);
nand U18316 (N_18316,N_17684,N_17806);
nor U18317 (N_18317,N_17903,N_17235);
nand U18318 (N_18318,N_17448,N_17239);
and U18319 (N_18319,N_17279,N_17703);
nand U18320 (N_18320,N_17931,N_17420);
or U18321 (N_18321,N_17058,N_17999);
nor U18322 (N_18322,N_17199,N_17422);
nor U18323 (N_18323,N_17809,N_17035);
nor U18324 (N_18324,N_17925,N_17568);
and U18325 (N_18325,N_17529,N_17463);
nor U18326 (N_18326,N_17801,N_17112);
xor U18327 (N_18327,N_17882,N_17716);
nand U18328 (N_18328,N_17143,N_17132);
xnor U18329 (N_18329,N_17947,N_17086);
nor U18330 (N_18330,N_17557,N_17476);
and U18331 (N_18331,N_17004,N_17282);
or U18332 (N_18332,N_17445,N_17287);
nor U18333 (N_18333,N_17142,N_17687);
nand U18334 (N_18334,N_17190,N_17144);
nand U18335 (N_18335,N_17156,N_17301);
nor U18336 (N_18336,N_17330,N_17610);
or U18337 (N_18337,N_17400,N_17800);
xor U18338 (N_18338,N_17545,N_17123);
or U18339 (N_18339,N_17159,N_17725);
or U18340 (N_18340,N_17194,N_17819);
nor U18341 (N_18341,N_17900,N_17289);
or U18342 (N_18342,N_17564,N_17095);
or U18343 (N_18343,N_17181,N_17721);
and U18344 (N_18344,N_17961,N_17248);
nor U18345 (N_18345,N_17066,N_17119);
and U18346 (N_18346,N_17590,N_17296);
xnor U18347 (N_18347,N_17502,N_17370);
xor U18348 (N_18348,N_17025,N_17656);
and U18349 (N_18349,N_17544,N_17407);
xor U18350 (N_18350,N_17102,N_17249);
or U18351 (N_18351,N_17756,N_17225);
or U18352 (N_18352,N_17358,N_17106);
or U18353 (N_18353,N_17605,N_17892);
and U18354 (N_18354,N_17555,N_17858);
xor U18355 (N_18355,N_17995,N_17140);
nand U18356 (N_18356,N_17065,N_17751);
or U18357 (N_18357,N_17734,N_17782);
xnor U18358 (N_18358,N_17958,N_17748);
and U18359 (N_18359,N_17685,N_17050);
nand U18360 (N_18360,N_17886,N_17690);
and U18361 (N_18361,N_17278,N_17859);
and U18362 (N_18362,N_17166,N_17586);
nand U18363 (N_18363,N_17486,N_17742);
nor U18364 (N_18364,N_17959,N_17699);
or U18365 (N_18365,N_17423,N_17232);
xnor U18366 (N_18366,N_17898,N_17880);
or U18367 (N_18367,N_17623,N_17637);
nand U18368 (N_18368,N_17254,N_17600);
and U18369 (N_18369,N_17131,N_17740);
and U18370 (N_18370,N_17594,N_17867);
nor U18371 (N_18371,N_17197,N_17744);
xnor U18372 (N_18372,N_17295,N_17072);
xnor U18373 (N_18373,N_17133,N_17648);
xor U18374 (N_18374,N_17291,N_17260);
nand U18375 (N_18375,N_17700,N_17731);
or U18376 (N_18376,N_17366,N_17501);
xnor U18377 (N_18377,N_17386,N_17682);
nand U18378 (N_18378,N_17836,N_17264);
xor U18379 (N_18379,N_17206,N_17608);
or U18380 (N_18380,N_17012,N_17280);
or U18381 (N_18381,N_17269,N_17236);
or U18382 (N_18382,N_17795,N_17998);
xor U18383 (N_18383,N_17933,N_17220);
or U18384 (N_18384,N_17163,N_17485);
xnor U18385 (N_18385,N_17251,N_17161);
nor U18386 (N_18386,N_17506,N_17661);
nor U18387 (N_18387,N_17708,N_17994);
and U18388 (N_18388,N_17663,N_17256);
or U18389 (N_18389,N_17889,N_17621);
and U18390 (N_18390,N_17268,N_17978);
or U18391 (N_18391,N_17604,N_17390);
nand U18392 (N_18392,N_17729,N_17770);
xnor U18393 (N_18393,N_17070,N_17934);
or U18394 (N_18394,N_17943,N_17977);
nor U18395 (N_18395,N_17419,N_17293);
nand U18396 (N_18396,N_17589,N_17417);
and U18397 (N_18397,N_17714,N_17328);
and U18398 (N_18398,N_17885,N_17669);
xnor U18399 (N_18399,N_17111,N_17426);
nand U18400 (N_18400,N_17069,N_17963);
and U18401 (N_18401,N_17320,N_17215);
xor U18402 (N_18402,N_17191,N_17949);
and U18403 (N_18403,N_17735,N_17554);
xor U18404 (N_18404,N_17794,N_17458);
nand U18405 (N_18405,N_17811,N_17228);
or U18406 (N_18406,N_17067,N_17022);
xnor U18407 (N_18407,N_17945,N_17636);
xor U18408 (N_18408,N_17321,N_17139);
nand U18409 (N_18409,N_17387,N_17028);
or U18410 (N_18410,N_17777,N_17799);
nand U18411 (N_18411,N_17226,N_17559);
or U18412 (N_18412,N_17981,N_17924);
nand U18413 (N_18413,N_17814,N_17325);
xor U18414 (N_18414,N_17691,N_17129);
nor U18415 (N_18415,N_17056,N_17415);
and U18416 (N_18416,N_17037,N_17951);
xnor U18417 (N_18417,N_17241,N_17297);
nor U18418 (N_18418,N_17547,N_17516);
or U18419 (N_18419,N_17666,N_17561);
xor U18420 (N_18420,N_17272,N_17212);
xor U18421 (N_18421,N_17593,N_17991);
nor U18422 (N_18422,N_17989,N_17425);
nor U18423 (N_18423,N_17976,N_17309);
nand U18424 (N_18424,N_17578,N_17825);
nand U18425 (N_18425,N_17936,N_17259);
nand U18426 (N_18426,N_17722,N_17935);
nor U18427 (N_18427,N_17335,N_17477);
and U18428 (N_18428,N_17565,N_17304);
or U18429 (N_18429,N_17498,N_17810);
nand U18430 (N_18430,N_17572,N_17696);
and U18431 (N_18431,N_17134,N_17596);
nand U18432 (N_18432,N_17006,N_17726);
nor U18433 (N_18433,N_17753,N_17921);
nor U18434 (N_18434,N_17652,N_17389);
nand U18435 (N_18435,N_17895,N_17843);
nand U18436 (N_18436,N_17647,N_17631);
nor U18437 (N_18437,N_17484,N_17288);
nor U18438 (N_18438,N_17855,N_17174);
nor U18439 (N_18439,N_17850,N_17841);
or U18440 (N_18440,N_17060,N_17487);
nand U18441 (N_18441,N_17432,N_17003);
or U18442 (N_18442,N_17692,N_17718);
nor U18443 (N_18443,N_17505,N_17474);
or U18444 (N_18444,N_17064,N_17110);
and U18445 (N_18445,N_17884,N_17077);
and U18446 (N_18446,N_17862,N_17412);
or U18447 (N_18447,N_17312,N_17302);
xnor U18448 (N_18448,N_17323,N_17619);
xor U18449 (N_18449,N_17853,N_17611);
and U18450 (N_18450,N_17121,N_17284);
and U18451 (N_18451,N_17488,N_17041);
nor U18452 (N_18452,N_17640,N_17901);
xnor U18453 (N_18453,N_17245,N_17952);
xor U18454 (N_18454,N_17164,N_17073);
or U18455 (N_18455,N_17300,N_17707);
or U18456 (N_18456,N_17618,N_17926);
or U18457 (N_18457,N_17607,N_17953);
nand U18458 (N_18458,N_17240,N_17427);
or U18459 (N_18459,N_17775,N_17329);
nand U18460 (N_18460,N_17738,N_17038);
or U18461 (N_18461,N_17186,N_17303);
and U18462 (N_18462,N_17851,N_17397);
nand U18463 (N_18463,N_17946,N_17310);
nand U18464 (N_18464,N_17170,N_17406);
and U18465 (N_18465,N_17784,N_17034);
or U18466 (N_18466,N_17575,N_17638);
xnor U18467 (N_18467,N_17327,N_17266);
or U18468 (N_18468,N_17453,N_17347);
nand U18469 (N_18469,N_17246,N_17883);
or U18470 (N_18470,N_17032,N_17574);
and U18471 (N_18471,N_17373,N_17834);
nor U18472 (N_18472,N_17224,N_17063);
nor U18473 (N_18473,N_17779,N_17650);
or U18474 (N_18474,N_17078,N_17816);
and U18475 (N_18475,N_17750,N_17408);
and U18476 (N_18476,N_17525,N_17602);
and U18477 (N_18477,N_17152,N_17737);
and U18478 (N_18478,N_17749,N_17969);
xor U18479 (N_18479,N_17201,N_17182);
nor U18480 (N_18480,N_17361,N_17527);
xor U18481 (N_18481,N_17349,N_17878);
xnor U18482 (N_18482,N_17242,N_17362);
nor U18483 (N_18483,N_17380,N_17984);
nor U18484 (N_18484,N_17247,N_17556);
xnor U18485 (N_18485,N_17927,N_17444);
xor U18486 (N_18486,N_17054,N_17986);
and U18487 (N_18487,N_17286,N_17646);
or U18488 (N_18488,N_17165,N_17039);
nand U18489 (N_18489,N_17694,N_17178);
nor U18490 (N_18490,N_17979,N_17126);
nand U18491 (N_18491,N_17875,N_17010);
xnor U18492 (N_18492,N_17632,N_17207);
or U18493 (N_18493,N_17122,N_17252);
nor U18494 (N_18494,N_17688,N_17355);
or U18495 (N_18495,N_17276,N_17141);
xnor U18496 (N_18496,N_17188,N_17011);
or U18497 (N_18497,N_17847,N_17000);
nor U18498 (N_18498,N_17466,N_17897);
or U18499 (N_18499,N_17202,N_17710);
and U18500 (N_18500,N_17307,N_17856);
and U18501 (N_18501,N_17176,N_17492);
xnor U18502 (N_18502,N_17445,N_17921);
and U18503 (N_18503,N_17578,N_17537);
nand U18504 (N_18504,N_17988,N_17146);
or U18505 (N_18505,N_17026,N_17947);
and U18506 (N_18506,N_17584,N_17568);
and U18507 (N_18507,N_17523,N_17988);
xnor U18508 (N_18508,N_17738,N_17912);
xnor U18509 (N_18509,N_17669,N_17780);
nand U18510 (N_18510,N_17906,N_17495);
xnor U18511 (N_18511,N_17957,N_17636);
nand U18512 (N_18512,N_17183,N_17149);
or U18513 (N_18513,N_17357,N_17974);
and U18514 (N_18514,N_17313,N_17736);
or U18515 (N_18515,N_17343,N_17625);
or U18516 (N_18516,N_17510,N_17276);
xor U18517 (N_18517,N_17022,N_17336);
nand U18518 (N_18518,N_17545,N_17676);
nor U18519 (N_18519,N_17051,N_17845);
xnor U18520 (N_18520,N_17176,N_17110);
nand U18521 (N_18521,N_17740,N_17329);
nand U18522 (N_18522,N_17301,N_17925);
nand U18523 (N_18523,N_17665,N_17381);
xor U18524 (N_18524,N_17911,N_17453);
nand U18525 (N_18525,N_17668,N_17228);
nand U18526 (N_18526,N_17128,N_17116);
and U18527 (N_18527,N_17567,N_17017);
and U18528 (N_18528,N_17303,N_17053);
or U18529 (N_18529,N_17952,N_17351);
or U18530 (N_18530,N_17907,N_17510);
and U18531 (N_18531,N_17337,N_17693);
nand U18532 (N_18532,N_17177,N_17217);
xor U18533 (N_18533,N_17077,N_17769);
nor U18534 (N_18534,N_17644,N_17830);
xor U18535 (N_18535,N_17023,N_17933);
or U18536 (N_18536,N_17711,N_17659);
nor U18537 (N_18537,N_17986,N_17103);
and U18538 (N_18538,N_17800,N_17793);
xnor U18539 (N_18539,N_17588,N_17124);
xor U18540 (N_18540,N_17613,N_17773);
or U18541 (N_18541,N_17840,N_17922);
xor U18542 (N_18542,N_17103,N_17373);
nor U18543 (N_18543,N_17809,N_17231);
nand U18544 (N_18544,N_17024,N_17897);
nor U18545 (N_18545,N_17357,N_17593);
or U18546 (N_18546,N_17761,N_17010);
xnor U18547 (N_18547,N_17610,N_17847);
nand U18548 (N_18548,N_17693,N_17463);
nand U18549 (N_18549,N_17700,N_17594);
nor U18550 (N_18550,N_17322,N_17342);
or U18551 (N_18551,N_17117,N_17895);
and U18552 (N_18552,N_17801,N_17828);
and U18553 (N_18553,N_17946,N_17108);
or U18554 (N_18554,N_17853,N_17632);
nor U18555 (N_18555,N_17211,N_17479);
nand U18556 (N_18556,N_17044,N_17263);
nand U18557 (N_18557,N_17078,N_17824);
nor U18558 (N_18558,N_17952,N_17515);
or U18559 (N_18559,N_17131,N_17046);
nand U18560 (N_18560,N_17804,N_17615);
nor U18561 (N_18561,N_17089,N_17516);
nor U18562 (N_18562,N_17804,N_17825);
xor U18563 (N_18563,N_17006,N_17960);
nand U18564 (N_18564,N_17265,N_17245);
or U18565 (N_18565,N_17794,N_17571);
or U18566 (N_18566,N_17344,N_17599);
nand U18567 (N_18567,N_17510,N_17419);
nand U18568 (N_18568,N_17620,N_17358);
or U18569 (N_18569,N_17184,N_17360);
nor U18570 (N_18570,N_17403,N_17826);
and U18571 (N_18571,N_17387,N_17414);
and U18572 (N_18572,N_17438,N_17185);
xnor U18573 (N_18573,N_17381,N_17637);
nand U18574 (N_18574,N_17844,N_17317);
xnor U18575 (N_18575,N_17428,N_17314);
or U18576 (N_18576,N_17552,N_17121);
xnor U18577 (N_18577,N_17318,N_17391);
and U18578 (N_18578,N_17330,N_17563);
or U18579 (N_18579,N_17501,N_17809);
or U18580 (N_18580,N_17006,N_17669);
or U18581 (N_18581,N_17302,N_17948);
xor U18582 (N_18582,N_17191,N_17980);
nand U18583 (N_18583,N_17159,N_17959);
or U18584 (N_18584,N_17487,N_17458);
or U18585 (N_18585,N_17507,N_17185);
nor U18586 (N_18586,N_17746,N_17745);
or U18587 (N_18587,N_17177,N_17905);
nor U18588 (N_18588,N_17701,N_17089);
nand U18589 (N_18589,N_17672,N_17799);
nand U18590 (N_18590,N_17906,N_17714);
xor U18591 (N_18591,N_17830,N_17734);
and U18592 (N_18592,N_17366,N_17040);
xnor U18593 (N_18593,N_17729,N_17931);
nand U18594 (N_18594,N_17602,N_17121);
nor U18595 (N_18595,N_17470,N_17467);
nand U18596 (N_18596,N_17350,N_17689);
xnor U18597 (N_18597,N_17151,N_17847);
nor U18598 (N_18598,N_17564,N_17508);
xnor U18599 (N_18599,N_17658,N_17147);
and U18600 (N_18600,N_17729,N_17476);
nand U18601 (N_18601,N_17807,N_17225);
nand U18602 (N_18602,N_17207,N_17538);
xnor U18603 (N_18603,N_17978,N_17139);
nand U18604 (N_18604,N_17094,N_17619);
nor U18605 (N_18605,N_17206,N_17830);
and U18606 (N_18606,N_17151,N_17655);
or U18607 (N_18607,N_17753,N_17575);
xnor U18608 (N_18608,N_17049,N_17612);
nand U18609 (N_18609,N_17560,N_17365);
nor U18610 (N_18610,N_17395,N_17935);
nand U18611 (N_18611,N_17982,N_17813);
or U18612 (N_18612,N_17869,N_17331);
or U18613 (N_18613,N_17445,N_17346);
and U18614 (N_18614,N_17926,N_17923);
nand U18615 (N_18615,N_17913,N_17307);
nand U18616 (N_18616,N_17173,N_17546);
nand U18617 (N_18617,N_17080,N_17226);
xnor U18618 (N_18618,N_17933,N_17412);
and U18619 (N_18619,N_17679,N_17690);
or U18620 (N_18620,N_17711,N_17667);
nand U18621 (N_18621,N_17995,N_17863);
and U18622 (N_18622,N_17623,N_17493);
or U18623 (N_18623,N_17903,N_17470);
nand U18624 (N_18624,N_17558,N_17133);
xor U18625 (N_18625,N_17925,N_17142);
nor U18626 (N_18626,N_17402,N_17538);
xnor U18627 (N_18627,N_17093,N_17629);
nand U18628 (N_18628,N_17072,N_17242);
nand U18629 (N_18629,N_17109,N_17626);
xnor U18630 (N_18630,N_17075,N_17470);
or U18631 (N_18631,N_17469,N_17172);
and U18632 (N_18632,N_17935,N_17309);
nor U18633 (N_18633,N_17915,N_17079);
and U18634 (N_18634,N_17806,N_17420);
nand U18635 (N_18635,N_17210,N_17817);
nand U18636 (N_18636,N_17938,N_17154);
or U18637 (N_18637,N_17637,N_17979);
nor U18638 (N_18638,N_17160,N_17632);
or U18639 (N_18639,N_17294,N_17663);
or U18640 (N_18640,N_17520,N_17145);
and U18641 (N_18641,N_17355,N_17571);
xnor U18642 (N_18642,N_17161,N_17697);
xnor U18643 (N_18643,N_17474,N_17914);
or U18644 (N_18644,N_17577,N_17872);
or U18645 (N_18645,N_17104,N_17838);
nand U18646 (N_18646,N_17759,N_17173);
nor U18647 (N_18647,N_17546,N_17704);
xnor U18648 (N_18648,N_17946,N_17538);
xor U18649 (N_18649,N_17006,N_17648);
xor U18650 (N_18650,N_17787,N_17465);
or U18651 (N_18651,N_17416,N_17793);
nor U18652 (N_18652,N_17392,N_17686);
or U18653 (N_18653,N_17389,N_17745);
nand U18654 (N_18654,N_17252,N_17896);
nor U18655 (N_18655,N_17623,N_17619);
xor U18656 (N_18656,N_17445,N_17466);
nor U18657 (N_18657,N_17845,N_17718);
nor U18658 (N_18658,N_17379,N_17953);
nor U18659 (N_18659,N_17396,N_17702);
nand U18660 (N_18660,N_17460,N_17283);
xnor U18661 (N_18661,N_17206,N_17152);
xor U18662 (N_18662,N_17207,N_17703);
xor U18663 (N_18663,N_17464,N_17741);
nor U18664 (N_18664,N_17586,N_17115);
xnor U18665 (N_18665,N_17917,N_17970);
nand U18666 (N_18666,N_17652,N_17279);
and U18667 (N_18667,N_17266,N_17638);
nor U18668 (N_18668,N_17594,N_17222);
nor U18669 (N_18669,N_17137,N_17147);
and U18670 (N_18670,N_17332,N_17176);
nor U18671 (N_18671,N_17794,N_17417);
and U18672 (N_18672,N_17416,N_17898);
nor U18673 (N_18673,N_17891,N_17095);
and U18674 (N_18674,N_17922,N_17913);
xor U18675 (N_18675,N_17518,N_17610);
xor U18676 (N_18676,N_17142,N_17980);
nor U18677 (N_18677,N_17292,N_17262);
nand U18678 (N_18678,N_17505,N_17120);
and U18679 (N_18679,N_17267,N_17088);
or U18680 (N_18680,N_17466,N_17409);
or U18681 (N_18681,N_17148,N_17094);
or U18682 (N_18682,N_17718,N_17387);
nor U18683 (N_18683,N_17127,N_17252);
or U18684 (N_18684,N_17692,N_17133);
nor U18685 (N_18685,N_17061,N_17824);
nand U18686 (N_18686,N_17352,N_17438);
xnor U18687 (N_18687,N_17483,N_17193);
and U18688 (N_18688,N_17554,N_17062);
nand U18689 (N_18689,N_17007,N_17130);
nor U18690 (N_18690,N_17740,N_17224);
xnor U18691 (N_18691,N_17213,N_17287);
xor U18692 (N_18692,N_17971,N_17659);
nor U18693 (N_18693,N_17417,N_17379);
or U18694 (N_18694,N_17841,N_17847);
nand U18695 (N_18695,N_17960,N_17893);
nand U18696 (N_18696,N_17756,N_17036);
nand U18697 (N_18697,N_17568,N_17148);
nand U18698 (N_18698,N_17526,N_17888);
xor U18699 (N_18699,N_17635,N_17057);
nor U18700 (N_18700,N_17173,N_17484);
or U18701 (N_18701,N_17339,N_17600);
nand U18702 (N_18702,N_17546,N_17348);
or U18703 (N_18703,N_17176,N_17206);
and U18704 (N_18704,N_17875,N_17413);
or U18705 (N_18705,N_17912,N_17717);
or U18706 (N_18706,N_17379,N_17110);
xnor U18707 (N_18707,N_17876,N_17969);
or U18708 (N_18708,N_17508,N_17513);
nand U18709 (N_18709,N_17915,N_17786);
or U18710 (N_18710,N_17517,N_17352);
or U18711 (N_18711,N_17091,N_17891);
xor U18712 (N_18712,N_17281,N_17387);
and U18713 (N_18713,N_17907,N_17817);
nor U18714 (N_18714,N_17032,N_17009);
or U18715 (N_18715,N_17071,N_17193);
or U18716 (N_18716,N_17759,N_17749);
nor U18717 (N_18717,N_17427,N_17986);
and U18718 (N_18718,N_17677,N_17530);
nor U18719 (N_18719,N_17144,N_17674);
nor U18720 (N_18720,N_17525,N_17760);
or U18721 (N_18721,N_17267,N_17182);
nor U18722 (N_18722,N_17642,N_17632);
or U18723 (N_18723,N_17786,N_17791);
and U18724 (N_18724,N_17082,N_17923);
nand U18725 (N_18725,N_17053,N_17881);
xor U18726 (N_18726,N_17979,N_17257);
nand U18727 (N_18727,N_17330,N_17213);
and U18728 (N_18728,N_17211,N_17183);
nor U18729 (N_18729,N_17378,N_17087);
and U18730 (N_18730,N_17987,N_17939);
xor U18731 (N_18731,N_17296,N_17628);
xnor U18732 (N_18732,N_17407,N_17352);
nand U18733 (N_18733,N_17795,N_17754);
or U18734 (N_18734,N_17643,N_17655);
xor U18735 (N_18735,N_17993,N_17768);
or U18736 (N_18736,N_17968,N_17424);
nor U18737 (N_18737,N_17373,N_17211);
xnor U18738 (N_18738,N_17843,N_17148);
or U18739 (N_18739,N_17659,N_17876);
nand U18740 (N_18740,N_17001,N_17626);
nand U18741 (N_18741,N_17730,N_17414);
nor U18742 (N_18742,N_17164,N_17137);
xnor U18743 (N_18743,N_17408,N_17695);
or U18744 (N_18744,N_17581,N_17580);
nand U18745 (N_18745,N_17757,N_17714);
nor U18746 (N_18746,N_17135,N_17370);
or U18747 (N_18747,N_17530,N_17092);
xor U18748 (N_18748,N_17609,N_17543);
nor U18749 (N_18749,N_17176,N_17354);
and U18750 (N_18750,N_17980,N_17700);
or U18751 (N_18751,N_17691,N_17474);
or U18752 (N_18752,N_17822,N_17956);
and U18753 (N_18753,N_17342,N_17793);
nand U18754 (N_18754,N_17898,N_17953);
nor U18755 (N_18755,N_17733,N_17281);
nor U18756 (N_18756,N_17117,N_17607);
xor U18757 (N_18757,N_17372,N_17547);
nor U18758 (N_18758,N_17399,N_17587);
xor U18759 (N_18759,N_17386,N_17688);
xnor U18760 (N_18760,N_17951,N_17813);
xnor U18761 (N_18761,N_17963,N_17627);
xor U18762 (N_18762,N_17967,N_17532);
and U18763 (N_18763,N_17378,N_17485);
and U18764 (N_18764,N_17332,N_17288);
nand U18765 (N_18765,N_17221,N_17513);
nor U18766 (N_18766,N_17803,N_17660);
or U18767 (N_18767,N_17778,N_17963);
and U18768 (N_18768,N_17034,N_17683);
or U18769 (N_18769,N_17967,N_17143);
nand U18770 (N_18770,N_17825,N_17226);
nand U18771 (N_18771,N_17831,N_17004);
and U18772 (N_18772,N_17486,N_17318);
xor U18773 (N_18773,N_17778,N_17425);
or U18774 (N_18774,N_17090,N_17922);
and U18775 (N_18775,N_17460,N_17194);
or U18776 (N_18776,N_17251,N_17574);
or U18777 (N_18777,N_17296,N_17073);
or U18778 (N_18778,N_17711,N_17272);
nand U18779 (N_18779,N_17655,N_17547);
and U18780 (N_18780,N_17592,N_17446);
xor U18781 (N_18781,N_17412,N_17403);
nor U18782 (N_18782,N_17658,N_17169);
and U18783 (N_18783,N_17068,N_17173);
nand U18784 (N_18784,N_17642,N_17423);
and U18785 (N_18785,N_17036,N_17641);
and U18786 (N_18786,N_17086,N_17006);
nand U18787 (N_18787,N_17124,N_17116);
or U18788 (N_18788,N_17192,N_17096);
nor U18789 (N_18789,N_17574,N_17783);
xnor U18790 (N_18790,N_17749,N_17962);
nand U18791 (N_18791,N_17348,N_17664);
or U18792 (N_18792,N_17755,N_17015);
xor U18793 (N_18793,N_17103,N_17732);
or U18794 (N_18794,N_17810,N_17460);
nand U18795 (N_18795,N_17717,N_17287);
nand U18796 (N_18796,N_17250,N_17073);
nand U18797 (N_18797,N_17790,N_17593);
and U18798 (N_18798,N_17193,N_17506);
nand U18799 (N_18799,N_17922,N_17549);
and U18800 (N_18800,N_17427,N_17569);
xor U18801 (N_18801,N_17163,N_17053);
nor U18802 (N_18802,N_17861,N_17032);
nor U18803 (N_18803,N_17796,N_17139);
or U18804 (N_18804,N_17477,N_17479);
and U18805 (N_18805,N_17389,N_17184);
xor U18806 (N_18806,N_17850,N_17942);
nor U18807 (N_18807,N_17401,N_17649);
or U18808 (N_18808,N_17193,N_17464);
nand U18809 (N_18809,N_17308,N_17005);
nor U18810 (N_18810,N_17753,N_17162);
nand U18811 (N_18811,N_17458,N_17137);
or U18812 (N_18812,N_17707,N_17803);
nor U18813 (N_18813,N_17629,N_17503);
nand U18814 (N_18814,N_17932,N_17316);
nand U18815 (N_18815,N_17237,N_17654);
xnor U18816 (N_18816,N_17888,N_17153);
nand U18817 (N_18817,N_17889,N_17961);
or U18818 (N_18818,N_17241,N_17656);
nor U18819 (N_18819,N_17563,N_17995);
or U18820 (N_18820,N_17388,N_17381);
nor U18821 (N_18821,N_17223,N_17621);
and U18822 (N_18822,N_17745,N_17500);
and U18823 (N_18823,N_17992,N_17843);
or U18824 (N_18824,N_17488,N_17239);
and U18825 (N_18825,N_17824,N_17722);
or U18826 (N_18826,N_17208,N_17675);
or U18827 (N_18827,N_17070,N_17110);
xor U18828 (N_18828,N_17587,N_17372);
nand U18829 (N_18829,N_17411,N_17473);
nor U18830 (N_18830,N_17775,N_17830);
xor U18831 (N_18831,N_17131,N_17228);
and U18832 (N_18832,N_17933,N_17695);
nor U18833 (N_18833,N_17507,N_17669);
nor U18834 (N_18834,N_17608,N_17088);
xor U18835 (N_18835,N_17526,N_17521);
nor U18836 (N_18836,N_17374,N_17806);
nor U18837 (N_18837,N_17547,N_17626);
nand U18838 (N_18838,N_17806,N_17469);
xnor U18839 (N_18839,N_17568,N_17613);
xor U18840 (N_18840,N_17521,N_17439);
or U18841 (N_18841,N_17651,N_17655);
nor U18842 (N_18842,N_17123,N_17502);
xor U18843 (N_18843,N_17676,N_17199);
nor U18844 (N_18844,N_17725,N_17530);
xor U18845 (N_18845,N_17190,N_17976);
xor U18846 (N_18846,N_17484,N_17797);
xor U18847 (N_18847,N_17043,N_17774);
xnor U18848 (N_18848,N_17478,N_17001);
nor U18849 (N_18849,N_17045,N_17371);
and U18850 (N_18850,N_17937,N_17456);
or U18851 (N_18851,N_17715,N_17212);
xor U18852 (N_18852,N_17320,N_17090);
nand U18853 (N_18853,N_17151,N_17949);
nor U18854 (N_18854,N_17927,N_17097);
and U18855 (N_18855,N_17892,N_17415);
or U18856 (N_18856,N_17690,N_17439);
nand U18857 (N_18857,N_17584,N_17341);
nand U18858 (N_18858,N_17638,N_17375);
nor U18859 (N_18859,N_17506,N_17675);
and U18860 (N_18860,N_17762,N_17690);
or U18861 (N_18861,N_17846,N_17133);
xnor U18862 (N_18862,N_17449,N_17795);
nand U18863 (N_18863,N_17861,N_17689);
nor U18864 (N_18864,N_17174,N_17648);
xor U18865 (N_18865,N_17024,N_17534);
nand U18866 (N_18866,N_17672,N_17784);
nor U18867 (N_18867,N_17618,N_17171);
nor U18868 (N_18868,N_17491,N_17856);
or U18869 (N_18869,N_17020,N_17985);
nand U18870 (N_18870,N_17931,N_17702);
and U18871 (N_18871,N_17943,N_17383);
xor U18872 (N_18872,N_17836,N_17397);
and U18873 (N_18873,N_17644,N_17721);
and U18874 (N_18874,N_17917,N_17309);
xor U18875 (N_18875,N_17938,N_17338);
nor U18876 (N_18876,N_17304,N_17547);
or U18877 (N_18877,N_17207,N_17852);
and U18878 (N_18878,N_17576,N_17436);
nor U18879 (N_18879,N_17602,N_17159);
nand U18880 (N_18880,N_17744,N_17778);
nand U18881 (N_18881,N_17428,N_17606);
nand U18882 (N_18882,N_17681,N_17561);
and U18883 (N_18883,N_17037,N_17730);
xor U18884 (N_18884,N_17415,N_17272);
and U18885 (N_18885,N_17302,N_17730);
and U18886 (N_18886,N_17149,N_17937);
or U18887 (N_18887,N_17323,N_17948);
and U18888 (N_18888,N_17880,N_17577);
xnor U18889 (N_18889,N_17622,N_17376);
nor U18890 (N_18890,N_17487,N_17550);
and U18891 (N_18891,N_17158,N_17992);
nand U18892 (N_18892,N_17192,N_17261);
xnor U18893 (N_18893,N_17395,N_17717);
nand U18894 (N_18894,N_17958,N_17030);
and U18895 (N_18895,N_17819,N_17563);
nand U18896 (N_18896,N_17004,N_17472);
or U18897 (N_18897,N_17589,N_17765);
and U18898 (N_18898,N_17132,N_17709);
or U18899 (N_18899,N_17772,N_17220);
or U18900 (N_18900,N_17500,N_17561);
xor U18901 (N_18901,N_17958,N_17139);
nor U18902 (N_18902,N_17530,N_17529);
nor U18903 (N_18903,N_17991,N_17668);
nand U18904 (N_18904,N_17747,N_17466);
nor U18905 (N_18905,N_17637,N_17228);
nor U18906 (N_18906,N_17022,N_17832);
and U18907 (N_18907,N_17289,N_17754);
and U18908 (N_18908,N_17317,N_17240);
nand U18909 (N_18909,N_17615,N_17678);
xnor U18910 (N_18910,N_17712,N_17741);
nand U18911 (N_18911,N_17491,N_17502);
nand U18912 (N_18912,N_17808,N_17418);
xnor U18913 (N_18913,N_17702,N_17202);
and U18914 (N_18914,N_17321,N_17461);
nor U18915 (N_18915,N_17318,N_17844);
or U18916 (N_18916,N_17664,N_17784);
or U18917 (N_18917,N_17417,N_17813);
nor U18918 (N_18918,N_17370,N_17928);
and U18919 (N_18919,N_17056,N_17154);
and U18920 (N_18920,N_17428,N_17942);
nand U18921 (N_18921,N_17579,N_17982);
and U18922 (N_18922,N_17423,N_17713);
and U18923 (N_18923,N_17272,N_17917);
nand U18924 (N_18924,N_17495,N_17561);
nand U18925 (N_18925,N_17343,N_17274);
and U18926 (N_18926,N_17961,N_17694);
nor U18927 (N_18927,N_17598,N_17146);
and U18928 (N_18928,N_17895,N_17920);
and U18929 (N_18929,N_17659,N_17689);
or U18930 (N_18930,N_17811,N_17662);
nor U18931 (N_18931,N_17741,N_17788);
or U18932 (N_18932,N_17516,N_17832);
or U18933 (N_18933,N_17927,N_17483);
nor U18934 (N_18934,N_17815,N_17428);
nor U18935 (N_18935,N_17026,N_17794);
or U18936 (N_18936,N_17362,N_17204);
or U18937 (N_18937,N_17131,N_17307);
xor U18938 (N_18938,N_17859,N_17315);
or U18939 (N_18939,N_17480,N_17943);
nor U18940 (N_18940,N_17267,N_17174);
xor U18941 (N_18941,N_17898,N_17076);
nand U18942 (N_18942,N_17713,N_17021);
nand U18943 (N_18943,N_17849,N_17939);
nor U18944 (N_18944,N_17121,N_17425);
nor U18945 (N_18945,N_17377,N_17196);
and U18946 (N_18946,N_17785,N_17524);
nand U18947 (N_18947,N_17075,N_17522);
nor U18948 (N_18948,N_17615,N_17181);
nand U18949 (N_18949,N_17593,N_17033);
xnor U18950 (N_18950,N_17224,N_17950);
xnor U18951 (N_18951,N_17158,N_17990);
nand U18952 (N_18952,N_17120,N_17993);
xnor U18953 (N_18953,N_17002,N_17135);
nand U18954 (N_18954,N_17797,N_17582);
xnor U18955 (N_18955,N_17823,N_17313);
and U18956 (N_18956,N_17964,N_17263);
or U18957 (N_18957,N_17022,N_17413);
nand U18958 (N_18958,N_17427,N_17310);
or U18959 (N_18959,N_17829,N_17896);
or U18960 (N_18960,N_17200,N_17803);
nand U18961 (N_18961,N_17664,N_17811);
xnor U18962 (N_18962,N_17026,N_17856);
nor U18963 (N_18963,N_17380,N_17666);
or U18964 (N_18964,N_17354,N_17321);
and U18965 (N_18965,N_17247,N_17042);
xnor U18966 (N_18966,N_17698,N_17298);
nand U18967 (N_18967,N_17500,N_17662);
nand U18968 (N_18968,N_17092,N_17897);
or U18969 (N_18969,N_17523,N_17960);
nor U18970 (N_18970,N_17944,N_17565);
nand U18971 (N_18971,N_17101,N_17411);
nand U18972 (N_18972,N_17211,N_17336);
nand U18973 (N_18973,N_17603,N_17806);
and U18974 (N_18974,N_17261,N_17672);
xor U18975 (N_18975,N_17797,N_17883);
nand U18976 (N_18976,N_17253,N_17051);
or U18977 (N_18977,N_17413,N_17742);
xnor U18978 (N_18978,N_17015,N_17836);
nand U18979 (N_18979,N_17070,N_17213);
or U18980 (N_18980,N_17113,N_17609);
nand U18981 (N_18981,N_17028,N_17115);
xor U18982 (N_18982,N_17249,N_17367);
xor U18983 (N_18983,N_17130,N_17818);
nor U18984 (N_18984,N_17052,N_17198);
nor U18985 (N_18985,N_17115,N_17560);
or U18986 (N_18986,N_17747,N_17154);
nand U18987 (N_18987,N_17893,N_17767);
nor U18988 (N_18988,N_17359,N_17067);
nand U18989 (N_18989,N_17450,N_17113);
nand U18990 (N_18990,N_17096,N_17592);
nand U18991 (N_18991,N_17742,N_17747);
nor U18992 (N_18992,N_17870,N_17872);
and U18993 (N_18993,N_17202,N_17010);
nand U18994 (N_18994,N_17399,N_17471);
xnor U18995 (N_18995,N_17319,N_17353);
nor U18996 (N_18996,N_17738,N_17907);
xor U18997 (N_18997,N_17943,N_17767);
nand U18998 (N_18998,N_17614,N_17946);
nor U18999 (N_18999,N_17761,N_17651);
xnor U19000 (N_19000,N_18249,N_18301);
nor U19001 (N_19001,N_18983,N_18555);
nand U19002 (N_19002,N_18328,N_18210);
nor U19003 (N_19003,N_18081,N_18359);
nand U19004 (N_19004,N_18697,N_18561);
or U19005 (N_19005,N_18257,N_18919);
xor U19006 (N_19006,N_18025,N_18826);
nor U19007 (N_19007,N_18549,N_18295);
nand U19008 (N_19008,N_18197,N_18304);
or U19009 (N_19009,N_18052,N_18538);
nand U19010 (N_19010,N_18439,N_18226);
nor U19011 (N_19011,N_18221,N_18784);
nand U19012 (N_19012,N_18687,N_18120);
nor U19013 (N_19013,N_18125,N_18633);
or U19014 (N_19014,N_18253,N_18695);
and U19015 (N_19015,N_18181,N_18563);
or U19016 (N_19016,N_18230,N_18469);
nand U19017 (N_19017,N_18392,N_18461);
and U19018 (N_19018,N_18040,N_18757);
nand U19019 (N_19019,N_18817,N_18048);
xnor U19020 (N_19020,N_18338,N_18786);
nand U19021 (N_19021,N_18426,N_18487);
nor U19022 (N_19022,N_18551,N_18146);
nand U19023 (N_19023,N_18101,N_18660);
nand U19024 (N_19024,N_18476,N_18128);
xor U19025 (N_19025,N_18227,N_18195);
nand U19026 (N_19026,N_18175,N_18150);
nor U19027 (N_19027,N_18039,N_18132);
xor U19028 (N_19028,N_18577,N_18258);
xnor U19029 (N_19029,N_18051,N_18397);
nor U19030 (N_19030,N_18918,N_18155);
or U19031 (N_19031,N_18104,N_18030);
xnor U19032 (N_19032,N_18722,N_18746);
xor U19033 (N_19033,N_18365,N_18381);
nand U19034 (N_19034,N_18765,N_18739);
or U19035 (N_19035,N_18999,N_18590);
xnor U19036 (N_19036,N_18006,N_18431);
and U19037 (N_19037,N_18193,N_18570);
and U19038 (N_19038,N_18942,N_18066);
nor U19039 (N_19039,N_18761,N_18846);
xor U19040 (N_19040,N_18886,N_18848);
nand U19041 (N_19041,N_18485,N_18357);
and U19042 (N_19042,N_18941,N_18995);
xnor U19043 (N_19043,N_18454,N_18776);
and U19044 (N_19044,N_18812,N_18875);
xor U19045 (N_19045,N_18756,N_18018);
and U19046 (N_19046,N_18478,N_18882);
nor U19047 (N_19047,N_18803,N_18928);
nand U19048 (N_19048,N_18429,N_18562);
or U19049 (N_19049,N_18038,N_18837);
nor U19050 (N_19050,N_18732,N_18363);
xnor U19051 (N_19051,N_18893,N_18534);
or U19052 (N_19052,N_18185,N_18599);
nand U19053 (N_19053,N_18419,N_18537);
and U19054 (N_19054,N_18654,N_18109);
or U19055 (N_19055,N_18348,N_18289);
or U19056 (N_19056,N_18926,N_18573);
or U19057 (N_19057,N_18200,N_18134);
nor U19058 (N_19058,N_18143,N_18859);
nor U19059 (N_19059,N_18675,N_18007);
xor U19060 (N_19060,N_18266,N_18058);
nand U19061 (N_19061,N_18730,N_18307);
nor U19062 (N_19062,N_18644,N_18064);
nand U19063 (N_19063,N_18932,N_18208);
or U19064 (N_19064,N_18093,N_18901);
and U19065 (N_19065,N_18275,N_18750);
xor U19066 (N_19066,N_18914,N_18718);
xnor U19067 (N_19067,N_18661,N_18671);
or U19068 (N_19068,N_18530,N_18184);
nor U19069 (N_19069,N_18115,N_18147);
or U19070 (N_19070,N_18522,N_18892);
and U19071 (N_19071,N_18626,N_18499);
nand U19072 (N_19072,N_18246,N_18923);
or U19073 (N_19073,N_18665,N_18664);
or U19074 (N_19074,N_18311,N_18390);
nor U19075 (N_19075,N_18055,N_18690);
nor U19076 (N_19076,N_18020,N_18232);
and U19077 (N_19077,N_18323,N_18922);
or U19078 (N_19078,N_18380,N_18580);
nand U19079 (N_19079,N_18740,N_18993);
or U19080 (N_19080,N_18078,N_18717);
and U19081 (N_19081,N_18282,N_18008);
and U19082 (N_19082,N_18514,N_18989);
nor U19083 (N_19083,N_18847,N_18624);
xor U19084 (N_19084,N_18236,N_18736);
and U19085 (N_19085,N_18069,N_18996);
nand U19086 (N_19086,N_18327,N_18368);
nor U19087 (N_19087,N_18141,N_18828);
or U19088 (N_19088,N_18890,N_18685);
xor U19089 (N_19089,N_18871,N_18260);
nand U19090 (N_19090,N_18743,N_18910);
and U19091 (N_19091,N_18726,N_18869);
and U19092 (N_19092,N_18263,N_18900);
xor U19093 (N_19093,N_18261,N_18924);
or U19094 (N_19094,N_18938,N_18149);
or U19095 (N_19095,N_18474,N_18170);
xnor U19096 (N_19096,N_18374,N_18734);
xnor U19097 (N_19097,N_18558,N_18838);
xnor U19098 (N_19098,N_18477,N_18252);
xor U19099 (N_19099,N_18395,N_18744);
nand U19100 (N_19100,N_18254,N_18201);
or U19101 (N_19101,N_18383,N_18199);
nor U19102 (N_19102,N_18727,N_18242);
xnor U19103 (N_19103,N_18267,N_18724);
and U19104 (N_19104,N_18693,N_18192);
xnor U19105 (N_19105,N_18470,N_18532);
and U19106 (N_19106,N_18127,N_18519);
and U19107 (N_19107,N_18707,N_18105);
nand U19108 (N_19108,N_18572,N_18351);
nor U19109 (N_19109,N_18517,N_18417);
or U19110 (N_19110,N_18306,N_18659);
nor U19111 (N_19111,N_18858,N_18653);
nand U19112 (N_19112,N_18788,N_18895);
nand U19113 (N_19113,N_18962,N_18747);
or U19114 (N_19114,N_18407,N_18488);
nor U19115 (N_19115,N_18814,N_18314);
or U19116 (N_19116,N_18872,N_18000);
and U19117 (N_19117,N_18174,N_18436);
and U19118 (N_19118,N_18234,N_18421);
or U19119 (N_19119,N_18604,N_18600);
nand U19120 (N_19120,N_18523,N_18168);
or U19121 (N_19121,N_18832,N_18943);
nor U19122 (N_19122,N_18865,N_18703);
nor U19123 (N_19123,N_18864,N_18107);
and U19124 (N_19124,N_18513,N_18584);
and U19125 (N_19125,N_18643,N_18594);
nor U19126 (N_19126,N_18767,N_18940);
nor U19127 (N_19127,N_18984,N_18084);
xnor U19128 (N_19128,N_18879,N_18694);
nand U19129 (N_19129,N_18967,N_18949);
and U19130 (N_19130,N_18621,N_18585);
nand U19131 (N_19131,N_18638,N_18112);
or U19132 (N_19132,N_18632,N_18430);
nor U19133 (N_19133,N_18080,N_18033);
xor U19134 (N_19134,N_18162,N_18711);
or U19135 (N_19135,N_18974,N_18891);
nand U19136 (N_19136,N_18712,N_18557);
and U19137 (N_19137,N_18542,N_18404);
and U19138 (N_19138,N_18849,N_18804);
or U19139 (N_19139,N_18031,N_18535);
nand U19140 (N_19140,N_18823,N_18264);
nor U19141 (N_19141,N_18163,N_18219);
nor U19142 (N_19142,N_18507,N_18681);
nand U19143 (N_19143,N_18618,N_18937);
xor U19144 (N_19144,N_18623,N_18965);
or U19145 (N_19145,N_18027,N_18142);
xor U19146 (N_19146,N_18096,N_18516);
and U19147 (N_19147,N_18228,N_18936);
and U19148 (N_19148,N_18539,N_18198);
xor U19149 (N_19149,N_18686,N_18482);
nor U19150 (N_19150,N_18309,N_18220);
xnor U19151 (N_19151,N_18668,N_18673);
nor U19152 (N_19152,N_18370,N_18443);
or U19153 (N_19153,N_18355,N_18164);
nor U19154 (N_19154,N_18867,N_18586);
and U19155 (N_19155,N_18975,N_18795);
xnor U19156 (N_19156,N_18243,N_18369);
and U19157 (N_19157,N_18728,N_18953);
and U19158 (N_19158,N_18554,N_18990);
or U19159 (N_19159,N_18930,N_18769);
and U19160 (N_19160,N_18959,N_18830);
or U19161 (N_19161,N_18316,N_18777);
and U19162 (N_19162,N_18546,N_18839);
xor U19163 (N_19163,N_18315,N_18605);
xnor U19164 (N_19164,N_18427,N_18720);
or U19165 (N_19165,N_18280,N_18224);
and U19166 (N_19166,N_18362,N_18620);
nand U19167 (N_19167,N_18716,N_18509);
nand U19168 (N_19168,N_18933,N_18366);
nand U19169 (N_19169,N_18256,N_18160);
or U19170 (N_19170,N_18087,N_18899);
and U19171 (N_19171,N_18495,N_18816);
and U19172 (N_19172,N_18709,N_18334);
nor U19173 (N_19173,N_18097,N_18721);
nor U19174 (N_19174,N_18455,N_18272);
or U19175 (N_19175,N_18887,N_18708);
or U19176 (N_19176,N_18755,N_18475);
nor U19177 (N_19177,N_18944,N_18305);
nand U19178 (N_19178,N_18931,N_18980);
xor U19179 (N_19179,N_18001,N_18543);
nor U19180 (N_19180,N_18152,N_18131);
xnor U19181 (N_19181,N_18780,N_18925);
nor U19182 (N_19182,N_18836,N_18670);
nand U19183 (N_19183,N_18412,N_18528);
xnor U19184 (N_19184,N_18403,N_18428);
and U19185 (N_19185,N_18218,N_18679);
xnor U19186 (N_19186,N_18748,N_18606);
xor U19187 (N_19187,N_18733,N_18352);
nand U19188 (N_19188,N_18207,N_18715);
nor U19189 (N_19189,N_18462,N_18966);
nor U19190 (N_19190,N_18818,N_18731);
or U19191 (N_19191,N_18014,N_18157);
or U19192 (N_19192,N_18833,N_18229);
or U19193 (N_19193,N_18092,N_18138);
or U19194 (N_19194,N_18574,N_18285);
and U19195 (N_19195,N_18969,N_18636);
and U19196 (N_19196,N_18413,N_18973);
or U19197 (N_19197,N_18269,N_18647);
xor U19198 (N_19198,N_18122,N_18464);
and U19199 (N_19199,N_18987,N_18372);
nand U19200 (N_19200,N_18015,N_18388);
and U19201 (N_19201,N_18399,N_18217);
nand U19202 (N_19202,N_18408,N_18710);
nor U19203 (N_19203,N_18466,N_18345);
or U19204 (N_19204,N_18595,N_18432);
and U19205 (N_19205,N_18533,N_18287);
or U19206 (N_19206,N_18662,N_18531);
xnor U19207 (N_19207,N_18045,N_18753);
xnor U19208 (N_19208,N_18683,N_18335);
and U19209 (N_19209,N_18433,N_18524);
or U19210 (N_19210,N_18111,N_18460);
nor U19211 (N_19211,N_18054,N_18754);
xnor U19212 (N_19212,N_18552,N_18794);
nor U19213 (N_19213,N_18347,N_18920);
nand U19214 (N_19214,N_18159,N_18086);
xor U19215 (N_19215,N_18213,N_18515);
xor U19216 (N_19216,N_18855,N_18699);
nand U19217 (N_19217,N_18473,N_18298);
nor U19218 (N_19218,N_18332,N_18212);
or U19219 (N_19219,N_18801,N_18194);
and U19220 (N_19220,N_18401,N_18319);
nor U19221 (N_19221,N_18593,N_18829);
nand U19222 (N_19222,N_18284,N_18545);
or U19223 (N_19223,N_18077,N_18525);
or U19224 (N_19224,N_18023,N_18760);
and U19225 (N_19225,N_18103,N_18607);
or U19226 (N_19226,N_18279,N_18581);
nor U19227 (N_19227,N_18424,N_18738);
xor U19228 (N_19228,N_18073,N_18442);
nand U19229 (N_19229,N_18663,N_18119);
nand U19230 (N_19230,N_18021,N_18505);
or U19231 (N_19231,N_18290,N_18802);
and U19232 (N_19232,N_18402,N_18457);
and U19233 (N_19233,N_18070,N_18773);
and U19234 (N_19234,N_18050,N_18165);
nand U19235 (N_19235,N_18094,N_18028);
nor U19236 (N_19236,N_18610,N_18749);
and U19237 (N_19237,N_18915,N_18102);
xnor U19238 (N_19238,N_18321,N_18151);
nor U19239 (N_19239,N_18444,N_18735);
nand U19240 (N_19240,N_18797,N_18857);
nor U19241 (N_19241,N_18898,N_18467);
xnor U19242 (N_19242,N_18642,N_18917);
nand U19243 (N_19243,N_18459,N_18903);
nand U19244 (N_19244,N_18927,N_18674);
nor U19245 (N_19245,N_18682,N_18645);
nand U19246 (N_19246,N_18416,N_18972);
and U19247 (N_19247,N_18144,N_18587);
xnor U19248 (N_19248,N_18723,N_18011);
or U19249 (N_19249,N_18425,N_18214);
or U19250 (N_19250,N_18908,N_18768);
nor U19251 (N_19251,N_18579,N_18676);
or U19252 (N_19252,N_18393,N_18520);
nor U19253 (N_19253,N_18449,N_18637);
nor U19254 (N_19254,N_18954,N_18960);
xnor U19255 (N_19255,N_18382,N_18527);
or U19256 (N_19256,N_18188,N_18447);
xnor U19257 (N_19257,N_18405,N_18500);
or U19258 (N_19258,N_18597,N_18700);
or U19259 (N_19259,N_18622,N_18223);
nor U19260 (N_19260,N_18742,N_18751);
nor U19261 (N_19261,N_18190,N_18877);
nor U19262 (N_19262,N_18819,N_18056);
nand U19263 (N_19263,N_18759,N_18035);
nand U19264 (N_19264,N_18434,N_18880);
xnor U19265 (N_19265,N_18775,N_18089);
or U19266 (N_19266,N_18518,N_18592);
or U19267 (N_19267,N_18656,N_18613);
or U19268 (N_19268,N_18391,N_18822);
nand U19269 (N_19269,N_18815,N_18237);
nor U19270 (N_19270,N_18627,N_18982);
nor U19271 (N_19271,N_18608,N_18255);
and U19272 (N_19272,N_18293,N_18176);
or U19273 (N_19273,N_18696,N_18326);
and U19274 (N_19274,N_18386,N_18169);
nor U19275 (N_19275,N_18912,N_18963);
or U19276 (N_19276,N_18651,N_18688);
nand U19277 (N_19277,N_18994,N_18167);
nor U19278 (N_19278,N_18398,N_18484);
xor U19279 (N_19279,N_18649,N_18971);
xor U19280 (N_19280,N_18437,N_18781);
nand U19281 (N_19281,N_18772,N_18400);
nand U19282 (N_19282,N_18680,N_18807);
xor U19283 (N_19283,N_18344,N_18490);
xor U19284 (N_19284,N_18017,N_18059);
or U19285 (N_19285,N_18968,N_18079);
and U19286 (N_19286,N_18916,N_18019);
nand U19287 (N_19287,N_18281,N_18611);
or U19288 (N_19288,N_18379,N_18313);
or U19289 (N_19289,N_18512,N_18779);
nand U19290 (N_19290,N_18053,N_18265);
or U19291 (N_19291,N_18782,N_18043);
nor U19292 (N_19292,N_18706,N_18568);
xnor U19293 (N_19293,N_18148,N_18894);
nand U19294 (N_19294,N_18628,N_18583);
xor U19295 (N_19295,N_18046,N_18640);
or U19296 (N_19296,N_18438,N_18418);
xnor U19297 (N_19297,N_18560,N_18648);
nand U19298 (N_19298,N_18657,N_18248);
or U19299 (N_19299,N_18614,N_18133);
and U19300 (N_19300,N_18231,N_18906);
and U19301 (N_19301,N_18124,N_18286);
xnor U19302 (N_19302,N_18825,N_18114);
and U19303 (N_19303,N_18991,N_18881);
or U19304 (N_19304,N_18853,N_18251);
nand U19305 (N_19305,N_18929,N_18725);
xnor U19306 (N_19306,N_18322,N_18268);
nand U19307 (N_19307,N_18294,N_18835);
nor U19308 (N_19308,N_18299,N_18550);
and U19309 (N_19309,N_18737,N_18582);
nand U19310 (N_19310,N_18806,N_18486);
nor U19311 (N_19311,N_18870,N_18762);
nand U19312 (N_19312,N_18082,N_18354);
nor U19313 (N_19313,N_18451,N_18339);
xnor U19314 (N_19314,N_18126,N_18161);
nand U19315 (N_19315,N_18905,N_18153);
nor U19316 (N_19316,N_18129,N_18502);
xor U19317 (N_19317,N_18957,N_18186);
or U19318 (N_19318,N_18988,N_18576);
nor U19319 (N_19319,N_18396,N_18037);
or U19320 (N_19320,N_18448,N_18329);
and U19321 (N_19321,N_18420,N_18824);
nor U19322 (N_19322,N_18009,N_18571);
or U19323 (N_19323,N_18884,N_18625);
nand U19324 (N_19324,N_18778,N_18764);
or U19325 (N_19325,N_18808,N_18410);
nand U19326 (N_19326,N_18222,N_18866);
or U19327 (N_19327,N_18156,N_18456);
nor U19328 (N_19328,N_18977,N_18140);
and U19329 (N_19329,N_18446,N_18100);
nor U19330 (N_19330,N_18411,N_18377);
or U19331 (N_19331,N_18575,N_18095);
nor U19332 (N_19332,N_18805,N_18075);
and U19333 (N_19333,N_18445,N_18771);
and U19334 (N_19334,N_18068,N_18452);
and U19335 (N_19335,N_18591,N_18239);
nand U19336 (N_19336,N_18130,N_18791);
xor U19337 (N_19337,N_18787,N_18312);
or U19338 (N_19338,N_18308,N_18415);
nand U19339 (N_19339,N_18752,N_18116);
nand U19340 (N_19340,N_18353,N_18745);
and U19341 (N_19341,N_18209,N_18179);
nor U19342 (N_19342,N_18939,N_18024);
nand U19343 (N_19343,N_18841,N_18741);
or U19344 (N_19344,N_18216,N_18529);
xnor U19345 (N_19345,N_18360,N_18506);
xnor U19346 (N_19346,N_18854,N_18904);
nand U19347 (N_19347,N_18483,N_18758);
and U19348 (N_19348,N_18074,N_18330);
and U19349 (N_19349,N_18646,N_18278);
nor U19350 (N_19350,N_18985,N_18567);
nor U19351 (N_19351,N_18493,N_18851);
or U19352 (N_19352,N_18961,N_18876);
xor U19353 (N_19353,N_18336,N_18283);
xnor U19354 (N_19354,N_18986,N_18385);
and U19355 (N_19355,N_18811,N_18958);
and U19356 (N_19356,N_18564,N_18565);
xor U19357 (N_19357,N_18566,N_18123);
nand U19358 (N_19358,N_18701,N_18770);
xor U19359 (N_19359,N_18414,N_18145);
or U19360 (N_19360,N_18350,N_18501);
nor U19361 (N_19361,N_18106,N_18491);
and U19362 (N_19362,N_18245,N_18569);
or U19363 (N_19363,N_18800,N_18292);
nand U19364 (N_19364,N_18631,N_18809);
nor U19365 (N_19365,N_18384,N_18247);
xnor U19366 (N_19366,N_18076,N_18061);
and U19367 (N_19367,N_18856,N_18510);
or U19368 (N_19368,N_18541,N_18177);
nor U19369 (N_19369,N_18065,N_18511);
or U19370 (N_19370,N_18137,N_18719);
and U19371 (N_19371,N_18099,N_18827);
nor U19372 (N_19372,N_18793,N_18979);
or U19373 (N_19373,N_18154,N_18843);
nor U19374 (N_19374,N_18598,N_18766);
nand U19375 (N_19375,N_18652,N_18191);
or U19376 (N_19376,N_18296,N_18274);
nor U19377 (N_19377,N_18955,N_18845);
xor U19378 (N_19378,N_18303,N_18796);
nor U19379 (N_19379,N_18342,N_18612);
xor U19380 (N_19380,N_18083,N_18036);
nor U19381 (N_19381,N_18002,N_18005);
xnor U19382 (N_19382,N_18435,N_18003);
nor U19383 (N_19383,N_18998,N_18012);
and U19384 (N_19384,N_18792,N_18831);
xor U19385 (N_19385,N_18616,N_18375);
nand U19386 (N_19386,N_18602,N_18349);
nor U19387 (N_19387,N_18821,N_18799);
and U19388 (N_19388,N_18139,N_18536);
nand U19389 (N_19389,N_18136,N_18559);
xor U19390 (N_19390,N_18714,N_18885);
xnor U19391 (N_19391,N_18774,N_18356);
xor U19392 (N_19392,N_18063,N_18883);
nand U19393 (N_19393,N_18032,N_18049);
or U19394 (N_19394,N_18422,N_18698);
nor U19395 (N_19395,N_18238,N_18547);
nand U19396 (N_19396,N_18423,N_18911);
nand U19397 (N_19397,N_18324,N_18297);
nor U19398 (N_19398,N_18878,N_18964);
or U19399 (N_19399,N_18317,N_18763);
or U19400 (N_19400,N_18861,N_18970);
nor U19401 (N_19401,N_18783,N_18108);
xnor U19402 (N_19402,N_18183,N_18498);
nand U19403 (N_19403,N_18948,N_18166);
xor U19404 (N_19404,N_18158,N_18016);
and U19405 (N_19405,N_18704,N_18480);
nor U19406 (N_19406,N_18450,N_18113);
and U19407 (N_19407,N_18271,N_18333);
and U19408 (N_19408,N_18641,N_18067);
or U19409 (N_19409,N_18658,N_18098);
or U19410 (N_19410,N_18820,N_18540);
nand U19411 (N_19411,N_18041,N_18553);
nor U19412 (N_19412,N_18004,N_18609);
nand U19413 (N_19413,N_18376,N_18873);
nor U19414 (N_19414,N_18273,N_18496);
xnor U19415 (N_19415,N_18494,N_18178);
xnor U19416 (N_19416,N_18992,N_18601);
nand U19417 (N_19417,N_18182,N_18302);
and U19418 (N_19418,N_18172,N_18346);
and U19419 (N_19419,N_18010,N_18489);
nor U19420 (N_19420,N_18013,N_18318);
xor U19421 (N_19421,N_18276,N_18689);
xnor U19422 (N_19422,N_18913,N_18834);
nand U19423 (N_19423,N_18463,N_18952);
or U19424 (N_19424,N_18389,N_18981);
nor U19425 (N_19425,N_18578,N_18310);
nor U19426 (N_19426,N_18934,N_18852);
and U19427 (N_19427,N_18291,N_18902);
and U19428 (N_19428,N_18300,N_18888);
nand U19429 (N_19429,N_18202,N_18042);
nor U19430 (N_19430,N_18471,N_18072);
xnor U19431 (N_19431,N_18378,N_18874);
or U19432 (N_19432,N_18343,N_18785);
nor U19433 (N_19433,N_18364,N_18860);
or U19434 (N_19434,N_18135,N_18409);
and U19435 (N_19435,N_18225,N_18705);
xor U19436 (N_19436,N_18088,N_18241);
nand U19437 (N_19437,N_18341,N_18619);
or U19438 (N_19438,N_18026,N_18337);
xor U19439 (N_19439,N_18667,N_18947);
nor U19440 (N_19440,N_18526,N_18907);
or U19441 (N_19441,N_18203,N_18233);
xnor U19442 (N_19442,N_18548,N_18090);
xnor U19443 (N_19443,N_18672,N_18121);
and U19444 (N_19444,N_18367,N_18504);
or U19445 (N_19445,N_18863,N_18034);
xor U19446 (N_19446,N_18950,N_18118);
nand U19447 (N_19447,N_18503,N_18669);
nor U19448 (N_19448,N_18842,N_18521);
and U19449 (N_19449,N_18071,N_18085);
nor U19450 (N_19450,N_18173,N_18205);
and U19451 (N_19451,N_18394,N_18544);
or U19452 (N_19452,N_18277,N_18022);
xnor U19453 (N_19453,N_18492,N_18997);
xnor U19454 (N_19454,N_18889,N_18091);
or U19455 (N_19455,N_18588,N_18702);
xor U19456 (N_19456,N_18921,N_18897);
nor U19457 (N_19457,N_18684,N_18240);
and U19458 (N_19458,N_18691,N_18458);
nor U19459 (N_19459,N_18678,N_18713);
nand U19460 (N_19460,N_18187,N_18868);
or U19461 (N_19461,N_18655,N_18047);
xor U19462 (N_19462,N_18371,N_18262);
xnor U19463 (N_19463,N_18250,N_18320);
xor U19464 (N_19464,N_18044,N_18978);
and U19465 (N_19465,N_18850,N_18440);
nand U19466 (N_19466,N_18029,N_18196);
and U19467 (N_19467,N_18441,N_18617);
and U19468 (N_19468,N_18956,N_18589);
xnor U19469 (N_19469,N_18508,N_18813);
and U19470 (N_19470,N_18453,N_18946);
or U19471 (N_19471,N_18206,N_18840);
nor U19472 (N_19472,N_18789,N_18945);
and U19473 (N_19473,N_18639,N_18692);
nor U19474 (N_19474,N_18634,N_18331);
nand U19475 (N_19475,N_18615,N_18060);
or U19476 (N_19476,N_18896,N_18057);
xor U19477 (N_19477,N_18810,N_18976);
xor U19478 (N_19478,N_18288,N_18117);
and U19479 (N_19479,N_18481,N_18666);
and U19480 (N_19480,N_18215,N_18497);
xor U19481 (N_19481,N_18235,N_18259);
nor U19482 (N_19482,N_18180,N_18630);
xnor U19483 (N_19483,N_18479,N_18189);
and U19484 (N_19484,N_18244,N_18556);
xnor U19485 (N_19485,N_18862,N_18650);
xor U19486 (N_19486,N_18270,N_18677);
nand U19487 (N_19487,N_18110,N_18472);
xor U19488 (N_19488,N_18909,N_18629);
xor U19489 (N_19489,N_18635,N_18171);
nand U19490 (N_19490,N_18844,N_18361);
nand U19491 (N_19491,N_18465,N_18204);
or U19492 (N_19492,N_18596,N_18406);
and U19493 (N_19493,N_18373,N_18790);
xor U19494 (N_19494,N_18935,N_18340);
or U19495 (N_19495,N_18387,N_18062);
nand U19496 (N_19496,N_18325,N_18468);
or U19497 (N_19497,N_18729,N_18603);
nor U19498 (N_19498,N_18951,N_18358);
nor U19499 (N_19499,N_18798,N_18211);
xnor U19500 (N_19500,N_18222,N_18728);
or U19501 (N_19501,N_18325,N_18418);
xor U19502 (N_19502,N_18724,N_18387);
nand U19503 (N_19503,N_18966,N_18747);
and U19504 (N_19504,N_18677,N_18832);
and U19505 (N_19505,N_18377,N_18662);
nand U19506 (N_19506,N_18349,N_18497);
nor U19507 (N_19507,N_18584,N_18858);
and U19508 (N_19508,N_18601,N_18836);
nor U19509 (N_19509,N_18343,N_18095);
xnor U19510 (N_19510,N_18670,N_18472);
xor U19511 (N_19511,N_18230,N_18140);
or U19512 (N_19512,N_18142,N_18950);
nand U19513 (N_19513,N_18596,N_18444);
xor U19514 (N_19514,N_18279,N_18309);
nor U19515 (N_19515,N_18347,N_18002);
and U19516 (N_19516,N_18936,N_18708);
or U19517 (N_19517,N_18024,N_18917);
and U19518 (N_19518,N_18062,N_18310);
nand U19519 (N_19519,N_18887,N_18005);
and U19520 (N_19520,N_18028,N_18735);
or U19521 (N_19521,N_18213,N_18696);
or U19522 (N_19522,N_18068,N_18920);
nand U19523 (N_19523,N_18325,N_18702);
or U19524 (N_19524,N_18879,N_18969);
and U19525 (N_19525,N_18891,N_18366);
nand U19526 (N_19526,N_18864,N_18527);
or U19527 (N_19527,N_18977,N_18159);
or U19528 (N_19528,N_18215,N_18881);
or U19529 (N_19529,N_18166,N_18042);
or U19530 (N_19530,N_18570,N_18320);
and U19531 (N_19531,N_18547,N_18464);
nand U19532 (N_19532,N_18961,N_18674);
nand U19533 (N_19533,N_18005,N_18282);
nor U19534 (N_19534,N_18815,N_18321);
nand U19535 (N_19535,N_18760,N_18234);
or U19536 (N_19536,N_18531,N_18151);
xor U19537 (N_19537,N_18781,N_18644);
nand U19538 (N_19538,N_18281,N_18711);
nand U19539 (N_19539,N_18974,N_18076);
xor U19540 (N_19540,N_18080,N_18174);
and U19541 (N_19541,N_18199,N_18738);
and U19542 (N_19542,N_18038,N_18573);
and U19543 (N_19543,N_18943,N_18882);
nor U19544 (N_19544,N_18577,N_18051);
and U19545 (N_19545,N_18609,N_18321);
nor U19546 (N_19546,N_18583,N_18313);
or U19547 (N_19547,N_18487,N_18909);
and U19548 (N_19548,N_18505,N_18089);
and U19549 (N_19549,N_18505,N_18871);
nor U19550 (N_19550,N_18555,N_18833);
and U19551 (N_19551,N_18166,N_18285);
xor U19552 (N_19552,N_18010,N_18156);
or U19553 (N_19553,N_18420,N_18255);
xnor U19554 (N_19554,N_18853,N_18655);
xnor U19555 (N_19555,N_18021,N_18739);
nor U19556 (N_19556,N_18521,N_18823);
xnor U19557 (N_19557,N_18126,N_18645);
nand U19558 (N_19558,N_18718,N_18116);
or U19559 (N_19559,N_18997,N_18941);
nor U19560 (N_19560,N_18191,N_18855);
nor U19561 (N_19561,N_18062,N_18281);
nor U19562 (N_19562,N_18071,N_18533);
xor U19563 (N_19563,N_18878,N_18972);
nand U19564 (N_19564,N_18571,N_18665);
nand U19565 (N_19565,N_18124,N_18855);
nand U19566 (N_19566,N_18650,N_18299);
and U19567 (N_19567,N_18098,N_18496);
xnor U19568 (N_19568,N_18064,N_18048);
or U19569 (N_19569,N_18767,N_18904);
xnor U19570 (N_19570,N_18025,N_18085);
nand U19571 (N_19571,N_18491,N_18851);
or U19572 (N_19572,N_18568,N_18735);
nor U19573 (N_19573,N_18095,N_18678);
nand U19574 (N_19574,N_18957,N_18776);
nor U19575 (N_19575,N_18389,N_18041);
or U19576 (N_19576,N_18970,N_18997);
xor U19577 (N_19577,N_18723,N_18116);
xnor U19578 (N_19578,N_18071,N_18545);
and U19579 (N_19579,N_18392,N_18779);
or U19580 (N_19580,N_18067,N_18146);
nand U19581 (N_19581,N_18665,N_18542);
nand U19582 (N_19582,N_18088,N_18433);
and U19583 (N_19583,N_18395,N_18712);
nor U19584 (N_19584,N_18326,N_18858);
and U19585 (N_19585,N_18423,N_18310);
nand U19586 (N_19586,N_18925,N_18544);
and U19587 (N_19587,N_18998,N_18381);
xor U19588 (N_19588,N_18331,N_18480);
or U19589 (N_19589,N_18497,N_18214);
xor U19590 (N_19590,N_18504,N_18862);
or U19591 (N_19591,N_18705,N_18265);
xor U19592 (N_19592,N_18992,N_18085);
xor U19593 (N_19593,N_18688,N_18329);
nand U19594 (N_19594,N_18876,N_18767);
nand U19595 (N_19595,N_18846,N_18111);
xnor U19596 (N_19596,N_18953,N_18895);
xor U19597 (N_19597,N_18772,N_18105);
and U19598 (N_19598,N_18466,N_18467);
nor U19599 (N_19599,N_18439,N_18521);
nor U19600 (N_19600,N_18888,N_18085);
nor U19601 (N_19601,N_18238,N_18432);
or U19602 (N_19602,N_18915,N_18594);
nor U19603 (N_19603,N_18518,N_18122);
and U19604 (N_19604,N_18519,N_18827);
xor U19605 (N_19605,N_18590,N_18218);
xor U19606 (N_19606,N_18428,N_18347);
nand U19607 (N_19607,N_18330,N_18670);
xnor U19608 (N_19608,N_18600,N_18033);
xnor U19609 (N_19609,N_18300,N_18880);
and U19610 (N_19610,N_18743,N_18160);
and U19611 (N_19611,N_18961,N_18840);
nand U19612 (N_19612,N_18408,N_18801);
nand U19613 (N_19613,N_18306,N_18848);
or U19614 (N_19614,N_18753,N_18008);
nor U19615 (N_19615,N_18422,N_18677);
or U19616 (N_19616,N_18373,N_18197);
xnor U19617 (N_19617,N_18723,N_18052);
nor U19618 (N_19618,N_18936,N_18583);
xor U19619 (N_19619,N_18667,N_18676);
xnor U19620 (N_19620,N_18208,N_18725);
or U19621 (N_19621,N_18086,N_18352);
xor U19622 (N_19622,N_18441,N_18645);
and U19623 (N_19623,N_18317,N_18938);
xor U19624 (N_19624,N_18235,N_18811);
and U19625 (N_19625,N_18047,N_18451);
nand U19626 (N_19626,N_18682,N_18397);
xor U19627 (N_19627,N_18661,N_18163);
nor U19628 (N_19628,N_18307,N_18768);
and U19629 (N_19629,N_18577,N_18136);
nand U19630 (N_19630,N_18955,N_18827);
and U19631 (N_19631,N_18090,N_18844);
and U19632 (N_19632,N_18133,N_18544);
nand U19633 (N_19633,N_18512,N_18095);
nand U19634 (N_19634,N_18012,N_18336);
and U19635 (N_19635,N_18101,N_18771);
and U19636 (N_19636,N_18572,N_18888);
and U19637 (N_19637,N_18951,N_18599);
nand U19638 (N_19638,N_18384,N_18091);
xor U19639 (N_19639,N_18945,N_18495);
xnor U19640 (N_19640,N_18505,N_18435);
nand U19641 (N_19641,N_18076,N_18398);
xnor U19642 (N_19642,N_18706,N_18552);
nand U19643 (N_19643,N_18563,N_18939);
nor U19644 (N_19644,N_18598,N_18493);
xor U19645 (N_19645,N_18422,N_18876);
or U19646 (N_19646,N_18847,N_18705);
or U19647 (N_19647,N_18360,N_18882);
or U19648 (N_19648,N_18146,N_18717);
xnor U19649 (N_19649,N_18914,N_18736);
xnor U19650 (N_19650,N_18717,N_18033);
or U19651 (N_19651,N_18953,N_18082);
and U19652 (N_19652,N_18228,N_18646);
and U19653 (N_19653,N_18950,N_18810);
nor U19654 (N_19654,N_18524,N_18633);
nand U19655 (N_19655,N_18243,N_18521);
nand U19656 (N_19656,N_18605,N_18491);
or U19657 (N_19657,N_18904,N_18846);
xor U19658 (N_19658,N_18464,N_18373);
xnor U19659 (N_19659,N_18524,N_18069);
xor U19660 (N_19660,N_18971,N_18740);
xnor U19661 (N_19661,N_18850,N_18809);
and U19662 (N_19662,N_18339,N_18981);
nand U19663 (N_19663,N_18296,N_18605);
nor U19664 (N_19664,N_18672,N_18263);
nor U19665 (N_19665,N_18494,N_18268);
nand U19666 (N_19666,N_18012,N_18209);
xnor U19667 (N_19667,N_18819,N_18205);
and U19668 (N_19668,N_18942,N_18383);
nand U19669 (N_19669,N_18125,N_18899);
and U19670 (N_19670,N_18199,N_18802);
nor U19671 (N_19671,N_18994,N_18636);
and U19672 (N_19672,N_18259,N_18262);
and U19673 (N_19673,N_18444,N_18132);
nand U19674 (N_19674,N_18946,N_18269);
nand U19675 (N_19675,N_18025,N_18236);
nor U19676 (N_19676,N_18761,N_18525);
nor U19677 (N_19677,N_18791,N_18661);
xnor U19678 (N_19678,N_18290,N_18642);
or U19679 (N_19679,N_18585,N_18266);
nand U19680 (N_19680,N_18061,N_18876);
and U19681 (N_19681,N_18080,N_18038);
and U19682 (N_19682,N_18465,N_18740);
nor U19683 (N_19683,N_18895,N_18080);
and U19684 (N_19684,N_18361,N_18163);
or U19685 (N_19685,N_18263,N_18372);
nand U19686 (N_19686,N_18582,N_18921);
nor U19687 (N_19687,N_18927,N_18852);
nand U19688 (N_19688,N_18080,N_18195);
and U19689 (N_19689,N_18872,N_18737);
nor U19690 (N_19690,N_18005,N_18833);
nand U19691 (N_19691,N_18096,N_18375);
nor U19692 (N_19692,N_18964,N_18722);
xor U19693 (N_19693,N_18776,N_18361);
or U19694 (N_19694,N_18530,N_18728);
nand U19695 (N_19695,N_18547,N_18855);
or U19696 (N_19696,N_18610,N_18144);
or U19697 (N_19697,N_18070,N_18990);
or U19698 (N_19698,N_18204,N_18196);
or U19699 (N_19699,N_18616,N_18467);
or U19700 (N_19700,N_18656,N_18724);
nor U19701 (N_19701,N_18233,N_18958);
and U19702 (N_19702,N_18356,N_18686);
and U19703 (N_19703,N_18014,N_18586);
nor U19704 (N_19704,N_18955,N_18609);
xnor U19705 (N_19705,N_18540,N_18237);
and U19706 (N_19706,N_18742,N_18791);
and U19707 (N_19707,N_18311,N_18546);
xor U19708 (N_19708,N_18915,N_18097);
nand U19709 (N_19709,N_18617,N_18516);
nor U19710 (N_19710,N_18707,N_18710);
xor U19711 (N_19711,N_18210,N_18031);
and U19712 (N_19712,N_18568,N_18627);
xor U19713 (N_19713,N_18265,N_18535);
and U19714 (N_19714,N_18845,N_18659);
nand U19715 (N_19715,N_18036,N_18019);
xor U19716 (N_19716,N_18369,N_18542);
or U19717 (N_19717,N_18070,N_18097);
nand U19718 (N_19718,N_18683,N_18505);
or U19719 (N_19719,N_18330,N_18662);
nand U19720 (N_19720,N_18833,N_18241);
nor U19721 (N_19721,N_18978,N_18120);
and U19722 (N_19722,N_18328,N_18497);
nand U19723 (N_19723,N_18715,N_18890);
and U19724 (N_19724,N_18803,N_18411);
xor U19725 (N_19725,N_18328,N_18560);
or U19726 (N_19726,N_18014,N_18425);
or U19727 (N_19727,N_18479,N_18137);
xnor U19728 (N_19728,N_18786,N_18942);
nand U19729 (N_19729,N_18070,N_18325);
nor U19730 (N_19730,N_18048,N_18130);
xnor U19731 (N_19731,N_18347,N_18360);
and U19732 (N_19732,N_18377,N_18260);
xnor U19733 (N_19733,N_18555,N_18815);
xnor U19734 (N_19734,N_18228,N_18266);
xnor U19735 (N_19735,N_18079,N_18329);
xnor U19736 (N_19736,N_18162,N_18274);
or U19737 (N_19737,N_18225,N_18317);
and U19738 (N_19738,N_18706,N_18763);
nor U19739 (N_19739,N_18067,N_18201);
and U19740 (N_19740,N_18708,N_18620);
nand U19741 (N_19741,N_18208,N_18720);
xor U19742 (N_19742,N_18592,N_18582);
and U19743 (N_19743,N_18834,N_18982);
xnor U19744 (N_19744,N_18366,N_18887);
and U19745 (N_19745,N_18417,N_18940);
or U19746 (N_19746,N_18326,N_18887);
and U19747 (N_19747,N_18193,N_18372);
or U19748 (N_19748,N_18521,N_18289);
nand U19749 (N_19749,N_18290,N_18837);
nor U19750 (N_19750,N_18046,N_18210);
nand U19751 (N_19751,N_18985,N_18923);
and U19752 (N_19752,N_18277,N_18731);
xnor U19753 (N_19753,N_18156,N_18105);
or U19754 (N_19754,N_18864,N_18264);
nor U19755 (N_19755,N_18468,N_18510);
nand U19756 (N_19756,N_18783,N_18047);
and U19757 (N_19757,N_18973,N_18039);
nand U19758 (N_19758,N_18467,N_18654);
nand U19759 (N_19759,N_18090,N_18778);
or U19760 (N_19760,N_18836,N_18076);
nand U19761 (N_19761,N_18549,N_18327);
and U19762 (N_19762,N_18462,N_18061);
and U19763 (N_19763,N_18597,N_18554);
or U19764 (N_19764,N_18691,N_18370);
and U19765 (N_19765,N_18328,N_18498);
nor U19766 (N_19766,N_18902,N_18761);
or U19767 (N_19767,N_18391,N_18153);
nor U19768 (N_19768,N_18398,N_18560);
and U19769 (N_19769,N_18648,N_18089);
nor U19770 (N_19770,N_18426,N_18355);
xnor U19771 (N_19771,N_18221,N_18760);
or U19772 (N_19772,N_18366,N_18983);
nand U19773 (N_19773,N_18204,N_18968);
nand U19774 (N_19774,N_18682,N_18067);
or U19775 (N_19775,N_18297,N_18458);
and U19776 (N_19776,N_18624,N_18096);
xnor U19777 (N_19777,N_18208,N_18573);
and U19778 (N_19778,N_18943,N_18388);
nor U19779 (N_19779,N_18924,N_18542);
nand U19780 (N_19780,N_18877,N_18134);
xor U19781 (N_19781,N_18074,N_18312);
nand U19782 (N_19782,N_18445,N_18637);
and U19783 (N_19783,N_18752,N_18271);
or U19784 (N_19784,N_18709,N_18864);
nand U19785 (N_19785,N_18332,N_18073);
and U19786 (N_19786,N_18447,N_18087);
and U19787 (N_19787,N_18386,N_18350);
nand U19788 (N_19788,N_18171,N_18728);
nor U19789 (N_19789,N_18452,N_18035);
nor U19790 (N_19790,N_18247,N_18979);
xor U19791 (N_19791,N_18963,N_18734);
and U19792 (N_19792,N_18913,N_18565);
nand U19793 (N_19793,N_18121,N_18397);
nor U19794 (N_19794,N_18861,N_18209);
or U19795 (N_19795,N_18759,N_18942);
nor U19796 (N_19796,N_18195,N_18618);
nand U19797 (N_19797,N_18766,N_18623);
nor U19798 (N_19798,N_18504,N_18029);
xor U19799 (N_19799,N_18845,N_18853);
and U19800 (N_19800,N_18084,N_18546);
xnor U19801 (N_19801,N_18330,N_18829);
nor U19802 (N_19802,N_18305,N_18797);
xor U19803 (N_19803,N_18239,N_18392);
and U19804 (N_19804,N_18853,N_18113);
nor U19805 (N_19805,N_18234,N_18432);
or U19806 (N_19806,N_18693,N_18788);
nor U19807 (N_19807,N_18440,N_18531);
or U19808 (N_19808,N_18313,N_18064);
nor U19809 (N_19809,N_18526,N_18056);
and U19810 (N_19810,N_18269,N_18856);
nor U19811 (N_19811,N_18892,N_18521);
xor U19812 (N_19812,N_18785,N_18416);
nand U19813 (N_19813,N_18506,N_18621);
nand U19814 (N_19814,N_18543,N_18569);
or U19815 (N_19815,N_18778,N_18903);
and U19816 (N_19816,N_18166,N_18902);
or U19817 (N_19817,N_18656,N_18372);
and U19818 (N_19818,N_18111,N_18865);
nor U19819 (N_19819,N_18227,N_18296);
nor U19820 (N_19820,N_18065,N_18564);
xnor U19821 (N_19821,N_18238,N_18799);
or U19822 (N_19822,N_18326,N_18724);
nand U19823 (N_19823,N_18686,N_18663);
nor U19824 (N_19824,N_18853,N_18240);
or U19825 (N_19825,N_18215,N_18554);
nor U19826 (N_19826,N_18185,N_18866);
nor U19827 (N_19827,N_18356,N_18677);
xnor U19828 (N_19828,N_18295,N_18575);
nor U19829 (N_19829,N_18524,N_18511);
and U19830 (N_19830,N_18780,N_18745);
nand U19831 (N_19831,N_18610,N_18731);
nand U19832 (N_19832,N_18232,N_18547);
nand U19833 (N_19833,N_18425,N_18342);
and U19834 (N_19834,N_18118,N_18676);
xnor U19835 (N_19835,N_18819,N_18016);
xnor U19836 (N_19836,N_18796,N_18571);
and U19837 (N_19837,N_18633,N_18878);
nand U19838 (N_19838,N_18362,N_18904);
or U19839 (N_19839,N_18458,N_18196);
nor U19840 (N_19840,N_18779,N_18702);
and U19841 (N_19841,N_18687,N_18090);
and U19842 (N_19842,N_18622,N_18340);
xor U19843 (N_19843,N_18792,N_18316);
xnor U19844 (N_19844,N_18957,N_18189);
nor U19845 (N_19845,N_18359,N_18758);
nor U19846 (N_19846,N_18586,N_18500);
and U19847 (N_19847,N_18547,N_18017);
nor U19848 (N_19848,N_18652,N_18271);
xor U19849 (N_19849,N_18134,N_18477);
nand U19850 (N_19850,N_18536,N_18894);
and U19851 (N_19851,N_18719,N_18412);
xnor U19852 (N_19852,N_18344,N_18383);
and U19853 (N_19853,N_18112,N_18207);
nand U19854 (N_19854,N_18252,N_18562);
nand U19855 (N_19855,N_18284,N_18509);
and U19856 (N_19856,N_18523,N_18021);
nor U19857 (N_19857,N_18491,N_18311);
xor U19858 (N_19858,N_18646,N_18025);
xor U19859 (N_19859,N_18002,N_18857);
nand U19860 (N_19860,N_18642,N_18212);
nand U19861 (N_19861,N_18238,N_18444);
nand U19862 (N_19862,N_18015,N_18353);
or U19863 (N_19863,N_18462,N_18736);
nand U19864 (N_19864,N_18877,N_18346);
nor U19865 (N_19865,N_18885,N_18777);
nor U19866 (N_19866,N_18251,N_18913);
or U19867 (N_19867,N_18260,N_18580);
xor U19868 (N_19868,N_18151,N_18045);
xor U19869 (N_19869,N_18103,N_18631);
nor U19870 (N_19870,N_18837,N_18686);
nand U19871 (N_19871,N_18716,N_18826);
nand U19872 (N_19872,N_18323,N_18861);
nand U19873 (N_19873,N_18808,N_18046);
nor U19874 (N_19874,N_18540,N_18324);
and U19875 (N_19875,N_18880,N_18394);
nor U19876 (N_19876,N_18818,N_18749);
nor U19877 (N_19877,N_18933,N_18993);
nand U19878 (N_19878,N_18521,N_18590);
or U19879 (N_19879,N_18186,N_18580);
nor U19880 (N_19880,N_18717,N_18160);
nor U19881 (N_19881,N_18656,N_18228);
nand U19882 (N_19882,N_18784,N_18423);
or U19883 (N_19883,N_18186,N_18413);
and U19884 (N_19884,N_18005,N_18051);
or U19885 (N_19885,N_18285,N_18874);
and U19886 (N_19886,N_18819,N_18169);
nor U19887 (N_19887,N_18541,N_18730);
xor U19888 (N_19888,N_18250,N_18019);
xor U19889 (N_19889,N_18696,N_18710);
xnor U19890 (N_19890,N_18976,N_18815);
and U19891 (N_19891,N_18563,N_18587);
nand U19892 (N_19892,N_18238,N_18179);
nand U19893 (N_19893,N_18436,N_18101);
or U19894 (N_19894,N_18947,N_18868);
nor U19895 (N_19895,N_18029,N_18177);
nor U19896 (N_19896,N_18513,N_18797);
nand U19897 (N_19897,N_18653,N_18282);
nor U19898 (N_19898,N_18554,N_18211);
or U19899 (N_19899,N_18539,N_18850);
or U19900 (N_19900,N_18501,N_18339);
nand U19901 (N_19901,N_18331,N_18965);
and U19902 (N_19902,N_18336,N_18334);
nand U19903 (N_19903,N_18728,N_18733);
nor U19904 (N_19904,N_18192,N_18965);
nand U19905 (N_19905,N_18405,N_18842);
xnor U19906 (N_19906,N_18668,N_18704);
nor U19907 (N_19907,N_18100,N_18262);
and U19908 (N_19908,N_18682,N_18052);
nor U19909 (N_19909,N_18904,N_18732);
or U19910 (N_19910,N_18855,N_18751);
xor U19911 (N_19911,N_18531,N_18937);
or U19912 (N_19912,N_18782,N_18729);
or U19913 (N_19913,N_18040,N_18581);
nor U19914 (N_19914,N_18137,N_18229);
nand U19915 (N_19915,N_18254,N_18277);
or U19916 (N_19916,N_18880,N_18472);
xor U19917 (N_19917,N_18326,N_18138);
and U19918 (N_19918,N_18452,N_18977);
xnor U19919 (N_19919,N_18695,N_18438);
and U19920 (N_19920,N_18428,N_18540);
and U19921 (N_19921,N_18694,N_18067);
xnor U19922 (N_19922,N_18443,N_18630);
nor U19923 (N_19923,N_18064,N_18188);
and U19924 (N_19924,N_18629,N_18808);
xor U19925 (N_19925,N_18907,N_18157);
xnor U19926 (N_19926,N_18878,N_18718);
xnor U19927 (N_19927,N_18958,N_18294);
nor U19928 (N_19928,N_18841,N_18343);
nor U19929 (N_19929,N_18175,N_18078);
or U19930 (N_19930,N_18662,N_18397);
nand U19931 (N_19931,N_18031,N_18349);
xnor U19932 (N_19932,N_18490,N_18975);
xnor U19933 (N_19933,N_18525,N_18356);
nand U19934 (N_19934,N_18421,N_18547);
nor U19935 (N_19935,N_18049,N_18070);
xnor U19936 (N_19936,N_18575,N_18302);
xnor U19937 (N_19937,N_18132,N_18677);
xnor U19938 (N_19938,N_18753,N_18089);
xnor U19939 (N_19939,N_18516,N_18152);
xnor U19940 (N_19940,N_18815,N_18032);
xor U19941 (N_19941,N_18975,N_18521);
or U19942 (N_19942,N_18386,N_18906);
xnor U19943 (N_19943,N_18962,N_18903);
or U19944 (N_19944,N_18712,N_18748);
and U19945 (N_19945,N_18392,N_18676);
and U19946 (N_19946,N_18262,N_18809);
or U19947 (N_19947,N_18260,N_18003);
and U19948 (N_19948,N_18330,N_18824);
and U19949 (N_19949,N_18914,N_18398);
nand U19950 (N_19950,N_18186,N_18937);
xnor U19951 (N_19951,N_18205,N_18014);
and U19952 (N_19952,N_18636,N_18560);
nor U19953 (N_19953,N_18270,N_18778);
and U19954 (N_19954,N_18771,N_18383);
nor U19955 (N_19955,N_18976,N_18338);
nand U19956 (N_19956,N_18568,N_18940);
or U19957 (N_19957,N_18510,N_18302);
or U19958 (N_19958,N_18085,N_18398);
nor U19959 (N_19959,N_18574,N_18360);
or U19960 (N_19960,N_18412,N_18592);
nand U19961 (N_19961,N_18432,N_18465);
and U19962 (N_19962,N_18381,N_18751);
nor U19963 (N_19963,N_18409,N_18578);
nor U19964 (N_19964,N_18980,N_18371);
xor U19965 (N_19965,N_18843,N_18972);
nor U19966 (N_19966,N_18320,N_18101);
xor U19967 (N_19967,N_18095,N_18046);
nor U19968 (N_19968,N_18146,N_18430);
and U19969 (N_19969,N_18238,N_18157);
and U19970 (N_19970,N_18543,N_18414);
nand U19971 (N_19971,N_18296,N_18761);
nor U19972 (N_19972,N_18844,N_18780);
nor U19973 (N_19973,N_18030,N_18797);
nor U19974 (N_19974,N_18605,N_18854);
nor U19975 (N_19975,N_18046,N_18666);
xor U19976 (N_19976,N_18408,N_18086);
nor U19977 (N_19977,N_18067,N_18447);
nor U19978 (N_19978,N_18884,N_18405);
nand U19979 (N_19979,N_18107,N_18513);
or U19980 (N_19980,N_18272,N_18324);
or U19981 (N_19981,N_18923,N_18089);
and U19982 (N_19982,N_18102,N_18706);
nand U19983 (N_19983,N_18191,N_18434);
and U19984 (N_19984,N_18638,N_18714);
nor U19985 (N_19985,N_18898,N_18201);
or U19986 (N_19986,N_18976,N_18893);
or U19987 (N_19987,N_18908,N_18474);
xor U19988 (N_19988,N_18013,N_18146);
or U19989 (N_19989,N_18522,N_18820);
xnor U19990 (N_19990,N_18716,N_18879);
and U19991 (N_19991,N_18125,N_18658);
xor U19992 (N_19992,N_18495,N_18080);
nor U19993 (N_19993,N_18359,N_18198);
nand U19994 (N_19994,N_18806,N_18666);
nand U19995 (N_19995,N_18884,N_18447);
nand U19996 (N_19996,N_18736,N_18640);
nand U19997 (N_19997,N_18762,N_18858);
xnor U19998 (N_19998,N_18898,N_18512);
nor U19999 (N_19999,N_18111,N_18408);
nor UO_0 (O_0,N_19738,N_19710);
nand UO_1 (O_1,N_19639,N_19648);
or UO_2 (O_2,N_19553,N_19592);
nand UO_3 (O_3,N_19248,N_19962);
nand UO_4 (O_4,N_19767,N_19845);
xnor UO_5 (O_5,N_19799,N_19785);
and UO_6 (O_6,N_19963,N_19159);
xor UO_7 (O_7,N_19319,N_19964);
nand UO_8 (O_8,N_19714,N_19961);
and UO_9 (O_9,N_19383,N_19076);
nand UO_10 (O_10,N_19158,N_19462);
or UO_11 (O_11,N_19361,N_19720);
or UO_12 (O_12,N_19184,N_19444);
xnor UO_13 (O_13,N_19906,N_19100);
and UO_14 (O_14,N_19448,N_19751);
xnor UO_15 (O_15,N_19627,N_19487);
xor UO_16 (O_16,N_19849,N_19669);
nor UO_17 (O_17,N_19632,N_19951);
xor UO_18 (O_18,N_19792,N_19994);
or UO_19 (O_19,N_19607,N_19441);
nor UO_20 (O_20,N_19117,N_19514);
nand UO_21 (O_21,N_19629,N_19063);
nand UO_22 (O_22,N_19736,N_19716);
nand UO_23 (O_23,N_19612,N_19346);
and UO_24 (O_24,N_19357,N_19491);
or UO_25 (O_25,N_19153,N_19301);
or UO_26 (O_26,N_19608,N_19379);
nand UO_27 (O_27,N_19615,N_19650);
nor UO_28 (O_28,N_19231,N_19304);
or UO_29 (O_29,N_19257,N_19925);
and UO_30 (O_30,N_19399,N_19011);
nand UO_31 (O_31,N_19423,N_19705);
nand UO_32 (O_32,N_19679,N_19960);
and UO_33 (O_33,N_19474,N_19932);
xor UO_34 (O_34,N_19801,N_19146);
nand UO_35 (O_35,N_19056,N_19111);
and UO_36 (O_36,N_19038,N_19182);
xor UO_37 (O_37,N_19277,N_19136);
or UO_38 (O_38,N_19032,N_19835);
or UO_39 (O_39,N_19765,N_19978);
or UO_40 (O_40,N_19531,N_19701);
and UO_41 (O_41,N_19034,N_19311);
or UO_42 (O_42,N_19074,N_19019);
and UO_43 (O_43,N_19559,N_19855);
and UO_44 (O_44,N_19786,N_19910);
or UO_45 (O_45,N_19838,N_19299);
and UO_46 (O_46,N_19478,N_19308);
nand UO_47 (O_47,N_19846,N_19413);
xor UO_48 (O_48,N_19393,N_19348);
nand UO_49 (O_49,N_19293,N_19740);
and UO_50 (O_50,N_19505,N_19524);
nor UO_51 (O_51,N_19519,N_19349);
nor UO_52 (O_52,N_19713,N_19689);
xor UO_53 (O_53,N_19094,N_19986);
xor UO_54 (O_54,N_19848,N_19018);
and UO_55 (O_55,N_19582,N_19195);
or UO_56 (O_56,N_19270,N_19084);
xor UO_57 (O_57,N_19120,N_19709);
nand UO_58 (O_58,N_19633,N_19587);
and UO_59 (O_59,N_19722,N_19321);
nand UO_60 (O_60,N_19699,N_19000);
and UO_61 (O_61,N_19567,N_19667);
nand UO_62 (O_62,N_19224,N_19946);
and UO_63 (O_63,N_19661,N_19354);
and UO_64 (O_64,N_19427,N_19678);
and UO_65 (O_65,N_19563,N_19013);
xor UO_66 (O_66,N_19671,N_19461);
xor UO_67 (O_67,N_19764,N_19598);
xor UO_68 (O_68,N_19175,N_19205);
nor UO_69 (O_69,N_19398,N_19258);
or UO_70 (O_70,N_19930,N_19316);
nor UO_71 (O_71,N_19318,N_19768);
and UO_72 (O_72,N_19261,N_19766);
or UO_73 (O_73,N_19918,N_19334);
xor UO_74 (O_74,N_19203,N_19305);
and UO_75 (O_75,N_19450,N_19811);
xnor UO_76 (O_76,N_19174,N_19275);
xnor UO_77 (O_77,N_19233,N_19818);
and UO_78 (O_78,N_19244,N_19538);
nand UO_79 (O_79,N_19754,N_19351);
nor UO_80 (O_80,N_19565,N_19700);
nor UO_81 (O_81,N_19337,N_19602);
and UO_82 (O_82,N_19280,N_19437);
nand UO_83 (O_83,N_19016,N_19603);
or UO_84 (O_84,N_19359,N_19360);
nand UO_85 (O_85,N_19472,N_19414);
nor UO_86 (O_86,N_19186,N_19228);
and UO_87 (O_87,N_19167,N_19252);
nand UO_88 (O_88,N_19358,N_19924);
or UO_89 (O_89,N_19036,N_19073);
xor UO_90 (O_90,N_19396,N_19495);
xor UO_91 (O_91,N_19421,N_19613);
nor UO_92 (O_92,N_19080,N_19193);
or UO_93 (O_93,N_19243,N_19665);
and UO_94 (O_94,N_19861,N_19515);
nand UO_95 (O_95,N_19901,N_19520);
nand UO_96 (O_96,N_19759,N_19870);
or UO_97 (O_97,N_19366,N_19571);
or UO_98 (O_98,N_19131,N_19529);
and UO_99 (O_99,N_19498,N_19057);
nor UO_100 (O_100,N_19171,N_19546);
xor UO_101 (O_101,N_19002,N_19819);
and UO_102 (O_102,N_19580,N_19331);
or UO_103 (O_103,N_19757,N_19353);
nor UO_104 (O_104,N_19206,N_19152);
xor UO_105 (O_105,N_19548,N_19105);
and UO_106 (O_106,N_19099,N_19109);
or UO_107 (O_107,N_19418,N_19187);
nor UO_108 (O_108,N_19460,N_19232);
nand UO_109 (O_109,N_19822,N_19770);
and UO_110 (O_110,N_19547,N_19616);
xor UO_111 (O_111,N_19513,N_19047);
nand UO_112 (O_112,N_19813,N_19126);
nor UO_113 (O_113,N_19226,N_19332);
and UO_114 (O_114,N_19464,N_19691);
or UO_115 (O_115,N_19907,N_19431);
xnor UO_116 (O_116,N_19343,N_19771);
nor UO_117 (O_117,N_19997,N_19688);
nor UO_118 (O_118,N_19412,N_19726);
and UO_119 (O_119,N_19895,N_19268);
nor UO_120 (O_120,N_19509,N_19935);
nand UO_121 (O_121,N_19637,N_19375);
and UO_122 (O_122,N_19718,N_19336);
xor UO_123 (O_123,N_19079,N_19255);
nor UO_124 (O_124,N_19609,N_19492);
or UO_125 (O_125,N_19055,N_19647);
or UO_126 (O_126,N_19941,N_19769);
nand UO_127 (O_127,N_19237,N_19267);
xnor UO_128 (O_128,N_19512,N_19338);
nor UO_129 (O_129,N_19683,N_19664);
or UO_130 (O_130,N_19292,N_19116);
and UO_131 (O_131,N_19342,N_19972);
nor UO_132 (O_132,N_19216,N_19752);
nand UO_133 (O_133,N_19622,N_19614);
or UO_134 (O_134,N_19674,N_19681);
or UO_135 (O_135,N_19842,N_19004);
nand UO_136 (O_136,N_19409,N_19408);
nand UO_137 (O_137,N_19090,N_19516);
xor UO_138 (O_138,N_19108,N_19863);
and UO_139 (O_139,N_19922,N_19411);
nor UO_140 (O_140,N_19455,N_19912);
or UO_141 (O_141,N_19287,N_19154);
or UO_142 (O_142,N_19178,N_19776);
nand UO_143 (O_143,N_19051,N_19536);
or UO_144 (O_144,N_19077,N_19052);
nor UO_145 (O_145,N_19724,N_19812);
and UO_146 (O_146,N_19115,N_19630);
xnor UO_147 (O_147,N_19191,N_19298);
or UO_148 (O_148,N_19641,N_19549);
xnor UO_149 (O_149,N_19953,N_19033);
xor UO_150 (O_150,N_19163,N_19254);
xor UO_151 (O_151,N_19217,N_19003);
nand UO_152 (O_152,N_19269,N_19352);
or UO_153 (O_153,N_19875,N_19309);
and UO_154 (O_154,N_19715,N_19561);
or UO_155 (O_155,N_19528,N_19939);
or UO_156 (O_156,N_19410,N_19943);
nor UO_157 (O_157,N_19112,N_19893);
or UO_158 (O_158,N_19753,N_19075);
nor UO_159 (O_159,N_19887,N_19458);
nor UO_160 (O_160,N_19852,N_19646);
or UO_161 (O_161,N_19314,N_19282);
and UO_162 (O_162,N_19839,N_19834);
and UO_163 (O_163,N_19285,N_19824);
or UO_164 (O_164,N_19929,N_19390);
or UO_165 (O_165,N_19795,N_19595);
nor UO_166 (O_166,N_19170,N_19235);
and UO_167 (O_167,N_19685,N_19222);
or UO_168 (O_168,N_19263,N_19329);
or UO_169 (O_169,N_19374,N_19067);
xor UO_170 (O_170,N_19728,N_19467);
and UO_171 (O_171,N_19434,N_19151);
xor UO_172 (O_172,N_19281,N_19921);
nor UO_173 (O_173,N_19804,N_19327);
nand UO_174 (O_174,N_19082,N_19652);
nand UO_175 (O_175,N_19485,N_19101);
xnor UO_176 (O_176,N_19891,N_19162);
and UO_177 (O_177,N_19212,N_19307);
or UO_178 (O_178,N_19843,N_19750);
and UO_179 (O_179,N_19719,N_19916);
nor UO_180 (O_180,N_19208,N_19310);
nor UO_181 (O_181,N_19578,N_19975);
and UO_182 (O_182,N_19706,N_19790);
and UO_183 (O_183,N_19594,N_19266);
nor UO_184 (O_184,N_19695,N_19827);
xor UO_185 (O_185,N_19289,N_19473);
xor UO_186 (O_186,N_19980,N_19059);
nand UO_187 (O_187,N_19847,N_19982);
and UO_188 (O_188,N_19430,N_19103);
nand UO_189 (O_189,N_19780,N_19676);
xnor UO_190 (O_190,N_19241,N_19959);
and UO_191 (O_191,N_19940,N_19821);
or UO_192 (O_192,N_19831,N_19890);
nor UO_193 (O_193,N_19976,N_19139);
or UO_194 (O_194,N_19783,N_19039);
or UO_195 (O_195,N_19405,N_19143);
nand UO_196 (O_196,N_19942,N_19800);
nor UO_197 (O_197,N_19370,N_19569);
and UO_198 (O_198,N_19755,N_19192);
nand UO_199 (O_199,N_19945,N_19868);
nand UO_200 (O_200,N_19885,N_19954);
or UO_201 (O_201,N_19356,N_19742);
nor UO_202 (O_202,N_19197,N_19570);
and UO_203 (O_203,N_19137,N_19601);
nand UO_204 (O_204,N_19198,N_19554);
and UO_205 (O_205,N_19294,N_19808);
or UO_206 (O_206,N_19006,N_19113);
nor UO_207 (O_207,N_19948,N_19576);
or UO_208 (O_208,N_19897,N_19588);
nor UO_209 (O_209,N_19042,N_19325);
nor UO_210 (O_210,N_19854,N_19097);
or UO_211 (O_211,N_19867,N_19172);
or UO_212 (O_212,N_19523,N_19482);
nand UO_213 (O_213,N_19905,N_19904);
or UO_214 (O_214,N_19892,N_19522);
and UO_215 (O_215,N_19560,N_19256);
or UO_216 (O_216,N_19881,N_19210);
nor UO_217 (O_217,N_19746,N_19617);
nand UO_218 (O_218,N_19017,N_19511);
xor UO_219 (O_219,N_19551,N_19864);
nor UO_220 (O_220,N_19107,N_19322);
nand UO_221 (O_221,N_19218,N_19748);
nor UO_222 (O_222,N_19062,N_19694);
nand UO_223 (O_223,N_19541,N_19635);
and UO_224 (O_224,N_19010,N_19704);
xor UO_225 (O_225,N_19335,N_19072);
or UO_226 (O_226,N_19979,N_19091);
nor UO_227 (O_227,N_19734,N_19283);
nor UO_228 (O_228,N_19250,N_19466);
xor UO_229 (O_229,N_19973,N_19631);
or UO_230 (O_230,N_19532,N_19568);
nor UO_231 (O_231,N_19687,N_19138);
xor UO_232 (O_232,N_19230,N_19401);
or UO_233 (O_233,N_19686,N_19121);
and UO_234 (O_234,N_19447,N_19376);
nor UO_235 (O_235,N_19628,N_19653);
nand UO_236 (O_236,N_19106,N_19562);
xnor UO_237 (O_237,N_19791,N_19542);
nand UO_238 (O_238,N_19046,N_19775);
or UO_239 (O_239,N_19911,N_19341);
and UO_240 (O_240,N_19128,N_19773);
and UO_241 (O_241,N_19041,N_19874);
nor UO_242 (O_242,N_19851,N_19435);
and UO_243 (O_243,N_19898,N_19219);
or UO_244 (O_244,N_19288,N_19150);
and UO_245 (O_245,N_19001,N_19480);
and UO_246 (O_246,N_19324,N_19225);
and UO_247 (O_247,N_19098,N_19213);
or UO_248 (O_248,N_19087,N_19284);
nand UO_249 (O_249,N_19659,N_19952);
xor UO_250 (O_250,N_19050,N_19733);
or UO_251 (O_251,N_19988,N_19276);
and UO_252 (O_252,N_19415,N_19499);
nand UO_253 (O_253,N_19645,N_19806);
and UO_254 (O_254,N_19272,N_19743);
nor UO_255 (O_255,N_19265,N_19672);
nand UO_256 (O_256,N_19832,N_19888);
or UO_257 (O_257,N_19428,N_19995);
xnor UO_258 (O_258,N_19816,N_19999);
nand UO_259 (O_259,N_19744,N_19302);
nor UO_260 (O_260,N_19496,N_19802);
nand UO_261 (O_261,N_19957,N_19749);
xnor UO_262 (O_262,N_19481,N_19558);
nor UO_263 (O_263,N_19488,N_19774);
nand UO_264 (O_264,N_19841,N_19596);
xor UO_265 (O_265,N_19389,N_19955);
nor UO_266 (O_266,N_19692,N_19384);
nor UO_267 (O_267,N_19229,N_19015);
xnor UO_268 (O_268,N_19909,N_19782);
and UO_269 (O_269,N_19573,N_19610);
nor UO_270 (O_270,N_19456,N_19236);
or UO_271 (O_271,N_19419,N_19820);
nor UO_272 (O_272,N_19539,N_19618);
and UO_273 (O_273,N_19031,N_19371);
xnor UO_274 (O_274,N_19798,N_19054);
nand UO_275 (O_275,N_19443,N_19395);
nand UO_276 (O_276,N_19971,N_19833);
nand UO_277 (O_277,N_19142,N_19040);
nor UO_278 (O_278,N_19998,N_19853);
nand UO_279 (O_279,N_19927,N_19703);
xor UO_280 (O_280,N_19424,N_19966);
nor UO_281 (O_281,N_19214,N_19459);
or UO_282 (O_282,N_19914,N_19134);
or UO_283 (O_283,N_19871,N_19970);
nand UO_284 (O_284,N_19166,N_19027);
nor UO_285 (O_285,N_19735,N_19044);
nor UO_286 (O_286,N_19207,N_19124);
or UO_287 (O_287,N_19673,N_19660);
xor UO_288 (O_288,N_19234,N_19894);
or UO_289 (O_289,N_19949,N_19240);
nand UO_290 (O_290,N_19259,N_19974);
nand UO_291 (O_291,N_19920,N_19081);
nand UO_292 (O_292,N_19968,N_19156);
or UO_293 (O_293,N_19944,N_19586);
xor UO_294 (O_294,N_19119,N_19312);
and UO_295 (O_295,N_19506,N_19446);
or UO_296 (O_296,N_19037,N_19377);
nor UO_297 (O_297,N_19278,N_19862);
and UO_298 (O_298,N_19026,N_19525);
and UO_299 (O_299,N_19540,N_19707);
or UO_300 (O_300,N_19494,N_19741);
nand UO_301 (O_301,N_19526,N_19860);
or UO_302 (O_302,N_19756,N_19879);
xnor UO_303 (O_303,N_19391,N_19527);
nand UO_304 (O_304,N_19344,N_19043);
nand UO_305 (O_305,N_19656,N_19597);
xnor UO_306 (O_306,N_19083,N_19378);
or UO_307 (O_307,N_19130,N_19238);
nand UO_308 (O_308,N_19577,N_19271);
or UO_309 (O_309,N_19157,N_19878);
nand UO_310 (O_310,N_19303,N_19828);
nand UO_311 (O_311,N_19385,N_19684);
nor UO_312 (O_312,N_19199,N_19859);
nand UO_313 (O_313,N_19876,N_19696);
nand UO_314 (O_314,N_19347,N_19449);
nor UO_315 (O_315,N_19809,N_19711);
xnor UO_316 (O_316,N_19295,N_19552);
xor UO_317 (O_317,N_19251,N_19877);
xor UO_318 (O_318,N_19457,N_19717);
or UO_319 (O_319,N_19416,N_19122);
and UO_320 (O_320,N_19028,N_19145);
and UO_321 (O_321,N_19938,N_19535);
nand UO_322 (O_322,N_19165,N_19180);
or UO_323 (O_323,N_19179,N_19368);
or UO_324 (O_324,N_19024,N_19127);
and UO_325 (O_325,N_19865,N_19593);
or UO_326 (O_326,N_19844,N_19397);
or UO_327 (O_327,N_19173,N_19500);
and UO_328 (O_328,N_19483,N_19135);
xor UO_329 (O_329,N_19566,N_19432);
xnor UO_330 (O_330,N_19005,N_19814);
or UO_331 (O_331,N_19984,N_19758);
nor UO_332 (O_332,N_19697,N_19985);
xnor UO_333 (O_333,N_19078,N_19950);
xor UO_334 (O_334,N_19315,N_19731);
and UO_335 (O_335,N_19185,N_19260);
nor UO_336 (O_336,N_19221,N_19992);
xor UO_337 (O_337,N_19089,N_19297);
nor UO_338 (O_338,N_19947,N_19682);
and UO_339 (O_339,N_19463,N_19917);
and UO_340 (O_340,N_19708,N_19453);
or UO_341 (O_341,N_19339,N_19320);
nand UO_342 (O_342,N_19058,N_19903);
nand UO_343 (O_343,N_19247,N_19658);
nand UO_344 (O_344,N_19147,N_19407);
xnor UO_345 (O_345,N_19246,N_19438);
xnor UO_346 (O_346,N_19784,N_19330);
or UO_347 (O_347,N_19702,N_19977);
or UO_348 (O_348,N_19468,N_19636);
and UO_349 (O_349,N_19118,N_19189);
xnor UO_350 (O_350,N_19394,N_19886);
nor UO_351 (O_351,N_19279,N_19923);
and UO_352 (O_352,N_19388,N_19882);
or UO_353 (O_353,N_19584,N_19557);
and UO_354 (O_354,N_19404,N_19729);
and UO_355 (O_355,N_19837,N_19555);
and UO_356 (O_356,N_19023,N_19521);
nand UO_357 (O_357,N_19045,N_19144);
nor UO_358 (O_358,N_19326,N_19534);
nor UO_359 (O_359,N_19363,N_19095);
or UO_360 (O_360,N_19429,N_19132);
xor UO_361 (O_361,N_19902,N_19096);
xor UO_362 (O_362,N_19274,N_19110);
xnor UO_363 (O_363,N_19591,N_19958);
nand UO_364 (O_364,N_19967,N_19668);
nor UO_365 (O_365,N_19889,N_19012);
and UO_366 (O_366,N_19605,N_19915);
and UO_367 (O_367,N_19008,N_19931);
nor UO_368 (O_368,N_19620,N_19657);
and UO_369 (O_369,N_19933,N_19747);
nor UO_370 (O_370,N_19623,N_19850);
and UO_371 (O_371,N_19544,N_19662);
nand UO_372 (O_372,N_19543,N_19392);
and UO_373 (O_373,N_19956,N_19402);
xor UO_374 (O_374,N_19919,N_19670);
or UO_375 (O_375,N_19497,N_19666);
and UO_376 (O_376,N_19085,N_19486);
nand UO_377 (O_377,N_19066,N_19493);
or UO_378 (O_378,N_19009,N_19989);
nand UO_379 (O_379,N_19102,N_19264);
or UO_380 (O_380,N_19723,N_19872);
and UO_381 (O_381,N_19209,N_19680);
nand UO_382 (O_382,N_19510,N_19417);
nand UO_383 (O_383,N_19638,N_19364);
nor UO_384 (O_384,N_19420,N_19725);
nand UO_385 (O_385,N_19440,N_19590);
nand UO_386 (O_386,N_19869,N_19654);
nor UO_387 (O_387,N_19634,N_19550);
and UO_388 (O_388,N_19760,N_19796);
xor UO_389 (O_389,N_19857,N_19690);
nor UO_390 (O_390,N_19899,N_19426);
and UO_391 (O_391,N_19065,N_19140);
nor UO_392 (O_392,N_19035,N_19323);
and UO_393 (O_393,N_19369,N_19655);
nand UO_394 (O_394,N_19200,N_19503);
xnor UO_395 (O_395,N_19161,N_19141);
and UO_396 (O_396,N_19245,N_19908);
xor UO_397 (O_397,N_19425,N_19183);
or UO_398 (O_398,N_19242,N_19778);
xor UO_399 (O_399,N_19149,N_19965);
nand UO_400 (O_400,N_19625,N_19204);
or UO_401 (O_401,N_19517,N_19489);
nand UO_402 (O_402,N_19007,N_19061);
xor UO_403 (O_403,N_19380,N_19333);
xnor UO_404 (O_404,N_19730,N_19502);
nor UO_405 (O_405,N_19169,N_19317);
nand UO_406 (O_406,N_19433,N_19470);
xnor UO_407 (O_407,N_19286,N_19585);
or UO_408 (O_408,N_19788,N_19781);
or UO_409 (O_409,N_19693,N_19545);
and UO_410 (O_410,N_19442,N_19249);
xor UO_411 (O_411,N_19640,N_19934);
nand UO_412 (O_412,N_19350,N_19196);
or UO_413 (O_413,N_19574,N_19779);
nand UO_414 (O_414,N_19190,N_19148);
and UO_415 (O_415,N_19880,N_19340);
xnor UO_416 (O_416,N_19807,N_19365);
and UO_417 (O_417,N_19611,N_19518);
xnor UO_418 (O_418,N_19530,N_19194);
nor UO_419 (O_419,N_19070,N_19300);
and UO_420 (O_420,N_19030,N_19589);
xnor UO_421 (O_421,N_19600,N_19712);
and UO_422 (O_422,N_19581,N_19291);
xnor UO_423 (O_423,N_19188,N_19071);
and UO_424 (O_424,N_19793,N_19810);
xor UO_425 (O_425,N_19465,N_19490);
xor UO_426 (O_426,N_19983,N_19176);
nand UO_427 (O_427,N_19858,N_19677);
xnor UO_428 (O_428,N_19129,N_19884);
nor UO_429 (O_429,N_19104,N_19092);
nand UO_430 (O_430,N_19387,N_19164);
nor UO_431 (O_431,N_19619,N_19533);
nor UO_432 (O_432,N_19866,N_19313);
nor UO_433 (O_433,N_19829,N_19762);
or UO_434 (O_434,N_19475,N_19649);
and UO_435 (O_435,N_19290,N_19406);
or UO_436 (O_436,N_19823,N_19020);
nor UO_437 (O_437,N_19403,N_19471);
or UO_438 (O_438,N_19201,N_19202);
or UO_439 (O_439,N_19996,N_19022);
or UO_440 (O_440,N_19926,N_19991);
and UO_441 (O_441,N_19830,N_19761);
and UO_442 (O_442,N_19123,N_19273);
and UO_443 (O_443,N_19355,N_19873);
or UO_444 (O_444,N_19896,N_19064);
or UO_445 (O_445,N_19732,N_19160);
nor UO_446 (O_446,N_19253,N_19797);
nand UO_447 (O_447,N_19624,N_19721);
nor UO_448 (O_448,N_19069,N_19382);
nand UO_449 (O_449,N_19088,N_19981);
xor UO_450 (O_450,N_19029,N_19501);
nand UO_451 (O_451,N_19439,N_19060);
xnor UO_452 (O_452,N_19227,N_19599);
and UO_453 (O_453,N_19913,N_19476);
nor UO_454 (O_454,N_19579,N_19386);
nand UO_455 (O_455,N_19133,N_19987);
nor UO_456 (O_456,N_19651,N_19296);
or UO_457 (O_457,N_19445,N_19928);
xnor UO_458 (O_458,N_19817,N_19484);
or UO_459 (O_459,N_19177,N_19025);
or UO_460 (O_460,N_19422,N_19239);
nand UO_461 (O_461,N_19990,N_19621);
xnor UO_462 (O_462,N_19815,N_19745);
or UO_463 (O_463,N_19936,N_19373);
nor UO_464 (O_464,N_19727,N_19856);
nor UO_465 (O_465,N_19763,N_19805);
xnor UO_466 (O_466,N_19572,N_19093);
and UO_467 (O_467,N_19479,N_19372);
or UO_468 (O_468,N_19737,N_19537);
nand UO_469 (O_469,N_19504,N_19086);
xnor UO_470 (O_470,N_19223,N_19606);
nor UO_471 (O_471,N_19789,N_19068);
nor UO_472 (O_472,N_19211,N_19826);
nand UO_473 (O_473,N_19626,N_19168);
nor UO_474 (O_474,N_19400,N_19803);
and UO_475 (O_475,N_19675,N_19306);
and UO_476 (O_476,N_19114,N_19739);
xor UO_477 (O_477,N_19698,N_19825);
or UO_478 (O_478,N_19345,N_19155);
xor UO_479 (O_479,N_19993,N_19049);
or UO_480 (O_480,N_19508,N_19794);
and UO_481 (O_481,N_19014,N_19181);
or UO_482 (O_482,N_19452,N_19469);
nand UO_483 (O_483,N_19937,N_19777);
and UO_484 (O_484,N_19215,N_19836);
or UO_485 (O_485,N_19787,N_19642);
or UO_486 (O_486,N_19840,N_19556);
xor UO_487 (O_487,N_19772,N_19575);
nor UO_488 (O_488,N_19564,N_19262);
or UO_489 (O_489,N_19604,N_19644);
nor UO_490 (O_490,N_19436,N_19381);
nor UO_491 (O_491,N_19477,N_19900);
or UO_492 (O_492,N_19583,N_19328);
nor UO_493 (O_493,N_19507,N_19048);
nand UO_494 (O_494,N_19663,N_19220);
or UO_495 (O_495,N_19053,N_19367);
and UO_496 (O_496,N_19969,N_19021);
nor UO_497 (O_497,N_19125,N_19454);
xor UO_498 (O_498,N_19451,N_19883);
nand UO_499 (O_499,N_19643,N_19362);
nor UO_500 (O_500,N_19999,N_19118);
and UO_501 (O_501,N_19099,N_19674);
xor UO_502 (O_502,N_19456,N_19202);
and UO_503 (O_503,N_19638,N_19601);
nand UO_504 (O_504,N_19547,N_19899);
or UO_505 (O_505,N_19028,N_19529);
xor UO_506 (O_506,N_19680,N_19232);
or UO_507 (O_507,N_19917,N_19999);
nor UO_508 (O_508,N_19468,N_19894);
and UO_509 (O_509,N_19652,N_19411);
nor UO_510 (O_510,N_19166,N_19047);
xor UO_511 (O_511,N_19012,N_19284);
xnor UO_512 (O_512,N_19910,N_19075);
nor UO_513 (O_513,N_19610,N_19715);
nand UO_514 (O_514,N_19298,N_19949);
xnor UO_515 (O_515,N_19100,N_19772);
xor UO_516 (O_516,N_19796,N_19622);
nand UO_517 (O_517,N_19328,N_19155);
nand UO_518 (O_518,N_19899,N_19792);
nand UO_519 (O_519,N_19532,N_19262);
xnor UO_520 (O_520,N_19613,N_19266);
nand UO_521 (O_521,N_19016,N_19643);
nand UO_522 (O_522,N_19217,N_19480);
nand UO_523 (O_523,N_19296,N_19336);
and UO_524 (O_524,N_19083,N_19040);
nand UO_525 (O_525,N_19571,N_19216);
nor UO_526 (O_526,N_19826,N_19633);
or UO_527 (O_527,N_19791,N_19550);
nor UO_528 (O_528,N_19318,N_19365);
nor UO_529 (O_529,N_19731,N_19206);
nand UO_530 (O_530,N_19456,N_19828);
xor UO_531 (O_531,N_19558,N_19820);
or UO_532 (O_532,N_19679,N_19156);
nor UO_533 (O_533,N_19093,N_19868);
xnor UO_534 (O_534,N_19470,N_19471);
nand UO_535 (O_535,N_19271,N_19198);
nor UO_536 (O_536,N_19896,N_19447);
xnor UO_537 (O_537,N_19256,N_19450);
and UO_538 (O_538,N_19379,N_19242);
xnor UO_539 (O_539,N_19988,N_19824);
nor UO_540 (O_540,N_19033,N_19551);
nand UO_541 (O_541,N_19028,N_19604);
nor UO_542 (O_542,N_19840,N_19915);
nand UO_543 (O_543,N_19277,N_19222);
or UO_544 (O_544,N_19323,N_19389);
and UO_545 (O_545,N_19102,N_19448);
xnor UO_546 (O_546,N_19959,N_19942);
nor UO_547 (O_547,N_19649,N_19557);
xor UO_548 (O_548,N_19543,N_19986);
or UO_549 (O_549,N_19038,N_19796);
or UO_550 (O_550,N_19221,N_19597);
or UO_551 (O_551,N_19394,N_19763);
and UO_552 (O_552,N_19546,N_19015);
nand UO_553 (O_553,N_19882,N_19633);
nand UO_554 (O_554,N_19073,N_19575);
xnor UO_555 (O_555,N_19884,N_19276);
and UO_556 (O_556,N_19773,N_19216);
or UO_557 (O_557,N_19577,N_19920);
nand UO_558 (O_558,N_19676,N_19038);
nor UO_559 (O_559,N_19815,N_19114);
nand UO_560 (O_560,N_19333,N_19797);
and UO_561 (O_561,N_19371,N_19364);
and UO_562 (O_562,N_19064,N_19357);
or UO_563 (O_563,N_19213,N_19673);
xor UO_564 (O_564,N_19811,N_19896);
nor UO_565 (O_565,N_19888,N_19635);
or UO_566 (O_566,N_19061,N_19377);
or UO_567 (O_567,N_19294,N_19721);
and UO_568 (O_568,N_19606,N_19357);
and UO_569 (O_569,N_19396,N_19169);
nand UO_570 (O_570,N_19775,N_19418);
xor UO_571 (O_571,N_19504,N_19838);
nor UO_572 (O_572,N_19080,N_19887);
xnor UO_573 (O_573,N_19603,N_19879);
xnor UO_574 (O_574,N_19876,N_19361);
and UO_575 (O_575,N_19906,N_19786);
or UO_576 (O_576,N_19278,N_19307);
nand UO_577 (O_577,N_19581,N_19549);
xor UO_578 (O_578,N_19313,N_19325);
nor UO_579 (O_579,N_19367,N_19972);
nor UO_580 (O_580,N_19705,N_19246);
nand UO_581 (O_581,N_19579,N_19707);
xor UO_582 (O_582,N_19347,N_19673);
nand UO_583 (O_583,N_19378,N_19100);
and UO_584 (O_584,N_19158,N_19805);
or UO_585 (O_585,N_19705,N_19133);
and UO_586 (O_586,N_19441,N_19239);
and UO_587 (O_587,N_19507,N_19804);
or UO_588 (O_588,N_19180,N_19621);
and UO_589 (O_589,N_19474,N_19246);
and UO_590 (O_590,N_19246,N_19609);
xnor UO_591 (O_591,N_19185,N_19327);
nor UO_592 (O_592,N_19798,N_19918);
nand UO_593 (O_593,N_19176,N_19953);
or UO_594 (O_594,N_19191,N_19301);
and UO_595 (O_595,N_19157,N_19191);
nor UO_596 (O_596,N_19806,N_19925);
xnor UO_597 (O_597,N_19615,N_19279);
xor UO_598 (O_598,N_19513,N_19870);
nor UO_599 (O_599,N_19946,N_19581);
xnor UO_600 (O_600,N_19672,N_19858);
or UO_601 (O_601,N_19586,N_19530);
nand UO_602 (O_602,N_19835,N_19678);
nor UO_603 (O_603,N_19021,N_19232);
nand UO_604 (O_604,N_19862,N_19161);
nor UO_605 (O_605,N_19472,N_19882);
nand UO_606 (O_606,N_19321,N_19565);
xnor UO_607 (O_607,N_19612,N_19095);
nand UO_608 (O_608,N_19889,N_19534);
nor UO_609 (O_609,N_19431,N_19333);
or UO_610 (O_610,N_19356,N_19721);
and UO_611 (O_611,N_19766,N_19539);
nand UO_612 (O_612,N_19584,N_19667);
and UO_613 (O_613,N_19761,N_19770);
or UO_614 (O_614,N_19760,N_19900);
nor UO_615 (O_615,N_19785,N_19493);
and UO_616 (O_616,N_19052,N_19081);
xor UO_617 (O_617,N_19809,N_19389);
or UO_618 (O_618,N_19727,N_19358);
and UO_619 (O_619,N_19770,N_19875);
nor UO_620 (O_620,N_19044,N_19182);
nor UO_621 (O_621,N_19415,N_19352);
and UO_622 (O_622,N_19418,N_19206);
nor UO_623 (O_623,N_19823,N_19799);
nand UO_624 (O_624,N_19909,N_19620);
nand UO_625 (O_625,N_19727,N_19233);
xnor UO_626 (O_626,N_19122,N_19307);
nand UO_627 (O_627,N_19070,N_19280);
xor UO_628 (O_628,N_19395,N_19303);
nand UO_629 (O_629,N_19752,N_19419);
and UO_630 (O_630,N_19767,N_19630);
xor UO_631 (O_631,N_19342,N_19693);
xor UO_632 (O_632,N_19196,N_19071);
or UO_633 (O_633,N_19063,N_19087);
and UO_634 (O_634,N_19454,N_19819);
and UO_635 (O_635,N_19932,N_19864);
and UO_636 (O_636,N_19649,N_19555);
or UO_637 (O_637,N_19987,N_19681);
and UO_638 (O_638,N_19896,N_19791);
nand UO_639 (O_639,N_19953,N_19100);
or UO_640 (O_640,N_19859,N_19652);
nand UO_641 (O_641,N_19522,N_19429);
nor UO_642 (O_642,N_19125,N_19057);
and UO_643 (O_643,N_19419,N_19340);
xnor UO_644 (O_644,N_19575,N_19741);
nand UO_645 (O_645,N_19717,N_19516);
or UO_646 (O_646,N_19071,N_19978);
nor UO_647 (O_647,N_19190,N_19045);
or UO_648 (O_648,N_19742,N_19309);
xnor UO_649 (O_649,N_19277,N_19766);
nor UO_650 (O_650,N_19331,N_19643);
and UO_651 (O_651,N_19356,N_19033);
nor UO_652 (O_652,N_19088,N_19001);
xor UO_653 (O_653,N_19506,N_19026);
and UO_654 (O_654,N_19856,N_19875);
or UO_655 (O_655,N_19586,N_19388);
xor UO_656 (O_656,N_19799,N_19654);
and UO_657 (O_657,N_19171,N_19330);
nor UO_658 (O_658,N_19618,N_19068);
nand UO_659 (O_659,N_19608,N_19593);
nor UO_660 (O_660,N_19368,N_19026);
or UO_661 (O_661,N_19655,N_19732);
or UO_662 (O_662,N_19334,N_19176);
nor UO_663 (O_663,N_19328,N_19486);
xor UO_664 (O_664,N_19732,N_19120);
and UO_665 (O_665,N_19346,N_19272);
or UO_666 (O_666,N_19547,N_19189);
xnor UO_667 (O_667,N_19066,N_19896);
nor UO_668 (O_668,N_19317,N_19552);
xnor UO_669 (O_669,N_19829,N_19411);
or UO_670 (O_670,N_19667,N_19938);
or UO_671 (O_671,N_19290,N_19997);
xor UO_672 (O_672,N_19554,N_19959);
xor UO_673 (O_673,N_19051,N_19282);
or UO_674 (O_674,N_19322,N_19311);
nor UO_675 (O_675,N_19401,N_19346);
xnor UO_676 (O_676,N_19515,N_19423);
nand UO_677 (O_677,N_19746,N_19649);
or UO_678 (O_678,N_19386,N_19768);
or UO_679 (O_679,N_19690,N_19720);
nor UO_680 (O_680,N_19100,N_19984);
xor UO_681 (O_681,N_19878,N_19908);
and UO_682 (O_682,N_19084,N_19676);
and UO_683 (O_683,N_19375,N_19379);
xnor UO_684 (O_684,N_19448,N_19594);
nor UO_685 (O_685,N_19011,N_19599);
and UO_686 (O_686,N_19298,N_19744);
nand UO_687 (O_687,N_19877,N_19192);
nand UO_688 (O_688,N_19351,N_19070);
or UO_689 (O_689,N_19452,N_19604);
xor UO_690 (O_690,N_19642,N_19375);
xor UO_691 (O_691,N_19415,N_19509);
nor UO_692 (O_692,N_19881,N_19456);
nor UO_693 (O_693,N_19024,N_19215);
nor UO_694 (O_694,N_19068,N_19663);
xnor UO_695 (O_695,N_19867,N_19544);
xor UO_696 (O_696,N_19613,N_19645);
xor UO_697 (O_697,N_19667,N_19921);
xnor UO_698 (O_698,N_19144,N_19242);
nand UO_699 (O_699,N_19058,N_19191);
and UO_700 (O_700,N_19089,N_19925);
nor UO_701 (O_701,N_19633,N_19560);
nand UO_702 (O_702,N_19270,N_19082);
xor UO_703 (O_703,N_19548,N_19601);
nand UO_704 (O_704,N_19571,N_19122);
xor UO_705 (O_705,N_19264,N_19633);
nand UO_706 (O_706,N_19525,N_19927);
nand UO_707 (O_707,N_19405,N_19590);
nand UO_708 (O_708,N_19313,N_19104);
nand UO_709 (O_709,N_19599,N_19822);
or UO_710 (O_710,N_19035,N_19398);
or UO_711 (O_711,N_19437,N_19943);
xor UO_712 (O_712,N_19902,N_19968);
nand UO_713 (O_713,N_19899,N_19919);
xor UO_714 (O_714,N_19209,N_19553);
and UO_715 (O_715,N_19454,N_19700);
and UO_716 (O_716,N_19892,N_19639);
nand UO_717 (O_717,N_19869,N_19283);
nor UO_718 (O_718,N_19622,N_19979);
xnor UO_719 (O_719,N_19346,N_19448);
or UO_720 (O_720,N_19862,N_19532);
or UO_721 (O_721,N_19704,N_19772);
nor UO_722 (O_722,N_19155,N_19043);
nor UO_723 (O_723,N_19245,N_19818);
xor UO_724 (O_724,N_19193,N_19544);
nor UO_725 (O_725,N_19936,N_19260);
nand UO_726 (O_726,N_19024,N_19919);
and UO_727 (O_727,N_19216,N_19016);
nand UO_728 (O_728,N_19783,N_19406);
xor UO_729 (O_729,N_19866,N_19713);
nor UO_730 (O_730,N_19894,N_19212);
nand UO_731 (O_731,N_19527,N_19290);
nor UO_732 (O_732,N_19738,N_19495);
and UO_733 (O_733,N_19735,N_19112);
or UO_734 (O_734,N_19444,N_19984);
and UO_735 (O_735,N_19375,N_19277);
or UO_736 (O_736,N_19568,N_19174);
xor UO_737 (O_737,N_19489,N_19881);
and UO_738 (O_738,N_19129,N_19336);
and UO_739 (O_739,N_19885,N_19156);
nand UO_740 (O_740,N_19456,N_19823);
xor UO_741 (O_741,N_19939,N_19951);
xnor UO_742 (O_742,N_19217,N_19477);
nand UO_743 (O_743,N_19797,N_19164);
nor UO_744 (O_744,N_19880,N_19266);
or UO_745 (O_745,N_19790,N_19567);
xor UO_746 (O_746,N_19085,N_19123);
xor UO_747 (O_747,N_19005,N_19733);
and UO_748 (O_748,N_19472,N_19063);
or UO_749 (O_749,N_19796,N_19572);
and UO_750 (O_750,N_19463,N_19170);
nand UO_751 (O_751,N_19943,N_19032);
nor UO_752 (O_752,N_19095,N_19155);
or UO_753 (O_753,N_19139,N_19988);
and UO_754 (O_754,N_19026,N_19981);
xnor UO_755 (O_755,N_19064,N_19732);
xnor UO_756 (O_756,N_19583,N_19371);
or UO_757 (O_757,N_19345,N_19427);
nand UO_758 (O_758,N_19374,N_19161);
nand UO_759 (O_759,N_19371,N_19956);
or UO_760 (O_760,N_19942,N_19214);
or UO_761 (O_761,N_19903,N_19069);
and UO_762 (O_762,N_19637,N_19201);
and UO_763 (O_763,N_19335,N_19839);
nand UO_764 (O_764,N_19384,N_19357);
or UO_765 (O_765,N_19916,N_19749);
xor UO_766 (O_766,N_19842,N_19673);
or UO_767 (O_767,N_19221,N_19314);
xor UO_768 (O_768,N_19644,N_19738);
nor UO_769 (O_769,N_19065,N_19096);
or UO_770 (O_770,N_19516,N_19357);
xor UO_771 (O_771,N_19438,N_19893);
and UO_772 (O_772,N_19769,N_19343);
or UO_773 (O_773,N_19469,N_19608);
nand UO_774 (O_774,N_19987,N_19263);
or UO_775 (O_775,N_19679,N_19012);
or UO_776 (O_776,N_19167,N_19007);
nor UO_777 (O_777,N_19013,N_19891);
nor UO_778 (O_778,N_19814,N_19380);
xor UO_779 (O_779,N_19420,N_19517);
nor UO_780 (O_780,N_19498,N_19127);
and UO_781 (O_781,N_19015,N_19381);
and UO_782 (O_782,N_19877,N_19091);
xor UO_783 (O_783,N_19858,N_19025);
nand UO_784 (O_784,N_19175,N_19419);
nor UO_785 (O_785,N_19641,N_19466);
nor UO_786 (O_786,N_19019,N_19706);
or UO_787 (O_787,N_19819,N_19309);
and UO_788 (O_788,N_19771,N_19354);
or UO_789 (O_789,N_19774,N_19509);
xnor UO_790 (O_790,N_19498,N_19036);
nand UO_791 (O_791,N_19027,N_19051);
xor UO_792 (O_792,N_19764,N_19879);
xnor UO_793 (O_793,N_19359,N_19220);
nor UO_794 (O_794,N_19432,N_19172);
and UO_795 (O_795,N_19592,N_19295);
and UO_796 (O_796,N_19867,N_19912);
xor UO_797 (O_797,N_19130,N_19284);
nor UO_798 (O_798,N_19478,N_19241);
nor UO_799 (O_799,N_19277,N_19749);
nand UO_800 (O_800,N_19781,N_19557);
and UO_801 (O_801,N_19902,N_19005);
nor UO_802 (O_802,N_19996,N_19435);
and UO_803 (O_803,N_19745,N_19829);
xnor UO_804 (O_804,N_19747,N_19472);
and UO_805 (O_805,N_19231,N_19718);
nand UO_806 (O_806,N_19199,N_19548);
nor UO_807 (O_807,N_19379,N_19121);
and UO_808 (O_808,N_19860,N_19954);
or UO_809 (O_809,N_19325,N_19391);
xnor UO_810 (O_810,N_19285,N_19427);
nor UO_811 (O_811,N_19755,N_19204);
xor UO_812 (O_812,N_19631,N_19808);
nand UO_813 (O_813,N_19571,N_19416);
xor UO_814 (O_814,N_19934,N_19880);
nand UO_815 (O_815,N_19226,N_19882);
nor UO_816 (O_816,N_19228,N_19790);
nor UO_817 (O_817,N_19509,N_19630);
nor UO_818 (O_818,N_19153,N_19726);
nand UO_819 (O_819,N_19729,N_19141);
and UO_820 (O_820,N_19797,N_19808);
nand UO_821 (O_821,N_19983,N_19450);
nor UO_822 (O_822,N_19960,N_19895);
and UO_823 (O_823,N_19863,N_19978);
or UO_824 (O_824,N_19219,N_19340);
nand UO_825 (O_825,N_19317,N_19250);
xor UO_826 (O_826,N_19239,N_19638);
xor UO_827 (O_827,N_19954,N_19701);
nand UO_828 (O_828,N_19466,N_19691);
nor UO_829 (O_829,N_19901,N_19618);
and UO_830 (O_830,N_19848,N_19904);
or UO_831 (O_831,N_19794,N_19359);
nand UO_832 (O_832,N_19328,N_19683);
nand UO_833 (O_833,N_19137,N_19422);
nand UO_834 (O_834,N_19227,N_19664);
and UO_835 (O_835,N_19653,N_19333);
or UO_836 (O_836,N_19487,N_19392);
xor UO_837 (O_837,N_19329,N_19915);
xnor UO_838 (O_838,N_19034,N_19078);
nand UO_839 (O_839,N_19459,N_19393);
nand UO_840 (O_840,N_19262,N_19852);
and UO_841 (O_841,N_19865,N_19820);
nand UO_842 (O_842,N_19490,N_19176);
or UO_843 (O_843,N_19463,N_19202);
xnor UO_844 (O_844,N_19068,N_19564);
xnor UO_845 (O_845,N_19682,N_19893);
xor UO_846 (O_846,N_19543,N_19726);
and UO_847 (O_847,N_19902,N_19079);
and UO_848 (O_848,N_19013,N_19910);
or UO_849 (O_849,N_19725,N_19722);
or UO_850 (O_850,N_19855,N_19646);
nand UO_851 (O_851,N_19762,N_19232);
and UO_852 (O_852,N_19696,N_19577);
and UO_853 (O_853,N_19137,N_19684);
nor UO_854 (O_854,N_19099,N_19532);
nand UO_855 (O_855,N_19267,N_19853);
or UO_856 (O_856,N_19078,N_19265);
and UO_857 (O_857,N_19492,N_19566);
nor UO_858 (O_858,N_19156,N_19515);
nand UO_859 (O_859,N_19289,N_19389);
nand UO_860 (O_860,N_19227,N_19417);
xor UO_861 (O_861,N_19358,N_19140);
xnor UO_862 (O_862,N_19186,N_19749);
xor UO_863 (O_863,N_19893,N_19100);
nor UO_864 (O_864,N_19330,N_19967);
and UO_865 (O_865,N_19968,N_19983);
and UO_866 (O_866,N_19141,N_19207);
nand UO_867 (O_867,N_19676,N_19743);
nand UO_868 (O_868,N_19598,N_19905);
nor UO_869 (O_869,N_19728,N_19047);
and UO_870 (O_870,N_19350,N_19027);
xnor UO_871 (O_871,N_19789,N_19931);
and UO_872 (O_872,N_19230,N_19327);
nor UO_873 (O_873,N_19278,N_19374);
nor UO_874 (O_874,N_19122,N_19166);
xnor UO_875 (O_875,N_19653,N_19738);
and UO_876 (O_876,N_19600,N_19592);
nor UO_877 (O_877,N_19928,N_19818);
nor UO_878 (O_878,N_19978,N_19298);
or UO_879 (O_879,N_19889,N_19631);
nor UO_880 (O_880,N_19187,N_19410);
and UO_881 (O_881,N_19834,N_19588);
or UO_882 (O_882,N_19598,N_19086);
nor UO_883 (O_883,N_19044,N_19858);
xor UO_884 (O_884,N_19622,N_19438);
nand UO_885 (O_885,N_19346,N_19204);
xor UO_886 (O_886,N_19568,N_19185);
and UO_887 (O_887,N_19213,N_19879);
nand UO_888 (O_888,N_19092,N_19586);
xor UO_889 (O_889,N_19450,N_19608);
nand UO_890 (O_890,N_19074,N_19031);
nand UO_891 (O_891,N_19819,N_19991);
or UO_892 (O_892,N_19067,N_19013);
or UO_893 (O_893,N_19530,N_19024);
nand UO_894 (O_894,N_19266,N_19022);
or UO_895 (O_895,N_19781,N_19521);
nand UO_896 (O_896,N_19749,N_19010);
or UO_897 (O_897,N_19086,N_19402);
nand UO_898 (O_898,N_19643,N_19961);
xnor UO_899 (O_899,N_19878,N_19637);
and UO_900 (O_900,N_19494,N_19470);
nand UO_901 (O_901,N_19166,N_19314);
or UO_902 (O_902,N_19531,N_19850);
xor UO_903 (O_903,N_19037,N_19102);
or UO_904 (O_904,N_19253,N_19016);
and UO_905 (O_905,N_19877,N_19061);
nand UO_906 (O_906,N_19249,N_19336);
nand UO_907 (O_907,N_19847,N_19644);
and UO_908 (O_908,N_19679,N_19696);
nand UO_909 (O_909,N_19534,N_19458);
or UO_910 (O_910,N_19699,N_19344);
xnor UO_911 (O_911,N_19173,N_19558);
xnor UO_912 (O_912,N_19367,N_19411);
and UO_913 (O_913,N_19934,N_19946);
and UO_914 (O_914,N_19466,N_19418);
and UO_915 (O_915,N_19690,N_19778);
and UO_916 (O_916,N_19897,N_19227);
xor UO_917 (O_917,N_19225,N_19298);
nand UO_918 (O_918,N_19402,N_19457);
nand UO_919 (O_919,N_19333,N_19924);
nand UO_920 (O_920,N_19658,N_19447);
or UO_921 (O_921,N_19606,N_19631);
nand UO_922 (O_922,N_19574,N_19773);
or UO_923 (O_923,N_19377,N_19639);
nand UO_924 (O_924,N_19301,N_19376);
and UO_925 (O_925,N_19805,N_19428);
or UO_926 (O_926,N_19976,N_19062);
nor UO_927 (O_927,N_19123,N_19919);
or UO_928 (O_928,N_19789,N_19549);
and UO_929 (O_929,N_19510,N_19562);
and UO_930 (O_930,N_19808,N_19400);
or UO_931 (O_931,N_19565,N_19434);
or UO_932 (O_932,N_19440,N_19067);
or UO_933 (O_933,N_19963,N_19051);
and UO_934 (O_934,N_19338,N_19480);
and UO_935 (O_935,N_19766,N_19545);
nand UO_936 (O_936,N_19579,N_19838);
and UO_937 (O_937,N_19597,N_19528);
or UO_938 (O_938,N_19381,N_19175);
nor UO_939 (O_939,N_19798,N_19500);
nand UO_940 (O_940,N_19174,N_19893);
nand UO_941 (O_941,N_19572,N_19313);
nor UO_942 (O_942,N_19773,N_19097);
or UO_943 (O_943,N_19569,N_19174);
and UO_944 (O_944,N_19156,N_19227);
nand UO_945 (O_945,N_19489,N_19895);
and UO_946 (O_946,N_19506,N_19286);
nor UO_947 (O_947,N_19081,N_19201);
and UO_948 (O_948,N_19380,N_19444);
or UO_949 (O_949,N_19837,N_19812);
or UO_950 (O_950,N_19164,N_19887);
xor UO_951 (O_951,N_19273,N_19929);
nor UO_952 (O_952,N_19152,N_19618);
nand UO_953 (O_953,N_19752,N_19894);
nand UO_954 (O_954,N_19813,N_19963);
xor UO_955 (O_955,N_19488,N_19462);
and UO_956 (O_956,N_19385,N_19874);
and UO_957 (O_957,N_19987,N_19547);
nand UO_958 (O_958,N_19344,N_19873);
xor UO_959 (O_959,N_19832,N_19777);
nor UO_960 (O_960,N_19415,N_19469);
nand UO_961 (O_961,N_19982,N_19067);
or UO_962 (O_962,N_19067,N_19825);
nand UO_963 (O_963,N_19760,N_19180);
xnor UO_964 (O_964,N_19606,N_19275);
nor UO_965 (O_965,N_19657,N_19439);
nand UO_966 (O_966,N_19686,N_19910);
and UO_967 (O_967,N_19539,N_19818);
nor UO_968 (O_968,N_19855,N_19342);
nand UO_969 (O_969,N_19111,N_19599);
or UO_970 (O_970,N_19348,N_19738);
nor UO_971 (O_971,N_19361,N_19504);
nor UO_972 (O_972,N_19368,N_19710);
nor UO_973 (O_973,N_19347,N_19604);
or UO_974 (O_974,N_19906,N_19327);
and UO_975 (O_975,N_19075,N_19474);
nor UO_976 (O_976,N_19109,N_19421);
nor UO_977 (O_977,N_19010,N_19492);
xnor UO_978 (O_978,N_19774,N_19347);
nand UO_979 (O_979,N_19399,N_19880);
xnor UO_980 (O_980,N_19236,N_19632);
and UO_981 (O_981,N_19789,N_19878);
xnor UO_982 (O_982,N_19286,N_19818);
and UO_983 (O_983,N_19241,N_19112);
xor UO_984 (O_984,N_19671,N_19448);
nor UO_985 (O_985,N_19697,N_19988);
or UO_986 (O_986,N_19489,N_19416);
xor UO_987 (O_987,N_19039,N_19479);
nor UO_988 (O_988,N_19253,N_19662);
nor UO_989 (O_989,N_19115,N_19775);
or UO_990 (O_990,N_19409,N_19107);
and UO_991 (O_991,N_19766,N_19534);
nand UO_992 (O_992,N_19320,N_19856);
xnor UO_993 (O_993,N_19695,N_19661);
xnor UO_994 (O_994,N_19021,N_19202);
nand UO_995 (O_995,N_19181,N_19584);
nand UO_996 (O_996,N_19996,N_19260);
nand UO_997 (O_997,N_19406,N_19179);
xnor UO_998 (O_998,N_19004,N_19739);
nand UO_999 (O_999,N_19907,N_19801);
or UO_1000 (O_1000,N_19219,N_19992);
nand UO_1001 (O_1001,N_19183,N_19472);
nor UO_1002 (O_1002,N_19980,N_19865);
and UO_1003 (O_1003,N_19951,N_19849);
and UO_1004 (O_1004,N_19728,N_19552);
nand UO_1005 (O_1005,N_19910,N_19210);
nand UO_1006 (O_1006,N_19045,N_19035);
and UO_1007 (O_1007,N_19284,N_19608);
or UO_1008 (O_1008,N_19080,N_19258);
nor UO_1009 (O_1009,N_19148,N_19129);
xnor UO_1010 (O_1010,N_19331,N_19794);
xnor UO_1011 (O_1011,N_19443,N_19978);
xnor UO_1012 (O_1012,N_19458,N_19666);
nand UO_1013 (O_1013,N_19487,N_19014);
xor UO_1014 (O_1014,N_19100,N_19010);
nor UO_1015 (O_1015,N_19679,N_19722);
nor UO_1016 (O_1016,N_19303,N_19810);
and UO_1017 (O_1017,N_19033,N_19168);
nor UO_1018 (O_1018,N_19334,N_19593);
or UO_1019 (O_1019,N_19303,N_19611);
nor UO_1020 (O_1020,N_19476,N_19917);
xnor UO_1021 (O_1021,N_19427,N_19368);
xor UO_1022 (O_1022,N_19007,N_19733);
xnor UO_1023 (O_1023,N_19326,N_19178);
xnor UO_1024 (O_1024,N_19174,N_19033);
and UO_1025 (O_1025,N_19064,N_19235);
and UO_1026 (O_1026,N_19835,N_19097);
xor UO_1027 (O_1027,N_19757,N_19664);
nor UO_1028 (O_1028,N_19753,N_19723);
nand UO_1029 (O_1029,N_19752,N_19407);
nor UO_1030 (O_1030,N_19266,N_19846);
xnor UO_1031 (O_1031,N_19986,N_19239);
nor UO_1032 (O_1032,N_19274,N_19664);
and UO_1033 (O_1033,N_19787,N_19781);
nor UO_1034 (O_1034,N_19877,N_19265);
nand UO_1035 (O_1035,N_19959,N_19622);
nand UO_1036 (O_1036,N_19306,N_19715);
xor UO_1037 (O_1037,N_19951,N_19622);
or UO_1038 (O_1038,N_19026,N_19516);
xnor UO_1039 (O_1039,N_19204,N_19058);
nor UO_1040 (O_1040,N_19332,N_19881);
or UO_1041 (O_1041,N_19588,N_19785);
nor UO_1042 (O_1042,N_19455,N_19018);
or UO_1043 (O_1043,N_19887,N_19833);
nor UO_1044 (O_1044,N_19240,N_19019);
and UO_1045 (O_1045,N_19440,N_19945);
and UO_1046 (O_1046,N_19735,N_19039);
or UO_1047 (O_1047,N_19547,N_19332);
xnor UO_1048 (O_1048,N_19457,N_19364);
nand UO_1049 (O_1049,N_19394,N_19052);
and UO_1050 (O_1050,N_19880,N_19910);
xnor UO_1051 (O_1051,N_19724,N_19582);
or UO_1052 (O_1052,N_19240,N_19919);
or UO_1053 (O_1053,N_19646,N_19000);
xor UO_1054 (O_1054,N_19646,N_19356);
nand UO_1055 (O_1055,N_19184,N_19732);
and UO_1056 (O_1056,N_19041,N_19219);
nor UO_1057 (O_1057,N_19947,N_19421);
and UO_1058 (O_1058,N_19620,N_19781);
xor UO_1059 (O_1059,N_19177,N_19570);
and UO_1060 (O_1060,N_19175,N_19772);
xor UO_1061 (O_1061,N_19452,N_19140);
nor UO_1062 (O_1062,N_19876,N_19125);
xor UO_1063 (O_1063,N_19864,N_19293);
or UO_1064 (O_1064,N_19804,N_19704);
or UO_1065 (O_1065,N_19302,N_19309);
and UO_1066 (O_1066,N_19608,N_19831);
nor UO_1067 (O_1067,N_19416,N_19202);
or UO_1068 (O_1068,N_19365,N_19301);
or UO_1069 (O_1069,N_19404,N_19689);
and UO_1070 (O_1070,N_19115,N_19273);
or UO_1071 (O_1071,N_19433,N_19575);
nor UO_1072 (O_1072,N_19271,N_19742);
nor UO_1073 (O_1073,N_19146,N_19992);
xor UO_1074 (O_1074,N_19966,N_19531);
or UO_1075 (O_1075,N_19721,N_19130);
nor UO_1076 (O_1076,N_19372,N_19617);
and UO_1077 (O_1077,N_19472,N_19702);
or UO_1078 (O_1078,N_19784,N_19585);
or UO_1079 (O_1079,N_19237,N_19034);
xor UO_1080 (O_1080,N_19585,N_19480);
nand UO_1081 (O_1081,N_19685,N_19364);
nand UO_1082 (O_1082,N_19840,N_19167);
and UO_1083 (O_1083,N_19150,N_19513);
xnor UO_1084 (O_1084,N_19700,N_19946);
xnor UO_1085 (O_1085,N_19398,N_19902);
nand UO_1086 (O_1086,N_19855,N_19258);
or UO_1087 (O_1087,N_19089,N_19610);
or UO_1088 (O_1088,N_19878,N_19573);
xor UO_1089 (O_1089,N_19657,N_19226);
xnor UO_1090 (O_1090,N_19936,N_19170);
or UO_1091 (O_1091,N_19905,N_19168);
xor UO_1092 (O_1092,N_19905,N_19562);
and UO_1093 (O_1093,N_19377,N_19257);
xnor UO_1094 (O_1094,N_19048,N_19635);
xnor UO_1095 (O_1095,N_19558,N_19213);
xor UO_1096 (O_1096,N_19863,N_19190);
and UO_1097 (O_1097,N_19201,N_19068);
nand UO_1098 (O_1098,N_19817,N_19296);
nand UO_1099 (O_1099,N_19779,N_19086);
xnor UO_1100 (O_1100,N_19840,N_19176);
and UO_1101 (O_1101,N_19235,N_19158);
xnor UO_1102 (O_1102,N_19735,N_19616);
xnor UO_1103 (O_1103,N_19495,N_19211);
and UO_1104 (O_1104,N_19643,N_19474);
xnor UO_1105 (O_1105,N_19579,N_19410);
xor UO_1106 (O_1106,N_19452,N_19149);
or UO_1107 (O_1107,N_19679,N_19427);
or UO_1108 (O_1108,N_19078,N_19977);
xnor UO_1109 (O_1109,N_19120,N_19026);
nand UO_1110 (O_1110,N_19843,N_19594);
nor UO_1111 (O_1111,N_19989,N_19099);
nor UO_1112 (O_1112,N_19507,N_19509);
xor UO_1113 (O_1113,N_19632,N_19873);
nor UO_1114 (O_1114,N_19219,N_19897);
nand UO_1115 (O_1115,N_19806,N_19205);
xnor UO_1116 (O_1116,N_19875,N_19456);
nor UO_1117 (O_1117,N_19610,N_19058);
or UO_1118 (O_1118,N_19521,N_19093);
and UO_1119 (O_1119,N_19777,N_19686);
xor UO_1120 (O_1120,N_19526,N_19162);
nand UO_1121 (O_1121,N_19873,N_19943);
nor UO_1122 (O_1122,N_19046,N_19297);
nand UO_1123 (O_1123,N_19093,N_19266);
and UO_1124 (O_1124,N_19480,N_19873);
and UO_1125 (O_1125,N_19612,N_19655);
or UO_1126 (O_1126,N_19818,N_19479);
and UO_1127 (O_1127,N_19401,N_19719);
xnor UO_1128 (O_1128,N_19098,N_19672);
xor UO_1129 (O_1129,N_19381,N_19123);
xnor UO_1130 (O_1130,N_19220,N_19611);
nor UO_1131 (O_1131,N_19188,N_19690);
xnor UO_1132 (O_1132,N_19294,N_19638);
nand UO_1133 (O_1133,N_19549,N_19121);
or UO_1134 (O_1134,N_19792,N_19515);
nor UO_1135 (O_1135,N_19694,N_19302);
xnor UO_1136 (O_1136,N_19806,N_19138);
nand UO_1137 (O_1137,N_19310,N_19356);
and UO_1138 (O_1138,N_19229,N_19013);
nand UO_1139 (O_1139,N_19345,N_19047);
and UO_1140 (O_1140,N_19239,N_19416);
and UO_1141 (O_1141,N_19745,N_19057);
xnor UO_1142 (O_1142,N_19619,N_19187);
and UO_1143 (O_1143,N_19111,N_19626);
nand UO_1144 (O_1144,N_19330,N_19338);
nor UO_1145 (O_1145,N_19576,N_19198);
and UO_1146 (O_1146,N_19701,N_19580);
nand UO_1147 (O_1147,N_19892,N_19282);
and UO_1148 (O_1148,N_19657,N_19842);
nand UO_1149 (O_1149,N_19533,N_19833);
and UO_1150 (O_1150,N_19589,N_19685);
and UO_1151 (O_1151,N_19082,N_19789);
nand UO_1152 (O_1152,N_19448,N_19242);
nand UO_1153 (O_1153,N_19911,N_19500);
and UO_1154 (O_1154,N_19688,N_19970);
xor UO_1155 (O_1155,N_19195,N_19876);
and UO_1156 (O_1156,N_19116,N_19460);
and UO_1157 (O_1157,N_19058,N_19618);
nor UO_1158 (O_1158,N_19389,N_19547);
nor UO_1159 (O_1159,N_19570,N_19967);
or UO_1160 (O_1160,N_19793,N_19304);
and UO_1161 (O_1161,N_19092,N_19634);
and UO_1162 (O_1162,N_19729,N_19950);
or UO_1163 (O_1163,N_19710,N_19821);
nand UO_1164 (O_1164,N_19097,N_19900);
or UO_1165 (O_1165,N_19608,N_19268);
and UO_1166 (O_1166,N_19453,N_19062);
or UO_1167 (O_1167,N_19239,N_19523);
nand UO_1168 (O_1168,N_19478,N_19620);
nor UO_1169 (O_1169,N_19834,N_19927);
and UO_1170 (O_1170,N_19951,N_19080);
and UO_1171 (O_1171,N_19142,N_19175);
xnor UO_1172 (O_1172,N_19153,N_19466);
or UO_1173 (O_1173,N_19257,N_19721);
nor UO_1174 (O_1174,N_19816,N_19127);
and UO_1175 (O_1175,N_19329,N_19975);
nand UO_1176 (O_1176,N_19526,N_19896);
and UO_1177 (O_1177,N_19176,N_19757);
xor UO_1178 (O_1178,N_19580,N_19542);
xor UO_1179 (O_1179,N_19682,N_19333);
xnor UO_1180 (O_1180,N_19862,N_19877);
xor UO_1181 (O_1181,N_19467,N_19782);
nand UO_1182 (O_1182,N_19684,N_19129);
nor UO_1183 (O_1183,N_19558,N_19938);
nand UO_1184 (O_1184,N_19052,N_19605);
nor UO_1185 (O_1185,N_19705,N_19276);
xor UO_1186 (O_1186,N_19148,N_19265);
nand UO_1187 (O_1187,N_19447,N_19000);
nor UO_1188 (O_1188,N_19358,N_19165);
xnor UO_1189 (O_1189,N_19559,N_19521);
nor UO_1190 (O_1190,N_19370,N_19102);
and UO_1191 (O_1191,N_19521,N_19089);
xnor UO_1192 (O_1192,N_19951,N_19458);
and UO_1193 (O_1193,N_19417,N_19859);
nor UO_1194 (O_1194,N_19854,N_19443);
xnor UO_1195 (O_1195,N_19490,N_19063);
nor UO_1196 (O_1196,N_19389,N_19831);
or UO_1197 (O_1197,N_19257,N_19962);
and UO_1198 (O_1198,N_19678,N_19828);
xor UO_1199 (O_1199,N_19295,N_19409);
xnor UO_1200 (O_1200,N_19961,N_19218);
and UO_1201 (O_1201,N_19300,N_19963);
nor UO_1202 (O_1202,N_19590,N_19531);
and UO_1203 (O_1203,N_19581,N_19925);
nor UO_1204 (O_1204,N_19122,N_19261);
nand UO_1205 (O_1205,N_19346,N_19557);
and UO_1206 (O_1206,N_19093,N_19752);
nor UO_1207 (O_1207,N_19860,N_19148);
or UO_1208 (O_1208,N_19740,N_19457);
and UO_1209 (O_1209,N_19511,N_19315);
or UO_1210 (O_1210,N_19685,N_19601);
and UO_1211 (O_1211,N_19876,N_19621);
xnor UO_1212 (O_1212,N_19216,N_19431);
nor UO_1213 (O_1213,N_19751,N_19153);
or UO_1214 (O_1214,N_19427,N_19909);
or UO_1215 (O_1215,N_19832,N_19013);
nand UO_1216 (O_1216,N_19143,N_19309);
nand UO_1217 (O_1217,N_19648,N_19435);
xnor UO_1218 (O_1218,N_19322,N_19104);
nand UO_1219 (O_1219,N_19365,N_19642);
nand UO_1220 (O_1220,N_19315,N_19445);
nand UO_1221 (O_1221,N_19961,N_19913);
nand UO_1222 (O_1222,N_19769,N_19225);
and UO_1223 (O_1223,N_19133,N_19453);
and UO_1224 (O_1224,N_19840,N_19796);
and UO_1225 (O_1225,N_19679,N_19438);
nor UO_1226 (O_1226,N_19488,N_19337);
or UO_1227 (O_1227,N_19655,N_19197);
and UO_1228 (O_1228,N_19555,N_19742);
nand UO_1229 (O_1229,N_19228,N_19039);
nor UO_1230 (O_1230,N_19842,N_19667);
xnor UO_1231 (O_1231,N_19763,N_19036);
or UO_1232 (O_1232,N_19150,N_19116);
nor UO_1233 (O_1233,N_19127,N_19873);
or UO_1234 (O_1234,N_19638,N_19009);
and UO_1235 (O_1235,N_19715,N_19885);
nand UO_1236 (O_1236,N_19293,N_19857);
xor UO_1237 (O_1237,N_19207,N_19016);
or UO_1238 (O_1238,N_19636,N_19056);
nor UO_1239 (O_1239,N_19738,N_19584);
and UO_1240 (O_1240,N_19329,N_19642);
nand UO_1241 (O_1241,N_19890,N_19734);
or UO_1242 (O_1242,N_19860,N_19881);
xor UO_1243 (O_1243,N_19243,N_19870);
nor UO_1244 (O_1244,N_19566,N_19510);
xnor UO_1245 (O_1245,N_19524,N_19460);
xor UO_1246 (O_1246,N_19811,N_19316);
xnor UO_1247 (O_1247,N_19404,N_19430);
and UO_1248 (O_1248,N_19389,N_19599);
nor UO_1249 (O_1249,N_19338,N_19062);
and UO_1250 (O_1250,N_19657,N_19043);
nand UO_1251 (O_1251,N_19305,N_19733);
nor UO_1252 (O_1252,N_19271,N_19568);
nand UO_1253 (O_1253,N_19800,N_19721);
xor UO_1254 (O_1254,N_19135,N_19360);
or UO_1255 (O_1255,N_19295,N_19067);
nand UO_1256 (O_1256,N_19300,N_19341);
nand UO_1257 (O_1257,N_19721,N_19873);
xor UO_1258 (O_1258,N_19074,N_19009);
or UO_1259 (O_1259,N_19855,N_19586);
nand UO_1260 (O_1260,N_19525,N_19332);
xor UO_1261 (O_1261,N_19271,N_19809);
or UO_1262 (O_1262,N_19370,N_19426);
xor UO_1263 (O_1263,N_19262,N_19300);
and UO_1264 (O_1264,N_19415,N_19127);
or UO_1265 (O_1265,N_19577,N_19127);
or UO_1266 (O_1266,N_19616,N_19109);
xor UO_1267 (O_1267,N_19792,N_19701);
nand UO_1268 (O_1268,N_19049,N_19320);
nand UO_1269 (O_1269,N_19637,N_19391);
and UO_1270 (O_1270,N_19439,N_19675);
or UO_1271 (O_1271,N_19230,N_19493);
nand UO_1272 (O_1272,N_19344,N_19717);
nor UO_1273 (O_1273,N_19801,N_19989);
and UO_1274 (O_1274,N_19199,N_19819);
and UO_1275 (O_1275,N_19112,N_19218);
xnor UO_1276 (O_1276,N_19650,N_19336);
nor UO_1277 (O_1277,N_19453,N_19091);
or UO_1278 (O_1278,N_19336,N_19192);
nor UO_1279 (O_1279,N_19934,N_19211);
or UO_1280 (O_1280,N_19572,N_19846);
xnor UO_1281 (O_1281,N_19695,N_19474);
nand UO_1282 (O_1282,N_19000,N_19385);
nor UO_1283 (O_1283,N_19590,N_19414);
nand UO_1284 (O_1284,N_19262,N_19651);
xnor UO_1285 (O_1285,N_19223,N_19705);
or UO_1286 (O_1286,N_19597,N_19414);
and UO_1287 (O_1287,N_19398,N_19628);
or UO_1288 (O_1288,N_19580,N_19743);
nand UO_1289 (O_1289,N_19706,N_19745);
xnor UO_1290 (O_1290,N_19928,N_19601);
nor UO_1291 (O_1291,N_19105,N_19772);
nor UO_1292 (O_1292,N_19264,N_19288);
or UO_1293 (O_1293,N_19656,N_19893);
nor UO_1294 (O_1294,N_19532,N_19602);
nand UO_1295 (O_1295,N_19525,N_19386);
and UO_1296 (O_1296,N_19113,N_19088);
or UO_1297 (O_1297,N_19187,N_19532);
or UO_1298 (O_1298,N_19780,N_19118);
or UO_1299 (O_1299,N_19877,N_19523);
or UO_1300 (O_1300,N_19667,N_19000);
nand UO_1301 (O_1301,N_19593,N_19523);
or UO_1302 (O_1302,N_19177,N_19768);
nand UO_1303 (O_1303,N_19289,N_19243);
nand UO_1304 (O_1304,N_19249,N_19023);
or UO_1305 (O_1305,N_19537,N_19888);
nand UO_1306 (O_1306,N_19812,N_19814);
and UO_1307 (O_1307,N_19175,N_19490);
or UO_1308 (O_1308,N_19239,N_19841);
and UO_1309 (O_1309,N_19048,N_19362);
or UO_1310 (O_1310,N_19043,N_19863);
xor UO_1311 (O_1311,N_19831,N_19330);
and UO_1312 (O_1312,N_19977,N_19782);
nand UO_1313 (O_1313,N_19124,N_19611);
xor UO_1314 (O_1314,N_19668,N_19479);
and UO_1315 (O_1315,N_19426,N_19586);
or UO_1316 (O_1316,N_19754,N_19551);
xnor UO_1317 (O_1317,N_19955,N_19022);
or UO_1318 (O_1318,N_19374,N_19325);
nand UO_1319 (O_1319,N_19426,N_19237);
and UO_1320 (O_1320,N_19999,N_19312);
or UO_1321 (O_1321,N_19345,N_19601);
nor UO_1322 (O_1322,N_19121,N_19342);
or UO_1323 (O_1323,N_19337,N_19519);
nor UO_1324 (O_1324,N_19473,N_19506);
and UO_1325 (O_1325,N_19957,N_19584);
xnor UO_1326 (O_1326,N_19816,N_19669);
nand UO_1327 (O_1327,N_19340,N_19229);
or UO_1328 (O_1328,N_19973,N_19050);
or UO_1329 (O_1329,N_19576,N_19245);
nor UO_1330 (O_1330,N_19169,N_19322);
and UO_1331 (O_1331,N_19026,N_19644);
and UO_1332 (O_1332,N_19039,N_19355);
xor UO_1333 (O_1333,N_19521,N_19334);
nor UO_1334 (O_1334,N_19342,N_19998);
nor UO_1335 (O_1335,N_19867,N_19205);
or UO_1336 (O_1336,N_19815,N_19876);
and UO_1337 (O_1337,N_19559,N_19383);
or UO_1338 (O_1338,N_19638,N_19763);
xor UO_1339 (O_1339,N_19294,N_19004);
nor UO_1340 (O_1340,N_19731,N_19829);
and UO_1341 (O_1341,N_19913,N_19099);
and UO_1342 (O_1342,N_19464,N_19154);
and UO_1343 (O_1343,N_19373,N_19995);
xor UO_1344 (O_1344,N_19548,N_19966);
and UO_1345 (O_1345,N_19551,N_19529);
or UO_1346 (O_1346,N_19172,N_19990);
and UO_1347 (O_1347,N_19138,N_19202);
nand UO_1348 (O_1348,N_19377,N_19193);
nor UO_1349 (O_1349,N_19003,N_19429);
or UO_1350 (O_1350,N_19726,N_19738);
nor UO_1351 (O_1351,N_19498,N_19623);
xnor UO_1352 (O_1352,N_19498,N_19576);
or UO_1353 (O_1353,N_19435,N_19957);
and UO_1354 (O_1354,N_19147,N_19237);
nand UO_1355 (O_1355,N_19542,N_19050);
xor UO_1356 (O_1356,N_19161,N_19451);
and UO_1357 (O_1357,N_19758,N_19487);
and UO_1358 (O_1358,N_19609,N_19320);
xor UO_1359 (O_1359,N_19866,N_19933);
nor UO_1360 (O_1360,N_19708,N_19864);
or UO_1361 (O_1361,N_19663,N_19935);
or UO_1362 (O_1362,N_19843,N_19392);
or UO_1363 (O_1363,N_19347,N_19522);
xor UO_1364 (O_1364,N_19377,N_19153);
nor UO_1365 (O_1365,N_19436,N_19938);
nand UO_1366 (O_1366,N_19788,N_19503);
or UO_1367 (O_1367,N_19540,N_19011);
nor UO_1368 (O_1368,N_19793,N_19101);
nor UO_1369 (O_1369,N_19739,N_19534);
xor UO_1370 (O_1370,N_19094,N_19976);
xnor UO_1371 (O_1371,N_19885,N_19232);
nand UO_1372 (O_1372,N_19696,N_19012);
nand UO_1373 (O_1373,N_19512,N_19117);
and UO_1374 (O_1374,N_19552,N_19687);
or UO_1375 (O_1375,N_19816,N_19203);
nor UO_1376 (O_1376,N_19603,N_19897);
nand UO_1377 (O_1377,N_19135,N_19861);
nor UO_1378 (O_1378,N_19147,N_19256);
or UO_1379 (O_1379,N_19987,N_19659);
or UO_1380 (O_1380,N_19638,N_19126);
xnor UO_1381 (O_1381,N_19080,N_19943);
nor UO_1382 (O_1382,N_19843,N_19950);
nand UO_1383 (O_1383,N_19279,N_19945);
nor UO_1384 (O_1384,N_19008,N_19723);
or UO_1385 (O_1385,N_19684,N_19737);
nor UO_1386 (O_1386,N_19321,N_19479);
nor UO_1387 (O_1387,N_19837,N_19081);
and UO_1388 (O_1388,N_19811,N_19483);
or UO_1389 (O_1389,N_19090,N_19308);
nor UO_1390 (O_1390,N_19150,N_19205);
nor UO_1391 (O_1391,N_19525,N_19865);
xnor UO_1392 (O_1392,N_19956,N_19880);
nor UO_1393 (O_1393,N_19939,N_19819);
or UO_1394 (O_1394,N_19112,N_19588);
xnor UO_1395 (O_1395,N_19421,N_19932);
xnor UO_1396 (O_1396,N_19552,N_19339);
or UO_1397 (O_1397,N_19286,N_19456);
nor UO_1398 (O_1398,N_19113,N_19320);
and UO_1399 (O_1399,N_19389,N_19820);
nor UO_1400 (O_1400,N_19910,N_19034);
nor UO_1401 (O_1401,N_19671,N_19581);
and UO_1402 (O_1402,N_19157,N_19353);
and UO_1403 (O_1403,N_19334,N_19126);
xor UO_1404 (O_1404,N_19156,N_19543);
nand UO_1405 (O_1405,N_19628,N_19890);
and UO_1406 (O_1406,N_19829,N_19318);
xnor UO_1407 (O_1407,N_19931,N_19898);
xnor UO_1408 (O_1408,N_19736,N_19097);
xor UO_1409 (O_1409,N_19955,N_19520);
or UO_1410 (O_1410,N_19279,N_19404);
xnor UO_1411 (O_1411,N_19388,N_19848);
nor UO_1412 (O_1412,N_19879,N_19948);
nor UO_1413 (O_1413,N_19050,N_19659);
nor UO_1414 (O_1414,N_19762,N_19507);
or UO_1415 (O_1415,N_19518,N_19988);
or UO_1416 (O_1416,N_19147,N_19196);
xor UO_1417 (O_1417,N_19209,N_19465);
or UO_1418 (O_1418,N_19974,N_19191);
and UO_1419 (O_1419,N_19251,N_19617);
nor UO_1420 (O_1420,N_19772,N_19874);
nand UO_1421 (O_1421,N_19792,N_19744);
and UO_1422 (O_1422,N_19338,N_19644);
nand UO_1423 (O_1423,N_19517,N_19841);
xnor UO_1424 (O_1424,N_19157,N_19219);
or UO_1425 (O_1425,N_19731,N_19101);
nor UO_1426 (O_1426,N_19049,N_19006);
nand UO_1427 (O_1427,N_19784,N_19778);
nand UO_1428 (O_1428,N_19797,N_19550);
nor UO_1429 (O_1429,N_19097,N_19869);
xnor UO_1430 (O_1430,N_19145,N_19031);
nor UO_1431 (O_1431,N_19907,N_19212);
nand UO_1432 (O_1432,N_19159,N_19219);
nand UO_1433 (O_1433,N_19233,N_19905);
xor UO_1434 (O_1434,N_19408,N_19140);
or UO_1435 (O_1435,N_19240,N_19738);
or UO_1436 (O_1436,N_19502,N_19710);
and UO_1437 (O_1437,N_19857,N_19621);
nand UO_1438 (O_1438,N_19826,N_19452);
nand UO_1439 (O_1439,N_19381,N_19344);
xor UO_1440 (O_1440,N_19993,N_19344);
xnor UO_1441 (O_1441,N_19946,N_19158);
nand UO_1442 (O_1442,N_19220,N_19487);
nor UO_1443 (O_1443,N_19127,N_19779);
and UO_1444 (O_1444,N_19919,N_19929);
nand UO_1445 (O_1445,N_19249,N_19823);
nand UO_1446 (O_1446,N_19687,N_19737);
or UO_1447 (O_1447,N_19429,N_19426);
xnor UO_1448 (O_1448,N_19929,N_19870);
nor UO_1449 (O_1449,N_19105,N_19390);
nand UO_1450 (O_1450,N_19091,N_19233);
and UO_1451 (O_1451,N_19670,N_19952);
nor UO_1452 (O_1452,N_19170,N_19062);
xnor UO_1453 (O_1453,N_19484,N_19754);
nor UO_1454 (O_1454,N_19484,N_19315);
and UO_1455 (O_1455,N_19088,N_19844);
and UO_1456 (O_1456,N_19730,N_19843);
or UO_1457 (O_1457,N_19204,N_19104);
or UO_1458 (O_1458,N_19509,N_19323);
or UO_1459 (O_1459,N_19187,N_19275);
nand UO_1460 (O_1460,N_19597,N_19789);
xor UO_1461 (O_1461,N_19726,N_19595);
xnor UO_1462 (O_1462,N_19720,N_19265);
nor UO_1463 (O_1463,N_19786,N_19015);
xor UO_1464 (O_1464,N_19709,N_19961);
and UO_1465 (O_1465,N_19000,N_19868);
nand UO_1466 (O_1466,N_19705,N_19953);
nor UO_1467 (O_1467,N_19575,N_19078);
nor UO_1468 (O_1468,N_19728,N_19665);
or UO_1469 (O_1469,N_19608,N_19220);
and UO_1470 (O_1470,N_19202,N_19333);
or UO_1471 (O_1471,N_19639,N_19283);
and UO_1472 (O_1472,N_19463,N_19112);
or UO_1473 (O_1473,N_19865,N_19940);
nor UO_1474 (O_1474,N_19955,N_19756);
nand UO_1475 (O_1475,N_19713,N_19227);
or UO_1476 (O_1476,N_19400,N_19902);
xnor UO_1477 (O_1477,N_19245,N_19749);
or UO_1478 (O_1478,N_19011,N_19846);
or UO_1479 (O_1479,N_19615,N_19130);
and UO_1480 (O_1480,N_19920,N_19267);
xor UO_1481 (O_1481,N_19633,N_19691);
nand UO_1482 (O_1482,N_19462,N_19727);
and UO_1483 (O_1483,N_19497,N_19950);
or UO_1484 (O_1484,N_19243,N_19876);
nor UO_1485 (O_1485,N_19463,N_19796);
xor UO_1486 (O_1486,N_19596,N_19759);
nand UO_1487 (O_1487,N_19656,N_19062);
xor UO_1488 (O_1488,N_19404,N_19446);
nand UO_1489 (O_1489,N_19526,N_19571);
nor UO_1490 (O_1490,N_19315,N_19828);
and UO_1491 (O_1491,N_19897,N_19383);
xnor UO_1492 (O_1492,N_19283,N_19584);
nand UO_1493 (O_1493,N_19698,N_19010);
nor UO_1494 (O_1494,N_19830,N_19614);
xnor UO_1495 (O_1495,N_19307,N_19290);
or UO_1496 (O_1496,N_19722,N_19931);
and UO_1497 (O_1497,N_19665,N_19486);
nand UO_1498 (O_1498,N_19202,N_19786);
xnor UO_1499 (O_1499,N_19658,N_19912);
nor UO_1500 (O_1500,N_19273,N_19116);
xnor UO_1501 (O_1501,N_19344,N_19611);
and UO_1502 (O_1502,N_19184,N_19007);
nor UO_1503 (O_1503,N_19736,N_19820);
and UO_1504 (O_1504,N_19579,N_19675);
and UO_1505 (O_1505,N_19801,N_19064);
or UO_1506 (O_1506,N_19139,N_19890);
or UO_1507 (O_1507,N_19245,N_19442);
nand UO_1508 (O_1508,N_19372,N_19375);
nor UO_1509 (O_1509,N_19927,N_19820);
xnor UO_1510 (O_1510,N_19158,N_19187);
or UO_1511 (O_1511,N_19783,N_19582);
and UO_1512 (O_1512,N_19708,N_19489);
xor UO_1513 (O_1513,N_19954,N_19747);
or UO_1514 (O_1514,N_19355,N_19172);
and UO_1515 (O_1515,N_19456,N_19398);
nand UO_1516 (O_1516,N_19115,N_19358);
nand UO_1517 (O_1517,N_19195,N_19514);
nor UO_1518 (O_1518,N_19836,N_19954);
nor UO_1519 (O_1519,N_19718,N_19459);
nor UO_1520 (O_1520,N_19038,N_19640);
nor UO_1521 (O_1521,N_19013,N_19925);
nand UO_1522 (O_1522,N_19750,N_19051);
xor UO_1523 (O_1523,N_19797,N_19917);
and UO_1524 (O_1524,N_19999,N_19252);
xnor UO_1525 (O_1525,N_19120,N_19004);
nand UO_1526 (O_1526,N_19530,N_19480);
nor UO_1527 (O_1527,N_19672,N_19807);
or UO_1528 (O_1528,N_19009,N_19022);
and UO_1529 (O_1529,N_19338,N_19746);
or UO_1530 (O_1530,N_19525,N_19885);
xor UO_1531 (O_1531,N_19540,N_19071);
nand UO_1532 (O_1532,N_19063,N_19701);
xnor UO_1533 (O_1533,N_19695,N_19126);
xnor UO_1534 (O_1534,N_19858,N_19113);
nor UO_1535 (O_1535,N_19819,N_19844);
and UO_1536 (O_1536,N_19587,N_19766);
nor UO_1537 (O_1537,N_19237,N_19071);
nand UO_1538 (O_1538,N_19409,N_19369);
nand UO_1539 (O_1539,N_19375,N_19190);
xor UO_1540 (O_1540,N_19162,N_19488);
nand UO_1541 (O_1541,N_19525,N_19812);
xor UO_1542 (O_1542,N_19326,N_19006);
and UO_1543 (O_1543,N_19429,N_19700);
xnor UO_1544 (O_1544,N_19425,N_19905);
and UO_1545 (O_1545,N_19447,N_19084);
nand UO_1546 (O_1546,N_19223,N_19520);
or UO_1547 (O_1547,N_19353,N_19418);
nand UO_1548 (O_1548,N_19530,N_19690);
xnor UO_1549 (O_1549,N_19614,N_19493);
or UO_1550 (O_1550,N_19335,N_19556);
nor UO_1551 (O_1551,N_19231,N_19406);
or UO_1552 (O_1552,N_19120,N_19560);
nand UO_1553 (O_1553,N_19123,N_19270);
nand UO_1554 (O_1554,N_19600,N_19697);
and UO_1555 (O_1555,N_19038,N_19525);
or UO_1556 (O_1556,N_19982,N_19641);
or UO_1557 (O_1557,N_19819,N_19250);
and UO_1558 (O_1558,N_19609,N_19453);
nor UO_1559 (O_1559,N_19713,N_19459);
nor UO_1560 (O_1560,N_19203,N_19417);
nand UO_1561 (O_1561,N_19095,N_19211);
and UO_1562 (O_1562,N_19052,N_19643);
and UO_1563 (O_1563,N_19528,N_19861);
xor UO_1564 (O_1564,N_19408,N_19721);
and UO_1565 (O_1565,N_19692,N_19426);
nand UO_1566 (O_1566,N_19093,N_19789);
xor UO_1567 (O_1567,N_19941,N_19178);
and UO_1568 (O_1568,N_19374,N_19238);
nor UO_1569 (O_1569,N_19933,N_19472);
and UO_1570 (O_1570,N_19687,N_19484);
xnor UO_1571 (O_1571,N_19261,N_19751);
or UO_1572 (O_1572,N_19553,N_19046);
and UO_1573 (O_1573,N_19784,N_19677);
or UO_1574 (O_1574,N_19678,N_19890);
nand UO_1575 (O_1575,N_19065,N_19842);
nor UO_1576 (O_1576,N_19176,N_19454);
xor UO_1577 (O_1577,N_19153,N_19187);
nor UO_1578 (O_1578,N_19827,N_19205);
nand UO_1579 (O_1579,N_19434,N_19693);
xor UO_1580 (O_1580,N_19239,N_19068);
and UO_1581 (O_1581,N_19561,N_19110);
xor UO_1582 (O_1582,N_19281,N_19955);
nor UO_1583 (O_1583,N_19884,N_19188);
or UO_1584 (O_1584,N_19943,N_19775);
and UO_1585 (O_1585,N_19216,N_19494);
xnor UO_1586 (O_1586,N_19998,N_19757);
nand UO_1587 (O_1587,N_19841,N_19442);
nor UO_1588 (O_1588,N_19294,N_19026);
and UO_1589 (O_1589,N_19523,N_19857);
xor UO_1590 (O_1590,N_19044,N_19060);
or UO_1591 (O_1591,N_19216,N_19702);
nor UO_1592 (O_1592,N_19589,N_19661);
xor UO_1593 (O_1593,N_19968,N_19180);
nand UO_1594 (O_1594,N_19396,N_19458);
and UO_1595 (O_1595,N_19308,N_19390);
nor UO_1596 (O_1596,N_19154,N_19928);
xor UO_1597 (O_1597,N_19546,N_19933);
xor UO_1598 (O_1598,N_19284,N_19585);
nor UO_1599 (O_1599,N_19344,N_19044);
and UO_1600 (O_1600,N_19044,N_19546);
and UO_1601 (O_1601,N_19677,N_19949);
nor UO_1602 (O_1602,N_19961,N_19502);
nor UO_1603 (O_1603,N_19366,N_19600);
xnor UO_1604 (O_1604,N_19867,N_19339);
or UO_1605 (O_1605,N_19318,N_19878);
xor UO_1606 (O_1606,N_19345,N_19638);
nor UO_1607 (O_1607,N_19599,N_19152);
xnor UO_1608 (O_1608,N_19551,N_19153);
nand UO_1609 (O_1609,N_19664,N_19422);
nor UO_1610 (O_1610,N_19079,N_19035);
and UO_1611 (O_1611,N_19908,N_19482);
nor UO_1612 (O_1612,N_19966,N_19206);
nand UO_1613 (O_1613,N_19153,N_19053);
xnor UO_1614 (O_1614,N_19848,N_19508);
and UO_1615 (O_1615,N_19084,N_19590);
nand UO_1616 (O_1616,N_19598,N_19423);
nand UO_1617 (O_1617,N_19508,N_19024);
xnor UO_1618 (O_1618,N_19772,N_19151);
xnor UO_1619 (O_1619,N_19484,N_19291);
nand UO_1620 (O_1620,N_19937,N_19439);
or UO_1621 (O_1621,N_19757,N_19064);
nor UO_1622 (O_1622,N_19311,N_19014);
nand UO_1623 (O_1623,N_19950,N_19773);
xor UO_1624 (O_1624,N_19001,N_19360);
xnor UO_1625 (O_1625,N_19033,N_19954);
nand UO_1626 (O_1626,N_19267,N_19086);
nor UO_1627 (O_1627,N_19150,N_19948);
or UO_1628 (O_1628,N_19155,N_19809);
nor UO_1629 (O_1629,N_19995,N_19638);
nand UO_1630 (O_1630,N_19335,N_19099);
and UO_1631 (O_1631,N_19626,N_19011);
xnor UO_1632 (O_1632,N_19323,N_19881);
nor UO_1633 (O_1633,N_19237,N_19251);
xnor UO_1634 (O_1634,N_19877,N_19690);
xnor UO_1635 (O_1635,N_19993,N_19740);
xor UO_1636 (O_1636,N_19153,N_19098);
and UO_1637 (O_1637,N_19975,N_19356);
or UO_1638 (O_1638,N_19349,N_19407);
nand UO_1639 (O_1639,N_19324,N_19899);
xnor UO_1640 (O_1640,N_19472,N_19002);
xor UO_1641 (O_1641,N_19764,N_19087);
nor UO_1642 (O_1642,N_19696,N_19252);
xnor UO_1643 (O_1643,N_19322,N_19555);
and UO_1644 (O_1644,N_19492,N_19877);
or UO_1645 (O_1645,N_19598,N_19728);
or UO_1646 (O_1646,N_19866,N_19687);
xnor UO_1647 (O_1647,N_19196,N_19433);
and UO_1648 (O_1648,N_19497,N_19873);
and UO_1649 (O_1649,N_19514,N_19220);
nand UO_1650 (O_1650,N_19308,N_19150);
nand UO_1651 (O_1651,N_19350,N_19975);
nand UO_1652 (O_1652,N_19937,N_19824);
nor UO_1653 (O_1653,N_19989,N_19541);
xnor UO_1654 (O_1654,N_19128,N_19762);
or UO_1655 (O_1655,N_19461,N_19171);
nor UO_1656 (O_1656,N_19155,N_19646);
nand UO_1657 (O_1657,N_19054,N_19026);
or UO_1658 (O_1658,N_19635,N_19352);
and UO_1659 (O_1659,N_19519,N_19774);
and UO_1660 (O_1660,N_19630,N_19306);
or UO_1661 (O_1661,N_19616,N_19684);
xnor UO_1662 (O_1662,N_19549,N_19396);
or UO_1663 (O_1663,N_19322,N_19308);
nor UO_1664 (O_1664,N_19319,N_19004);
and UO_1665 (O_1665,N_19473,N_19574);
and UO_1666 (O_1666,N_19191,N_19786);
and UO_1667 (O_1667,N_19641,N_19459);
or UO_1668 (O_1668,N_19758,N_19451);
or UO_1669 (O_1669,N_19669,N_19922);
and UO_1670 (O_1670,N_19458,N_19087);
xnor UO_1671 (O_1671,N_19539,N_19167);
xor UO_1672 (O_1672,N_19135,N_19173);
and UO_1673 (O_1673,N_19888,N_19915);
and UO_1674 (O_1674,N_19554,N_19812);
nand UO_1675 (O_1675,N_19284,N_19458);
nor UO_1676 (O_1676,N_19736,N_19805);
xor UO_1677 (O_1677,N_19331,N_19691);
or UO_1678 (O_1678,N_19528,N_19236);
nor UO_1679 (O_1679,N_19280,N_19151);
xnor UO_1680 (O_1680,N_19583,N_19725);
and UO_1681 (O_1681,N_19851,N_19997);
nand UO_1682 (O_1682,N_19431,N_19676);
and UO_1683 (O_1683,N_19570,N_19249);
nor UO_1684 (O_1684,N_19225,N_19356);
nor UO_1685 (O_1685,N_19260,N_19731);
xnor UO_1686 (O_1686,N_19681,N_19741);
and UO_1687 (O_1687,N_19907,N_19254);
or UO_1688 (O_1688,N_19544,N_19542);
or UO_1689 (O_1689,N_19783,N_19677);
or UO_1690 (O_1690,N_19923,N_19833);
nor UO_1691 (O_1691,N_19744,N_19321);
or UO_1692 (O_1692,N_19927,N_19308);
nand UO_1693 (O_1693,N_19248,N_19401);
or UO_1694 (O_1694,N_19003,N_19835);
nand UO_1695 (O_1695,N_19500,N_19438);
nor UO_1696 (O_1696,N_19259,N_19794);
nor UO_1697 (O_1697,N_19287,N_19020);
or UO_1698 (O_1698,N_19170,N_19336);
or UO_1699 (O_1699,N_19760,N_19861);
and UO_1700 (O_1700,N_19444,N_19611);
nand UO_1701 (O_1701,N_19323,N_19755);
nand UO_1702 (O_1702,N_19576,N_19614);
nor UO_1703 (O_1703,N_19668,N_19991);
nand UO_1704 (O_1704,N_19010,N_19895);
or UO_1705 (O_1705,N_19459,N_19136);
xnor UO_1706 (O_1706,N_19322,N_19800);
xnor UO_1707 (O_1707,N_19295,N_19170);
nand UO_1708 (O_1708,N_19138,N_19503);
nand UO_1709 (O_1709,N_19489,N_19798);
xnor UO_1710 (O_1710,N_19966,N_19181);
or UO_1711 (O_1711,N_19656,N_19626);
nor UO_1712 (O_1712,N_19422,N_19883);
or UO_1713 (O_1713,N_19563,N_19301);
xor UO_1714 (O_1714,N_19597,N_19102);
nor UO_1715 (O_1715,N_19814,N_19417);
nor UO_1716 (O_1716,N_19886,N_19665);
and UO_1717 (O_1717,N_19225,N_19574);
xor UO_1718 (O_1718,N_19504,N_19511);
nand UO_1719 (O_1719,N_19400,N_19923);
or UO_1720 (O_1720,N_19197,N_19444);
nand UO_1721 (O_1721,N_19899,N_19209);
nor UO_1722 (O_1722,N_19708,N_19320);
or UO_1723 (O_1723,N_19855,N_19606);
nor UO_1724 (O_1724,N_19045,N_19518);
nand UO_1725 (O_1725,N_19262,N_19705);
xor UO_1726 (O_1726,N_19007,N_19550);
nor UO_1727 (O_1727,N_19387,N_19625);
nor UO_1728 (O_1728,N_19814,N_19317);
xnor UO_1729 (O_1729,N_19521,N_19671);
nand UO_1730 (O_1730,N_19902,N_19275);
xnor UO_1731 (O_1731,N_19933,N_19079);
nor UO_1732 (O_1732,N_19898,N_19194);
nor UO_1733 (O_1733,N_19630,N_19557);
and UO_1734 (O_1734,N_19674,N_19791);
nand UO_1735 (O_1735,N_19727,N_19910);
nor UO_1736 (O_1736,N_19236,N_19405);
and UO_1737 (O_1737,N_19939,N_19947);
or UO_1738 (O_1738,N_19006,N_19766);
or UO_1739 (O_1739,N_19686,N_19391);
nand UO_1740 (O_1740,N_19107,N_19774);
xor UO_1741 (O_1741,N_19612,N_19669);
and UO_1742 (O_1742,N_19724,N_19141);
nand UO_1743 (O_1743,N_19261,N_19267);
and UO_1744 (O_1744,N_19059,N_19656);
and UO_1745 (O_1745,N_19289,N_19029);
and UO_1746 (O_1746,N_19060,N_19900);
nand UO_1747 (O_1747,N_19838,N_19903);
nand UO_1748 (O_1748,N_19506,N_19230);
and UO_1749 (O_1749,N_19594,N_19824);
xnor UO_1750 (O_1750,N_19223,N_19018);
or UO_1751 (O_1751,N_19786,N_19468);
and UO_1752 (O_1752,N_19304,N_19770);
or UO_1753 (O_1753,N_19611,N_19747);
nand UO_1754 (O_1754,N_19679,N_19976);
and UO_1755 (O_1755,N_19958,N_19237);
or UO_1756 (O_1756,N_19664,N_19845);
nand UO_1757 (O_1757,N_19404,N_19061);
nor UO_1758 (O_1758,N_19081,N_19554);
and UO_1759 (O_1759,N_19923,N_19157);
xor UO_1760 (O_1760,N_19569,N_19860);
or UO_1761 (O_1761,N_19659,N_19274);
nand UO_1762 (O_1762,N_19598,N_19435);
xnor UO_1763 (O_1763,N_19069,N_19983);
and UO_1764 (O_1764,N_19678,N_19983);
and UO_1765 (O_1765,N_19495,N_19290);
and UO_1766 (O_1766,N_19652,N_19775);
and UO_1767 (O_1767,N_19323,N_19851);
nor UO_1768 (O_1768,N_19748,N_19758);
nor UO_1769 (O_1769,N_19769,N_19373);
or UO_1770 (O_1770,N_19659,N_19253);
or UO_1771 (O_1771,N_19558,N_19727);
nand UO_1772 (O_1772,N_19189,N_19206);
nand UO_1773 (O_1773,N_19149,N_19559);
and UO_1774 (O_1774,N_19804,N_19076);
xor UO_1775 (O_1775,N_19497,N_19783);
nand UO_1776 (O_1776,N_19890,N_19728);
nor UO_1777 (O_1777,N_19850,N_19118);
nor UO_1778 (O_1778,N_19490,N_19839);
xnor UO_1779 (O_1779,N_19927,N_19078);
and UO_1780 (O_1780,N_19939,N_19054);
nand UO_1781 (O_1781,N_19042,N_19961);
nor UO_1782 (O_1782,N_19114,N_19770);
xnor UO_1783 (O_1783,N_19343,N_19410);
xnor UO_1784 (O_1784,N_19741,N_19644);
or UO_1785 (O_1785,N_19420,N_19243);
nand UO_1786 (O_1786,N_19221,N_19155);
or UO_1787 (O_1787,N_19036,N_19467);
xor UO_1788 (O_1788,N_19002,N_19611);
and UO_1789 (O_1789,N_19512,N_19207);
xnor UO_1790 (O_1790,N_19527,N_19176);
xnor UO_1791 (O_1791,N_19996,N_19718);
nand UO_1792 (O_1792,N_19541,N_19091);
or UO_1793 (O_1793,N_19515,N_19005);
xnor UO_1794 (O_1794,N_19905,N_19307);
or UO_1795 (O_1795,N_19247,N_19833);
xor UO_1796 (O_1796,N_19071,N_19158);
and UO_1797 (O_1797,N_19674,N_19962);
or UO_1798 (O_1798,N_19276,N_19390);
and UO_1799 (O_1799,N_19380,N_19815);
nor UO_1800 (O_1800,N_19023,N_19038);
or UO_1801 (O_1801,N_19402,N_19698);
xnor UO_1802 (O_1802,N_19937,N_19286);
nand UO_1803 (O_1803,N_19821,N_19810);
and UO_1804 (O_1804,N_19014,N_19047);
and UO_1805 (O_1805,N_19970,N_19259);
nor UO_1806 (O_1806,N_19671,N_19272);
and UO_1807 (O_1807,N_19910,N_19238);
xor UO_1808 (O_1808,N_19094,N_19463);
nor UO_1809 (O_1809,N_19636,N_19013);
xor UO_1810 (O_1810,N_19330,N_19488);
or UO_1811 (O_1811,N_19261,N_19674);
and UO_1812 (O_1812,N_19705,N_19878);
xor UO_1813 (O_1813,N_19039,N_19590);
and UO_1814 (O_1814,N_19863,N_19807);
or UO_1815 (O_1815,N_19894,N_19549);
or UO_1816 (O_1816,N_19181,N_19069);
nor UO_1817 (O_1817,N_19118,N_19814);
xor UO_1818 (O_1818,N_19510,N_19652);
nor UO_1819 (O_1819,N_19990,N_19063);
xor UO_1820 (O_1820,N_19017,N_19669);
nand UO_1821 (O_1821,N_19484,N_19861);
nor UO_1822 (O_1822,N_19101,N_19085);
xor UO_1823 (O_1823,N_19720,N_19281);
xor UO_1824 (O_1824,N_19198,N_19936);
or UO_1825 (O_1825,N_19650,N_19128);
xor UO_1826 (O_1826,N_19238,N_19721);
nor UO_1827 (O_1827,N_19283,N_19987);
xnor UO_1828 (O_1828,N_19646,N_19704);
nand UO_1829 (O_1829,N_19397,N_19616);
or UO_1830 (O_1830,N_19974,N_19418);
xnor UO_1831 (O_1831,N_19403,N_19528);
and UO_1832 (O_1832,N_19179,N_19045);
nand UO_1833 (O_1833,N_19522,N_19286);
or UO_1834 (O_1834,N_19268,N_19720);
nor UO_1835 (O_1835,N_19925,N_19912);
nor UO_1836 (O_1836,N_19001,N_19524);
and UO_1837 (O_1837,N_19272,N_19124);
nand UO_1838 (O_1838,N_19399,N_19467);
nor UO_1839 (O_1839,N_19346,N_19237);
and UO_1840 (O_1840,N_19122,N_19721);
nand UO_1841 (O_1841,N_19738,N_19396);
nor UO_1842 (O_1842,N_19223,N_19862);
nand UO_1843 (O_1843,N_19730,N_19164);
or UO_1844 (O_1844,N_19778,N_19125);
xnor UO_1845 (O_1845,N_19649,N_19963);
nand UO_1846 (O_1846,N_19096,N_19246);
nor UO_1847 (O_1847,N_19011,N_19966);
nand UO_1848 (O_1848,N_19654,N_19947);
nand UO_1849 (O_1849,N_19588,N_19885);
nand UO_1850 (O_1850,N_19166,N_19134);
or UO_1851 (O_1851,N_19976,N_19043);
xnor UO_1852 (O_1852,N_19658,N_19012);
nor UO_1853 (O_1853,N_19977,N_19380);
xor UO_1854 (O_1854,N_19548,N_19516);
or UO_1855 (O_1855,N_19850,N_19342);
nand UO_1856 (O_1856,N_19603,N_19375);
nand UO_1857 (O_1857,N_19747,N_19696);
nand UO_1858 (O_1858,N_19638,N_19585);
or UO_1859 (O_1859,N_19186,N_19632);
nor UO_1860 (O_1860,N_19065,N_19631);
nor UO_1861 (O_1861,N_19456,N_19083);
xnor UO_1862 (O_1862,N_19747,N_19520);
or UO_1863 (O_1863,N_19082,N_19253);
xnor UO_1864 (O_1864,N_19610,N_19499);
xnor UO_1865 (O_1865,N_19446,N_19026);
and UO_1866 (O_1866,N_19540,N_19956);
and UO_1867 (O_1867,N_19711,N_19457);
and UO_1868 (O_1868,N_19206,N_19557);
xor UO_1869 (O_1869,N_19624,N_19193);
and UO_1870 (O_1870,N_19138,N_19097);
nand UO_1871 (O_1871,N_19466,N_19834);
or UO_1872 (O_1872,N_19423,N_19065);
and UO_1873 (O_1873,N_19865,N_19658);
xor UO_1874 (O_1874,N_19420,N_19358);
xor UO_1875 (O_1875,N_19892,N_19390);
nand UO_1876 (O_1876,N_19608,N_19114);
nor UO_1877 (O_1877,N_19335,N_19763);
and UO_1878 (O_1878,N_19485,N_19956);
and UO_1879 (O_1879,N_19829,N_19241);
and UO_1880 (O_1880,N_19758,N_19222);
and UO_1881 (O_1881,N_19288,N_19272);
nor UO_1882 (O_1882,N_19735,N_19231);
or UO_1883 (O_1883,N_19612,N_19391);
nor UO_1884 (O_1884,N_19338,N_19934);
and UO_1885 (O_1885,N_19657,N_19832);
nor UO_1886 (O_1886,N_19196,N_19157);
and UO_1887 (O_1887,N_19774,N_19789);
xnor UO_1888 (O_1888,N_19656,N_19020);
or UO_1889 (O_1889,N_19106,N_19783);
nand UO_1890 (O_1890,N_19926,N_19139);
or UO_1891 (O_1891,N_19196,N_19904);
and UO_1892 (O_1892,N_19301,N_19935);
nand UO_1893 (O_1893,N_19679,N_19920);
xnor UO_1894 (O_1894,N_19839,N_19415);
and UO_1895 (O_1895,N_19380,N_19997);
xor UO_1896 (O_1896,N_19938,N_19758);
nand UO_1897 (O_1897,N_19024,N_19259);
xor UO_1898 (O_1898,N_19890,N_19754);
xnor UO_1899 (O_1899,N_19367,N_19574);
nor UO_1900 (O_1900,N_19212,N_19140);
nand UO_1901 (O_1901,N_19139,N_19948);
xnor UO_1902 (O_1902,N_19274,N_19082);
or UO_1903 (O_1903,N_19464,N_19576);
nand UO_1904 (O_1904,N_19204,N_19833);
nor UO_1905 (O_1905,N_19035,N_19104);
or UO_1906 (O_1906,N_19541,N_19008);
nor UO_1907 (O_1907,N_19992,N_19881);
and UO_1908 (O_1908,N_19836,N_19226);
nand UO_1909 (O_1909,N_19193,N_19646);
and UO_1910 (O_1910,N_19616,N_19198);
and UO_1911 (O_1911,N_19023,N_19820);
and UO_1912 (O_1912,N_19211,N_19790);
nand UO_1913 (O_1913,N_19841,N_19238);
xnor UO_1914 (O_1914,N_19277,N_19734);
nor UO_1915 (O_1915,N_19202,N_19995);
nand UO_1916 (O_1916,N_19788,N_19404);
xnor UO_1917 (O_1917,N_19448,N_19975);
nor UO_1918 (O_1918,N_19347,N_19880);
and UO_1919 (O_1919,N_19707,N_19975);
nand UO_1920 (O_1920,N_19946,N_19053);
xnor UO_1921 (O_1921,N_19256,N_19155);
xor UO_1922 (O_1922,N_19661,N_19768);
nand UO_1923 (O_1923,N_19939,N_19776);
nor UO_1924 (O_1924,N_19655,N_19044);
nand UO_1925 (O_1925,N_19534,N_19008);
xnor UO_1926 (O_1926,N_19672,N_19304);
and UO_1927 (O_1927,N_19041,N_19172);
xnor UO_1928 (O_1928,N_19435,N_19810);
xnor UO_1929 (O_1929,N_19398,N_19516);
xor UO_1930 (O_1930,N_19440,N_19941);
nand UO_1931 (O_1931,N_19246,N_19391);
or UO_1932 (O_1932,N_19096,N_19229);
xnor UO_1933 (O_1933,N_19908,N_19326);
or UO_1934 (O_1934,N_19468,N_19341);
nand UO_1935 (O_1935,N_19140,N_19417);
nor UO_1936 (O_1936,N_19543,N_19457);
nand UO_1937 (O_1937,N_19056,N_19211);
or UO_1938 (O_1938,N_19531,N_19645);
and UO_1939 (O_1939,N_19639,N_19337);
and UO_1940 (O_1940,N_19221,N_19366);
and UO_1941 (O_1941,N_19657,N_19614);
nor UO_1942 (O_1942,N_19927,N_19095);
xnor UO_1943 (O_1943,N_19092,N_19182);
xor UO_1944 (O_1944,N_19556,N_19062);
nand UO_1945 (O_1945,N_19082,N_19495);
or UO_1946 (O_1946,N_19223,N_19361);
nand UO_1947 (O_1947,N_19956,N_19026);
nand UO_1948 (O_1948,N_19176,N_19378);
xnor UO_1949 (O_1949,N_19144,N_19273);
nor UO_1950 (O_1950,N_19574,N_19402);
nor UO_1951 (O_1951,N_19679,N_19115);
xor UO_1952 (O_1952,N_19106,N_19707);
xnor UO_1953 (O_1953,N_19929,N_19118);
or UO_1954 (O_1954,N_19455,N_19210);
or UO_1955 (O_1955,N_19539,N_19268);
and UO_1956 (O_1956,N_19828,N_19403);
xor UO_1957 (O_1957,N_19556,N_19967);
xor UO_1958 (O_1958,N_19790,N_19069);
nand UO_1959 (O_1959,N_19101,N_19803);
or UO_1960 (O_1960,N_19973,N_19835);
or UO_1961 (O_1961,N_19782,N_19757);
and UO_1962 (O_1962,N_19468,N_19686);
nand UO_1963 (O_1963,N_19255,N_19023);
xor UO_1964 (O_1964,N_19880,N_19198);
xor UO_1965 (O_1965,N_19959,N_19186);
or UO_1966 (O_1966,N_19682,N_19128);
xnor UO_1967 (O_1967,N_19196,N_19059);
xor UO_1968 (O_1968,N_19284,N_19022);
nand UO_1969 (O_1969,N_19658,N_19698);
and UO_1970 (O_1970,N_19611,N_19719);
or UO_1971 (O_1971,N_19996,N_19094);
or UO_1972 (O_1972,N_19709,N_19567);
and UO_1973 (O_1973,N_19339,N_19660);
nand UO_1974 (O_1974,N_19946,N_19501);
nand UO_1975 (O_1975,N_19666,N_19300);
xor UO_1976 (O_1976,N_19905,N_19677);
or UO_1977 (O_1977,N_19629,N_19103);
or UO_1978 (O_1978,N_19157,N_19705);
or UO_1979 (O_1979,N_19925,N_19665);
and UO_1980 (O_1980,N_19169,N_19069);
nor UO_1981 (O_1981,N_19146,N_19467);
or UO_1982 (O_1982,N_19180,N_19601);
nand UO_1983 (O_1983,N_19148,N_19364);
or UO_1984 (O_1984,N_19435,N_19033);
nor UO_1985 (O_1985,N_19422,N_19834);
nand UO_1986 (O_1986,N_19310,N_19800);
xnor UO_1987 (O_1987,N_19208,N_19440);
xor UO_1988 (O_1988,N_19095,N_19816);
nor UO_1989 (O_1989,N_19833,N_19423);
nor UO_1990 (O_1990,N_19732,N_19331);
nand UO_1991 (O_1991,N_19113,N_19508);
or UO_1992 (O_1992,N_19780,N_19008);
and UO_1993 (O_1993,N_19071,N_19889);
or UO_1994 (O_1994,N_19437,N_19413);
or UO_1995 (O_1995,N_19723,N_19012);
and UO_1996 (O_1996,N_19723,N_19986);
xnor UO_1997 (O_1997,N_19550,N_19844);
nand UO_1998 (O_1998,N_19787,N_19969);
nor UO_1999 (O_1999,N_19493,N_19782);
or UO_2000 (O_2000,N_19988,N_19032);
or UO_2001 (O_2001,N_19364,N_19335);
or UO_2002 (O_2002,N_19893,N_19971);
xnor UO_2003 (O_2003,N_19351,N_19137);
or UO_2004 (O_2004,N_19028,N_19796);
xor UO_2005 (O_2005,N_19032,N_19227);
nand UO_2006 (O_2006,N_19595,N_19238);
and UO_2007 (O_2007,N_19740,N_19152);
xor UO_2008 (O_2008,N_19713,N_19361);
nand UO_2009 (O_2009,N_19675,N_19120);
nand UO_2010 (O_2010,N_19354,N_19526);
xor UO_2011 (O_2011,N_19816,N_19086);
nor UO_2012 (O_2012,N_19837,N_19272);
nor UO_2013 (O_2013,N_19524,N_19756);
xnor UO_2014 (O_2014,N_19551,N_19091);
xor UO_2015 (O_2015,N_19997,N_19078);
nand UO_2016 (O_2016,N_19949,N_19252);
or UO_2017 (O_2017,N_19332,N_19379);
nor UO_2018 (O_2018,N_19817,N_19115);
xor UO_2019 (O_2019,N_19186,N_19343);
or UO_2020 (O_2020,N_19787,N_19726);
and UO_2021 (O_2021,N_19797,N_19059);
nand UO_2022 (O_2022,N_19599,N_19460);
xnor UO_2023 (O_2023,N_19796,N_19373);
xor UO_2024 (O_2024,N_19344,N_19745);
nand UO_2025 (O_2025,N_19478,N_19049);
nor UO_2026 (O_2026,N_19821,N_19626);
and UO_2027 (O_2027,N_19074,N_19174);
nor UO_2028 (O_2028,N_19775,N_19851);
nand UO_2029 (O_2029,N_19935,N_19097);
or UO_2030 (O_2030,N_19562,N_19021);
xor UO_2031 (O_2031,N_19044,N_19725);
or UO_2032 (O_2032,N_19199,N_19450);
and UO_2033 (O_2033,N_19191,N_19990);
or UO_2034 (O_2034,N_19124,N_19671);
xnor UO_2035 (O_2035,N_19908,N_19597);
and UO_2036 (O_2036,N_19402,N_19673);
nor UO_2037 (O_2037,N_19834,N_19115);
or UO_2038 (O_2038,N_19491,N_19153);
nand UO_2039 (O_2039,N_19802,N_19178);
or UO_2040 (O_2040,N_19608,N_19443);
xor UO_2041 (O_2041,N_19368,N_19042);
nand UO_2042 (O_2042,N_19241,N_19761);
or UO_2043 (O_2043,N_19270,N_19980);
and UO_2044 (O_2044,N_19334,N_19437);
xor UO_2045 (O_2045,N_19363,N_19677);
xnor UO_2046 (O_2046,N_19824,N_19709);
or UO_2047 (O_2047,N_19545,N_19163);
xor UO_2048 (O_2048,N_19437,N_19166);
nand UO_2049 (O_2049,N_19013,N_19444);
nor UO_2050 (O_2050,N_19499,N_19364);
nor UO_2051 (O_2051,N_19680,N_19098);
nand UO_2052 (O_2052,N_19013,N_19575);
nand UO_2053 (O_2053,N_19597,N_19040);
xor UO_2054 (O_2054,N_19149,N_19839);
or UO_2055 (O_2055,N_19274,N_19397);
xor UO_2056 (O_2056,N_19426,N_19127);
nand UO_2057 (O_2057,N_19229,N_19665);
xnor UO_2058 (O_2058,N_19475,N_19844);
xnor UO_2059 (O_2059,N_19043,N_19400);
or UO_2060 (O_2060,N_19219,N_19060);
and UO_2061 (O_2061,N_19013,N_19429);
nand UO_2062 (O_2062,N_19532,N_19221);
nor UO_2063 (O_2063,N_19759,N_19996);
nand UO_2064 (O_2064,N_19281,N_19901);
nor UO_2065 (O_2065,N_19464,N_19036);
nand UO_2066 (O_2066,N_19523,N_19638);
xnor UO_2067 (O_2067,N_19344,N_19602);
xnor UO_2068 (O_2068,N_19523,N_19904);
nor UO_2069 (O_2069,N_19789,N_19281);
xor UO_2070 (O_2070,N_19438,N_19522);
or UO_2071 (O_2071,N_19697,N_19477);
nand UO_2072 (O_2072,N_19939,N_19193);
nand UO_2073 (O_2073,N_19037,N_19411);
xnor UO_2074 (O_2074,N_19396,N_19583);
or UO_2075 (O_2075,N_19131,N_19175);
and UO_2076 (O_2076,N_19301,N_19107);
xnor UO_2077 (O_2077,N_19672,N_19486);
and UO_2078 (O_2078,N_19913,N_19151);
xor UO_2079 (O_2079,N_19032,N_19622);
nor UO_2080 (O_2080,N_19363,N_19107);
and UO_2081 (O_2081,N_19347,N_19543);
or UO_2082 (O_2082,N_19540,N_19070);
xor UO_2083 (O_2083,N_19850,N_19627);
or UO_2084 (O_2084,N_19384,N_19561);
nand UO_2085 (O_2085,N_19322,N_19472);
nor UO_2086 (O_2086,N_19573,N_19438);
xor UO_2087 (O_2087,N_19211,N_19627);
nand UO_2088 (O_2088,N_19038,N_19509);
or UO_2089 (O_2089,N_19516,N_19867);
nor UO_2090 (O_2090,N_19540,N_19709);
nor UO_2091 (O_2091,N_19515,N_19114);
nand UO_2092 (O_2092,N_19767,N_19331);
nor UO_2093 (O_2093,N_19971,N_19341);
or UO_2094 (O_2094,N_19014,N_19951);
and UO_2095 (O_2095,N_19101,N_19249);
nor UO_2096 (O_2096,N_19832,N_19944);
nor UO_2097 (O_2097,N_19912,N_19756);
nand UO_2098 (O_2098,N_19588,N_19032);
nor UO_2099 (O_2099,N_19203,N_19717);
xor UO_2100 (O_2100,N_19797,N_19276);
xnor UO_2101 (O_2101,N_19309,N_19197);
or UO_2102 (O_2102,N_19469,N_19062);
nor UO_2103 (O_2103,N_19615,N_19716);
and UO_2104 (O_2104,N_19144,N_19135);
and UO_2105 (O_2105,N_19114,N_19639);
xnor UO_2106 (O_2106,N_19964,N_19617);
and UO_2107 (O_2107,N_19117,N_19632);
nand UO_2108 (O_2108,N_19472,N_19111);
or UO_2109 (O_2109,N_19366,N_19857);
and UO_2110 (O_2110,N_19333,N_19686);
or UO_2111 (O_2111,N_19120,N_19536);
and UO_2112 (O_2112,N_19576,N_19122);
nand UO_2113 (O_2113,N_19682,N_19549);
or UO_2114 (O_2114,N_19168,N_19308);
nand UO_2115 (O_2115,N_19913,N_19832);
and UO_2116 (O_2116,N_19910,N_19580);
or UO_2117 (O_2117,N_19849,N_19418);
and UO_2118 (O_2118,N_19397,N_19293);
nor UO_2119 (O_2119,N_19628,N_19829);
or UO_2120 (O_2120,N_19389,N_19378);
or UO_2121 (O_2121,N_19651,N_19216);
and UO_2122 (O_2122,N_19151,N_19871);
nand UO_2123 (O_2123,N_19464,N_19639);
nor UO_2124 (O_2124,N_19335,N_19120);
and UO_2125 (O_2125,N_19954,N_19626);
and UO_2126 (O_2126,N_19759,N_19189);
and UO_2127 (O_2127,N_19420,N_19553);
or UO_2128 (O_2128,N_19311,N_19672);
nand UO_2129 (O_2129,N_19430,N_19700);
or UO_2130 (O_2130,N_19394,N_19560);
and UO_2131 (O_2131,N_19664,N_19819);
nand UO_2132 (O_2132,N_19467,N_19654);
nor UO_2133 (O_2133,N_19688,N_19101);
xnor UO_2134 (O_2134,N_19703,N_19955);
nor UO_2135 (O_2135,N_19603,N_19623);
or UO_2136 (O_2136,N_19375,N_19087);
or UO_2137 (O_2137,N_19638,N_19510);
xnor UO_2138 (O_2138,N_19227,N_19797);
nand UO_2139 (O_2139,N_19339,N_19896);
and UO_2140 (O_2140,N_19651,N_19010);
xor UO_2141 (O_2141,N_19445,N_19551);
nand UO_2142 (O_2142,N_19295,N_19384);
nand UO_2143 (O_2143,N_19449,N_19064);
nor UO_2144 (O_2144,N_19141,N_19329);
nor UO_2145 (O_2145,N_19960,N_19397);
nor UO_2146 (O_2146,N_19641,N_19843);
nand UO_2147 (O_2147,N_19899,N_19923);
xor UO_2148 (O_2148,N_19723,N_19333);
or UO_2149 (O_2149,N_19640,N_19460);
or UO_2150 (O_2150,N_19392,N_19530);
nand UO_2151 (O_2151,N_19563,N_19537);
and UO_2152 (O_2152,N_19112,N_19144);
or UO_2153 (O_2153,N_19696,N_19968);
and UO_2154 (O_2154,N_19331,N_19416);
nor UO_2155 (O_2155,N_19564,N_19135);
or UO_2156 (O_2156,N_19551,N_19393);
xor UO_2157 (O_2157,N_19682,N_19448);
and UO_2158 (O_2158,N_19433,N_19878);
nor UO_2159 (O_2159,N_19212,N_19489);
or UO_2160 (O_2160,N_19690,N_19140);
and UO_2161 (O_2161,N_19324,N_19042);
or UO_2162 (O_2162,N_19491,N_19296);
nand UO_2163 (O_2163,N_19721,N_19595);
nand UO_2164 (O_2164,N_19567,N_19699);
nand UO_2165 (O_2165,N_19943,N_19334);
or UO_2166 (O_2166,N_19575,N_19916);
or UO_2167 (O_2167,N_19992,N_19913);
or UO_2168 (O_2168,N_19558,N_19928);
or UO_2169 (O_2169,N_19209,N_19645);
and UO_2170 (O_2170,N_19499,N_19984);
and UO_2171 (O_2171,N_19756,N_19741);
nand UO_2172 (O_2172,N_19171,N_19479);
nor UO_2173 (O_2173,N_19945,N_19987);
nand UO_2174 (O_2174,N_19900,N_19242);
or UO_2175 (O_2175,N_19791,N_19970);
and UO_2176 (O_2176,N_19039,N_19728);
or UO_2177 (O_2177,N_19973,N_19781);
and UO_2178 (O_2178,N_19422,N_19904);
or UO_2179 (O_2179,N_19483,N_19129);
nand UO_2180 (O_2180,N_19369,N_19311);
or UO_2181 (O_2181,N_19697,N_19386);
nor UO_2182 (O_2182,N_19961,N_19848);
nor UO_2183 (O_2183,N_19393,N_19291);
xnor UO_2184 (O_2184,N_19476,N_19136);
or UO_2185 (O_2185,N_19166,N_19712);
nand UO_2186 (O_2186,N_19961,N_19931);
xor UO_2187 (O_2187,N_19647,N_19199);
xnor UO_2188 (O_2188,N_19107,N_19473);
or UO_2189 (O_2189,N_19067,N_19023);
or UO_2190 (O_2190,N_19151,N_19720);
and UO_2191 (O_2191,N_19149,N_19664);
nor UO_2192 (O_2192,N_19875,N_19792);
nand UO_2193 (O_2193,N_19226,N_19327);
nand UO_2194 (O_2194,N_19439,N_19096);
xor UO_2195 (O_2195,N_19844,N_19746);
or UO_2196 (O_2196,N_19620,N_19003);
xnor UO_2197 (O_2197,N_19620,N_19555);
or UO_2198 (O_2198,N_19131,N_19297);
or UO_2199 (O_2199,N_19049,N_19083);
nand UO_2200 (O_2200,N_19110,N_19218);
xnor UO_2201 (O_2201,N_19315,N_19253);
nand UO_2202 (O_2202,N_19612,N_19824);
nand UO_2203 (O_2203,N_19730,N_19488);
nor UO_2204 (O_2204,N_19810,N_19005);
nor UO_2205 (O_2205,N_19957,N_19919);
xor UO_2206 (O_2206,N_19881,N_19816);
or UO_2207 (O_2207,N_19720,N_19547);
nor UO_2208 (O_2208,N_19623,N_19270);
and UO_2209 (O_2209,N_19504,N_19503);
nor UO_2210 (O_2210,N_19200,N_19913);
or UO_2211 (O_2211,N_19262,N_19315);
nor UO_2212 (O_2212,N_19313,N_19253);
nand UO_2213 (O_2213,N_19647,N_19252);
nor UO_2214 (O_2214,N_19816,N_19644);
nand UO_2215 (O_2215,N_19198,N_19647);
nor UO_2216 (O_2216,N_19916,N_19908);
nand UO_2217 (O_2217,N_19425,N_19919);
nand UO_2218 (O_2218,N_19694,N_19113);
nand UO_2219 (O_2219,N_19389,N_19854);
nor UO_2220 (O_2220,N_19149,N_19413);
nor UO_2221 (O_2221,N_19918,N_19367);
and UO_2222 (O_2222,N_19067,N_19910);
and UO_2223 (O_2223,N_19244,N_19085);
or UO_2224 (O_2224,N_19666,N_19329);
nand UO_2225 (O_2225,N_19409,N_19604);
and UO_2226 (O_2226,N_19410,N_19558);
nor UO_2227 (O_2227,N_19412,N_19270);
or UO_2228 (O_2228,N_19519,N_19064);
nand UO_2229 (O_2229,N_19683,N_19607);
and UO_2230 (O_2230,N_19391,N_19947);
nand UO_2231 (O_2231,N_19012,N_19627);
and UO_2232 (O_2232,N_19896,N_19769);
nand UO_2233 (O_2233,N_19268,N_19069);
and UO_2234 (O_2234,N_19781,N_19564);
nor UO_2235 (O_2235,N_19933,N_19994);
nand UO_2236 (O_2236,N_19386,N_19512);
nor UO_2237 (O_2237,N_19184,N_19903);
nor UO_2238 (O_2238,N_19081,N_19586);
xnor UO_2239 (O_2239,N_19018,N_19806);
and UO_2240 (O_2240,N_19769,N_19040);
and UO_2241 (O_2241,N_19493,N_19911);
or UO_2242 (O_2242,N_19286,N_19242);
xnor UO_2243 (O_2243,N_19788,N_19518);
nand UO_2244 (O_2244,N_19033,N_19913);
xnor UO_2245 (O_2245,N_19687,N_19457);
xor UO_2246 (O_2246,N_19152,N_19150);
xor UO_2247 (O_2247,N_19185,N_19655);
nor UO_2248 (O_2248,N_19995,N_19161);
and UO_2249 (O_2249,N_19408,N_19184);
or UO_2250 (O_2250,N_19837,N_19271);
nand UO_2251 (O_2251,N_19729,N_19334);
nand UO_2252 (O_2252,N_19069,N_19779);
or UO_2253 (O_2253,N_19551,N_19970);
nor UO_2254 (O_2254,N_19906,N_19089);
and UO_2255 (O_2255,N_19714,N_19254);
nand UO_2256 (O_2256,N_19684,N_19630);
and UO_2257 (O_2257,N_19041,N_19545);
or UO_2258 (O_2258,N_19494,N_19132);
nand UO_2259 (O_2259,N_19750,N_19228);
and UO_2260 (O_2260,N_19488,N_19007);
nand UO_2261 (O_2261,N_19998,N_19626);
and UO_2262 (O_2262,N_19090,N_19708);
nor UO_2263 (O_2263,N_19046,N_19583);
nor UO_2264 (O_2264,N_19403,N_19583);
nand UO_2265 (O_2265,N_19352,N_19208);
xnor UO_2266 (O_2266,N_19846,N_19836);
or UO_2267 (O_2267,N_19826,N_19048);
and UO_2268 (O_2268,N_19570,N_19086);
or UO_2269 (O_2269,N_19963,N_19003);
or UO_2270 (O_2270,N_19008,N_19451);
xor UO_2271 (O_2271,N_19011,N_19158);
and UO_2272 (O_2272,N_19262,N_19972);
and UO_2273 (O_2273,N_19028,N_19375);
and UO_2274 (O_2274,N_19850,N_19478);
xnor UO_2275 (O_2275,N_19158,N_19918);
and UO_2276 (O_2276,N_19277,N_19773);
nor UO_2277 (O_2277,N_19069,N_19947);
and UO_2278 (O_2278,N_19617,N_19412);
nand UO_2279 (O_2279,N_19122,N_19116);
nor UO_2280 (O_2280,N_19603,N_19589);
nor UO_2281 (O_2281,N_19870,N_19707);
xor UO_2282 (O_2282,N_19940,N_19334);
or UO_2283 (O_2283,N_19493,N_19599);
or UO_2284 (O_2284,N_19894,N_19820);
nand UO_2285 (O_2285,N_19816,N_19115);
nand UO_2286 (O_2286,N_19663,N_19276);
nand UO_2287 (O_2287,N_19083,N_19777);
nor UO_2288 (O_2288,N_19253,N_19644);
and UO_2289 (O_2289,N_19604,N_19020);
nand UO_2290 (O_2290,N_19491,N_19787);
nor UO_2291 (O_2291,N_19246,N_19821);
nor UO_2292 (O_2292,N_19160,N_19571);
nor UO_2293 (O_2293,N_19197,N_19541);
nor UO_2294 (O_2294,N_19087,N_19267);
nand UO_2295 (O_2295,N_19337,N_19612);
nor UO_2296 (O_2296,N_19190,N_19663);
and UO_2297 (O_2297,N_19692,N_19467);
or UO_2298 (O_2298,N_19296,N_19414);
nor UO_2299 (O_2299,N_19497,N_19269);
nand UO_2300 (O_2300,N_19610,N_19779);
and UO_2301 (O_2301,N_19387,N_19837);
nor UO_2302 (O_2302,N_19211,N_19709);
nor UO_2303 (O_2303,N_19761,N_19528);
nor UO_2304 (O_2304,N_19275,N_19890);
or UO_2305 (O_2305,N_19322,N_19523);
nand UO_2306 (O_2306,N_19329,N_19380);
xor UO_2307 (O_2307,N_19730,N_19994);
and UO_2308 (O_2308,N_19946,N_19575);
nor UO_2309 (O_2309,N_19296,N_19960);
nor UO_2310 (O_2310,N_19969,N_19186);
and UO_2311 (O_2311,N_19099,N_19835);
or UO_2312 (O_2312,N_19197,N_19049);
nor UO_2313 (O_2313,N_19928,N_19879);
and UO_2314 (O_2314,N_19726,N_19040);
nand UO_2315 (O_2315,N_19973,N_19429);
and UO_2316 (O_2316,N_19446,N_19340);
xor UO_2317 (O_2317,N_19054,N_19315);
and UO_2318 (O_2318,N_19878,N_19748);
or UO_2319 (O_2319,N_19397,N_19071);
and UO_2320 (O_2320,N_19560,N_19639);
nor UO_2321 (O_2321,N_19701,N_19260);
nand UO_2322 (O_2322,N_19326,N_19469);
nor UO_2323 (O_2323,N_19652,N_19228);
or UO_2324 (O_2324,N_19326,N_19945);
nor UO_2325 (O_2325,N_19391,N_19737);
nand UO_2326 (O_2326,N_19357,N_19276);
and UO_2327 (O_2327,N_19368,N_19077);
or UO_2328 (O_2328,N_19443,N_19009);
nor UO_2329 (O_2329,N_19044,N_19611);
xor UO_2330 (O_2330,N_19390,N_19398);
nand UO_2331 (O_2331,N_19907,N_19995);
nor UO_2332 (O_2332,N_19097,N_19828);
and UO_2333 (O_2333,N_19832,N_19928);
nor UO_2334 (O_2334,N_19177,N_19758);
or UO_2335 (O_2335,N_19803,N_19523);
nor UO_2336 (O_2336,N_19367,N_19245);
xnor UO_2337 (O_2337,N_19711,N_19098);
nand UO_2338 (O_2338,N_19280,N_19522);
nand UO_2339 (O_2339,N_19169,N_19460);
and UO_2340 (O_2340,N_19457,N_19849);
nor UO_2341 (O_2341,N_19494,N_19975);
and UO_2342 (O_2342,N_19563,N_19039);
nor UO_2343 (O_2343,N_19083,N_19625);
nor UO_2344 (O_2344,N_19921,N_19710);
nand UO_2345 (O_2345,N_19414,N_19198);
or UO_2346 (O_2346,N_19333,N_19234);
xnor UO_2347 (O_2347,N_19294,N_19086);
nand UO_2348 (O_2348,N_19893,N_19369);
and UO_2349 (O_2349,N_19284,N_19554);
or UO_2350 (O_2350,N_19415,N_19085);
or UO_2351 (O_2351,N_19557,N_19009);
nor UO_2352 (O_2352,N_19130,N_19120);
and UO_2353 (O_2353,N_19343,N_19511);
or UO_2354 (O_2354,N_19177,N_19415);
or UO_2355 (O_2355,N_19442,N_19610);
xnor UO_2356 (O_2356,N_19158,N_19579);
xor UO_2357 (O_2357,N_19703,N_19664);
nand UO_2358 (O_2358,N_19280,N_19018);
or UO_2359 (O_2359,N_19447,N_19400);
nor UO_2360 (O_2360,N_19960,N_19838);
or UO_2361 (O_2361,N_19865,N_19268);
and UO_2362 (O_2362,N_19131,N_19363);
nor UO_2363 (O_2363,N_19307,N_19421);
xnor UO_2364 (O_2364,N_19922,N_19544);
nand UO_2365 (O_2365,N_19763,N_19695);
or UO_2366 (O_2366,N_19449,N_19504);
or UO_2367 (O_2367,N_19228,N_19368);
nor UO_2368 (O_2368,N_19684,N_19665);
or UO_2369 (O_2369,N_19554,N_19180);
or UO_2370 (O_2370,N_19913,N_19676);
or UO_2371 (O_2371,N_19063,N_19948);
or UO_2372 (O_2372,N_19803,N_19996);
or UO_2373 (O_2373,N_19026,N_19985);
nand UO_2374 (O_2374,N_19100,N_19508);
or UO_2375 (O_2375,N_19070,N_19922);
or UO_2376 (O_2376,N_19247,N_19718);
xnor UO_2377 (O_2377,N_19485,N_19951);
xnor UO_2378 (O_2378,N_19534,N_19447);
xor UO_2379 (O_2379,N_19620,N_19614);
xnor UO_2380 (O_2380,N_19212,N_19582);
nor UO_2381 (O_2381,N_19156,N_19373);
and UO_2382 (O_2382,N_19324,N_19011);
and UO_2383 (O_2383,N_19139,N_19842);
xnor UO_2384 (O_2384,N_19245,N_19744);
nand UO_2385 (O_2385,N_19751,N_19860);
nand UO_2386 (O_2386,N_19040,N_19333);
or UO_2387 (O_2387,N_19665,N_19324);
xnor UO_2388 (O_2388,N_19198,N_19285);
or UO_2389 (O_2389,N_19350,N_19105);
nand UO_2390 (O_2390,N_19655,N_19906);
or UO_2391 (O_2391,N_19197,N_19652);
xnor UO_2392 (O_2392,N_19147,N_19341);
nand UO_2393 (O_2393,N_19288,N_19499);
nor UO_2394 (O_2394,N_19934,N_19499);
xnor UO_2395 (O_2395,N_19731,N_19961);
nor UO_2396 (O_2396,N_19548,N_19197);
xor UO_2397 (O_2397,N_19888,N_19495);
xnor UO_2398 (O_2398,N_19641,N_19795);
nand UO_2399 (O_2399,N_19410,N_19188);
nand UO_2400 (O_2400,N_19259,N_19968);
or UO_2401 (O_2401,N_19360,N_19607);
and UO_2402 (O_2402,N_19531,N_19145);
and UO_2403 (O_2403,N_19679,N_19771);
and UO_2404 (O_2404,N_19542,N_19904);
nor UO_2405 (O_2405,N_19861,N_19482);
xnor UO_2406 (O_2406,N_19833,N_19747);
nand UO_2407 (O_2407,N_19413,N_19143);
xor UO_2408 (O_2408,N_19456,N_19424);
nand UO_2409 (O_2409,N_19686,N_19976);
nand UO_2410 (O_2410,N_19704,N_19966);
nor UO_2411 (O_2411,N_19377,N_19353);
xnor UO_2412 (O_2412,N_19906,N_19949);
or UO_2413 (O_2413,N_19367,N_19018);
nor UO_2414 (O_2414,N_19550,N_19071);
nand UO_2415 (O_2415,N_19089,N_19843);
nand UO_2416 (O_2416,N_19497,N_19545);
nor UO_2417 (O_2417,N_19321,N_19817);
xor UO_2418 (O_2418,N_19793,N_19811);
nor UO_2419 (O_2419,N_19758,N_19221);
and UO_2420 (O_2420,N_19421,N_19183);
xor UO_2421 (O_2421,N_19563,N_19248);
or UO_2422 (O_2422,N_19693,N_19305);
nand UO_2423 (O_2423,N_19810,N_19229);
nand UO_2424 (O_2424,N_19863,N_19400);
nor UO_2425 (O_2425,N_19133,N_19673);
xnor UO_2426 (O_2426,N_19965,N_19664);
nor UO_2427 (O_2427,N_19322,N_19147);
nand UO_2428 (O_2428,N_19863,N_19595);
or UO_2429 (O_2429,N_19168,N_19688);
or UO_2430 (O_2430,N_19515,N_19662);
xor UO_2431 (O_2431,N_19966,N_19988);
xnor UO_2432 (O_2432,N_19321,N_19475);
or UO_2433 (O_2433,N_19534,N_19812);
or UO_2434 (O_2434,N_19500,N_19055);
and UO_2435 (O_2435,N_19572,N_19759);
xnor UO_2436 (O_2436,N_19084,N_19086);
nand UO_2437 (O_2437,N_19451,N_19220);
or UO_2438 (O_2438,N_19254,N_19820);
nor UO_2439 (O_2439,N_19200,N_19579);
nand UO_2440 (O_2440,N_19646,N_19919);
nand UO_2441 (O_2441,N_19985,N_19147);
and UO_2442 (O_2442,N_19668,N_19036);
xnor UO_2443 (O_2443,N_19036,N_19948);
nor UO_2444 (O_2444,N_19534,N_19728);
or UO_2445 (O_2445,N_19003,N_19082);
nand UO_2446 (O_2446,N_19099,N_19054);
nor UO_2447 (O_2447,N_19593,N_19357);
xnor UO_2448 (O_2448,N_19821,N_19714);
xor UO_2449 (O_2449,N_19509,N_19949);
nor UO_2450 (O_2450,N_19553,N_19628);
xor UO_2451 (O_2451,N_19702,N_19100);
xnor UO_2452 (O_2452,N_19182,N_19090);
nor UO_2453 (O_2453,N_19675,N_19602);
nand UO_2454 (O_2454,N_19739,N_19359);
nor UO_2455 (O_2455,N_19098,N_19473);
xnor UO_2456 (O_2456,N_19542,N_19218);
or UO_2457 (O_2457,N_19065,N_19100);
or UO_2458 (O_2458,N_19295,N_19444);
or UO_2459 (O_2459,N_19199,N_19947);
nand UO_2460 (O_2460,N_19374,N_19917);
nor UO_2461 (O_2461,N_19031,N_19635);
nand UO_2462 (O_2462,N_19288,N_19918);
nand UO_2463 (O_2463,N_19566,N_19244);
nand UO_2464 (O_2464,N_19389,N_19133);
or UO_2465 (O_2465,N_19898,N_19866);
nand UO_2466 (O_2466,N_19937,N_19892);
nand UO_2467 (O_2467,N_19014,N_19055);
nor UO_2468 (O_2468,N_19328,N_19353);
nor UO_2469 (O_2469,N_19359,N_19131);
nand UO_2470 (O_2470,N_19020,N_19086);
nor UO_2471 (O_2471,N_19429,N_19464);
nor UO_2472 (O_2472,N_19160,N_19651);
xor UO_2473 (O_2473,N_19595,N_19948);
xor UO_2474 (O_2474,N_19974,N_19617);
and UO_2475 (O_2475,N_19950,N_19838);
nor UO_2476 (O_2476,N_19846,N_19863);
nor UO_2477 (O_2477,N_19517,N_19831);
and UO_2478 (O_2478,N_19821,N_19751);
and UO_2479 (O_2479,N_19206,N_19344);
nand UO_2480 (O_2480,N_19180,N_19319);
or UO_2481 (O_2481,N_19854,N_19467);
nor UO_2482 (O_2482,N_19509,N_19301);
and UO_2483 (O_2483,N_19672,N_19857);
xor UO_2484 (O_2484,N_19343,N_19744);
nand UO_2485 (O_2485,N_19124,N_19799);
nand UO_2486 (O_2486,N_19761,N_19308);
nand UO_2487 (O_2487,N_19384,N_19901);
or UO_2488 (O_2488,N_19436,N_19727);
xor UO_2489 (O_2489,N_19527,N_19289);
xor UO_2490 (O_2490,N_19740,N_19904);
or UO_2491 (O_2491,N_19565,N_19281);
xor UO_2492 (O_2492,N_19845,N_19627);
and UO_2493 (O_2493,N_19459,N_19505);
nand UO_2494 (O_2494,N_19567,N_19146);
xor UO_2495 (O_2495,N_19933,N_19218);
xnor UO_2496 (O_2496,N_19768,N_19913);
nor UO_2497 (O_2497,N_19737,N_19787);
and UO_2498 (O_2498,N_19397,N_19599);
or UO_2499 (O_2499,N_19179,N_19302);
endmodule