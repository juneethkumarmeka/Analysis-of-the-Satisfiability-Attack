module basic_1000_10000_1500_5_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_715,In_905);
nand U1 (N_1,In_970,In_76);
nand U2 (N_2,In_925,In_12);
and U3 (N_3,In_588,In_286);
nand U4 (N_4,In_277,In_834);
nand U5 (N_5,In_274,In_315);
or U6 (N_6,In_882,In_42);
xnor U7 (N_7,In_46,In_309);
nor U8 (N_8,In_145,In_654);
or U9 (N_9,In_320,In_785);
or U10 (N_10,In_541,In_466);
and U11 (N_11,In_267,In_125);
nand U12 (N_12,In_199,In_17);
nand U13 (N_13,In_531,In_305);
nor U14 (N_14,In_36,In_415);
or U15 (N_15,In_604,In_405);
and U16 (N_16,In_381,In_816);
and U17 (N_17,In_867,In_573);
or U18 (N_18,In_741,In_49);
nand U19 (N_19,In_656,In_845);
xor U20 (N_20,In_175,In_211);
nand U21 (N_21,In_689,In_294);
and U22 (N_22,In_410,In_234);
or U23 (N_23,In_28,In_404);
or U24 (N_24,In_943,In_120);
nand U25 (N_25,In_424,In_457);
nor U26 (N_26,In_141,In_701);
or U27 (N_27,In_92,In_853);
xnor U28 (N_28,In_321,In_215);
nand U29 (N_29,In_40,In_184);
nor U30 (N_30,In_408,In_1);
and U31 (N_31,In_505,In_468);
or U32 (N_32,In_190,In_124);
and U33 (N_33,In_583,In_868);
or U34 (N_34,In_13,In_712);
nor U35 (N_35,In_345,In_978);
and U36 (N_36,In_461,In_403);
or U37 (N_37,In_479,In_940);
nand U38 (N_38,In_959,In_126);
nand U39 (N_39,In_751,In_709);
nor U40 (N_40,In_729,In_929);
nor U41 (N_41,In_714,In_795);
nor U42 (N_42,In_976,In_284);
and U43 (N_43,In_969,In_987);
and U44 (N_44,In_744,In_938);
nand U45 (N_45,In_891,In_365);
nand U46 (N_46,In_792,In_26);
nor U47 (N_47,In_844,In_396);
and U48 (N_48,In_972,In_140);
and U49 (N_49,In_734,In_310);
or U50 (N_50,In_39,In_19);
nor U51 (N_51,In_463,In_643);
and U52 (N_52,In_576,In_172);
nand U53 (N_53,In_551,In_133);
nand U54 (N_54,In_559,In_219);
nor U55 (N_55,In_149,In_524);
and U56 (N_56,In_10,In_776);
nor U57 (N_57,In_870,In_808);
or U58 (N_58,In_176,In_766);
xor U59 (N_59,In_979,In_961);
and U60 (N_60,In_733,In_653);
nor U61 (N_61,In_83,In_798);
or U62 (N_62,In_630,In_183);
nor U63 (N_63,In_813,In_455);
nand U64 (N_64,In_991,In_413);
xnor U65 (N_65,In_349,In_809);
and U66 (N_66,In_241,In_258);
and U67 (N_67,In_333,In_409);
or U68 (N_68,In_150,In_567);
and U69 (N_69,In_535,In_691);
or U70 (N_70,In_862,In_412);
xor U71 (N_71,In_780,In_803);
and U72 (N_72,In_562,In_717);
nor U73 (N_73,In_248,In_121);
nand U74 (N_74,In_693,In_949);
or U75 (N_75,In_101,In_810);
and U76 (N_76,In_486,In_429);
and U77 (N_77,In_113,In_936);
nor U78 (N_78,In_552,In_253);
or U79 (N_79,In_600,In_962);
and U80 (N_80,In_406,In_569);
and U81 (N_81,In_871,In_740);
nor U82 (N_82,In_617,In_446);
nor U83 (N_83,In_613,In_843);
or U84 (N_84,In_932,In_484);
nand U85 (N_85,In_30,In_492);
nor U86 (N_86,In_330,In_865);
nand U87 (N_87,In_671,In_584);
and U88 (N_88,In_655,In_433);
nor U89 (N_89,In_638,In_912);
nor U90 (N_90,In_303,In_883);
and U91 (N_91,In_119,In_922);
nand U92 (N_92,In_517,In_821);
nand U93 (N_93,In_84,In_478);
or U94 (N_94,In_47,In_591);
or U95 (N_95,In_775,In_243);
nor U96 (N_96,In_346,In_550);
and U97 (N_97,In_289,In_366);
nand U98 (N_98,In_35,In_516);
nor U99 (N_99,In_34,In_580);
nor U100 (N_100,In_112,In_157);
nor U101 (N_101,In_33,In_896);
nand U102 (N_102,In_635,In_364);
nand U103 (N_103,In_271,In_755);
nand U104 (N_104,In_933,In_449);
and U105 (N_105,In_759,In_279);
or U106 (N_106,In_828,In_838);
nand U107 (N_107,In_38,In_168);
xor U108 (N_108,In_518,In_439);
or U109 (N_109,In_702,In_213);
nand U110 (N_110,In_134,In_687);
and U111 (N_111,In_207,In_866);
or U112 (N_112,In_238,In_898);
nand U113 (N_113,In_308,In_826);
and U114 (N_114,In_765,In_422);
nand U115 (N_115,In_787,In_437);
nor U116 (N_116,In_166,In_363);
and U117 (N_117,In_615,In_908);
or U118 (N_118,In_41,In_391);
nor U119 (N_119,In_738,In_37);
nand U120 (N_120,In_859,In_779);
xor U121 (N_121,In_358,In_87);
nand U122 (N_122,In_105,In_444);
or U123 (N_123,In_226,In_489);
and U124 (N_124,In_512,In_95);
nand U125 (N_125,In_343,In_244);
xnor U126 (N_126,In_189,In_103);
nor U127 (N_127,In_490,In_454);
and U128 (N_128,In_980,In_863);
and U129 (N_129,In_0,In_957);
xor U130 (N_130,In_616,In_416);
and U131 (N_131,In_662,In_470);
nor U132 (N_132,In_778,In_414);
nor U133 (N_133,In_235,In_262);
xor U134 (N_134,In_706,In_43);
nand U135 (N_135,In_663,In_532);
or U136 (N_136,In_625,In_677);
and U137 (N_137,In_388,In_137);
or U138 (N_138,In_963,In_22);
or U139 (N_139,In_692,In_476);
and U140 (N_140,In_749,In_132);
nor U141 (N_141,In_228,In_748);
or U142 (N_142,In_138,In_621);
and U143 (N_143,In_839,In_440);
nand U144 (N_144,In_469,In_370);
or U145 (N_145,In_68,In_288);
xnor U146 (N_146,In_220,In_678);
nand U147 (N_147,In_180,In_682);
or U148 (N_148,In_475,In_393);
or U149 (N_149,In_57,In_864);
or U150 (N_150,In_283,In_32);
or U151 (N_151,In_306,In_993);
nand U152 (N_152,In_718,In_764);
nand U153 (N_153,In_716,In_769);
nand U154 (N_154,In_254,In_328);
and U155 (N_155,In_231,In_597);
and U156 (N_156,In_911,In_639);
or U157 (N_157,In_300,In_148);
nand U158 (N_158,In_225,In_118);
or U159 (N_159,In_102,In_699);
nand U160 (N_160,In_667,In_688);
nand U161 (N_161,In_886,In_135);
xor U162 (N_162,In_571,In_165);
xor U163 (N_163,In_216,In_392);
xor U164 (N_164,In_452,In_467);
and U165 (N_165,In_772,In_472);
nand U166 (N_166,In_601,In_144);
nor U167 (N_167,In_881,In_955);
and U168 (N_168,In_636,In_272);
nand U169 (N_169,In_160,In_934);
nand U170 (N_170,In_623,In_572);
nor U171 (N_171,In_298,In_61);
xor U172 (N_172,In_106,In_739);
xnor U173 (N_173,In_510,In_622);
and U174 (N_174,In_927,In_494);
nor U175 (N_175,In_21,In_768);
or U176 (N_176,In_992,In_669);
nor U177 (N_177,In_756,In_852);
nand U178 (N_178,In_163,In_586);
nand U179 (N_179,In_158,In_182);
or U180 (N_180,In_773,In_265);
nand U181 (N_181,In_177,In_117);
nor U182 (N_182,In_425,In_256);
nor U183 (N_183,In_534,In_435);
nand U184 (N_184,In_607,In_958);
xnor U185 (N_185,In_214,In_337);
xor U186 (N_186,In_703,In_338);
or U187 (N_187,In_450,In_673);
or U188 (N_188,In_371,In_218);
nand U189 (N_189,In_782,In_788);
and U190 (N_190,In_200,In_944);
nand U191 (N_191,In_27,In_194);
nand U192 (N_192,In_796,In_115);
xor U193 (N_193,In_626,In_841);
or U194 (N_194,In_89,In_602);
nand U195 (N_195,In_201,In_317);
nor U196 (N_196,In_998,In_760);
nand U197 (N_197,In_546,In_947);
and U198 (N_198,In_67,In_640);
nand U199 (N_199,In_974,In_694);
nand U200 (N_200,In_786,In_418);
nand U201 (N_201,In_167,In_5);
nand U202 (N_202,In_523,In_227);
nand U203 (N_203,In_842,In_521);
and U204 (N_204,In_916,In_423);
or U205 (N_205,In_316,In_445);
or U206 (N_206,In_268,In_743);
and U207 (N_207,In_977,In_155);
nand U208 (N_208,In_64,In_968);
or U209 (N_209,In_975,In_665);
and U210 (N_210,In_335,In_884);
nand U211 (N_211,In_185,In_456);
nand U212 (N_212,In_192,In_65);
or U213 (N_213,In_649,In_372);
or U214 (N_214,In_173,In_915);
nor U215 (N_215,In_686,In_252);
nand U216 (N_216,In_221,In_637);
nand U217 (N_217,In_924,In_985);
nand U218 (N_218,In_417,In_605);
nor U219 (N_219,In_910,In_889);
or U220 (N_220,In_606,In_77);
or U221 (N_221,In_98,In_485);
nor U222 (N_222,In_246,In_250);
nor U223 (N_223,In_156,In_731);
xor U224 (N_224,In_100,In_645);
nand U225 (N_225,In_596,In_614);
and U226 (N_226,In_983,In_350);
or U227 (N_227,In_685,In_483);
xnor U228 (N_228,In_697,In_888);
nor U229 (N_229,In_368,In_251);
nand U230 (N_230,In_984,In_212);
or U231 (N_231,In_432,In_539);
nor U232 (N_232,In_402,In_482);
or U233 (N_233,In_362,In_502);
or U234 (N_234,In_641,In_946);
nor U235 (N_235,In_698,In_63);
or U236 (N_236,In_754,In_202);
and U237 (N_237,In_887,In_96);
or U238 (N_238,In_585,In_179);
or U239 (N_239,In_762,In_874);
and U240 (N_240,In_619,In_610);
or U241 (N_241,In_812,In_836);
nand U242 (N_242,In_942,In_847);
nand U243 (N_243,In_726,In_644);
nor U244 (N_244,In_81,In_4);
and U245 (N_245,In_603,In_59);
and U246 (N_246,In_442,In_544);
nor U247 (N_247,In_509,In_123);
and U248 (N_248,In_728,In_264);
nand U249 (N_249,In_428,In_334);
nor U250 (N_250,In_147,In_481);
nor U251 (N_251,In_507,In_823);
xor U252 (N_252,In_477,In_579);
nand U253 (N_253,In_713,In_761);
and U254 (N_254,In_263,In_259);
xor U255 (N_255,In_835,In_690);
or U256 (N_256,In_837,In_822);
xor U257 (N_257,In_914,In_491);
and U258 (N_258,In_127,In_290);
nor U259 (N_259,In_909,In_831);
xnor U260 (N_260,In_131,In_169);
nor U261 (N_261,In_570,In_74);
nor U262 (N_262,In_850,In_727);
or U263 (N_263,In_892,In_800);
nor U264 (N_264,In_462,In_648);
or U265 (N_265,In_58,In_496);
xor U266 (N_266,In_849,In_400);
or U267 (N_267,In_876,In_598);
nand U268 (N_268,In_820,In_797);
nor U269 (N_269,In_608,In_854);
or U270 (N_270,In_878,In_783);
nand U271 (N_271,In_520,In_275);
and U272 (N_272,In_632,In_558);
nor U273 (N_273,In_53,In_599);
nor U274 (N_274,In_767,In_758);
or U275 (N_275,In_564,In_695);
and U276 (N_276,In_210,In_443);
nand U277 (N_277,In_893,In_676);
or U278 (N_278,In_497,In_3);
nor U279 (N_279,In_356,In_411);
and U280 (N_280,In_390,In_270);
or U281 (N_281,In_198,In_23);
and U282 (N_282,In_581,In_860);
or U283 (N_283,In_229,In_15);
or U284 (N_284,In_178,In_730);
nand U285 (N_285,In_122,In_487);
nand U286 (N_286,In_965,In_735);
and U287 (N_287,In_8,In_378);
and U288 (N_288,In_500,In_331);
and U289 (N_289,In_661,In_668);
xor U290 (N_290,In_872,In_217);
or U291 (N_291,In_186,In_276);
nor U292 (N_292,In_561,In_858);
xnor U293 (N_293,In_273,In_143);
and U294 (N_294,In_926,In_170);
or U295 (N_295,In_672,In_151);
xor U296 (N_296,In_574,In_78);
or U297 (N_297,In_825,In_548);
nand U298 (N_298,In_397,In_684);
or U299 (N_299,In_436,In_700);
and U300 (N_300,In_827,In_664);
and U301 (N_301,In_931,In_139);
or U302 (N_302,In_318,In_856);
and U303 (N_303,In_563,In_543);
nand U304 (N_304,In_832,In_913);
or U305 (N_305,In_249,In_312);
xor U306 (N_306,In_746,In_997);
nand U307 (N_307,In_204,In_376);
and U308 (N_308,In_20,In_332);
nand U309 (N_309,In_257,In_447);
xnor U310 (N_310,In_503,In_181);
or U311 (N_311,In_973,In_385);
xor U312 (N_312,In_811,In_285);
xor U313 (N_313,In_994,In_611);
or U314 (N_314,In_361,In_110);
nand U315 (N_315,In_819,In_879);
nand U316 (N_316,In_996,In_995);
and U317 (N_317,In_594,In_681);
nor U318 (N_318,In_593,In_885);
nand U319 (N_319,In_899,In_73);
or U320 (N_320,In_56,In_195);
or U321 (N_321,In_525,In_627);
and U322 (N_322,In_794,In_419);
nand U323 (N_323,In_880,In_79);
nor U324 (N_324,In_162,In_322);
and U325 (N_325,In_116,In_130);
or U326 (N_326,In_399,In_292);
or U327 (N_327,In_154,In_287);
or U328 (N_328,In_960,In_474);
and U329 (N_329,In_624,In_986);
and U330 (N_330,In_651,In_80);
nor U331 (N_331,In_679,In_398);
or U332 (N_332,In_86,In_919);
nand U333 (N_333,In_2,In_725);
and U334 (N_334,In_302,In_982);
nand U335 (N_335,In_193,In_945);
and U336 (N_336,In_347,In_242);
and U337 (N_337,In_777,In_704);
nor U338 (N_338,In_557,In_519);
nor U339 (N_339,In_556,In_451);
nand U340 (N_340,In_367,In_774);
and U341 (N_341,In_107,In_565);
nor U342 (N_342,In_188,In_353);
or U343 (N_343,In_595,In_465);
nand U344 (N_344,In_72,In_511);
or U345 (N_345,In_705,In_950);
or U346 (N_346,In_935,In_266);
or U347 (N_347,In_784,In_757);
xnor U348 (N_348,In_25,In_920);
and U349 (N_349,In_325,In_815);
nor U350 (N_350,In_314,In_374);
and U351 (N_351,In_848,In_710);
xor U352 (N_352,In_747,In_501);
or U353 (N_353,In_642,In_51);
and U354 (N_354,In_473,In_69);
nor U355 (N_355,In_869,In_24);
or U356 (N_356,In_395,In_989);
nand U357 (N_357,In_97,In_877);
nand U358 (N_358,In_171,In_261);
nor U359 (N_359,In_537,In_71);
xnor U360 (N_360,In_904,In_545);
or U361 (N_361,In_313,In_458);
nand U362 (N_362,In_952,In_14);
nand U363 (N_363,In_939,In_953);
nand U364 (N_364,In_895,In_508);
or U365 (N_365,In_634,In_674);
nor U366 (N_366,In_921,In_568);
nor U367 (N_367,In_438,In_504);
and U368 (N_368,In_205,In_352);
and U369 (N_369,In_209,In_297);
and U370 (N_370,In_658,In_902);
nand U371 (N_371,In_917,In_354);
nor U372 (N_372,In_951,In_401);
xnor U373 (N_373,In_90,In_582);
nor U374 (N_374,In_633,In_529);
and U375 (N_375,In_357,In_964);
and U376 (N_376,In_805,In_708);
and U377 (N_377,In_351,In_495);
nand U378 (N_378,In_384,In_675);
xor U379 (N_379,In_722,In_488);
nand U380 (N_380,In_480,In_434);
and U381 (N_381,In_161,In_324);
nor U382 (N_382,In_631,In_136);
or U383 (N_383,In_245,In_196);
or U384 (N_384,In_441,In_281);
nand U385 (N_385,In_814,In_799);
nand U386 (N_386,In_628,In_377);
nor U387 (N_387,In_99,In_547);
and U388 (N_388,In_301,In_382);
or U389 (N_389,In_818,In_29);
xnor U390 (N_390,In_319,In_577);
nor U391 (N_391,In_829,In_471);
nor U392 (N_392,In_732,In_903);
and U393 (N_393,In_430,In_770);
and U394 (N_394,In_590,In_239);
xor U395 (N_395,In_514,In_55);
or U396 (N_396,In_533,In_60);
or U397 (N_397,In_720,In_724);
nor U398 (N_398,In_420,In_52);
and U399 (N_399,In_174,In_538);
and U400 (N_400,In_612,In_719);
nor U401 (N_401,In_326,In_448);
or U402 (N_402,In_129,In_379);
nor U403 (N_403,In_223,In_191);
and U404 (N_404,In_578,In_652);
or U405 (N_405,In_875,In_793);
or U406 (N_406,In_269,In_230);
nand U407 (N_407,In_114,In_293);
and U408 (N_408,In_146,In_344);
and U409 (N_409,In_683,In_790);
or U410 (N_410,In_620,In_203);
nor U411 (N_411,In_967,In_498);
nor U412 (N_412,In_70,In_506);
or U413 (N_413,In_771,In_373);
or U414 (N_414,In_948,In_901);
nand U415 (N_415,In_7,In_990);
or U416 (N_416,In_359,In_336);
or U417 (N_417,In_781,In_108);
xor U418 (N_418,In_526,In_791);
nand U419 (N_419,In_629,In_890);
nor U420 (N_420,In_50,In_907);
nor U421 (N_421,In_680,In_342);
and U422 (N_422,In_459,In_530);
or U423 (N_423,In_88,In_369);
nor U424 (N_424,In_553,In_804);
nor U425 (N_425,In_45,In_923);
and U426 (N_426,In_307,In_427);
nor U427 (N_427,In_109,In_763);
or U428 (N_428,In_560,In_752);
or U429 (N_429,In_91,In_299);
xnor U430 (N_430,In_536,In_657);
or U431 (N_431,In_801,In_383);
or U432 (N_432,In_421,In_9);
nand U433 (N_433,In_527,In_515);
or U434 (N_434,In_589,In_240);
nand U435 (N_435,In_966,In_540);
or U436 (N_436,In_522,In_232);
or U437 (N_437,In_750,In_956);
nand U438 (N_438,In_807,In_988);
and U439 (N_439,In_153,In_296);
nand U440 (N_440,In_327,In_855);
or U441 (N_441,In_918,In_295);
or U442 (N_442,In_954,In_873);
or U443 (N_443,In_464,In_206);
nor U444 (N_444,In_111,In_128);
and U445 (N_445,In_493,In_528);
nor U446 (N_446,In_830,In_93);
or U447 (N_447,In_900,In_311);
nor U448 (N_448,In_208,In_609);
or U449 (N_449,In_894,In_360);
nand U450 (N_450,In_387,In_453);
or U451 (N_451,In_44,In_647);
nor U452 (N_452,In_431,In_355);
nand U453 (N_453,In_75,In_670);
nand U454 (N_454,In_971,In_802);
and U455 (N_455,In_696,In_928);
and U456 (N_456,In_164,In_291);
nand U457 (N_457,In_82,In_11);
or U458 (N_458,In_941,In_906);
and U459 (N_459,In_340,In_742);
nand U460 (N_460,In_846,In_323);
or U461 (N_461,In_660,In_85);
xor U462 (N_462,In_389,In_236);
or U463 (N_463,In_566,In_721);
and U464 (N_464,In_280,In_499);
or U465 (N_465,In_260,In_18);
nor U466 (N_466,In_278,In_187);
nor U467 (N_467,In_659,In_426);
xnor U468 (N_468,In_224,In_304);
nand U469 (N_469,In_255,In_375);
and U470 (N_470,In_646,In_618);
or U471 (N_471,In_31,In_861);
and U472 (N_472,In_817,In_66);
or U473 (N_473,In_94,In_6);
or U474 (N_474,In_575,In_897);
or U475 (N_475,In_587,In_407);
and U476 (N_476,In_341,In_937);
nand U477 (N_477,In_753,In_723);
and U478 (N_478,In_707,In_233);
nand U479 (N_479,In_857,In_833);
or U480 (N_480,In_222,In_592);
or U481 (N_481,In_142,In_711);
nand U482 (N_482,In_247,In_999);
and U483 (N_483,In_554,In_48);
and U484 (N_484,In_666,In_197);
or U485 (N_485,In_789,In_394);
or U486 (N_486,In_806,In_650);
nor U487 (N_487,In_62,In_840);
nor U488 (N_488,In_555,In_736);
nor U489 (N_489,In_549,In_851);
or U490 (N_490,In_237,In_930);
and U491 (N_491,In_348,In_339);
or U492 (N_492,In_513,In_824);
or U493 (N_493,In_386,In_104);
xor U494 (N_494,In_16,In_737);
and U495 (N_495,In_542,In_329);
nor U496 (N_496,In_159,In_152);
and U497 (N_497,In_460,In_380);
and U498 (N_498,In_282,In_745);
nor U499 (N_499,In_54,In_981);
or U500 (N_500,In_768,In_263);
or U501 (N_501,In_536,In_464);
and U502 (N_502,In_893,In_456);
xor U503 (N_503,In_690,In_186);
or U504 (N_504,In_378,In_889);
or U505 (N_505,In_453,In_400);
or U506 (N_506,In_293,In_178);
nor U507 (N_507,In_907,In_875);
nand U508 (N_508,In_788,In_266);
nor U509 (N_509,In_580,In_923);
nand U510 (N_510,In_680,In_203);
nor U511 (N_511,In_699,In_42);
nor U512 (N_512,In_525,In_453);
nor U513 (N_513,In_176,In_707);
nor U514 (N_514,In_944,In_1);
and U515 (N_515,In_177,In_681);
or U516 (N_516,In_230,In_853);
and U517 (N_517,In_785,In_560);
nor U518 (N_518,In_743,In_445);
and U519 (N_519,In_2,In_923);
and U520 (N_520,In_827,In_324);
nor U521 (N_521,In_854,In_637);
and U522 (N_522,In_979,In_546);
or U523 (N_523,In_263,In_292);
nand U524 (N_524,In_534,In_390);
nor U525 (N_525,In_618,In_255);
nand U526 (N_526,In_939,In_581);
nand U527 (N_527,In_578,In_317);
nand U528 (N_528,In_458,In_760);
nand U529 (N_529,In_242,In_525);
and U530 (N_530,In_841,In_998);
nor U531 (N_531,In_508,In_699);
or U532 (N_532,In_563,In_222);
and U533 (N_533,In_854,In_503);
or U534 (N_534,In_450,In_415);
nand U535 (N_535,In_385,In_357);
nor U536 (N_536,In_447,In_688);
or U537 (N_537,In_644,In_950);
or U538 (N_538,In_133,In_282);
nor U539 (N_539,In_768,In_104);
and U540 (N_540,In_318,In_198);
nand U541 (N_541,In_712,In_199);
nand U542 (N_542,In_895,In_180);
and U543 (N_543,In_112,In_390);
xor U544 (N_544,In_822,In_916);
or U545 (N_545,In_656,In_749);
and U546 (N_546,In_722,In_729);
and U547 (N_547,In_973,In_410);
xor U548 (N_548,In_958,In_423);
nor U549 (N_549,In_168,In_807);
or U550 (N_550,In_245,In_26);
xnor U551 (N_551,In_741,In_691);
nor U552 (N_552,In_1,In_428);
and U553 (N_553,In_348,In_463);
and U554 (N_554,In_108,In_767);
nor U555 (N_555,In_450,In_355);
nor U556 (N_556,In_348,In_743);
and U557 (N_557,In_118,In_638);
xor U558 (N_558,In_198,In_62);
nand U559 (N_559,In_585,In_702);
nor U560 (N_560,In_983,In_967);
nand U561 (N_561,In_250,In_314);
or U562 (N_562,In_291,In_643);
or U563 (N_563,In_906,In_510);
or U564 (N_564,In_636,In_453);
nand U565 (N_565,In_988,In_303);
or U566 (N_566,In_383,In_701);
and U567 (N_567,In_14,In_374);
nand U568 (N_568,In_889,In_618);
xor U569 (N_569,In_679,In_93);
nand U570 (N_570,In_940,In_204);
or U571 (N_571,In_399,In_177);
or U572 (N_572,In_30,In_218);
or U573 (N_573,In_402,In_822);
nand U574 (N_574,In_762,In_300);
nand U575 (N_575,In_960,In_393);
nand U576 (N_576,In_712,In_768);
and U577 (N_577,In_625,In_757);
nor U578 (N_578,In_578,In_527);
or U579 (N_579,In_132,In_198);
xnor U580 (N_580,In_835,In_4);
nand U581 (N_581,In_779,In_816);
nor U582 (N_582,In_952,In_386);
nand U583 (N_583,In_773,In_936);
or U584 (N_584,In_620,In_709);
nor U585 (N_585,In_58,In_988);
or U586 (N_586,In_65,In_194);
nor U587 (N_587,In_578,In_803);
nor U588 (N_588,In_932,In_202);
nand U589 (N_589,In_34,In_378);
nor U590 (N_590,In_426,In_747);
nor U591 (N_591,In_874,In_636);
and U592 (N_592,In_523,In_826);
nor U593 (N_593,In_529,In_150);
nor U594 (N_594,In_902,In_456);
or U595 (N_595,In_895,In_175);
nor U596 (N_596,In_862,In_765);
nor U597 (N_597,In_744,In_546);
nand U598 (N_598,In_412,In_863);
xor U599 (N_599,In_820,In_560);
nor U600 (N_600,In_318,In_87);
nand U601 (N_601,In_853,In_632);
nand U602 (N_602,In_803,In_705);
nor U603 (N_603,In_494,In_737);
xor U604 (N_604,In_442,In_645);
nand U605 (N_605,In_296,In_387);
xnor U606 (N_606,In_513,In_404);
and U607 (N_607,In_24,In_58);
or U608 (N_608,In_371,In_7);
nand U609 (N_609,In_425,In_460);
nand U610 (N_610,In_414,In_328);
and U611 (N_611,In_296,In_260);
and U612 (N_612,In_908,In_424);
and U613 (N_613,In_830,In_424);
nand U614 (N_614,In_760,In_697);
nand U615 (N_615,In_97,In_186);
nand U616 (N_616,In_749,In_195);
nor U617 (N_617,In_184,In_663);
nand U618 (N_618,In_825,In_64);
nor U619 (N_619,In_768,In_814);
or U620 (N_620,In_552,In_27);
or U621 (N_621,In_641,In_238);
nor U622 (N_622,In_814,In_800);
nand U623 (N_623,In_517,In_355);
or U624 (N_624,In_750,In_726);
nand U625 (N_625,In_372,In_972);
nand U626 (N_626,In_514,In_29);
nand U627 (N_627,In_963,In_609);
nand U628 (N_628,In_286,In_662);
nand U629 (N_629,In_268,In_40);
or U630 (N_630,In_162,In_602);
xor U631 (N_631,In_164,In_223);
and U632 (N_632,In_698,In_821);
nor U633 (N_633,In_441,In_471);
nand U634 (N_634,In_519,In_651);
or U635 (N_635,In_305,In_102);
or U636 (N_636,In_343,In_332);
nand U637 (N_637,In_645,In_293);
or U638 (N_638,In_70,In_690);
nand U639 (N_639,In_258,In_317);
nand U640 (N_640,In_314,In_819);
nand U641 (N_641,In_188,In_336);
nor U642 (N_642,In_911,In_361);
and U643 (N_643,In_984,In_670);
nor U644 (N_644,In_357,In_335);
nor U645 (N_645,In_433,In_521);
and U646 (N_646,In_335,In_529);
or U647 (N_647,In_806,In_415);
nor U648 (N_648,In_97,In_14);
nand U649 (N_649,In_113,In_436);
nand U650 (N_650,In_932,In_13);
nor U651 (N_651,In_508,In_830);
nand U652 (N_652,In_784,In_120);
xor U653 (N_653,In_106,In_627);
nor U654 (N_654,In_411,In_73);
nand U655 (N_655,In_722,In_174);
xor U656 (N_656,In_998,In_27);
and U657 (N_657,In_174,In_252);
or U658 (N_658,In_805,In_656);
nand U659 (N_659,In_579,In_213);
nand U660 (N_660,In_38,In_521);
nor U661 (N_661,In_942,In_296);
or U662 (N_662,In_227,In_54);
and U663 (N_663,In_873,In_264);
nand U664 (N_664,In_156,In_539);
or U665 (N_665,In_598,In_542);
or U666 (N_666,In_309,In_127);
or U667 (N_667,In_864,In_952);
or U668 (N_668,In_355,In_553);
or U669 (N_669,In_817,In_769);
xor U670 (N_670,In_592,In_298);
or U671 (N_671,In_138,In_17);
or U672 (N_672,In_84,In_825);
and U673 (N_673,In_27,In_499);
nor U674 (N_674,In_114,In_667);
nor U675 (N_675,In_797,In_69);
or U676 (N_676,In_686,In_916);
nor U677 (N_677,In_827,In_800);
nor U678 (N_678,In_906,In_896);
or U679 (N_679,In_919,In_79);
and U680 (N_680,In_709,In_546);
and U681 (N_681,In_674,In_834);
and U682 (N_682,In_369,In_709);
or U683 (N_683,In_402,In_731);
and U684 (N_684,In_397,In_452);
nand U685 (N_685,In_115,In_899);
or U686 (N_686,In_503,In_303);
nor U687 (N_687,In_118,In_906);
and U688 (N_688,In_152,In_493);
nor U689 (N_689,In_926,In_814);
or U690 (N_690,In_710,In_284);
nand U691 (N_691,In_896,In_341);
nor U692 (N_692,In_17,In_2);
and U693 (N_693,In_493,In_652);
or U694 (N_694,In_599,In_768);
xor U695 (N_695,In_70,In_855);
and U696 (N_696,In_4,In_600);
or U697 (N_697,In_886,In_679);
nor U698 (N_698,In_630,In_61);
nand U699 (N_699,In_115,In_575);
nand U700 (N_700,In_387,In_898);
nor U701 (N_701,In_976,In_986);
nor U702 (N_702,In_503,In_102);
nand U703 (N_703,In_853,In_356);
nor U704 (N_704,In_346,In_606);
nand U705 (N_705,In_600,In_105);
or U706 (N_706,In_192,In_187);
or U707 (N_707,In_716,In_937);
nand U708 (N_708,In_321,In_199);
or U709 (N_709,In_958,In_155);
or U710 (N_710,In_965,In_333);
nor U711 (N_711,In_71,In_964);
nor U712 (N_712,In_170,In_954);
xor U713 (N_713,In_476,In_264);
or U714 (N_714,In_816,In_416);
or U715 (N_715,In_970,In_239);
nand U716 (N_716,In_891,In_657);
and U717 (N_717,In_115,In_164);
and U718 (N_718,In_70,In_530);
xor U719 (N_719,In_690,In_959);
nand U720 (N_720,In_475,In_455);
or U721 (N_721,In_271,In_576);
xnor U722 (N_722,In_366,In_219);
and U723 (N_723,In_372,In_186);
nor U724 (N_724,In_471,In_487);
or U725 (N_725,In_146,In_709);
nand U726 (N_726,In_184,In_177);
nor U727 (N_727,In_224,In_13);
and U728 (N_728,In_501,In_924);
and U729 (N_729,In_856,In_132);
nor U730 (N_730,In_479,In_531);
nor U731 (N_731,In_811,In_313);
and U732 (N_732,In_715,In_588);
and U733 (N_733,In_998,In_618);
or U734 (N_734,In_629,In_300);
nand U735 (N_735,In_339,In_458);
xor U736 (N_736,In_745,In_450);
nor U737 (N_737,In_834,In_176);
and U738 (N_738,In_929,In_765);
nand U739 (N_739,In_681,In_985);
or U740 (N_740,In_649,In_418);
nand U741 (N_741,In_584,In_545);
nor U742 (N_742,In_79,In_930);
or U743 (N_743,In_489,In_869);
xnor U744 (N_744,In_574,In_285);
and U745 (N_745,In_557,In_242);
nor U746 (N_746,In_106,In_154);
xnor U747 (N_747,In_121,In_739);
xor U748 (N_748,In_953,In_912);
and U749 (N_749,In_292,In_286);
nand U750 (N_750,In_68,In_261);
nor U751 (N_751,In_341,In_153);
and U752 (N_752,In_870,In_273);
nor U753 (N_753,In_221,In_228);
nand U754 (N_754,In_691,In_984);
nand U755 (N_755,In_38,In_772);
or U756 (N_756,In_622,In_131);
and U757 (N_757,In_325,In_185);
nor U758 (N_758,In_468,In_35);
and U759 (N_759,In_689,In_878);
xor U760 (N_760,In_1,In_89);
and U761 (N_761,In_743,In_373);
nand U762 (N_762,In_255,In_729);
and U763 (N_763,In_504,In_155);
nor U764 (N_764,In_614,In_700);
xor U765 (N_765,In_250,In_470);
nand U766 (N_766,In_412,In_263);
or U767 (N_767,In_109,In_837);
nor U768 (N_768,In_319,In_514);
or U769 (N_769,In_562,In_947);
nand U770 (N_770,In_588,In_19);
and U771 (N_771,In_107,In_784);
nor U772 (N_772,In_624,In_662);
or U773 (N_773,In_135,In_597);
nor U774 (N_774,In_187,In_431);
nand U775 (N_775,In_101,In_18);
and U776 (N_776,In_899,In_202);
xor U777 (N_777,In_663,In_880);
nor U778 (N_778,In_387,In_989);
nor U779 (N_779,In_821,In_925);
or U780 (N_780,In_340,In_307);
or U781 (N_781,In_317,In_91);
or U782 (N_782,In_55,In_955);
xnor U783 (N_783,In_339,In_409);
nand U784 (N_784,In_796,In_792);
nor U785 (N_785,In_812,In_135);
and U786 (N_786,In_392,In_124);
nor U787 (N_787,In_46,In_732);
and U788 (N_788,In_328,In_7);
nor U789 (N_789,In_971,In_681);
and U790 (N_790,In_530,In_380);
nor U791 (N_791,In_238,In_91);
nand U792 (N_792,In_426,In_170);
nor U793 (N_793,In_391,In_600);
nor U794 (N_794,In_741,In_622);
nand U795 (N_795,In_34,In_679);
nor U796 (N_796,In_70,In_170);
nand U797 (N_797,In_945,In_24);
nand U798 (N_798,In_628,In_544);
nor U799 (N_799,In_300,In_574);
xnor U800 (N_800,In_80,In_595);
nor U801 (N_801,In_524,In_585);
nor U802 (N_802,In_577,In_387);
and U803 (N_803,In_102,In_141);
nand U804 (N_804,In_948,In_750);
nand U805 (N_805,In_445,In_655);
or U806 (N_806,In_719,In_94);
or U807 (N_807,In_942,In_133);
or U808 (N_808,In_742,In_917);
nand U809 (N_809,In_526,In_230);
or U810 (N_810,In_10,In_317);
and U811 (N_811,In_483,In_506);
or U812 (N_812,In_508,In_562);
and U813 (N_813,In_632,In_68);
or U814 (N_814,In_513,In_782);
and U815 (N_815,In_758,In_214);
xnor U816 (N_816,In_387,In_809);
nor U817 (N_817,In_802,In_767);
nand U818 (N_818,In_351,In_411);
and U819 (N_819,In_348,In_457);
or U820 (N_820,In_166,In_711);
nor U821 (N_821,In_169,In_439);
or U822 (N_822,In_337,In_162);
nand U823 (N_823,In_554,In_529);
nor U824 (N_824,In_582,In_850);
and U825 (N_825,In_189,In_45);
nand U826 (N_826,In_740,In_233);
nand U827 (N_827,In_112,In_284);
nand U828 (N_828,In_428,In_358);
or U829 (N_829,In_644,In_843);
and U830 (N_830,In_902,In_749);
nand U831 (N_831,In_925,In_421);
nand U832 (N_832,In_541,In_393);
or U833 (N_833,In_517,In_60);
and U834 (N_834,In_174,In_508);
or U835 (N_835,In_896,In_506);
nand U836 (N_836,In_324,In_435);
and U837 (N_837,In_226,In_77);
and U838 (N_838,In_772,In_909);
nor U839 (N_839,In_552,In_733);
and U840 (N_840,In_239,In_204);
nor U841 (N_841,In_107,In_115);
nand U842 (N_842,In_898,In_488);
and U843 (N_843,In_696,In_411);
or U844 (N_844,In_66,In_634);
and U845 (N_845,In_627,In_734);
and U846 (N_846,In_602,In_104);
and U847 (N_847,In_27,In_186);
and U848 (N_848,In_857,In_898);
nand U849 (N_849,In_724,In_568);
nor U850 (N_850,In_704,In_758);
or U851 (N_851,In_102,In_323);
and U852 (N_852,In_24,In_0);
nor U853 (N_853,In_919,In_603);
nor U854 (N_854,In_23,In_483);
nand U855 (N_855,In_452,In_193);
nor U856 (N_856,In_228,In_581);
and U857 (N_857,In_709,In_667);
nand U858 (N_858,In_988,In_319);
and U859 (N_859,In_411,In_927);
xnor U860 (N_860,In_299,In_227);
xnor U861 (N_861,In_661,In_440);
nand U862 (N_862,In_566,In_883);
and U863 (N_863,In_440,In_349);
and U864 (N_864,In_950,In_882);
or U865 (N_865,In_224,In_77);
or U866 (N_866,In_348,In_323);
or U867 (N_867,In_278,In_501);
nand U868 (N_868,In_355,In_663);
or U869 (N_869,In_218,In_732);
and U870 (N_870,In_730,In_530);
or U871 (N_871,In_893,In_694);
nor U872 (N_872,In_63,In_357);
or U873 (N_873,In_202,In_643);
and U874 (N_874,In_130,In_420);
or U875 (N_875,In_201,In_153);
nor U876 (N_876,In_415,In_432);
or U877 (N_877,In_964,In_689);
or U878 (N_878,In_26,In_153);
xor U879 (N_879,In_429,In_595);
or U880 (N_880,In_285,In_645);
nand U881 (N_881,In_335,In_417);
and U882 (N_882,In_413,In_65);
xor U883 (N_883,In_555,In_857);
nand U884 (N_884,In_647,In_933);
nor U885 (N_885,In_131,In_160);
nor U886 (N_886,In_699,In_539);
or U887 (N_887,In_256,In_387);
xnor U888 (N_888,In_706,In_228);
or U889 (N_889,In_814,In_441);
or U890 (N_890,In_296,In_900);
or U891 (N_891,In_114,In_179);
and U892 (N_892,In_4,In_104);
nand U893 (N_893,In_694,In_294);
xnor U894 (N_894,In_897,In_166);
nor U895 (N_895,In_841,In_260);
nand U896 (N_896,In_503,In_401);
xor U897 (N_897,In_801,In_565);
and U898 (N_898,In_686,In_229);
or U899 (N_899,In_416,In_40);
or U900 (N_900,In_582,In_159);
and U901 (N_901,In_911,In_347);
or U902 (N_902,In_103,In_641);
or U903 (N_903,In_261,In_642);
nor U904 (N_904,In_836,In_571);
and U905 (N_905,In_267,In_843);
xor U906 (N_906,In_548,In_729);
and U907 (N_907,In_677,In_813);
nor U908 (N_908,In_253,In_44);
nor U909 (N_909,In_718,In_496);
or U910 (N_910,In_523,In_105);
or U911 (N_911,In_102,In_665);
and U912 (N_912,In_887,In_413);
or U913 (N_913,In_7,In_931);
xnor U914 (N_914,In_407,In_137);
and U915 (N_915,In_397,In_111);
nand U916 (N_916,In_434,In_916);
nand U917 (N_917,In_621,In_635);
and U918 (N_918,In_521,In_758);
nand U919 (N_919,In_54,In_671);
and U920 (N_920,In_621,In_912);
nor U921 (N_921,In_565,In_918);
xor U922 (N_922,In_776,In_430);
and U923 (N_923,In_918,In_741);
or U924 (N_924,In_443,In_347);
nor U925 (N_925,In_205,In_289);
or U926 (N_926,In_459,In_736);
nand U927 (N_927,In_810,In_918);
nand U928 (N_928,In_655,In_582);
nand U929 (N_929,In_544,In_935);
and U930 (N_930,In_429,In_288);
nor U931 (N_931,In_973,In_258);
nand U932 (N_932,In_698,In_553);
nand U933 (N_933,In_895,In_466);
nand U934 (N_934,In_758,In_873);
nand U935 (N_935,In_966,In_677);
nand U936 (N_936,In_698,In_278);
xor U937 (N_937,In_853,In_995);
and U938 (N_938,In_760,In_44);
and U939 (N_939,In_524,In_829);
nor U940 (N_940,In_315,In_235);
and U941 (N_941,In_963,In_173);
and U942 (N_942,In_111,In_483);
and U943 (N_943,In_228,In_213);
nor U944 (N_944,In_859,In_940);
or U945 (N_945,In_979,In_912);
and U946 (N_946,In_186,In_192);
nand U947 (N_947,In_88,In_569);
nor U948 (N_948,In_141,In_84);
nor U949 (N_949,In_310,In_376);
nor U950 (N_950,In_729,In_511);
nand U951 (N_951,In_58,In_671);
or U952 (N_952,In_199,In_856);
nand U953 (N_953,In_904,In_655);
nor U954 (N_954,In_306,In_523);
and U955 (N_955,In_287,In_454);
and U956 (N_956,In_148,In_544);
nor U957 (N_957,In_171,In_3);
nand U958 (N_958,In_912,In_407);
and U959 (N_959,In_112,In_742);
nor U960 (N_960,In_983,In_623);
nand U961 (N_961,In_622,In_250);
and U962 (N_962,In_629,In_353);
nor U963 (N_963,In_782,In_351);
and U964 (N_964,In_553,In_923);
nor U965 (N_965,In_182,In_963);
or U966 (N_966,In_557,In_856);
nor U967 (N_967,In_964,In_569);
and U968 (N_968,In_261,In_704);
or U969 (N_969,In_963,In_131);
nand U970 (N_970,In_842,In_809);
nand U971 (N_971,In_50,In_516);
nand U972 (N_972,In_580,In_913);
and U973 (N_973,In_100,In_793);
xnor U974 (N_974,In_210,In_766);
nand U975 (N_975,In_929,In_744);
nor U976 (N_976,In_724,In_772);
nand U977 (N_977,In_748,In_392);
xnor U978 (N_978,In_498,In_40);
xnor U979 (N_979,In_225,In_550);
xor U980 (N_980,In_417,In_407);
nor U981 (N_981,In_263,In_367);
nand U982 (N_982,In_31,In_799);
and U983 (N_983,In_902,In_160);
and U984 (N_984,In_310,In_665);
or U985 (N_985,In_80,In_448);
xnor U986 (N_986,In_199,In_874);
and U987 (N_987,In_61,In_897);
xnor U988 (N_988,In_59,In_264);
xnor U989 (N_989,In_220,In_684);
and U990 (N_990,In_279,In_814);
or U991 (N_991,In_112,In_4);
and U992 (N_992,In_636,In_806);
xnor U993 (N_993,In_409,In_773);
or U994 (N_994,In_647,In_361);
or U995 (N_995,In_728,In_625);
or U996 (N_996,In_581,In_942);
nor U997 (N_997,In_170,In_7);
nand U998 (N_998,In_43,In_785);
and U999 (N_999,In_309,In_750);
nand U1000 (N_1000,In_625,In_825);
and U1001 (N_1001,In_368,In_830);
and U1002 (N_1002,In_938,In_319);
and U1003 (N_1003,In_854,In_616);
nor U1004 (N_1004,In_956,In_1);
and U1005 (N_1005,In_587,In_695);
nor U1006 (N_1006,In_203,In_946);
nand U1007 (N_1007,In_161,In_782);
or U1008 (N_1008,In_76,In_950);
nor U1009 (N_1009,In_577,In_658);
nand U1010 (N_1010,In_308,In_32);
or U1011 (N_1011,In_717,In_586);
and U1012 (N_1012,In_624,In_328);
xnor U1013 (N_1013,In_617,In_712);
or U1014 (N_1014,In_865,In_687);
and U1015 (N_1015,In_938,In_913);
nor U1016 (N_1016,In_795,In_369);
or U1017 (N_1017,In_422,In_151);
nand U1018 (N_1018,In_236,In_401);
and U1019 (N_1019,In_639,In_727);
and U1020 (N_1020,In_650,In_95);
and U1021 (N_1021,In_841,In_828);
nor U1022 (N_1022,In_777,In_448);
xor U1023 (N_1023,In_868,In_557);
or U1024 (N_1024,In_849,In_988);
xnor U1025 (N_1025,In_848,In_885);
nand U1026 (N_1026,In_891,In_258);
nand U1027 (N_1027,In_40,In_168);
nand U1028 (N_1028,In_471,In_513);
xnor U1029 (N_1029,In_719,In_861);
xnor U1030 (N_1030,In_311,In_967);
nor U1031 (N_1031,In_558,In_650);
nor U1032 (N_1032,In_758,In_85);
or U1033 (N_1033,In_623,In_372);
or U1034 (N_1034,In_423,In_657);
or U1035 (N_1035,In_70,In_350);
nand U1036 (N_1036,In_232,In_190);
or U1037 (N_1037,In_376,In_34);
or U1038 (N_1038,In_300,In_761);
and U1039 (N_1039,In_658,In_842);
xor U1040 (N_1040,In_751,In_735);
nor U1041 (N_1041,In_172,In_771);
xnor U1042 (N_1042,In_732,In_733);
or U1043 (N_1043,In_168,In_396);
nor U1044 (N_1044,In_613,In_293);
nor U1045 (N_1045,In_304,In_499);
nand U1046 (N_1046,In_716,In_390);
nand U1047 (N_1047,In_482,In_995);
nand U1048 (N_1048,In_770,In_404);
nand U1049 (N_1049,In_551,In_404);
or U1050 (N_1050,In_761,In_629);
nor U1051 (N_1051,In_342,In_320);
and U1052 (N_1052,In_363,In_127);
nand U1053 (N_1053,In_45,In_478);
or U1054 (N_1054,In_111,In_265);
nand U1055 (N_1055,In_836,In_768);
nand U1056 (N_1056,In_743,In_412);
nor U1057 (N_1057,In_523,In_961);
nand U1058 (N_1058,In_877,In_756);
and U1059 (N_1059,In_601,In_991);
and U1060 (N_1060,In_626,In_890);
or U1061 (N_1061,In_861,In_264);
nor U1062 (N_1062,In_314,In_321);
and U1063 (N_1063,In_778,In_62);
and U1064 (N_1064,In_50,In_142);
xor U1065 (N_1065,In_447,In_829);
nand U1066 (N_1066,In_851,In_916);
xnor U1067 (N_1067,In_800,In_795);
nor U1068 (N_1068,In_605,In_588);
nand U1069 (N_1069,In_296,In_429);
xor U1070 (N_1070,In_229,In_42);
nor U1071 (N_1071,In_637,In_11);
and U1072 (N_1072,In_869,In_813);
nand U1073 (N_1073,In_480,In_162);
nor U1074 (N_1074,In_350,In_926);
nor U1075 (N_1075,In_692,In_191);
nand U1076 (N_1076,In_301,In_75);
nor U1077 (N_1077,In_782,In_38);
and U1078 (N_1078,In_201,In_109);
and U1079 (N_1079,In_548,In_835);
nand U1080 (N_1080,In_557,In_531);
nor U1081 (N_1081,In_415,In_513);
and U1082 (N_1082,In_446,In_153);
xor U1083 (N_1083,In_867,In_920);
or U1084 (N_1084,In_219,In_162);
or U1085 (N_1085,In_294,In_134);
nand U1086 (N_1086,In_789,In_505);
and U1087 (N_1087,In_960,In_594);
nor U1088 (N_1088,In_387,In_997);
or U1089 (N_1089,In_123,In_723);
nand U1090 (N_1090,In_154,In_16);
xor U1091 (N_1091,In_640,In_806);
and U1092 (N_1092,In_673,In_14);
or U1093 (N_1093,In_366,In_320);
nor U1094 (N_1094,In_83,In_841);
nand U1095 (N_1095,In_908,In_71);
or U1096 (N_1096,In_418,In_545);
nand U1097 (N_1097,In_470,In_219);
nor U1098 (N_1098,In_794,In_29);
and U1099 (N_1099,In_96,In_405);
and U1100 (N_1100,In_547,In_167);
xnor U1101 (N_1101,In_516,In_354);
and U1102 (N_1102,In_34,In_918);
or U1103 (N_1103,In_893,In_439);
nand U1104 (N_1104,In_828,In_244);
nand U1105 (N_1105,In_153,In_760);
and U1106 (N_1106,In_85,In_299);
nor U1107 (N_1107,In_507,In_667);
or U1108 (N_1108,In_275,In_858);
or U1109 (N_1109,In_968,In_457);
nand U1110 (N_1110,In_500,In_268);
xor U1111 (N_1111,In_790,In_728);
and U1112 (N_1112,In_711,In_578);
and U1113 (N_1113,In_348,In_905);
or U1114 (N_1114,In_230,In_656);
and U1115 (N_1115,In_235,In_712);
and U1116 (N_1116,In_246,In_177);
and U1117 (N_1117,In_232,In_749);
nor U1118 (N_1118,In_119,In_286);
nor U1119 (N_1119,In_821,In_581);
nand U1120 (N_1120,In_413,In_781);
and U1121 (N_1121,In_174,In_893);
xor U1122 (N_1122,In_956,In_735);
nor U1123 (N_1123,In_389,In_395);
nor U1124 (N_1124,In_693,In_799);
nand U1125 (N_1125,In_172,In_132);
xor U1126 (N_1126,In_490,In_12);
nor U1127 (N_1127,In_466,In_79);
or U1128 (N_1128,In_885,In_524);
or U1129 (N_1129,In_684,In_147);
nor U1130 (N_1130,In_455,In_90);
or U1131 (N_1131,In_545,In_896);
nand U1132 (N_1132,In_70,In_688);
or U1133 (N_1133,In_580,In_270);
nor U1134 (N_1134,In_105,In_594);
and U1135 (N_1135,In_833,In_332);
nand U1136 (N_1136,In_935,In_104);
and U1137 (N_1137,In_404,In_344);
and U1138 (N_1138,In_285,In_999);
or U1139 (N_1139,In_268,In_44);
or U1140 (N_1140,In_501,In_426);
and U1141 (N_1141,In_681,In_585);
nor U1142 (N_1142,In_38,In_723);
or U1143 (N_1143,In_352,In_388);
nand U1144 (N_1144,In_127,In_953);
xor U1145 (N_1145,In_768,In_749);
and U1146 (N_1146,In_351,In_825);
nor U1147 (N_1147,In_532,In_78);
xnor U1148 (N_1148,In_426,In_508);
and U1149 (N_1149,In_455,In_429);
nor U1150 (N_1150,In_503,In_626);
nor U1151 (N_1151,In_140,In_980);
and U1152 (N_1152,In_849,In_465);
nand U1153 (N_1153,In_130,In_687);
and U1154 (N_1154,In_423,In_435);
nor U1155 (N_1155,In_574,In_32);
nand U1156 (N_1156,In_924,In_689);
or U1157 (N_1157,In_431,In_254);
nor U1158 (N_1158,In_544,In_233);
or U1159 (N_1159,In_352,In_982);
xor U1160 (N_1160,In_979,In_767);
or U1161 (N_1161,In_25,In_850);
nand U1162 (N_1162,In_760,In_854);
or U1163 (N_1163,In_817,In_127);
nand U1164 (N_1164,In_390,In_492);
xnor U1165 (N_1165,In_770,In_806);
nand U1166 (N_1166,In_696,In_427);
or U1167 (N_1167,In_582,In_740);
or U1168 (N_1168,In_314,In_931);
nor U1169 (N_1169,In_592,In_145);
nor U1170 (N_1170,In_24,In_572);
and U1171 (N_1171,In_264,In_644);
nor U1172 (N_1172,In_360,In_150);
nor U1173 (N_1173,In_266,In_523);
nor U1174 (N_1174,In_573,In_119);
xnor U1175 (N_1175,In_614,In_934);
xor U1176 (N_1176,In_324,In_113);
or U1177 (N_1177,In_599,In_117);
and U1178 (N_1178,In_76,In_899);
nand U1179 (N_1179,In_471,In_822);
nand U1180 (N_1180,In_264,In_760);
and U1181 (N_1181,In_432,In_352);
or U1182 (N_1182,In_152,In_849);
or U1183 (N_1183,In_494,In_52);
nor U1184 (N_1184,In_571,In_233);
or U1185 (N_1185,In_654,In_622);
or U1186 (N_1186,In_864,In_382);
xor U1187 (N_1187,In_797,In_653);
or U1188 (N_1188,In_36,In_654);
nor U1189 (N_1189,In_663,In_228);
nand U1190 (N_1190,In_763,In_136);
and U1191 (N_1191,In_415,In_192);
xnor U1192 (N_1192,In_577,In_864);
nand U1193 (N_1193,In_534,In_197);
nor U1194 (N_1194,In_280,In_304);
xnor U1195 (N_1195,In_224,In_328);
nand U1196 (N_1196,In_685,In_506);
and U1197 (N_1197,In_838,In_579);
or U1198 (N_1198,In_882,In_66);
nor U1199 (N_1199,In_712,In_456);
and U1200 (N_1200,In_628,In_336);
and U1201 (N_1201,In_621,In_747);
nor U1202 (N_1202,In_539,In_685);
nand U1203 (N_1203,In_563,In_494);
xnor U1204 (N_1204,In_953,In_172);
or U1205 (N_1205,In_882,In_688);
nand U1206 (N_1206,In_677,In_652);
nand U1207 (N_1207,In_908,In_241);
nor U1208 (N_1208,In_360,In_701);
nor U1209 (N_1209,In_5,In_85);
nand U1210 (N_1210,In_301,In_626);
nand U1211 (N_1211,In_962,In_845);
and U1212 (N_1212,In_951,In_735);
nand U1213 (N_1213,In_294,In_326);
or U1214 (N_1214,In_88,In_309);
and U1215 (N_1215,In_310,In_890);
nand U1216 (N_1216,In_576,In_427);
and U1217 (N_1217,In_699,In_13);
and U1218 (N_1218,In_280,In_712);
nand U1219 (N_1219,In_819,In_930);
nand U1220 (N_1220,In_794,In_757);
nor U1221 (N_1221,In_546,In_723);
nand U1222 (N_1222,In_568,In_134);
and U1223 (N_1223,In_840,In_140);
nand U1224 (N_1224,In_205,In_824);
and U1225 (N_1225,In_369,In_3);
nor U1226 (N_1226,In_22,In_5);
nand U1227 (N_1227,In_840,In_27);
nor U1228 (N_1228,In_797,In_53);
and U1229 (N_1229,In_924,In_769);
or U1230 (N_1230,In_424,In_47);
xnor U1231 (N_1231,In_94,In_811);
nand U1232 (N_1232,In_362,In_553);
or U1233 (N_1233,In_47,In_293);
and U1234 (N_1234,In_869,In_194);
nand U1235 (N_1235,In_753,In_391);
nand U1236 (N_1236,In_718,In_594);
nor U1237 (N_1237,In_492,In_256);
nand U1238 (N_1238,In_394,In_162);
nand U1239 (N_1239,In_778,In_160);
nor U1240 (N_1240,In_712,In_573);
xor U1241 (N_1241,In_943,In_51);
or U1242 (N_1242,In_498,In_689);
or U1243 (N_1243,In_512,In_192);
or U1244 (N_1244,In_466,In_223);
nor U1245 (N_1245,In_508,In_59);
and U1246 (N_1246,In_614,In_472);
or U1247 (N_1247,In_166,In_127);
nand U1248 (N_1248,In_911,In_925);
nor U1249 (N_1249,In_232,In_607);
and U1250 (N_1250,In_191,In_435);
nand U1251 (N_1251,In_436,In_782);
or U1252 (N_1252,In_613,In_139);
nand U1253 (N_1253,In_455,In_300);
nand U1254 (N_1254,In_376,In_546);
nand U1255 (N_1255,In_537,In_761);
nor U1256 (N_1256,In_251,In_853);
or U1257 (N_1257,In_514,In_460);
and U1258 (N_1258,In_472,In_343);
or U1259 (N_1259,In_897,In_790);
or U1260 (N_1260,In_152,In_576);
nor U1261 (N_1261,In_268,In_299);
nand U1262 (N_1262,In_200,In_708);
or U1263 (N_1263,In_212,In_224);
nor U1264 (N_1264,In_135,In_499);
nor U1265 (N_1265,In_484,In_412);
nand U1266 (N_1266,In_143,In_964);
and U1267 (N_1267,In_490,In_365);
or U1268 (N_1268,In_54,In_563);
and U1269 (N_1269,In_989,In_99);
or U1270 (N_1270,In_559,In_981);
nor U1271 (N_1271,In_133,In_545);
nor U1272 (N_1272,In_446,In_906);
xnor U1273 (N_1273,In_902,In_387);
and U1274 (N_1274,In_74,In_64);
or U1275 (N_1275,In_237,In_849);
nor U1276 (N_1276,In_402,In_875);
nand U1277 (N_1277,In_536,In_895);
nor U1278 (N_1278,In_893,In_440);
or U1279 (N_1279,In_105,In_29);
xnor U1280 (N_1280,In_766,In_603);
nor U1281 (N_1281,In_928,In_400);
or U1282 (N_1282,In_365,In_186);
or U1283 (N_1283,In_696,In_715);
nor U1284 (N_1284,In_758,In_539);
nor U1285 (N_1285,In_712,In_513);
or U1286 (N_1286,In_52,In_922);
or U1287 (N_1287,In_541,In_484);
nand U1288 (N_1288,In_731,In_677);
and U1289 (N_1289,In_497,In_314);
or U1290 (N_1290,In_555,In_91);
nand U1291 (N_1291,In_882,In_939);
and U1292 (N_1292,In_225,In_510);
and U1293 (N_1293,In_181,In_743);
xor U1294 (N_1294,In_302,In_930);
and U1295 (N_1295,In_923,In_72);
or U1296 (N_1296,In_216,In_441);
and U1297 (N_1297,In_325,In_548);
and U1298 (N_1298,In_204,In_48);
and U1299 (N_1299,In_435,In_247);
nor U1300 (N_1300,In_286,In_766);
and U1301 (N_1301,In_132,In_587);
or U1302 (N_1302,In_761,In_779);
nor U1303 (N_1303,In_681,In_886);
xnor U1304 (N_1304,In_467,In_159);
or U1305 (N_1305,In_657,In_250);
nand U1306 (N_1306,In_666,In_805);
nor U1307 (N_1307,In_815,In_231);
nor U1308 (N_1308,In_653,In_349);
xor U1309 (N_1309,In_993,In_963);
xnor U1310 (N_1310,In_5,In_388);
nor U1311 (N_1311,In_772,In_956);
nor U1312 (N_1312,In_896,In_898);
xor U1313 (N_1313,In_124,In_141);
nand U1314 (N_1314,In_701,In_960);
and U1315 (N_1315,In_481,In_965);
xnor U1316 (N_1316,In_555,In_70);
and U1317 (N_1317,In_410,In_948);
or U1318 (N_1318,In_861,In_799);
nand U1319 (N_1319,In_102,In_149);
nand U1320 (N_1320,In_557,In_815);
nand U1321 (N_1321,In_455,In_826);
nand U1322 (N_1322,In_689,In_11);
and U1323 (N_1323,In_328,In_460);
and U1324 (N_1324,In_142,In_726);
or U1325 (N_1325,In_464,In_605);
or U1326 (N_1326,In_160,In_90);
nor U1327 (N_1327,In_557,In_349);
and U1328 (N_1328,In_673,In_472);
or U1329 (N_1329,In_204,In_319);
or U1330 (N_1330,In_537,In_845);
and U1331 (N_1331,In_359,In_431);
nor U1332 (N_1332,In_163,In_439);
nor U1333 (N_1333,In_165,In_68);
and U1334 (N_1334,In_87,In_887);
and U1335 (N_1335,In_62,In_804);
or U1336 (N_1336,In_196,In_780);
and U1337 (N_1337,In_774,In_331);
and U1338 (N_1338,In_154,In_139);
nand U1339 (N_1339,In_320,In_201);
nor U1340 (N_1340,In_164,In_782);
or U1341 (N_1341,In_524,In_907);
or U1342 (N_1342,In_906,In_337);
or U1343 (N_1343,In_276,In_882);
nand U1344 (N_1344,In_468,In_917);
nand U1345 (N_1345,In_576,In_870);
nand U1346 (N_1346,In_335,In_610);
nor U1347 (N_1347,In_319,In_209);
xor U1348 (N_1348,In_872,In_508);
and U1349 (N_1349,In_468,In_771);
or U1350 (N_1350,In_370,In_403);
and U1351 (N_1351,In_891,In_121);
nand U1352 (N_1352,In_944,In_788);
or U1353 (N_1353,In_178,In_585);
nand U1354 (N_1354,In_216,In_457);
and U1355 (N_1355,In_653,In_357);
nor U1356 (N_1356,In_384,In_776);
or U1357 (N_1357,In_315,In_298);
nand U1358 (N_1358,In_734,In_513);
nor U1359 (N_1359,In_158,In_434);
or U1360 (N_1360,In_649,In_509);
nand U1361 (N_1361,In_150,In_478);
xor U1362 (N_1362,In_829,In_942);
and U1363 (N_1363,In_937,In_840);
or U1364 (N_1364,In_524,In_221);
nor U1365 (N_1365,In_261,In_873);
nand U1366 (N_1366,In_747,In_663);
nor U1367 (N_1367,In_460,In_60);
and U1368 (N_1368,In_649,In_171);
and U1369 (N_1369,In_990,In_271);
nor U1370 (N_1370,In_965,In_272);
or U1371 (N_1371,In_486,In_557);
nand U1372 (N_1372,In_413,In_993);
nor U1373 (N_1373,In_672,In_859);
and U1374 (N_1374,In_596,In_479);
nand U1375 (N_1375,In_773,In_924);
or U1376 (N_1376,In_36,In_862);
or U1377 (N_1377,In_851,In_608);
or U1378 (N_1378,In_814,In_335);
xor U1379 (N_1379,In_743,In_720);
and U1380 (N_1380,In_590,In_643);
and U1381 (N_1381,In_551,In_618);
and U1382 (N_1382,In_808,In_482);
and U1383 (N_1383,In_553,In_450);
and U1384 (N_1384,In_918,In_170);
or U1385 (N_1385,In_429,In_113);
nand U1386 (N_1386,In_170,In_671);
nand U1387 (N_1387,In_591,In_569);
nand U1388 (N_1388,In_269,In_47);
xnor U1389 (N_1389,In_924,In_13);
or U1390 (N_1390,In_328,In_476);
nor U1391 (N_1391,In_19,In_682);
or U1392 (N_1392,In_904,In_874);
or U1393 (N_1393,In_924,In_881);
nor U1394 (N_1394,In_291,In_570);
nor U1395 (N_1395,In_965,In_86);
or U1396 (N_1396,In_500,In_519);
xor U1397 (N_1397,In_890,In_995);
xor U1398 (N_1398,In_669,In_807);
nand U1399 (N_1399,In_544,In_987);
xor U1400 (N_1400,In_179,In_766);
nor U1401 (N_1401,In_886,In_677);
xor U1402 (N_1402,In_445,In_309);
nor U1403 (N_1403,In_532,In_50);
nor U1404 (N_1404,In_366,In_89);
nand U1405 (N_1405,In_340,In_568);
nor U1406 (N_1406,In_529,In_487);
or U1407 (N_1407,In_888,In_348);
and U1408 (N_1408,In_708,In_251);
xnor U1409 (N_1409,In_971,In_172);
or U1410 (N_1410,In_234,In_194);
or U1411 (N_1411,In_412,In_248);
or U1412 (N_1412,In_457,In_370);
or U1413 (N_1413,In_380,In_169);
nand U1414 (N_1414,In_582,In_538);
or U1415 (N_1415,In_150,In_640);
nor U1416 (N_1416,In_195,In_483);
or U1417 (N_1417,In_702,In_266);
nand U1418 (N_1418,In_54,In_216);
or U1419 (N_1419,In_442,In_18);
and U1420 (N_1420,In_650,In_471);
nor U1421 (N_1421,In_894,In_879);
and U1422 (N_1422,In_591,In_519);
nand U1423 (N_1423,In_107,In_79);
nand U1424 (N_1424,In_34,In_909);
nor U1425 (N_1425,In_328,In_751);
nor U1426 (N_1426,In_230,In_668);
and U1427 (N_1427,In_136,In_772);
xor U1428 (N_1428,In_540,In_193);
and U1429 (N_1429,In_866,In_456);
and U1430 (N_1430,In_987,In_527);
or U1431 (N_1431,In_582,In_827);
and U1432 (N_1432,In_354,In_601);
nand U1433 (N_1433,In_948,In_929);
or U1434 (N_1434,In_80,In_42);
or U1435 (N_1435,In_445,In_669);
nand U1436 (N_1436,In_372,In_232);
nand U1437 (N_1437,In_75,In_151);
and U1438 (N_1438,In_428,In_635);
nor U1439 (N_1439,In_944,In_480);
nand U1440 (N_1440,In_502,In_379);
and U1441 (N_1441,In_727,In_18);
nor U1442 (N_1442,In_614,In_453);
and U1443 (N_1443,In_623,In_366);
nand U1444 (N_1444,In_768,In_793);
or U1445 (N_1445,In_60,In_511);
nor U1446 (N_1446,In_840,In_884);
and U1447 (N_1447,In_410,In_595);
or U1448 (N_1448,In_730,In_241);
and U1449 (N_1449,In_686,In_388);
nand U1450 (N_1450,In_767,In_454);
nand U1451 (N_1451,In_801,In_599);
nor U1452 (N_1452,In_242,In_326);
nor U1453 (N_1453,In_963,In_220);
and U1454 (N_1454,In_27,In_112);
nand U1455 (N_1455,In_661,In_618);
nand U1456 (N_1456,In_95,In_210);
nor U1457 (N_1457,In_982,In_425);
and U1458 (N_1458,In_640,In_811);
and U1459 (N_1459,In_944,In_848);
and U1460 (N_1460,In_553,In_421);
and U1461 (N_1461,In_899,In_310);
or U1462 (N_1462,In_52,In_992);
and U1463 (N_1463,In_277,In_987);
and U1464 (N_1464,In_678,In_2);
xnor U1465 (N_1465,In_646,In_927);
or U1466 (N_1466,In_791,In_302);
xnor U1467 (N_1467,In_475,In_564);
nand U1468 (N_1468,In_175,In_208);
nor U1469 (N_1469,In_526,In_80);
and U1470 (N_1470,In_35,In_512);
xor U1471 (N_1471,In_384,In_946);
nor U1472 (N_1472,In_441,In_550);
nor U1473 (N_1473,In_456,In_359);
nor U1474 (N_1474,In_909,In_257);
or U1475 (N_1475,In_482,In_590);
and U1476 (N_1476,In_774,In_952);
or U1477 (N_1477,In_375,In_755);
nor U1478 (N_1478,In_391,In_916);
nand U1479 (N_1479,In_121,In_72);
or U1480 (N_1480,In_250,In_993);
nor U1481 (N_1481,In_427,In_734);
nand U1482 (N_1482,In_501,In_928);
and U1483 (N_1483,In_186,In_927);
xnor U1484 (N_1484,In_248,In_234);
nand U1485 (N_1485,In_669,In_279);
nor U1486 (N_1486,In_321,In_675);
or U1487 (N_1487,In_128,In_313);
xor U1488 (N_1488,In_751,In_707);
and U1489 (N_1489,In_677,In_998);
nand U1490 (N_1490,In_202,In_910);
nand U1491 (N_1491,In_594,In_144);
nand U1492 (N_1492,In_479,In_670);
or U1493 (N_1493,In_648,In_734);
and U1494 (N_1494,In_127,In_228);
or U1495 (N_1495,In_743,In_345);
or U1496 (N_1496,In_597,In_592);
or U1497 (N_1497,In_813,In_843);
nor U1498 (N_1498,In_157,In_540);
and U1499 (N_1499,In_701,In_915);
and U1500 (N_1500,In_532,In_614);
nand U1501 (N_1501,In_109,In_165);
nand U1502 (N_1502,In_210,In_613);
nor U1503 (N_1503,In_180,In_397);
and U1504 (N_1504,In_289,In_868);
xnor U1505 (N_1505,In_309,In_436);
nor U1506 (N_1506,In_57,In_0);
or U1507 (N_1507,In_272,In_620);
and U1508 (N_1508,In_465,In_277);
nor U1509 (N_1509,In_963,In_828);
or U1510 (N_1510,In_239,In_798);
nand U1511 (N_1511,In_40,In_165);
and U1512 (N_1512,In_336,In_1);
or U1513 (N_1513,In_835,In_673);
xor U1514 (N_1514,In_948,In_914);
xor U1515 (N_1515,In_718,In_562);
and U1516 (N_1516,In_33,In_275);
nor U1517 (N_1517,In_579,In_424);
nand U1518 (N_1518,In_842,In_201);
or U1519 (N_1519,In_153,In_14);
nand U1520 (N_1520,In_704,In_298);
nor U1521 (N_1521,In_494,In_978);
and U1522 (N_1522,In_128,In_934);
and U1523 (N_1523,In_3,In_440);
nor U1524 (N_1524,In_273,In_232);
nand U1525 (N_1525,In_78,In_512);
or U1526 (N_1526,In_106,In_364);
nand U1527 (N_1527,In_539,In_225);
or U1528 (N_1528,In_289,In_712);
nor U1529 (N_1529,In_345,In_473);
and U1530 (N_1530,In_381,In_737);
and U1531 (N_1531,In_155,In_378);
nor U1532 (N_1532,In_198,In_263);
or U1533 (N_1533,In_897,In_927);
nand U1534 (N_1534,In_942,In_520);
nand U1535 (N_1535,In_906,In_128);
and U1536 (N_1536,In_214,In_584);
or U1537 (N_1537,In_598,In_430);
nor U1538 (N_1538,In_438,In_96);
or U1539 (N_1539,In_701,In_794);
nand U1540 (N_1540,In_172,In_322);
xnor U1541 (N_1541,In_942,In_779);
and U1542 (N_1542,In_298,In_100);
nor U1543 (N_1543,In_994,In_343);
and U1544 (N_1544,In_299,In_1);
nor U1545 (N_1545,In_374,In_522);
and U1546 (N_1546,In_432,In_268);
or U1547 (N_1547,In_102,In_439);
nand U1548 (N_1548,In_460,In_416);
nor U1549 (N_1549,In_127,In_704);
or U1550 (N_1550,In_726,In_21);
nand U1551 (N_1551,In_922,In_828);
and U1552 (N_1552,In_86,In_725);
and U1553 (N_1553,In_167,In_186);
and U1554 (N_1554,In_444,In_634);
and U1555 (N_1555,In_44,In_423);
nand U1556 (N_1556,In_122,In_489);
xor U1557 (N_1557,In_932,In_697);
and U1558 (N_1558,In_707,In_515);
and U1559 (N_1559,In_634,In_828);
nor U1560 (N_1560,In_228,In_370);
and U1561 (N_1561,In_6,In_662);
nand U1562 (N_1562,In_369,In_54);
nor U1563 (N_1563,In_413,In_753);
or U1564 (N_1564,In_392,In_922);
nor U1565 (N_1565,In_58,In_191);
or U1566 (N_1566,In_863,In_192);
and U1567 (N_1567,In_805,In_388);
nand U1568 (N_1568,In_302,In_843);
or U1569 (N_1569,In_657,In_291);
nor U1570 (N_1570,In_74,In_311);
or U1571 (N_1571,In_4,In_561);
nor U1572 (N_1572,In_148,In_404);
or U1573 (N_1573,In_950,In_973);
nor U1574 (N_1574,In_326,In_69);
xor U1575 (N_1575,In_69,In_653);
nor U1576 (N_1576,In_883,In_891);
nand U1577 (N_1577,In_664,In_536);
nand U1578 (N_1578,In_372,In_194);
nand U1579 (N_1579,In_481,In_105);
or U1580 (N_1580,In_902,In_620);
nor U1581 (N_1581,In_384,In_262);
nand U1582 (N_1582,In_786,In_740);
nand U1583 (N_1583,In_920,In_749);
nor U1584 (N_1584,In_30,In_16);
xnor U1585 (N_1585,In_625,In_693);
nand U1586 (N_1586,In_311,In_680);
or U1587 (N_1587,In_625,In_660);
or U1588 (N_1588,In_867,In_860);
xnor U1589 (N_1589,In_508,In_153);
nor U1590 (N_1590,In_734,In_681);
nor U1591 (N_1591,In_949,In_218);
nand U1592 (N_1592,In_204,In_398);
and U1593 (N_1593,In_828,In_589);
or U1594 (N_1594,In_802,In_861);
nor U1595 (N_1595,In_580,In_668);
nand U1596 (N_1596,In_208,In_86);
nor U1597 (N_1597,In_909,In_829);
or U1598 (N_1598,In_39,In_85);
and U1599 (N_1599,In_578,In_477);
nor U1600 (N_1600,In_210,In_148);
and U1601 (N_1601,In_177,In_436);
nor U1602 (N_1602,In_576,In_734);
nor U1603 (N_1603,In_172,In_850);
nand U1604 (N_1604,In_157,In_996);
and U1605 (N_1605,In_887,In_687);
nor U1606 (N_1606,In_486,In_678);
nand U1607 (N_1607,In_696,In_371);
and U1608 (N_1608,In_774,In_975);
or U1609 (N_1609,In_322,In_383);
and U1610 (N_1610,In_134,In_582);
nand U1611 (N_1611,In_720,In_721);
or U1612 (N_1612,In_70,In_48);
nand U1613 (N_1613,In_455,In_490);
and U1614 (N_1614,In_912,In_170);
or U1615 (N_1615,In_117,In_221);
and U1616 (N_1616,In_213,In_601);
nor U1617 (N_1617,In_85,In_333);
xor U1618 (N_1618,In_6,In_419);
nand U1619 (N_1619,In_543,In_332);
or U1620 (N_1620,In_169,In_336);
and U1621 (N_1621,In_42,In_185);
nor U1622 (N_1622,In_351,In_378);
nor U1623 (N_1623,In_18,In_567);
or U1624 (N_1624,In_370,In_281);
and U1625 (N_1625,In_530,In_687);
nand U1626 (N_1626,In_189,In_672);
nand U1627 (N_1627,In_195,In_169);
or U1628 (N_1628,In_948,In_363);
nand U1629 (N_1629,In_941,In_623);
nand U1630 (N_1630,In_340,In_639);
nor U1631 (N_1631,In_532,In_38);
nor U1632 (N_1632,In_966,In_651);
xor U1633 (N_1633,In_545,In_389);
or U1634 (N_1634,In_68,In_6);
or U1635 (N_1635,In_137,In_592);
xor U1636 (N_1636,In_728,In_605);
or U1637 (N_1637,In_772,In_199);
or U1638 (N_1638,In_117,In_302);
nor U1639 (N_1639,In_309,In_209);
nor U1640 (N_1640,In_549,In_8);
and U1641 (N_1641,In_734,In_598);
or U1642 (N_1642,In_687,In_387);
nand U1643 (N_1643,In_613,In_356);
nand U1644 (N_1644,In_848,In_101);
xnor U1645 (N_1645,In_535,In_375);
nor U1646 (N_1646,In_656,In_815);
and U1647 (N_1647,In_264,In_894);
nand U1648 (N_1648,In_866,In_749);
nand U1649 (N_1649,In_888,In_511);
nor U1650 (N_1650,In_424,In_521);
nor U1651 (N_1651,In_554,In_510);
or U1652 (N_1652,In_346,In_136);
xnor U1653 (N_1653,In_731,In_824);
or U1654 (N_1654,In_835,In_504);
nor U1655 (N_1655,In_758,In_462);
nand U1656 (N_1656,In_4,In_823);
xnor U1657 (N_1657,In_944,In_488);
or U1658 (N_1658,In_205,In_425);
xor U1659 (N_1659,In_32,In_746);
and U1660 (N_1660,In_328,In_43);
nand U1661 (N_1661,In_592,In_843);
nand U1662 (N_1662,In_894,In_259);
nor U1663 (N_1663,In_800,In_579);
nor U1664 (N_1664,In_273,In_641);
and U1665 (N_1665,In_416,In_56);
and U1666 (N_1666,In_964,In_19);
nand U1667 (N_1667,In_733,In_86);
nor U1668 (N_1668,In_215,In_293);
or U1669 (N_1669,In_249,In_851);
or U1670 (N_1670,In_548,In_412);
nor U1671 (N_1671,In_549,In_984);
nand U1672 (N_1672,In_125,In_843);
or U1673 (N_1673,In_523,In_311);
xnor U1674 (N_1674,In_912,In_399);
nand U1675 (N_1675,In_478,In_180);
nand U1676 (N_1676,In_290,In_83);
or U1677 (N_1677,In_795,In_237);
and U1678 (N_1678,In_453,In_745);
or U1679 (N_1679,In_754,In_94);
and U1680 (N_1680,In_102,In_317);
nor U1681 (N_1681,In_718,In_780);
nand U1682 (N_1682,In_448,In_811);
or U1683 (N_1683,In_13,In_240);
xnor U1684 (N_1684,In_502,In_841);
and U1685 (N_1685,In_690,In_385);
nor U1686 (N_1686,In_606,In_532);
or U1687 (N_1687,In_855,In_333);
nor U1688 (N_1688,In_451,In_382);
xor U1689 (N_1689,In_610,In_475);
nand U1690 (N_1690,In_983,In_233);
nand U1691 (N_1691,In_427,In_293);
nor U1692 (N_1692,In_401,In_43);
and U1693 (N_1693,In_814,In_164);
nor U1694 (N_1694,In_886,In_261);
or U1695 (N_1695,In_99,In_632);
nor U1696 (N_1696,In_791,In_427);
and U1697 (N_1697,In_308,In_604);
and U1698 (N_1698,In_157,In_789);
and U1699 (N_1699,In_407,In_164);
nor U1700 (N_1700,In_212,In_466);
or U1701 (N_1701,In_437,In_451);
and U1702 (N_1702,In_829,In_246);
and U1703 (N_1703,In_370,In_332);
or U1704 (N_1704,In_311,In_878);
and U1705 (N_1705,In_839,In_291);
nand U1706 (N_1706,In_189,In_153);
nand U1707 (N_1707,In_237,In_964);
xor U1708 (N_1708,In_595,In_228);
nor U1709 (N_1709,In_498,In_593);
nand U1710 (N_1710,In_357,In_302);
nand U1711 (N_1711,In_661,In_524);
nand U1712 (N_1712,In_920,In_839);
or U1713 (N_1713,In_97,In_789);
nand U1714 (N_1714,In_993,In_973);
and U1715 (N_1715,In_986,In_439);
nor U1716 (N_1716,In_804,In_993);
nor U1717 (N_1717,In_391,In_429);
or U1718 (N_1718,In_187,In_732);
nor U1719 (N_1719,In_711,In_14);
nor U1720 (N_1720,In_365,In_902);
or U1721 (N_1721,In_929,In_277);
and U1722 (N_1722,In_343,In_896);
nand U1723 (N_1723,In_33,In_296);
or U1724 (N_1724,In_548,In_782);
or U1725 (N_1725,In_282,In_687);
nand U1726 (N_1726,In_571,In_939);
or U1727 (N_1727,In_589,In_447);
xnor U1728 (N_1728,In_901,In_946);
nor U1729 (N_1729,In_331,In_954);
xor U1730 (N_1730,In_42,In_753);
nand U1731 (N_1731,In_906,In_815);
nor U1732 (N_1732,In_231,In_274);
or U1733 (N_1733,In_623,In_625);
and U1734 (N_1734,In_872,In_833);
nand U1735 (N_1735,In_669,In_751);
nand U1736 (N_1736,In_296,In_163);
nand U1737 (N_1737,In_175,In_729);
nand U1738 (N_1738,In_221,In_523);
nand U1739 (N_1739,In_630,In_686);
nor U1740 (N_1740,In_560,In_786);
and U1741 (N_1741,In_802,In_247);
nand U1742 (N_1742,In_483,In_858);
nor U1743 (N_1743,In_32,In_874);
or U1744 (N_1744,In_770,In_631);
nand U1745 (N_1745,In_386,In_906);
nand U1746 (N_1746,In_697,In_674);
nand U1747 (N_1747,In_47,In_607);
nor U1748 (N_1748,In_879,In_0);
xnor U1749 (N_1749,In_591,In_515);
nor U1750 (N_1750,In_177,In_794);
or U1751 (N_1751,In_605,In_770);
nor U1752 (N_1752,In_343,In_649);
nor U1753 (N_1753,In_386,In_512);
or U1754 (N_1754,In_443,In_361);
nand U1755 (N_1755,In_941,In_956);
or U1756 (N_1756,In_492,In_576);
or U1757 (N_1757,In_876,In_143);
or U1758 (N_1758,In_359,In_386);
nor U1759 (N_1759,In_424,In_446);
and U1760 (N_1760,In_473,In_323);
nand U1761 (N_1761,In_438,In_289);
and U1762 (N_1762,In_516,In_992);
nor U1763 (N_1763,In_830,In_415);
or U1764 (N_1764,In_832,In_105);
and U1765 (N_1765,In_817,In_855);
or U1766 (N_1766,In_344,In_578);
nor U1767 (N_1767,In_806,In_912);
nor U1768 (N_1768,In_37,In_36);
nand U1769 (N_1769,In_998,In_25);
nand U1770 (N_1770,In_169,In_161);
or U1771 (N_1771,In_609,In_440);
and U1772 (N_1772,In_218,In_134);
and U1773 (N_1773,In_116,In_13);
nor U1774 (N_1774,In_839,In_604);
xor U1775 (N_1775,In_266,In_955);
and U1776 (N_1776,In_646,In_499);
nor U1777 (N_1777,In_33,In_382);
or U1778 (N_1778,In_13,In_52);
and U1779 (N_1779,In_771,In_145);
and U1780 (N_1780,In_641,In_467);
nand U1781 (N_1781,In_554,In_226);
nand U1782 (N_1782,In_89,In_855);
nand U1783 (N_1783,In_387,In_874);
nor U1784 (N_1784,In_217,In_202);
and U1785 (N_1785,In_907,In_893);
or U1786 (N_1786,In_542,In_486);
or U1787 (N_1787,In_713,In_836);
nor U1788 (N_1788,In_680,In_966);
xnor U1789 (N_1789,In_999,In_347);
xor U1790 (N_1790,In_637,In_979);
or U1791 (N_1791,In_48,In_439);
nand U1792 (N_1792,In_422,In_925);
xnor U1793 (N_1793,In_616,In_714);
or U1794 (N_1794,In_960,In_958);
nor U1795 (N_1795,In_385,In_937);
and U1796 (N_1796,In_484,In_530);
and U1797 (N_1797,In_61,In_283);
or U1798 (N_1798,In_950,In_898);
and U1799 (N_1799,In_381,In_757);
nand U1800 (N_1800,In_113,In_194);
and U1801 (N_1801,In_924,In_151);
xor U1802 (N_1802,In_832,In_999);
nand U1803 (N_1803,In_612,In_395);
nand U1804 (N_1804,In_514,In_670);
nor U1805 (N_1805,In_992,In_535);
xnor U1806 (N_1806,In_604,In_548);
or U1807 (N_1807,In_694,In_115);
or U1808 (N_1808,In_672,In_166);
and U1809 (N_1809,In_68,In_903);
or U1810 (N_1810,In_137,In_544);
nor U1811 (N_1811,In_532,In_836);
nand U1812 (N_1812,In_902,In_572);
nand U1813 (N_1813,In_833,In_952);
nor U1814 (N_1814,In_752,In_132);
xor U1815 (N_1815,In_373,In_400);
nand U1816 (N_1816,In_648,In_611);
nand U1817 (N_1817,In_208,In_326);
xor U1818 (N_1818,In_851,In_901);
nor U1819 (N_1819,In_601,In_372);
nand U1820 (N_1820,In_699,In_382);
nor U1821 (N_1821,In_78,In_398);
and U1822 (N_1822,In_68,In_283);
and U1823 (N_1823,In_354,In_355);
and U1824 (N_1824,In_619,In_792);
nor U1825 (N_1825,In_810,In_215);
xnor U1826 (N_1826,In_903,In_282);
or U1827 (N_1827,In_846,In_49);
and U1828 (N_1828,In_416,In_678);
nor U1829 (N_1829,In_584,In_291);
nand U1830 (N_1830,In_369,In_694);
or U1831 (N_1831,In_307,In_699);
xnor U1832 (N_1832,In_252,In_109);
or U1833 (N_1833,In_339,In_404);
and U1834 (N_1834,In_488,In_582);
nor U1835 (N_1835,In_893,In_78);
and U1836 (N_1836,In_481,In_811);
nor U1837 (N_1837,In_333,In_461);
xnor U1838 (N_1838,In_483,In_740);
nand U1839 (N_1839,In_626,In_506);
nand U1840 (N_1840,In_575,In_852);
xnor U1841 (N_1841,In_466,In_815);
and U1842 (N_1842,In_339,In_549);
nand U1843 (N_1843,In_546,In_62);
or U1844 (N_1844,In_125,In_270);
and U1845 (N_1845,In_651,In_144);
nor U1846 (N_1846,In_109,In_204);
or U1847 (N_1847,In_376,In_884);
xor U1848 (N_1848,In_799,In_198);
and U1849 (N_1849,In_506,In_538);
nor U1850 (N_1850,In_956,In_932);
xnor U1851 (N_1851,In_785,In_871);
or U1852 (N_1852,In_653,In_882);
nor U1853 (N_1853,In_166,In_58);
xor U1854 (N_1854,In_875,In_441);
nand U1855 (N_1855,In_466,In_571);
nor U1856 (N_1856,In_507,In_567);
or U1857 (N_1857,In_828,In_398);
nand U1858 (N_1858,In_242,In_141);
or U1859 (N_1859,In_154,In_195);
nand U1860 (N_1860,In_447,In_411);
nand U1861 (N_1861,In_794,In_750);
xor U1862 (N_1862,In_181,In_321);
or U1863 (N_1863,In_216,In_127);
xor U1864 (N_1864,In_651,In_194);
and U1865 (N_1865,In_214,In_244);
nand U1866 (N_1866,In_451,In_395);
nand U1867 (N_1867,In_293,In_484);
nor U1868 (N_1868,In_883,In_448);
nor U1869 (N_1869,In_295,In_690);
or U1870 (N_1870,In_91,In_437);
nand U1871 (N_1871,In_49,In_178);
nor U1872 (N_1872,In_448,In_167);
or U1873 (N_1873,In_190,In_824);
and U1874 (N_1874,In_470,In_780);
nand U1875 (N_1875,In_379,In_453);
or U1876 (N_1876,In_273,In_629);
nor U1877 (N_1877,In_990,In_190);
nor U1878 (N_1878,In_323,In_41);
or U1879 (N_1879,In_520,In_915);
xnor U1880 (N_1880,In_652,In_442);
and U1881 (N_1881,In_499,In_601);
xnor U1882 (N_1882,In_808,In_868);
or U1883 (N_1883,In_568,In_720);
or U1884 (N_1884,In_556,In_957);
or U1885 (N_1885,In_375,In_618);
or U1886 (N_1886,In_71,In_365);
or U1887 (N_1887,In_188,In_863);
and U1888 (N_1888,In_578,In_931);
xnor U1889 (N_1889,In_15,In_582);
or U1890 (N_1890,In_969,In_73);
or U1891 (N_1891,In_645,In_68);
and U1892 (N_1892,In_592,In_938);
nand U1893 (N_1893,In_496,In_758);
xnor U1894 (N_1894,In_119,In_141);
nor U1895 (N_1895,In_782,In_607);
nor U1896 (N_1896,In_292,In_246);
or U1897 (N_1897,In_721,In_768);
nand U1898 (N_1898,In_575,In_0);
nand U1899 (N_1899,In_332,In_586);
and U1900 (N_1900,In_705,In_9);
nand U1901 (N_1901,In_724,In_964);
or U1902 (N_1902,In_325,In_92);
nand U1903 (N_1903,In_842,In_239);
or U1904 (N_1904,In_621,In_650);
nor U1905 (N_1905,In_727,In_974);
or U1906 (N_1906,In_413,In_253);
and U1907 (N_1907,In_810,In_314);
nor U1908 (N_1908,In_333,In_843);
nand U1909 (N_1909,In_171,In_606);
or U1910 (N_1910,In_182,In_243);
or U1911 (N_1911,In_711,In_584);
and U1912 (N_1912,In_262,In_329);
xnor U1913 (N_1913,In_882,In_865);
nand U1914 (N_1914,In_959,In_631);
nand U1915 (N_1915,In_882,In_523);
and U1916 (N_1916,In_588,In_281);
nor U1917 (N_1917,In_127,In_945);
nand U1918 (N_1918,In_668,In_129);
nor U1919 (N_1919,In_279,In_570);
nand U1920 (N_1920,In_73,In_872);
and U1921 (N_1921,In_916,In_821);
nor U1922 (N_1922,In_726,In_193);
nor U1923 (N_1923,In_115,In_856);
nor U1924 (N_1924,In_942,In_666);
and U1925 (N_1925,In_64,In_993);
or U1926 (N_1926,In_601,In_998);
nor U1927 (N_1927,In_869,In_809);
nor U1928 (N_1928,In_186,In_484);
nor U1929 (N_1929,In_857,In_247);
nand U1930 (N_1930,In_634,In_490);
xor U1931 (N_1931,In_537,In_308);
nand U1932 (N_1932,In_250,In_549);
nand U1933 (N_1933,In_588,In_274);
and U1934 (N_1934,In_754,In_367);
nand U1935 (N_1935,In_594,In_346);
or U1936 (N_1936,In_901,In_828);
nand U1937 (N_1937,In_931,In_642);
nor U1938 (N_1938,In_872,In_589);
nor U1939 (N_1939,In_548,In_24);
and U1940 (N_1940,In_840,In_646);
or U1941 (N_1941,In_937,In_782);
nand U1942 (N_1942,In_801,In_264);
or U1943 (N_1943,In_400,In_581);
xor U1944 (N_1944,In_237,In_921);
and U1945 (N_1945,In_149,In_462);
nand U1946 (N_1946,In_898,In_984);
nand U1947 (N_1947,In_953,In_270);
nand U1948 (N_1948,In_513,In_245);
and U1949 (N_1949,In_384,In_923);
and U1950 (N_1950,In_153,In_942);
and U1951 (N_1951,In_881,In_905);
and U1952 (N_1952,In_300,In_127);
nor U1953 (N_1953,In_988,In_27);
and U1954 (N_1954,In_613,In_687);
and U1955 (N_1955,In_515,In_425);
and U1956 (N_1956,In_197,In_337);
xor U1957 (N_1957,In_697,In_351);
nor U1958 (N_1958,In_181,In_508);
nand U1959 (N_1959,In_203,In_189);
and U1960 (N_1960,In_858,In_233);
or U1961 (N_1961,In_514,In_660);
and U1962 (N_1962,In_994,In_383);
xor U1963 (N_1963,In_892,In_78);
nor U1964 (N_1964,In_424,In_26);
nor U1965 (N_1965,In_227,In_737);
nor U1966 (N_1966,In_765,In_861);
and U1967 (N_1967,In_253,In_62);
nand U1968 (N_1968,In_415,In_600);
nand U1969 (N_1969,In_213,In_638);
and U1970 (N_1970,In_534,In_967);
and U1971 (N_1971,In_499,In_683);
nand U1972 (N_1972,In_369,In_880);
or U1973 (N_1973,In_317,In_987);
or U1974 (N_1974,In_306,In_416);
nor U1975 (N_1975,In_388,In_487);
and U1976 (N_1976,In_733,In_450);
and U1977 (N_1977,In_39,In_372);
nor U1978 (N_1978,In_785,In_1);
and U1979 (N_1979,In_392,In_887);
and U1980 (N_1980,In_810,In_848);
and U1981 (N_1981,In_847,In_707);
and U1982 (N_1982,In_339,In_15);
xor U1983 (N_1983,In_707,In_997);
nand U1984 (N_1984,In_813,In_84);
nor U1985 (N_1985,In_359,In_838);
nor U1986 (N_1986,In_272,In_973);
xnor U1987 (N_1987,In_462,In_515);
nand U1988 (N_1988,In_269,In_250);
or U1989 (N_1989,In_424,In_328);
nor U1990 (N_1990,In_383,In_70);
and U1991 (N_1991,In_539,In_531);
nor U1992 (N_1992,In_922,In_293);
xor U1993 (N_1993,In_286,In_480);
and U1994 (N_1994,In_731,In_363);
and U1995 (N_1995,In_403,In_50);
and U1996 (N_1996,In_735,In_501);
or U1997 (N_1997,In_809,In_55);
nor U1998 (N_1998,In_560,In_768);
nor U1999 (N_1999,In_701,In_966);
and U2000 (N_2000,N_1367,N_1762);
or U2001 (N_2001,N_632,N_1606);
xnor U2002 (N_2002,N_1843,N_1288);
xnor U2003 (N_2003,N_1764,N_1754);
nor U2004 (N_2004,N_194,N_806);
or U2005 (N_2005,N_214,N_746);
nand U2006 (N_2006,N_534,N_1516);
xnor U2007 (N_2007,N_441,N_6);
nor U2008 (N_2008,N_825,N_267);
nor U2009 (N_2009,N_1482,N_329);
nand U2010 (N_2010,N_1401,N_968);
nor U2011 (N_2011,N_1144,N_49);
or U2012 (N_2012,N_1410,N_203);
nor U2013 (N_2013,N_683,N_1308);
nor U2014 (N_2014,N_1155,N_409);
nor U2015 (N_2015,N_826,N_1396);
and U2016 (N_2016,N_1445,N_1848);
nand U2017 (N_2017,N_452,N_107);
or U2018 (N_2018,N_1858,N_708);
nor U2019 (N_2019,N_1815,N_1374);
and U2020 (N_2020,N_1122,N_1102);
nor U2021 (N_2021,N_1197,N_30);
nor U2022 (N_2022,N_1636,N_1924);
and U2023 (N_2023,N_323,N_741);
nand U2024 (N_2024,N_456,N_1560);
xor U2025 (N_2025,N_1439,N_1430);
nand U2026 (N_2026,N_927,N_1538);
nand U2027 (N_2027,N_1822,N_569);
or U2028 (N_2028,N_475,N_988);
nor U2029 (N_2029,N_1300,N_282);
and U2030 (N_2030,N_1025,N_1687);
nor U2031 (N_2031,N_258,N_778);
or U2032 (N_2032,N_419,N_1635);
and U2033 (N_2033,N_1472,N_1404);
or U2034 (N_2034,N_1906,N_1685);
xor U2035 (N_2035,N_748,N_706);
and U2036 (N_2036,N_1782,N_1909);
and U2037 (N_2037,N_223,N_1292);
nand U2038 (N_2038,N_805,N_1739);
nand U2039 (N_2039,N_1831,N_577);
xnor U2040 (N_2040,N_1798,N_410);
and U2041 (N_2041,N_400,N_813);
or U2042 (N_2042,N_909,N_1420);
and U2043 (N_2043,N_235,N_642);
and U2044 (N_2044,N_721,N_1012);
or U2045 (N_2045,N_1515,N_809);
nor U2046 (N_2046,N_336,N_870);
nor U2047 (N_2047,N_474,N_1281);
or U2048 (N_2048,N_956,N_690);
or U2049 (N_2049,N_60,N_1097);
or U2050 (N_2050,N_510,N_357);
or U2051 (N_2051,N_123,N_782);
or U2052 (N_2052,N_1605,N_566);
and U2053 (N_2053,N_627,N_1252);
nand U2054 (N_2054,N_1215,N_532);
or U2055 (N_2055,N_354,N_815);
nor U2056 (N_2056,N_148,N_159);
or U2057 (N_2057,N_662,N_1266);
nor U2058 (N_2058,N_1552,N_149);
and U2059 (N_2059,N_1674,N_747);
nor U2060 (N_2060,N_1403,N_919);
nor U2061 (N_2061,N_140,N_614);
nand U2062 (N_2062,N_1968,N_1640);
or U2063 (N_2063,N_346,N_1608);
nor U2064 (N_2064,N_508,N_402);
xor U2065 (N_2065,N_1612,N_433);
or U2066 (N_2066,N_78,N_1461);
and U2067 (N_2067,N_1573,N_1361);
nand U2068 (N_2068,N_1774,N_378);
or U2069 (N_2069,N_1956,N_177);
nand U2070 (N_2070,N_1167,N_91);
nor U2071 (N_2071,N_1239,N_687);
or U2072 (N_2072,N_290,N_602);
and U2073 (N_2073,N_596,N_1362);
nor U2074 (N_2074,N_1826,N_1448);
and U2075 (N_2075,N_1451,N_133);
and U2076 (N_2076,N_1898,N_1865);
and U2077 (N_2077,N_1223,N_1655);
and U2078 (N_2078,N_95,N_1354);
nand U2079 (N_2079,N_44,N_929);
and U2080 (N_2080,N_794,N_1489);
or U2081 (N_2081,N_920,N_786);
or U2082 (N_2082,N_166,N_1123);
xor U2083 (N_2083,N_617,N_857);
and U2084 (N_2084,N_57,N_976);
nor U2085 (N_2085,N_574,N_73);
nor U2086 (N_2086,N_1184,N_1153);
nor U2087 (N_2087,N_1305,N_1969);
or U2088 (N_2088,N_1264,N_1158);
nand U2089 (N_2089,N_442,N_603);
nand U2090 (N_2090,N_1648,N_657);
and U2091 (N_2091,N_545,N_1381);
nand U2092 (N_2092,N_29,N_1501);
or U2093 (N_2093,N_1991,N_685);
nand U2094 (N_2094,N_891,N_144);
and U2095 (N_2095,N_1716,N_397);
nor U2096 (N_2096,N_276,N_1022);
nand U2097 (N_2097,N_186,N_420);
and U2098 (N_2098,N_430,N_1806);
nand U2099 (N_2099,N_1047,N_62);
and U2100 (N_2100,N_1370,N_616);
and U2101 (N_2101,N_1033,N_1183);
nand U2102 (N_2102,N_444,N_306);
or U2103 (N_2103,N_496,N_878);
and U2104 (N_2104,N_833,N_608);
and U2105 (N_2105,N_1170,N_1690);
nand U2106 (N_2106,N_1205,N_549);
nand U2107 (N_2107,N_1903,N_155);
nand U2108 (N_2108,N_1103,N_1624);
nor U2109 (N_2109,N_190,N_607);
or U2110 (N_2110,N_831,N_1411);
nand U2111 (N_2111,N_218,N_379);
or U2112 (N_2112,N_983,N_1468);
and U2113 (N_2113,N_376,N_345);
or U2114 (N_2114,N_1057,N_1712);
xor U2115 (N_2115,N_1582,N_189);
nand U2116 (N_2116,N_1957,N_256);
or U2117 (N_2117,N_36,N_1455);
and U2118 (N_2118,N_1156,N_967);
and U2119 (N_2119,N_1632,N_331);
and U2120 (N_2120,N_1509,N_1176);
nand U2121 (N_2121,N_856,N_1457);
and U2122 (N_2122,N_307,N_269);
xnor U2123 (N_2123,N_246,N_471);
or U2124 (N_2124,N_658,N_160);
and U2125 (N_2125,N_1980,N_399);
nor U2126 (N_2126,N_1079,N_992);
xor U2127 (N_2127,N_362,N_1295);
nor U2128 (N_2128,N_1888,N_202);
xnor U2129 (N_2129,N_482,N_559);
or U2130 (N_2130,N_671,N_1916);
xor U2131 (N_2131,N_668,N_588);
and U2132 (N_2132,N_1673,N_1614);
nor U2133 (N_2133,N_1729,N_1793);
or U2134 (N_2134,N_1702,N_161);
nor U2135 (N_2135,N_743,N_460);
and U2136 (N_2136,N_908,N_277);
and U2137 (N_2137,N_1009,N_758);
nand U2138 (N_2138,N_1817,N_546);
and U2139 (N_2139,N_892,N_355);
or U2140 (N_2140,N_772,N_461);
or U2141 (N_2141,N_1778,N_1399);
nor U2142 (N_2142,N_75,N_1830);
and U2143 (N_2143,N_1050,N_1409);
nand U2144 (N_2144,N_1010,N_1091);
xor U2145 (N_2145,N_1100,N_1626);
xnor U2146 (N_2146,N_673,N_486);
nor U2147 (N_2147,N_1657,N_311);
or U2148 (N_2148,N_249,N_953);
or U2149 (N_2149,N_726,N_492);
and U2150 (N_2150,N_618,N_1602);
nor U2151 (N_2151,N_134,N_23);
nor U2152 (N_2152,N_15,N_1819);
nand U2153 (N_2153,N_684,N_1449);
nor U2154 (N_2154,N_9,N_936);
and U2155 (N_2155,N_1920,N_1678);
and U2156 (N_2156,N_1821,N_1355);
and U2157 (N_2157,N_1684,N_562);
nand U2158 (N_2158,N_1519,N_139);
nand U2159 (N_2159,N_1530,N_1611);
xnor U2160 (N_2160,N_1628,N_1023);
and U2161 (N_2161,N_639,N_1651);
nor U2162 (N_2162,N_780,N_1856);
and U2163 (N_2163,N_383,N_583);
nor U2164 (N_2164,N_1125,N_226);
or U2165 (N_2165,N_1915,N_1303);
and U2166 (N_2166,N_284,N_1928);
nand U2167 (N_2167,N_1026,N_1034);
nor U2168 (N_2168,N_917,N_429);
nand U2169 (N_2169,N_470,N_1485);
and U2170 (N_2170,N_1788,N_1293);
nor U2171 (N_2171,N_476,N_1595);
xor U2172 (N_2172,N_2,N_334);
and U2173 (N_2173,N_1376,N_1311);
nor U2174 (N_2174,N_434,N_1832);
nand U2175 (N_2175,N_1005,N_1593);
nand U2176 (N_2176,N_328,N_184);
or U2177 (N_2177,N_63,N_1761);
and U2178 (N_2178,N_453,N_1384);
and U2179 (N_2179,N_1201,N_222);
nand U2180 (N_2180,N_1571,N_972);
and U2181 (N_2181,N_1352,N_1564);
xor U2182 (N_2182,N_1203,N_915);
or U2183 (N_2183,N_1621,N_304);
or U2184 (N_2184,N_1836,N_1180);
and U2185 (N_2185,N_1524,N_1255);
nor U2186 (N_2186,N_1336,N_118);
nor U2187 (N_2187,N_1586,N_459);
or U2188 (N_2188,N_1443,N_1043);
and U2189 (N_2189,N_886,N_1109);
or U2190 (N_2190,N_1108,N_1488);
nor U2191 (N_2191,N_423,N_1329);
nor U2192 (N_2192,N_1795,N_1583);
nor U2193 (N_2193,N_787,N_1864);
nand U2194 (N_2194,N_146,N_655);
nor U2195 (N_2195,N_1507,N_1032);
and U2196 (N_2196,N_624,N_1060);
xnor U2197 (N_2197,N_1545,N_180);
nor U2198 (N_2198,N_941,N_1977);
xor U2199 (N_2199,N_1995,N_612);
xor U2200 (N_2200,N_1557,N_1174);
or U2201 (N_2201,N_1569,N_1412);
nor U2202 (N_2202,N_100,N_1610);
or U2203 (N_2203,N_1699,N_403);
nor U2204 (N_2204,N_414,N_197);
nor U2205 (N_2205,N_517,N_1900);
nor U2206 (N_2206,N_902,N_1724);
nand U2207 (N_2207,N_493,N_871);
and U2208 (N_2208,N_1017,N_255);
xor U2209 (N_2209,N_582,N_1850);
or U2210 (N_2210,N_1715,N_206);
and U2211 (N_2211,N_696,N_339);
and U2212 (N_2212,N_1555,N_1398);
nor U2213 (N_2213,N_1084,N_145);
xor U2214 (N_2214,N_827,N_1905);
nand U2215 (N_2215,N_1157,N_117);
or U2216 (N_2216,N_873,N_183);
and U2217 (N_2217,N_1578,N_46);
and U2218 (N_2218,N_436,N_1733);
and U2219 (N_2219,N_254,N_1659);
xor U2220 (N_2220,N_904,N_274);
xnor U2221 (N_2221,N_736,N_1750);
or U2222 (N_2222,N_1315,N_1853);
and U2223 (N_2223,N_1820,N_11);
and U2224 (N_2224,N_1475,N_1181);
xor U2225 (N_2225,N_1901,N_800);
nor U2226 (N_2226,N_1914,N_1723);
nand U2227 (N_2227,N_820,N_61);
nand U2228 (N_2228,N_1711,N_439);
and U2229 (N_2229,N_1378,N_1718);
nand U2230 (N_2230,N_1607,N_1946);
nor U2231 (N_2231,N_702,N_1868);
and U2232 (N_2232,N_1649,N_727);
and U2233 (N_2233,N_544,N_1707);
nor U2234 (N_2234,N_248,N_1587);
nand U2235 (N_2235,N_849,N_1664);
nor U2236 (N_2236,N_1114,N_1392);
nor U2237 (N_2237,N_413,N_1134);
nor U2238 (N_2238,N_1751,N_1139);
xor U2239 (N_2239,N_645,N_1693);
or U2240 (N_2240,N_1780,N_1141);
nand U2241 (N_2241,N_1280,N_765);
nor U2242 (N_2242,N_350,N_1747);
nand U2243 (N_2243,N_1600,N_205);
nand U2244 (N_2244,N_1497,N_1386);
nor U2245 (N_2245,N_1120,N_1414);
nor U2246 (N_2246,N_600,N_862);
or U2247 (N_2247,N_447,N_670);
nand U2248 (N_2248,N_554,N_1741);
nor U2249 (N_2249,N_384,N_636);
and U2250 (N_2250,N_349,N_543);
or U2251 (N_2251,N_1880,N_868);
xnor U2252 (N_2252,N_1435,N_259);
and U2253 (N_2253,N_744,N_335);
or U2254 (N_2254,N_1616,N_796);
or U2255 (N_2255,N_565,N_1537);
nand U2256 (N_2256,N_722,N_1302);
or U2257 (N_2257,N_1550,N_784);
xnor U2258 (N_2258,N_585,N_666);
and U2259 (N_2259,N_1558,N_1278);
nor U2260 (N_2260,N_1121,N_982);
nand U2261 (N_2261,N_279,N_253);
or U2262 (N_2262,N_652,N_922);
nand U2263 (N_2263,N_714,N_1510);
nand U2264 (N_2264,N_1163,N_1596);
and U2265 (N_2265,N_1147,N_1949);
nand U2266 (N_2266,N_392,N_1385);
and U2267 (N_2267,N_381,N_1979);
nor U2268 (N_2268,N_1294,N_74);
or U2269 (N_2269,N_1230,N_215);
nor U2270 (N_2270,N_1846,N_1382);
and U2271 (N_2271,N_960,N_1543);
or U2272 (N_2272,N_1040,N_188);
nand U2273 (N_2273,N_244,N_83);
xor U2274 (N_2274,N_1695,N_1907);
nor U2275 (N_2275,N_1471,N_1743);
xnor U2276 (N_2276,N_1663,N_387);
and U2277 (N_2277,N_753,N_28);
or U2278 (N_2278,N_1634,N_1881);
or U2279 (N_2279,N_701,N_834);
and U2280 (N_2280,N_1656,N_978);
or U2281 (N_2281,N_239,N_1938);
and U2282 (N_2282,N_321,N_1601);
xor U2283 (N_2283,N_1814,N_790);
nor U2284 (N_2284,N_1188,N_730);
or U2285 (N_2285,N_373,N_654);
nor U2286 (N_2286,N_1185,N_664);
nand U2287 (N_2287,N_1225,N_232);
and U2288 (N_2288,N_369,N_237);
nand U2289 (N_2289,N_360,N_1375);
nor U2290 (N_2290,N_70,N_513);
or U2291 (N_2291,N_219,N_1581);
xnor U2292 (N_2292,N_212,N_1683);
nand U2293 (N_2293,N_1958,N_1345);
or U2294 (N_2294,N_1087,N_47);
and U2295 (N_2295,N_1368,N_961);
nor U2296 (N_2296,N_405,N_332);
or U2297 (N_2297,N_681,N_644);
and U2298 (N_2298,N_1927,N_943);
and U2299 (N_2299,N_84,N_634);
or U2300 (N_2300,N_1000,N_1011);
nand U2301 (N_2301,N_1929,N_1923);
or U2302 (N_2302,N_693,N_71);
nor U2303 (N_2303,N_175,N_557);
nor U2304 (N_2304,N_368,N_754);
and U2305 (N_2305,N_1861,N_1740);
and U2306 (N_2306,N_224,N_342);
or U2307 (N_2307,N_720,N_599);
or U2308 (N_2308,N_1479,N_750);
nor U2309 (N_2309,N_1243,N_1776);
xnor U2310 (N_2310,N_380,N_1348);
xnor U2311 (N_2311,N_126,N_217);
nand U2312 (N_2312,N_1811,N_506);
nor U2313 (N_2313,N_1085,N_1356);
and U2314 (N_2314,N_337,N_1785);
or U2315 (N_2315,N_167,N_1459);
nor U2316 (N_2316,N_1823,N_1541);
nand U2317 (N_2317,N_1494,N_649);
and U2318 (N_2318,N_114,N_851);
xor U2319 (N_2319,N_17,N_1129);
and U2320 (N_2320,N_821,N_1737);
nor U2321 (N_2321,N_1997,N_1189);
or U2322 (N_2322,N_1146,N_814);
nand U2323 (N_2323,N_1941,N_1062);
nor U2324 (N_2324,N_1574,N_1682);
or U2325 (N_2325,N_556,N_1970);
nor U2326 (N_2326,N_1127,N_121);
or U2327 (N_2327,N_1708,N_85);
or U2328 (N_2328,N_1713,N_1604);
nand U2329 (N_2329,N_1705,N_725);
nor U2330 (N_2330,N_1879,N_287);
or U2331 (N_2331,N_90,N_310);
nor U2332 (N_2332,N_1646,N_299);
and U2333 (N_2333,N_1171,N_1887);
or U2334 (N_2334,N_1267,N_531);
nor U2335 (N_2335,N_1766,N_1234);
nor U2336 (N_2336,N_1789,N_1452);
nor U2337 (N_2337,N_1116,N_1990);
nor U2338 (N_2338,N_521,N_1554);
or U2339 (N_2339,N_467,N_12);
nand U2340 (N_2340,N_1745,N_643);
and U2341 (N_2341,N_789,N_1250);
or U2342 (N_2342,N_1787,N_391);
or U2343 (N_2343,N_1801,N_1769);
nor U2344 (N_2344,N_533,N_1758);
nor U2345 (N_2345,N_1742,N_152);
nand U2346 (N_2346,N_1617,N_1366);
or U2347 (N_2347,N_548,N_1502);
nand U2348 (N_2348,N_724,N_443);
nand U2349 (N_2349,N_1099,N_1372);
nor U2350 (N_2350,N_1306,N_358);
or U2351 (N_2351,N_1013,N_1512);
xor U2352 (N_2352,N_1478,N_942);
or U2353 (N_2353,N_1818,N_1453);
and U2354 (N_2354,N_385,N_1592);
nand U2355 (N_2355,N_1679,N_1505);
nor U2356 (N_2356,N_330,N_1442);
xnor U2357 (N_2357,N_382,N_1492);
or U2358 (N_2358,N_1508,N_209);
and U2359 (N_2359,N_515,N_717);
and U2360 (N_2360,N_56,N_704);
nand U2361 (N_2361,N_623,N_42);
or U2362 (N_2362,N_1466,N_1535);
or U2363 (N_2363,N_567,N_650);
or U2364 (N_2364,N_1481,N_903);
nand U2365 (N_2365,N_637,N_1187);
or U2366 (N_2366,N_1021,N_552);
xnor U2367 (N_2367,N_689,N_1642);
and U2368 (N_2368,N_1214,N_289);
or U2369 (N_2369,N_1248,N_247);
xor U2370 (N_2370,N_1987,N_739);
or U2371 (N_2371,N_1534,N_728);
nor U2372 (N_2372,N_930,N_1775);
nand U2373 (N_2373,N_1413,N_1698);
or U2374 (N_2374,N_1931,N_997);
and U2375 (N_2375,N_1397,N_265);
and U2376 (N_2376,N_1588,N_1897);
or U2377 (N_2377,N_1809,N_1473);
or U2378 (N_2378,N_1474,N_498);
nand U2379 (N_2379,N_1433,N_1018);
nand U2380 (N_2380,N_1661,N_1675);
nand U2381 (N_2381,N_322,N_1178);
nand U2382 (N_2382,N_1186,N_611);
nand U2383 (N_2383,N_783,N_1567);
or U2384 (N_2384,N_1719,N_966);
nand U2385 (N_2385,N_937,N_1283);
and U2386 (N_2386,N_416,N_1458);
or U2387 (N_2387,N_1867,N_415);
and U2388 (N_2388,N_575,N_847);
nand U2389 (N_2389,N_1738,N_846);
or U2390 (N_2390,N_1198,N_1316);
or U2391 (N_2391,N_905,N_1944);
and U2392 (N_2392,N_101,N_1553);
nor U2393 (N_2393,N_523,N_314);
nand U2394 (N_2394,N_1947,N_1173);
or U2395 (N_2395,N_449,N_170);
nand U2396 (N_2396,N_676,N_1427);
and U2397 (N_2397,N_1262,N_1067);
or U2398 (N_2398,N_1194,N_1111);
nor U2399 (N_2399,N_934,N_458);
and U2400 (N_2400,N_1734,N_987);
nand U2401 (N_2401,N_1273,N_1432);
nor U2402 (N_2402,N_1556,N_869);
or U2403 (N_2403,N_1589,N_715);
and U2404 (N_2404,N_1835,N_1299);
xnor U2405 (N_2405,N_1770,N_876);
or U2406 (N_2406,N_773,N_1531);
nand U2407 (N_2407,N_1598,N_1963);
or U2408 (N_2408,N_16,N_1562);
or U2409 (N_2409,N_45,N_1222);
xor U2410 (N_2410,N_1772,N_483);
and U2411 (N_2411,N_351,N_1086);
nand U2412 (N_2412,N_807,N_867);
or U2413 (N_2413,N_305,N_980);
or U2414 (N_2414,N_1756,N_386);
nor U2415 (N_2415,N_751,N_699);
xnor U2416 (N_2416,N_529,N_1644);
nor U2417 (N_2417,N_938,N_1996);
and U2418 (N_2418,N_396,N_1030);
and U2419 (N_2419,N_200,N_1862);
xnor U2420 (N_2420,N_1059,N_948);
or U2421 (N_2421,N_1387,N_418);
or U2422 (N_2422,N_480,N_1200);
nor U2423 (N_2423,N_791,N_984);
and U2424 (N_2424,N_1055,N_842);
or U2425 (N_2425,N_1975,N_1866);
nor U2426 (N_2426,N_64,N_1135);
and U2427 (N_2427,N_723,N_464);
and U2428 (N_2428,N_516,N_1726);
or U2429 (N_2429,N_425,N_312);
nor U2430 (N_2430,N_740,N_1837);
nor U2431 (N_2431,N_7,N_1042);
or U2432 (N_2432,N_113,N_479);
nand U2433 (N_2433,N_48,N_974);
nand U2434 (N_2434,N_77,N_950);
nor U2435 (N_2435,N_1454,N_1217);
nand U2436 (N_2436,N_1703,N_877);
and U2437 (N_2437,N_169,N_1480);
nor U2438 (N_2438,N_893,N_522);
and U2439 (N_2439,N_769,N_1104);
nand U2440 (N_2440,N_1575,N_1429);
and U2441 (N_2441,N_1694,N_989);
and U2442 (N_2442,N_1282,N_1256);
or U2443 (N_2443,N_367,N_1643);
or U2444 (N_2444,N_537,N_1549);
nand U2445 (N_2445,N_854,N_530);
nand U2446 (N_2446,N_1752,N_1343);
nor U2447 (N_2447,N_958,N_932);
nor U2448 (N_2448,N_1670,N_547);
or U2449 (N_2449,N_500,N_1686);
and U2450 (N_2450,N_865,N_1160);
nand U2451 (N_2451,N_1857,N_1730);
and U2452 (N_2452,N_977,N_1048);
and U2453 (N_2453,N_1195,N_1031);
xor U2454 (N_2454,N_949,N_1052);
xor U2455 (N_2455,N_1212,N_1523);
and U2456 (N_2456,N_1755,N_271);
nand U2457 (N_2457,N_263,N_315);
nor U2458 (N_2458,N_185,N_1464);
nand U2459 (N_2459,N_250,N_1999);
nor U2460 (N_2460,N_802,N_1204);
and U2461 (N_2461,N_946,N_1658);
nand U2462 (N_2462,N_1165,N_795);
xnor U2463 (N_2463,N_1072,N_120);
and U2464 (N_2464,N_1520,N_1419);
or U2465 (N_2465,N_707,N_275);
nand U2466 (N_2466,N_944,N_648);
nand U2467 (N_2467,N_288,N_211);
and U2468 (N_2468,N_885,N_1800);
or U2469 (N_2469,N_1889,N_1090);
and U2470 (N_2470,N_76,N_27);
and U2471 (N_2471,N_931,N_1838);
or U2472 (N_2472,N_526,N_626);
and U2473 (N_2473,N_1051,N_1095);
nor U2474 (N_2474,N_686,N_918);
nor U2475 (N_2475,N_1622,N_1877);
nor U2476 (N_2476,N_1808,N_88);
and U2477 (N_2477,N_996,N_604);
and U2478 (N_2478,N_551,N_438);
nor U2479 (N_2479,N_38,N_127);
or U2480 (N_2480,N_1312,N_1006);
and U2481 (N_2481,N_656,N_1007);
or U2482 (N_2482,N_435,N_1077);
or U2483 (N_2483,N_238,N_124);
nand U2484 (N_2484,N_1563,N_66);
xnor U2485 (N_2485,N_220,N_1532);
or U2486 (N_2486,N_1105,N_1117);
xor U2487 (N_2487,N_1681,N_595);
nand U2488 (N_2488,N_50,N_804);
and U2489 (N_2489,N_1263,N_1493);
nand U2490 (N_2490,N_573,N_1882);
nand U2491 (N_2491,N_864,N_641);
or U2492 (N_2492,N_1191,N_1771);
nand U2493 (N_2493,N_1620,N_674);
or U2494 (N_2494,N_182,N_103);
nand U2495 (N_2495,N_233,N_1922);
or U2496 (N_2496,N_1717,N_1842);
nor U2497 (N_2497,N_561,N_1894);
nor U2498 (N_2498,N_1318,N_347);
or U2499 (N_2499,N_1962,N_1744);
or U2500 (N_2500,N_1169,N_875);
nand U2501 (N_2501,N_756,N_1498);
nand U2502 (N_2502,N_41,N_964);
and U2503 (N_2503,N_1319,N_866);
nand U2504 (N_2504,N_1691,N_1101);
nor U2505 (N_2505,N_25,N_581);
nor U2506 (N_2506,N_733,N_503);
nand U2507 (N_2507,N_35,N_1229);
nor U2508 (N_2508,N_261,N_1346);
nor U2509 (N_2509,N_19,N_951);
nand U2510 (N_2510,N_793,N_620);
xnor U2511 (N_2511,N_981,N_990);
and U2512 (N_2512,N_1335,N_799);
nor U2513 (N_2513,N_1015,N_906);
and U2514 (N_2514,N_757,N_1383);
or U2515 (N_2515,N_466,N_1297);
or U2516 (N_2516,N_504,N_995);
nor U2517 (N_2517,N_1049,N_1511);
nand U2518 (N_2518,N_518,N_1314);
nand U2519 (N_2519,N_1008,N_1089);
nor U2520 (N_2520,N_659,N_116);
and U2521 (N_2521,N_1525,N_1393);
nand U2522 (N_2522,N_297,N_268);
nand U2523 (N_2523,N_72,N_525);
nand U2524 (N_2524,N_1613,N_431);
or U2525 (N_2525,N_640,N_1504);
nor U2526 (N_2526,N_558,N_729);
and U2527 (N_2527,N_234,N_859);
nor U2528 (N_2528,N_1885,N_1344);
and U2529 (N_2529,N_841,N_1065);
nand U2530 (N_2530,N_1797,N_213);
and U2531 (N_2531,N_1910,N_779);
nor U2532 (N_2532,N_363,N_1166);
xor U2533 (N_2533,N_171,N_499);
nor U2534 (N_2534,N_1580,N_1112);
nand U2535 (N_2535,N_1773,N_147);
and U2536 (N_2536,N_755,N_317);
or U2537 (N_2537,N_352,N_375);
and U2538 (N_2538,N_852,N_925);
or U2539 (N_2539,N_1896,N_286);
or U2540 (N_2540,N_718,N_1175);
or U2541 (N_2541,N_294,N_1330);
xor U2542 (N_2542,N_1279,N_571);
and U2543 (N_2543,N_1063,N_1839);
nand U2544 (N_2544,N_1965,N_1365);
nor U2545 (N_2545,N_1037,N_539);
and U2546 (N_2546,N_774,N_462);
nand U2547 (N_2547,N_1447,N_1886);
nor U2548 (N_2548,N_1075,N_1542);
nor U2549 (N_2549,N_1937,N_450);
and U2550 (N_2550,N_933,N_1873);
nand U2551 (N_2551,N_1207,N_1572);
nor U2552 (N_2552,N_863,N_251);
nand U2553 (N_2553,N_1746,N_10);
nor U2554 (N_2554,N_973,N_1003);
or U2555 (N_2555,N_564,N_164);
nand U2556 (N_2556,N_481,N_485);
or U2557 (N_2557,N_1662,N_625);
nor U2558 (N_2558,N_1465,N_1310);
nand U2559 (N_2559,N_1389,N_240);
nand U2560 (N_2560,N_344,N_965);
and U2561 (N_2561,N_395,N_389);
xnor U2562 (N_2562,N_1218,N_80);
or U2563 (N_2563,N_1076,N_1945);
and U2564 (N_2564,N_1014,N_828);
or U2565 (N_2565,N_536,N_850);
or U2566 (N_2566,N_55,N_911);
and U2567 (N_2567,N_1805,N_1342);
nor U2568 (N_2568,N_594,N_1470);
and U2569 (N_2569,N_731,N_1487);
or U2570 (N_2570,N_463,N_572);
or U2571 (N_2571,N_1148,N_491);
and U2572 (N_2572,N_291,N_125);
nor U2573 (N_2573,N_563,N_33);
and U2574 (N_2574,N_1847,N_1757);
or U2575 (N_2575,N_1841,N_1298);
nor U2576 (N_2576,N_162,N_132);
xor U2577 (N_2577,N_1441,N_92);
xnor U2578 (N_2578,N_440,N_1599);
nor U2579 (N_2579,N_93,N_1477);
nor U2580 (N_2580,N_698,N_176);
and U2581 (N_2581,N_1667,N_1036);
and U2582 (N_2582,N_609,N_1669);
or U2583 (N_2583,N_762,N_192);
and U2584 (N_2584,N_1988,N_678);
xor U2585 (N_2585,N_1869,N_1113);
or U2586 (N_2586,N_1093,N_1016);
nor U2587 (N_2587,N_660,N_894);
or U2588 (N_2588,N_1145,N_954);
nor U2589 (N_2589,N_1619,N_1467);
or U2590 (N_2590,N_528,N_1235);
nor U2591 (N_2591,N_1164,N_1456);
nor U2592 (N_2592,N_1136,N_998);
nor U2593 (N_2593,N_1638,N_129);
and U2594 (N_2594,N_1307,N_1400);
nand U2595 (N_2595,N_79,N_204);
or U2596 (N_2596,N_1998,N_427);
nor U2597 (N_2597,N_822,N_1227);
xnor U2598 (N_2598,N_1138,N_488);
nor U2599 (N_2599,N_1001,N_411);
nor U2600 (N_2600,N_1641,N_494);
nand U2601 (N_2601,N_901,N_1096);
nand U2602 (N_2602,N_1211,N_1486);
or U2603 (N_2603,N_1221,N_1921);
xnor U2604 (N_2604,N_1182,N_18);
nand U2605 (N_2605,N_1871,N_1024);
nand U2606 (N_2606,N_1506,N_1749);
nor U2607 (N_2607,N_1816,N_1844);
nor U2608 (N_2608,N_1660,N_1926);
xnor U2609 (N_2609,N_1296,N_59);
nor U2610 (N_2610,N_1834,N_764);
nor U2611 (N_2611,N_32,N_712);
or U2612 (N_2612,N_1630,N_1259);
or U2613 (N_2613,N_1625,N_1154);
nand U2614 (N_2614,N_1631,N_1973);
xnor U2615 (N_2615,N_1251,N_67);
nand U2616 (N_2616,N_1417,N_1199);
and U2617 (N_2617,N_719,N_1275);
nand U2618 (N_2618,N_1978,N_501);
nand U2619 (N_2619,N_1561,N_1364);
or U2620 (N_2620,N_775,N_1106);
xnor U2621 (N_2621,N_986,N_131);
nor U2622 (N_2622,N_1483,N_1484);
and U2623 (N_2623,N_1518,N_1615);
and U2624 (N_2624,N_231,N_1540);
or U2625 (N_2625,N_576,N_888);
nor U2626 (N_2626,N_1943,N_601);
or U2627 (N_2627,N_880,N_1426);
nand U2628 (N_2628,N_1781,N_1045);
nand U2629 (N_2629,N_1349,N_1904);
and U2630 (N_2630,N_1168,N_165);
nand U2631 (N_2631,N_316,N_792);
xnor U2632 (N_2632,N_1064,N_605);
nor U2633 (N_2633,N_553,N_406);
or U2634 (N_2634,N_1993,N_808);
nor U2635 (N_2635,N_1233,N_104);
and U2636 (N_2636,N_1246,N_1513);
xnor U2637 (N_2637,N_763,N_540);
or U2638 (N_2638,N_811,N_1895);
nand U2639 (N_2639,N_1891,N_1238);
and U2640 (N_2640,N_1035,N_1402);
and U2641 (N_2641,N_1380,N_1849);
nor U2642 (N_2642,N_454,N_1131);
nor U2643 (N_2643,N_1727,N_398);
nor U2644 (N_2644,N_1056,N_622);
xor U2645 (N_2645,N_1829,N_1313);
nand U2646 (N_2646,N_697,N_1714);
nor U2647 (N_2647,N_1359,N_1078);
nor U2648 (N_2648,N_1992,N_207);
nor U2649 (N_2649,N_445,N_1132);
or U2650 (N_2650,N_58,N_5);
nor U2651 (N_2651,N_1768,N_1875);
nor U2652 (N_2652,N_884,N_325);
nand U2653 (N_2653,N_816,N_560);
nor U2654 (N_2654,N_1653,N_122);
and U2655 (N_2655,N_1870,N_446);
nand U2656 (N_2656,N_333,N_318);
or U2657 (N_2657,N_1786,N_1377);
nand U2658 (N_2658,N_108,N_1363);
and U2659 (N_2659,N_1824,N_874);
nand U2660 (N_2660,N_705,N_1753);
or U2661 (N_2661,N_343,N_1254);
and U2662 (N_2662,N_710,N_327);
nor U2663 (N_2663,N_797,N_1088);
nand U2664 (N_2664,N_677,N_1124);
and U2665 (N_2665,N_830,N_1514);
or U2666 (N_2666,N_136,N_798);
and U2667 (N_2667,N_579,N_1731);
xor U2668 (N_2668,N_3,N_1236);
or U2669 (N_2669,N_777,N_421);
nand U2670 (N_2670,N_487,N_1286);
or U2671 (N_2671,N_109,N_975);
or U2672 (N_2672,N_1416,N_1645);
nor U2673 (N_2673,N_1369,N_691);
or U2674 (N_2674,N_1765,N_86);
nor U2675 (N_2675,N_994,N_1942);
nor U2676 (N_2676,N_613,N_128);
or U2677 (N_2677,N_228,N_1917);
or U2678 (N_2678,N_102,N_422);
or U2679 (N_2679,N_1902,N_1701);
or U2680 (N_2680,N_1568,N_1807);
and U2681 (N_2681,N_667,N_555);
and U2682 (N_2682,N_1245,N_1083);
xnor U2683 (N_2683,N_914,N_53);
or U2684 (N_2684,N_635,N_1434);
and U2685 (N_2685,N_1650,N_262);
and U2686 (N_2686,N_1799,N_1276);
and U2687 (N_2687,N_1274,N_631);
xnor U2688 (N_2688,N_497,N_26);
and U2689 (N_2689,N_1597,N_1536);
nand U2690 (N_2690,N_1812,N_1019);
or U2691 (N_2691,N_1721,N_1982);
nand U2692 (N_2692,N_1038,N_663);
nand U2693 (N_2693,N_65,N_348);
nor U2694 (N_2694,N_907,N_591);
nor U2695 (N_2695,N_887,N_1883);
nor U2696 (N_2696,N_1517,N_1428);
nor U2697 (N_2697,N_340,N_285);
or U2698 (N_2698,N_22,N_1317);
or U2699 (N_2699,N_511,N_1119);
and U2700 (N_2700,N_653,N_883);
nand U2701 (N_2701,N_947,N_143);
nor U2702 (N_2702,N_970,N_1859);
xor U2703 (N_2703,N_836,N_292);
and U2704 (N_2704,N_178,N_1845);
or U2705 (N_2705,N_87,N_1950);
nand U2706 (N_2706,N_1825,N_1046);
nor U2707 (N_2707,N_138,N_1618);
and U2708 (N_2708,N_1689,N_1028);
nor U2709 (N_2709,N_230,N_1258);
nor U2710 (N_2710,N_858,N_1341);
nand U2711 (N_2711,N_1964,N_848);
xnor U2712 (N_2712,N_437,N_82);
and U2713 (N_2713,N_1271,N_570);
nand U2714 (N_2714,N_1725,N_319);
or U2715 (N_2715,N_1784,N_527);
or U2716 (N_2716,N_243,N_1224);
xnor U2717 (N_2717,N_835,N_818);
nor U2718 (N_2718,N_195,N_1490);
nand U2719 (N_2719,N_1340,N_1668);
or U2720 (N_2720,N_8,N_1261);
or U2721 (N_2721,N_1130,N_156);
or U2722 (N_2722,N_952,N_1706);
and U2723 (N_2723,N_1436,N_955);
or U2724 (N_2724,N_1529,N_817);
xnor U2725 (N_2725,N_1955,N_1763);
nor U2726 (N_2726,N_1732,N_1469);
and U2727 (N_2727,N_621,N_308);
or U2728 (N_2728,N_1952,N_1637);
and U2729 (N_2729,N_1810,N_519);
and U2730 (N_2730,N_1268,N_1863);
nand U2731 (N_2731,N_408,N_732);
or U2732 (N_2732,N_1081,N_1357);
nand U2733 (N_2733,N_1424,N_926);
or U2734 (N_2734,N_1700,N_1347);
nand U2735 (N_2735,N_300,N_241);
nand U2736 (N_2736,N_1908,N_1395);
and U2737 (N_2737,N_638,N_1860);
nor U2738 (N_2738,N_860,N_473);
nand U2739 (N_2739,N_1672,N_1591);
or U2740 (N_2740,N_1804,N_374);
and U2741 (N_2741,N_1939,N_1566);
nor U2742 (N_2742,N_252,N_1333);
nor U2743 (N_2743,N_771,N_1351);
and U2744 (N_2744,N_1783,N_1985);
nor U2745 (N_2745,N_1720,N_338);
nand U2746 (N_2746,N_1803,N_1463);
or U2747 (N_2747,N_130,N_1688);
xor U2748 (N_2748,N_844,N_606);
nor U2749 (N_2749,N_945,N_1321);
or U2750 (N_2750,N_507,N_1584);
nor U2751 (N_2751,N_302,N_54);
and U2752 (N_2752,N_150,N_838);
and U2753 (N_2753,N_1704,N_1110);
nand U2754 (N_2754,N_1893,N_1603);
nor U2755 (N_2755,N_1406,N_1149);
nand U2756 (N_2756,N_1226,N_840);
or U2757 (N_2757,N_1020,N_619);
nand U2758 (N_2758,N_912,N_524);
nand U2759 (N_2759,N_959,N_309);
nor U2760 (N_2760,N_455,N_1912);
xnor U2761 (N_2761,N_1967,N_1665);
or U2762 (N_2762,N_153,N_1876);
or U2763 (N_2763,N_361,N_13);
nor U2764 (N_2764,N_264,N_1633);
nand U2765 (N_2765,N_1760,N_1546);
nand U2766 (N_2766,N_97,N_520);
and U2767 (N_2767,N_1647,N_734);
and U2768 (N_2768,N_1337,N_110);
nand U2769 (N_2769,N_1966,N_1976);
nand U2770 (N_2770,N_760,N_69);
or U2771 (N_2771,N_1986,N_1373);
or U2772 (N_2772,N_21,N_1981);
and U2773 (N_2773,N_1654,N_1162);
and U2774 (N_2774,N_4,N_266);
nand U2775 (N_2775,N_713,N_1231);
or U2776 (N_2776,N_417,N_812);
xor U2777 (N_2777,N_580,N_1209);
nand U2778 (N_2778,N_759,N_1759);
nand U2779 (N_2779,N_1247,N_1551);
and U2780 (N_2780,N_320,N_1462);
and U2781 (N_2781,N_372,N_81);
nand U2782 (N_2782,N_1709,N_281);
xnor U2783 (N_2783,N_1159,N_939);
nand U2784 (N_2784,N_749,N_225);
and U2785 (N_2785,N_590,N_985);
nand U2786 (N_2786,N_1192,N_770);
or U2787 (N_2787,N_1450,N_776);
nand U2788 (N_2788,N_1802,N_1069);
nand U2789 (N_2789,N_141,N_1629);
and U2790 (N_2790,N_709,N_1527);
or U2791 (N_2791,N_928,N_688);
nor U2792 (N_2792,N_301,N_924);
nor U2793 (N_2793,N_694,N_633);
or U2794 (N_2794,N_628,N_1972);
xor U2795 (N_2795,N_897,N_514);
nand U2796 (N_2796,N_236,N_829);
nand U2797 (N_2797,N_1521,N_1228);
and U2798 (N_2798,N_1671,N_1107);
and U2799 (N_2799,N_1140,N_1394);
or U2800 (N_2800,N_1379,N_1577);
nor U2801 (N_2801,N_1852,N_1098);
or U2802 (N_2802,N_432,N_682);
or U2803 (N_2803,N_1405,N_1440);
nand U2804 (N_2804,N_923,N_767);
nor U2805 (N_2805,N_168,N_711);
nand U2806 (N_2806,N_1444,N_158);
nand U2807 (N_2807,N_505,N_969);
or U2808 (N_2808,N_598,N_1935);
nand U2809 (N_2809,N_1202,N_1027);
and U2810 (N_2810,N_1994,N_1270);
nor U2811 (N_2811,N_1533,N_535);
xnor U2812 (N_2812,N_1548,N_1940);
nand U2813 (N_2813,N_1918,N_163);
and U2814 (N_2814,N_889,N_963);
or U2815 (N_2815,N_1044,N_1039);
and U2816 (N_2816,N_1080,N_651);
or U2817 (N_2817,N_1495,N_999);
or U2818 (N_2818,N_1152,N_1179);
nand U2819 (N_2819,N_1196,N_752);
and U2820 (N_2820,N_1913,N_819);
nor U2821 (N_2821,N_448,N_1748);
or U2822 (N_2822,N_629,N_1539);
and U2823 (N_2823,N_1265,N_669);
or U2824 (N_2824,N_910,N_472);
nand U2825 (N_2825,N_502,N_1639);
xor U2826 (N_2826,N_89,N_587);
xor U2827 (N_2827,N_1041,N_1220);
nor U2828 (N_2828,N_1137,N_1899);
or U2829 (N_2829,N_1415,N_68);
nand U2830 (N_2830,N_1260,N_1094);
or U2831 (N_2831,N_801,N_1813);
or U2832 (N_2832,N_1325,N_1422);
or U2833 (N_2833,N_940,N_364);
xor U2834 (N_2834,N_1974,N_1796);
nor U2835 (N_2835,N_1073,N_881);
nand U2836 (N_2836,N_1331,N_993);
or U2837 (N_2837,N_823,N_1161);
and U2838 (N_2838,N_353,N_1590);
or U2839 (N_2839,N_584,N_359);
and U2840 (N_2840,N_489,N_1054);
and U2841 (N_2841,N_1332,N_1503);
nand U2842 (N_2842,N_1358,N_845);
nor U2843 (N_2843,N_393,N_99);
nor U2844 (N_2844,N_181,N_916);
xor U2845 (N_2845,N_401,N_921);
and U2846 (N_2846,N_1948,N_119);
xnor U2847 (N_2847,N_356,N_115);
nand U2848 (N_2848,N_1425,N_1237);
nor U2849 (N_2849,N_0,N_1071);
and U2850 (N_2850,N_221,N_1219);
and U2851 (N_2851,N_1058,N_703);
or U2852 (N_2852,N_1269,N_957);
and U2853 (N_2853,N_1792,N_1623);
xnor U2854 (N_2854,N_1884,N_1118);
or U2855 (N_2855,N_210,N_1827);
or U2856 (N_2856,N_1208,N_151);
or U2857 (N_2857,N_278,N_1984);
or U2858 (N_2858,N_495,N_1890);
or U2859 (N_2859,N_1971,N_593);
and U2860 (N_2860,N_1253,N_366);
or U2861 (N_2861,N_280,N_173);
nand U2862 (N_2862,N_568,N_1143);
xnor U2863 (N_2863,N_198,N_370);
or U2864 (N_2864,N_647,N_201);
xor U2865 (N_2865,N_270,N_550);
or U2866 (N_2866,N_890,N_1115);
or U2867 (N_2867,N_1241,N_738);
or U2868 (N_2868,N_1526,N_1959);
nor U2869 (N_2869,N_1326,N_20);
nand U2870 (N_2870,N_187,N_646);
nor U2871 (N_2871,N_37,N_1559);
nor U2872 (N_2872,N_853,N_227);
nor U2873 (N_2873,N_839,N_1840);
or U2874 (N_2874,N_900,N_1585);
or U2875 (N_2875,N_1068,N_1092);
or U2876 (N_2876,N_592,N_1855);
and U2877 (N_2877,N_672,N_326);
nand U2878 (N_2878,N_742,N_761);
and U2879 (N_2879,N_1878,N_1833);
and U2880 (N_2880,N_457,N_1431);
and U2881 (N_2881,N_1954,N_1);
and U2882 (N_2882,N_1579,N_1053);
or U2883 (N_2883,N_1082,N_468);
and U2884 (N_2884,N_979,N_1960);
or U2885 (N_2885,N_1418,N_43);
nor U2886 (N_2886,N_1932,N_191);
xnor U2887 (N_2887,N_1277,N_196);
nand U2888 (N_2888,N_451,N_1609);
or U2889 (N_2889,N_1677,N_1476);
and U2890 (N_2890,N_1460,N_1338);
nand U2891 (N_2891,N_245,N_94);
or U2892 (N_2892,N_855,N_154);
or U2893 (N_2893,N_1722,N_1301);
nand U2894 (N_2894,N_1323,N_1522);
nor U2895 (N_2895,N_1126,N_578);
and U2896 (N_2896,N_843,N_1828);
or U2897 (N_2897,N_1133,N_179);
and U2898 (N_2898,N_1289,N_1874);
nand U2899 (N_2899,N_296,N_465);
or U2900 (N_2900,N_1790,N_509);
nor U2901 (N_2901,N_1290,N_1528);
or U2902 (N_2902,N_1791,N_1350);
and U2903 (N_2903,N_1029,N_512);
nor U2904 (N_2904,N_1547,N_1360);
nor U2905 (N_2905,N_962,N_1491);
xnor U2906 (N_2906,N_469,N_216);
nand U2907 (N_2907,N_1735,N_260);
xor U2908 (N_2908,N_1892,N_1172);
or U2909 (N_2909,N_781,N_1213);
and U2910 (N_2910,N_879,N_1794);
or U2911 (N_2911,N_1696,N_1232);
nor U2912 (N_2912,N_538,N_1257);
nor U2913 (N_2913,N_1151,N_737);
xnor U2914 (N_2914,N_1371,N_680);
or U2915 (N_2915,N_283,N_766);
nor U2916 (N_2916,N_394,N_1594);
nor U2917 (N_2917,N_1438,N_1309);
and U2918 (N_2918,N_257,N_1983);
xor U2919 (N_2919,N_40,N_412);
nand U2920 (N_2920,N_1499,N_1951);
or U2921 (N_2921,N_1767,N_1576);
nand U2922 (N_2922,N_1339,N_1961);
nand U2923 (N_2923,N_1933,N_1322);
and U2924 (N_2924,N_788,N_229);
nor U2925 (N_2925,N_1002,N_1652);
nor U2926 (N_2926,N_1206,N_735);
nor U2927 (N_2927,N_695,N_1728);
nand U2928 (N_2928,N_872,N_407);
nand U2929 (N_2929,N_1930,N_1779);
and U2930 (N_2930,N_478,N_586);
or U2931 (N_2931,N_1074,N_541);
and U2932 (N_2932,N_193,N_1190);
nor U2933 (N_2933,N_424,N_199);
nor U2934 (N_2934,N_785,N_174);
nand U2935 (N_2935,N_589,N_768);
nor U2936 (N_2936,N_208,N_1710);
nand U2937 (N_2937,N_135,N_1421);
nor U2938 (N_2938,N_1066,N_1249);
or U2939 (N_2939,N_991,N_1242);
or U2940 (N_2940,N_837,N_1320);
or U2941 (N_2941,N_1150,N_39);
xnor U2942 (N_2942,N_1284,N_896);
xnor U2943 (N_2943,N_1388,N_1697);
or U2944 (N_2944,N_1070,N_630);
nand U2945 (N_2945,N_615,N_1570);
nand U2946 (N_2946,N_112,N_388);
nor U2947 (N_2947,N_371,N_913);
nor U2948 (N_2948,N_1911,N_810);
or U2949 (N_2949,N_242,N_1872);
nand U2950 (N_2950,N_1272,N_1953);
xnor U2951 (N_2951,N_1177,N_610);
xor U2952 (N_2952,N_824,N_1544);
nor U2953 (N_2953,N_679,N_1142);
nor U2954 (N_2954,N_157,N_428);
nor U2955 (N_2955,N_324,N_898);
nand U2956 (N_2956,N_1936,N_1240);
nor U2957 (N_2957,N_1692,N_96);
or U2958 (N_2958,N_1328,N_832);
or U2959 (N_2959,N_390,N_1736);
or U2960 (N_2960,N_1500,N_1210);
or U2961 (N_2961,N_1004,N_700);
nor U2962 (N_2962,N_661,N_1353);
or U2963 (N_2963,N_273,N_404);
nand U2964 (N_2964,N_861,N_803);
nor U2965 (N_2965,N_597,N_675);
xnor U2966 (N_2966,N_1128,N_1565);
and U2967 (N_2967,N_137,N_1408);
and U2968 (N_2968,N_1390,N_105);
nor U2969 (N_2969,N_1304,N_1989);
nor U2970 (N_2970,N_1407,N_1925);
or U2971 (N_2971,N_484,N_1437);
and U2972 (N_2972,N_365,N_899);
nor U2973 (N_2973,N_14,N_142);
nor U2974 (N_2974,N_477,N_1680);
xnor U2975 (N_2975,N_895,N_313);
and U2976 (N_2976,N_1777,N_745);
and U2977 (N_2977,N_1423,N_98);
and U2978 (N_2978,N_426,N_1334);
nor U2979 (N_2979,N_272,N_542);
or U2980 (N_2980,N_1327,N_1919);
xor U2981 (N_2981,N_111,N_1324);
and U2982 (N_2982,N_1216,N_882);
and U2983 (N_2983,N_1666,N_298);
and U2984 (N_2984,N_1193,N_341);
or U2985 (N_2985,N_172,N_490);
xnor U2986 (N_2986,N_106,N_1391);
or U2987 (N_2987,N_1854,N_31);
and U2988 (N_2988,N_1934,N_295);
and U2989 (N_2989,N_51,N_24);
or U2990 (N_2990,N_1285,N_692);
or U2991 (N_2991,N_1851,N_1446);
and U2992 (N_2992,N_971,N_1287);
and U2993 (N_2993,N_1061,N_935);
or U2994 (N_2994,N_716,N_303);
xnor U2995 (N_2995,N_1627,N_293);
or U2996 (N_2996,N_1496,N_665);
and U2997 (N_2997,N_1244,N_1291);
nand U2998 (N_2998,N_377,N_52);
nor U2999 (N_2999,N_1676,N_34);
and U3000 (N_3000,N_754,N_957);
and U3001 (N_3001,N_997,N_1956);
or U3002 (N_3002,N_1453,N_433);
nand U3003 (N_3003,N_38,N_1598);
and U3004 (N_3004,N_1804,N_709);
and U3005 (N_3005,N_1548,N_1129);
xor U3006 (N_3006,N_1826,N_1582);
nand U3007 (N_3007,N_911,N_577);
nor U3008 (N_3008,N_1698,N_1974);
nand U3009 (N_3009,N_1236,N_1020);
nor U3010 (N_3010,N_1887,N_724);
xor U3011 (N_3011,N_1744,N_1882);
and U3012 (N_3012,N_978,N_1595);
nor U3013 (N_3013,N_871,N_1006);
nor U3014 (N_3014,N_326,N_1270);
xor U3015 (N_3015,N_1771,N_1809);
or U3016 (N_3016,N_865,N_1912);
and U3017 (N_3017,N_1489,N_483);
or U3018 (N_3018,N_1694,N_427);
xor U3019 (N_3019,N_480,N_1669);
nor U3020 (N_3020,N_340,N_94);
nand U3021 (N_3021,N_325,N_335);
and U3022 (N_3022,N_1097,N_1161);
and U3023 (N_3023,N_742,N_763);
xnor U3024 (N_3024,N_601,N_1532);
or U3025 (N_3025,N_1603,N_334);
or U3026 (N_3026,N_1494,N_1009);
nand U3027 (N_3027,N_231,N_1811);
and U3028 (N_3028,N_352,N_1734);
and U3029 (N_3029,N_1322,N_33);
or U3030 (N_3030,N_573,N_1051);
or U3031 (N_3031,N_338,N_1844);
nor U3032 (N_3032,N_301,N_1725);
and U3033 (N_3033,N_1948,N_1458);
and U3034 (N_3034,N_23,N_1707);
or U3035 (N_3035,N_1933,N_700);
nand U3036 (N_3036,N_350,N_242);
nand U3037 (N_3037,N_1346,N_1133);
or U3038 (N_3038,N_982,N_1469);
or U3039 (N_3039,N_520,N_60);
or U3040 (N_3040,N_782,N_1754);
or U3041 (N_3041,N_618,N_1592);
nor U3042 (N_3042,N_1455,N_1298);
nor U3043 (N_3043,N_366,N_359);
or U3044 (N_3044,N_586,N_144);
nand U3045 (N_3045,N_1323,N_307);
nand U3046 (N_3046,N_757,N_60);
or U3047 (N_3047,N_550,N_1312);
nand U3048 (N_3048,N_52,N_1199);
or U3049 (N_3049,N_550,N_815);
and U3050 (N_3050,N_698,N_612);
or U3051 (N_3051,N_1512,N_237);
and U3052 (N_3052,N_421,N_295);
xor U3053 (N_3053,N_36,N_1068);
nand U3054 (N_3054,N_1557,N_1257);
xor U3055 (N_3055,N_896,N_614);
nand U3056 (N_3056,N_882,N_254);
or U3057 (N_3057,N_571,N_1925);
or U3058 (N_3058,N_784,N_653);
or U3059 (N_3059,N_1475,N_513);
and U3060 (N_3060,N_279,N_679);
nand U3061 (N_3061,N_139,N_1928);
xnor U3062 (N_3062,N_1202,N_1581);
nor U3063 (N_3063,N_1010,N_1051);
nor U3064 (N_3064,N_40,N_1362);
xnor U3065 (N_3065,N_1429,N_1372);
or U3066 (N_3066,N_1456,N_1436);
and U3067 (N_3067,N_859,N_791);
and U3068 (N_3068,N_642,N_280);
nand U3069 (N_3069,N_1968,N_916);
nand U3070 (N_3070,N_647,N_278);
nand U3071 (N_3071,N_493,N_460);
nand U3072 (N_3072,N_1979,N_891);
or U3073 (N_3073,N_1012,N_1904);
and U3074 (N_3074,N_153,N_627);
nor U3075 (N_3075,N_1042,N_1076);
and U3076 (N_3076,N_950,N_387);
and U3077 (N_3077,N_890,N_814);
nand U3078 (N_3078,N_1401,N_722);
and U3079 (N_3079,N_1243,N_783);
or U3080 (N_3080,N_1203,N_1577);
or U3081 (N_3081,N_376,N_1363);
nand U3082 (N_3082,N_1999,N_18);
nor U3083 (N_3083,N_263,N_1097);
and U3084 (N_3084,N_1165,N_1985);
xor U3085 (N_3085,N_1109,N_573);
nor U3086 (N_3086,N_1043,N_457);
nor U3087 (N_3087,N_604,N_270);
or U3088 (N_3088,N_1996,N_667);
nand U3089 (N_3089,N_1210,N_1374);
or U3090 (N_3090,N_1352,N_1649);
or U3091 (N_3091,N_1117,N_1334);
or U3092 (N_3092,N_1027,N_870);
nand U3093 (N_3093,N_442,N_1592);
and U3094 (N_3094,N_937,N_1998);
nor U3095 (N_3095,N_297,N_1761);
and U3096 (N_3096,N_828,N_1675);
nor U3097 (N_3097,N_1020,N_671);
nor U3098 (N_3098,N_370,N_853);
or U3099 (N_3099,N_905,N_1316);
nand U3100 (N_3100,N_1613,N_764);
nor U3101 (N_3101,N_1107,N_439);
nand U3102 (N_3102,N_943,N_664);
nor U3103 (N_3103,N_962,N_498);
and U3104 (N_3104,N_1331,N_1934);
and U3105 (N_3105,N_54,N_234);
nand U3106 (N_3106,N_500,N_1333);
and U3107 (N_3107,N_1769,N_461);
nor U3108 (N_3108,N_1196,N_417);
and U3109 (N_3109,N_76,N_524);
xnor U3110 (N_3110,N_1764,N_1847);
nand U3111 (N_3111,N_1331,N_1349);
nand U3112 (N_3112,N_523,N_1564);
nand U3113 (N_3113,N_1835,N_735);
or U3114 (N_3114,N_1216,N_588);
nor U3115 (N_3115,N_1113,N_1737);
nand U3116 (N_3116,N_1540,N_471);
nor U3117 (N_3117,N_1992,N_1137);
nor U3118 (N_3118,N_448,N_1702);
or U3119 (N_3119,N_269,N_1524);
and U3120 (N_3120,N_1390,N_759);
xor U3121 (N_3121,N_520,N_1317);
nand U3122 (N_3122,N_1368,N_1106);
nand U3123 (N_3123,N_917,N_1534);
nand U3124 (N_3124,N_1370,N_804);
or U3125 (N_3125,N_881,N_817);
and U3126 (N_3126,N_1401,N_1820);
or U3127 (N_3127,N_478,N_419);
nor U3128 (N_3128,N_990,N_1399);
or U3129 (N_3129,N_102,N_1829);
nor U3130 (N_3130,N_1386,N_149);
nor U3131 (N_3131,N_92,N_1871);
nand U3132 (N_3132,N_341,N_1992);
or U3133 (N_3133,N_1412,N_628);
or U3134 (N_3134,N_806,N_504);
nor U3135 (N_3135,N_1169,N_640);
nand U3136 (N_3136,N_1489,N_864);
xor U3137 (N_3137,N_1612,N_584);
and U3138 (N_3138,N_1558,N_415);
nor U3139 (N_3139,N_350,N_1641);
nor U3140 (N_3140,N_285,N_1586);
nand U3141 (N_3141,N_1703,N_933);
nand U3142 (N_3142,N_1710,N_928);
nor U3143 (N_3143,N_406,N_729);
nor U3144 (N_3144,N_1565,N_588);
or U3145 (N_3145,N_851,N_118);
nand U3146 (N_3146,N_1984,N_1541);
nand U3147 (N_3147,N_1681,N_980);
or U3148 (N_3148,N_1150,N_968);
nand U3149 (N_3149,N_178,N_802);
nor U3150 (N_3150,N_1371,N_1218);
or U3151 (N_3151,N_1643,N_1259);
and U3152 (N_3152,N_677,N_790);
and U3153 (N_3153,N_63,N_202);
or U3154 (N_3154,N_1578,N_1432);
and U3155 (N_3155,N_1461,N_867);
nand U3156 (N_3156,N_1138,N_611);
nand U3157 (N_3157,N_1747,N_1750);
nand U3158 (N_3158,N_1105,N_717);
nand U3159 (N_3159,N_1750,N_645);
nor U3160 (N_3160,N_1328,N_1639);
or U3161 (N_3161,N_602,N_1810);
nor U3162 (N_3162,N_953,N_1852);
nor U3163 (N_3163,N_622,N_1202);
nand U3164 (N_3164,N_1489,N_1142);
nand U3165 (N_3165,N_837,N_1440);
or U3166 (N_3166,N_948,N_783);
or U3167 (N_3167,N_1014,N_1142);
nand U3168 (N_3168,N_1110,N_1274);
and U3169 (N_3169,N_1496,N_984);
nand U3170 (N_3170,N_955,N_630);
xnor U3171 (N_3171,N_1733,N_582);
and U3172 (N_3172,N_735,N_854);
nand U3173 (N_3173,N_811,N_1308);
nor U3174 (N_3174,N_59,N_1245);
nor U3175 (N_3175,N_902,N_424);
or U3176 (N_3176,N_911,N_1633);
nand U3177 (N_3177,N_549,N_1641);
or U3178 (N_3178,N_1608,N_778);
nand U3179 (N_3179,N_1019,N_214);
and U3180 (N_3180,N_588,N_1026);
nand U3181 (N_3181,N_474,N_937);
nand U3182 (N_3182,N_1323,N_214);
and U3183 (N_3183,N_1911,N_1920);
nor U3184 (N_3184,N_746,N_1388);
nor U3185 (N_3185,N_224,N_656);
or U3186 (N_3186,N_798,N_1792);
and U3187 (N_3187,N_580,N_182);
nand U3188 (N_3188,N_1469,N_1369);
and U3189 (N_3189,N_192,N_1945);
nor U3190 (N_3190,N_394,N_319);
or U3191 (N_3191,N_1110,N_1036);
or U3192 (N_3192,N_1534,N_362);
or U3193 (N_3193,N_427,N_607);
nand U3194 (N_3194,N_1866,N_1795);
and U3195 (N_3195,N_1266,N_1035);
nor U3196 (N_3196,N_1449,N_37);
and U3197 (N_3197,N_343,N_1407);
nand U3198 (N_3198,N_55,N_668);
nor U3199 (N_3199,N_466,N_604);
nor U3200 (N_3200,N_1621,N_1003);
or U3201 (N_3201,N_240,N_1044);
nand U3202 (N_3202,N_1967,N_1950);
nor U3203 (N_3203,N_309,N_1363);
xnor U3204 (N_3204,N_1973,N_253);
or U3205 (N_3205,N_651,N_614);
and U3206 (N_3206,N_1193,N_698);
nor U3207 (N_3207,N_8,N_1522);
nand U3208 (N_3208,N_1114,N_40);
nor U3209 (N_3209,N_942,N_1777);
xor U3210 (N_3210,N_211,N_411);
and U3211 (N_3211,N_155,N_1460);
nor U3212 (N_3212,N_1756,N_706);
nand U3213 (N_3213,N_923,N_614);
nand U3214 (N_3214,N_1210,N_561);
or U3215 (N_3215,N_1917,N_486);
or U3216 (N_3216,N_215,N_131);
nor U3217 (N_3217,N_1090,N_1697);
xor U3218 (N_3218,N_1928,N_1011);
nor U3219 (N_3219,N_1809,N_1335);
or U3220 (N_3220,N_357,N_1186);
and U3221 (N_3221,N_794,N_1917);
or U3222 (N_3222,N_1613,N_1424);
and U3223 (N_3223,N_31,N_1575);
and U3224 (N_3224,N_1675,N_968);
nand U3225 (N_3225,N_575,N_1691);
and U3226 (N_3226,N_1289,N_1213);
nand U3227 (N_3227,N_707,N_643);
or U3228 (N_3228,N_1701,N_20);
or U3229 (N_3229,N_1940,N_1790);
nand U3230 (N_3230,N_367,N_742);
or U3231 (N_3231,N_1903,N_550);
or U3232 (N_3232,N_76,N_917);
nand U3233 (N_3233,N_879,N_748);
nor U3234 (N_3234,N_535,N_1395);
and U3235 (N_3235,N_1204,N_468);
or U3236 (N_3236,N_1061,N_1338);
or U3237 (N_3237,N_1234,N_793);
nor U3238 (N_3238,N_446,N_1660);
xnor U3239 (N_3239,N_1907,N_985);
or U3240 (N_3240,N_635,N_1088);
and U3241 (N_3241,N_733,N_747);
or U3242 (N_3242,N_1805,N_1271);
and U3243 (N_3243,N_772,N_1409);
nor U3244 (N_3244,N_315,N_705);
xor U3245 (N_3245,N_227,N_1928);
xnor U3246 (N_3246,N_644,N_720);
or U3247 (N_3247,N_471,N_428);
or U3248 (N_3248,N_443,N_1732);
nor U3249 (N_3249,N_1515,N_200);
and U3250 (N_3250,N_1468,N_1622);
nand U3251 (N_3251,N_1550,N_177);
nor U3252 (N_3252,N_1651,N_1262);
nand U3253 (N_3253,N_152,N_1623);
nand U3254 (N_3254,N_547,N_933);
nor U3255 (N_3255,N_1192,N_686);
or U3256 (N_3256,N_1731,N_1264);
and U3257 (N_3257,N_544,N_372);
or U3258 (N_3258,N_1842,N_1822);
nor U3259 (N_3259,N_894,N_108);
or U3260 (N_3260,N_730,N_519);
and U3261 (N_3261,N_1408,N_1608);
nand U3262 (N_3262,N_868,N_1938);
nor U3263 (N_3263,N_1169,N_1031);
and U3264 (N_3264,N_1639,N_250);
nand U3265 (N_3265,N_1693,N_322);
and U3266 (N_3266,N_1047,N_1719);
and U3267 (N_3267,N_1754,N_419);
or U3268 (N_3268,N_963,N_227);
or U3269 (N_3269,N_1285,N_133);
or U3270 (N_3270,N_1518,N_1780);
and U3271 (N_3271,N_1529,N_544);
or U3272 (N_3272,N_16,N_1773);
nor U3273 (N_3273,N_280,N_1656);
nor U3274 (N_3274,N_551,N_128);
nor U3275 (N_3275,N_89,N_1903);
nor U3276 (N_3276,N_627,N_487);
nor U3277 (N_3277,N_608,N_589);
and U3278 (N_3278,N_836,N_1211);
or U3279 (N_3279,N_355,N_99);
and U3280 (N_3280,N_960,N_1851);
nand U3281 (N_3281,N_661,N_1087);
or U3282 (N_3282,N_540,N_1371);
nor U3283 (N_3283,N_1613,N_200);
nor U3284 (N_3284,N_526,N_415);
xnor U3285 (N_3285,N_1540,N_1967);
and U3286 (N_3286,N_1739,N_927);
nand U3287 (N_3287,N_292,N_271);
nand U3288 (N_3288,N_1941,N_8);
and U3289 (N_3289,N_569,N_823);
or U3290 (N_3290,N_1423,N_936);
nor U3291 (N_3291,N_167,N_664);
nor U3292 (N_3292,N_1923,N_204);
and U3293 (N_3293,N_1817,N_1140);
and U3294 (N_3294,N_1240,N_253);
xnor U3295 (N_3295,N_730,N_710);
and U3296 (N_3296,N_665,N_729);
or U3297 (N_3297,N_23,N_443);
and U3298 (N_3298,N_920,N_29);
or U3299 (N_3299,N_1380,N_1217);
nor U3300 (N_3300,N_224,N_693);
nor U3301 (N_3301,N_752,N_762);
or U3302 (N_3302,N_1476,N_277);
or U3303 (N_3303,N_1133,N_1897);
nor U3304 (N_3304,N_1592,N_219);
or U3305 (N_3305,N_1946,N_680);
nand U3306 (N_3306,N_1433,N_210);
nand U3307 (N_3307,N_574,N_426);
or U3308 (N_3308,N_1361,N_1693);
or U3309 (N_3309,N_1436,N_0);
and U3310 (N_3310,N_527,N_875);
nand U3311 (N_3311,N_1910,N_1577);
or U3312 (N_3312,N_1224,N_714);
nor U3313 (N_3313,N_272,N_1674);
nor U3314 (N_3314,N_1629,N_1650);
or U3315 (N_3315,N_17,N_1280);
nand U3316 (N_3316,N_654,N_670);
or U3317 (N_3317,N_557,N_1385);
or U3318 (N_3318,N_729,N_974);
nand U3319 (N_3319,N_1734,N_737);
and U3320 (N_3320,N_1367,N_111);
nand U3321 (N_3321,N_1415,N_918);
nand U3322 (N_3322,N_779,N_1912);
or U3323 (N_3323,N_1889,N_45);
and U3324 (N_3324,N_1548,N_1979);
or U3325 (N_3325,N_1731,N_648);
nand U3326 (N_3326,N_94,N_551);
nand U3327 (N_3327,N_347,N_1251);
xor U3328 (N_3328,N_1405,N_1739);
xor U3329 (N_3329,N_1488,N_208);
nand U3330 (N_3330,N_1286,N_1987);
nand U3331 (N_3331,N_1495,N_1975);
nand U3332 (N_3332,N_545,N_1481);
and U3333 (N_3333,N_1220,N_972);
nand U3334 (N_3334,N_751,N_1752);
nand U3335 (N_3335,N_1766,N_1496);
and U3336 (N_3336,N_662,N_1170);
and U3337 (N_3337,N_112,N_606);
nand U3338 (N_3338,N_897,N_314);
nor U3339 (N_3339,N_1869,N_1616);
or U3340 (N_3340,N_1487,N_1087);
and U3341 (N_3341,N_656,N_1174);
nand U3342 (N_3342,N_588,N_927);
nand U3343 (N_3343,N_847,N_618);
xnor U3344 (N_3344,N_1454,N_589);
or U3345 (N_3345,N_943,N_1240);
nor U3346 (N_3346,N_1060,N_205);
or U3347 (N_3347,N_238,N_1917);
or U3348 (N_3348,N_817,N_1069);
nor U3349 (N_3349,N_553,N_1886);
or U3350 (N_3350,N_919,N_1690);
nor U3351 (N_3351,N_570,N_744);
nor U3352 (N_3352,N_770,N_117);
nor U3353 (N_3353,N_1177,N_186);
or U3354 (N_3354,N_645,N_1280);
nand U3355 (N_3355,N_1045,N_667);
nor U3356 (N_3356,N_1136,N_1126);
and U3357 (N_3357,N_1671,N_757);
and U3358 (N_3358,N_1471,N_1021);
or U3359 (N_3359,N_7,N_1996);
nor U3360 (N_3360,N_1665,N_682);
xnor U3361 (N_3361,N_287,N_896);
nand U3362 (N_3362,N_1180,N_496);
xor U3363 (N_3363,N_1176,N_619);
nor U3364 (N_3364,N_1315,N_934);
nor U3365 (N_3365,N_1197,N_96);
nor U3366 (N_3366,N_124,N_1036);
nor U3367 (N_3367,N_338,N_110);
nor U3368 (N_3368,N_433,N_1818);
and U3369 (N_3369,N_799,N_905);
and U3370 (N_3370,N_1623,N_954);
nor U3371 (N_3371,N_128,N_1569);
or U3372 (N_3372,N_417,N_313);
nor U3373 (N_3373,N_908,N_280);
xor U3374 (N_3374,N_1686,N_1420);
nand U3375 (N_3375,N_1326,N_1742);
xor U3376 (N_3376,N_597,N_97);
and U3377 (N_3377,N_1469,N_1122);
nand U3378 (N_3378,N_841,N_1718);
xor U3379 (N_3379,N_836,N_83);
and U3380 (N_3380,N_1,N_729);
nor U3381 (N_3381,N_975,N_658);
or U3382 (N_3382,N_529,N_37);
nor U3383 (N_3383,N_730,N_890);
xor U3384 (N_3384,N_733,N_1266);
and U3385 (N_3385,N_1581,N_1919);
or U3386 (N_3386,N_1753,N_32);
or U3387 (N_3387,N_1121,N_1375);
nand U3388 (N_3388,N_475,N_954);
nor U3389 (N_3389,N_733,N_722);
nor U3390 (N_3390,N_317,N_1811);
or U3391 (N_3391,N_136,N_169);
or U3392 (N_3392,N_350,N_1653);
nor U3393 (N_3393,N_488,N_453);
xnor U3394 (N_3394,N_1244,N_308);
and U3395 (N_3395,N_952,N_965);
xor U3396 (N_3396,N_1267,N_1055);
nand U3397 (N_3397,N_1156,N_1260);
nor U3398 (N_3398,N_1148,N_1415);
nor U3399 (N_3399,N_964,N_350);
and U3400 (N_3400,N_602,N_1580);
or U3401 (N_3401,N_1958,N_996);
and U3402 (N_3402,N_1820,N_199);
nand U3403 (N_3403,N_556,N_179);
nor U3404 (N_3404,N_28,N_1022);
nor U3405 (N_3405,N_289,N_1816);
or U3406 (N_3406,N_1379,N_860);
nor U3407 (N_3407,N_1395,N_1377);
or U3408 (N_3408,N_1084,N_1071);
xor U3409 (N_3409,N_1271,N_1607);
and U3410 (N_3410,N_1546,N_107);
or U3411 (N_3411,N_118,N_614);
and U3412 (N_3412,N_1249,N_357);
xor U3413 (N_3413,N_1398,N_1705);
nor U3414 (N_3414,N_778,N_561);
or U3415 (N_3415,N_1215,N_1480);
nand U3416 (N_3416,N_1445,N_1399);
and U3417 (N_3417,N_225,N_197);
nand U3418 (N_3418,N_883,N_1154);
and U3419 (N_3419,N_46,N_997);
nor U3420 (N_3420,N_774,N_881);
or U3421 (N_3421,N_1381,N_1200);
or U3422 (N_3422,N_1474,N_1343);
and U3423 (N_3423,N_650,N_636);
and U3424 (N_3424,N_1108,N_1470);
nor U3425 (N_3425,N_100,N_1560);
and U3426 (N_3426,N_773,N_108);
and U3427 (N_3427,N_1212,N_540);
nand U3428 (N_3428,N_420,N_1796);
and U3429 (N_3429,N_268,N_886);
nor U3430 (N_3430,N_1454,N_1765);
or U3431 (N_3431,N_75,N_265);
and U3432 (N_3432,N_798,N_909);
nand U3433 (N_3433,N_58,N_1519);
nand U3434 (N_3434,N_1624,N_1613);
nor U3435 (N_3435,N_813,N_1817);
nor U3436 (N_3436,N_651,N_1886);
nand U3437 (N_3437,N_1019,N_483);
nand U3438 (N_3438,N_934,N_171);
nor U3439 (N_3439,N_1532,N_629);
or U3440 (N_3440,N_1333,N_1769);
and U3441 (N_3441,N_1668,N_725);
nand U3442 (N_3442,N_614,N_1056);
nor U3443 (N_3443,N_1961,N_800);
nand U3444 (N_3444,N_1609,N_470);
nor U3445 (N_3445,N_801,N_1077);
and U3446 (N_3446,N_1332,N_1382);
and U3447 (N_3447,N_491,N_427);
or U3448 (N_3448,N_1298,N_660);
or U3449 (N_3449,N_225,N_951);
and U3450 (N_3450,N_1669,N_47);
nor U3451 (N_3451,N_442,N_1323);
and U3452 (N_3452,N_1391,N_1113);
nand U3453 (N_3453,N_1127,N_1460);
nor U3454 (N_3454,N_494,N_584);
or U3455 (N_3455,N_342,N_1814);
nand U3456 (N_3456,N_736,N_1744);
or U3457 (N_3457,N_673,N_589);
xnor U3458 (N_3458,N_1790,N_1236);
or U3459 (N_3459,N_604,N_1697);
nand U3460 (N_3460,N_1881,N_535);
and U3461 (N_3461,N_232,N_202);
or U3462 (N_3462,N_1832,N_106);
nor U3463 (N_3463,N_402,N_1215);
or U3464 (N_3464,N_607,N_1394);
or U3465 (N_3465,N_1107,N_1649);
or U3466 (N_3466,N_719,N_1651);
or U3467 (N_3467,N_310,N_917);
nand U3468 (N_3468,N_945,N_409);
xor U3469 (N_3469,N_488,N_529);
nand U3470 (N_3470,N_1619,N_1204);
or U3471 (N_3471,N_513,N_1833);
nand U3472 (N_3472,N_120,N_1000);
or U3473 (N_3473,N_1654,N_216);
nand U3474 (N_3474,N_383,N_1486);
nand U3475 (N_3475,N_1760,N_493);
nand U3476 (N_3476,N_1401,N_292);
nand U3477 (N_3477,N_334,N_973);
xnor U3478 (N_3478,N_183,N_25);
or U3479 (N_3479,N_1819,N_1172);
and U3480 (N_3480,N_28,N_1814);
nor U3481 (N_3481,N_900,N_800);
and U3482 (N_3482,N_321,N_1823);
or U3483 (N_3483,N_360,N_1798);
or U3484 (N_3484,N_1276,N_858);
nor U3485 (N_3485,N_1293,N_1618);
or U3486 (N_3486,N_1907,N_659);
nand U3487 (N_3487,N_717,N_1769);
and U3488 (N_3488,N_313,N_1479);
and U3489 (N_3489,N_943,N_78);
xnor U3490 (N_3490,N_1415,N_692);
nand U3491 (N_3491,N_1076,N_1432);
or U3492 (N_3492,N_147,N_133);
and U3493 (N_3493,N_1336,N_1338);
nand U3494 (N_3494,N_1449,N_764);
and U3495 (N_3495,N_1737,N_310);
nand U3496 (N_3496,N_1670,N_1304);
and U3497 (N_3497,N_1542,N_767);
nand U3498 (N_3498,N_480,N_1364);
and U3499 (N_3499,N_1140,N_340);
nor U3500 (N_3500,N_924,N_471);
and U3501 (N_3501,N_1057,N_738);
nor U3502 (N_3502,N_554,N_945);
nor U3503 (N_3503,N_68,N_1654);
or U3504 (N_3504,N_998,N_1685);
nand U3505 (N_3505,N_1972,N_1520);
xor U3506 (N_3506,N_989,N_1737);
nand U3507 (N_3507,N_1890,N_688);
and U3508 (N_3508,N_1207,N_422);
nor U3509 (N_3509,N_1956,N_1917);
or U3510 (N_3510,N_1712,N_1982);
nand U3511 (N_3511,N_821,N_1840);
nand U3512 (N_3512,N_107,N_1897);
nand U3513 (N_3513,N_354,N_627);
or U3514 (N_3514,N_1008,N_423);
nor U3515 (N_3515,N_559,N_371);
or U3516 (N_3516,N_1284,N_818);
nor U3517 (N_3517,N_932,N_1100);
or U3518 (N_3518,N_548,N_149);
nand U3519 (N_3519,N_1627,N_1144);
nor U3520 (N_3520,N_1152,N_971);
and U3521 (N_3521,N_725,N_935);
or U3522 (N_3522,N_1023,N_516);
nor U3523 (N_3523,N_723,N_1051);
xnor U3524 (N_3524,N_1418,N_867);
and U3525 (N_3525,N_1428,N_1068);
nand U3526 (N_3526,N_1375,N_133);
nand U3527 (N_3527,N_207,N_14);
nor U3528 (N_3528,N_1515,N_1405);
nor U3529 (N_3529,N_562,N_783);
nor U3530 (N_3530,N_501,N_1186);
nor U3531 (N_3531,N_1002,N_593);
nand U3532 (N_3532,N_228,N_1922);
nor U3533 (N_3533,N_671,N_536);
and U3534 (N_3534,N_1946,N_1125);
nor U3535 (N_3535,N_1151,N_1802);
or U3536 (N_3536,N_1771,N_808);
nor U3537 (N_3537,N_1315,N_687);
nor U3538 (N_3538,N_470,N_188);
nor U3539 (N_3539,N_670,N_1152);
or U3540 (N_3540,N_1490,N_1507);
nand U3541 (N_3541,N_961,N_686);
and U3542 (N_3542,N_127,N_1854);
nand U3543 (N_3543,N_1376,N_402);
nor U3544 (N_3544,N_677,N_564);
and U3545 (N_3545,N_598,N_179);
nor U3546 (N_3546,N_823,N_898);
nor U3547 (N_3547,N_372,N_237);
nand U3548 (N_3548,N_1764,N_555);
nor U3549 (N_3549,N_1556,N_1056);
or U3550 (N_3550,N_807,N_1334);
or U3551 (N_3551,N_1063,N_1142);
and U3552 (N_3552,N_1152,N_64);
and U3553 (N_3553,N_340,N_143);
nand U3554 (N_3554,N_1894,N_246);
xor U3555 (N_3555,N_1291,N_1799);
nand U3556 (N_3556,N_1727,N_433);
nand U3557 (N_3557,N_553,N_1826);
nor U3558 (N_3558,N_1036,N_508);
xnor U3559 (N_3559,N_1933,N_496);
nand U3560 (N_3560,N_581,N_1809);
nand U3561 (N_3561,N_29,N_508);
xor U3562 (N_3562,N_681,N_960);
or U3563 (N_3563,N_222,N_14);
nand U3564 (N_3564,N_1855,N_1833);
xnor U3565 (N_3565,N_1336,N_1671);
nor U3566 (N_3566,N_1071,N_117);
nor U3567 (N_3567,N_50,N_1867);
or U3568 (N_3568,N_1288,N_690);
or U3569 (N_3569,N_764,N_768);
nand U3570 (N_3570,N_1697,N_932);
nor U3571 (N_3571,N_1177,N_1343);
nand U3572 (N_3572,N_536,N_18);
or U3573 (N_3573,N_437,N_986);
nor U3574 (N_3574,N_702,N_1523);
nor U3575 (N_3575,N_43,N_415);
and U3576 (N_3576,N_629,N_1213);
nor U3577 (N_3577,N_727,N_1212);
nor U3578 (N_3578,N_1105,N_1962);
nand U3579 (N_3579,N_1267,N_1070);
or U3580 (N_3580,N_791,N_894);
nor U3581 (N_3581,N_136,N_1245);
nor U3582 (N_3582,N_1371,N_712);
nor U3583 (N_3583,N_1761,N_940);
nor U3584 (N_3584,N_51,N_1524);
nor U3585 (N_3585,N_1336,N_627);
nor U3586 (N_3586,N_271,N_87);
or U3587 (N_3587,N_1518,N_835);
nor U3588 (N_3588,N_1060,N_919);
or U3589 (N_3589,N_835,N_137);
or U3590 (N_3590,N_1707,N_334);
and U3591 (N_3591,N_658,N_1290);
nand U3592 (N_3592,N_232,N_1391);
nand U3593 (N_3593,N_1121,N_502);
or U3594 (N_3594,N_1132,N_727);
nor U3595 (N_3595,N_1266,N_1067);
xnor U3596 (N_3596,N_1901,N_1213);
nand U3597 (N_3597,N_787,N_378);
and U3598 (N_3598,N_779,N_288);
or U3599 (N_3599,N_819,N_331);
or U3600 (N_3600,N_1827,N_494);
or U3601 (N_3601,N_481,N_1830);
xor U3602 (N_3602,N_208,N_1825);
xnor U3603 (N_3603,N_2,N_1408);
or U3604 (N_3604,N_1248,N_11);
or U3605 (N_3605,N_1733,N_980);
or U3606 (N_3606,N_1008,N_678);
and U3607 (N_3607,N_1445,N_1567);
nand U3608 (N_3608,N_1768,N_465);
nand U3609 (N_3609,N_284,N_581);
or U3610 (N_3610,N_1874,N_1588);
or U3611 (N_3611,N_379,N_1956);
and U3612 (N_3612,N_91,N_1392);
nor U3613 (N_3613,N_618,N_496);
nor U3614 (N_3614,N_1081,N_1308);
nor U3615 (N_3615,N_13,N_720);
or U3616 (N_3616,N_468,N_89);
nand U3617 (N_3617,N_1353,N_735);
or U3618 (N_3618,N_1475,N_1095);
and U3619 (N_3619,N_1782,N_1954);
and U3620 (N_3620,N_65,N_1682);
or U3621 (N_3621,N_1538,N_1088);
xnor U3622 (N_3622,N_1843,N_1805);
and U3623 (N_3623,N_1154,N_452);
and U3624 (N_3624,N_225,N_528);
nor U3625 (N_3625,N_1980,N_1716);
nand U3626 (N_3626,N_613,N_106);
nand U3627 (N_3627,N_1886,N_1907);
xnor U3628 (N_3628,N_809,N_724);
and U3629 (N_3629,N_642,N_1903);
nor U3630 (N_3630,N_883,N_387);
nor U3631 (N_3631,N_563,N_1986);
or U3632 (N_3632,N_1142,N_1506);
nor U3633 (N_3633,N_1783,N_217);
nand U3634 (N_3634,N_984,N_1100);
nor U3635 (N_3635,N_1069,N_1221);
and U3636 (N_3636,N_632,N_566);
nor U3637 (N_3637,N_1607,N_238);
nand U3638 (N_3638,N_1832,N_587);
and U3639 (N_3639,N_1023,N_1599);
nor U3640 (N_3640,N_38,N_478);
and U3641 (N_3641,N_1127,N_139);
and U3642 (N_3642,N_963,N_709);
and U3643 (N_3643,N_1619,N_1140);
and U3644 (N_3644,N_1089,N_380);
or U3645 (N_3645,N_102,N_1311);
and U3646 (N_3646,N_1400,N_1246);
xor U3647 (N_3647,N_985,N_278);
or U3648 (N_3648,N_258,N_1351);
nor U3649 (N_3649,N_1401,N_1275);
and U3650 (N_3650,N_119,N_1694);
nand U3651 (N_3651,N_52,N_1051);
nor U3652 (N_3652,N_537,N_1215);
or U3653 (N_3653,N_1344,N_1057);
and U3654 (N_3654,N_1694,N_1940);
and U3655 (N_3655,N_1633,N_1562);
nand U3656 (N_3656,N_1977,N_548);
and U3657 (N_3657,N_1708,N_1588);
and U3658 (N_3658,N_1835,N_1186);
or U3659 (N_3659,N_490,N_1276);
xnor U3660 (N_3660,N_1298,N_212);
and U3661 (N_3661,N_280,N_935);
nand U3662 (N_3662,N_1204,N_1490);
or U3663 (N_3663,N_1973,N_1290);
nand U3664 (N_3664,N_1232,N_460);
or U3665 (N_3665,N_1167,N_594);
nand U3666 (N_3666,N_1048,N_1411);
or U3667 (N_3667,N_1135,N_488);
and U3668 (N_3668,N_562,N_334);
nor U3669 (N_3669,N_1051,N_492);
or U3670 (N_3670,N_702,N_283);
or U3671 (N_3671,N_1592,N_1663);
and U3672 (N_3672,N_1440,N_1502);
or U3673 (N_3673,N_484,N_804);
or U3674 (N_3674,N_15,N_1645);
nand U3675 (N_3675,N_1821,N_943);
nand U3676 (N_3676,N_1229,N_552);
and U3677 (N_3677,N_346,N_987);
nor U3678 (N_3678,N_1864,N_1550);
nand U3679 (N_3679,N_779,N_255);
and U3680 (N_3680,N_655,N_1022);
or U3681 (N_3681,N_859,N_1885);
nand U3682 (N_3682,N_561,N_952);
and U3683 (N_3683,N_755,N_611);
nor U3684 (N_3684,N_841,N_451);
nor U3685 (N_3685,N_793,N_381);
or U3686 (N_3686,N_170,N_700);
nor U3687 (N_3687,N_1244,N_187);
nand U3688 (N_3688,N_500,N_1981);
xnor U3689 (N_3689,N_964,N_1781);
or U3690 (N_3690,N_815,N_371);
or U3691 (N_3691,N_375,N_1423);
nor U3692 (N_3692,N_1837,N_1952);
or U3693 (N_3693,N_54,N_1981);
or U3694 (N_3694,N_181,N_3);
xnor U3695 (N_3695,N_1736,N_886);
nand U3696 (N_3696,N_964,N_1763);
or U3697 (N_3697,N_271,N_555);
and U3698 (N_3698,N_302,N_1053);
nor U3699 (N_3699,N_17,N_148);
nand U3700 (N_3700,N_1979,N_345);
and U3701 (N_3701,N_1866,N_722);
or U3702 (N_3702,N_1950,N_317);
and U3703 (N_3703,N_1765,N_1108);
and U3704 (N_3704,N_17,N_90);
nor U3705 (N_3705,N_1980,N_1414);
or U3706 (N_3706,N_1111,N_1098);
and U3707 (N_3707,N_1690,N_687);
nor U3708 (N_3708,N_107,N_1158);
or U3709 (N_3709,N_205,N_375);
xor U3710 (N_3710,N_850,N_1369);
nand U3711 (N_3711,N_893,N_409);
nor U3712 (N_3712,N_458,N_1220);
nand U3713 (N_3713,N_705,N_1179);
nor U3714 (N_3714,N_1329,N_1423);
and U3715 (N_3715,N_640,N_1613);
or U3716 (N_3716,N_606,N_1502);
or U3717 (N_3717,N_842,N_1652);
and U3718 (N_3718,N_326,N_191);
or U3719 (N_3719,N_456,N_616);
and U3720 (N_3720,N_1861,N_117);
nor U3721 (N_3721,N_728,N_934);
nor U3722 (N_3722,N_632,N_513);
xor U3723 (N_3723,N_1103,N_870);
nand U3724 (N_3724,N_1814,N_32);
nor U3725 (N_3725,N_1830,N_1182);
and U3726 (N_3726,N_402,N_1670);
or U3727 (N_3727,N_1094,N_1224);
nand U3728 (N_3728,N_60,N_98);
and U3729 (N_3729,N_1093,N_134);
or U3730 (N_3730,N_1466,N_187);
or U3731 (N_3731,N_810,N_1954);
nand U3732 (N_3732,N_1282,N_40);
and U3733 (N_3733,N_132,N_641);
nor U3734 (N_3734,N_419,N_1099);
or U3735 (N_3735,N_880,N_1781);
nand U3736 (N_3736,N_245,N_1857);
and U3737 (N_3737,N_1307,N_610);
nand U3738 (N_3738,N_1875,N_713);
nor U3739 (N_3739,N_345,N_1600);
and U3740 (N_3740,N_113,N_1248);
or U3741 (N_3741,N_1340,N_1176);
or U3742 (N_3742,N_798,N_1153);
and U3743 (N_3743,N_1923,N_510);
nor U3744 (N_3744,N_151,N_844);
or U3745 (N_3745,N_584,N_1784);
xnor U3746 (N_3746,N_120,N_732);
nand U3747 (N_3747,N_1633,N_1901);
nand U3748 (N_3748,N_1544,N_387);
nand U3749 (N_3749,N_529,N_1887);
or U3750 (N_3750,N_17,N_361);
nor U3751 (N_3751,N_1951,N_1070);
or U3752 (N_3752,N_1882,N_422);
and U3753 (N_3753,N_99,N_1273);
xnor U3754 (N_3754,N_316,N_1219);
nand U3755 (N_3755,N_1172,N_1335);
or U3756 (N_3756,N_1472,N_887);
nand U3757 (N_3757,N_1012,N_494);
nor U3758 (N_3758,N_757,N_1691);
or U3759 (N_3759,N_417,N_327);
and U3760 (N_3760,N_1766,N_1870);
xor U3761 (N_3761,N_1561,N_899);
nand U3762 (N_3762,N_1614,N_871);
or U3763 (N_3763,N_849,N_472);
and U3764 (N_3764,N_1985,N_1945);
nand U3765 (N_3765,N_340,N_1838);
nand U3766 (N_3766,N_408,N_1560);
nand U3767 (N_3767,N_1891,N_549);
or U3768 (N_3768,N_602,N_154);
nor U3769 (N_3769,N_1829,N_13);
nand U3770 (N_3770,N_247,N_398);
xor U3771 (N_3771,N_181,N_1647);
nand U3772 (N_3772,N_1169,N_617);
and U3773 (N_3773,N_1059,N_617);
or U3774 (N_3774,N_1685,N_1919);
nand U3775 (N_3775,N_95,N_1300);
nand U3776 (N_3776,N_1960,N_434);
or U3777 (N_3777,N_1924,N_1063);
or U3778 (N_3778,N_201,N_440);
nand U3779 (N_3779,N_1949,N_81);
nor U3780 (N_3780,N_1707,N_662);
and U3781 (N_3781,N_96,N_822);
nor U3782 (N_3782,N_557,N_1654);
or U3783 (N_3783,N_192,N_1878);
or U3784 (N_3784,N_130,N_431);
nand U3785 (N_3785,N_1730,N_1557);
or U3786 (N_3786,N_641,N_1696);
or U3787 (N_3787,N_1965,N_924);
or U3788 (N_3788,N_813,N_705);
nand U3789 (N_3789,N_1441,N_184);
nand U3790 (N_3790,N_269,N_998);
or U3791 (N_3791,N_1655,N_643);
nor U3792 (N_3792,N_232,N_1075);
or U3793 (N_3793,N_1187,N_1971);
or U3794 (N_3794,N_1495,N_6);
nand U3795 (N_3795,N_1524,N_1898);
nand U3796 (N_3796,N_1131,N_1251);
nor U3797 (N_3797,N_171,N_684);
nand U3798 (N_3798,N_1952,N_1367);
nor U3799 (N_3799,N_1789,N_964);
nor U3800 (N_3800,N_993,N_1571);
nand U3801 (N_3801,N_224,N_1481);
and U3802 (N_3802,N_682,N_1103);
nor U3803 (N_3803,N_821,N_278);
nor U3804 (N_3804,N_1558,N_1336);
nand U3805 (N_3805,N_1204,N_1527);
nor U3806 (N_3806,N_1651,N_510);
or U3807 (N_3807,N_1961,N_719);
nor U3808 (N_3808,N_1076,N_237);
nand U3809 (N_3809,N_338,N_1187);
nand U3810 (N_3810,N_1323,N_1168);
or U3811 (N_3811,N_1502,N_1490);
or U3812 (N_3812,N_1337,N_933);
or U3813 (N_3813,N_1974,N_177);
or U3814 (N_3814,N_968,N_114);
nor U3815 (N_3815,N_900,N_1352);
nor U3816 (N_3816,N_1550,N_315);
or U3817 (N_3817,N_1799,N_1598);
and U3818 (N_3818,N_390,N_1393);
nand U3819 (N_3819,N_1888,N_1148);
nor U3820 (N_3820,N_1356,N_1502);
nand U3821 (N_3821,N_1107,N_21);
nor U3822 (N_3822,N_666,N_1398);
xor U3823 (N_3823,N_1563,N_556);
or U3824 (N_3824,N_1497,N_1901);
nand U3825 (N_3825,N_755,N_307);
or U3826 (N_3826,N_1222,N_471);
or U3827 (N_3827,N_212,N_1514);
and U3828 (N_3828,N_1818,N_413);
and U3829 (N_3829,N_356,N_1810);
xor U3830 (N_3830,N_395,N_1805);
and U3831 (N_3831,N_713,N_1230);
and U3832 (N_3832,N_144,N_254);
or U3833 (N_3833,N_1141,N_185);
nand U3834 (N_3834,N_1631,N_877);
nand U3835 (N_3835,N_1667,N_1191);
and U3836 (N_3836,N_1321,N_1850);
and U3837 (N_3837,N_1053,N_1151);
nand U3838 (N_3838,N_1513,N_1111);
nand U3839 (N_3839,N_1661,N_1534);
or U3840 (N_3840,N_1455,N_576);
or U3841 (N_3841,N_1147,N_1921);
nand U3842 (N_3842,N_835,N_1305);
and U3843 (N_3843,N_18,N_1794);
xnor U3844 (N_3844,N_410,N_839);
and U3845 (N_3845,N_1395,N_170);
nor U3846 (N_3846,N_720,N_636);
or U3847 (N_3847,N_220,N_460);
or U3848 (N_3848,N_682,N_1849);
or U3849 (N_3849,N_246,N_1630);
xor U3850 (N_3850,N_1002,N_615);
or U3851 (N_3851,N_564,N_301);
and U3852 (N_3852,N_158,N_847);
or U3853 (N_3853,N_1699,N_1901);
and U3854 (N_3854,N_418,N_663);
and U3855 (N_3855,N_1262,N_1507);
or U3856 (N_3856,N_1017,N_1002);
or U3857 (N_3857,N_1158,N_287);
or U3858 (N_3858,N_1159,N_1431);
nand U3859 (N_3859,N_1981,N_738);
and U3860 (N_3860,N_1694,N_592);
nor U3861 (N_3861,N_1138,N_1842);
or U3862 (N_3862,N_1239,N_1985);
nand U3863 (N_3863,N_339,N_391);
nor U3864 (N_3864,N_658,N_1225);
and U3865 (N_3865,N_945,N_21);
nand U3866 (N_3866,N_1374,N_589);
and U3867 (N_3867,N_39,N_1209);
nor U3868 (N_3868,N_1853,N_47);
or U3869 (N_3869,N_1207,N_325);
xnor U3870 (N_3870,N_626,N_897);
or U3871 (N_3871,N_452,N_1196);
or U3872 (N_3872,N_799,N_1627);
or U3873 (N_3873,N_1180,N_860);
nor U3874 (N_3874,N_1137,N_573);
nor U3875 (N_3875,N_994,N_93);
or U3876 (N_3876,N_1882,N_1664);
nand U3877 (N_3877,N_737,N_1968);
and U3878 (N_3878,N_550,N_1885);
and U3879 (N_3879,N_862,N_139);
or U3880 (N_3880,N_1750,N_159);
or U3881 (N_3881,N_1772,N_1795);
nor U3882 (N_3882,N_524,N_617);
nor U3883 (N_3883,N_1268,N_1408);
and U3884 (N_3884,N_782,N_484);
and U3885 (N_3885,N_1419,N_843);
xor U3886 (N_3886,N_479,N_1127);
nand U3887 (N_3887,N_989,N_1156);
or U3888 (N_3888,N_1102,N_1020);
nor U3889 (N_3889,N_1959,N_1658);
and U3890 (N_3890,N_648,N_460);
and U3891 (N_3891,N_796,N_112);
nor U3892 (N_3892,N_1692,N_1317);
nor U3893 (N_3893,N_198,N_742);
and U3894 (N_3894,N_1742,N_1948);
and U3895 (N_3895,N_1723,N_47);
nand U3896 (N_3896,N_584,N_464);
nor U3897 (N_3897,N_69,N_1734);
nand U3898 (N_3898,N_1859,N_1338);
nand U3899 (N_3899,N_1448,N_644);
nor U3900 (N_3900,N_308,N_422);
nor U3901 (N_3901,N_1062,N_201);
and U3902 (N_3902,N_1677,N_1846);
nor U3903 (N_3903,N_1883,N_1539);
nor U3904 (N_3904,N_900,N_410);
nand U3905 (N_3905,N_10,N_1079);
and U3906 (N_3906,N_1645,N_1474);
nand U3907 (N_3907,N_852,N_965);
or U3908 (N_3908,N_1977,N_439);
and U3909 (N_3909,N_83,N_1542);
or U3910 (N_3910,N_745,N_1361);
and U3911 (N_3911,N_1756,N_1585);
nor U3912 (N_3912,N_1390,N_451);
nand U3913 (N_3913,N_1436,N_1480);
nand U3914 (N_3914,N_394,N_946);
nor U3915 (N_3915,N_481,N_1922);
nor U3916 (N_3916,N_811,N_312);
or U3917 (N_3917,N_904,N_1135);
or U3918 (N_3918,N_1306,N_1197);
and U3919 (N_3919,N_914,N_918);
or U3920 (N_3920,N_824,N_1758);
xnor U3921 (N_3921,N_546,N_1872);
nand U3922 (N_3922,N_609,N_688);
nand U3923 (N_3923,N_1160,N_1826);
nand U3924 (N_3924,N_977,N_1847);
xnor U3925 (N_3925,N_598,N_1495);
and U3926 (N_3926,N_234,N_1425);
nor U3927 (N_3927,N_738,N_1542);
or U3928 (N_3928,N_1333,N_1205);
and U3929 (N_3929,N_993,N_687);
nand U3930 (N_3930,N_1786,N_1992);
and U3931 (N_3931,N_392,N_1206);
or U3932 (N_3932,N_424,N_1093);
nand U3933 (N_3933,N_1845,N_744);
nor U3934 (N_3934,N_1506,N_484);
nor U3935 (N_3935,N_1883,N_832);
and U3936 (N_3936,N_366,N_1053);
and U3937 (N_3937,N_1176,N_1610);
or U3938 (N_3938,N_744,N_1969);
and U3939 (N_3939,N_1114,N_822);
and U3940 (N_3940,N_672,N_1682);
or U3941 (N_3941,N_997,N_1545);
or U3942 (N_3942,N_155,N_834);
and U3943 (N_3943,N_1640,N_1874);
or U3944 (N_3944,N_846,N_867);
and U3945 (N_3945,N_1912,N_1091);
nor U3946 (N_3946,N_1158,N_211);
or U3947 (N_3947,N_1891,N_1838);
and U3948 (N_3948,N_912,N_1956);
or U3949 (N_3949,N_216,N_1418);
and U3950 (N_3950,N_1030,N_242);
or U3951 (N_3951,N_753,N_1571);
or U3952 (N_3952,N_1504,N_301);
and U3953 (N_3953,N_1607,N_982);
nor U3954 (N_3954,N_1138,N_1024);
nor U3955 (N_3955,N_1701,N_401);
nor U3956 (N_3956,N_270,N_1451);
nor U3957 (N_3957,N_1069,N_1828);
and U3958 (N_3958,N_713,N_314);
xor U3959 (N_3959,N_685,N_1360);
and U3960 (N_3960,N_712,N_297);
nand U3961 (N_3961,N_696,N_45);
nor U3962 (N_3962,N_25,N_1242);
nand U3963 (N_3963,N_372,N_743);
or U3964 (N_3964,N_1943,N_839);
and U3965 (N_3965,N_468,N_1839);
xnor U3966 (N_3966,N_900,N_1499);
and U3967 (N_3967,N_661,N_100);
xor U3968 (N_3968,N_109,N_1006);
nand U3969 (N_3969,N_1866,N_801);
xnor U3970 (N_3970,N_1809,N_693);
and U3971 (N_3971,N_1157,N_948);
nor U3972 (N_3972,N_1404,N_50);
or U3973 (N_3973,N_885,N_253);
xnor U3974 (N_3974,N_981,N_1003);
and U3975 (N_3975,N_761,N_168);
nor U3976 (N_3976,N_413,N_1903);
and U3977 (N_3977,N_1113,N_1894);
nand U3978 (N_3978,N_1294,N_817);
or U3979 (N_3979,N_656,N_1728);
and U3980 (N_3980,N_1315,N_527);
and U3981 (N_3981,N_1406,N_540);
or U3982 (N_3982,N_1905,N_1647);
nand U3983 (N_3983,N_1942,N_1455);
or U3984 (N_3984,N_336,N_685);
nor U3985 (N_3985,N_685,N_1500);
and U3986 (N_3986,N_1437,N_82);
and U3987 (N_3987,N_1709,N_508);
nor U3988 (N_3988,N_1664,N_71);
and U3989 (N_3989,N_1384,N_814);
or U3990 (N_3990,N_270,N_131);
or U3991 (N_3991,N_1409,N_1044);
and U3992 (N_3992,N_404,N_328);
and U3993 (N_3993,N_1648,N_676);
or U3994 (N_3994,N_1319,N_757);
nor U3995 (N_3995,N_616,N_1309);
nor U3996 (N_3996,N_965,N_1324);
or U3997 (N_3997,N_32,N_275);
xor U3998 (N_3998,N_323,N_1069);
or U3999 (N_3999,N_291,N_1253);
and U4000 (N_4000,N_2299,N_3340);
nor U4001 (N_4001,N_2088,N_3290);
or U4002 (N_4002,N_3672,N_3287);
nand U4003 (N_4003,N_2631,N_2650);
nor U4004 (N_4004,N_2349,N_2228);
xor U4005 (N_4005,N_2147,N_2905);
nor U4006 (N_4006,N_2948,N_2420);
and U4007 (N_4007,N_2259,N_2310);
nand U4008 (N_4008,N_3766,N_3241);
nand U4009 (N_4009,N_2790,N_2331);
or U4010 (N_4010,N_3623,N_2380);
or U4011 (N_4011,N_2745,N_2936);
nand U4012 (N_4012,N_3940,N_2467);
xor U4013 (N_4013,N_2158,N_2181);
nor U4014 (N_4014,N_2030,N_3110);
nor U4015 (N_4015,N_2061,N_2086);
nor U4016 (N_4016,N_3432,N_3419);
or U4017 (N_4017,N_3436,N_3918);
nand U4018 (N_4018,N_2332,N_2084);
nor U4019 (N_4019,N_3178,N_3488);
nand U4020 (N_4020,N_2895,N_2796);
nor U4021 (N_4021,N_3261,N_3701);
nor U4022 (N_4022,N_3602,N_3556);
xor U4023 (N_4023,N_2763,N_2060);
and U4024 (N_4024,N_2369,N_2969);
nor U4025 (N_4025,N_3197,N_3743);
and U4026 (N_4026,N_2643,N_2987);
nor U4027 (N_4027,N_3509,N_3513);
xnor U4028 (N_4028,N_3267,N_3729);
or U4029 (N_4029,N_2548,N_3664);
or U4030 (N_4030,N_3221,N_2012);
and U4031 (N_4031,N_3304,N_3062);
and U4032 (N_4032,N_2191,N_3022);
and U4033 (N_4033,N_3656,N_2511);
nor U4034 (N_4034,N_3210,N_2142);
or U4035 (N_4035,N_2924,N_3390);
or U4036 (N_4036,N_3652,N_2862);
nor U4037 (N_4037,N_2661,N_2907);
and U4038 (N_4038,N_2094,N_3228);
or U4039 (N_4039,N_2351,N_2381);
or U4040 (N_4040,N_3712,N_2513);
nor U4041 (N_4041,N_2001,N_2446);
nand U4042 (N_4042,N_3620,N_2937);
nand U4043 (N_4043,N_3342,N_2676);
nand U4044 (N_4044,N_2684,N_2805);
or U4045 (N_4045,N_2041,N_3675);
nand U4046 (N_4046,N_3421,N_2536);
or U4047 (N_4047,N_3187,N_2405);
nand U4048 (N_4048,N_3280,N_3470);
nor U4049 (N_4049,N_3885,N_3552);
or U4050 (N_4050,N_3506,N_3038);
nor U4051 (N_4051,N_3866,N_3102);
or U4052 (N_4052,N_3154,N_2305);
or U4053 (N_4053,N_2664,N_3025);
and U4054 (N_4054,N_2209,N_2524);
nand U4055 (N_4055,N_2187,N_3821);
nor U4056 (N_4056,N_3942,N_2478);
and U4057 (N_4057,N_2154,N_2584);
and U4058 (N_4058,N_3747,N_3951);
nand U4059 (N_4059,N_2180,N_2560);
or U4060 (N_4060,N_3739,N_3580);
nor U4061 (N_4061,N_2927,N_3968);
or U4062 (N_4062,N_3435,N_3200);
xor U4063 (N_4063,N_3379,N_2260);
and U4064 (N_4064,N_3984,N_2338);
or U4065 (N_4065,N_3808,N_3558);
and U4066 (N_4066,N_2667,N_3910);
or U4067 (N_4067,N_2668,N_3817);
xnor U4068 (N_4068,N_3216,N_3055);
xnor U4069 (N_4069,N_2497,N_2779);
or U4070 (N_4070,N_3430,N_2639);
nor U4071 (N_4071,N_3936,N_2294);
or U4072 (N_4072,N_3970,N_2199);
nor U4073 (N_4073,N_3655,N_2838);
nor U4074 (N_4074,N_2889,N_3682);
and U4075 (N_4075,N_2922,N_3935);
and U4076 (N_4076,N_2892,N_3735);
xor U4077 (N_4077,N_2742,N_3969);
nand U4078 (N_4078,N_2344,N_3531);
nand U4079 (N_4079,N_3986,N_3741);
nand U4080 (N_4080,N_2329,N_3777);
nand U4081 (N_4081,N_2770,N_2984);
or U4082 (N_4082,N_2975,N_2270);
nor U4083 (N_4083,N_3472,N_3478);
or U4084 (N_4084,N_2235,N_3779);
nor U4085 (N_4085,N_3526,N_3281);
nor U4086 (N_4086,N_2098,N_2883);
and U4087 (N_4087,N_2938,N_3730);
or U4088 (N_4088,N_2500,N_3897);
xnor U4089 (N_4089,N_3431,N_2978);
or U4090 (N_4090,N_3560,N_3172);
and U4091 (N_4091,N_2352,N_2050);
and U4092 (N_4092,N_2469,N_2174);
nor U4093 (N_4093,N_3718,N_2034);
nor U4094 (N_4094,N_2404,N_2823);
or U4095 (N_4095,N_2722,N_3857);
nor U4096 (N_4096,N_2652,N_3871);
and U4097 (N_4097,N_2029,N_3246);
nor U4098 (N_4098,N_2445,N_2635);
xnor U4099 (N_4099,N_3155,N_2470);
and U4100 (N_4100,N_3151,N_3691);
nor U4101 (N_4101,N_2637,N_3294);
and U4102 (N_4102,N_2778,N_3394);
and U4103 (N_4103,N_3574,N_2241);
nor U4104 (N_4104,N_3893,N_2026);
and U4105 (N_4105,N_2509,N_3829);
nand U4106 (N_4106,N_3875,N_2909);
or U4107 (N_4107,N_2399,N_2249);
or U4108 (N_4108,N_3532,N_3310);
and U4109 (N_4109,N_3673,N_3939);
and U4110 (N_4110,N_3086,N_2256);
nand U4111 (N_4111,N_3768,N_3257);
nand U4112 (N_4112,N_3400,N_3322);
or U4113 (N_4113,N_2562,N_3818);
nor U4114 (N_4114,N_3794,N_3859);
nor U4115 (N_4115,N_2550,N_2786);
or U4116 (N_4116,N_2646,N_2946);
nor U4117 (N_4117,N_2741,N_2456);
and U4118 (N_4118,N_2616,N_3147);
or U4119 (N_4119,N_2426,N_3750);
nor U4120 (N_4120,N_2375,N_2833);
xnor U4121 (N_4121,N_3189,N_2910);
and U4122 (N_4122,N_2366,N_3649);
nand U4123 (N_4123,N_3359,N_2760);
nor U4124 (N_4124,N_3492,N_3996);
or U4125 (N_4125,N_2119,N_3567);
xor U4126 (N_4126,N_3402,N_3783);
and U4127 (N_4127,N_2649,N_2049);
nor U4128 (N_4128,N_3639,N_2554);
nor U4129 (N_4129,N_2950,N_3778);
xor U4130 (N_4130,N_2710,N_3813);
or U4131 (N_4131,N_3186,N_2755);
or U4132 (N_4132,N_2165,N_3529);
and U4133 (N_4133,N_3796,N_3111);
nor U4134 (N_4134,N_3719,N_3380);
or U4135 (N_4135,N_2401,N_3406);
nor U4136 (N_4136,N_3598,N_3021);
nand U4137 (N_4137,N_3165,N_2015);
nand U4138 (N_4138,N_2171,N_3654);
nand U4139 (N_4139,N_2611,N_2698);
nor U4140 (N_4140,N_2312,N_2377);
or U4141 (N_4141,N_2433,N_2874);
or U4142 (N_4142,N_2185,N_2683);
xor U4143 (N_4143,N_3047,N_3272);
nor U4144 (N_4144,N_2159,N_2289);
or U4145 (N_4145,N_3355,N_3923);
nand U4146 (N_4146,N_2286,N_3106);
or U4147 (N_4147,N_3895,N_2091);
or U4148 (N_4148,N_3120,N_2170);
nor U4149 (N_4149,N_2920,N_2148);
nor U4150 (N_4150,N_3301,N_3208);
or U4151 (N_4151,N_2901,N_2320);
nor U4152 (N_4152,N_2687,N_3067);
and U4153 (N_4153,N_2935,N_2085);
nand U4154 (N_4154,N_2977,N_2493);
or U4155 (N_4155,N_2854,N_3133);
nand U4156 (N_4156,N_3028,N_2781);
xnor U4157 (N_4157,N_3225,N_3125);
nand U4158 (N_4158,N_3103,N_2971);
or U4159 (N_4159,N_3037,N_3149);
nand U4160 (N_4160,N_2184,N_2864);
nand U4161 (N_4161,N_3901,N_3388);
nor U4162 (N_4162,N_3298,N_3651);
nand U4163 (N_4163,N_2557,N_2443);
nand U4164 (N_4164,N_2829,N_3722);
nand U4165 (N_4165,N_2339,N_2983);
nor U4166 (N_4166,N_3997,N_2402);
or U4167 (N_4167,N_2169,N_3925);
and U4168 (N_4168,N_2675,N_2032);
or U4169 (N_4169,N_2240,N_2578);
nor U4170 (N_4170,N_3467,N_2655);
nand U4171 (N_4171,N_2038,N_3095);
nand U4172 (N_4172,N_3156,N_2168);
nor U4173 (N_4173,N_3896,N_3934);
or U4174 (N_4174,N_2859,N_3587);
nand U4175 (N_4175,N_2737,N_3653);
nand U4176 (N_4176,N_2634,N_3306);
xor U4177 (N_4177,N_2138,N_2630);
and U4178 (N_4178,N_2725,N_3459);
nand U4179 (N_4179,N_3019,N_2832);
nor U4180 (N_4180,N_3029,N_3787);
or U4181 (N_4181,N_3792,N_2265);
and U4182 (N_4182,N_2048,N_3373);
or U4183 (N_4183,N_2113,N_2843);
and U4184 (N_4184,N_3592,N_2765);
nor U4185 (N_4185,N_2510,N_2163);
nor U4186 (N_4186,N_2886,N_2746);
or U4187 (N_4187,N_2997,N_3445);
xor U4188 (N_4188,N_2313,N_2441);
xnor U4189 (N_4189,N_2089,N_3590);
or U4190 (N_4190,N_2897,N_3677);
and U4191 (N_4191,N_2822,N_2943);
nor U4192 (N_4192,N_3305,N_3776);
and U4193 (N_4193,N_3563,N_3130);
nor U4194 (N_4194,N_2272,N_2047);
nor U4195 (N_4195,N_3692,N_3374);
xnor U4196 (N_4196,N_3076,N_2201);
xor U4197 (N_4197,N_2186,N_2821);
and U4198 (N_4198,N_3721,N_2330);
or U4199 (N_4199,N_3321,N_2237);
and U4200 (N_4200,N_2413,N_2553);
nand U4201 (N_4201,N_2880,N_3239);
xor U4202 (N_4202,N_2728,N_2274);
nor U4203 (N_4203,N_2111,N_3256);
or U4204 (N_4204,N_3457,N_2257);
nor U4205 (N_4205,N_3503,N_2852);
nor U4206 (N_4206,N_2136,N_3959);
and U4207 (N_4207,N_3898,N_3217);
or U4208 (N_4208,N_3632,N_3919);
xor U4209 (N_4209,N_3081,N_3209);
or U4210 (N_4210,N_2820,N_2143);
and U4211 (N_4211,N_3903,N_3686);
xor U4212 (N_4212,N_2112,N_3370);
or U4213 (N_4213,N_2617,N_2930);
xnor U4214 (N_4214,N_2870,N_2956);
and U4215 (N_4215,N_3279,N_2754);
and U4216 (N_4216,N_3605,N_3657);
or U4217 (N_4217,N_3284,N_3372);
and U4218 (N_4218,N_2678,N_3520);
and U4219 (N_4219,N_3364,N_2428);
nor U4220 (N_4220,N_3960,N_2198);
nor U4221 (N_4221,N_2387,N_3411);
nand U4222 (N_4222,N_2220,N_3980);
nand U4223 (N_4223,N_3058,N_3113);
nor U4224 (N_4224,N_3444,N_3150);
or U4225 (N_4225,N_2602,N_2613);
nand U4226 (N_4226,N_3108,N_3224);
and U4227 (N_4227,N_3732,N_2403);
nand U4228 (N_4228,N_2819,N_2262);
and U4229 (N_4229,N_2271,N_2979);
nor U4230 (N_4230,N_3845,N_3064);
nand U4231 (N_4231,N_3158,N_3736);
xnor U4232 (N_4232,N_2176,N_3480);
nand U4233 (N_4233,N_2110,N_3755);
and U4234 (N_4234,N_3823,N_3738);
nand U4235 (N_4235,N_3754,N_3414);
and U4236 (N_4236,N_3827,N_3625);
nor U4237 (N_4237,N_3873,N_2016);
xor U4238 (N_4238,N_3894,N_2504);
or U4239 (N_4239,N_2238,N_2000);
nor U4240 (N_4240,N_3912,N_3853);
or U4241 (N_4241,N_2083,N_3157);
and U4242 (N_4242,N_2690,N_3616);
or U4243 (N_4243,N_2847,N_2303);
or U4244 (N_4244,N_2723,N_2477);
or U4245 (N_4245,N_3589,N_2712);
and U4246 (N_4246,N_3990,N_3798);
nand U4247 (N_4247,N_2716,N_2534);
nand U4248 (N_4248,N_3035,N_3733);
nand U4249 (N_4249,N_2255,N_3769);
or U4250 (N_4250,N_3425,N_3391);
nand U4251 (N_4251,N_2783,N_3785);
xnor U4252 (N_4252,N_3879,N_2980);
xnor U4253 (N_4253,N_3698,N_3127);
or U4254 (N_4254,N_2252,N_2587);
or U4255 (N_4255,N_3293,N_3799);
nor U4256 (N_4256,N_3618,N_2431);
nor U4257 (N_4257,N_2591,N_2551);
nand U4258 (N_4258,N_3100,N_3099);
and U4259 (N_4259,N_3410,N_2985);
and U4260 (N_4260,N_2998,N_3689);
or U4261 (N_4261,N_3448,N_3326);
nor U4262 (N_4262,N_3336,N_2757);
or U4263 (N_4263,N_2435,N_3586);
nor U4264 (N_4264,N_3356,N_2654);
nand U4265 (N_4265,N_2475,N_3679);
or U4266 (N_4266,N_2498,N_2748);
nand U4267 (N_4267,N_3737,N_3123);
xor U4268 (N_4268,N_2776,N_3039);
nor U4269 (N_4269,N_3504,N_3824);
or U4270 (N_4270,N_2632,N_2989);
xnor U4271 (N_4271,N_3665,N_3114);
nor U4272 (N_4272,N_2721,N_2869);
nand U4273 (N_4273,N_3045,N_3196);
nand U4274 (N_4274,N_3170,N_3433);
nor U4275 (N_4275,N_2797,N_3027);
nor U4276 (N_4276,N_3536,N_3518);
nand U4277 (N_4277,N_2769,N_3198);
or U4278 (N_4278,N_3214,N_2005);
nor U4279 (N_4279,N_3763,N_3077);
and U4280 (N_4280,N_2014,N_3059);
or U4281 (N_4281,N_3481,N_3202);
nand U4282 (N_4282,N_3351,N_3804);
or U4283 (N_4283,N_2549,N_2628);
or U4284 (N_4284,N_3748,N_2058);
nor U4285 (N_4285,N_3191,N_3915);
nand U4286 (N_4286,N_3384,N_2590);
and U4287 (N_4287,N_3948,N_3668);
or U4288 (N_4288,N_3302,N_3704);
nand U4289 (N_4289,N_2245,N_2296);
nor U4290 (N_4290,N_3933,N_2368);
nor U4291 (N_4291,N_2348,N_2440);
nor U4292 (N_4292,N_2474,N_2659);
nand U4293 (N_4293,N_2868,N_2472);
and U4294 (N_4294,N_2100,N_3757);
and U4295 (N_4295,N_2193,N_3463);
nor U4296 (N_4296,N_3323,N_2844);
nand U4297 (N_4297,N_2853,N_3159);
and U4298 (N_4298,N_3311,N_2028);
nor U4299 (N_4299,N_3597,N_2319);
and U4300 (N_4300,N_2610,N_2693);
nor U4301 (N_4301,N_2495,N_2020);
or U4302 (N_4302,N_2968,N_3348);
and U4303 (N_4303,N_2103,N_3759);
nor U4304 (N_4304,N_2818,N_2166);
or U4305 (N_4305,N_3052,N_2127);
and U4306 (N_4306,N_3723,N_2124);
nand U4307 (N_4307,N_3498,N_2738);
or U4308 (N_4308,N_2382,N_2093);
nand U4309 (N_4309,N_2782,N_3690);
nor U4310 (N_4310,N_3703,N_3801);
xnor U4311 (N_4311,N_2814,N_3450);
or U4312 (N_4312,N_3874,N_2116);
nand U4313 (N_4313,N_3115,N_3717);
nand U4314 (N_4314,N_3429,N_3146);
nor U4315 (N_4315,N_2718,N_3485);
xor U4316 (N_4316,N_3884,N_3815);
nand U4317 (N_4317,N_3013,N_2515);
nor U4318 (N_4318,N_3510,N_3858);
nand U4319 (N_4319,N_3848,N_3017);
xor U4320 (N_4320,N_3253,N_2066);
and U4321 (N_4321,N_2809,N_3337);
and U4322 (N_4322,N_3167,N_2359);
or U4323 (N_4323,N_3088,N_3661);
or U4324 (N_4324,N_3222,N_2452);
nand U4325 (N_4325,N_2502,N_2916);
xor U4326 (N_4326,N_2799,N_2882);
nor U4327 (N_4327,N_2106,N_2134);
or U4328 (N_4328,N_2523,N_3387);
or U4329 (N_4329,N_3211,N_2307);
xor U4330 (N_4330,N_3469,N_2720);
nand U4331 (N_4331,N_3285,N_2932);
xnor U4332 (N_4332,N_2246,N_2466);
and U4333 (N_4333,N_3004,N_3631);
or U4334 (N_4334,N_3584,N_2940);
and U4335 (N_4335,N_3144,N_3927);
nand U4336 (N_4336,N_2999,N_2660);
and U4337 (N_4337,N_3206,N_3568);
and U4338 (N_4338,N_2218,N_2273);
nand U4339 (N_4339,N_2599,N_3476);
or U4340 (N_4340,N_2561,N_3188);
nand U4341 (N_4341,N_3350,N_3606);
and U4342 (N_4342,N_3867,N_3637);
or U4343 (N_4343,N_2689,N_3882);
nor U4344 (N_4344,N_3300,N_2629);
nor U4345 (N_4345,N_2161,N_3524);
xor U4346 (N_4346,N_3579,N_2115);
nand U4347 (N_4347,N_2057,N_3258);
xnor U4348 (N_4348,N_3954,N_2207);
or U4349 (N_4349,N_2327,N_3040);
or U4350 (N_4350,N_2749,N_3494);
and U4351 (N_4351,N_3118,N_3439);
or U4352 (N_4352,N_2538,N_3963);
xor U4353 (N_4353,N_2539,N_3192);
nand U4354 (N_4354,N_3343,N_2333);
xnor U4355 (N_4355,N_3325,N_3424);
nor U4356 (N_4356,N_2415,N_3036);
or U4357 (N_4357,N_3345,N_2345);
nor U4358 (N_4358,N_3385,N_2959);
xor U4359 (N_4359,N_2597,N_2045);
nor U4360 (N_4360,N_3015,N_2276);
and U4361 (N_4361,N_2640,N_3569);
nand U4362 (N_4362,N_3989,N_3521);
xor U4363 (N_4363,N_2311,N_2037);
and U4364 (N_4364,N_3877,N_3112);
nor U4365 (N_4365,N_3163,N_3810);
or U4366 (N_4366,N_2496,N_2701);
nand U4367 (N_4367,N_3193,N_3837);
nor U4368 (N_4368,N_2295,N_2644);
and U4369 (N_4369,N_2473,N_2826);
nand U4370 (N_4370,N_3352,N_3561);
or U4371 (N_4371,N_3002,N_2827);
nand U4372 (N_4372,N_3985,N_2063);
and U4373 (N_4373,N_2771,N_3595);
nor U4374 (N_4374,N_3277,N_3836);
or U4375 (N_4375,N_2577,N_2335);
nand U4376 (N_4376,N_2817,N_2266);
nor U4377 (N_4377,N_2202,N_3212);
nand U4378 (N_4378,N_2347,N_3617);
or U4379 (N_4379,N_3608,N_3807);
nor U4380 (N_4380,N_2713,N_3514);
xor U4381 (N_4381,N_3502,N_3994);
nand U4382 (N_4382,N_3409,N_3423);
and U4383 (N_4383,N_3987,N_3262);
nor U4384 (N_4384,N_3057,N_3462);
xnor U4385 (N_4385,N_3681,N_2102);
or U4386 (N_4386,N_2623,N_3443);
and U4387 (N_4387,N_2321,N_3931);
or U4388 (N_4388,N_3964,N_3880);
nor U4389 (N_4389,N_3018,N_2806);
nor U4390 (N_4390,N_2200,N_3397);
nand U4391 (N_4391,N_3454,N_3068);
xor U4392 (N_4392,N_3440,N_2356);
and U4393 (N_4393,N_2429,N_3773);
nand U4394 (N_4394,N_3628,N_2263);
nor U4395 (N_4395,N_2455,N_3138);
nor U4396 (N_4396,N_3642,N_3696);
nand U4397 (N_4397,N_3800,N_2444);
or U4398 (N_4398,N_3962,N_3864);
xnor U4399 (N_4399,N_2318,N_2866);
or U4400 (N_4400,N_3713,N_2114);
nor U4401 (N_4401,N_2691,N_3947);
or U4402 (N_4402,N_3072,N_2811);
nor U4403 (N_4403,N_3236,N_2939);
and U4404 (N_4404,N_3647,N_3338);
nand U4405 (N_4405,N_3700,N_3501);
or U4406 (N_4406,N_3447,N_3268);
and U4407 (N_4407,N_2952,N_2747);
or U4408 (N_4408,N_2494,N_3876);
or U4409 (N_4409,N_2145,N_2278);
or U4410 (N_4410,N_2314,N_2665);
nand U4411 (N_4411,N_2485,N_2899);
nand U4412 (N_4412,N_3640,N_2688);
xor U4413 (N_4413,N_3288,N_2195);
nand U4414 (N_4414,N_3244,N_3441);
and U4415 (N_4415,N_2961,N_3053);
xnor U4416 (N_4416,N_2575,N_3603);
or U4417 (N_4417,N_3797,N_2958);
or U4418 (N_4418,N_3407,N_3972);
or U4419 (N_4419,N_2288,N_3822);
or U4420 (N_4420,N_3033,N_3548);
nor U4421 (N_4421,N_2283,N_2267);
or U4422 (N_4422,N_2068,N_2316);
and U4423 (N_4423,N_2626,N_3107);
or U4424 (N_4424,N_3243,N_3060);
nor U4425 (N_4425,N_3557,N_2400);
or U4426 (N_4426,N_2964,N_2537);
nor U4427 (N_4427,N_3137,N_2357);
nor U4428 (N_4428,N_2662,N_2911);
or U4429 (N_4429,N_2324,N_3795);
xor U4430 (N_4430,N_3865,N_3263);
or U4431 (N_4431,N_3975,N_2543);
xor U4432 (N_4432,N_3816,N_3734);
or U4433 (N_4433,N_2231,N_3596);
or U4434 (N_4434,N_2379,N_3533);
and U4435 (N_4435,N_2619,N_3341);
or U4436 (N_4436,N_3839,N_2394);
nand U4437 (N_4437,N_3886,N_3255);
and U4438 (N_4438,N_2605,N_3260);
or U4439 (N_4439,N_3909,N_2842);
xnor U4440 (N_4440,N_3405,N_2846);
and U4441 (N_4441,N_3361,N_2393);
nand U4442 (N_4442,N_2371,N_3767);
nand U4443 (N_4443,N_2077,N_3803);
nor U4444 (N_4444,N_3226,N_3073);
xor U4445 (N_4445,N_3075,N_2807);
nor U4446 (N_4446,N_2601,N_3740);
or U4447 (N_4447,N_3965,N_2285);
nand U4448 (N_4448,N_3599,N_3889);
nand U4449 (N_4449,N_2604,N_3296);
and U4450 (N_4450,N_3066,N_3709);
and U4451 (N_4451,N_2593,N_2653);
or U4452 (N_4452,N_2530,N_2559);
nand U4453 (N_4453,N_2700,N_3314);
nand U4454 (N_4454,N_3054,N_3852);
nor U4455 (N_4455,N_2923,N_3645);
nor U4456 (N_4456,N_2242,N_2007);
nand U4457 (N_4457,N_3660,N_2934);
nor U4458 (N_4458,N_2603,N_3995);
and U4459 (N_4459,N_2501,N_3937);
and U4460 (N_4460,N_2099,N_3522);
xor U4461 (N_4461,N_3791,N_3334);
xnor U4462 (N_4462,N_3559,N_2419);
or U4463 (N_4463,N_3530,N_3550);
and U4464 (N_4464,N_2579,N_2904);
and U4465 (N_4465,N_3046,N_3674);
nand U4466 (N_4466,N_2881,N_3840);
nand U4467 (N_4467,N_2123,N_3535);
nor U4468 (N_4468,N_2740,N_2913);
or U4469 (N_4469,N_2759,N_2052);
and U4470 (N_4470,N_3781,N_3339);
nand U4471 (N_4471,N_3276,N_3511);
or U4472 (N_4472,N_2645,N_3953);
and U4473 (N_4473,N_2677,N_3269);
nor U4474 (N_4474,N_3184,N_2993);
or U4475 (N_4475,N_3418,N_3644);
xor U4476 (N_4476,N_2566,N_2766);
nand U4477 (N_4477,N_3327,N_2160);
xnor U4478 (N_4478,N_2837,N_3201);
and U4479 (N_4479,N_3977,N_2418);
nor U4480 (N_4480,N_3000,N_2460);
and U4481 (N_4481,N_2175,N_2606);
nor U4482 (N_4482,N_3141,N_2824);
and U4483 (N_4483,N_2558,N_2608);
nor U4484 (N_4484,N_3128,N_3612);
and U4485 (N_4485,N_2096,N_2533);
and U4486 (N_4486,N_2442,N_2043);
nor U4487 (N_4487,N_3842,N_3104);
nor U4488 (N_4488,N_2297,N_2751);
nand U4489 (N_4489,N_2081,N_3475);
xnor U4490 (N_4490,N_2078,N_3451);
or U4491 (N_4491,N_3292,N_3122);
and U4492 (N_4492,N_2526,N_2232);
and U4493 (N_4493,N_2762,N_2731);
or U4494 (N_4494,N_2830,N_2322);
and U4495 (N_4495,N_2595,N_3973);
and U4496 (N_4496,N_2370,N_2768);
xnor U4497 (N_4497,N_3929,N_2222);
nor U4498 (N_4498,N_2035,N_2795);
nor U4499 (N_4499,N_3009,N_3160);
nor U4500 (N_4500,N_3168,N_3376);
and U4501 (N_4501,N_3838,N_3638);
or U4502 (N_4502,N_2850,N_2902);
nand U4503 (N_4503,N_2407,N_2621);
nand U4504 (N_4504,N_3134,N_2073);
xor U4505 (N_4505,N_3403,N_3667);
or U4506 (N_4506,N_3868,N_3992);
or U4507 (N_4507,N_3636,N_3860);
nor U4508 (N_4508,N_3694,N_2674);
nand U4509 (N_4509,N_3274,N_3544);
or U4510 (N_4510,N_3621,N_2743);
xor U4511 (N_4511,N_3952,N_2070);
and U4512 (N_4512,N_3487,N_3979);
nor U4513 (N_4513,N_2641,N_2484);
nand U4514 (N_4514,N_2416,N_2459);
nand U4515 (N_4515,N_3164,N_2618);
nand U4516 (N_4516,N_2507,N_3266);
nand U4517 (N_4517,N_2933,N_3949);
and U4518 (N_4518,N_2293,N_2908);
or U4519 (N_4519,N_3249,N_2552);
xnor U4520 (N_4520,N_3820,N_2825);
or U4521 (N_4521,N_3684,N_2520);
and U4522 (N_4522,N_3887,N_2926);
nor U4523 (N_4523,N_2337,N_2173);
nand U4524 (N_4524,N_3482,N_2010);
and U4525 (N_4525,N_2858,N_2839);
and U4526 (N_4526,N_3540,N_2921);
nand U4527 (N_4527,N_2210,N_2421);
xor U4528 (N_4528,N_2615,N_3109);
xnor U4529 (N_4529,N_3588,N_2574);
and U4530 (N_4530,N_3219,N_2849);
nor U4531 (N_4531,N_2216,N_2620);
nand U4532 (N_4532,N_3720,N_3207);
or U4533 (N_4533,N_2929,N_3240);
or U4534 (N_4534,N_3090,N_2162);
nor U4535 (N_4535,N_3676,N_2251);
or U4536 (N_4536,N_3659,N_3050);
or U4537 (N_4537,N_2075,N_3941);
nand U4538 (N_4538,N_3899,N_3551);
nor U4539 (N_4539,N_2828,N_3378);
nand U4540 (N_4540,N_3437,N_3982);
or U4541 (N_4541,N_3371,N_2125);
xor U4542 (N_4542,N_3687,N_3085);
xor U4543 (N_4543,N_2736,N_3014);
xor U4544 (N_4544,N_2965,N_2845);
and U4545 (N_4545,N_3041,N_2009);
and U4546 (N_4546,N_2519,N_2588);
nor U4547 (N_4547,N_3140,N_2682);
and U4548 (N_4548,N_2206,N_3591);
or U4549 (N_4549,N_2600,N_3926);
nand U4550 (N_4550,N_3145,N_3347);
nand U4551 (N_4551,N_2917,N_3581);
xor U4552 (N_4552,N_2126,N_2107);
and U4553 (N_4553,N_2062,N_3474);
nand U4554 (N_4554,N_2236,N_2801);
or U4555 (N_4555,N_3252,N_3790);
or U4556 (N_4556,N_3609,N_2439);
nor U4557 (N_4557,N_3650,N_3854);
xor U4558 (N_4558,N_3863,N_2141);
and U4559 (N_4559,N_2353,N_2563);
or U4560 (N_4560,N_3515,N_3199);
and U4561 (N_4561,N_2914,N_2258);
and U4562 (N_4562,N_2522,N_2080);
or U4563 (N_4563,N_3578,N_2178);
nand U4564 (N_4564,N_2981,N_2487);
or U4565 (N_4565,N_3966,N_2006);
nand U4566 (N_4566,N_2638,N_2019);
and U4567 (N_4567,N_2960,N_2364);
nand U4568 (N_4568,N_2915,N_2571);
and U4569 (N_4569,N_2027,N_3042);
nand U4570 (N_4570,N_3920,N_2951);
and U4571 (N_4571,N_2503,N_3010);
and U4572 (N_4572,N_3758,N_3699);
nand U4573 (N_4573,N_2135,N_3319);
nand U4574 (N_4574,N_2900,N_2931);
or U4575 (N_4575,N_2212,N_3538);
and U4576 (N_4576,N_3600,N_3490);
nand U4577 (N_4577,N_3495,N_3049);
and U4578 (N_4578,N_3297,N_3507);
nand U4579 (N_4579,N_2287,N_2248);
or U4580 (N_4580,N_2018,N_3749);
nor U4581 (N_4581,N_3685,N_2894);
nand U4582 (N_4582,N_2150,N_2733);
and U4583 (N_4583,N_3819,N_2994);
nand U4584 (N_4584,N_3744,N_2957);
xor U4585 (N_4585,N_2840,N_2449);
or U4586 (N_4586,N_2264,N_3762);
nand U4587 (N_4587,N_2430,N_2476);
nand U4588 (N_4588,N_2244,N_2692);
or U4589 (N_4589,N_2205,N_3555);
nand U4590 (N_4590,N_2966,N_3043);
and U4591 (N_4591,N_3126,N_3412);
and U4592 (N_4592,N_3007,N_3627);
or U4593 (N_4593,N_2482,N_2791);
or U4594 (N_4594,N_2681,N_3945);
nor U4595 (N_4595,N_2447,N_2156);
nor U4596 (N_4596,N_2872,N_3135);
nor U4597 (N_4597,N_3404,N_3428);
or U4598 (N_4598,N_2792,N_3888);
and U4599 (N_4599,N_2082,N_3862);
nand U4600 (N_4600,N_2481,N_2417);
or U4601 (N_4601,N_2573,N_3215);
nand U4602 (N_4602,N_2545,N_3528);
or U4603 (N_4603,N_2857,N_2919);
nand U4604 (N_4604,N_2298,N_2383);
nor U4605 (N_4605,N_3183,N_3231);
or U4606 (N_4606,N_3950,N_2149);
nor U4607 (N_4607,N_2261,N_2540);
and U4608 (N_4608,N_3611,N_2188);
xnor U4609 (N_4609,N_2483,N_2315);
or U4610 (N_4610,N_2925,N_3745);
nor U4611 (N_4611,N_2179,N_3174);
or U4612 (N_4612,N_2773,N_2727);
nor U4613 (N_4613,N_2157,N_3237);
nand U4614 (N_4614,N_3971,N_3802);
nand U4615 (N_4615,N_3230,N_3093);
or U4616 (N_4616,N_3139,N_3542);
and U4617 (N_4617,N_3547,N_3166);
or U4618 (N_4618,N_3101,N_3275);
nor U4619 (N_4619,N_3782,N_2326);
or U4620 (N_4620,N_2277,N_3087);
and U4621 (N_4621,N_3786,N_2039);
nor U4622 (N_4622,N_2250,N_2717);
nor U4623 (N_4623,N_3074,N_3031);
or U4624 (N_4624,N_3583,N_2992);
nand U4625 (N_4625,N_2384,N_2309);
or U4626 (N_4626,N_2719,N_2022);
or U4627 (N_4627,N_3153,N_2409);
nor U4628 (N_4628,N_3479,N_2896);
nor U4629 (N_4629,N_2777,N_2758);
and U4630 (N_4630,N_2053,N_3978);
or U4631 (N_4631,N_3185,N_2734);
xor U4632 (N_4632,N_2453,N_3930);
nand U4633 (N_4633,N_2813,N_3026);
or U4634 (N_4634,N_2121,N_3678);
nor U4635 (N_4635,N_3295,N_3223);
or U4636 (N_4636,N_2432,N_3333);
or U4637 (N_4637,N_2967,N_2508);
nand U4638 (N_4638,N_2183,N_2622);
xnor U4639 (N_4639,N_3944,N_3291);
nand U4640 (N_4640,N_3265,N_3905);
nand U4641 (N_4641,N_2219,N_3731);
and U4642 (N_4642,N_3011,N_3413);
nand U4643 (N_4643,N_3383,N_2586);
xor U4644 (N_4644,N_2592,N_2970);
nor U4645 (N_4645,N_3916,N_3283);
nor U4646 (N_4646,N_3233,N_2358);
nand U4647 (N_4647,N_2764,N_2253);
nand U4648 (N_4648,N_2323,N_3349);
and U4649 (N_4649,N_2233,N_3344);
or U4650 (N_4650,N_2463,N_2986);
nand U4651 (N_4651,N_2529,N_2651);
and U4652 (N_4652,N_2340,N_2017);
nand U4653 (N_4653,N_2568,N_2396);
or U4654 (N_4654,N_2949,N_3248);
and U4655 (N_4655,N_2282,N_3771);
nor U4656 (N_4656,N_3051,N_3727);
nor U4657 (N_4657,N_3900,N_3726);
or U4658 (N_4658,N_3999,N_2679);
or U4659 (N_4659,N_3707,N_3911);
nor U4660 (N_4660,N_2406,N_2594);
nor U4661 (N_4661,N_2131,N_2317);
nand U4662 (N_4662,N_3641,N_2412);
and U4663 (N_4663,N_2726,N_3332);
xor U4664 (N_4664,N_2812,N_3136);
nor U4665 (N_4665,N_2750,N_2197);
nand U4666 (N_4666,N_3835,N_2877);
or U4667 (N_4667,N_2151,N_3554);
nand U4668 (N_4668,N_3282,N_3205);
nand U4669 (N_4669,N_2172,N_3643);
and U4670 (N_4670,N_3182,N_2024);
nor U4671 (N_4671,N_2424,N_2385);
nor U4672 (N_4672,N_2451,N_3855);
or U4673 (N_4673,N_2614,N_3030);
and U4674 (N_4674,N_2087,N_3020);
nor U4675 (N_4675,N_3299,N_3572);
xnor U4676 (N_4676,N_3924,N_2425);
nand U4677 (N_4677,N_3805,N_3396);
nor U4678 (N_4678,N_2567,N_3670);
xnor U4679 (N_4679,N_2702,N_3368);
or U4680 (N_4680,N_3497,N_2468);
xnor U4681 (N_4681,N_2546,N_3851);
and U4682 (N_4682,N_3575,N_3534);
and U4683 (N_4683,N_3811,N_3065);
xor U4684 (N_4684,N_3577,N_3613);
and U4685 (N_4685,N_2815,N_3921);
and U4686 (N_4686,N_2011,N_3826);
nor U4687 (N_4687,N_3213,N_2398);
and U4688 (N_4688,N_2104,N_3516);
nand U4689 (N_4689,N_3500,N_2800);
nand U4690 (N_4690,N_2855,N_2301);
nor U4691 (N_4691,N_2144,N_3446);
and U4692 (N_4692,N_2564,N_3247);
or U4693 (N_4693,N_3195,N_3220);
nand U4694 (N_4694,N_3317,N_2517);
nand U4695 (N_4695,N_2673,N_2505);
nand U4696 (N_4696,N_3615,N_2064);
nand U4697 (N_4697,N_3229,N_2890);
or U4698 (N_4698,N_2879,N_3523);
nor U4699 (N_4699,N_3377,N_2697);
nor U4700 (N_4700,N_3218,N_2450);
nor U4701 (N_4701,N_3746,N_3680);
xnor U4702 (N_4702,N_3789,N_3465);
or U4703 (N_4703,N_3708,N_3242);
and U4704 (N_4704,N_2670,N_3119);
nand U4705 (N_4705,N_3753,N_2003);
or U4706 (N_4706,N_2648,N_3286);
nand U4707 (N_4707,N_3834,N_2389);
and U4708 (N_4708,N_2281,N_2471);
nor U4709 (N_4709,N_2906,N_2972);
and U4710 (N_4710,N_2013,N_3830);
nand U4711 (N_4711,N_3728,N_3132);
nand U4712 (N_4712,N_2302,N_2040);
nor U4713 (N_4713,N_2486,N_3307);
nor U4714 (N_4714,N_3142,N_3016);
nand U4715 (N_4715,N_2669,N_3422);
xnor U4716 (N_4716,N_3398,N_2709);
or U4717 (N_4717,N_2798,N_2269);
or U4718 (N_4718,N_2204,N_2196);
nor U4719 (N_4719,N_2194,N_2774);
or U4720 (N_4720,N_3955,N_2190);
or U4721 (N_4721,N_2589,N_2438);
nand U4722 (N_4722,N_2836,N_3671);
and U4723 (N_4723,N_2873,N_2525);
or U4724 (N_4724,N_2576,N_2891);
or U4725 (N_4725,N_2065,N_3083);
nor U4726 (N_4726,N_2076,N_3991);
or U4727 (N_4727,N_2658,N_2397);
nand U4728 (N_4728,N_3071,N_2962);
and U4729 (N_4729,N_3082,N_3254);
or U4730 (N_4730,N_3711,N_2544);
nand U4731 (N_4731,N_2954,N_2023);
nand U4732 (N_4732,N_3784,N_2942);
nor U4733 (N_4733,N_2137,N_3245);
xor U4734 (N_4734,N_2753,N_3129);
and U4735 (N_4735,N_2696,N_2097);
or U4736 (N_4736,N_2275,N_2627);
and U4737 (N_4737,N_3869,N_3079);
nand U4738 (N_4738,N_3358,N_3716);
or U4739 (N_4739,N_3330,N_2213);
nand U4740 (N_4740,N_3566,N_3693);
nand U4741 (N_4741,N_3204,N_3375);
and U4742 (N_4742,N_2521,N_3190);
and U4743 (N_4743,N_2656,N_2598);
or U4744 (N_4744,N_3957,N_2056);
nor U4745 (N_4745,N_3607,N_2234);
and U4746 (N_4746,N_2875,N_2373);
nand U4747 (N_4747,N_2991,N_3981);
nor U4748 (N_4748,N_3594,N_3008);
nand U4749 (N_4749,N_2871,N_2941);
nand U4750 (N_4750,N_3324,N_3034);
or U4751 (N_4751,N_2856,N_3760);
and U4752 (N_4752,N_3148,N_2885);
nand U4753 (N_4753,N_2362,N_2512);
nand U4754 (N_4754,N_2325,N_2390);
nor U4755 (N_4755,N_3455,N_3604);
nand U4756 (N_4756,N_2350,N_3097);
or U4757 (N_4757,N_2767,N_2004);
xnor U4758 (N_4758,N_3250,N_3539);
nand U4759 (N_4759,N_3308,N_2118);
nor U4760 (N_4760,N_2848,N_2531);
or U4761 (N_4761,N_3774,N_3943);
nor U4762 (N_4762,N_3032,N_3234);
or U4763 (N_4763,N_3922,N_2247);
nor U4764 (N_4764,N_3491,N_2334);
nor U4765 (N_4765,N_3849,N_3562);
and U4766 (N_4766,N_2704,N_2528);
nand U4767 (N_4767,N_2422,N_2152);
or U4768 (N_4768,N_3271,N_3576);
nand U4769 (N_4769,N_2514,N_2306);
nor U4770 (N_4770,N_2680,N_3329);
nand U4771 (N_4771,N_2794,N_2203);
or U4772 (N_4772,N_3902,N_2328);
or U4773 (N_4773,N_3001,N_2336);
and U4774 (N_4774,N_2146,N_3369);
nand U4775 (N_4775,N_2376,N_2489);
or U4776 (N_4776,N_3362,N_2780);
xor U4777 (N_4777,N_2752,N_2414);
and U4778 (N_4778,N_3938,N_3565);
nand U4779 (N_4779,N_2192,N_2947);
nand U4780 (N_4780,N_2355,N_3289);
nand U4781 (N_4781,N_3365,N_2189);
nor U4782 (N_4782,N_3715,N_3788);
xnor U4783 (N_4783,N_2878,N_3772);
nor U4784 (N_4784,N_3382,N_3751);
or U4785 (N_4785,N_3303,N_2211);
nor U4786 (N_4786,N_2739,N_3725);
and U4787 (N_4787,N_3173,N_3505);
nor U4788 (N_4788,N_2887,N_2427);
nand U4789 (N_4789,N_3662,N_2912);
or U4790 (N_4790,N_3683,N_2793);
and U4791 (N_4791,N_2609,N_3496);
nor U4792 (N_4792,N_2128,N_3814);
or U4793 (N_4793,N_3499,N_2109);
and U4794 (N_4794,N_3084,N_2214);
or U4795 (N_4795,N_2480,N_2542);
nor U4796 (N_4796,N_2518,N_3702);
nor U4797 (N_4797,N_2071,N_3143);
or U4798 (N_4798,N_3890,N_2711);
or U4799 (N_4799,N_3360,N_2706);
xor U4800 (N_4800,N_2129,N_2724);
nor U4801 (N_4801,N_3582,N_2863);
xor U4802 (N_4802,N_2117,N_3493);
nand U4803 (N_4803,N_3564,N_2974);
and U4804 (N_4804,N_2457,N_2666);
and U4805 (N_4805,N_3328,N_3658);
or U4806 (N_4806,N_3044,N_3124);
or U4807 (N_4807,N_3417,N_2290);
nand U4808 (N_4808,N_2230,N_3235);
and U4809 (N_4809,N_3131,N_2021);
and U4810 (N_4810,N_3426,N_2243);
or U4811 (N_4811,N_3318,N_3315);
or U4812 (N_4812,N_3688,N_2488);
and U4813 (N_4813,N_3434,N_2025);
nor U4814 (N_4814,N_3466,N_2031);
and U4815 (N_4815,N_3092,N_2580);
and U4816 (N_4816,N_2945,N_2982);
nor U4817 (N_4817,N_2410,N_2672);
nand U4818 (N_4818,N_3761,N_2816);
or U4819 (N_4819,N_2079,N_2499);
and U4820 (N_4820,N_3048,N_3812);
xnor U4821 (N_4821,N_2434,N_2042);
and U4822 (N_4822,N_3780,N_2120);
and U4823 (N_4823,N_3633,N_2582);
or U4824 (N_4824,N_2069,N_3363);
nor U4825 (N_4825,N_3232,N_2239);
nor U4826 (N_4826,N_3161,N_3714);
or U4827 (N_4827,N_2454,N_3483);
and U4828 (N_4828,N_3056,N_2884);
nand U4829 (N_4829,N_3395,N_2686);
nand U4830 (N_4830,N_2732,N_3458);
or U4831 (N_4831,N_2583,N_3914);
or U4832 (N_4832,N_3408,N_2841);
or U4833 (N_4833,N_2343,N_2122);
nand U4834 (N_4834,N_3527,N_2408);
and U4835 (N_4835,N_2167,N_2944);
nand U4836 (N_4836,N_2002,N_2851);
and U4837 (N_4837,N_2105,N_3648);
and U4838 (N_4838,N_3517,N_2130);
or U4839 (N_4839,N_3841,N_3833);
nand U4840 (N_4840,N_3393,N_3389);
and U4841 (N_4841,N_2304,N_3278);
nand U4842 (N_4842,N_2995,N_3619);
nand U4843 (N_4843,N_2367,N_2555);
and U4844 (N_4844,N_3116,N_2803);
and U4845 (N_4845,N_3831,N_2067);
and U4846 (N_4846,N_3227,N_3152);
and U4847 (N_4847,N_2715,N_3453);
xor U4848 (N_4848,N_3705,N_2280);
nand U4849 (N_4849,N_2292,N_2955);
nor U4850 (N_4850,N_2217,N_3069);
and U4851 (N_4851,N_2268,N_3194);
and U4852 (N_4852,N_2625,N_3828);
nand U4853 (N_4853,N_3063,N_2585);
and U4854 (N_4854,N_2996,N_3177);
nand U4855 (N_4855,N_2108,N_3313);
or U4856 (N_4856,N_2834,N_2893);
nor U4857 (N_4857,N_3907,N_3891);
or U4858 (N_4858,N_3626,N_3180);
or U4859 (N_4859,N_3357,N_2565);
nand U4860 (N_4860,N_3367,N_2072);
nor U4861 (N_4861,N_3775,N_3974);
or U4862 (N_4862,N_2918,N_2372);
nor U4863 (N_4863,N_3171,N_3806);
nand U4864 (N_4864,N_3946,N_2458);
nor U4865 (N_4865,N_3622,N_3003);
or U4866 (N_4866,N_3908,N_2182);
nand U4867 (N_4867,N_2729,N_2090);
xor U4868 (N_4868,N_2506,N_2642);
and U4869 (N_4869,N_2860,N_2541);
nand U4870 (N_4870,N_3541,N_2363);
nand U4871 (N_4871,N_3471,N_2888);
and U4872 (N_4872,N_2378,N_3346);
nand U4873 (N_4873,N_3449,N_3203);
xnor U4874 (N_4874,N_3264,N_3416);
or U4875 (N_4875,N_2547,N_3438);
nor U4876 (N_4876,N_2527,N_3765);
xnor U4877 (N_4877,N_3913,N_3169);
nor U4878 (N_4878,N_3988,N_2423);
and U4879 (N_4879,N_3872,N_3844);
nand U4880 (N_4880,N_2036,N_3553);
or U4881 (N_4881,N_2008,N_2788);
and U4882 (N_4882,N_2569,N_3460);
xnor U4883 (N_4883,N_2225,N_2361);
nor U4884 (N_4884,N_3850,N_2059);
and U4885 (N_4885,N_2789,N_3098);
or U4886 (N_4886,N_3427,N_2744);
and U4887 (N_4887,N_3630,N_3353);
nand U4888 (N_4888,N_3917,N_2101);
nand U4889 (N_4889,N_2810,N_3956);
nor U4890 (N_4890,N_3666,N_3601);
and U4891 (N_4891,N_3270,N_2988);
nand U4892 (N_4892,N_2535,N_3706);
and U4893 (N_4893,N_2976,N_2772);
nor U4894 (N_4894,N_3585,N_2092);
and U4895 (N_4895,N_2607,N_2227);
nor U4896 (N_4896,N_2705,N_3825);
nor U4897 (N_4897,N_2215,N_3525);
nand U4898 (N_4898,N_3121,N_2572);
nor U4899 (N_4899,N_3473,N_2224);
and U4900 (N_4900,N_3181,N_2436);
and U4901 (N_4901,N_3316,N_3259);
xnor U4902 (N_4902,N_3251,N_2492);
nor U4903 (N_4903,N_3629,N_3399);
nand U4904 (N_4904,N_3484,N_3967);
or U4905 (N_4905,N_3238,N_3742);
and U4906 (N_4906,N_3634,N_3832);
or U4907 (N_4907,N_3005,N_3331);
or U4908 (N_4908,N_2570,N_2624);
xnor U4909 (N_4909,N_3546,N_2155);
nor U4910 (N_4910,N_3663,N_2802);
nand U4911 (N_4911,N_2636,N_3928);
or U4912 (N_4912,N_2462,N_3710);
or U4913 (N_4913,N_3078,N_3537);
xnor U4914 (N_4914,N_2229,N_2291);
nand U4915 (N_4915,N_3309,N_3646);
or U4916 (N_4916,N_3080,N_2133);
nor U4917 (N_4917,N_2095,N_2903);
and U4918 (N_4918,N_2532,N_3091);
nor U4919 (N_4919,N_2464,N_2647);
or U4920 (N_4920,N_3366,N_2360);
nor U4921 (N_4921,N_2707,N_2761);
nand U4922 (N_4922,N_3442,N_3695);
or U4923 (N_4923,N_3061,N_2208);
and U4924 (N_4924,N_2735,N_3096);
or U4925 (N_4925,N_2054,N_2300);
or U4926 (N_4926,N_2411,N_3468);
nor U4927 (N_4927,N_3976,N_3105);
and U4928 (N_4928,N_3415,N_3983);
nand U4929 (N_4929,N_3958,N_3175);
nor U4930 (N_4930,N_2074,N_2861);
nor U4931 (N_4931,N_3846,N_3420);
nor U4932 (N_4932,N_2835,N_3614);
and U4933 (N_4933,N_2804,N_2308);
nand U4934 (N_4934,N_3861,N_3669);
nor U4935 (N_4935,N_2374,N_2395);
xnor U4936 (N_4936,N_3519,N_3635);
and U4937 (N_4937,N_2437,N_2279);
and U4938 (N_4938,N_3883,N_3549);
nand U4939 (N_4939,N_2596,N_3070);
nand U4940 (N_4940,N_2787,N_3335);
and U4941 (N_4941,N_2055,N_2973);
nor U4942 (N_4942,N_2671,N_3486);
and U4943 (N_4943,N_2657,N_3464);
and U4944 (N_4944,N_3624,N_3024);
nand U4945 (N_4945,N_2044,N_3843);
nor U4946 (N_4946,N_3006,N_3878);
nand U4947 (N_4947,N_3770,N_2865);
nor U4948 (N_4948,N_3756,N_3456);
and U4949 (N_4949,N_2831,N_2963);
nor U4950 (N_4950,N_3545,N_3904);
nand U4951 (N_4951,N_2386,N_2775);
nand U4952 (N_4952,N_3697,N_2556);
or U4953 (N_4953,N_2341,N_3461);
nand U4954 (N_4954,N_2284,N_2346);
nand U4955 (N_4955,N_2784,N_2342);
or U4956 (N_4956,N_3906,N_2046);
nor U4957 (N_4957,N_2448,N_3401);
and U4958 (N_4958,N_2491,N_2365);
xnor U4959 (N_4959,N_2785,N_3354);
or U4960 (N_4960,N_2388,N_3961);
and U4961 (N_4961,N_3162,N_2461);
and U4962 (N_4962,N_2695,N_2479);
nand U4963 (N_4963,N_3856,N_3179);
nand U4964 (N_4964,N_3809,N_3392);
or U4965 (N_4965,N_2663,N_3932);
and U4966 (N_4966,N_2699,N_3508);
nand U4967 (N_4967,N_3571,N_3094);
nand U4968 (N_4968,N_2808,N_2221);
and U4969 (N_4969,N_2867,N_2226);
or U4970 (N_4970,N_2465,N_2876);
nor U4971 (N_4971,N_3573,N_2633);
nor U4972 (N_4972,N_3570,N_2164);
nor U4973 (N_4973,N_3881,N_2730);
xnor U4974 (N_4974,N_2140,N_3386);
or U4975 (N_4975,N_2254,N_3793);
nor U4976 (N_4976,N_3543,N_2685);
nor U4977 (N_4977,N_2990,N_2612);
and U4978 (N_4978,N_2177,N_3610);
nand U4979 (N_4979,N_3993,N_3764);
nand U4980 (N_4980,N_3512,N_2132);
nor U4981 (N_4981,N_3998,N_3489);
nor U4982 (N_4982,N_3176,N_2694);
nand U4983 (N_4983,N_3381,N_2928);
nor U4984 (N_4984,N_2139,N_3452);
and U4985 (N_4985,N_2756,N_3012);
and U4986 (N_4986,N_2490,N_2953);
and U4987 (N_4987,N_3089,N_2581);
nor U4988 (N_4988,N_2153,N_2516);
xnor U4989 (N_4989,N_3847,N_2223);
xor U4990 (N_4990,N_3320,N_3724);
nand U4991 (N_4991,N_3870,N_3892);
xor U4992 (N_4992,N_2051,N_2703);
and U4993 (N_4993,N_2898,N_2391);
nand U4994 (N_4994,N_2714,N_3273);
nor U4995 (N_4995,N_3023,N_2033);
nor U4996 (N_4996,N_3117,N_2354);
xnor U4997 (N_4997,N_3752,N_3477);
or U4998 (N_4998,N_2392,N_2708);
nand U4999 (N_4999,N_3593,N_3312);
nor U5000 (N_5000,N_3912,N_3824);
or U5001 (N_5001,N_2706,N_2446);
nand U5002 (N_5002,N_2348,N_2436);
nand U5003 (N_5003,N_2445,N_3738);
nand U5004 (N_5004,N_2417,N_2921);
or U5005 (N_5005,N_3564,N_3989);
xnor U5006 (N_5006,N_2189,N_2791);
xnor U5007 (N_5007,N_2646,N_2859);
or U5008 (N_5008,N_2819,N_2102);
nand U5009 (N_5009,N_2791,N_3569);
nand U5010 (N_5010,N_2675,N_3916);
nand U5011 (N_5011,N_3796,N_3984);
nor U5012 (N_5012,N_3257,N_2563);
and U5013 (N_5013,N_3582,N_3202);
and U5014 (N_5014,N_2513,N_2246);
xnor U5015 (N_5015,N_2609,N_3738);
and U5016 (N_5016,N_2260,N_3327);
nor U5017 (N_5017,N_2963,N_2634);
or U5018 (N_5018,N_3333,N_2649);
and U5019 (N_5019,N_2176,N_3082);
or U5020 (N_5020,N_3616,N_3209);
nand U5021 (N_5021,N_2749,N_3074);
nor U5022 (N_5022,N_3244,N_2807);
or U5023 (N_5023,N_3795,N_3629);
nand U5024 (N_5024,N_3984,N_3382);
nor U5025 (N_5025,N_3332,N_3506);
or U5026 (N_5026,N_2161,N_2811);
or U5027 (N_5027,N_2165,N_3410);
or U5028 (N_5028,N_3657,N_3778);
or U5029 (N_5029,N_3311,N_2027);
xnor U5030 (N_5030,N_3918,N_2985);
or U5031 (N_5031,N_2544,N_3133);
nor U5032 (N_5032,N_2582,N_3936);
nand U5033 (N_5033,N_2809,N_3500);
nor U5034 (N_5034,N_2270,N_3873);
xor U5035 (N_5035,N_3466,N_2183);
and U5036 (N_5036,N_2677,N_2226);
nand U5037 (N_5037,N_2049,N_2008);
nor U5038 (N_5038,N_3157,N_2738);
nand U5039 (N_5039,N_2902,N_3401);
nand U5040 (N_5040,N_2468,N_2314);
and U5041 (N_5041,N_2924,N_2021);
xor U5042 (N_5042,N_3794,N_2550);
nand U5043 (N_5043,N_3098,N_2472);
nand U5044 (N_5044,N_3982,N_2423);
and U5045 (N_5045,N_2790,N_2910);
nand U5046 (N_5046,N_2735,N_2311);
and U5047 (N_5047,N_3519,N_3099);
xor U5048 (N_5048,N_2885,N_2850);
xor U5049 (N_5049,N_3455,N_2768);
or U5050 (N_5050,N_2305,N_3089);
or U5051 (N_5051,N_2690,N_3154);
and U5052 (N_5052,N_2925,N_3983);
nor U5053 (N_5053,N_2521,N_2374);
nor U5054 (N_5054,N_3689,N_3843);
xnor U5055 (N_5055,N_3308,N_3728);
and U5056 (N_5056,N_3120,N_3515);
nor U5057 (N_5057,N_2090,N_3340);
or U5058 (N_5058,N_3486,N_3378);
nor U5059 (N_5059,N_3209,N_3174);
or U5060 (N_5060,N_2236,N_3982);
nand U5061 (N_5061,N_3284,N_2912);
nor U5062 (N_5062,N_2294,N_3996);
or U5063 (N_5063,N_3902,N_3188);
and U5064 (N_5064,N_2822,N_2654);
or U5065 (N_5065,N_3972,N_2160);
nand U5066 (N_5066,N_2079,N_3981);
and U5067 (N_5067,N_3707,N_3708);
nand U5068 (N_5068,N_2449,N_3055);
nor U5069 (N_5069,N_2010,N_2555);
nor U5070 (N_5070,N_3676,N_2271);
and U5071 (N_5071,N_2069,N_2942);
nor U5072 (N_5072,N_3358,N_3791);
or U5073 (N_5073,N_3114,N_2912);
and U5074 (N_5074,N_2825,N_3122);
xor U5075 (N_5075,N_2081,N_2519);
and U5076 (N_5076,N_3425,N_3430);
nand U5077 (N_5077,N_3191,N_2598);
xor U5078 (N_5078,N_3002,N_2341);
nand U5079 (N_5079,N_2609,N_3867);
nor U5080 (N_5080,N_2434,N_3261);
or U5081 (N_5081,N_2737,N_3805);
nor U5082 (N_5082,N_2772,N_3245);
nand U5083 (N_5083,N_3906,N_2852);
nor U5084 (N_5084,N_2193,N_3009);
nor U5085 (N_5085,N_2378,N_3357);
nor U5086 (N_5086,N_3705,N_2391);
nor U5087 (N_5087,N_2804,N_3869);
nand U5088 (N_5088,N_2703,N_3207);
or U5089 (N_5089,N_2698,N_2020);
or U5090 (N_5090,N_2420,N_2646);
nor U5091 (N_5091,N_3844,N_2690);
nand U5092 (N_5092,N_2768,N_3169);
nor U5093 (N_5093,N_2700,N_3471);
nor U5094 (N_5094,N_2915,N_3932);
and U5095 (N_5095,N_2455,N_2757);
and U5096 (N_5096,N_3410,N_3209);
nor U5097 (N_5097,N_2672,N_3252);
and U5098 (N_5098,N_2515,N_2237);
nand U5099 (N_5099,N_2840,N_3803);
nor U5100 (N_5100,N_2399,N_3609);
nor U5101 (N_5101,N_2253,N_3045);
xnor U5102 (N_5102,N_3969,N_2406);
nor U5103 (N_5103,N_3510,N_2082);
nor U5104 (N_5104,N_3397,N_3447);
nand U5105 (N_5105,N_2086,N_2548);
nor U5106 (N_5106,N_2021,N_3166);
nand U5107 (N_5107,N_3141,N_2932);
nand U5108 (N_5108,N_2687,N_3556);
or U5109 (N_5109,N_3169,N_3187);
nand U5110 (N_5110,N_3814,N_2794);
or U5111 (N_5111,N_2328,N_2433);
and U5112 (N_5112,N_2787,N_3204);
and U5113 (N_5113,N_3664,N_2945);
nand U5114 (N_5114,N_2104,N_2653);
nand U5115 (N_5115,N_3637,N_3589);
nor U5116 (N_5116,N_2920,N_2195);
or U5117 (N_5117,N_3455,N_3259);
nand U5118 (N_5118,N_2337,N_2461);
and U5119 (N_5119,N_2501,N_3496);
nand U5120 (N_5120,N_3469,N_2279);
nand U5121 (N_5121,N_2220,N_3064);
and U5122 (N_5122,N_2254,N_3946);
nor U5123 (N_5123,N_3912,N_2002);
nand U5124 (N_5124,N_2220,N_3198);
nor U5125 (N_5125,N_3146,N_3221);
or U5126 (N_5126,N_3092,N_2907);
or U5127 (N_5127,N_3615,N_2066);
nor U5128 (N_5128,N_2919,N_3010);
nor U5129 (N_5129,N_3552,N_2803);
nand U5130 (N_5130,N_2045,N_2858);
or U5131 (N_5131,N_2595,N_3265);
nand U5132 (N_5132,N_2526,N_3901);
or U5133 (N_5133,N_2671,N_3999);
or U5134 (N_5134,N_2610,N_3269);
nand U5135 (N_5135,N_2402,N_2152);
and U5136 (N_5136,N_3810,N_2572);
nor U5137 (N_5137,N_3234,N_2042);
nand U5138 (N_5138,N_3303,N_2545);
nor U5139 (N_5139,N_2231,N_2363);
nor U5140 (N_5140,N_2931,N_2670);
and U5141 (N_5141,N_2438,N_3017);
nand U5142 (N_5142,N_3134,N_3713);
xor U5143 (N_5143,N_3430,N_3882);
nand U5144 (N_5144,N_2678,N_3282);
or U5145 (N_5145,N_3250,N_2337);
nand U5146 (N_5146,N_2816,N_2455);
nor U5147 (N_5147,N_3044,N_2705);
nor U5148 (N_5148,N_2813,N_3839);
or U5149 (N_5149,N_3907,N_3969);
xor U5150 (N_5150,N_3841,N_2978);
nor U5151 (N_5151,N_3836,N_2601);
and U5152 (N_5152,N_3466,N_3443);
nand U5153 (N_5153,N_3972,N_3911);
nor U5154 (N_5154,N_3644,N_3205);
nand U5155 (N_5155,N_2637,N_3620);
nor U5156 (N_5156,N_2693,N_3437);
nand U5157 (N_5157,N_2748,N_3268);
or U5158 (N_5158,N_2610,N_2687);
or U5159 (N_5159,N_2951,N_3184);
nand U5160 (N_5160,N_2867,N_3813);
nor U5161 (N_5161,N_2292,N_2899);
xnor U5162 (N_5162,N_2974,N_2059);
nor U5163 (N_5163,N_2443,N_3010);
or U5164 (N_5164,N_2419,N_2874);
or U5165 (N_5165,N_3822,N_2385);
xnor U5166 (N_5166,N_3328,N_3994);
nand U5167 (N_5167,N_3914,N_2009);
or U5168 (N_5168,N_2899,N_2856);
nand U5169 (N_5169,N_3266,N_3253);
nand U5170 (N_5170,N_3534,N_2306);
nor U5171 (N_5171,N_2675,N_3740);
nand U5172 (N_5172,N_3369,N_3729);
and U5173 (N_5173,N_2743,N_3449);
nor U5174 (N_5174,N_2229,N_3389);
nor U5175 (N_5175,N_2069,N_3454);
and U5176 (N_5176,N_2982,N_2248);
and U5177 (N_5177,N_2671,N_3543);
xor U5178 (N_5178,N_2549,N_3906);
nor U5179 (N_5179,N_3151,N_2002);
nand U5180 (N_5180,N_3036,N_3694);
nor U5181 (N_5181,N_3212,N_3214);
and U5182 (N_5182,N_2627,N_2211);
or U5183 (N_5183,N_2305,N_3439);
and U5184 (N_5184,N_3873,N_3285);
or U5185 (N_5185,N_3548,N_2167);
nand U5186 (N_5186,N_2984,N_3308);
and U5187 (N_5187,N_3528,N_2318);
or U5188 (N_5188,N_2832,N_2848);
xor U5189 (N_5189,N_3687,N_3285);
nor U5190 (N_5190,N_2099,N_3142);
and U5191 (N_5191,N_2531,N_3778);
nand U5192 (N_5192,N_2490,N_3675);
nand U5193 (N_5193,N_3695,N_3943);
nand U5194 (N_5194,N_2587,N_2617);
nand U5195 (N_5195,N_3683,N_2094);
nand U5196 (N_5196,N_2721,N_3318);
and U5197 (N_5197,N_2760,N_2186);
xor U5198 (N_5198,N_2008,N_3079);
nor U5199 (N_5199,N_3035,N_2177);
nor U5200 (N_5200,N_3641,N_2927);
and U5201 (N_5201,N_2768,N_3134);
or U5202 (N_5202,N_2275,N_2804);
nand U5203 (N_5203,N_3126,N_2357);
or U5204 (N_5204,N_3189,N_3611);
xnor U5205 (N_5205,N_3824,N_2960);
and U5206 (N_5206,N_2152,N_2053);
and U5207 (N_5207,N_3135,N_2969);
or U5208 (N_5208,N_2080,N_2036);
nor U5209 (N_5209,N_2557,N_2908);
and U5210 (N_5210,N_2044,N_3592);
nand U5211 (N_5211,N_3972,N_3483);
nand U5212 (N_5212,N_2070,N_3484);
and U5213 (N_5213,N_2034,N_2573);
nand U5214 (N_5214,N_2522,N_2690);
nand U5215 (N_5215,N_3056,N_2647);
and U5216 (N_5216,N_2439,N_2243);
xnor U5217 (N_5217,N_2131,N_3996);
nor U5218 (N_5218,N_3145,N_3004);
and U5219 (N_5219,N_3464,N_3028);
and U5220 (N_5220,N_2466,N_3765);
and U5221 (N_5221,N_2313,N_3437);
nor U5222 (N_5222,N_3461,N_2283);
nor U5223 (N_5223,N_3349,N_3269);
or U5224 (N_5224,N_2042,N_3721);
nor U5225 (N_5225,N_3027,N_3063);
and U5226 (N_5226,N_2257,N_2774);
or U5227 (N_5227,N_3355,N_2146);
or U5228 (N_5228,N_3154,N_3560);
nor U5229 (N_5229,N_3222,N_3443);
and U5230 (N_5230,N_3572,N_3598);
or U5231 (N_5231,N_3645,N_2334);
xor U5232 (N_5232,N_2259,N_2494);
nand U5233 (N_5233,N_2560,N_2340);
or U5234 (N_5234,N_2519,N_3429);
or U5235 (N_5235,N_2970,N_3838);
nand U5236 (N_5236,N_2304,N_3142);
and U5237 (N_5237,N_2647,N_2593);
nor U5238 (N_5238,N_2600,N_2458);
nand U5239 (N_5239,N_2158,N_3417);
or U5240 (N_5240,N_2218,N_3761);
or U5241 (N_5241,N_2537,N_2283);
or U5242 (N_5242,N_2399,N_2531);
and U5243 (N_5243,N_2638,N_3887);
xor U5244 (N_5244,N_2605,N_3268);
nand U5245 (N_5245,N_2679,N_2814);
and U5246 (N_5246,N_3434,N_2920);
and U5247 (N_5247,N_3077,N_2140);
nand U5248 (N_5248,N_2057,N_2809);
nand U5249 (N_5249,N_2165,N_3129);
nor U5250 (N_5250,N_2682,N_2901);
or U5251 (N_5251,N_3751,N_3957);
nor U5252 (N_5252,N_3193,N_2443);
xnor U5253 (N_5253,N_3645,N_2474);
and U5254 (N_5254,N_2191,N_3584);
nor U5255 (N_5255,N_3418,N_3214);
or U5256 (N_5256,N_3732,N_2694);
and U5257 (N_5257,N_3201,N_3621);
and U5258 (N_5258,N_3599,N_3516);
xor U5259 (N_5259,N_3464,N_2012);
nand U5260 (N_5260,N_3824,N_2160);
or U5261 (N_5261,N_2185,N_3650);
or U5262 (N_5262,N_3932,N_2879);
xor U5263 (N_5263,N_3898,N_2228);
nand U5264 (N_5264,N_2300,N_2634);
xor U5265 (N_5265,N_2156,N_3114);
or U5266 (N_5266,N_3426,N_3271);
and U5267 (N_5267,N_2005,N_2695);
nor U5268 (N_5268,N_3130,N_3192);
or U5269 (N_5269,N_2608,N_2154);
and U5270 (N_5270,N_2226,N_2116);
nor U5271 (N_5271,N_2599,N_3331);
nand U5272 (N_5272,N_2147,N_3090);
nor U5273 (N_5273,N_2183,N_3680);
nand U5274 (N_5274,N_2255,N_2818);
nand U5275 (N_5275,N_3038,N_2247);
or U5276 (N_5276,N_2159,N_2751);
or U5277 (N_5277,N_3153,N_2897);
nand U5278 (N_5278,N_2263,N_2886);
and U5279 (N_5279,N_3799,N_3958);
and U5280 (N_5280,N_2411,N_3816);
nand U5281 (N_5281,N_2591,N_2652);
nand U5282 (N_5282,N_2548,N_3967);
or U5283 (N_5283,N_3861,N_3125);
and U5284 (N_5284,N_2347,N_3307);
and U5285 (N_5285,N_3938,N_3626);
nand U5286 (N_5286,N_3384,N_3493);
or U5287 (N_5287,N_3947,N_2055);
or U5288 (N_5288,N_2696,N_2856);
nand U5289 (N_5289,N_2351,N_3483);
nor U5290 (N_5290,N_3760,N_2249);
nand U5291 (N_5291,N_2895,N_2917);
nand U5292 (N_5292,N_2363,N_3232);
nor U5293 (N_5293,N_3618,N_3578);
xor U5294 (N_5294,N_3032,N_3899);
or U5295 (N_5295,N_2611,N_2503);
nand U5296 (N_5296,N_3931,N_2699);
nor U5297 (N_5297,N_2539,N_2903);
nand U5298 (N_5298,N_2668,N_2690);
nand U5299 (N_5299,N_2381,N_2714);
or U5300 (N_5300,N_2253,N_3137);
nand U5301 (N_5301,N_2667,N_3490);
or U5302 (N_5302,N_2239,N_2249);
and U5303 (N_5303,N_3637,N_2338);
nand U5304 (N_5304,N_2818,N_2796);
xor U5305 (N_5305,N_2172,N_3018);
nand U5306 (N_5306,N_2878,N_3629);
nor U5307 (N_5307,N_3802,N_3548);
nor U5308 (N_5308,N_2415,N_2658);
or U5309 (N_5309,N_2538,N_3189);
or U5310 (N_5310,N_3246,N_2901);
and U5311 (N_5311,N_2053,N_2541);
or U5312 (N_5312,N_2712,N_3943);
xnor U5313 (N_5313,N_3443,N_3208);
and U5314 (N_5314,N_2312,N_3145);
nor U5315 (N_5315,N_2757,N_3666);
nor U5316 (N_5316,N_3365,N_2075);
or U5317 (N_5317,N_3370,N_2966);
or U5318 (N_5318,N_3793,N_3599);
or U5319 (N_5319,N_3506,N_2271);
nor U5320 (N_5320,N_2742,N_2112);
and U5321 (N_5321,N_3231,N_3427);
nand U5322 (N_5322,N_3204,N_3198);
nand U5323 (N_5323,N_3022,N_3821);
nand U5324 (N_5324,N_3289,N_2544);
nand U5325 (N_5325,N_2364,N_2664);
nor U5326 (N_5326,N_3784,N_2628);
nor U5327 (N_5327,N_3443,N_3420);
nand U5328 (N_5328,N_3839,N_2865);
nand U5329 (N_5329,N_2585,N_2623);
or U5330 (N_5330,N_2601,N_3134);
xnor U5331 (N_5331,N_2916,N_2037);
nand U5332 (N_5332,N_2756,N_2815);
and U5333 (N_5333,N_2822,N_3397);
or U5334 (N_5334,N_3896,N_3819);
and U5335 (N_5335,N_2300,N_3554);
and U5336 (N_5336,N_2678,N_3576);
nor U5337 (N_5337,N_2412,N_3708);
xor U5338 (N_5338,N_3110,N_2374);
nor U5339 (N_5339,N_3698,N_3801);
or U5340 (N_5340,N_3206,N_3919);
and U5341 (N_5341,N_3348,N_2481);
xnor U5342 (N_5342,N_3539,N_2461);
nor U5343 (N_5343,N_2809,N_3469);
nor U5344 (N_5344,N_2155,N_3230);
nor U5345 (N_5345,N_2399,N_3953);
or U5346 (N_5346,N_2382,N_2635);
and U5347 (N_5347,N_3195,N_3849);
and U5348 (N_5348,N_2964,N_3373);
and U5349 (N_5349,N_3469,N_3939);
or U5350 (N_5350,N_3899,N_2499);
nor U5351 (N_5351,N_2813,N_3271);
and U5352 (N_5352,N_3133,N_2724);
and U5353 (N_5353,N_3491,N_3200);
xor U5354 (N_5354,N_3148,N_2305);
and U5355 (N_5355,N_2221,N_3233);
and U5356 (N_5356,N_3050,N_2189);
xor U5357 (N_5357,N_3136,N_3917);
or U5358 (N_5358,N_2870,N_3908);
and U5359 (N_5359,N_3987,N_3738);
or U5360 (N_5360,N_3695,N_2227);
nor U5361 (N_5361,N_2979,N_2946);
or U5362 (N_5362,N_2561,N_2259);
xnor U5363 (N_5363,N_3819,N_2879);
or U5364 (N_5364,N_3985,N_3553);
xor U5365 (N_5365,N_3248,N_3831);
and U5366 (N_5366,N_2367,N_3651);
nand U5367 (N_5367,N_2277,N_2394);
and U5368 (N_5368,N_2440,N_3300);
nand U5369 (N_5369,N_2136,N_3493);
or U5370 (N_5370,N_3132,N_3457);
nand U5371 (N_5371,N_3449,N_3699);
and U5372 (N_5372,N_2782,N_2944);
and U5373 (N_5373,N_2964,N_3289);
nor U5374 (N_5374,N_3579,N_3683);
nor U5375 (N_5375,N_3110,N_2669);
nand U5376 (N_5376,N_2692,N_2689);
nor U5377 (N_5377,N_2359,N_3544);
nor U5378 (N_5378,N_3087,N_3067);
xor U5379 (N_5379,N_2984,N_3824);
nor U5380 (N_5380,N_3773,N_2259);
xnor U5381 (N_5381,N_2802,N_2428);
or U5382 (N_5382,N_2278,N_3779);
nand U5383 (N_5383,N_3043,N_3500);
nor U5384 (N_5384,N_3443,N_2116);
nor U5385 (N_5385,N_3429,N_2167);
or U5386 (N_5386,N_3581,N_3977);
xnor U5387 (N_5387,N_3359,N_3441);
or U5388 (N_5388,N_2143,N_2855);
nor U5389 (N_5389,N_2849,N_2183);
or U5390 (N_5390,N_3713,N_3159);
or U5391 (N_5391,N_2982,N_3180);
and U5392 (N_5392,N_2264,N_3669);
or U5393 (N_5393,N_3845,N_3502);
nor U5394 (N_5394,N_3680,N_2302);
nor U5395 (N_5395,N_3659,N_3015);
nor U5396 (N_5396,N_2427,N_2146);
or U5397 (N_5397,N_2442,N_3262);
xor U5398 (N_5398,N_2253,N_3397);
nor U5399 (N_5399,N_3297,N_3901);
and U5400 (N_5400,N_3451,N_3137);
and U5401 (N_5401,N_3028,N_3027);
nand U5402 (N_5402,N_2887,N_2938);
nand U5403 (N_5403,N_2879,N_2369);
xor U5404 (N_5404,N_3146,N_2918);
and U5405 (N_5405,N_2017,N_2533);
nor U5406 (N_5406,N_3718,N_3460);
and U5407 (N_5407,N_3939,N_3501);
and U5408 (N_5408,N_2504,N_2070);
and U5409 (N_5409,N_2805,N_2816);
nand U5410 (N_5410,N_3809,N_3041);
nor U5411 (N_5411,N_2140,N_3254);
and U5412 (N_5412,N_2015,N_2629);
or U5413 (N_5413,N_3395,N_2219);
nor U5414 (N_5414,N_2222,N_2708);
nor U5415 (N_5415,N_3402,N_2743);
nand U5416 (N_5416,N_3240,N_3015);
nor U5417 (N_5417,N_2177,N_2633);
and U5418 (N_5418,N_3477,N_3664);
or U5419 (N_5419,N_3295,N_2862);
or U5420 (N_5420,N_2828,N_3037);
and U5421 (N_5421,N_3962,N_2240);
nand U5422 (N_5422,N_3672,N_3081);
nand U5423 (N_5423,N_3679,N_3855);
nand U5424 (N_5424,N_2057,N_2601);
or U5425 (N_5425,N_2995,N_2243);
or U5426 (N_5426,N_3817,N_2823);
xnor U5427 (N_5427,N_3801,N_2257);
or U5428 (N_5428,N_2080,N_2932);
or U5429 (N_5429,N_2972,N_3085);
nand U5430 (N_5430,N_2083,N_3110);
and U5431 (N_5431,N_3618,N_3694);
nand U5432 (N_5432,N_3724,N_2694);
or U5433 (N_5433,N_3642,N_2580);
nand U5434 (N_5434,N_3624,N_3864);
xnor U5435 (N_5435,N_3914,N_3374);
nor U5436 (N_5436,N_3434,N_3651);
and U5437 (N_5437,N_3848,N_2288);
nor U5438 (N_5438,N_3281,N_2525);
and U5439 (N_5439,N_3042,N_3852);
nor U5440 (N_5440,N_2983,N_2363);
nand U5441 (N_5441,N_2175,N_3210);
or U5442 (N_5442,N_2808,N_2046);
and U5443 (N_5443,N_2462,N_3434);
or U5444 (N_5444,N_2617,N_2746);
nor U5445 (N_5445,N_2987,N_2348);
or U5446 (N_5446,N_2158,N_2681);
nand U5447 (N_5447,N_3011,N_2007);
or U5448 (N_5448,N_2691,N_3453);
and U5449 (N_5449,N_3041,N_2456);
nand U5450 (N_5450,N_2444,N_3943);
or U5451 (N_5451,N_3367,N_3668);
or U5452 (N_5452,N_2942,N_3495);
or U5453 (N_5453,N_2665,N_2597);
nor U5454 (N_5454,N_3798,N_2140);
nor U5455 (N_5455,N_3010,N_2600);
nor U5456 (N_5456,N_2190,N_2075);
and U5457 (N_5457,N_3146,N_3616);
and U5458 (N_5458,N_2985,N_3796);
nand U5459 (N_5459,N_2899,N_3607);
nor U5460 (N_5460,N_2083,N_2345);
and U5461 (N_5461,N_3295,N_3424);
xor U5462 (N_5462,N_2785,N_2177);
nand U5463 (N_5463,N_3258,N_3323);
or U5464 (N_5464,N_2416,N_2261);
nand U5465 (N_5465,N_3779,N_3222);
and U5466 (N_5466,N_2738,N_3580);
nor U5467 (N_5467,N_2122,N_3784);
nand U5468 (N_5468,N_2533,N_2781);
nand U5469 (N_5469,N_3038,N_2335);
and U5470 (N_5470,N_3427,N_3051);
or U5471 (N_5471,N_2120,N_3880);
xor U5472 (N_5472,N_2277,N_3600);
and U5473 (N_5473,N_2112,N_3345);
nor U5474 (N_5474,N_2543,N_3067);
and U5475 (N_5475,N_3754,N_2878);
nor U5476 (N_5476,N_2605,N_2094);
and U5477 (N_5477,N_3931,N_3249);
xor U5478 (N_5478,N_2291,N_3040);
and U5479 (N_5479,N_3657,N_2296);
and U5480 (N_5480,N_2985,N_3813);
nand U5481 (N_5481,N_2768,N_3353);
nor U5482 (N_5482,N_2687,N_3390);
nand U5483 (N_5483,N_2679,N_2357);
nand U5484 (N_5484,N_2465,N_3913);
nor U5485 (N_5485,N_3286,N_2255);
xnor U5486 (N_5486,N_3818,N_2769);
and U5487 (N_5487,N_2834,N_3463);
nand U5488 (N_5488,N_2987,N_3291);
nand U5489 (N_5489,N_3475,N_2470);
and U5490 (N_5490,N_3907,N_3693);
or U5491 (N_5491,N_2744,N_3625);
and U5492 (N_5492,N_2042,N_3224);
and U5493 (N_5493,N_2231,N_2222);
and U5494 (N_5494,N_2655,N_3274);
nor U5495 (N_5495,N_3511,N_3249);
or U5496 (N_5496,N_2339,N_2328);
nand U5497 (N_5497,N_3829,N_3318);
and U5498 (N_5498,N_3409,N_3048);
nor U5499 (N_5499,N_2520,N_3149);
xnor U5500 (N_5500,N_2941,N_3657);
nor U5501 (N_5501,N_3720,N_3174);
nand U5502 (N_5502,N_2698,N_3513);
or U5503 (N_5503,N_2418,N_3886);
or U5504 (N_5504,N_2299,N_2685);
or U5505 (N_5505,N_3626,N_3928);
nor U5506 (N_5506,N_3225,N_3405);
nand U5507 (N_5507,N_3590,N_2524);
nor U5508 (N_5508,N_2394,N_2237);
or U5509 (N_5509,N_3074,N_3973);
xnor U5510 (N_5510,N_2240,N_3978);
and U5511 (N_5511,N_2438,N_2762);
nand U5512 (N_5512,N_3019,N_2157);
and U5513 (N_5513,N_2090,N_3785);
or U5514 (N_5514,N_3498,N_2311);
or U5515 (N_5515,N_2366,N_2451);
and U5516 (N_5516,N_2544,N_2470);
nor U5517 (N_5517,N_2019,N_3992);
xor U5518 (N_5518,N_3313,N_3684);
and U5519 (N_5519,N_3554,N_3804);
and U5520 (N_5520,N_3004,N_2711);
and U5521 (N_5521,N_3126,N_3413);
nor U5522 (N_5522,N_2148,N_2624);
and U5523 (N_5523,N_3015,N_2914);
and U5524 (N_5524,N_3682,N_3324);
and U5525 (N_5525,N_2665,N_2988);
nand U5526 (N_5526,N_2056,N_3751);
nor U5527 (N_5527,N_3432,N_2688);
nor U5528 (N_5528,N_3479,N_3869);
nand U5529 (N_5529,N_3136,N_3390);
or U5530 (N_5530,N_3736,N_2427);
and U5531 (N_5531,N_2394,N_2685);
nand U5532 (N_5532,N_3926,N_2647);
and U5533 (N_5533,N_2110,N_3472);
nand U5534 (N_5534,N_2249,N_2497);
and U5535 (N_5535,N_2570,N_2029);
and U5536 (N_5536,N_2271,N_3628);
and U5537 (N_5537,N_2724,N_3299);
nand U5538 (N_5538,N_3166,N_3782);
nor U5539 (N_5539,N_2785,N_3628);
and U5540 (N_5540,N_3795,N_2561);
or U5541 (N_5541,N_2101,N_2814);
nand U5542 (N_5542,N_3353,N_3117);
and U5543 (N_5543,N_2796,N_3039);
and U5544 (N_5544,N_2961,N_3493);
nand U5545 (N_5545,N_3377,N_2142);
or U5546 (N_5546,N_3218,N_2859);
or U5547 (N_5547,N_2169,N_2249);
nor U5548 (N_5548,N_3549,N_2766);
xor U5549 (N_5549,N_2543,N_3805);
nor U5550 (N_5550,N_2193,N_3655);
xor U5551 (N_5551,N_2318,N_3717);
or U5552 (N_5552,N_3559,N_2384);
xnor U5553 (N_5553,N_2840,N_3412);
and U5554 (N_5554,N_2031,N_3164);
and U5555 (N_5555,N_2908,N_3067);
nor U5556 (N_5556,N_3483,N_2621);
and U5557 (N_5557,N_2934,N_2748);
xnor U5558 (N_5558,N_3349,N_3540);
xnor U5559 (N_5559,N_3686,N_2609);
nor U5560 (N_5560,N_2395,N_3926);
or U5561 (N_5561,N_2291,N_3912);
nor U5562 (N_5562,N_3754,N_2031);
nor U5563 (N_5563,N_3361,N_3168);
nand U5564 (N_5564,N_2896,N_3297);
or U5565 (N_5565,N_2164,N_3037);
and U5566 (N_5566,N_2776,N_3808);
xnor U5567 (N_5567,N_2942,N_2391);
nor U5568 (N_5568,N_2238,N_2421);
nor U5569 (N_5569,N_2231,N_3787);
nand U5570 (N_5570,N_2183,N_2343);
nand U5571 (N_5571,N_2888,N_2569);
nor U5572 (N_5572,N_3975,N_2899);
or U5573 (N_5573,N_2680,N_3760);
nand U5574 (N_5574,N_3875,N_2710);
and U5575 (N_5575,N_3171,N_3122);
and U5576 (N_5576,N_2312,N_3076);
nand U5577 (N_5577,N_3044,N_3730);
nor U5578 (N_5578,N_2014,N_3230);
nor U5579 (N_5579,N_3625,N_3993);
nor U5580 (N_5580,N_3661,N_2399);
nor U5581 (N_5581,N_3787,N_3958);
nand U5582 (N_5582,N_2257,N_3442);
nor U5583 (N_5583,N_3691,N_2603);
or U5584 (N_5584,N_3630,N_2525);
or U5585 (N_5585,N_2189,N_3864);
or U5586 (N_5586,N_3894,N_2459);
xor U5587 (N_5587,N_2726,N_2593);
xor U5588 (N_5588,N_2091,N_2110);
and U5589 (N_5589,N_3864,N_3749);
nor U5590 (N_5590,N_2969,N_3750);
nand U5591 (N_5591,N_2878,N_2114);
and U5592 (N_5592,N_3855,N_2427);
or U5593 (N_5593,N_2095,N_3234);
nand U5594 (N_5594,N_2964,N_3065);
nor U5595 (N_5595,N_2930,N_2278);
or U5596 (N_5596,N_2608,N_2891);
or U5597 (N_5597,N_3637,N_2560);
xor U5598 (N_5598,N_2285,N_2429);
nand U5599 (N_5599,N_2537,N_2584);
nand U5600 (N_5600,N_3748,N_3001);
nand U5601 (N_5601,N_2968,N_2170);
or U5602 (N_5602,N_2854,N_3428);
and U5603 (N_5603,N_3142,N_3988);
nand U5604 (N_5604,N_3904,N_3190);
nand U5605 (N_5605,N_2140,N_3278);
and U5606 (N_5606,N_2090,N_3204);
nand U5607 (N_5607,N_2286,N_2223);
or U5608 (N_5608,N_3728,N_3578);
or U5609 (N_5609,N_3121,N_3048);
and U5610 (N_5610,N_3891,N_2533);
nor U5611 (N_5611,N_2713,N_2593);
nor U5612 (N_5612,N_2796,N_3144);
nor U5613 (N_5613,N_2257,N_2816);
or U5614 (N_5614,N_2103,N_3020);
nand U5615 (N_5615,N_2442,N_3944);
nand U5616 (N_5616,N_3200,N_2135);
or U5617 (N_5617,N_2794,N_3396);
and U5618 (N_5618,N_2776,N_3730);
nand U5619 (N_5619,N_2933,N_2224);
nor U5620 (N_5620,N_3743,N_2002);
and U5621 (N_5621,N_3187,N_3244);
or U5622 (N_5622,N_2819,N_3952);
nor U5623 (N_5623,N_2046,N_2873);
and U5624 (N_5624,N_3641,N_3735);
nand U5625 (N_5625,N_2044,N_3305);
nand U5626 (N_5626,N_3071,N_2126);
or U5627 (N_5627,N_2797,N_2676);
nor U5628 (N_5628,N_2747,N_3250);
nor U5629 (N_5629,N_3650,N_2143);
xor U5630 (N_5630,N_3274,N_2821);
nor U5631 (N_5631,N_3357,N_2224);
nor U5632 (N_5632,N_2119,N_3611);
or U5633 (N_5633,N_2066,N_2405);
nor U5634 (N_5634,N_3869,N_3581);
nor U5635 (N_5635,N_3217,N_3973);
and U5636 (N_5636,N_2539,N_3995);
nor U5637 (N_5637,N_2581,N_2818);
nor U5638 (N_5638,N_2057,N_3499);
nand U5639 (N_5639,N_3667,N_2082);
nor U5640 (N_5640,N_2303,N_2471);
or U5641 (N_5641,N_2438,N_2993);
and U5642 (N_5642,N_2508,N_2526);
nor U5643 (N_5643,N_2580,N_3870);
and U5644 (N_5644,N_2026,N_2663);
nor U5645 (N_5645,N_3318,N_3851);
or U5646 (N_5646,N_2344,N_2174);
and U5647 (N_5647,N_3609,N_2236);
nor U5648 (N_5648,N_2898,N_3442);
nand U5649 (N_5649,N_2255,N_3129);
nand U5650 (N_5650,N_2965,N_3028);
or U5651 (N_5651,N_2713,N_2947);
nand U5652 (N_5652,N_3080,N_2245);
nand U5653 (N_5653,N_2592,N_2234);
and U5654 (N_5654,N_3161,N_3449);
or U5655 (N_5655,N_2463,N_2153);
or U5656 (N_5656,N_3886,N_2550);
or U5657 (N_5657,N_3705,N_3791);
and U5658 (N_5658,N_3173,N_2511);
or U5659 (N_5659,N_2440,N_3464);
and U5660 (N_5660,N_2912,N_3682);
nand U5661 (N_5661,N_3133,N_3391);
xor U5662 (N_5662,N_3486,N_3921);
or U5663 (N_5663,N_3621,N_2362);
nand U5664 (N_5664,N_2902,N_2814);
nand U5665 (N_5665,N_3675,N_3201);
or U5666 (N_5666,N_2649,N_2067);
or U5667 (N_5667,N_2160,N_3242);
nor U5668 (N_5668,N_3889,N_3894);
and U5669 (N_5669,N_3117,N_3842);
or U5670 (N_5670,N_2164,N_2737);
nand U5671 (N_5671,N_3914,N_3220);
nor U5672 (N_5672,N_2056,N_2982);
nor U5673 (N_5673,N_3272,N_3469);
and U5674 (N_5674,N_2635,N_2638);
or U5675 (N_5675,N_3931,N_2893);
nand U5676 (N_5676,N_3223,N_3196);
nand U5677 (N_5677,N_2793,N_2608);
and U5678 (N_5678,N_3693,N_2350);
nand U5679 (N_5679,N_3780,N_3764);
and U5680 (N_5680,N_2316,N_2930);
nand U5681 (N_5681,N_2440,N_3772);
and U5682 (N_5682,N_2978,N_3781);
or U5683 (N_5683,N_2141,N_2739);
nor U5684 (N_5684,N_3487,N_3983);
and U5685 (N_5685,N_3608,N_3095);
and U5686 (N_5686,N_3837,N_2804);
nor U5687 (N_5687,N_3390,N_3129);
nor U5688 (N_5688,N_2145,N_3564);
nand U5689 (N_5689,N_2146,N_2637);
nor U5690 (N_5690,N_3994,N_2318);
nor U5691 (N_5691,N_3446,N_2190);
or U5692 (N_5692,N_3551,N_3002);
or U5693 (N_5693,N_3535,N_2462);
or U5694 (N_5694,N_3834,N_2169);
or U5695 (N_5695,N_3340,N_3127);
and U5696 (N_5696,N_2152,N_3244);
or U5697 (N_5697,N_3196,N_3494);
nor U5698 (N_5698,N_3802,N_2922);
and U5699 (N_5699,N_2040,N_3150);
or U5700 (N_5700,N_2850,N_2234);
nor U5701 (N_5701,N_3859,N_3402);
and U5702 (N_5702,N_2726,N_3898);
nand U5703 (N_5703,N_3105,N_3613);
xnor U5704 (N_5704,N_3592,N_3881);
xnor U5705 (N_5705,N_3105,N_3289);
and U5706 (N_5706,N_2729,N_3164);
or U5707 (N_5707,N_2665,N_3775);
and U5708 (N_5708,N_3619,N_2306);
and U5709 (N_5709,N_2565,N_2748);
nand U5710 (N_5710,N_3143,N_3502);
and U5711 (N_5711,N_2305,N_3663);
nand U5712 (N_5712,N_3408,N_2441);
nand U5713 (N_5713,N_2470,N_2069);
nor U5714 (N_5714,N_2090,N_2661);
or U5715 (N_5715,N_2516,N_3779);
or U5716 (N_5716,N_3291,N_3519);
nor U5717 (N_5717,N_3896,N_3494);
or U5718 (N_5718,N_2741,N_2868);
xnor U5719 (N_5719,N_2335,N_2043);
nor U5720 (N_5720,N_3865,N_3702);
and U5721 (N_5721,N_2378,N_3685);
and U5722 (N_5722,N_3250,N_3430);
nor U5723 (N_5723,N_2259,N_3169);
xor U5724 (N_5724,N_3938,N_2821);
nand U5725 (N_5725,N_3505,N_3756);
xor U5726 (N_5726,N_2867,N_2263);
nor U5727 (N_5727,N_3643,N_3726);
and U5728 (N_5728,N_3672,N_3445);
or U5729 (N_5729,N_3362,N_2078);
nand U5730 (N_5730,N_3073,N_2974);
xor U5731 (N_5731,N_2803,N_3528);
or U5732 (N_5732,N_3772,N_3130);
and U5733 (N_5733,N_3434,N_2835);
nor U5734 (N_5734,N_2320,N_2401);
or U5735 (N_5735,N_2530,N_2426);
and U5736 (N_5736,N_3328,N_3333);
or U5737 (N_5737,N_2860,N_2639);
nand U5738 (N_5738,N_3346,N_2802);
or U5739 (N_5739,N_3629,N_2746);
or U5740 (N_5740,N_3380,N_3122);
nand U5741 (N_5741,N_2266,N_3624);
nand U5742 (N_5742,N_2165,N_2102);
nor U5743 (N_5743,N_2128,N_3969);
or U5744 (N_5744,N_2489,N_2353);
nand U5745 (N_5745,N_3821,N_3503);
or U5746 (N_5746,N_3918,N_3143);
or U5747 (N_5747,N_3356,N_3479);
and U5748 (N_5748,N_2333,N_2327);
or U5749 (N_5749,N_2077,N_3617);
and U5750 (N_5750,N_3210,N_3708);
nand U5751 (N_5751,N_2865,N_2788);
nand U5752 (N_5752,N_3204,N_3174);
and U5753 (N_5753,N_3576,N_2650);
and U5754 (N_5754,N_3439,N_2005);
nand U5755 (N_5755,N_2613,N_3921);
nor U5756 (N_5756,N_2948,N_2545);
and U5757 (N_5757,N_3629,N_2604);
or U5758 (N_5758,N_2112,N_2972);
or U5759 (N_5759,N_2687,N_2505);
nand U5760 (N_5760,N_2417,N_2933);
nor U5761 (N_5761,N_3364,N_3971);
and U5762 (N_5762,N_2648,N_2545);
or U5763 (N_5763,N_2186,N_2074);
nand U5764 (N_5764,N_2611,N_3005);
or U5765 (N_5765,N_2262,N_3164);
xnor U5766 (N_5766,N_2725,N_3092);
or U5767 (N_5767,N_2765,N_3167);
and U5768 (N_5768,N_2655,N_2272);
xnor U5769 (N_5769,N_3178,N_3565);
nand U5770 (N_5770,N_3210,N_3389);
and U5771 (N_5771,N_3802,N_2103);
nand U5772 (N_5772,N_3550,N_2713);
and U5773 (N_5773,N_2349,N_3352);
and U5774 (N_5774,N_3813,N_3613);
nor U5775 (N_5775,N_3921,N_3980);
and U5776 (N_5776,N_2181,N_3101);
or U5777 (N_5777,N_2421,N_2810);
and U5778 (N_5778,N_3094,N_3972);
and U5779 (N_5779,N_3012,N_3837);
xor U5780 (N_5780,N_3174,N_2500);
nand U5781 (N_5781,N_2538,N_3102);
and U5782 (N_5782,N_2402,N_2753);
nor U5783 (N_5783,N_3609,N_2469);
xor U5784 (N_5784,N_2756,N_2269);
or U5785 (N_5785,N_2225,N_3488);
nor U5786 (N_5786,N_3179,N_2822);
and U5787 (N_5787,N_3585,N_3498);
and U5788 (N_5788,N_2034,N_2390);
and U5789 (N_5789,N_2908,N_2221);
nand U5790 (N_5790,N_3947,N_3870);
nand U5791 (N_5791,N_2618,N_2226);
or U5792 (N_5792,N_3337,N_3945);
or U5793 (N_5793,N_2933,N_3572);
nor U5794 (N_5794,N_2091,N_3574);
nor U5795 (N_5795,N_3420,N_3686);
nand U5796 (N_5796,N_2709,N_3279);
or U5797 (N_5797,N_2317,N_3936);
and U5798 (N_5798,N_2851,N_3857);
nor U5799 (N_5799,N_3389,N_2464);
nor U5800 (N_5800,N_3316,N_2358);
xnor U5801 (N_5801,N_3797,N_2461);
or U5802 (N_5802,N_3156,N_3187);
and U5803 (N_5803,N_3747,N_2959);
or U5804 (N_5804,N_2172,N_3806);
nor U5805 (N_5805,N_3140,N_3772);
or U5806 (N_5806,N_2857,N_3893);
or U5807 (N_5807,N_3004,N_2325);
or U5808 (N_5808,N_3437,N_3501);
nor U5809 (N_5809,N_3253,N_2622);
or U5810 (N_5810,N_3632,N_3223);
nand U5811 (N_5811,N_3371,N_2109);
nor U5812 (N_5812,N_2512,N_3996);
or U5813 (N_5813,N_2089,N_2670);
xnor U5814 (N_5814,N_3094,N_3750);
or U5815 (N_5815,N_3649,N_2906);
xnor U5816 (N_5816,N_3889,N_2660);
and U5817 (N_5817,N_2810,N_2412);
and U5818 (N_5818,N_2089,N_2550);
nor U5819 (N_5819,N_3622,N_3322);
or U5820 (N_5820,N_3829,N_2648);
and U5821 (N_5821,N_2567,N_2865);
or U5822 (N_5822,N_2499,N_2397);
or U5823 (N_5823,N_2625,N_2650);
or U5824 (N_5824,N_3376,N_2778);
and U5825 (N_5825,N_2780,N_2578);
nand U5826 (N_5826,N_3397,N_2370);
and U5827 (N_5827,N_3715,N_3713);
and U5828 (N_5828,N_2519,N_2556);
nand U5829 (N_5829,N_3649,N_3530);
nand U5830 (N_5830,N_3870,N_2125);
nor U5831 (N_5831,N_3085,N_2828);
xnor U5832 (N_5832,N_2034,N_3938);
nor U5833 (N_5833,N_3305,N_2829);
or U5834 (N_5834,N_2189,N_3925);
nor U5835 (N_5835,N_2968,N_3541);
nand U5836 (N_5836,N_3122,N_2777);
or U5837 (N_5837,N_2414,N_2891);
nor U5838 (N_5838,N_2982,N_3942);
nand U5839 (N_5839,N_3649,N_3875);
and U5840 (N_5840,N_3383,N_2086);
nor U5841 (N_5841,N_2702,N_3365);
nand U5842 (N_5842,N_2292,N_3567);
and U5843 (N_5843,N_2031,N_3137);
nand U5844 (N_5844,N_3004,N_2578);
nor U5845 (N_5845,N_3317,N_3137);
nor U5846 (N_5846,N_3313,N_2940);
nor U5847 (N_5847,N_2138,N_2795);
and U5848 (N_5848,N_2295,N_2240);
and U5849 (N_5849,N_2903,N_3534);
xor U5850 (N_5850,N_2855,N_2603);
xor U5851 (N_5851,N_2800,N_2809);
xor U5852 (N_5852,N_3214,N_2645);
and U5853 (N_5853,N_2250,N_3675);
or U5854 (N_5854,N_2928,N_3393);
nor U5855 (N_5855,N_2737,N_2096);
xnor U5856 (N_5856,N_3030,N_2443);
and U5857 (N_5857,N_2988,N_3997);
or U5858 (N_5858,N_3240,N_2506);
nand U5859 (N_5859,N_2433,N_3783);
nor U5860 (N_5860,N_2004,N_2355);
or U5861 (N_5861,N_2934,N_3072);
and U5862 (N_5862,N_3238,N_2550);
nand U5863 (N_5863,N_2081,N_3814);
and U5864 (N_5864,N_3900,N_3589);
nor U5865 (N_5865,N_2304,N_3195);
nand U5866 (N_5866,N_2947,N_3215);
and U5867 (N_5867,N_2339,N_3802);
and U5868 (N_5868,N_3757,N_2857);
and U5869 (N_5869,N_3049,N_3507);
xnor U5870 (N_5870,N_2694,N_3909);
xor U5871 (N_5871,N_3113,N_2223);
nand U5872 (N_5872,N_2076,N_3645);
or U5873 (N_5873,N_2414,N_3071);
or U5874 (N_5874,N_2033,N_2369);
and U5875 (N_5875,N_2000,N_3711);
and U5876 (N_5876,N_2653,N_2128);
or U5877 (N_5877,N_3878,N_2070);
nor U5878 (N_5878,N_2868,N_2408);
nor U5879 (N_5879,N_3835,N_3154);
nand U5880 (N_5880,N_2906,N_3271);
or U5881 (N_5881,N_3050,N_3185);
nand U5882 (N_5882,N_3951,N_3960);
and U5883 (N_5883,N_2844,N_3776);
xnor U5884 (N_5884,N_3054,N_3845);
nand U5885 (N_5885,N_2924,N_2608);
and U5886 (N_5886,N_3327,N_3968);
or U5887 (N_5887,N_3513,N_2253);
xnor U5888 (N_5888,N_3640,N_2365);
nor U5889 (N_5889,N_3530,N_3427);
or U5890 (N_5890,N_3224,N_2586);
or U5891 (N_5891,N_2690,N_2922);
nor U5892 (N_5892,N_2955,N_2699);
xnor U5893 (N_5893,N_2665,N_3132);
or U5894 (N_5894,N_2167,N_2254);
nor U5895 (N_5895,N_3556,N_2674);
and U5896 (N_5896,N_2510,N_3707);
nor U5897 (N_5897,N_3735,N_2128);
xnor U5898 (N_5898,N_2630,N_2478);
and U5899 (N_5899,N_3992,N_2629);
xor U5900 (N_5900,N_2646,N_2272);
nand U5901 (N_5901,N_3792,N_3872);
and U5902 (N_5902,N_2111,N_3924);
nor U5903 (N_5903,N_2868,N_2274);
nor U5904 (N_5904,N_2629,N_3521);
and U5905 (N_5905,N_3121,N_2289);
or U5906 (N_5906,N_3894,N_2373);
or U5907 (N_5907,N_2155,N_2548);
and U5908 (N_5908,N_3260,N_2404);
and U5909 (N_5909,N_2366,N_3482);
nand U5910 (N_5910,N_3758,N_3087);
xor U5911 (N_5911,N_3554,N_3147);
nand U5912 (N_5912,N_2532,N_3147);
or U5913 (N_5913,N_3875,N_2028);
and U5914 (N_5914,N_3650,N_2930);
and U5915 (N_5915,N_3142,N_3923);
nor U5916 (N_5916,N_3036,N_3426);
nand U5917 (N_5917,N_2126,N_2400);
nor U5918 (N_5918,N_2764,N_2814);
nor U5919 (N_5919,N_2766,N_2138);
nand U5920 (N_5920,N_3240,N_2366);
and U5921 (N_5921,N_3923,N_2377);
and U5922 (N_5922,N_3387,N_3429);
and U5923 (N_5923,N_3955,N_3651);
or U5924 (N_5924,N_2202,N_3144);
xor U5925 (N_5925,N_2206,N_2422);
nand U5926 (N_5926,N_3497,N_2865);
or U5927 (N_5927,N_2837,N_3428);
nand U5928 (N_5928,N_3197,N_2938);
or U5929 (N_5929,N_2805,N_2141);
nor U5930 (N_5930,N_2552,N_3894);
nand U5931 (N_5931,N_3941,N_2957);
nor U5932 (N_5932,N_2698,N_3643);
nand U5933 (N_5933,N_2985,N_3371);
nand U5934 (N_5934,N_2240,N_2770);
and U5935 (N_5935,N_3738,N_3471);
or U5936 (N_5936,N_2268,N_3965);
or U5937 (N_5937,N_2593,N_3389);
or U5938 (N_5938,N_3779,N_3378);
or U5939 (N_5939,N_2614,N_3804);
or U5940 (N_5940,N_3673,N_3506);
nor U5941 (N_5941,N_2181,N_3977);
or U5942 (N_5942,N_2827,N_2077);
nand U5943 (N_5943,N_3616,N_2310);
nor U5944 (N_5944,N_3318,N_3344);
and U5945 (N_5945,N_2095,N_2768);
nand U5946 (N_5946,N_2692,N_2306);
or U5947 (N_5947,N_2181,N_3002);
nand U5948 (N_5948,N_2521,N_2916);
or U5949 (N_5949,N_3560,N_3898);
nand U5950 (N_5950,N_3121,N_3175);
nand U5951 (N_5951,N_2368,N_2126);
nand U5952 (N_5952,N_3629,N_2369);
or U5953 (N_5953,N_2573,N_3224);
nor U5954 (N_5954,N_2686,N_2258);
nor U5955 (N_5955,N_2700,N_3004);
nand U5956 (N_5956,N_2670,N_3023);
and U5957 (N_5957,N_2476,N_2127);
nand U5958 (N_5958,N_3028,N_3862);
or U5959 (N_5959,N_2012,N_3797);
nand U5960 (N_5960,N_2279,N_3036);
nand U5961 (N_5961,N_3519,N_3214);
nand U5962 (N_5962,N_3737,N_2696);
nand U5963 (N_5963,N_2130,N_3765);
nor U5964 (N_5964,N_2289,N_3165);
xnor U5965 (N_5965,N_3584,N_3762);
nand U5966 (N_5966,N_3170,N_3199);
xnor U5967 (N_5967,N_3780,N_2688);
xor U5968 (N_5968,N_2964,N_3571);
and U5969 (N_5969,N_2697,N_3347);
or U5970 (N_5970,N_3690,N_3382);
and U5971 (N_5971,N_2908,N_3822);
or U5972 (N_5972,N_2428,N_3345);
nand U5973 (N_5973,N_3530,N_3455);
nand U5974 (N_5974,N_2827,N_3206);
xor U5975 (N_5975,N_3271,N_2019);
nor U5976 (N_5976,N_3551,N_2017);
and U5977 (N_5977,N_3085,N_3538);
and U5978 (N_5978,N_2615,N_3589);
nand U5979 (N_5979,N_3751,N_3091);
or U5980 (N_5980,N_2380,N_3194);
and U5981 (N_5981,N_3128,N_2710);
nor U5982 (N_5982,N_3680,N_2380);
and U5983 (N_5983,N_3009,N_3760);
and U5984 (N_5984,N_2419,N_3004);
or U5985 (N_5985,N_2264,N_3053);
or U5986 (N_5986,N_2924,N_3275);
and U5987 (N_5987,N_2998,N_3052);
nor U5988 (N_5988,N_3093,N_2407);
nand U5989 (N_5989,N_3422,N_2773);
nand U5990 (N_5990,N_3696,N_3788);
xor U5991 (N_5991,N_3639,N_3028);
and U5992 (N_5992,N_3734,N_3580);
and U5993 (N_5993,N_3997,N_3321);
or U5994 (N_5994,N_2840,N_3052);
nand U5995 (N_5995,N_2486,N_3403);
nor U5996 (N_5996,N_2975,N_2389);
nor U5997 (N_5997,N_3682,N_2654);
and U5998 (N_5998,N_2831,N_2741);
nor U5999 (N_5999,N_3879,N_3684);
and U6000 (N_6000,N_4090,N_4366);
nor U6001 (N_6001,N_5077,N_5605);
and U6002 (N_6002,N_5143,N_4442);
or U6003 (N_6003,N_5619,N_5924);
or U6004 (N_6004,N_5758,N_4082);
or U6005 (N_6005,N_4353,N_5005);
nor U6006 (N_6006,N_5611,N_4563);
or U6007 (N_6007,N_4581,N_5125);
nor U6008 (N_6008,N_5505,N_4264);
nor U6009 (N_6009,N_5108,N_4315);
or U6010 (N_6010,N_4232,N_4772);
or U6011 (N_6011,N_4673,N_5399);
nand U6012 (N_6012,N_4964,N_5989);
nor U6013 (N_6013,N_5579,N_4074);
nor U6014 (N_6014,N_4378,N_4329);
nor U6015 (N_6015,N_5227,N_4922);
nand U6016 (N_6016,N_5095,N_5506);
nand U6017 (N_6017,N_4101,N_5603);
nand U6018 (N_6018,N_5326,N_4534);
nor U6019 (N_6019,N_5219,N_4761);
xnor U6020 (N_6020,N_5766,N_5024);
nor U6021 (N_6021,N_5297,N_4757);
nand U6022 (N_6022,N_5867,N_5244);
or U6023 (N_6023,N_4413,N_4499);
nor U6024 (N_6024,N_5713,N_5952);
nor U6025 (N_6025,N_4991,N_5184);
or U6026 (N_6026,N_5870,N_4094);
and U6027 (N_6027,N_4398,N_4656);
nand U6028 (N_6028,N_4619,N_5463);
and U6029 (N_6029,N_5013,N_5616);
nor U6030 (N_6030,N_4701,N_4115);
and U6031 (N_6031,N_5906,N_5478);
nor U6032 (N_6032,N_5567,N_5073);
nor U6033 (N_6033,N_4308,N_5654);
or U6034 (N_6034,N_5601,N_4351);
or U6035 (N_6035,N_5561,N_5979);
nor U6036 (N_6036,N_4405,N_4186);
or U6037 (N_6037,N_5759,N_4750);
xnor U6038 (N_6038,N_4356,N_5753);
nand U6039 (N_6039,N_5522,N_4244);
nand U6040 (N_6040,N_5688,N_4902);
and U6041 (N_6041,N_4173,N_5599);
and U6042 (N_6042,N_4475,N_4859);
or U6043 (N_6043,N_5692,N_4560);
nor U6044 (N_6044,N_5813,N_4763);
and U6045 (N_6045,N_5784,N_5763);
or U6046 (N_6046,N_5846,N_4609);
nor U6047 (N_6047,N_4449,N_5205);
nand U6048 (N_6048,N_5332,N_5464);
nor U6049 (N_6049,N_4660,N_5173);
xor U6050 (N_6050,N_5221,N_4272);
nand U6051 (N_6051,N_5861,N_4259);
or U6052 (N_6052,N_4995,N_4128);
or U6053 (N_6053,N_4179,N_5771);
nand U6054 (N_6054,N_5600,N_4407);
nand U6055 (N_6055,N_5944,N_5899);
and U6056 (N_6056,N_5860,N_5613);
nand U6057 (N_6057,N_5290,N_4450);
or U6058 (N_6058,N_4374,N_5903);
or U6059 (N_6059,N_4337,N_4939);
or U6060 (N_6060,N_5090,N_4530);
and U6061 (N_6061,N_4169,N_5345);
nand U6062 (N_6062,N_4154,N_5652);
or U6063 (N_6063,N_4292,N_4565);
xnor U6064 (N_6064,N_5696,N_4429);
nand U6065 (N_6065,N_4759,N_5118);
nand U6066 (N_6066,N_4219,N_5527);
xor U6067 (N_6067,N_4228,N_5637);
or U6068 (N_6068,N_4009,N_4653);
or U6069 (N_6069,N_5590,N_4392);
nand U6070 (N_6070,N_4735,N_4994);
nand U6071 (N_6071,N_5953,N_5190);
nand U6072 (N_6072,N_5974,N_4057);
nor U6073 (N_6073,N_4233,N_4410);
nand U6074 (N_6074,N_5673,N_5859);
nand U6075 (N_6075,N_4391,N_4835);
or U6076 (N_6076,N_4175,N_4245);
xor U6077 (N_6077,N_4302,N_5355);
or U6078 (N_6078,N_4016,N_4503);
nor U6079 (N_6079,N_4976,N_4348);
nand U6080 (N_6080,N_4945,N_4506);
nand U6081 (N_6081,N_4171,N_4519);
or U6082 (N_6082,N_4388,N_4222);
nand U6083 (N_6083,N_5742,N_4849);
nand U6084 (N_6084,N_4526,N_4518);
or U6085 (N_6085,N_4202,N_4040);
nand U6086 (N_6086,N_5514,N_5727);
nand U6087 (N_6087,N_4806,N_4580);
xor U6088 (N_6088,N_4185,N_5946);
xor U6089 (N_6089,N_5341,N_4894);
nor U6090 (N_6090,N_4345,N_4980);
nor U6091 (N_6091,N_5700,N_4646);
nand U6092 (N_6092,N_5898,N_5553);
and U6093 (N_6093,N_4961,N_5820);
xnor U6094 (N_6094,N_5022,N_5206);
xor U6095 (N_6095,N_5307,N_5113);
and U6096 (N_6096,N_4797,N_4114);
or U6097 (N_6097,N_4816,N_4511);
nand U6098 (N_6098,N_4866,N_4411);
nand U6099 (N_6099,N_4088,N_4042);
and U6100 (N_6100,N_5398,N_4212);
or U6101 (N_6101,N_5035,N_4958);
nand U6102 (N_6102,N_4885,N_4397);
or U6103 (N_6103,N_4722,N_4294);
and U6104 (N_6104,N_5680,N_4531);
or U6105 (N_6105,N_4313,N_4711);
or U6106 (N_6106,N_4207,N_4118);
nand U6107 (N_6107,N_5292,N_4149);
nand U6108 (N_6108,N_5550,N_4102);
nor U6109 (N_6109,N_5558,N_4028);
or U6110 (N_6110,N_5214,N_5381);
and U6111 (N_6111,N_5996,N_4886);
nor U6112 (N_6112,N_4807,N_4617);
and U6113 (N_6113,N_4936,N_4390);
nand U6114 (N_6114,N_5897,N_5793);
nand U6115 (N_6115,N_4818,N_4923);
xnor U6116 (N_6116,N_5009,N_5854);
or U6117 (N_6117,N_5481,N_4645);
nor U6118 (N_6118,N_5490,N_5783);
nand U6119 (N_6119,N_5821,N_5280);
xnor U6120 (N_6120,N_4508,N_5644);
nor U6121 (N_6121,N_5177,N_4963);
or U6122 (N_6122,N_5155,N_5299);
xnor U6123 (N_6123,N_4256,N_4426);
or U6124 (N_6124,N_4003,N_5532);
nand U6125 (N_6125,N_4664,N_4780);
nor U6126 (N_6126,N_5352,N_5656);
nand U6127 (N_6127,N_5218,N_4109);
or U6128 (N_6128,N_5868,N_5123);
and U6129 (N_6129,N_5126,N_4472);
nor U6130 (N_6130,N_5698,N_5706);
xnor U6131 (N_6131,N_4672,N_5800);
nand U6132 (N_6132,N_4605,N_4596);
nor U6133 (N_6133,N_5811,N_5887);
nand U6134 (N_6134,N_5919,N_4239);
nor U6135 (N_6135,N_4196,N_4773);
or U6136 (N_6136,N_4822,N_5675);
nand U6137 (N_6137,N_5195,N_4817);
and U6138 (N_6138,N_5866,N_4384);
nor U6139 (N_6139,N_5995,N_4748);
nand U6140 (N_6140,N_5436,N_4685);
nand U6141 (N_6141,N_4273,N_5954);
nand U6142 (N_6142,N_5740,N_5395);
and U6143 (N_6143,N_4951,N_5083);
nand U6144 (N_6144,N_4968,N_5743);
nand U6145 (N_6145,N_4703,N_4791);
nor U6146 (N_6146,N_5520,N_5094);
nand U6147 (N_6147,N_5351,N_5098);
and U6148 (N_6148,N_4373,N_4485);
nand U6149 (N_6149,N_4121,N_5283);
nand U6150 (N_6150,N_5911,N_5955);
and U6151 (N_6151,N_5138,N_5294);
or U6152 (N_6152,N_5962,N_5229);
nor U6153 (N_6153,N_4015,N_4423);
nand U6154 (N_6154,N_4532,N_5255);
or U6155 (N_6155,N_5267,N_5468);
and U6156 (N_6156,N_5382,N_5327);
nor U6157 (N_6157,N_4227,N_5609);
nor U6158 (N_6158,N_4887,N_5477);
nor U6159 (N_6159,N_4238,N_5862);
or U6160 (N_6160,N_5140,N_5475);
and U6161 (N_6161,N_5818,N_4547);
and U6162 (N_6162,N_4896,N_4744);
nand U6163 (N_6163,N_5983,N_5548);
nor U6164 (N_6164,N_4970,N_5985);
nor U6165 (N_6165,N_5970,N_5980);
xnor U6166 (N_6166,N_4269,N_4971);
nand U6167 (N_6167,N_5792,N_4717);
and U6168 (N_6168,N_4068,N_4357);
or U6169 (N_6169,N_4035,N_4603);
nand U6170 (N_6170,N_5354,N_4151);
nand U6171 (N_6171,N_5650,N_5245);
nand U6172 (N_6172,N_5466,N_5281);
and U6173 (N_6173,N_4361,N_4721);
xor U6174 (N_6174,N_4837,N_4047);
nand U6175 (N_6175,N_4841,N_4303);
nor U6176 (N_6176,N_4176,N_5660);
and U6177 (N_6177,N_5856,N_5316);
nand U6178 (N_6178,N_5851,N_4104);
nor U6179 (N_6179,N_5358,N_4189);
xor U6180 (N_6180,N_5390,N_4811);
and U6181 (N_6181,N_5584,N_5836);
nand U6182 (N_6182,N_5422,N_4898);
nor U6183 (N_6183,N_4507,N_4138);
and U6184 (N_6184,N_5757,N_4274);
nor U6185 (N_6185,N_5342,N_4631);
or U6186 (N_6186,N_4350,N_5849);
or U6187 (N_6187,N_4793,N_5623);
or U6188 (N_6188,N_4174,N_5444);
or U6189 (N_6189,N_5699,N_5006);
or U6190 (N_6190,N_4237,N_4871);
xor U6191 (N_6191,N_4172,N_4576);
nand U6192 (N_6192,N_5804,N_4979);
nand U6193 (N_6193,N_5088,N_5470);
nand U6194 (N_6194,N_4640,N_4081);
nand U6195 (N_6195,N_4491,N_4786);
or U6196 (N_6196,N_5391,N_4824);
and U6197 (N_6197,N_5701,N_5032);
and U6198 (N_6198,N_5936,N_4271);
xor U6199 (N_6199,N_5581,N_4462);
and U6200 (N_6200,N_5314,N_5311);
and U6201 (N_6201,N_4572,N_5597);
nand U6202 (N_6202,N_4714,N_4105);
nand U6203 (N_6203,N_5751,N_5797);
or U6204 (N_6204,N_5714,N_5693);
and U6205 (N_6205,N_4328,N_4952);
nor U6206 (N_6206,N_5993,N_5659);
and U6207 (N_6207,N_5106,N_4493);
nor U6208 (N_6208,N_4826,N_4247);
and U6209 (N_6209,N_4144,N_5423);
nor U6210 (N_6210,N_5272,N_4771);
or U6211 (N_6211,N_4086,N_4062);
or U6212 (N_6212,N_5614,N_4148);
nor U6213 (N_6213,N_4064,N_5733);
nor U6214 (N_6214,N_4095,N_5394);
or U6215 (N_6215,N_4665,N_4908);
nor U6216 (N_6216,N_5511,N_5872);
and U6217 (N_6217,N_4589,N_5932);
and U6218 (N_6218,N_5193,N_5356);
nand U6219 (N_6219,N_4561,N_4451);
nand U6220 (N_6220,N_5164,N_5990);
and U6221 (N_6221,N_5238,N_5034);
xor U6222 (N_6222,N_5641,N_4000);
xnor U6223 (N_6223,N_5869,N_5788);
nor U6224 (N_6224,N_4467,N_5149);
nor U6225 (N_6225,N_5072,N_5796);
nor U6226 (N_6226,N_5521,N_5273);
and U6227 (N_6227,N_5829,N_5531);
and U6228 (N_6228,N_5662,N_5877);
or U6229 (N_6229,N_4632,N_4891);
nand U6230 (N_6230,N_4260,N_5460);
or U6231 (N_6231,N_4618,N_4119);
or U6232 (N_6232,N_4371,N_5883);
nand U6233 (N_6233,N_5051,N_5384);
nand U6234 (N_6234,N_5669,N_5334);
nand U6235 (N_6235,N_5596,N_5534);
xor U6236 (N_6236,N_4844,N_4008);
and U6237 (N_6237,N_5837,N_5257);
or U6238 (N_6238,N_4027,N_4320);
nor U6239 (N_6239,N_4550,N_4856);
nand U6240 (N_6240,N_5943,N_4488);
nand U6241 (N_6241,N_4928,N_5428);
and U6242 (N_6242,N_4687,N_4395);
nand U6243 (N_6243,N_4882,N_4428);
and U6244 (N_6244,N_4156,N_5805);
and U6245 (N_6245,N_4498,N_5594);
and U6246 (N_6246,N_4230,N_4682);
and U6247 (N_6247,N_4728,N_4986);
and U6248 (N_6248,N_5170,N_5554);
and U6249 (N_6249,N_4425,N_4539);
nand U6250 (N_6250,N_4178,N_4624);
xor U6251 (N_6251,N_4033,N_4677);
nand U6252 (N_6252,N_5949,N_5808);
nand U6253 (N_6253,N_4610,N_5144);
or U6254 (N_6254,N_5736,N_5730);
and U6255 (N_6255,N_5201,N_4076);
nand U6256 (N_6256,N_4180,N_5902);
xnor U6257 (N_6257,N_5920,N_5237);
or U6258 (N_6258,N_5573,N_4988);
or U6259 (N_6259,N_5528,N_5535);
and U6260 (N_6260,N_4892,N_5159);
or U6261 (N_6261,N_5055,N_5810);
or U6262 (N_6262,N_5657,N_5066);
nor U6263 (N_6263,N_5518,N_4688);
nand U6264 (N_6264,N_4990,N_4888);
nand U6265 (N_6265,N_4385,N_5031);
nand U6266 (N_6266,N_5529,N_4681);
and U6267 (N_6267,N_5212,N_4341);
and U6268 (N_6268,N_5449,N_4203);
nand U6269 (N_6269,N_4683,N_5541);
nand U6270 (N_6270,N_4235,N_4920);
nor U6271 (N_6271,N_4497,N_4344);
or U6272 (N_6272,N_5779,N_5973);
nor U6273 (N_6273,N_4365,N_5588);
and U6274 (N_6274,N_4045,N_4020);
nand U6275 (N_6275,N_5152,N_5265);
nand U6276 (N_6276,N_5415,N_4433);
nand U6277 (N_6277,N_5402,N_4279);
and U6278 (N_6278,N_5674,N_5277);
or U6279 (N_6279,N_5411,N_4133);
nor U6280 (N_6280,N_4085,N_4782);
nand U6281 (N_6281,N_5064,N_5141);
and U6282 (N_6282,N_4134,N_5617);
nand U6283 (N_6283,N_5723,N_4960);
or U6284 (N_6284,N_5647,N_5412);
or U6285 (N_6285,N_4661,N_5802);
nand U6286 (N_6286,N_5117,N_5270);
or U6287 (N_6287,N_4715,N_5293);
or U6288 (N_6288,N_5653,N_5357);
nand U6289 (N_6289,N_4324,N_4457);
or U6290 (N_6290,N_4477,N_5348);
nor U6291 (N_6291,N_5110,N_4868);
nand U6292 (N_6292,N_4443,N_5719);
or U6293 (N_6293,N_5089,N_4860);
nor U6294 (N_6294,N_4049,N_4827);
and U6295 (N_6295,N_4460,N_5480);
or U6296 (N_6296,N_4608,N_5430);
or U6297 (N_6297,N_4018,N_5069);
nor U6298 (N_6298,N_5695,N_5607);
and U6299 (N_6299,N_5947,N_4476);
and U6300 (N_6300,N_5775,N_4774);
nand U6301 (N_6301,N_4043,N_4766);
or U6302 (N_6302,N_4347,N_5582);
nor U6303 (N_6303,N_5732,N_5204);
nand U6304 (N_6304,N_4162,N_5180);
or U6305 (N_6305,N_5340,N_5798);
or U6306 (N_6306,N_5366,N_4921);
nor U6307 (N_6307,N_4249,N_5023);
or U6308 (N_6308,N_5000,N_5927);
xor U6309 (N_6309,N_4730,N_5183);
nor U6310 (N_6310,N_4193,N_4283);
or U6311 (N_6311,N_5703,N_5426);
or U6312 (N_6312,N_4097,N_4427);
nand U6313 (N_6313,N_4358,N_5433);
and U6314 (N_6314,N_4157,N_5879);
and U6315 (N_6315,N_5039,N_4041);
and U6316 (N_6316,N_5991,N_5346);
nand U6317 (N_6317,N_5377,N_5344);
or U6318 (N_6318,N_5044,N_4335);
nor U6319 (N_6319,N_5216,N_4767);
nand U6320 (N_6320,N_5543,N_5418);
and U6321 (N_6321,N_5574,N_5217);
or U6322 (N_6322,N_5645,N_4599);
and U6323 (N_6323,N_4087,N_4931);
nand U6324 (N_6324,N_5258,N_5365);
or U6325 (N_6325,N_4103,N_5857);
or U6326 (N_6326,N_5078,N_5547);
nor U6327 (N_6327,N_4117,N_4517);
and U6328 (N_6328,N_5852,N_5410);
nand U6329 (N_6329,N_5835,N_4598);
xor U6330 (N_6330,N_4557,N_5047);
nor U6331 (N_6331,N_5592,N_5658);
nor U6332 (N_6332,N_5296,N_4832);
and U6333 (N_6333,N_4808,N_5233);
or U6334 (N_6334,N_4368,N_5665);
nand U6335 (N_6335,N_4977,N_4216);
xnor U6336 (N_6336,N_4326,N_5571);
nor U6337 (N_6337,N_4742,N_5003);
nand U6338 (N_6338,N_5263,N_5266);
nor U6339 (N_6339,N_4510,N_5969);
nand U6340 (N_6340,N_4819,N_5168);
or U6341 (N_6341,N_4456,N_5538);
or U6342 (N_6342,N_4342,N_4304);
or U6343 (N_6343,N_4708,N_5323);
nand U6344 (N_6344,N_4336,N_5832);
xor U6345 (N_6345,N_4267,N_5071);
and U6346 (N_6346,N_4039,N_4635);
or U6347 (N_6347,N_4270,N_5997);
nor U6348 (N_6348,N_5011,N_4718);
nor U6349 (N_6349,N_5303,N_4501);
and U6350 (N_6350,N_4593,N_5812);
nor U6351 (N_6351,N_4323,N_5685);
or U6352 (N_6352,N_5838,N_4288);
or U6353 (N_6353,N_5087,N_5749);
nor U6354 (N_6354,N_5101,N_5400);
xnor U6355 (N_6355,N_5577,N_5228);
or U6356 (N_6356,N_5819,N_5814);
nor U6357 (N_6357,N_5236,N_4402);
nor U6358 (N_6358,N_5642,N_5112);
nand U6359 (N_6359,N_4438,N_4876);
or U6360 (N_6360,N_5729,N_5151);
nor U6361 (N_6361,N_5530,N_5994);
and U6362 (N_6362,N_4762,N_4845);
nor U6363 (N_6363,N_4083,N_4021);
nand U6364 (N_6364,N_4248,N_5791);
xor U6365 (N_6365,N_5509,N_4355);
nor U6366 (N_6366,N_4224,N_4933);
or U6367 (N_6367,N_5492,N_5200);
nand U6368 (N_6368,N_5278,N_4291);
and U6369 (N_6369,N_4437,N_5794);
and U6370 (N_6370,N_5199,N_5350);
and U6371 (N_6371,N_4556,N_4017);
xor U6372 (N_6372,N_5904,N_4719);
xor U6373 (N_6373,N_5191,N_5586);
nand U6374 (N_6374,N_5157,N_5568);
xnor U6375 (N_6375,N_4419,N_5604);
nand U6376 (N_6376,N_5122,N_5526);
or U6377 (N_6377,N_4627,N_4712);
or U6378 (N_6378,N_4551,N_5499);
xnor U6379 (N_6379,N_5968,N_5431);
or U6380 (N_6380,N_4187,N_4192);
xor U6381 (N_6381,N_5459,N_5304);
or U6382 (N_6382,N_4959,N_5376);
nand U6383 (N_6383,N_4482,N_5343);
nand U6384 (N_6384,N_4091,N_4657);
nor U6385 (N_6385,N_4025,N_5655);
nor U6386 (N_6386,N_4604,N_4246);
and U6387 (N_6387,N_4658,N_5153);
and U6388 (N_6388,N_4465,N_4536);
or U6389 (N_6389,N_5720,N_5638);
and U6390 (N_6390,N_5401,N_4676);
nand U6391 (N_6391,N_4883,N_5361);
or U6392 (N_6392,N_5243,N_5926);
xnor U6393 (N_6393,N_4542,N_5930);
nor U6394 (N_6394,N_5145,N_5682);
and U6395 (N_6395,N_4300,N_5052);
nor U6396 (N_6396,N_4029,N_5171);
nand U6397 (N_6397,N_4842,N_4515);
nand U6398 (N_6398,N_5606,N_5891);
nor U6399 (N_6399,N_5487,N_4792);
or U6400 (N_6400,N_5407,N_5785);
nand U6401 (N_6401,N_5131,N_4622);
xnor U6402 (N_6402,N_5918,N_5049);
xor U6403 (N_6403,N_4236,N_5300);
nand U6404 (N_6404,N_5182,N_4521);
or U6405 (N_6405,N_4843,N_5964);
or U6406 (N_6406,N_4798,N_4597);
and U6407 (N_6407,N_5988,N_4127);
and U6408 (N_6408,N_5754,N_5100);
nand U6409 (N_6409,N_5239,N_4092);
nor U6410 (N_6410,N_4785,N_4299);
nor U6411 (N_6411,N_4112,N_5485);
xor U6412 (N_6412,N_4862,N_5065);
nand U6413 (N_6413,N_5709,N_4700);
nor U6414 (N_6414,N_4654,N_4191);
nor U6415 (N_6415,N_5331,N_5322);
nand U6416 (N_6416,N_5246,N_5062);
nor U6417 (N_6417,N_5678,N_4639);
or U6418 (N_6418,N_5416,N_4295);
and U6419 (N_6419,N_4258,N_5724);
nor U6420 (N_6420,N_5166,N_4559);
nor U6421 (N_6421,N_5916,N_5546);
and U6422 (N_6422,N_4689,N_4644);
xnor U6423 (N_6423,N_5830,N_5704);
and U6424 (N_6424,N_5938,N_5747);
or U6425 (N_6425,N_5711,N_5012);
and U6426 (N_6426,N_5396,N_4659);
nand U6427 (N_6427,N_4571,N_4120);
or U6428 (N_6428,N_5080,N_5959);
and U6429 (N_6429,N_4881,N_4743);
nand U6430 (N_6430,N_5315,N_4825);
and U6431 (N_6431,N_4974,N_4403);
and U6432 (N_6432,N_5484,N_5172);
nor U6433 (N_6433,N_4099,N_5374);
nor U6434 (N_6434,N_5050,N_5276);
and U6435 (N_6435,N_4732,N_4067);
and U6436 (N_6436,N_4387,N_4929);
nand U6437 (N_6437,N_4549,N_4197);
and U6438 (N_6438,N_4278,N_5824);
nor U6439 (N_6439,N_4409,N_4864);
or U6440 (N_6440,N_4434,N_5163);
or U6441 (N_6441,N_5963,N_5741);
nand U6442 (N_6442,N_5966,N_4481);
and U6443 (N_6443,N_5556,N_4814);
nor U6444 (N_6444,N_5441,N_5207);
nor U6445 (N_6445,N_4445,N_5461);
nand U6446 (N_6446,N_5765,N_4975);
nand U6447 (N_6447,N_4262,N_5096);
or U6448 (N_6448,N_4590,N_4194);
nand U6449 (N_6449,N_5386,N_5786);
and U6450 (N_6450,N_5271,N_4254);
or U6451 (N_6451,N_5542,N_5807);
and U6452 (N_6452,N_4394,N_5620);
xnor U6453 (N_6453,N_4261,N_5249);
and U6454 (N_6454,N_4006,N_5458);
and U6455 (N_6455,N_4878,N_4367);
nand U6456 (N_6456,N_5687,N_5670);
nor U6457 (N_6457,N_5847,N_4932);
and U6458 (N_6458,N_4901,N_4486);
or U6459 (N_6459,N_5027,N_4126);
nand U6460 (N_6460,N_5942,N_5683);
nor U6461 (N_6461,N_4470,N_5795);
nor U6462 (N_6462,N_5744,N_5211);
nand U6463 (N_6463,N_4496,N_4552);
xnor U6464 (N_6464,N_5465,N_4788);
or U6465 (N_6465,N_4854,N_5137);
and U6466 (N_6466,N_4587,N_5907);
and U6467 (N_6467,N_5774,N_4381);
nand U6468 (N_6468,N_4941,N_5443);
or U6469 (N_6469,N_4048,N_5893);
nand U6470 (N_6470,N_5222,N_4217);
nor U6471 (N_6471,N_5998,N_5309);
or U6472 (N_6472,N_5482,N_4877);
or U6473 (N_6473,N_4942,N_5651);
or U6474 (N_6474,N_4838,N_5397);
nor U6475 (N_6475,N_5439,N_5372);
and U6476 (N_6476,N_5923,N_4399);
or U6477 (N_6477,N_4430,N_5841);
nor U6478 (N_6478,N_5434,N_5473);
and U6479 (N_6479,N_5640,N_4492);
nor U6480 (N_6480,N_5984,N_4143);
or U6481 (N_6481,N_5777,N_4161);
nand U6482 (N_6482,N_5892,N_4023);
nand U6483 (N_6483,N_4543,N_4024);
or U6484 (N_6484,N_5941,N_4787);
nor U6485 (N_6485,N_4240,N_5301);
or U6486 (N_6486,N_4012,N_5259);
or U6487 (N_6487,N_5209,N_4606);
nor U6488 (N_6488,N_4206,N_4781);
nor U6489 (N_6489,N_4795,N_4641);
or U6490 (N_6490,N_4937,N_5583);
nor U6491 (N_6491,N_4828,N_4211);
and U6492 (N_6492,N_5451,N_4875);
nor U6493 (N_6493,N_4312,N_5677);
and U6494 (N_6494,N_4541,N_5362);
nand U6495 (N_6495,N_4764,N_5223);
nor U6496 (N_6496,N_5068,N_5612);
xor U6497 (N_6497,N_4679,N_4981);
and U6498 (N_6498,N_5148,N_4626);
xnor U6499 (N_6499,N_4564,N_4046);
and U6500 (N_6500,N_5070,N_5587);
nor U6501 (N_6501,N_5565,N_5540);
or U6502 (N_6502,N_5076,N_4113);
and U6503 (N_6503,N_4935,N_4452);
nand U6504 (N_6504,N_5746,N_4123);
nor U6505 (N_6505,N_5524,N_4965);
nand U6506 (N_6506,N_4284,N_4075);
xnor U6507 (N_6507,N_5663,N_5544);
nand U6508 (N_6508,N_5756,N_4625);
nand U6509 (N_6509,N_5092,N_5578);
and U6510 (N_6510,N_5773,N_5186);
and U6511 (N_6511,N_4967,N_4796);
nor U6512 (N_6512,N_4642,N_4803);
and U6513 (N_6513,N_4812,N_4544);
and U6514 (N_6514,N_5737,N_5452);
and U6515 (N_6515,N_4418,N_4918);
nor U6516 (N_6516,N_4513,N_4277);
nor U6517 (N_6517,N_4802,N_4504);
nand U6518 (N_6518,N_5103,N_4904);
nand U6519 (N_6519,N_4070,N_4516);
or U6520 (N_6520,N_5863,N_4372);
nand U6521 (N_6521,N_5053,N_4648);
nand U6522 (N_6522,N_4301,N_5728);
and U6523 (N_6523,N_4032,N_5018);
or U6524 (N_6524,N_5510,N_5373);
or U6525 (N_6525,N_4383,N_4415);
or U6526 (N_6526,N_5371,N_5901);
nor U6527 (N_6527,N_4066,N_5162);
nor U6528 (N_6528,N_4989,N_4184);
and U6529 (N_6529,N_4458,N_5406);
and U6530 (N_6530,N_4674,N_5387);
nor U6531 (N_6531,N_5133,N_4110);
and U6532 (N_6532,N_5445,N_5215);
or U6533 (N_6533,N_5147,N_5254);
or U6534 (N_6534,N_5636,N_4997);
nand U6535 (N_6535,N_4234,N_4753);
or U6536 (N_6536,N_5427,N_5282);
xnor U6537 (N_6537,N_4140,N_5250);
and U6538 (N_6538,N_5033,N_5150);
or U6539 (N_6539,N_4690,N_4364);
nand U6540 (N_6540,N_5956,N_4713);
nand U6541 (N_6541,N_4160,N_4215);
and U6542 (N_6542,N_5041,N_4139);
nand U6543 (N_6543,N_5462,N_5850);
nor U6544 (N_6544,N_5745,N_4870);
or U6545 (N_6545,N_4930,N_4737);
and U6546 (N_6546,N_5404,N_5099);
and U6547 (N_6547,N_5085,N_4480);
nand U6548 (N_6548,N_4890,N_5825);
nor U6549 (N_6549,N_5982,N_4698);
nor U6550 (N_6550,N_4809,N_4071);
or U6551 (N_6551,N_5232,N_4170);
and U6552 (N_6552,N_5776,N_4494);
and U6553 (N_6553,N_5718,N_5061);
nor U6554 (N_6554,N_4266,N_4111);
nor U6555 (N_6555,N_5189,N_5888);
xor U6556 (N_6556,N_4389,N_4582);
xnor U6557 (N_6557,N_5324,N_4691);
nor U6558 (N_6558,N_4694,N_5336);
or U6559 (N_6559,N_4448,N_4984);
or U6560 (N_6560,N_4073,N_5248);
nand U6561 (N_6561,N_5417,N_5871);
xor U6562 (N_6562,N_5648,N_4600);
nor U6563 (N_6563,N_5353,N_4836);
and U6564 (N_6564,N_5450,N_4080);
nor U6565 (N_6565,N_4463,N_4897);
nor U6566 (N_6566,N_5909,N_5210);
or U6567 (N_6567,N_5202,N_5536);
or U6568 (N_6568,N_4408,N_5127);
nand U6569 (N_6569,N_5501,N_5457);
xnor U6570 (N_6570,N_4296,N_5067);
and U6571 (N_6571,N_4833,N_5317);
and U6572 (N_6572,N_4416,N_5306);
or U6573 (N_6573,N_5537,N_4122);
nor U6574 (N_6574,N_5500,N_4276);
nand U6575 (N_6575,N_5102,N_5516);
nand U6576 (N_6576,N_5684,N_5921);
and U6577 (N_6577,N_4079,N_4281);
or U6578 (N_6578,N_5338,N_5555);
nand U6579 (N_6579,N_4054,N_5424);
nor U6580 (N_6580,N_4400,N_4540);
nor U6581 (N_6581,N_4242,N_4943);
xor U6582 (N_6582,N_5562,N_4727);
or U6583 (N_6583,N_4096,N_4950);
and U6584 (N_6584,N_4848,N_5935);
xnor U6585 (N_6585,N_4725,N_4620);
nand U6586 (N_6586,N_4765,N_5933);
nand U6587 (N_6587,N_4089,N_4310);
and U6588 (N_6588,N_4693,N_5119);
nand U6589 (N_6589,N_4574,N_5945);
xnor U6590 (N_6590,N_4545,N_5632);
nand U6591 (N_6591,N_5816,N_5764);
nor U6592 (N_6592,N_5885,N_5021);
and U6593 (N_6593,N_5497,N_4915);
or U6594 (N_6594,N_4327,N_4483);
nand U6595 (N_6595,N_4275,N_4478);
or U6596 (N_6596,N_4268,N_4243);
nor U6597 (N_6597,N_5716,N_5036);
nand U6598 (N_6598,N_5347,N_4436);
and U6599 (N_6599,N_5030,N_4340);
and U6600 (N_6600,N_4314,N_4699);
or U6601 (N_6601,N_5513,N_5799);
nand U6602 (N_6602,N_4252,N_4790);
xor U6603 (N_6603,N_4223,N_4570);
nor U6604 (N_6604,N_4061,N_4583);
nor U6605 (N_6605,N_5999,N_5486);
and U6606 (N_6606,N_4846,N_4421);
and U6607 (N_6607,N_4910,N_5261);
xor U6608 (N_6608,N_4804,N_4037);
and U6609 (N_6609,N_5016,N_4716);
or U6610 (N_6610,N_4962,N_4982);
xor U6611 (N_6611,N_5330,N_5697);
and U6612 (N_6612,N_5010,N_5975);
xor U6613 (N_6613,N_5557,N_4459);
or U6614 (N_6614,N_4629,N_4591);
or U6615 (N_6615,N_4810,N_4778);
or U6616 (N_6616,N_5672,N_5922);
and U6617 (N_6617,N_4829,N_4022);
nor U6618 (N_6618,N_5624,N_5054);
xor U6619 (N_6619,N_4607,N_5167);
nand U6620 (N_6620,N_5875,N_4198);
nand U6621 (N_6621,N_4575,N_5978);
nor U6622 (N_6622,N_5158,N_5889);
nor U6623 (N_6623,N_4704,N_4396);
nor U6624 (N_6624,N_4137,N_5169);
or U6625 (N_6625,N_4038,N_5840);
nor U6626 (N_6626,N_4649,N_4229);
and U6627 (N_6627,N_4741,N_4821);
nor U6628 (N_6628,N_4996,N_4905);
and U6629 (N_6629,N_4731,N_4509);
nor U6630 (N_6630,N_4053,N_5447);
and U6631 (N_6631,N_4758,N_4720);
or U6632 (N_6632,N_5972,N_5681);
or U6633 (N_6633,N_4695,N_5007);
nor U6634 (N_6634,N_5308,N_5735);
and U6635 (N_6635,N_4853,N_4188);
nand U6636 (N_6636,N_5337,N_4668);
xor U6637 (N_6637,N_4615,N_5048);
and U6638 (N_6638,N_4406,N_4051);
xnor U6639 (N_6639,N_5413,N_4740);
nor U6640 (N_6640,N_4132,N_4265);
or U6641 (N_6641,N_4473,N_5801);
and U6642 (N_6642,N_5312,N_5086);
nand U6643 (N_6643,N_4471,N_4424);
or U6644 (N_6644,N_5251,N_4663);
nand U6645 (N_6645,N_5392,N_4455);
or U6646 (N_6646,N_4709,N_4895);
nor U6647 (N_6647,N_4056,N_5895);
nand U6648 (N_6648,N_5380,N_5161);
xor U6649 (N_6649,N_5507,N_4055);
nor U6650 (N_6650,N_4966,N_4004);
or U6651 (N_6651,N_4621,N_5175);
or U6652 (N_6652,N_5806,N_4538);
nand U6653 (N_6653,N_4623,N_4760);
and U6654 (N_6654,N_5987,N_4005);
xor U6655 (N_6655,N_4142,N_5625);
or U6656 (N_6656,N_5408,N_4464);
or U6657 (N_6657,N_4613,N_4044);
and U6658 (N_6658,N_4783,N_5865);
or U6659 (N_6659,N_4359,N_5453);
and U6660 (N_6660,N_5738,N_4146);
xnor U6661 (N_6661,N_4669,N_5967);
xnor U6662 (N_6662,N_4059,N_4052);
nor U6663 (N_6663,N_5363,N_5734);
and U6664 (N_6664,N_4072,N_5074);
and U6665 (N_6665,N_5057,N_5762);
nor U6666 (N_6666,N_4584,N_4321);
nor U6667 (N_6667,N_4857,N_4562);
or U6668 (N_6668,N_4777,N_5707);
or U6669 (N_6669,N_4333,N_4667);
nor U6670 (N_6670,N_4872,N_4749);
and U6671 (N_6671,N_5960,N_5174);
and U6672 (N_6672,N_5679,N_5004);
nand U6673 (N_6673,N_5178,N_4177);
and U6674 (N_6674,N_5726,N_4680);
and U6675 (N_6675,N_5002,N_5873);
and U6676 (N_6676,N_4221,N_4724);
nor U6677 (N_6677,N_5593,N_4447);
or U6678 (N_6678,N_4282,N_5627);
nand U6679 (N_6679,N_4010,N_4370);
nand U6680 (N_6680,N_5634,N_4461);
or U6681 (N_6681,N_4490,N_4671);
nor U6682 (N_6682,N_4001,N_5671);
nand U6683 (N_6683,N_5772,N_4141);
and U6684 (N_6684,N_4190,N_4729);
or U6685 (N_6685,N_5313,N_5855);
or U6686 (N_6686,N_4263,N_5780);
xor U6687 (N_6687,N_5185,N_4697);
and U6688 (N_6688,N_5971,N_5559);
nand U6689 (N_6689,N_4537,N_5442);
and U6690 (N_6690,N_5843,N_4352);
nand U6691 (N_6691,N_5639,N_5105);
and U6692 (N_6692,N_4289,N_5748);
nor U6693 (N_6693,N_5708,N_5950);
or U6694 (N_6694,N_5213,N_4647);
nor U6695 (N_6695,N_4136,N_4241);
and U6696 (N_6696,N_4666,N_4734);
or U6697 (N_6697,N_4938,N_4573);
nor U6698 (N_6698,N_4058,N_4992);
nor U6699 (N_6699,N_5479,N_4723);
nand U6700 (N_6700,N_5136,N_4946);
nor U6701 (N_6701,N_4339,N_5104);
and U6702 (N_6702,N_5360,N_4469);
nor U6703 (N_6703,N_4325,N_5114);
and U6704 (N_6704,N_4985,N_4726);
nor U6705 (N_6705,N_5325,N_4948);
and U6706 (N_6706,N_5197,N_5121);
nand U6707 (N_6707,N_4745,N_4776);
nand U6708 (N_6708,N_4290,N_4514);
or U6709 (N_6709,N_5437,N_5284);
xor U6710 (N_6710,N_5498,N_5752);
and U6711 (N_6711,N_5474,N_4874);
or U6712 (N_6712,N_5815,N_4919);
nor U6713 (N_6713,N_5710,N_5389);
nor U6714 (N_6714,N_5414,N_5512);
nor U6715 (N_6715,N_4678,N_4354);
xnor U6716 (N_6716,N_5285,N_4949);
or U6717 (N_6717,N_5809,N_5690);
or U6718 (N_6718,N_4401,N_5508);
nand U6719 (N_6719,N_4850,N_4675);
xor U6720 (N_6720,N_4611,N_5042);
and U6721 (N_6721,N_4555,N_5881);
or U6722 (N_6722,N_5635,N_5549);
nor U6723 (N_6723,N_4746,N_4225);
nand U6724 (N_6724,N_5469,N_4911);
or U6725 (N_6725,N_4546,N_5517);
or U6726 (N_6726,N_4655,N_4906);
or U6727 (N_6727,N_5705,N_5425);
nand U6728 (N_6728,N_5038,N_5664);
and U6729 (N_6729,N_4019,N_5992);
nor U6730 (N_6730,N_5196,N_4026);
xnor U6731 (N_6731,N_4739,N_4643);
nand U6732 (N_6732,N_5302,N_4375);
or U6733 (N_6733,N_4286,N_4209);
or U6734 (N_6734,N_5194,N_5234);
and U6735 (N_6735,N_5598,N_5502);
nor U6736 (N_6736,N_4998,N_5483);
or U6737 (N_6737,N_4567,N_5181);
and U6738 (N_6738,N_5731,N_5493);
nor U6739 (N_6739,N_4393,N_4441);
and U6740 (N_6740,N_4250,N_4338);
or U6741 (N_6741,N_5712,N_4914);
nand U6742 (N_6742,N_4414,N_4612);
and U6743 (N_6743,N_4955,N_4889);
nand U6744 (N_6744,N_4130,N_4297);
nor U6745 (N_6745,N_4331,N_5977);
nor U6746 (N_6746,N_4684,N_4034);
or U6747 (N_6747,N_5310,N_4311);
and U6748 (N_6748,N_4084,N_4852);
nand U6749 (N_6749,N_5160,N_4349);
xor U6750 (N_6750,N_4322,N_4050);
or U6751 (N_6751,N_4893,N_4226);
nand U6752 (N_6752,N_4007,N_4309);
or U6753 (N_6753,N_4638,N_5504);
nand U6754 (N_6754,N_4662,N_4578);
nand U6755 (N_6755,N_5615,N_4417);
and U6756 (N_6756,N_5913,N_4168);
nand U6757 (N_6757,N_4670,N_4210);
or U6758 (N_6758,N_4155,N_5097);
nor U6759 (N_6759,N_5563,N_5488);
or U6760 (N_6760,N_4182,N_5288);
nand U6761 (N_6761,N_4529,N_4444);
or U6762 (N_6762,N_5091,N_5770);
and U6763 (N_6763,N_5580,N_5359);
nor U6764 (N_6764,N_5264,N_4495);
nor U6765 (N_6765,N_5551,N_5291);
nor U6766 (N_6766,N_4956,N_5001);
nor U6767 (N_6767,N_4363,N_5610);
and U6768 (N_6768,N_4512,N_4116);
and U6769 (N_6769,N_5128,N_4446);
nand U6770 (N_6770,N_5025,N_4316);
and U6771 (N_6771,N_5575,N_4863);
nor U6772 (N_6772,N_5385,N_4484);
or U6773 (N_6773,N_5934,N_5715);
nor U6774 (N_6774,N_5939,N_5912);
and U6775 (N_6775,N_4013,N_5130);
and U6776 (N_6776,N_5231,N_4738);
or U6777 (N_6777,N_4900,N_5014);
or U6778 (N_6778,N_5739,N_4307);
nand U6779 (N_6779,N_4831,N_5421);
nand U6780 (N_6780,N_4208,N_4861);
xnor U6781 (N_6781,N_5876,N_5621);
nand U6782 (N_6782,N_5109,N_5379);
and U6783 (N_6783,N_4628,N_4947);
xnor U6784 (N_6784,N_5188,N_4858);
or U6785 (N_6785,N_5643,N_4479);
and U6786 (N_6786,N_5154,N_4251);
and U6787 (N_6787,N_4577,N_4030);
or U6788 (N_6788,N_5252,N_5570);
or U6789 (N_6789,N_4983,N_4135);
nand U6790 (N_6790,N_4978,N_5321);
nor U6791 (N_6791,N_4002,N_5491);
nor U6792 (N_6792,N_4069,N_5489);
and U6793 (N_6793,N_4926,N_5629);
or U6794 (N_6794,N_4220,N_4257);
xnor U6795 (N_6795,N_5828,N_4696);
nand U6796 (N_6796,N_4318,N_5241);
and U6797 (N_6797,N_4957,N_5778);
or U6798 (N_6798,N_5059,N_4830);
xnor U6799 (N_6799,N_4751,N_5958);
nand U6800 (N_6800,N_5328,N_4487);
and U6801 (N_6801,N_5686,N_5937);
and U6802 (N_6802,N_5124,N_5220);
and U6803 (N_6803,N_4706,N_5274);
xor U6804 (N_6804,N_4586,N_4412);
and U6805 (N_6805,N_5787,N_4431);
xor U6806 (N_6806,N_4195,N_5910);
nand U6807 (N_6807,N_5595,N_5721);
or U6808 (N_6808,N_4754,N_4306);
nand U6809 (N_6809,N_4707,N_4454);
and U6810 (N_6810,N_4523,N_4554);
and U6811 (N_6811,N_5349,N_5063);
or U6812 (N_6812,N_4601,N_5503);
and U6813 (N_6813,N_4736,N_4106);
and U6814 (N_6814,N_4362,N_5370);
and U6815 (N_6815,N_4869,N_4747);
or U6816 (N_6816,N_5900,N_5471);
xnor U6817 (N_6817,N_4692,N_5722);
xor U6818 (N_6818,N_5769,N_4376);
or U6819 (N_6819,N_5020,N_5914);
and U6820 (N_6820,N_4820,N_4768);
and U6821 (N_6821,N_5225,N_4287);
xnor U6822 (N_6822,N_5060,N_4987);
nand U6823 (N_6823,N_4334,N_5335);
or U6824 (N_6824,N_5760,N_4592);
nand U6825 (N_6825,N_5240,N_5448);
or U6826 (N_6826,N_5198,N_4183);
nand U6827 (N_6827,N_4533,N_5908);
and U6828 (N_6828,N_4524,N_4107);
or U6829 (N_6829,N_5208,N_4636);
nor U6830 (N_6830,N_5409,N_5295);
nor U6831 (N_6831,N_4163,N_5965);
nor U6832 (N_6832,N_4060,N_5017);
or U6833 (N_6833,N_5831,N_5226);
nand U6834 (N_6834,N_5134,N_5925);
xor U6835 (N_6835,N_5156,N_4468);
xnor U6836 (N_6836,N_4595,N_5628);
and U6837 (N_6837,N_5262,N_4527);
and U6838 (N_6838,N_4386,N_5056);
and U6839 (N_6839,N_4907,N_5844);
nand U6840 (N_6840,N_5931,N_5915);
or U6841 (N_6841,N_5874,N_4633);
or U6842 (N_6842,N_4733,N_5545);
or U6843 (N_6843,N_5589,N_5569);
and U6844 (N_6844,N_5079,N_5882);
and U6845 (N_6845,N_4873,N_4953);
or U6846 (N_6846,N_4972,N_5378);
nor U6847 (N_6847,N_4834,N_5456);
nor U6848 (N_6848,N_5405,N_4380);
nand U6849 (N_6849,N_5694,N_4218);
xor U6850 (N_6850,N_5986,N_5455);
and U6851 (N_6851,N_5435,N_5116);
xor U6852 (N_6852,N_4466,N_4851);
or U6853 (N_6853,N_5279,N_4823);
and U6854 (N_6854,N_5268,N_4131);
nor U6855 (N_6855,N_5058,N_5256);
and U6856 (N_6856,N_4917,N_5608);
or U6857 (N_6857,N_5957,N_5253);
nand U6858 (N_6858,N_4879,N_4789);
or U6859 (N_6859,N_4944,N_5082);
nand U6860 (N_6860,N_5026,N_5129);
nor U6861 (N_6861,N_5107,N_5319);
and U6862 (N_6862,N_4779,N_5630);
nand U6863 (N_6863,N_4588,N_5823);
or U6864 (N_6864,N_5075,N_5626);
or U6865 (N_6865,N_5467,N_4568);
nand U6866 (N_6866,N_5472,N_4011);
or U6867 (N_6867,N_4129,N_5242);
or U6868 (N_6868,N_4145,N_4014);
nor U6869 (N_6869,N_4201,N_5192);
or U6870 (N_6870,N_4969,N_5781);
nor U6871 (N_6871,N_5318,N_5440);
nor U6872 (N_6872,N_5622,N_4770);
and U6873 (N_6873,N_5717,N_5928);
and U6874 (N_6874,N_4839,N_5135);
or U6875 (N_6875,N_4098,N_5691);
nor U6876 (N_6876,N_4916,N_5454);
and U6877 (N_6877,N_5446,N_4382);
or U6878 (N_6878,N_5111,N_5203);
and U6879 (N_6879,N_5120,N_4379);
nand U6880 (N_6880,N_4031,N_5834);
nand U6881 (N_6881,N_4553,N_4973);
nand U6882 (N_6882,N_5247,N_4705);
or U6883 (N_6883,N_4100,N_5649);
nor U6884 (N_6884,N_4614,N_5827);
and U6885 (N_6885,N_5287,N_5564);
nor U6886 (N_6886,N_4940,N_5853);
nand U6887 (N_6887,N_4404,N_5822);
nand U6888 (N_6888,N_4805,N_5585);
or U6889 (N_6889,N_5019,N_4794);
xnor U6890 (N_6890,N_5275,N_5298);
nor U6891 (N_6891,N_4330,N_5896);
or U6892 (N_6892,N_5419,N_5368);
nor U6893 (N_6893,N_5494,N_5403);
nand U6894 (N_6894,N_5750,N_4769);
nand U6895 (N_6895,N_4439,N_4855);
xor U6896 (N_6896,N_5008,N_5948);
nand U6897 (N_6897,N_4280,N_5523);
nand U6898 (N_6898,N_4253,N_5789);
nor U6899 (N_6899,N_4204,N_5519);
and U6900 (N_6900,N_4594,N_4813);
or U6901 (N_6901,N_5539,N_4317);
or U6902 (N_6902,N_5224,N_4651);
nand U6903 (N_6903,N_5369,N_4867);
or U6904 (N_6904,N_4630,N_5826);
nor U6905 (N_6905,N_5878,N_5552);
nor U6906 (N_6906,N_4924,N_5367);
xor U6907 (N_6907,N_5666,N_4925);
nand U6908 (N_6908,N_4159,N_5420);
nand U6909 (N_6909,N_4865,N_5375);
or U6910 (N_6910,N_5045,N_4909);
and U6911 (N_6911,N_5676,N_4903);
xor U6912 (N_6912,N_5761,N_5755);
or U6913 (N_6913,N_4293,N_4637);
or U6914 (N_6914,N_4702,N_4585);
and U6915 (N_6915,N_5476,N_5817);
and U6916 (N_6916,N_5858,N_5393);
and U6917 (N_6917,N_5329,N_4332);
nand U6918 (N_6918,N_5496,N_5230);
and U6919 (N_6919,N_5333,N_5289);
or U6920 (N_6920,N_5132,N_4569);
nor U6921 (N_6921,N_5364,N_4535);
xnor U6922 (N_6922,N_4305,N_5702);
nand U6923 (N_6923,N_5661,N_4167);
or U6924 (N_6924,N_4558,N_4153);
and U6925 (N_6925,N_4152,N_4360);
nor U6926 (N_6926,N_5845,N_5560);
or U6927 (N_6927,N_5176,N_5917);
nand U6928 (N_6928,N_5438,N_4520);
or U6929 (N_6929,N_5046,N_4927);
nor U6930 (N_6930,N_4420,N_5146);
nor U6931 (N_6931,N_5631,N_5081);
or U6932 (N_6932,N_4505,N_4063);
and U6933 (N_6933,N_5139,N_5429);
and U6934 (N_6934,N_4602,N_4343);
nor U6935 (N_6935,N_5890,N_5905);
xnor U6936 (N_6936,N_4913,N_4755);
nor U6937 (N_6937,N_4616,N_5029);
or U6938 (N_6938,N_5668,N_4285);
nor U6939 (N_6939,N_4899,N_5576);
and U6940 (N_6940,N_5235,N_4784);
or U6941 (N_6941,N_4147,N_4093);
nor U6942 (N_6942,N_4164,N_5305);
nor U6943 (N_6943,N_4710,N_5833);
or U6944 (N_6944,N_4108,N_4346);
and U6945 (N_6945,N_4840,N_4566);
and U6946 (N_6946,N_4502,N_4440);
xnor U6947 (N_6947,N_4165,N_4884);
nor U6948 (N_6948,N_4205,N_4453);
nor U6949 (N_6949,N_5976,N_5040);
nand U6950 (N_6950,N_5667,N_4158);
and U6951 (N_6951,N_5848,N_5842);
nand U6952 (N_6952,N_4124,N_4686);
and U6953 (N_6953,N_4435,N_4213);
or U6954 (N_6954,N_5602,N_5782);
nand U6955 (N_6955,N_4319,N_4634);
nor U6956 (N_6956,N_4775,N_5015);
and U6957 (N_6957,N_5320,N_5115);
and U6958 (N_6958,N_4801,N_4756);
or U6959 (N_6959,N_5566,N_4500);
and U6960 (N_6960,N_4799,N_5043);
nor U6961 (N_6961,N_4847,N_4525);
and U6962 (N_6962,N_5533,N_5618);
or U6963 (N_6963,N_4474,N_4150);
nor U6964 (N_6964,N_4200,N_5864);
and U6965 (N_6965,N_4298,N_4934);
nor U6966 (N_6966,N_5165,N_4255);
nor U6967 (N_6967,N_5894,N_4432);
nand U6968 (N_6968,N_5495,N_5037);
nor U6969 (N_6969,N_4912,N_4369);
nand U6970 (N_6970,N_4579,N_5187);
nor U6971 (N_6971,N_4954,N_5884);
and U6972 (N_6972,N_4522,N_5260);
xor U6973 (N_6973,N_4231,N_5142);
nor U6974 (N_6974,N_5768,N_5388);
or U6975 (N_6975,N_5961,N_5880);
nand U6976 (N_6976,N_5286,N_4800);
nand U6977 (N_6977,N_5179,N_5646);
or U6978 (N_6978,N_5525,N_5790);
nor U6979 (N_6979,N_5084,N_5572);
nand U6980 (N_6980,N_4078,N_4993);
and U6981 (N_6981,N_5929,N_5725);
nor U6982 (N_6982,N_5339,N_5028);
nor U6983 (N_6983,N_4181,N_4077);
or U6984 (N_6984,N_5981,N_4422);
nor U6985 (N_6985,N_4999,N_4528);
nor U6986 (N_6986,N_5767,N_4377);
xor U6987 (N_6987,N_5269,N_4036);
nand U6988 (N_6988,N_5591,N_5886);
or U6989 (N_6989,N_5951,N_4125);
nand U6990 (N_6990,N_4548,N_5689);
xor U6991 (N_6991,N_5093,N_5839);
or U6992 (N_6992,N_5940,N_4214);
nand U6993 (N_6993,N_4489,N_4166);
nor U6994 (N_6994,N_4752,N_4815);
nor U6995 (N_6995,N_4650,N_5515);
and U6996 (N_6996,N_5432,N_4652);
nor U6997 (N_6997,N_5383,N_5633);
xor U6998 (N_6998,N_4065,N_4199);
or U6999 (N_6999,N_4880,N_5803);
nor U7000 (N_7000,N_5378,N_5629);
nand U7001 (N_7001,N_5341,N_5502);
and U7002 (N_7002,N_5476,N_4126);
or U7003 (N_7003,N_5554,N_5534);
nor U7004 (N_7004,N_4179,N_4774);
and U7005 (N_7005,N_5702,N_5834);
or U7006 (N_7006,N_5798,N_4626);
and U7007 (N_7007,N_5894,N_5564);
nand U7008 (N_7008,N_5239,N_4158);
nor U7009 (N_7009,N_4666,N_5723);
or U7010 (N_7010,N_5248,N_5912);
nor U7011 (N_7011,N_4066,N_5262);
and U7012 (N_7012,N_5796,N_4861);
nand U7013 (N_7013,N_4204,N_4547);
nor U7014 (N_7014,N_4855,N_5670);
or U7015 (N_7015,N_5528,N_5879);
nor U7016 (N_7016,N_5356,N_4394);
xor U7017 (N_7017,N_5928,N_4686);
nand U7018 (N_7018,N_4367,N_4317);
and U7019 (N_7019,N_5713,N_4462);
xnor U7020 (N_7020,N_4176,N_5037);
nand U7021 (N_7021,N_4421,N_5548);
or U7022 (N_7022,N_5426,N_4608);
xor U7023 (N_7023,N_5411,N_4475);
nand U7024 (N_7024,N_4730,N_4991);
nand U7025 (N_7025,N_5955,N_5414);
and U7026 (N_7026,N_4724,N_5251);
nand U7027 (N_7027,N_5061,N_4342);
and U7028 (N_7028,N_4075,N_4704);
nand U7029 (N_7029,N_4157,N_4855);
or U7030 (N_7030,N_5723,N_4965);
and U7031 (N_7031,N_4046,N_5024);
or U7032 (N_7032,N_5264,N_5021);
nand U7033 (N_7033,N_4015,N_4824);
or U7034 (N_7034,N_4367,N_4416);
xnor U7035 (N_7035,N_4594,N_4738);
nor U7036 (N_7036,N_5162,N_4792);
nand U7037 (N_7037,N_5792,N_5359);
and U7038 (N_7038,N_4128,N_5098);
nand U7039 (N_7039,N_4121,N_5783);
nor U7040 (N_7040,N_5787,N_4785);
nor U7041 (N_7041,N_4306,N_4378);
xnor U7042 (N_7042,N_4320,N_4525);
nor U7043 (N_7043,N_5679,N_4402);
nor U7044 (N_7044,N_4150,N_5358);
nor U7045 (N_7045,N_5369,N_5982);
and U7046 (N_7046,N_4926,N_4339);
xnor U7047 (N_7047,N_5709,N_5133);
and U7048 (N_7048,N_4366,N_4916);
and U7049 (N_7049,N_5607,N_5820);
and U7050 (N_7050,N_4614,N_4048);
xnor U7051 (N_7051,N_5261,N_5240);
nor U7052 (N_7052,N_5739,N_4666);
nor U7053 (N_7053,N_5564,N_5616);
nand U7054 (N_7054,N_5460,N_4747);
nand U7055 (N_7055,N_4373,N_4305);
or U7056 (N_7056,N_4654,N_4534);
or U7057 (N_7057,N_4244,N_4084);
or U7058 (N_7058,N_4226,N_5787);
and U7059 (N_7059,N_5062,N_5580);
or U7060 (N_7060,N_5744,N_4915);
nand U7061 (N_7061,N_5693,N_5334);
or U7062 (N_7062,N_5510,N_5234);
nor U7063 (N_7063,N_4255,N_5018);
nor U7064 (N_7064,N_4039,N_4116);
nand U7065 (N_7065,N_5532,N_5245);
xnor U7066 (N_7066,N_4628,N_5269);
and U7067 (N_7067,N_5467,N_4271);
nand U7068 (N_7068,N_5196,N_4583);
nor U7069 (N_7069,N_5253,N_4064);
nor U7070 (N_7070,N_5221,N_5861);
and U7071 (N_7071,N_4194,N_5857);
or U7072 (N_7072,N_5904,N_4550);
or U7073 (N_7073,N_5988,N_5994);
nor U7074 (N_7074,N_5924,N_5288);
nor U7075 (N_7075,N_5754,N_4262);
nor U7076 (N_7076,N_5158,N_5194);
or U7077 (N_7077,N_5169,N_4709);
nand U7078 (N_7078,N_4717,N_5185);
nand U7079 (N_7079,N_5339,N_4862);
nor U7080 (N_7080,N_4337,N_4695);
and U7081 (N_7081,N_5207,N_4101);
and U7082 (N_7082,N_4299,N_5551);
nand U7083 (N_7083,N_5780,N_4476);
and U7084 (N_7084,N_4085,N_4454);
nand U7085 (N_7085,N_4419,N_5001);
nand U7086 (N_7086,N_4844,N_5568);
or U7087 (N_7087,N_5897,N_5021);
or U7088 (N_7088,N_4504,N_4824);
nor U7089 (N_7089,N_4269,N_4981);
xnor U7090 (N_7090,N_4539,N_4203);
and U7091 (N_7091,N_4193,N_4811);
nand U7092 (N_7092,N_5307,N_5418);
and U7093 (N_7093,N_5289,N_5497);
and U7094 (N_7094,N_4982,N_5549);
or U7095 (N_7095,N_5355,N_4256);
and U7096 (N_7096,N_5032,N_4381);
or U7097 (N_7097,N_4486,N_5660);
and U7098 (N_7098,N_5933,N_5844);
and U7099 (N_7099,N_4977,N_4726);
or U7100 (N_7100,N_4563,N_4223);
nor U7101 (N_7101,N_4703,N_4458);
xor U7102 (N_7102,N_4168,N_4846);
and U7103 (N_7103,N_4720,N_4835);
or U7104 (N_7104,N_5598,N_5196);
nand U7105 (N_7105,N_5984,N_5236);
or U7106 (N_7106,N_4281,N_4539);
or U7107 (N_7107,N_5895,N_4800);
or U7108 (N_7108,N_5564,N_4969);
or U7109 (N_7109,N_5556,N_5809);
nand U7110 (N_7110,N_4951,N_5046);
or U7111 (N_7111,N_4574,N_5489);
and U7112 (N_7112,N_5554,N_4613);
nand U7113 (N_7113,N_5018,N_5394);
nand U7114 (N_7114,N_4974,N_5198);
or U7115 (N_7115,N_5595,N_4149);
nor U7116 (N_7116,N_5119,N_4254);
and U7117 (N_7117,N_5864,N_4327);
or U7118 (N_7118,N_5203,N_4787);
xor U7119 (N_7119,N_5844,N_4575);
or U7120 (N_7120,N_4290,N_5605);
nand U7121 (N_7121,N_5828,N_5945);
xor U7122 (N_7122,N_5124,N_4424);
nand U7123 (N_7123,N_5888,N_5870);
and U7124 (N_7124,N_4111,N_5002);
nor U7125 (N_7125,N_4661,N_5664);
and U7126 (N_7126,N_4524,N_5287);
and U7127 (N_7127,N_4671,N_5844);
xor U7128 (N_7128,N_5487,N_5872);
and U7129 (N_7129,N_4947,N_5616);
nor U7130 (N_7130,N_4304,N_4101);
nand U7131 (N_7131,N_5259,N_5874);
or U7132 (N_7132,N_5952,N_5187);
or U7133 (N_7133,N_4015,N_4919);
nand U7134 (N_7134,N_4948,N_4939);
or U7135 (N_7135,N_5056,N_4381);
nor U7136 (N_7136,N_4957,N_4756);
xor U7137 (N_7137,N_4340,N_5979);
nand U7138 (N_7138,N_5518,N_5119);
or U7139 (N_7139,N_4310,N_4541);
nand U7140 (N_7140,N_5265,N_5395);
or U7141 (N_7141,N_5681,N_4145);
nand U7142 (N_7142,N_5131,N_4052);
xnor U7143 (N_7143,N_5773,N_4015);
nor U7144 (N_7144,N_5377,N_5880);
and U7145 (N_7145,N_4447,N_5985);
nand U7146 (N_7146,N_4638,N_5606);
nor U7147 (N_7147,N_4625,N_4864);
or U7148 (N_7148,N_5952,N_5179);
nand U7149 (N_7149,N_5819,N_5321);
nand U7150 (N_7150,N_4775,N_4687);
or U7151 (N_7151,N_5075,N_4940);
or U7152 (N_7152,N_5224,N_5333);
or U7153 (N_7153,N_5143,N_5028);
or U7154 (N_7154,N_4409,N_5533);
and U7155 (N_7155,N_4173,N_4285);
xor U7156 (N_7156,N_5147,N_5607);
or U7157 (N_7157,N_4547,N_4950);
and U7158 (N_7158,N_4201,N_4140);
or U7159 (N_7159,N_5295,N_4160);
and U7160 (N_7160,N_5547,N_4326);
nor U7161 (N_7161,N_5871,N_5433);
nand U7162 (N_7162,N_4957,N_5735);
or U7163 (N_7163,N_4530,N_5079);
xnor U7164 (N_7164,N_5964,N_4398);
and U7165 (N_7165,N_4999,N_4307);
nand U7166 (N_7166,N_4178,N_5640);
nor U7167 (N_7167,N_4548,N_5543);
nand U7168 (N_7168,N_5756,N_5584);
nor U7169 (N_7169,N_5718,N_4674);
or U7170 (N_7170,N_4554,N_5204);
nand U7171 (N_7171,N_4845,N_5486);
or U7172 (N_7172,N_4021,N_5955);
nand U7173 (N_7173,N_5239,N_4232);
or U7174 (N_7174,N_4171,N_4674);
nor U7175 (N_7175,N_4254,N_5199);
or U7176 (N_7176,N_4435,N_5849);
and U7177 (N_7177,N_5228,N_4148);
or U7178 (N_7178,N_5124,N_4383);
or U7179 (N_7179,N_5781,N_4813);
or U7180 (N_7180,N_4916,N_4417);
xor U7181 (N_7181,N_4879,N_4548);
or U7182 (N_7182,N_4973,N_4586);
and U7183 (N_7183,N_5176,N_5798);
nor U7184 (N_7184,N_4764,N_5557);
nor U7185 (N_7185,N_5569,N_5830);
nand U7186 (N_7186,N_5051,N_5387);
nand U7187 (N_7187,N_4352,N_5874);
or U7188 (N_7188,N_5755,N_5874);
nor U7189 (N_7189,N_5078,N_4225);
xnor U7190 (N_7190,N_5793,N_4811);
nand U7191 (N_7191,N_5427,N_4445);
nor U7192 (N_7192,N_4171,N_4641);
and U7193 (N_7193,N_4381,N_4188);
nor U7194 (N_7194,N_5671,N_5053);
or U7195 (N_7195,N_5611,N_5026);
and U7196 (N_7196,N_4661,N_5690);
and U7197 (N_7197,N_5373,N_4711);
xnor U7198 (N_7198,N_5769,N_5541);
or U7199 (N_7199,N_5011,N_5116);
nor U7200 (N_7200,N_4958,N_5795);
and U7201 (N_7201,N_5743,N_4414);
nand U7202 (N_7202,N_4689,N_4417);
nor U7203 (N_7203,N_4519,N_5143);
and U7204 (N_7204,N_5483,N_4019);
or U7205 (N_7205,N_5753,N_4297);
or U7206 (N_7206,N_4826,N_5589);
and U7207 (N_7207,N_4933,N_5418);
or U7208 (N_7208,N_4071,N_5196);
or U7209 (N_7209,N_4390,N_4272);
nand U7210 (N_7210,N_5070,N_4664);
or U7211 (N_7211,N_5891,N_4896);
xnor U7212 (N_7212,N_5129,N_4933);
nor U7213 (N_7213,N_5683,N_4560);
or U7214 (N_7214,N_4569,N_4177);
nand U7215 (N_7215,N_5094,N_5143);
nand U7216 (N_7216,N_5162,N_4965);
and U7217 (N_7217,N_5318,N_4382);
nand U7218 (N_7218,N_5507,N_4129);
nand U7219 (N_7219,N_4626,N_4309);
or U7220 (N_7220,N_4553,N_5436);
and U7221 (N_7221,N_4966,N_5118);
and U7222 (N_7222,N_4001,N_5316);
and U7223 (N_7223,N_5569,N_4960);
xnor U7224 (N_7224,N_4474,N_4930);
and U7225 (N_7225,N_4677,N_4745);
nand U7226 (N_7226,N_4145,N_5054);
nor U7227 (N_7227,N_4631,N_5102);
nand U7228 (N_7228,N_4773,N_4219);
and U7229 (N_7229,N_5106,N_4533);
xnor U7230 (N_7230,N_4101,N_4739);
nor U7231 (N_7231,N_5940,N_5549);
nand U7232 (N_7232,N_4456,N_4067);
or U7233 (N_7233,N_5565,N_5671);
nand U7234 (N_7234,N_4165,N_4309);
and U7235 (N_7235,N_5235,N_4957);
or U7236 (N_7236,N_4794,N_5066);
or U7237 (N_7237,N_5417,N_4402);
nor U7238 (N_7238,N_5498,N_5221);
or U7239 (N_7239,N_4072,N_5679);
nor U7240 (N_7240,N_4727,N_4536);
nor U7241 (N_7241,N_4118,N_4405);
nor U7242 (N_7242,N_5314,N_5682);
nor U7243 (N_7243,N_4026,N_4999);
and U7244 (N_7244,N_5345,N_5071);
nand U7245 (N_7245,N_5488,N_5067);
nor U7246 (N_7246,N_4945,N_5438);
nand U7247 (N_7247,N_4903,N_5392);
nand U7248 (N_7248,N_4221,N_4654);
nand U7249 (N_7249,N_5513,N_4352);
xnor U7250 (N_7250,N_4304,N_5289);
and U7251 (N_7251,N_5926,N_4075);
or U7252 (N_7252,N_5498,N_4146);
nor U7253 (N_7253,N_5048,N_5585);
nand U7254 (N_7254,N_4473,N_5373);
nor U7255 (N_7255,N_5272,N_4124);
and U7256 (N_7256,N_4773,N_5768);
xor U7257 (N_7257,N_4633,N_5953);
and U7258 (N_7258,N_5808,N_4311);
nand U7259 (N_7259,N_4268,N_5260);
or U7260 (N_7260,N_5466,N_5400);
nor U7261 (N_7261,N_5553,N_4678);
or U7262 (N_7262,N_4942,N_4452);
or U7263 (N_7263,N_4765,N_5547);
or U7264 (N_7264,N_4065,N_4623);
nor U7265 (N_7265,N_4947,N_4799);
xnor U7266 (N_7266,N_5806,N_4612);
xor U7267 (N_7267,N_4638,N_4635);
nand U7268 (N_7268,N_4277,N_5960);
or U7269 (N_7269,N_5201,N_4232);
and U7270 (N_7270,N_5742,N_5740);
nand U7271 (N_7271,N_5311,N_5044);
xor U7272 (N_7272,N_4840,N_5951);
or U7273 (N_7273,N_5522,N_5863);
and U7274 (N_7274,N_4963,N_5210);
nand U7275 (N_7275,N_4351,N_5183);
and U7276 (N_7276,N_5773,N_4251);
nor U7277 (N_7277,N_5410,N_4894);
nor U7278 (N_7278,N_4786,N_4368);
nand U7279 (N_7279,N_5136,N_4367);
nand U7280 (N_7280,N_4198,N_5292);
nor U7281 (N_7281,N_4597,N_5352);
nand U7282 (N_7282,N_5738,N_5265);
nor U7283 (N_7283,N_4795,N_4789);
nand U7284 (N_7284,N_4781,N_4965);
and U7285 (N_7285,N_4654,N_4665);
nand U7286 (N_7286,N_5400,N_5250);
xor U7287 (N_7287,N_5574,N_4812);
nand U7288 (N_7288,N_5285,N_4642);
nand U7289 (N_7289,N_5101,N_5737);
xor U7290 (N_7290,N_4217,N_5762);
xor U7291 (N_7291,N_5770,N_5170);
nand U7292 (N_7292,N_4238,N_4799);
xor U7293 (N_7293,N_5780,N_4857);
xnor U7294 (N_7294,N_5130,N_5571);
xnor U7295 (N_7295,N_4303,N_5294);
or U7296 (N_7296,N_4044,N_4961);
and U7297 (N_7297,N_5398,N_5394);
nor U7298 (N_7298,N_5251,N_5266);
nand U7299 (N_7299,N_4859,N_4345);
or U7300 (N_7300,N_4519,N_4777);
nor U7301 (N_7301,N_5918,N_4448);
and U7302 (N_7302,N_4371,N_4249);
and U7303 (N_7303,N_5375,N_4028);
nand U7304 (N_7304,N_5947,N_5221);
and U7305 (N_7305,N_5963,N_4359);
or U7306 (N_7306,N_4180,N_5879);
nor U7307 (N_7307,N_4227,N_4966);
or U7308 (N_7308,N_4149,N_4472);
xor U7309 (N_7309,N_5993,N_4364);
nor U7310 (N_7310,N_4171,N_5086);
nand U7311 (N_7311,N_5390,N_5511);
nor U7312 (N_7312,N_4432,N_4575);
nor U7313 (N_7313,N_4123,N_4327);
and U7314 (N_7314,N_4192,N_4938);
xor U7315 (N_7315,N_5090,N_5864);
nand U7316 (N_7316,N_5447,N_5810);
or U7317 (N_7317,N_4678,N_5963);
nand U7318 (N_7318,N_4633,N_4110);
and U7319 (N_7319,N_4824,N_4203);
and U7320 (N_7320,N_5928,N_5210);
and U7321 (N_7321,N_4553,N_4614);
and U7322 (N_7322,N_5393,N_4326);
or U7323 (N_7323,N_4332,N_5528);
xor U7324 (N_7324,N_4954,N_5630);
xnor U7325 (N_7325,N_5617,N_4778);
or U7326 (N_7326,N_4324,N_4287);
nand U7327 (N_7327,N_5910,N_5921);
and U7328 (N_7328,N_5690,N_5661);
nand U7329 (N_7329,N_4640,N_4109);
nor U7330 (N_7330,N_5757,N_5305);
nor U7331 (N_7331,N_5629,N_5693);
xnor U7332 (N_7332,N_4397,N_4050);
nand U7333 (N_7333,N_5773,N_4958);
nand U7334 (N_7334,N_5455,N_4361);
nand U7335 (N_7335,N_5605,N_5540);
nor U7336 (N_7336,N_5082,N_4778);
nor U7337 (N_7337,N_5026,N_4359);
or U7338 (N_7338,N_4693,N_4001);
xnor U7339 (N_7339,N_5743,N_5890);
and U7340 (N_7340,N_4052,N_5670);
nand U7341 (N_7341,N_5335,N_5143);
nor U7342 (N_7342,N_5157,N_5210);
nor U7343 (N_7343,N_4662,N_4279);
nand U7344 (N_7344,N_5184,N_5828);
and U7345 (N_7345,N_4470,N_4556);
and U7346 (N_7346,N_5330,N_4198);
nand U7347 (N_7347,N_5229,N_4616);
xnor U7348 (N_7348,N_4241,N_4994);
nor U7349 (N_7349,N_4158,N_4257);
and U7350 (N_7350,N_5128,N_5783);
xnor U7351 (N_7351,N_4950,N_5336);
nand U7352 (N_7352,N_5959,N_4535);
and U7353 (N_7353,N_5658,N_5053);
nand U7354 (N_7354,N_4175,N_4872);
nor U7355 (N_7355,N_5159,N_5298);
and U7356 (N_7356,N_5745,N_5172);
and U7357 (N_7357,N_4408,N_4340);
and U7358 (N_7358,N_5207,N_4052);
xor U7359 (N_7359,N_5374,N_4874);
and U7360 (N_7360,N_4511,N_5837);
nor U7361 (N_7361,N_4210,N_5611);
nand U7362 (N_7362,N_5246,N_4294);
nor U7363 (N_7363,N_5476,N_4487);
xnor U7364 (N_7364,N_5860,N_4422);
or U7365 (N_7365,N_4250,N_5685);
or U7366 (N_7366,N_4178,N_4828);
nand U7367 (N_7367,N_5526,N_4714);
or U7368 (N_7368,N_5065,N_5048);
nor U7369 (N_7369,N_5313,N_4776);
or U7370 (N_7370,N_4559,N_4896);
nor U7371 (N_7371,N_5804,N_5786);
or U7372 (N_7372,N_4613,N_4615);
nand U7373 (N_7373,N_4367,N_5458);
or U7374 (N_7374,N_4308,N_5494);
xnor U7375 (N_7375,N_5238,N_4699);
or U7376 (N_7376,N_5033,N_5716);
and U7377 (N_7377,N_5085,N_5966);
nor U7378 (N_7378,N_4565,N_5525);
or U7379 (N_7379,N_5633,N_4116);
and U7380 (N_7380,N_5535,N_5896);
nand U7381 (N_7381,N_4709,N_4785);
or U7382 (N_7382,N_4757,N_5560);
xnor U7383 (N_7383,N_4337,N_5783);
nor U7384 (N_7384,N_5267,N_4688);
and U7385 (N_7385,N_5105,N_4637);
nor U7386 (N_7386,N_4807,N_4796);
or U7387 (N_7387,N_5444,N_4954);
or U7388 (N_7388,N_5297,N_4467);
nor U7389 (N_7389,N_4403,N_5404);
xnor U7390 (N_7390,N_4104,N_5348);
or U7391 (N_7391,N_5270,N_5133);
nor U7392 (N_7392,N_4098,N_5434);
xnor U7393 (N_7393,N_4565,N_4874);
or U7394 (N_7394,N_4758,N_4584);
or U7395 (N_7395,N_5872,N_5136);
xor U7396 (N_7396,N_5752,N_4263);
nor U7397 (N_7397,N_4225,N_4301);
and U7398 (N_7398,N_5225,N_4361);
and U7399 (N_7399,N_5986,N_5677);
nand U7400 (N_7400,N_4569,N_5815);
nor U7401 (N_7401,N_4779,N_4839);
or U7402 (N_7402,N_5502,N_4604);
nor U7403 (N_7403,N_5830,N_4061);
and U7404 (N_7404,N_4874,N_4944);
nor U7405 (N_7405,N_5754,N_5820);
and U7406 (N_7406,N_4507,N_4173);
xnor U7407 (N_7407,N_4280,N_5515);
nand U7408 (N_7408,N_4108,N_5449);
and U7409 (N_7409,N_4518,N_4072);
xnor U7410 (N_7410,N_4190,N_4950);
and U7411 (N_7411,N_4561,N_4048);
and U7412 (N_7412,N_4820,N_5013);
or U7413 (N_7413,N_5520,N_5737);
or U7414 (N_7414,N_4898,N_4565);
nor U7415 (N_7415,N_4753,N_4847);
or U7416 (N_7416,N_5561,N_5222);
nor U7417 (N_7417,N_4774,N_4280);
nor U7418 (N_7418,N_5240,N_4475);
and U7419 (N_7419,N_5840,N_5576);
and U7420 (N_7420,N_5173,N_4581);
or U7421 (N_7421,N_4331,N_5088);
nand U7422 (N_7422,N_4735,N_5985);
and U7423 (N_7423,N_4283,N_5744);
nor U7424 (N_7424,N_4226,N_5775);
xor U7425 (N_7425,N_4562,N_5671);
nor U7426 (N_7426,N_4243,N_4589);
nor U7427 (N_7427,N_5926,N_5502);
nor U7428 (N_7428,N_5461,N_5554);
and U7429 (N_7429,N_4420,N_5558);
and U7430 (N_7430,N_5952,N_4117);
or U7431 (N_7431,N_5580,N_5123);
and U7432 (N_7432,N_4967,N_5112);
or U7433 (N_7433,N_5238,N_4227);
and U7434 (N_7434,N_4230,N_5089);
nand U7435 (N_7435,N_4177,N_4291);
xnor U7436 (N_7436,N_4714,N_5183);
and U7437 (N_7437,N_5846,N_4673);
nand U7438 (N_7438,N_4566,N_4904);
nand U7439 (N_7439,N_4319,N_5511);
or U7440 (N_7440,N_4144,N_5172);
nand U7441 (N_7441,N_4386,N_4718);
nor U7442 (N_7442,N_5319,N_4064);
nor U7443 (N_7443,N_4484,N_4138);
nand U7444 (N_7444,N_4516,N_5198);
nand U7445 (N_7445,N_5754,N_4142);
xnor U7446 (N_7446,N_4262,N_5409);
nand U7447 (N_7447,N_5385,N_4765);
xnor U7448 (N_7448,N_5279,N_5100);
nor U7449 (N_7449,N_5236,N_4093);
xnor U7450 (N_7450,N_5218,N_4948);
nand U7451 (N_7451,N_5066,N_4680);
xnor U7452 (N_7452,N_5622,N_5615);
nor U7453 (N_7453,N_4382,N_4000);
nand U7454 (N_7454,N_5347,N_4277);
and U7455 (N_7455,N_4166,N_5870);
nor U7456 (N_7456,N_5378,N_4497);
nand U7457 (N_7457,N_4625,N_4807);
or U7458 (N_7458,N_5873,N_4145);
and U7459 (N_7459,N_5525,N_5773);
and U7460 (N_7460,N_5942,N_5063);
nor U7461 (N_7461,N_5134,N_4689);
xnor U7462 (N_7462,N_5265,N_4740);
nand U7463 (N_7463,N_4026,N_4784);
nand U7464 (N_7464,N_4665,N_5981);
nand U7465 (N_7465,N_4228,N_5411);
or U7466 (N_7466,N_4059,N_4550);
or U7467 (N_7467,N_4319,N_4770);
and U7468 (N_7468,N_4113,N_5826);
or U7469 (N_7469,N_4474,N_4465);
nor U7470 (N_7470,N_4973,N_4889);
and U7471 (N_7471,N_4366,N_5752);
and U7472 (N_7472,N_4135,N_4989);
or U7473 (N_7473,N_4612,N_5344);
or U7474 (N_7474,N_5005,N_5892);
or U7475 (N_7475,N_5845,N_5909);
nand U7476 (N_7476,N_5721,N_5127);
nor U7477 (N_7477,N_4269,N_4916);
nor U7478 (N_7478,N_4882,N_4877);
xnor U7479 (N_7479,N_4671,N_5200);
and U7480 (N_7480,N_4707,N_5614);
nand U7481 (N_7481,N_5995,N_5963);
or U7482 (N_7482,N_4089,N_4628);
and U7483 (N_7483,N_4886,N_5768);
or U7484 (N_7484,N_4941,N_5176);
nand U7485 (N_7485,N_4813,N_5709);
xnor U7486 (N_7486,N_5308,N_5033);
or U7487 (N_7487,N_5747,N_5108);
and U7488 (N_7488,N_4296,N_4698);
and U7489 (N_7489,N_4850,N_4396);
nor U7490 (N_7490,N_5519,N_5297);
and U7491 (N_7491,N_4670,N_4957);
nand U7492 (N_7492,N_4399,N_4903);
and U7493 (N_7493,N_5261,N_4745);
or U7494 (N_7494,N_5169,N_4004);
nor U7495 (N_7495,N_5755,N_5446);
xor U7496 (N_7496,N_4795,N_4065);
xor U7497 (N_7497,N_4125,N_4989);
nand U7498 (N_7498,N_4948,N_4728);
nand U7499 (N_7499,N_4348,N_5206);
nor U7500 (N_7500,N_5551,N_4100);
nand U7501 (N_7501,N_4361,N_5941);
and U7502 (N_7502,N_5746,N_5740);
and U7503 (N_7503,N_5571,N_4650);
nand U7504 (N_7504,N_4289,N_5811);
xnor U7505 (N_7505,N_5525,N_4056);
nand U7506 (N_7506,N_4315,N_4146);
and U7507 (N_7507,N_5925,N_5613);
or U7508 (N_7508,N_4665,N_4870);
or U7509 (N_7509,N_5152,N_5390);
nand U7510 (N_7510,N_5832,N_4244);
nor U7511 (N_7511,N_5613,N_4064);
nand U7512 (N_7512,N_4824,N_4471);
nor U7513 (N_7513,N_4643,N_4390);
and U7514 (N_7514,N_4187,N_4851);
or U7515 (N_7515,N_5045,N_4613);
nor U7516 (N_7516,N_4277,N_5280);
and U7517 (N_7517,N_5177,N_4385);
nor U7518 (N_7518,N_5077,N_4039);
and U7519 (N_7519,N_5798,N_5393);
or U7520 (N_7520,N_4190,N_5302);
or U7521 (N_7521,N_4217,N_5345);
or U7522 (N_7522,N_4803,N_5528);
and U7523 (N_7523,N_5730,N_4880);
or U7524 (N_7524,N_5650,N_5065);
nand U7525 (N_7525,N_4653,N_4391);
nor U7526 (N_7526,N_5319,N_4129);
nand U7527 (N_7527,N_4453,N_5464);
nand U7528 (N_7528,N_5585,N_5655);
and U7529 (N_7529,N_5326,N_5109);
nand U7530 (N_7530,N_4960,N_4532);
nor U7531 (N_7531,N_5109,N_4507);
or U7532 (N_7532,N_5375,N_5193);
nand U7533 (N_7533,N_5047,N_4909);
or U7534 (N_7534,N_4540,N_4018);
or U7535 (N_7535,N_5709,N_5770);
or U7536 (N_7536,N_4134,N_5209);
nor U7537 (N_7537,N_5204,N_4283);
xnor U7538 (N_7538,N_4162,N_4321);
and U7539 (N_7539,N_5386,N_5637);
nor U7540 (N_7540,N_5906,N_5253);
nor U7541 (N_7541,N_5735,N_5055);
or U7542 (N_7542,N_4320,N_4591);
and U7543 (N_7543,N_4155,N_4790);
nand U7544 (N_7544,N_5608,N_4562);
nor U7545 (N_7545,N_4198,N_4815);
or U7546 (N_7546,N_4104,N_4666);
and U7547 (N_7547,N_5300,N_4013);
and U7548 (N_7548,N_4395,N_4526);
nand U7549 (N_7549,N_5408,N_5492);
or U7550 (N_7550,N_5425,N_4619);
or U7551 (N_7551,N_5480,N_4231);
and U7552 (N_7552,N_5093,N_5099);
or U7553 (N_7553,N_5270,N_5439);
nand U7554 (N_7554,N_5706,N_5047);
nor U7555 (N_7555,N_5285,N_4748);
or U7556 (N_7556,N_4397,N_4577);
nand U7557 (N_7557,N_5826,N_4412);
and U7558 (N_7558,N_4265,N_4563);
nor U7559 (N_7559,N_5604,N_4810);
nor U7560 (N_7560,N_5957,N_4776);
xnor U7561 (N_7561,N_5874,N_5104);
nand U7562 (N_7562,N_4061,N_4652);
nor U7563 (N_7563,N_4440,N_4421);
or U7564 (N_7564,N_4194,N_4588);
and U7565 (N_7565,N_5550,N_5162);
or U7566 (N_7566,N_5635,N_4810);
nor U7567 (N_7567,N_4477,N_4811);
nand U7568 (N_7568,N_5948,N_4472);
xor U7569 (N_7569,N_4785,N_4604);
and U7570 (N_7570,N_4884,N_5493);
nand U7571 (N_7571,N_4359,N_5027);
nand U7572 (N_7572,N_5523,N_5054);
nor U7573 (N_7573,N_4924,N_5913);
nor U7574 (N_7574,N_4801,N_4959);
or U7575 (N_7575,N_5009,N_4889);
and U7576 (N_7576,N_5548,N_4159);
or U7577 (N_7577,N_5831,N_4284);
nand U7578 (N_7578,N_4689,N_5352);
and U7579 (N_7579,N_4691,N_5798);
and U7580 (N_7580,N_4405,N_5594);
or U7581 (N_7581,N_4623,N_4039);
nor U7582 (N_7582,N_4473,N_5112);
nand U7583 (N_7583,N_5061,N_4282);
and U7584 (N_7584,N_5368,N_4165);
xor U7585 (N_7585,N_4785,N_4697);
nor U7586 (N_7586,N_5657,N_4192);
or U7587 (N_7587,N_4517,N_5836);
nor U7588 (N_7588,N_5731,N_5533);
nand U7589 (N_7589,N_5396,N_5383);
nand U7590 (N_7590,N_5865,N_5545);
nand U7591 (N_7591,N_4067,N_4794);
nor U7592 (N_7592,N_4163,N_4082);
xnor U7593 (N_7593,N_5064,N_5019);
nor U7594 (N_7594,N_4874,N_5077);
or U7595 (N_7595,N_4632,N_5632);
and U7596 (N_7596,N_4113,N_4491);
and U7597 (N_7597,N_5612,N_5683);
or U7598 (N_7598,N_4990,N_5056);
or U7599 (N_7599,N_5813,N_5877);
nor U7600 (N_7600,N_5615,N_4619);
or U7601 (N_7601,N_4763,N_5890);
nor U7602 (N_7602,N_5696,N_5593);
or U7603 (N_7603,N_4103,N_4778);
and U7604 (N_7604,N_5017,N_4656);
xor U7605 (N_7605,N_5790,N_4191);
nand U7606 (N_7606,N_5464,N_4610);
nor U7607 (N_7607,N_5762,N_4402);
or U7608 (N_7608,N_5527,N_5688);
nor U7609 (N_7609,N_4301,N_4427);
nand U7610 (N_7610,N_5564,N_4915);
nor U7611 (N_7611,N_4532,N_4335);
or U7612 (N_7612,N_4373,N_5329);
nor U7613 (N_7613,N_4926,N_5619);
nor U7614 (N_7614,N_5601,N_4580);
and U7615 (N_7615,N_4286,N_4588);
or U7616 (N_7616,N_4428,N_4280);
and U7617 (N_7617,N_5324,N_5508);
and U7618 (N_7618,N_4157,N_4291);
and U7619 (N_7619,N_4773,N_5952);
or U7620 (N_7620,N_4632,N_5689);
nor U7621 (N_7621,N_5512,N_5864);
xor U7622 (N_7622,N_5379,N_5210);
nor U7623 (N_7623,N_4168,N_4912);
xnor U7624 (N_7624,N_5833,N_5589);
nor U7625 (N_7625,N_4239,N_5883);
and U7626 (N_7626,N_4717,N_5375);
or U7627 (N_7627,N_4072,N_4024);
or U7628 (N_7628,N_4208,N_5251);
nand U7629 (N_7629,N_4752,N_4155);
and U7630 (N_7630,N_5684,N_5879);
and U7631 (N_7631,N_4401,N_4943);
and U7632 (N_7632,N_4426,N_5401);
or U7633 (N_7633,N_5577,N_4750);
nand U7634 (N_7634,N_5485,N_4301);
and U7635 (N_7635,N_4888,N_5789);
and U7636 (N_7636,N_5050,N_5716);
nor U7637 (N_7637,N_4707,N_5050);
and U7638 (N_7638,N_5944,N_5410);
and U7639 (N_7639,N_5905,N_5627);
or U7640 (N_7640,N_4576,N_4791);
nor U7641 (N_7641,N_5612,N_5232);
nand U7642 (N_7642,N_5658,N_5469);
or U7643 (N_7643,N_5415,N_4336);
nand U7644 (N_7644,N_5853,N_4484);
and U7645 (N_7645,N_4861,N_4799);
nand U7646 (N_7646,N_4936,N_5533);
nand U7647 (N_7647,N_4087,N_5395);
xor U7648 (N_7648,N_4243,N_5925);
nand U7649 (N_7649,N_5071,N_5990);
nand U7650 (N_7650,N_4908,N_4597);
nor U7651 (N_7651,N_4405,N_5797);
or U7652 (N_7652,N_5081,N_4868);
or U7653 (N_7653,N_4089,N_4314);
nand U7654 (N_7654,N_4497,N_5200);
nor U7655 (N_7655,N_4814,N_5812);
nand U7656 (N_7656,N_5836,N_5810);
nor U7657 (N_7657,N_5543,N_5229);
nand U7658 (N_7658,N_5027,N_5397);
nand U7659 (N_7659,N_4616,N_5051);
nor U7660 (N_7660,N_4367,N_5692);
xor U7661 (N_7661,N_4053,N_5504);
or U7662 (N_7662,N_4638,N_5491);
nand U7663 (N_7663,N_4421,N_4095);
nor U7664 (N_7664,N_5594,N_4710);
or U7665 (N_7665,N_4761,N_5101);
nor U7666 (N_7666,N_5973,N_4537);
or U7667 (N_7667,N_4538,N_4934);
nor U7668 (N_7668,N_4470,N_4846);
xnor U7669 (N_7669,N_4285,N_5933);
nor U7670 (N_7670,N_5864,N_5900);
or U7671 (N_7671,N_5183,N_4855);
and U7672 (N_7672,N_4375,N_5826);
nor U7673 (N_7673,N_5895,N_4821);
and U7674 (N_7674,N_5860,N_5457);
nor U7675 (N_7675,N_4416,N_4173);
nand U7676 (N_7676,N_4812,N_4951);
nand U7677 (N_7677,N_4601,N_5035);
nor U7678 (N_7678,N_4453,N_4897);
and U7679 (N_7679,N_5112,N_5629);
or U7680 (N_7680,N_4168,N_4260);
nand U7681 (N_7681,N_5694,N_5022);
or U7682 (N_7682,N_5581,N_5062);
or U7683 (N_7683,N_5113,N_4850);
nand U7684 (N_7684,N_4361,N_4281);
nand U7685 (N_7685,N_4509,N_4381);
xnor U7686 (N_7686,N_4296,N_4425);
nand U7687 (N_7687,N_5687,N_5354);
and U7688 (N_7688,N_5217,N_5408);
nor U7689 (N_7689,N_5378,N_4704);
nor U7690 (N_7690,N_5047,N_5656);
nor U7691 (N_7691,N_5065,N_4271);
and U7692 (N_7692,N_4675,N_4333);
and U7693 (N_7693,N_4358,N_4381);
nor U7694 (N_7694,N_5318,N_5846);
nor U7695 (N_7695,N_4849,N_5214);
nand U7696 (N_7696,N_5032,N_4353);
xor U7697 (N_7697,N_4844,N_5384);
nor U7698 (N_7698,N_5214,N_4646);
nor U7699 (N_7699,N_4891,N_4512);
and U7700 (N_7700,N_5434,N_4858);
nand U7701 (N_7701,N_4919,N_5630);
nor U7702 (N_7702,N_5229,N_5843);
nor U7703 (N_7703,N_5018,N_5715);
nand U7704 (N_7704,N_5421,N_4167);
nand U7705 (N_7705,N_5341,N_4469);
and U7706 (N_7706,N_5219,N_5684);
and U7707 (N_7707,N_5896,N_5974);
or U7708 (N_7708,N_4472,N_5863);
xnor U7709 (N_7709,N_5983,N_5221);
nor U7710 (N_7710,N_4897,N_4494);
or U7711 (N_7711,N_4692,N_5613);
nor U7712 (N_7712,N_5679,N_5900);
and U7713 (N_7713,N_4699,N_5035);
nor U7714 (N_7714,N_5195,N_5861);
and U7715 (N_7715,N_5217,N_4941);
or U7716 (N_7716,N_5410,N_4057);
and U7717 (N_7717,N_5380,N_5345);
nand U7718 (N_7718,N_4320,N_5936);
or U7719 (N_7719,N_5242,N_4676);
and U7720 (N_7720,N_5029,N_4794);
or U7721 (N_7721,N_4518,N_4775);
nand U7722 (N_7722,N_4253,N_5636);
and U7723 (N_7723,N_5282,N_5216);
nor U7724 (N_7724,N_4555,N_4196);
nor U7725 (N_7725,N_5210,N_4734);
and U7726 (N_7726,N_5343,N_5328);
nor U7727 (N_7727,N_5701,N_5446);
or U7728 (N_7728,N_4937,N_5422);
nor U7729 (N_7729,N_5433,N_5738);
nand U7730 (N_7730,N_4873,N_4862);
or U7731 (N_7731,N_4991,N_4602);
and U7732 (N_7732,N_5736,N_4871);
nand U7733 (N_7733,N_4789,N_4465);
xnor U7734 (N_7734,N_5204,N_4876);
nand U7735 (N_7735,N_4584,N_5413);
and U7736 (N_7736,N_5585,N_4856);
or U7737 (N_7737,N_4698,N_5227);
nand U7738 (N_7738,N_5849,N_5648);
nand U7739 (N_7739,N_4757,N_5332);
or U7740 (N_7740,N_5844,N_4663);
nor U7741 (N_7741,N_4553,N_4036);
nand U7742 (N_7742,N_5724,N_5242);
or U7743 (N_7743,N_4667,N_5282);
or U7744 (N_7744,N_5921,N_4366);
xnor U7745 (N_7745,N_5404,N_5831);
and U7746 (N_7746,N_4213,N_5853);
nor U7747 (N_7747,N_4878,N_5596);
nand U7748 (N_7748,N_4509,N_4139);
nand U7749 (N_7749,N_5400,N_4666);
or U7750 (N_7750,N_4206,N_4084);
nor U7751 (N_7751,N_5634,N_4009);
nor U7752 (N_7752,N_5241,N_4892);
or U7753 (N_7753,N_4618,N_5222);
nor U7754 (N_7754,N_5584,N_5804);
nor U7755 (N_7755,N_4837,N_4769);
and U7756 (N_7756,N_5755,N_4739);
nand U7757 (N_7757,N_4502,N_5462);
nand U7758 (N_7758,N_4150,N_4214);
or U7759 (N_7759,N_4865,N_5034);
or U7760 (N_7760,N_5194,N_4265);
nand U7761 (N_7761,N_4053,N_5856);
or U7762 (N_7762,N_5066,N_4444);
nor U7763 (N_7763,N_5355,N_5362);
nand U7764 (N_7764,N_4072,N_4229);
nor U7765 (N_7765,N_4180,N_5979);
or U7766 (N_7766,N_5805,N_5283);
or U7767 (N_7767,N_4236,N_4016);
or U7768 (N_7768,N_4289,N_4578);
nor U7769 (N_7769,N_5074,N_4538);
or U7770 (N_7770,N_5211,N_5496);
nand U7771 (N_7771,N_4680,N_5187);
nand U7772 (N_7772,N_4599,N_4946);
nand U7773 (N_7773,N_5366,N_5959);
and U7774 (N_7774,N_5830,N_4103);
xnor U7775 (N_7775,N_4783,N_5536);
nand U7776 (N_7776,N_4773,N_4063);
xnor U7777 (N_7777,N_4771,N_5234);
nor U7778 (N_7778,N_5026,N_5700);
and U7779 (N_7779,N_5872,N_5512);
nand U7780 (N_7780,N_5136,N_4894);
nand U7781 (N_7781,N_5519,N_5918);
nor U7782 (N_7782,N_4052,N_5692);
nor U7783 (N_7783,N_5751,N_4454);
nand U7784 (N_7784,N_5907,N_4013);
and U7785 (N_7785,N_5226,N_5601);
nand U7786 (N_7786,N_4247,N_5152);
nor U7787 (N_7787,N_5704,N_5961);
nor U7788 (N_7788,N_4386,N_5713);
nor U7789 (N_7789,N_5325,N_5708);
and U7790 (N_7790,N_5997,N_4459);
or U7791 (N_7791,N_4046,N_5127);
and U7792 (N_7792,N_5084,N_5534);
and U7793 (N_7793,N_4589,N_5792);
nor U7794 (N_7794,N_5930,N_4798);
nand U7795 (N_7795,N_4515,N_4317);
or U7796 (N_7796,N_4394,N_4184);
and U7797 (N_7797,N_4344,N_4705);
or U7798 (N_7798,N_5326,N_5906);
and U7799 (N_7799,N_4066,N_5830);
nand U7800 (N_7800,N_5401,N_5687);
xnor U7801 (N_7801,N_4444,N_5561);
nor U7802 (N_7802,N_4619,N_4382);
nand U7803 (N_7803,N_5407,N_5873);
nor U7804 (N_7804,N_4166,N_5820);
nand U7805 (N_7805,N_4958,N_4205);
or U7806 (N_7806,N_5968,N_4166);
and U7807 (N_7807,N_4785,N_5852);
nor U7808 (N_7808,N_4525,N_4633);
or U7809 (N_7809,N_5918,N_4500);
and U7810 (N_7810,N_5416,N_5551);
and U7811 (N_7811,N_4858,N_5697);
nand U7812 (N_7812,N_5489,N_5278);
or U7813 (N_7813,N_5677,N_5245);
xor U7814 (N_7814,N_5676,N_4726);
xnor U7815 (N_7815,N_4526,N_4627);
nand U7816 (N_7816,N_4309,N_5588);
and U7817 (N_7817,N_5892,N_5216);
or U7818 (N_7818,N_5169,N_4405);
or U7819 (N_7819,N_4840,N_4258);
and U7820 (N_7820,N_4022,N_4273);
and U7821 (N_7821,N_5255,N_4905);
and U7822 (N_7822,N_5239,N_5449);
and U7823 (N_7823,N_5230,N_4205);
nor U7824 (N_7824,N_4312,N_5399);
xnor U7825 (N_7825,N_5116,N_4714);
nor U7826 (N_7826,N_5811,N_4238);
or U7827 (N_7827,N_4867,N_4499);
xnor U7828 (N_7828,N_4412,N_4478);
nor U7829 (N_7829,N_5407,N_5021);
nand U7830 (N_7830,N_4485,N_4110);
and U7831 (N_7831,N_4250,N_4747);
and U7832 (N_7832,N_5285,N_5570);
nand U7833 (N_7833,N_4040,N_5749);
nand U7834 (N_7834,N_5335,N_4395);
or U7835 (N_7835,N_4297,N_5917);
and U7836 (N_7836,N_5262,N_4491);
nand U7837 (N_7837,N_5490,N_4193);
xnor U7838 (N_7838,N_4255,N_4319);
and U7839 (N_7839,N_4164,N_5748);
and U7840 (N_7840,N_5175,N_4471);
nor U7841 (N_7841,N_4957,N_5055);
or U7842 (N_7842,N_5492,N_4836);
nand U7843 (N_7843,N_5485,N_4416);
nand U7844 (N_7844,N_4343,N_5869);
or U7845 (N_7845,N_5929,N_4612);
or U7846 (N_7846,N_4934,N_5481);
nand U7847 (N_7847,N_5233,N_5499);
and U7848 (N_7848,N_4052,N_4168);
nor U7849 (N_7849,N_4273,N_5093);
or U7850 (N_7850,N_4764,N_4448);
nand U7851 (N_7851,N_4670,N_5957);
nand U7852 (N_7852,N_5143,N_4215);
nand U7853 (N_7853,N_5362,N_4803);
nand U7854 (N_7854,N_4845,N_4364);
nor U7855 (N_7855,N_5972,N_5021);
nand U7856 (N_7856,N_4871,N_4829);
nand U7857 (N_7857,N_5478,N_4379);
and U7858 (N_7858,N_5178,N_4007);
and U7859 (N_7859,N_4681,N_4739);
nand U7860 (N_7860,N_4320,N_5188);
or U7861 (N_7861,N_5814,N_5253);
xor U7862 (N_7862,N_4279,N_5138);
nand U7863 (N_7863,N_4506,N_5797);
nor U7864 (N_7864,N_4088,N_5333);
and U7865 (N_7865,N_5717,N_5750);
xor U7866 (N_7866,N_5358,N_4061);
nand U7867 (N_7867,N_5470,N_5436);
nand U7868 (N_7868,N_4786,N_4500);
and U7869 (N_7869,N_4678,N_4939);
and U7870 (N_7870,N_5040,N_4833);
nand U7871 (N_7871,N_4556,N_5854);
nand U7872 (N_7872,N_4360,N_4088);
and U7873 (N_7873,N_4682,N_4572);
nand U7874 (N_7874,N_5501,N_5115);
and U7875 (N_7875,N_5293,N_5777);
or U7876 (N_7876,N_5912,N_4410);
nor U7877 (N_7877,N_4540,N_4460);
nand U7878 (N_7878,N_5239,N_5318);
nand U7879 (N_7879,N_5801,N_4162);
nor U7880 (N_7880,N_5580,N_4483);
and U7881 (N_7881,N_5325,N_5961);
and U7882 (N_7882,N_4667,N_4209);
and U7883 (N_7883,N_5744,N_5929);
nand U7884 (N_7884,N_4853,N_4010);
nor U7885 (N_7885,N_4897,N_4709);
nor U7886 (N_7886,N_5625,N_5518);
xor U7887 (N_7887,N_4446,N_4595);
nand U7888 (N_7888,N_5663,N_5482);
or U7889 (N_7889,N_4273,N_5978);
nor U7890 (N_7890,N_5301,N_4137);
xor U7891 (N_7891,N_5924,N_5837);
or U7892 (N_7892,N_5422,N_5299);
nor U7893 (N_7893,N_4927,N_4391);
and U7894 (N_7894,N_4329,N_5884);
nand U7895 (N_7895,N_4673,N_5992);
nor U7896 (N_7896,N_5110,N_5922);
nand U7897 (N_7897,N_5307,N_4090);
xor U7898 (N_7898,N_4599,N_4702);
nand U7899 (N_7899,N_4425,N_4345);
and U7900 (N_7900,N_5732,N_5626);
and U7901 (N_7901,N_4965,N_4602);
nor U7902 (N_7902,N_5346,N_4218);
nor U7903 (N_7903,N_5778,N_5870);
nor U7904 (N_7904,N_5994,N_5316);
xnor U7905 (N_7905,N_5700,N_4323);
or U7906 (N_7906,N_5010,N_5003);
nand U7907 (N_7907,N_4076,N_5166);
and U7908 (N_7908,N_5235,N_4649);
or U7909 (N_7909,N_5167,N_5537);
and U7910 (N_7910,N_5665,N_5127);
nand U7911 (N_7911,N_5949,N_4351);
and U7912 (N_7912,N_5813,N_5054);
nand U7913 (N_7913,N_5925,N_5760);
nor U7914 (N_7914,N_4953,N_5594);
nand U7915 (N_7915,N_4164,N_5311);
and U7916 (N_7916,N_4276,N_5399);
nor U7917 (N_7917,N_4306,N_5215);
and U7918 (N_7918,N_5336,N_4682);
nand U7919 (N_7919,N_5745,N_4988);
xor U7920 (N_7920,N_5190,N_4492);
nand U7921 (N_7921,N_5409,N_4997);
and U7922 (N_7922,N_5092,N_5805);
and U7923 (N_7923,N_5403,N_5237);
or U7924 (N_7924,N_5245,N_4301);
nor U7925 (N_7925,N_4144,N_5686);
nand U7926 (N_7926,N_4931,N_4359);
nand U7927 (N_7927,N_4262,N_4281);
nand U7928 (N_7928,N_4154,N_5201);
or U7929 (N_7929,N_5392,N_5655);
nand U7930 (N_7930,N_4421,N_4591);
or U7931 (N_7931,N_4169,N_4328);
xnor U7932 (N_7932,N_5925,N_5200);
nand U7933 (N_7933,N_5422,N_5606);
xor U7934 (N_7934,N_5521,N_4295);
and U7935 (N_7935,N_4322,N_4390);
and U7936 (N_7936,N_4910,N_5355);
nor U7937 (N_7937,N_5922,N_4743);
xnor U7938 (N_7938,N_5367,N_4976);
xnor U7939 (N_7939,N_5135,N_5303);
xor U7940 (N_7940,N_5082,N_5388);
or U7941 (N_7941,N_4495,N_5787);
nand U7942 (N_7942,N_5977,N_5840);
xor U7943 (N_7943,N_4738,N_5077);
nor U7944 (N_7944,N_5109,N_4087);
xnor U7945 (N_7945,N_4753,N_5170);
nor U7946 (N_7946,N_5257,N_5140);
nor U7947 (N_7947,N_5603,N_4982);
or U7948 (N_7948,N_4085,N_5772);
and U7949 (N_7949,N_4188,N_4079);
nor U7950 (N_7950,N_5449,N_5651);
nor U7951 (N_7951,N_5177,N_4051);
and U7952 (N_7952,N_5476,N_4402);
xor U7953 (N_7953,N_4053,N_4039);
nor U7954 (N_7954,N_4726,N_4652);
and U7955 (N_7955,N_5303,N_5008);
nor U7956 (N_7956,N_5168,N_4785);
nand U7957 (N_7957,N_5879,N_4830);
nand U7958 (N_7958,N_5732,N_4328);
nand U7959 (N_7959,N_4714,N_4095);
nand U7960 (N_7960,N_4246,N_5611);
or U7961 (N_7961,N_4313,N_5857);
or U7962 (N_7962,N_5116,N_5910);
nor U7963 (N_7963,N_4187,N_5856);
xor U7964 (N_7964,N_5911,N_4931);
and U7965 (N_7965,N_4129,N_4716);
and U7966 (N_7966,N_4706,N_4746);
nor U7967 (N_7967,N_4826,N_4151);
or U7968 (N_7968,N_5784,N_5021);
nand U7969 (N_7969,N_4424,N_5981);
nor U7970 (N_7970,N_4571,N_5934);
nor U7971 (N_7971,N_5062,N_5299);
and U7972 (N_7972,N_5778,N_4462);
and U7973 (N_7973,N_4950,N_4084);
and U7974 (N_7974,N_5959,N_5849);
or U7975 (N_7975,N_4527,N_4725);
or U7976 (N_7976,N_5829,N_5679);
nand U7977 (N_7977,N_4179,N_4293);
xor U7978 (N_7978,N_5211,N_5232);
nor U7979 (N_7979,N_5802,N_4668);
nor U7980 (N_7980,N_5783,N_5417);
and U7981 (N_7981,N_5548,N_5650);
nand U7982 (N_7982,N_4894,N_5531);
and U7983 (N_7983,N_4412,N_5701);
nand U7984 (N_7984,N_5776,N_4694);
nand U7985 (N_7985,N_5040,N_4243);
or U7986 (N_7986,N_5516,N_5950);
xnor U7987 (N_7987,N_4710,N_5377);
nand U7988 (N_7988,N_5889,N_4137);
or U7989 (N_7989,N_4116,N_4103);
nand U7990 (N_7990,N_4716,N_4832);
nand U7991 (N_7991,N_4996,N_4375);
or U7992 (N_7992,N_4931,N_5564);
nand U7993 (N_7993,N_5679,N_5376);
and U7994 (N_7994,N_4718,N_5254);
or U7995 (N_7995,N_4631,N_5804);
or U7996 (N_7996,N_5711,N_5078);
nand U7997 (N_7997,N_5684,N_4743);
nor U7998 (N_7998,N_4938,N_4253);
nand U7999 (N_7999,N_5697,N_5086);
and U8000 (N_8000,N_7872,N_7267);
xnor U8001 (N_8001,N_7830,N_7932);
nor U8002 (N_8002,N_7054,N_6027);
nor U8003 (N_8003,N_6530,N_6589);
and U8004 (N_8004,N_6470,N_6540);
xnor U8005 (N_8005,N_6856,N_7100);
or U8006 (N_8006,N_7404,N_7888);
nor U8007 (N_8007,N_7560,N_6384);
nor U8008 (N_8008,N_6817,N_6534);
nand U8009 (N_8009,N_6863,N_7575);
or U8010 (N_8010,N_6621,N_7491);
and U8011 (N_8011,N_7162,N_6999);
and U8012 (N_8012,N_6190,N_7539);
nand U8013 (N_8013,N_6899,N_6898);
xnor U8014 (N_8014,N_6580,N_7765);
or U8015 (N_8015,N_7989,N_7795);
or U8016 (N_8016,N_6373,N_6194);
or U8017 (N_8017,N_6598,N_6519);
or U8018 (N_8018,N_7704,N_6441);
and U8019 (N_8019,N_7327,N_6691);
or U8020 (N_8020,N_7648,N_6093);
and U8021 (N_8021,N_7150,N_7415);
xor U8022 (N_8022,N_7758,N_7687);
nor U8023 (N_8023,N_6121,N_6778);
nand U8024 (N_8024,N_6002,N_6904);
nand U8025 (N_8025,N_6884,N_6711);
nor U8026 (N_8026,N_6106,N_6088);
nor U8027 (N_8027,N_6791,N_6879);
nor U8028 (N_8028,N_6520,N_7558);
nand U8029 (N_8029,N_7483,N_7307);
and U8030 (N_8030,N_6703,N_6340);
or U8031 (N_8031,N_7818,N_6537);
nand U8032 (N_8032,N_7836,N_6498);
nand U8033 (N_8033,N_7445,N_6390);
or U8034 (N_8034,N_7835,N_7735);
and U8035 (N_8035,N_6684,N_7520);
or U8036 (N_8036,N_7407,N_7925);
and U8037 (N_8037,N_7416,N_6793);
or U8038 (N_8038,N_6569,N_6776);
and U8039 (N_8039,N_6171,N_6212);
and U8040 (N_8040,N_7188,N_7832);
nand U8041 (N_8041,N_7623,N_7330);
nor U8042 (N_8042,N_7079,N_6686);
nor U8043 (N_8043,N_6773,N_7695);
xor U8044 (N_8044,N_6451,N_6921);
xor U8045 (N_8045,N_7303,N_7672);
nand U8046 (N_8046,N_6262,N_7331);
or U8047 (N_8047,N_6085,N_6913);
nor U8048 (N_8048,N_6436,N_7196);
and U8049 (N_8049,N_7663,N_7841);
or U8050 (N_8050,N_7650,N_7442);
nand U8051 (N_8051,N_6582,N_7905);
nor U8052 (N_8052,N_7427,N_6414);
xor U8053 (N_8053,N_7502,N_7349);
nand U8054 (N_8054,N_6443,N_6374);
or U8055 (N_8055,N_7801,N_6061);
and U8056 (N_8056,N_6227,N_6766);
nor U8057 (N_8057,N_7897,N_7063);
or U8058 (N_8058,N_6523,N_6949);
or U8059 (N_8059,N_7840,N_7059);
nand U8060 (N_8060,N_7955,N_7958);
and U8061 (N_8061,N_7742,N_7856);
nor U8062 (N_8062,N_6463,N_6702);
nor U8063 (N_8063,N_7165,N_7454);
nand U8064 (N_8064,N_6077,N_7475);
and U8065 (N_8065,N_6364,N_6039);
nand U8066 (N_8066,N_7712,N_7133);
xor U8067 (N_8067,N_6597,N_6479);
and U8068 (N_8068,N_6063,N_7292);
or U8069 (N_8069,N_7459,N_7045);
nand U8070 (N_8070,N_7523,N_6885);
nor U8071 (N_8071,N_6539,N_6930);
nand U8072 (N_8072,N_7264,N_6031);
nor U8073 (N_8073,N_7305,N_6825);
and U8074 (N_8074,N_7018,N_7366);
or U8075 (N_8075,N_7394,N_7340);
and U8076 (N_8076,N_6193,N_7012);
nor U8077 (N_8077,N_6561,N_7437);
and U8078 (N_8078,N_6386,N_6416);
nand U8079 (N_8079,N_7392,N_6440);
or U8080 (N_8080,N_7641,N_6992);
or U8081 (N_8081,N_6634,N_6342);
nor U8082 (N_8082,N_6272,N_6016);
and U8083 (N_8083,N_6599,N_7482);
nor U8084 (N_8084,N_6465,N_6292);
or U8085 (N_8085,N_6152,N_7492);
or U8086 (N_8086,N_6348,N_7852);
and U8087 (N_8087,N_7291,N_7875);
nand U8088 (N_8088,N_6248,N_7730);
nor U8089 (N_8089,N_6285,N_6818);
nand U8090 (N_8090,N_7581,N_7721);
nor U8091 (N_8091,N_7511,N_7545);
nor U8092 (N_8092,N_7904,N_7250);
and U8093 (N_8093,N_7821,N_7791);
nor U8094 (N_8094,N_6464,N_6681);
nor U8095 (N_8095,N_7725,N_6835);
or U8096 (N_8096,N_6727,N_6293);
nand U8097 (N_8097,N_7919,N_7122);
or U8098 (N_8098,N_7660,N_7766);
nand U8099 (N_8099,N_7317,N_6758);
and U8100 (N_8100,N_6720,N_7943);
nor U8101 (N_8101,N_6586,N_7743);
nor U8102 (N_8102,N_7334,N_7974);
nand U8103 (N_8103,N_6795,N_7887);
and U8104 (N_8104,N_7049,N_7177);
or U8105 (N_8105,N_6485,N_6286);
xor U8106 (N_8106,N_6560,N_7175);
nor U8107 (N_8107,N_7803,N_6244);
nor U8108 (N_8108,N_7751,N_6705);
or U8109 (N_8109,N_7859,N_6455);
xor U8110 (N_8110,N_7684,N_7574);
and U8111 (N_8111,N_6779,N_6654);
or U8112 (N_8112,N_7044,N_7301);
or U8113 (N_8113,N_6546,N_6174);
and U8114 (N_8114,N_7608,N_7106);
or U8115 (N_8115,N_7253,N_6336);
nand U8116 (N_8116,N_6224,N_7813);
nand U8117 (N_8117,N_6626,N_6315);
xor U8118 (N_8118,N_7195,N_7135);
and U8119 (N_8119,N_7733,N_7024);
nand U8120 (N_8120,N_7249,N_7046);
nand U8121 (N_8121,N_6048,N_7233);
or U8122 (N_8122,N_6933,N_7970);
nand U8123 (N_8123,N_7453,N_6697);
and U8124 (N_8124,N_7134,N_6594);
xnor U8125 (N_8125,N_7747,N_6273);
or U8126 (N_8126,N_6247,N_7469);
and U8127 (N_8127,N_6263,N_7048);
nor U8128 (N_8128,N_7089,N_7361);
nand U8129 (N_8129,N_6944,N_6217);
nand U8130 (N_8130,N_7898,N_6346);
or U8131 (N_8131,N_6585,N_6721);
or U8132 (N_8132,N_7644,N_7076);
or U8133 (N_8133,N_7779,N_7972);
xor U8134 (N_8134,N_6310,N_7473);
nand U8135 (N_8135,N_7886,N_6046);
or U8136 (N_8136,N_7506,N_6158);
nand U8137 (N_8137,N_6764,N_7744);
nor U8138 (N_8138,N_6499,N_7908);
nand U8139 (N_8139,N_6723,N_6305);
nor U8140 (N_8140,N_6985,N_6869);
or U8141 (N_8141,N_7713,N_6641);
xor U8142 (N_8142,N_7971,N_6802);
xnor U8143 (N_8143,N_7153,N_6968);
nand U8144 (N_8144,N_7595,N_7983);
nand U8145 (N_8145,N_6090,N_7705);
nand U8146 (N_8146,N_7441,N_6735);
or U8147 (N_8147,N_7701,N_6369);
nor U8148 (N_8148,N_6919,N_7551);
nor U8149 (N_8149,N_7168,N_6494);
nor U8150 (N_8150,N_7975,N_7325);
or U8151 (N_8151,N_7164,N_6722);
nand U8152 (N_8152,N_6839,N_6553);
or U8153 (N_8153,N_7927,N_6145);
nor U8154 (N_8154,N_7521,N_7808);
or U8155 (N_8155,N_6394,N_6907);
nor U8156 (N_8156,N_6730,N_7239);
and U8157 (N_8157,N_7893,N_6886);
nand U8158 (N_8158,N_6640,N_7745);
and U8159 (N_8159,N_6562,N_6759);
nor U8160 (N_8160,N_7885,N_7774);
nand U8161 (N_8161,N_7834,N_7496);
and U8162 (N_8162,N_6089,N_6491);
nand U8163 (N_8163,N_7375,N_6118);
xnor U8164 (N_8164,N_6929,N_7771);
nand U8165 (N_8165,N_6945,N_7411);
nor U8166 (N_8166,N_7388,N_7959);
nand U8167 (N_8167,N_7238,N_7023);
nor U8168 (N_8168,N_6051,N_7467);
or U8169 (N_8169,N_6495,N_6125);
nor U8170 (N_8170,N_6277,N_7902);
nor U8171 (N_8171,N_6237,N_6922);
xor U8172 (N_8172,N_6829,N_6209);
or U8173 (N_8173,N_7583,N_6148);
nand U8174 (N_8174,N_6662,N_6876);
or U8175 (N_8175,N_7287,N_7103);
and U8176 (N_8176,N_7155,N_7259);
nor U8177 (N_8177,N_6325,N_6801);
nor U8178 (N_8178,N_6500,N_7444);
nor U8179 (N_8179,N_7058,N_7549);
or U8180 (N_8180,N_7669,N_6505);
nor U8181 (N_8181,N_6532,N_6117);
or U8182 (N_8182,N_7537,N_6830);
nor U8183 (N_8183,N_7617,N_6207);
nand U8184 (N_8184,N_6184,N_7866);
or U8185 (N_8185,N_6600,N_6350);
or U8186 (N_8186,N_6573,N_6756);
nor U8187 (N_8187,N_6476,N_7081);
nand U8188 (N_8188,N_7697,N_6630);
nand U8189 (N_8189,N_6814,N_7591);
and U8190 (N_8190,N_6317,N_6381);
and U8191 (N_8191,N_6078,N_6159);
or U8192 (N_8192,N_6535,N_7268);
nand U8193 (N_8193,N_6368,N_6412);
and U8194 (N_8194,N_7720,N_6484);
nand U8195 (N_8195,N_7215,N_7128);
nand U8196 (N_8196,N_6264,N_7376);
or U8197 (N_8197,N_6216,N_6055);
nand U8198 (N_8198,N_6322,N_7691);
nor U8199 (N_8199,N_7992,N_6877);
nor U8200 (N_8200,N_7481,N_6213);
nor U8201 (N_8201,N_7001,N_6983);
nor U8202 (N_8202,N_6805,N_6755);
and U8203 (N_8203,N_6139,N_6777);
nand U8204 (N_8204,N_6204,N_6775);
xnor U8205 (N_8205,N_6425,N_7082);
nor U8206 (N_8206,N_6229,N_7739);
and U8207 (N_8207,N_6618,N_7169);
xor U8208 (N_8208,N_7555,N_6417);
or U8209 (N_8209,N_7172,N_6296);
or U8210 (N_8210,N_7881,N_6780);
nor U8211 (N_8211,N_6220,N_7263);
nor U8212 (N_8212,N_6281,N_7039);
or U8213 (N_8213,N_7752,N_7759);
nand U8214 (N_8214,N_7967,N_6636);
or U8215 (N_8215,N_6757,N_7786);
xor U8216 (N_8216,N_7588,N_6896);
nand U8217 (N_8217,N_6187,N_7614);
or U8218 (N_8218,N_7863,N_7230);
nand U8219 (N_8219,N_6351,N_6150);
nor U8220 (N_8220,N_7200,N_6013);
and U8221 (N_8221,N_7719,N_7275);
and U8222 (N_8222,N_7677,N_7316);
and U8223 (N_8223,N_7220,N_6632);
nor U8224 (N_8224,N_7912,N_6864);
nor U8225 (N_8225,N_7027,N_7016);
nand U8226 (N_8226,N_6713,N_6254);
nor U8227 (N_8227,N_7569,N_7136);
nor U8228 (N_8228,N_6717,N_6897);
nand U8229 (N_8229,N_7386,N_6620);
and U8230 (N_8230,N_6076,N_6927);
nor U8231 (N_8231,N_7530,N_7903);
nand U8232 (N_8232,N_7728,N_6045);
nand U8233 (N_8233,N_7304,N_7393);
or U8234 (N_8234,N_6866,N_7116);
and U8235 (N_8235,N_6669,N_7013);
nand U8236 (N_8236,N_7084,N_7382);
nor U8237 (N_8237,N_7211,N_6134);
or U8238 (N_8238,N_6821,N_6307);
nor U8239 (N_8239,N_7668,N_7746);
or U8240 (N_8240,N_6813,N_7829);
xor U8241 (N_8241,N_6741,N_6496);
or U8242 (N_8242,N_6265,N_6136);
nor U8243 (N_8243,N_7201,N_7546);
or U8244 (N_8244,N_7618,N_6107);
nor U8245 (N_8245,N_7104,N_6306);
nand U8246 (N_8246,N_6564,N_7005);
nor U8247 (N_8247,N_7159,N_6060);
nand U8248 (N_8248,N_6257,N_6129);
nor U8249 (N_8249,N_6402,N_6453);
and U8250 (N_8250,N_7517,N_7942);
xor U8251 (N_8251,N_6643,N_7440);
nor U8252 (N_8252,N_6993,N_7675);
or U8253 (N_8253,N_7602,N_7237);
and U8254 (N_8254,N_6882,N_7525);
and U8255 (N_8255,N_6708,N_7399);
or U8256 (N_8256,N_6943,N_6393);
or U8257 (N_8257,N_7026,N_7799);
and U8258 (N_8258,N_7360,N_7065);
xor U8259 (N_8259,N_6043,N_7564);
nand U8260 (N_8260,N_6124,N_6831);
and U8261 (N_8261,N_7274,N_7861);
or U8262 (N_8262,N_6178,N_7205);
nand U8263 (N_8263,N_6895,N_7508);
nor U8264 (N_8264,N_6410,N_6951);
or U8265 (N_8265,N_7183,N_7993);
and U8266 (N_8266,N_6144,N_7251);
or U8267 (N_8267,N_7212,N_7838);
xor U8268 (N_8268,N_7086,N_7178);
or U8269 (N_8269,N_7369,N_6069);
nor U8270 (N_8270,N_7466,N_7014);
and U8271 (N_8271,N_6925,N_6177);
and U8272 (N_8272,N_7527,N_6682);
or U8273 (N_8273,N_6892,N_6788);
xnor U8274 (N_8274,N_6923,N_6784);
or U8275 (N_8275,N_7500,N_7718);
and U8276 (N_8276,N_6188,N_6131);
nand U8277 (N_8277,N_6047,N_7869);
nand U8278 (N_8278,N_7002,N_7882);
nand U8279 (N_8279,N_6926,N_6937);
or U8280 (N_8280,N_6415,N_7804);
xor U8281 (N_8281,N_6312,N_6575);
nand U8282 (N_8282,N_6473,N_6744);
or U8283 (N_8283,N_7649,N_7538);
or U8284 (N_8284,N_7413,N_7387);
or U8285 (N_8285,N_7101,N_7157);
or U8286 (N_8286,N_7348,N_6023);
nor U8287 (N_8287,N_6673,N_7810);
nor U8288 (N_8288,N_6460,N_6406);
nand U8289 (N_8289,N_7928,N_6710);
nand U8290 (N_8290,N_6041,N_7734);
and U8291 (N_8291,N_6649,N_6297);
nor U8292 (N_8292,N_6071,N_6628);
or U8293 (N_8293,N_7910,N_6541);
nand U8294 (N_8294,N_7278,N_7161);
nand U8295 (N_8295,N_7359,N_7607);
and U8296 (N_8296,N_6397,N_6311);
nand U8297 (N_8297,N_6001,N_6003);
and U8298 (N_8298,N_7221,N_7571);
or U8299 (N_8299,N_6309,N_6082);
nand U8300 (N_8300,N_7390,N_7032);
nand U8301 (N_8301,N_6872,N_7067);
or U8302 (N_8302,N_6400,N_6008);
xnor U8303 (N_8303,N_6672,N_7532);
nor U8304 (N_8304,N_6267,N_6080);
or U8305 (N_8305,N_6972,N_6854);
nor U8306 (N_8306,N_6555,N_6191);
nand U8307 (N_8307,N_7356,N_6276);
and U8308 (N_8308,N_7289,N_6081);
and U8309 (N_8309,N_7671,N_7290);
nand U8310 (N_8310,N_6870,N_6770);
and U8311 (N_8311,N_6005,N_7029);
or U8312 (N_8312,N_6957,N_6239);
and U8313 (N_8313,N_7916,N_6221);
nand U8314 (N_8314,N_6512,N_7339);
nand U8315 (N_8315,N_6631,N_7794);
and U8316 (N_8316,N_7884,N_7710);
nor U8317 (N_8317,N_7954,N_6963);
xnor U8318 (N_8318,N_6062,N_6798);
nand U8319 (N_8319,N_7913,N_7606);
nand U8320 (N_8320,N_7191,N_6362);
nor U8321 (N_8321,N_7722,N_7842);
nand U8322 (N_8322,N_7022,N_7812);
and U8323 (N_8323,N_6576,N_7590);
nand U8324 (N_8324,N_6889,N_6396);
or U8325 (N_8325,N_6423,N_6570);
or U8326 (N_8326,N_6344,N_7658);
nand U8327 (N_8327,N_7383,N_7900);
nor U8328 (N_8328,N_7344,N_6427);
and U8329 (N_8329,N_6568,N_6677);
nand U8330 (N_8330,N_6100,N_6235);
and U8331 (N_8331,N_6971,N_7978);
nand U8332 (N_8332,N_7341,N_7245);
nor U8333 (N_8333,N_7430,N_6616);
nand U8334 (N_8334,N_7034,N_6719);
nor U8335 (N_8335,N_6624,N_6210);
xor U8336 (N_8336,N_7934,N_6750);
and U8337 (N_8337,N_7613,N_6995);
nand U8338 (N_8338,N_7040,N_6301);
or U8339 (N_8339,N_7146,N_6444);
nor U8340 (N_8340,N_7503,N_6249);
nor U8341 (N_8341,N_6961,N_6280);
nand U8342 (N_8342,N_7306,N_7960);
xnor U8343 (N_8343,N_6429,N_6909);
and U8344 (N_8344,N_6170,N_6132);
nor U8345 (N_8345,N_7640,N_7938);
and U8346 (N_8346,N_6875,N_7909);
nor U8347 (N_8347,N_7347,N_6138);
or U8348 (N_8348,N_7137,N_7785);
nor U8349 (N_8349,N_7389,N_6675);
nor U8350 (N_8350,N_7541,N_6743);
xnor U8351 (N_8351,N_6493,N_7682);
xor U8352 (N_8352,N_7846,N_7163);
and U8353 (N_8353,N_7333,N_6180);
nand U8354 (N_8354,N_6695,N_6932);
and U8355 (N_8355,N_6371,N_6724);
nor U8356 (N_8356,N_6053,N_6327);
or U8357 (N_8357,N_7072,N_7624);
or U8358 (N_8358,N_7543,N_7561);
or U8359 (N_8359,N_7457,N_6516);
nor U8360 (N_8360,N_7255,N_7206);
and U8361 (N_8361,N_6857,N_6574);
xor U8362 (N_8362,N_7033,N_7901);
and U8363 (N_8363,N_7015,N_6940);
and U8364 (N_8364,N_6732,N_7055);
nand U8365 (N_8365,N_6075,N_6664);
nand U8366 (N_8366,N_6282,N_7185);
and U8367 (N_8367,N_6014,N_7851);
xor U8368 (N_8368,N_7513,N_6067);
and U8369 (N_8369,N_6608,N_7957);
and U8370 (N_8370,N_6915,N_7817);
xor U8371 (N_8371,N_7408,N_7228);
and U8372 (N_8372,N_6967,N_7160);
or U8373 (N_8373,N_7585,N_6647);
or U8374 (N_8374,N_6855,N_6324);
xor U8375 (N_8375,N_6328,N_7664);
and U8376 (N_8376,N_7662,N_6119);
or U8377 (N_8377,N_7035,N_6462);
or U8378 (N_8378,N_6948,N_6592);
nand U8379 (N_8379,N_7921,N_6823);
and U8380 (N_8380,N_6991,N_7401);
or U8381 (N_8381,N_7962,N_6611);
and U8382 (N_8382,N_7770,N_7936);
nand U8383 (N_8383,N_7423,N_6032);
nand U8384 (N_8384,N_7284,N_6827);
and U8385 (N_8385,N_7111,N_6038);
and U8386 (N_8386,N_6652,N_6973);
nand U8387 (N_8387,N_6057,N_6034);
nor U8388 (N_8388,N_6183,N_7659);
nand U8389 (N_8389,N_6728,N_6389);
and U8390 (N_8390,N_6116,N_7820);
or U8391 (N_8391,N_6469,N_6303);
nand U8392 (N_8392,N_6474,N_6467);
or U8393 (N_8393,N_7207,N_6753);
or U8394 (N_8394,N_7805,N_6841);
or U8395 (N_8395,N_7158,N_7777);
nand U8396 (N_8396,N_7793,N_6481);
nand U8397 (N_8397,N_7977,N_6054);
and U8398 (N_8398,N_7008,N_7519);
and U8399 (N_8399,N_6786,N_6357);
nor U8400 (N_8400,N_7850,N_6769);
or U8401 (N_8401,N_7980,N_6881);
nor U8402 (N_8402,N_6980,N_6650);
nor U8403 (N_8403,N_7198,N_6323);
nand U8404 (N_8404,N_6906,N_7999);
nand U8405 (N_8405,N_7688,N_6095);
or U8406 (N_8406,N_7295,N_7199);
and U8407 (N_8407,N_7933,N_7309);
xnor U8408 (N_8408,N_7748,N_7003);
xor U8409 (N_8409,N_6151,N_7286);
nand U8410 (N_8410,N_7764,N_7092);
and U8411 (N_8411,N_6147,N_7180);
or U8412 (N_8412,N_6782,N_7531);
nand U8413 (N_8413,N_7112,N_7579);
nor U8414 (N_8414,N_7935,N_6223);
nand U8415 (N_8415,N_6536,N_7406);
or U8416 (N_8416,N_7576,N_7000);
and U8417 (N_8417,N_7941,N_7709);
or U8418 (N_8418,N_7243,N_7310);
xnor U8419 (N_8419,N_6994,N_7918);
and U8420 (N_8420,N_6359,N_7378);
and U8421 (N_8421,N_6914,N_6517);
and U8422 (N_8422,N_7964,N_7920);
xnor U8423 (N_8423,N_6887,N_6299);
xnor U8424 (N_8424,N_7610,N_7297);
nor U8425 (N_8425,N_6800,N_7057);
xnor U8426 (N_8426,N_6487,N_6288);
xnor U8427 (N_8427,N_6928,N_6842);
nor U8428 (N_8428,N_6321,N_6326);
or U8429 (N_8429,N_7767,N_6225);
and U8430 (N_8430,N_7351,N_7593);
nor U8431 (N_8431,N_7984,N_7217);
nor U8432 (N_8432,N_7370,N_7109);
or U8433 (N_8433,N_7068,N_7654);
or U8434 (N_8434,N_7819,N_6851);
nor U8435 (N_8435,N_7468,N_6201);
or U8436 (N_8436,N_7418,N_6529);
and U8437 (N_8437,N_6514,N_6990);
or U8438 (N_8438,N_6007,N_7432);
or U8439 (N_8439,N_6847,N_6401);
nor U8440 (N_8440,N_7061,N_6349);
nand U8441 (N_8441,N_7768,N_7302);
or U8442 (N_8442,N_6458,N_6021);
or U8443 (N_8443,N_6736,N_7609);
or U8444 (N_8444,N_6737,N_6638);
nand U8445 (N_8445,N_7471,N_7584);
nand U8446 (N_8446,N_6143,N_7480);
nand U8447 (N_8447,N_6612,N_7434);
and U8448 (N_8448,N_7391,N_7802);
or U8449 (N_8449,N_6185,N_6482);
nand U8450 (N_8450,N_7184,N_6189);
nand U8451 (N_8451,N_6796,N_6206);
and U8452 (N_8452,N_7931,N_7796);
and U8453 (N_8453,N_7350,N_7629);
or U8454 (N_8454,N_6547,N_6421);
nor U8455 (N_8455,N_6867,N_7741);
xnor U8456 (N_8456,N_7486,N_7460);
or U8457 (N_8457,N_6004,N_6716);
nor U8458 (N_8458,N_6584,N_6409);
nand U8459 (N_8459,N_7945,N_7424);
or U8460 (N_8460,N_7108,N_7203);
and U8461 (N_8461,N_7843,N_7477);
and U8462 (N_8462,N_7526,N_6411);
and U8463 (N_8463,N_6356,N_7343);
or U8464 (N_8464,N_7338,N_6902);
or U8465 (N_8465,N_6567,N_6432);
nand U8466 (N_8466,N_6339,N_6557);
xor U8467 (N_8467,N_6483,N_6035);
nor U8468 (N_8468,N_6367,N_6581);
and U8469 (N_8469,N_7787,N_6284);
nor U8470 (N_8470,N_6578,N_6554);
or U8471 (N_8471,N_7451,N_7224);
xor U8472 (N_8472,N_7845,N_6619);
nand U8473 (N_8473,N_7880,N_7554);
and U8474 (N_8474,N_6941,N_6934);
or U8475 (N_8475,N_6316,N_6230);
nor U8476 (N_8476,N_7784,N_7176);
or U8477 (N_8477,N_6674,N_7154);
nand U8478 (N_8478,N_6527,N_6275);
and U8479 (N_8479,N_7328,N_7749);
nand U8480 (N_8480,N_6917,N_6338);
or U8481 (N_8481,N_6700,N_7071);
nor U8482 (N_8482,N_7498,N_7870);
nor U8483 (N_8483,N_7358,N_7951);
or U8484 (N_8484,N_7681,N_7949);
or U8485 (N_8485,N_6153,N_7438);
and U8486 (N_8486,N_7083,N_6072);
nand U8487 (N_8487,N_7354,N_7279);
nor U8488 (N_8488,N_6806,N_7123);
or U8489 (N_8489,N_7995,N_7105);
or U8490 (N_8490,N_6548,N_7011);
and U8491 (N_8491,N_6635,N_6011);
and U8492 (N_8492,N_7937,N_7098);
and U8493 (N_8493,N_7487,N_6228);
or U8494 (N_8494,N_6966,N_6203);
nor U8495 (N_8495,N_7070,N_7573);
or U8496 (N_8496,N_7277,N_7419);
xor U8497 (N_8497,N_6614,N_7547);
nand U8498 (N_8498,N_6883,N_7665);
or U8499 (N_8499,N_7877,N_7095);
nand U8500 (N_8500,N_7342,N_7956);
or U8501 (N_8501,N_6653,N_6765);
xor U8502 (N_8502,N_7113,N_7871);
and U8503 (N_8503,N_7472,N_6593);
or U8504 (N_8504,N_7950,N_7678);
or U8505 (N_8505,N_7627,N_6168);
or U8506 (N_8506,N_7944,N_7139);
nand U8507 (N_8507,N_6289,N_7099);
nor U8508 (N_8508,N_7269,N_6859);
and U8509 (N_8509,N_7711,N_7535);
xor U8510 (N_8510,N_7053,N_6693);
nor U8511 (N_8511,N_7876,N_7572);
xor U8512 (N_8512,N_7848,N_6231);
and U8513 (N_8513,N_7077,N_6953);
nand U8514 (N_8514,N_7559,N_6341);
or U8515 (N_8515,N_6114,N_6670);
and U8516 (N_8516,N_6278,N_7594);
nor U8517 (N_8517,N_7798,N_6712);
or U8518 (N_8518,N_6335,N_7652);
and U8519 (N_8519,N_6446,N_6550);
nor U8520 (N_8520,N_6361,N_6792);
or U8521 (N_8521,N_6916,N_7769);
nand U8522 (N_8522,N_6330,N_6918);
nor U8523 (N_8523,N_6513,N_7384);
and U8524 (N_8524,N_6113,N_6022);
nand U8525 (N_8525,N_6507,N_7216);
xnor U8526 (N_8526,N_7314,N_7816);
or U8527 (N_8527,N_6936,N_7315);
nor U8528 (N_8528,N_7647,N_6878);
and U8529 (N_8529,N_6111,N_7865);
nand U8530 (N_8530,N_6439,N_7449);
nor U8531 (N_8531,N_6435,N_7409);
or U8532 (N_8532,N_6510,N_7400);
nor U8533 (N_8533,N_7283,N_6009);
or U8534 (N_8534,N_6068,N_6492);
or U8535 (N_8535,N_6459,N_6094);
or U8536 (N_8536,N_6910,N_7398);
nand U8537 (N_8537,N_7948,N_6746);
nand U8538 (N_8538,N_6086,N_6372);
or U8539 (N_8539,N_7646,N_7761);
nor U8540 (N_8540,N_6566,N_6958);
nor U8541 (N_8541,N_7633,N_7655);
nor U8542 (N_8542,N_7320,N_7707);
nand U8543 (N_8543,N_6066,N_7186);
nor U8544 (N_8544,N_7947,N_7484);
nor U8545 (N_8545,N_7890,N_7611);
or U8546 (N_8546,N_6563,N_6549);
xnor U8547 (N_8547,N_7969,N_7042);
nand U8548 (N_8548,N_6156,N_6442);
nor U8549 (N_8549,N_7028,N_7009);
nor U8550 (N_8550,N_6250,N_7126);
and U8551 (N_8551,N_7825,N_6504);
or U8552 (N_8552,N_7855,N_7124);
or U8553 (N_8553,N_6154,N_7412);
nor U8554 (N_8554,N_6065,N_6232);
nor U8555 (N_8555,N_7926,N_6558);
xnor U8556 (N_8556,N_7476,N_6120);
nand U8557 (N_8557,N_7673,N_7849);
nor U8558 (N_8558,N_6271,N_6199);
and U8559 (N_8559,N_6480,N_6815);
or U8560 (N_8560,N_7698,N_7986);
and U8561 (N_8561,N_7661,N_6079);
nor U8562 (N_8562,N_7433,N_7740);
nand U8563 (N_8563,N_7857,N_7638);
nor U8564 (N_8564,N_6633,N_6318);
nor U8565 (N_8565,N_6583,N_7716);
nor U8566 (N_8566,N_7694,N_6538);
nor U8567 (N_8567,N_6761,N_6803);
nor U8568 (N_8568,N_6706,N_7036);
nor U8569 (N_8569,N_6329,N_7321);
nor U8570 (N_8570,N_6501,N_6287);
nand U8571 (N_8571,N_6165,N_6571);
nor U8572 (N_8572,N_7634,N_7130);
nand U8573 (N_8573,N_7929,N_6486);
and U8574 (N_8574,N_6182,N_7091);
xnor U8575 (N_8575,N_6754,N_6551);
nor U8576 (N_8576,N_6363,N_6333);
nor U8577 (N_8577,N_7296,N_6422);
and U8578 (N_8578,N_7729,N_7690);
nor U8579 (N_8579,N_7874,N_7078);
nor U8580 (N_8580,N_6380,N_7470);
and U8581 (N_8581,N_7425,N_6478);
or U8582 (N_8582,N_7187,N_6645);
nand U8583 (N_8583,N_7587,N_7019);
xor U8584 (N_8584,N_6767,N_7505);
and U8585 (N_8585,N_6261,N_7922);
and U8586 (N_8586,N_7166,N_7007);
xor U8587 (N_8587,N_7282,N_7421);
or U8588 (N_8588,N_7256,N_6676);
and U8589 (N_8589,N_7323,N_7988);
or U8590 (N_8590,N_6970,N_7381);
or U8591 (N_8591,N_6166,N_6893);
nor U8592 (N_8592,N_7414,N_7410);
or U8593 (N_8593,N_7565,N_6862);
nand U8594 (N_8594,N_7706,N_7429);
and U8595 (N_8595,N_6644,N_6370);
xor U8596 (N_8596,N_6685,N_6259);
and U8597 (N_8597,N_6092,N_7121);
nor U8598 (N_8598,N_7300,N_7998);
and U8599 (N_8599,N_6833,N_6572);
nor U8600 (N_8600,N_7868,N_6531);
and U8601 (N_8601,N_7417,N_6698);
xor U8602 (N_8602,N_6808,N_6506);
xnor U8603 (N_8603,N_7529,N_7147);
or U8604 (N_8604,N_6745,N_6101);
or U8605 (N_8605,N_6395,N_7010);
and U8606 (N_8606,N_6931,N_7173);
xnor U8607 (N_8607,N_6405,N_6202);
nand U8608 (N_8608,N_7385,N_7510);
nand U8609 (N_8609,N_7879,N_6434);
xor U8610 (N_8610,N_7515,N_7599);
nor U8611 (N_8611,N_7056,N_6610);
and U8612 (N_8612,N_6849,N_6748);
nand U8613 (N_8613,N_6601,N_7311);
or U8614 (N_8614,N_6714,N_6452);
nor U8615 (N_8615,N_7288,N_7374);
and U8616 (N_8616,N_6605,N_7262);
nand U8617 (N_8617,N_7127,N_6236);
nor U8618 (N_8618,N_7667,N_7426);
and U8619 (N_8619,N_6646,N_6173);
xor U8620 (N_8620,N_7110,N_6868);
and U8621 (N_8621,N_7604,N_6760);
and U8622 (N_8622,N_6590,N_7219);
nand U8623 (N_8623,N_7125,N_6874);
nor U8624 (N_8624,N_7474,N_7465);
and U8625 (N_8625,N_7152,N_7102);
and U8626 (N_8626,N_7276,N_7637);
and U8627 (N_8627,N_7676,N_7968);
and U8628 (N_8628,N_6822,N_7536);
and U8629 (N_8629,N_6018,N_6313);
and U8630 (N_8630,N_6383,N_6853);
or U8631 (N_8631,N_6924,N_6533);
nand U8632 (N_8632,N_7043,N_6903);
or U8633 (N_8633,N_7362,N_6087);
or U8634 (N_8634,N_6861,N_6214);
or U8635 (N_8635,N_6901,N_7911);
nor U8636 (N_8636,N_6378,N_7192);
nor U8637 (N_8637,N_7679,N_7352);
or U8638 (N_8638,N_6699,N_6098);
or U8639 (N_8639,N_7141,N_6097);
nor U8640 (N_8640,N_7755,N_7115);
or U8641 (N_8641,N_7428,N_6241);
or U8642 (N_8642,N_6687,N_6408);
nand U8643 (N_8643,N_7431,N_7462);
or U8644 (N_8644,N_6543,N_6771);
nand U8645 (N_8645,N_7504,N_7693);
nand U8646 (N_8646,N_6947,N_6477);
xor U8647 (N_8647,N_6420,N_6596);
nand U8648 (N_8648,N_6331,N_7732);
and U8649 (N_8649,N_6873,N_7257);
or U8650 (N_8650,N_7495,N_7952);
nor U8651 (N_8651,N_7373,N_7582);
nand U8652 (N_8652,N_7917,N_7864);
or U8653 (N_8653,N_6431,N_6167);
nand U8654 (N_8654,N_6648,N_7403);
and U8655 (N_8655,N_7680,N_6809);
nand U8656 (N_8656,N_7853,N_6515);
nand U8657 (N_8657,N_7463,N_7088);
or U8658 (N_8658,N_6300,N_6006);
xnor U8659 (N_8659,N_6376,N_6433);
or U8660 (N_8660,N_6126,N_7447);
nor U8661 (N_8661,N_6056,N_7578);
nand U8662 (N_8662,N_6064,N_6142);
nor U8663 (N_8663,N_7222,N_7509);
nor U8664 (N_8664,N_7140,N_7643);
nor U8665 (N_8665,N_6976,N_7456);
nor U8666 (N_8666,N_6939,N_7622);
or U8667 (N_8667,N_7540,N_7335);
nand U8668 (N_8668,N_7689,N_6651);
or U8669 (N_8669,N_6399,N_6314);
or U8670 (N_8670,N_7085,N_6683);
nor U8671 (N_8671,N_7612,N_6707);
xor U8672 (N_8672,N_7906,N_7731);
nor U8673 (N_8673,N_7522,N_6385);
nor U8674 (N_8674,N_6848,N_7246);
or U8675 (N_8675,N_7620,N_6366);
nor U8676 (N_8676,N_6445,N_7209);
nor U8677 (N_8677,N_7037,N_7118);
nand U8678 (N_8678,N_6334,N_6163);
nor U8679 (N_8679,N_7973,N_7299);
nand U8680 (N_8680,N_7548,N_6175);
nor U8681 (N_8681,N_6752,N_6595);
nor U8682 (N_8682,N_6627,N_7149);
xnor U8683 (N_8683,N_6471,N_6974);
and U8684 (N_8684,N_6198,N_6146);
or U8685 (N_8685,N_6000,N_7621);
or U8686 (N_8686,N_7708,N_7038);
or U8687 (N_8687,N_7093,N_7631);
nor U8688 (N_8688,N_7723,N_7990);
or U8689 (N_8689,N_6955,N_6988);
nand U8690 (N_8690,N_7772,N_7436);
or U8691 (N_8691,N_7653,N_7031);
nor U8692 (N_8692,N_6997,N_6556);
nor U8693 (N_8693,N_6457,N_7132);
and U8694 (N_8694,N_7080,N_7265);
nand U8695 (N_8695,N_7946,N_6475);
nor U8696 (N_8696,N_6810,N_7726);
and U8697 (N_8697,N_6617,N_6274);
or U8698 (N_8698,N_7336,N_6419);
or U8699 (N_8699,N_6387,N_6157);
and U8700 (N_8700,N_7923,N_7727);
xnor U8701 (N_8701,N_7254,N_7997);
nor U8702 (N_8702,N_7107,N_7225);
nand U8703 (N_8703,N_7966,N_7231);
and U8704 (N_8704,N_6836,N_6238);
nand U8705 (N_8705,N_6391,N_6242);
nand U8706 (N_8706,N_6828,N_7270);
or U8707 (N_8707,N_6603,N_7953);
or U8708 (N_8708,N_6542,N_6179);
nor U8709 (N_8709,N_7218,N_7422);
nor U8710 (N_8710,N_7174,N_6070);
nand U8711 (N_8711,N_7924,N_7156);
nor U8712 (N_8712,N_6379,N_7402);
and U8713 (N_8713,N_7982,N_6860);
nor U8714 (N_8714,N_7915,N_6962);
and U8715 (N_8715,N_7363,N_6219);
nand U8716 (N_8716,N_6489,N_6579);
nor U8717 (N_8717,N_6979,N_7489);
or U8718 (N_8718,N_6622,N_6783);
and U8719 (N_8719,N_7985,N_6602);
or U8720 (N_8720,N_6208,N_7326);
or U8721 (N_8721,N_7563,N_6797);
or U8722 (N_8722,N_7213,N_7223);
nor U8723 (N_8723,N_7148,N_7994);
or U8724 (N_8724,N_7736,N_7822);
and U8725 (N_8725,N_6522,N_6240);
or U8726 (N_8726,N_7685,N_6978);
or U8727 (N_8727,N_6059,N_6291);
nor U8728 (N_8728,N_6407,N_7144);
nand U8729 (N_8729,N_6290,N_6981);
or U8730 (N_8730,N_7312,N_7214);
and U8731 (N_8731,N_7756,N_7138);
or U8732 (N_8732,N_6840,N_7479);
and U8733 (N_8733,N_7151,N_7566);
or U8734 (N_8734,N_6528,N_7700);
and U8735 (N_8735,N_7051,N_7271);
or U8736 (N_8736,N_7189,N_7963);
and U8737 (N_8737,N_6105,N_7365);
or U8738 (N_8738,N_7397,N_7448);
nor U8739 (N_8739,N_6360,N_7656);
nor U8740 (N_8740,N_7455,N_6260);
or U8741 (N_8741,N_6975,N_7715);
nor U8742 (N_8742,N_6565,N_6858);
or U8743 (N_8743,N_6865,N_6704);
nor U8744 (N_8744,N_6781,N_6524);
nor U8745 (N_8745,N_6709,N_7789);
and U8746 (N_8746,N_6252,N_7094);
or U8747 (N_8747,N_6037,N_7811);
xnor U8748 (N_8748,N_7258,N_7858);
xnor U8749 (N_8749,N_6772,N_6074);
or U8750 (N_8750,N_6137,N_6160);
and U8751 (N_8751,N_6832,N_7603);
or U8752 (N_8752,N_7894,N_6666);
and U8753 (N_8753,N_7800,N_7247);
and U8754 (N_8754,N_7775,N_7616);
nand U8755 (N_8755,N_7760,N_6659);
and U8756 (N_8756,N_6679,N_7757);
nand U8757 (N_8757,N_6668,N_6701);
xor U8758 (N_8758,N_7395,N_7075);
and U8759 (N_8759,N_6657,N_6518);
nand U8760 (N_8760,N_7996,N_7261);
and U8761 (N_8761,N_6222,N_7976);
nand U8762 (N_8762,N_6112,N_7961);
nor U8763 (N_8763,N_6996,N_6108);
and U8764 (N_8764,N_7717,N_6040);
nor U8765 (N_8765,N_7670,N_7241);
nor U8766 (N_8766,N_6502,N_7940);
nor U8767 (N_8767,N_7273,N_6843);
and U8768 (N_8768,N_6790,N_6762);
or U8769 (N_8769,N_6197,N_7208);
nand U8770 (N_8770,N_6426,N_7589);
xnor U8771 (N_8771,N_6960,N_7202);
and U8772 (N_8772,N_7405,N_6667);
and U8773 (N_8773,N_6448,N_6656);
xor U8774 (N_8774,N_6811,N_7542);
nand U8775 (N_8775,N_6837,N_7782);
and U8776 (N_8776,N_7514,N_7597);
and U8777 (N_8777,N_7494,N_7773);
nand U8778 (N_8778,N_7272,N_7367);
nor U8779 (N_8779,N_6026,N_7194);
nor U8780 (N_8780,N_6233,N_6671);
and U8781 (N_8781,N_7142,N_7528);
nand U8782 (N_8782,N_6908,N_6161);
nor U8783 (N_8783,N_7580,N_6269);
nand U8784 (N_8784,N_6751,N_6984);
or U8785 (N_8785,N_7605,N_7332);
nor U8786 (N_8786,N_6911,N_6205);
or U8787 (N_8787,N_6696,N_6169);
nor U8788 (N_8788,N_6283,N_6826);
or U8789 (N_8789,N_6030,N_7981);
or U8790 (N_8790,N_6733,N_6033);
and U8791 (N_8791,N_7240,N_7556);
nor U8792 (N_8792,N_7226,N_7570);
nand U8793 (N_8793,N_6243,N_6785);
nand U8794 (N_8794,N_6680,N_6017);
and U8795 (N_8795,N_6998,N_7439);
or U8796 (N_8796,N_7281,N_7346);
and U8797 (N_8797,N_7488,N_7493);
and U8798 (N_8798,N_6320,N_6337);
nor U8799 (N_8799,N_6912,N_7702);
xor U8800 (N_8800,N_7878,N_7714);
nand U8801 (N_8801,N_7518,N_7377);
nand U8802 (N_8802,N_7242,N_6642);
xor U8803 (N_8803,N_6398,N_7171);
and U8804 (N_8804,N_7666,N_7167);
nand U8805 (N_8805,N_6258,N_6768);
nor U8806 (N_8806,N_6036,N_7809);
and U8807 (N_8807,N_7170,N_7557);
nor U8808 (N_8808,N_6552,N_7006);
and U8809 (N_8809,N_7143,N_6382);
or U8810 (N_8810,N_7499,N_7780);
nor U8811 (N_8811,N_6418,N_6128);
and U8812 (N_8812,N_7750,N_6319);
or U8813 (N_8813,N_6799,N_6715);
nor U8814 (N_8814,N_6019,N_6103);
or U8815 (N_8815,N_7552,N_6042);
xnor U8816 (N_8816,N_6688,N_6871);
nor U8817 (N_8817,N_7899,N_7831);
nand U8818 (N_8818,N_7244,N_6807);
nor U8819 (N_8819,N_6629,N_7737);
nand U8820 (N_8820,N_6430,N_7753);
or U8821 (N_8821,N_6742,N_7181);
or U8822 (N_8822,N_7232,N_7030);
nor U8823 (N_8823,N_7020,N_6804);
nand U8824 (N_8824,N_7443,N_6749);
nand U8825 (N_8825,N_7763,N_7464);
nor U8826 (N_8826,N_6456,N_6049);
nand U8827 (N_8827,N_6028,N_6545);
nand U8828 (N_8828,N_6200,N_7806);
and U8829 (N_8829,N_7345,N_7064);
nor U8830 (N_8830,N_7193,N_7050);
nand U8831 (N_8831,N_6774,N_7512);
and U8832 (N_8832,N_7478,N_6850);
xnor U8833 (N_8833,N_6977,N_6176);
nand U8834 (N_8834,N_6104,N_6155);
or U8835 (N_8835,N_7533,N_6964);
nor U8836 (N_8836,N_7844,N_7568);
and U8837 (N_8837,N_6526,N_7090);
xnor U8838 (N_8838,N_7210,N_7353);
nand U8839 (N_8839,N_7052,N_7754);
and U8840 (N_8840,N_7182,N_6607);
nor U8841 (N_8841,N_6447,N_7298);
and U8842 (N_8842,N_7266,N_7319);
nor U8843 (N_8843,N_6690,N_6591);
or U8844 (N_8844,N_7025,N_7069);
nor U8845 (N_8845,N_7657,N_6606);
nand U8846 (N_8846,N_6689,N_6141);
nand U8847 (N_8847,N_6989,N_6388);
or U8848 (N_8848,N_6133,N_6308);
nor U8849 (N_8849,N_7833,N_7260);
nand U8850 (N_8850,N_7826,N_7461);
or U8851 (N_8851,N_7600,N_6637);
nand U8852 (N_8852,N_7252,N_7889);
and U8853 (N_8853,N_6345,N_6509);
nand U8854 (N_8854,N_7131,N_7577);
nor U8855 (N_8855,N_7562,N_6900);
or U8856 (N_8856,N_7592,N_7814);
nor U8857 (N_8857,N_6099,N_7396);
nor U8858 (N_8858,N_6880,N_7724);
nor U8859 (N_8859,N_6268,N_6658);
or U8860 (N_8860,N_7883,N_6110);
nand U8861 (N_8861,N_7041,N_7524);
nand U8862 (N_8862,N_6353,N_7324);
xor U8863 (N_8863,N_7204,N_7516);
or U8864 (N_8864,N_7234,N_6403);
or U8865 (N_8865,N_7807,N_6130);
nor U8866 (N_8866,N_7114,N_7380);
xnor U8867 (N_8867,N_6834,N_6304);
and U8868 (N_8868,N_6195,N_7699);
nor U8869 (N_8869,N_6694,N_7987);
or U8870 (N_8870,N_7639,N_7308);
or U8871 (N_8871,N_7450,N_6218);
nand U8872 (N_8872,N_6365,N_6010);
or U8873 (N_8873,N_6819,N_6413);
or U8874 (N_8874,N_7119,N_6215);
and U8875 (N_8875,N_7435,N_6109);
nand U8876 (N_8876,N_6729,N_7357);
or U8877 (N_8877,N_7895,N_6279);
nand U8878 (N_8878,N_7632,N_7096);
nor U8879 (N_8879,N_6164,N_6096);
nand U8880 (N_8880,N_6588,N_7891);
nand U8881 (N_8881,N_6454,N_6211);
and U8882 (N_8882,N_7322,N_7651);
nand U8883 (N_8883,N_7021,N_6392);
nor U8884 (N_8884,N_6251,N_6816);
xor U8885 (N_8885,N_6625,N_6613);
and U8886 (N_8886,N_6965,N_7686);
nor U8887 (N_8887,N_7615,N_6950);
and U8888 (N_8888,N_7783,N_6734);
xnor U8889 (N_8889,N_6497,N_7372);
nor U8890 (N_8890,N_6295,N_6127);
nand U8891 (N_8891,N_7839,N_7619);
or U8892 (N_8892,N_7318,N_6890);
xnor U8893 (N_8893,N_7329,N_7642);
and U8894 (N_8894,N_6660,N_6352);
nor U8895 (N_8895,N_6544,N_6234);
xor U8896 (N_8896,N_6294,N_7630);
xor U8897 (N_8897,N_7120,N_6824);
xnor U8898 (N_8898,N_6838,N_6025);
and U8899 (N_8899,N_6852,N_6044);
and U8900 (N_8900,N_7074,N_7867);
nor U8901 (N_8901,N_6122,N_7507);
nand U8902 (N_8902,N_7097,N_7847);
nor U8903 (N_8903,N_6942,N_7823);
nand U8904 (N_8904,N_6946,N_6404);
or U8905 (N_8905,N_7873,N_7601);
xnor U8906 (N_8906,N_7896,N_7355);
nand U8907 (N_8907,N_6678,N_7062);
or U8908 (N_8908,N_7824,N_6196);
or U8909 (N_8909,N_6343,N_7776);
xnor U8910 (N_8910,N_7854,N_6969);
and U8911 (N_8911,N_6725,N_7907);
nand U8912 (N_8912,N_7129,N_6763);
and U8913 (N_8913,N_6718,N_6789);
nand U8914 (N_8914,N_6954,N_6490);
or U8915 (N_8915,N_7368,N_6083);
nor U8916 (N_8916,N_7683,N_6468);
nor U8917 (N_8917,N_7596,N_7364);
nand U8918 (N_8918,N_6787,N_6692);
nor U8919 (N_8919,N_7446,N_6461);
nor U8920 (N_8920,N_6952,N_6102);
or U8921 (N_8921,N_6058,N_6844);
nor U8922 (N_8922,N_6245,N_7066);
and U8923 (N_8923,N_7862,N_7452);
nand U8924 (N_8924,N_6466,N_6604);
nor U8925 (N_8925,N_7636,N_7190);
nand U8926 (N_8926,N_7781,N_6450);
or U8927 (N_8927,N_6149,N_6024);
xnor U8928 (N_8928,N_6358,N_6428);
and U8929 (N_8929,N_7598,N_6298);
and U8930 (N_8930,N_6521,N_6935);
nand U8931 (N_8931,N_6846,N_6256);
nor U8932 (N_8932,N_7379,N_7004);
nor U8933 (N_8933,N_6905,N_7197);
nand U8934 (N_8934,N_6665,N_6812);
or U8935 (N_8935,N_7567,N_6181);
or U8936 (N_8936,N_7229,N_6740);
or U8937 (N_8937,N_6140,N_6020);
nand U8938 (N_8938,N_7313,N_7490);
and U8939 (N_8939,N_6508,N_6449);
and U8940 (N_8940,N_6123,N_7073);
nor U8941 (N_8941,N_7047,N_7458);
nand U8942 (N_8942,N_7762,N_7645);
nand U8943 (N_8943,N_7586,N_6073);
xor U8944 (N_8944,N_7827,N_7626);
xor U8945 (N_8945,N_7930,N_7371);
nor U8946 (N_8946,N_6820,N_6726);
nor U8947 (N_8947,N_7635,N_6615);
nand U8948 (N_8948,N_6920,N_6559);
nor U8949 (N_8949,N_7017,N_7815);
nor U8950 (N_8950,N_6115,N_7294);
or U8951 (N_8951,N_7544,N_6663);
and U8952 (N_8952,N_6052,N_7280);
and U8953 (N_8953,N_6959,N_6739);
or U8954 (N_8954,N_6437,N_6891);
nor U8955 (N_8955,N_6091,N_7828);
or U8956 (N_8956,N_6587,N_6253);
nor U8957 (N_8957,N_6438,N_6354);
nand U8958 (N_8958,N_7628,N_6986);
nand U8959 (N_8959,N_6029,N_7227);
nor U8960 (N_8960,N_7797,N_7939);
nor U8961 (N_8961,N_7501,N_6015);
nor U8962 (N_8962,N_6302,N_6012);
nand U8963 (N_8963,N_6525,N_6794);
nand U8964 (N_8964,N_7788,N_6731);
xor U8965 (N_8965,N_6956,N_6255);
and U8966 (N_8966,N_6424,N_7914);
nor U8967 (N_8967,N_7860,N_6172);
or U8968 (N_8968,N_7337,N_6938);
or U8969 (N_8969,N_7790,N_6511);
or U8970 (N_8970,N_7692,N_7060);
nor U8971 (N_8971,N_7285,N_6135);
nor U8972 (N_8972,N_6982,N_6050);
nor U8973 (N_8973,N_7550,N_7087);
nand U8974 (N_8974,N_6347,N_7293);
and U8975 (N_8975,N_6488,N_6661);
xor U8976 (N_8976,N_7674,N_6655);
nand U8977 (N_8977,N_7248,N_6186);
nor U8978 (N_8978,N_7117,N_7145);
or U8979 (N_8979,N_6894,N_7553);
or U8980 (N_8980,N_6084,N_7792);
or U8981 (N_8981,N_7534,N_7965);
nor U8982 (N_8982,N_7991,N_7235);
or U8983 (N_8983,N_7420,N_6162);
or U8984 (N_8984,N_6503,N_6472);
and U8985 (N_8985,N_6192,N_7625);
xor U8986 (N_8986,N_6639,N_7979);
and U8987 (N_8987,N_7703,N_6845);
and U8988 (N_8988,N_6747,N_7778);
xor U8989 (N_8989,N_7497,N_7837);
or U8990 (N_8990,N_6375,N_7236);
nand U8991 (N_8991,N_6888,N_7696);
nand U8992 (N_8992,N_7485,N_6577);
or U8993 (N_8993,N_6266,N_6246);
and U8994 (N_8994,N_6738,N_7179);
nand U8995 (N_8995,N_6270,N_7738);
nor U8996 (N_8996,N_6332,N_6623);
nand U8997 (N_8997,N_6226,N_6355);
nor U8998 (N_8998,N_6609,N_6377);
or U8999 (N_8999,N_7892,N_6987);
and U9000 (N_9000,N_7385,N_6413);
nor U9001 (N_9001,N_7881,N_6267);
nand U9002 (N_9002,N_7339,N_6274);
nand U9003 (N_9003,N_6553,N_6633);
and U9004 (N_9004,N_6173,N_6140);
xnor U9005 (N_9005,N_6481,N_7679);
and U9006 (N_9006,N_7350,N_7299);
and U9007 (N_9007,N_6791,N_6182);
nor U9008 (N_9008,N_7033,N_6680);
xnor U9009 (N_9009,N_6863,N_6440);
nand U9010 (N_9010,N_6711,N_6914);
and U9011 (N_9011,N_6789,N_6393);
nand U9012 (N_9012,N_7485,N_6506);
nand U9013 (N_9013,N_6195,N_6096);
nand U9014 (N_9014,N_7327,N_6826);
nand U9015 (N_9015,N_6479,N_7655);
or U9016 (N_9016,N_7222,N_6950);
and U9017 (N_9017,N_6285,N_6814);
or U9018 (N_9018,N_6144,N_6298);
xor U9019 (N_9019,N_7156,N_6155);
or U9020 (N_9020,N_6978,N_6085);
nand U9021 (N_9021,N_6570,N_6601);
nand U9022 (N_9022,N_6657,N_6866);
or U9023 (N_9023,N_7621,N_7543);
xnor U9024 (N_9024,N_7414,N_6287);
nor U9025 (N_9025,N_6750,N_6453);
nand U9026 (N_9026,N_7183,N_7543);
nor U9027 (N_9027,N_6376,N_7019);
nand U9028 (N_9028,N_7464,N_6280);
nand U9029 (N_9029,N_7684,N_6602);
and U9030 (N_9030,N_6641,N_7803);
or U9031 (N_9031,N_7487,N_6787);
nor U9032 (N_9032,N_7945,N_6082);
xor U9033 (N_9033,N_6528,N_7970);
nand U9034 (N_9034,N_7689,N_6669);
or U9035 (N_9035,N_6163,N_7075);
and U9036 (N_9036,N_7872,N_6536);
and U9037 (N_9037,N_7501,N_7609);
xnor U9038 (N_9038,N_6022,N_7310);
nor U9039 (N_9039,N_7218,N_7241);
or U9040 (N_9040,N_6523,N_7169);
or U9041 (N_9041,N_7544,N_7610);
nor U9042 (N_9042,N_6237,N_7045);
nor U9043 (N_9043,N_7211,N_6990);
and U9044 (N_9044,N_7280,N_7140);
nor U9045 (N_9045,N_6914,N_7303);
nor U9046 (N_9046,N_7357,N_6138);
or U9047 (N_9047,N_6213,N_6138);
nor U9048 (N_9048,N_6857,N_7261);
and U9049 (N_9049,N_7857,N_7865);
or U9050 (N_9050,N_7967,N_6565);
xnor U9051 (N_9051,N_7705,N_6740);
nor U9052 (N_9052,N_7358,N_6810);
nand U9053 (N_9053,N_6101,N_7039);
or U9054 (N_9054,N_6534,N_6668);
or U9055 (N_9055,N_7166,N_7987);
nand U9056 (N_9056,N_6092,N_7712);
nand U9057 (N_9057,N_7764,N_7255);
nand U9058 (N_9058,N_6257,N_6749);
nor U9059 (N_9059,N_6546,N_7538);
nand U9060 (N_9060,N_6558,N_7932);
and U9061 (N_9061,N_7390,N_7523);
xor U9062 (N_9062,N_6788,N_6624);
nor U9063 (N_9063,N_7475,N_6434);
or U9064 (N_9064,N_7165,N_6839);
or U9065 (N_9065,N_6550,N_6843);
and U9066 (N_9066,N_6693,N_6232);
or U9067 (N_9067,N_6429,N_7817);
nand U9068 (N_9068,N_6583,N_6468);
and U9069 (N_9069,N_7443,N_6672);
xnor U9070 (N_9070,N_6472,N_7758);
nor U9071 (N_9071,N_6555,N_7533);
or U9072 (N_9072,N_6548,N_7810);
or U9073 (N_9073,N_6345,N_6440);
nand U9074 (N_9074,N_6451,N_7933);
or U9075 (N_9075,N_7203,N_6097);
nor U9076 (N_9076,N_7776,N_7439);
nor U9077 (N_9077,N_7931,N_7756);
nor U9078 (N_9078,N_6595,N_6161);
nand U9079 (N_9079,N_7920,N_6768);
and U9080 (N_9080,N_6816,N_6334);
nor U9081 (N_9081,N_7133,N_6702);
xnor U9082 (N_9082,N_6580,N_7175);
or U9083 (N_9083,N_7775,N_6441);
or U9084 (N_9084,N_6272,N_7617);
and U9085 (N_9085,N_7074,N_7449);
nand U9086 (N_9086,N_6267,N_7716);
nor U9087 (N_9087,N_6390,N_6355);
and U9088 (N_9088,N_6586,N_7690);
nand U9089 (N_9089,N_7282,N_7815);
nor U9090 (N_9090,N_7249,N_7960);
or U9091 (N_9091,N_6327,N_6523);
nand U9092 (N_9092,N_7019,N_6389);
and U9093 (N_9093,N_7590,N_7062);
nor U9094 (N_9094,N_7727,N_7517);
or U9095 (N_9095,N_6225,N_6663);
nor U9096 (N_9096,N_6170,N_6746);
nor U9097 (N_9097,N_6327,N_6866);
nand U9098 (N_9098,N_6681,N_6824);
nand U9099 (N_9099,N_6985,N_6571);
or U9100 (N_9100,N_7859,N_7475);
or U9101 (N_9101,N_6494,N_7507);
or U9102 (N_9102,N_7867,N_6481);
or U9103 (N_9103,N_7861,N_7446);
or U9104 (N_9104,N_6082,N_6035);
and U9105 (N_9105,N_7397,N_7598);
nor U9106 (N_9106,N_6521,N_7702);
nand U9107 (N_9107,N_6424,N_6877);
xor U9108 (N_9108,N_7184,N_7272);
nand U9109 (N_9109,N_7495,N_7927);
or U9110 (N_9110,N_6383,N_6975);
and U9111 (N_9111,N_7009,N_6039);
nand U9112 (N_9112,N_6807,N_7653);
or U9113 (N_9113,N_6006,N_6229);
nand U9114 (N_9114,N_6204,N_7827);
or U9115 (N_9115,N_6839,N_6498);
nor U9116 (N_9116,N_7054,N_6653);
or U9117 (N_9117,N_7410,N_7584);
nor U9118 (N_9118,N_7761,N_7862);
and U9119 (N_9119,N_7873,N_6386);
nor U9120 (N_9120,N_7354,N_7469);
nand U9121 (N_9121,N_7648,N_6362);
or U9122 (N_9122,N_6945,N_6343);
nand U9123 (N_9123,N_7109,N_6562);
nand U9124 (N_9124,N_6426,N_6512);
and U9125 (N_9125,N_7727,N_6949);
and U9126 (N_9126,N_7808,N_7852);
or U9127 (N_9127,N_7666,N_7488);
nor U9128 (N_9128,N_7781,N_6488);
nor U9129 (N_9129,N_7842,N_7017);
xor U9130 (N_9130,N_6983,N_7893);
or U9131 (N_9131,N_7516,N_7889);
nor U9132 (N_9132,N_6555,N_7187);
or U9133 (N_9133,N_6220,N_6329);
and U9134 (N_9134,N_7892,N_6600);
nand U9135 (N_9135,N_7868,N_6064);
and U9136 (N_9136,N_6501,N_6168);
nand U9137 (N_9137,N_7254,N_7293);
nand U9138 (N_9138,N_6604,N_7231);
nand U9139 (N_9139,N_6746,N_6275);
nand U9140 (N_9140,N_7129,N_7925);
nor U9141 (N_9141,N_6369,N_7462);
or U9142 (N_9142,N_7675,N_7360);
nor U9143 (N_9143,N_7573,N_7163);
nand U9144 (N_9144,N_6395,N_7394);
or U9145 (N_9145,N_7617,N_6727);
xor U9146 (N_9146,N_6630,N_7081);
nor U9147 (N_9147,N_7321,N_6312);
and U9148 (N_9148,N_6954,N_7920);
nor U9149 (N_9149,N_7031,N_6911);
xor U9150 (N_9150,N_7870,N_6906);
and U9151 (N_9151,N_7036,N_6068);
nand U9152 (N_9152,N_7479,N_7624);
or U9153 (N_9153,N_6572,N_6950);
or U9154 (N_9154,N_7695,N_6266);
and U9155 (N_9155,N_7281,N_7689);
nand U9156 (N_9156,N_7331,N_6568);
nand U9157 (N_9157,N_7552,N_6945);
nor U9158 (N_9158,N_7102,N_7405);
xnor U9159 (N_9159,N_7033,N_7571);
nor U9160 (N_9160,N_6321,N_6662);
and U9161 (N_9161,N_7688,N_6362);
and U9162 (N_9162,N_7110,N_7918);
nor U9163 (N_9163,N_7289,N_6246);
or U9164 (N_9164,N_7839,N_6586);
and U9165 (N_9165,N_6472,N_7879);
nand U9166 (N_9166,N_7278,N_7527);
nand U9167 (N_9167,N_6493,N_6654);
nor U9168 (N_9168,N_6620,N_6399);
nor U9169 (N_9169,N_7031,N_6929);
and U9170 (N_9170,N_6257,N_6641);
nor U9171 (N_9171,N_6579,N_7022);
and U9172 (N_9172,N_7033,N_7528);
or U9173 (N_9173,N_6059,N_6116);
nor U9174 (N_9174,N_6551,N_7066);
xor U9175 (N_9175,N_6062,N_7941);
nor U9176 (N_9176,N_7637,N_7894);
nand U9177 (N_9177,N_6240,N_7326);
xor U9178 (N_9178,N_6646,N_7540);
nor U9179 (N_9179,N_6961,N_6864);
or U9180 (N_9180,N_7720,N_6626);
nor U9181 (N_9181,N_6257,N_6315);
nand U9182 (N_9182,N_6629,N_6314);
nor U9183 (N_9183,N_6038,N_7654);
or U9184 (N_9184,N_6550,N_7486);
xnor U9185 (N_9185,N_7300,N_7839);
nand U9186 (N_9186,N_6494,N_7780);
nor U9187 (N_9187,N_6941,N_6637);
nand U9188 (N_9188,N_7029,N_6129);
and U9189 (N_9189,N_7838,N_6193);
and U9190 (N_9190,N_7953,N_6691);
and U9191 (N_9191,N_6597,N_7949);
nor U9192 (N_9192,N_7063,N_7363);
nor U9193 (N_9193,N_7565,N_7742);
or U9194 (N_9194,N_6994,N_6540);
nor U9195 (N_9195,N_6366,N_7711);
nand U9196 (N_9196,N_6349,N_6696);
and U9197 (N_9197,N_6429,N_7524);
and U9198 (N_9198,N_7941,N_7076);
or U9199 (N_9199,N_7445,N_6572);
or U9200 (N_9200,N_7105,N_6566);
or U9201 (N_9201,N_7710,N_7670);
nor U9202 (N_9202,N_7281,N_6745);
nand U9203 (N_9203,N_6376,N_7212);
nor U9204 (N_9204,N_7139,N_7546);
or U9205 (N_9205,N_6401,N_6313);
nor U9206 (N_9206,N_7016,N_7953);
or U9207 (N_9207,N_7774,N_7597);
nor U9208 (N_9208,N_7079,N_6685);
nand U9209 (N_9209,N_6891,N_6931);
and U9210 (N_9210,N_7252,N_6435);
or U9211 (N_9211,N_7485,N_7304);
nor U9212 (N_9212,N_7842,N_7532);
xor U9213 (N_9213,N_7668,N_7701);
nor U9214 (N_9214,N_6701,N_7506);
nor U9215 (N_9215,N_7908,N_7648);
and U9216 (N_9216,N_6389,N_6101);
nand U9217 (N_9217,N_6587,N_7987);
nand U9218 (N_9218,N_6475,N_7503);
nand U9219 (N_9219,N_6110,N_6425);
nor U9220 (N_9220,N_7583,N_7622);
and U9221 (N_9221,N_6379,N_7824);
or U9222 (N_9222,N_6078,N_7997);
or U9223 (N_9223,N_7194,N_7113);
xnor U9224 (N_9224,N_6606,N_6705);
nand U9225 (N_9225,N_7343,N_7851);
and U9226 (N_9226,N_7540,N_7735);
and U9227 (N_9227,N_7363,N_7991);
and U9228 (N_9228,N_6264,N_7545);
or U9229 (N_9229,N_7521,N_6529);
or U9230 (N_9230,N_6101,N_6193);
nor U9231 (N_9231,N_6289,N_6517);
and U9232 (N_9232,N_6463,N_6533);
nor U9233 (N_9233,N_6964,N_6724);
and U9234 (N_9234,N_6519,N_6143);
nand U9235 (N_9235,N_7225,N_6084);
nor U9236 (N_9236,N_6788,N_6449);
or U9237 (N_9237,N_7896,N_6266);
and U9238 (N_9238,N_6015,N_6183);
xor U9239 (N_9239,N_7710,N_7276);
nand U9240 (N_9240,N_7498,N_6812);
and U9241 (N_9241,N_6989,N_6709);
and U9242 (N_9242,N_7162,N_7950);
or U9243 (N_9243,N_6698,N_6977);
or U9244 (N_9244,N_7949,N_7633);
nor U9245 (N_9245,N_6688,N_7578);
or U9246 (N_9246,N_6732,N_6904);
or U9247 (N_9247,N_7302,N_7050);
and U9248 (N_9248,N_6589,N_7939);
or U9249 (N_9249,N_7252,N_7124);
and U9250 (N_9250,N_7901,N_7826);
or U9251 (N_9251,N_6850,N_6130);
or U9252 (N_9252,N_6727,N_6281);
nand U9253 (N_9253,N_6856,N_6320);
and U9254 (N_9254,N_6495,N_6241);
xor U9255 (N_9255,N_6361,N_7722);
nor U9256 (N_9256,N_7472,N_7320);
and U9257 (N_9257,N_7285,N_6628);
and U9258 (N_9258,N_7062,N_7074);
xor U9259 (N_9259,N_6990,N_7933);
and U9260 (N_9260,N_6584,N_7439);
or U9261 (N_9261,N_6134,N_7853);
or U9262 (N_9262,N_6025,N_7711);
nor U9263 (N_9263,N_7205,N_7890);
or U9264 (N_9264,N_6805,N_6809);
nand U9265 (N_9265,N_7318,N_7223);
or U9266 (N_9266,N_6486,N_6705);
xor U9267 (N_9267,N_6606,N_6810);
or U9268 (N_9268,N_6003,N_6620);
xor U9269 (N_9269,N_7997,N_6166);
nor U9270 (N_9270,N_6186,N_6479);
xor U9271 (N_9271,N_7988,N_6658);
xor U9272 (N_9272,N_7520,N_7027);
or U9273 (N_9273,N_6379,N_6911);
and U9274 (N_9274,N_7325,N_7540);
xnor U9275 (N_9275,N_7935,N_7971);
nor U9276 (N_9276,N_7955,N_6211);
nand U9277 (N_9277,N_6492,N_6986);
and U9278 (N_9278,N_7009,N_6450);
and U9279 (N_9279,N_7327,N_7133);
and U9280 (N_9280,N_6592,N_7445);
nand U9281 (N_9281,N_6745,N_6947);
nor U9282 (N_9282,N_7927,N_7172);
nand U9283 (N_9283,N_6043,N_7646);
and U9284 (N_9284,N_7130,N_6559);
nor U9285 (N_9285,N_6073,N_7209);
nand U9286 (N_9286,N_7144,N_7994);
and U9287 (N_9287,N_6681,N_6831);
or U9288 (N_9288,N_7452,N_7568);
xor U9289 (N_9289,N_7484,N_7115);
and U9290 (N_9290,N_7310,N_7262);
or U9291 (N_9291,N_6069,N_7081);
xnor U9292 (N_9292,N_7178,N_6524);
nand U9293 (N_9293,N_6779,N_6872);
and U9294 (N_9294,N_7874,N_7310);
or U9295 (N_9295,N_7308,N_7216);
or U9296 (N_9296,N_7671,N_6528);
xor U9297 (N_9297,N_6804,N_7326);
and U9298 (N_9298,N_7535,N_6818);
nor U9299 (N_9299,N_6950,N_6235);
nand U9300 (N_9300,N_6654,N_6244);
nor U9301 (N_9301,N_7890,N_6127);
nor U9302 (N_9302,N_6540,N_6373);
and U9303 (N_9303,N_7772,N_7922);
nor U9304 (N_9304,N_7366,N_7064);
nor U9305 (N_9305,N_7200,N_6399);
and U9306 (N_9306,N_7579,N_6874);
nor U9307 (N_9307,N_6786,N_6767);
and U9308 (N_9308,N_7901,N_7190);
xor U9309 (N_9309,N_7701,N_7383);
or U9310 (N_9310,N_6544,N_6096);
or U9311 (N_9311,N_6412,N_6319);
or U9312 (N_9312,N_6555,N_7461);
nand U9313 (N_9313,N_7598,N_6940);
nand U9314 (N_9314,N_6108,N_7413);
nor U9315 (N_9315,N_7324,N_6109);
nor U9316 (N_9316,N_7420,N_7362);
nor U9317 (N_9317,N_7496,N_6156);
nor U9318 (N_9318,N_7489,N_7755);
nand U9319 (N_9319,N_6818,N_7188);
nand U9320 (N_9320,N_7637,N_6854);
xnor U9321 (N_9321,N_7844,N_7729);
or U9322 (N_9322,N_7740,N_7394);
nor U9323 (N_9323,N_7467,N_6949);
nand U9324 (N_9324,N_6351,N_7041);
and U9325 (N_9325,N_6596,N_6535);
nand U9326 (N_9326,N_6948,N_6142);
and U9327 (N_9327,N_7476,N_7645);
nor U9328 (N_9328,N_7736,N_6873);
and U9329 (N_9329,N_6196,N_6278);
nor U9330 (N_9330,N_6481,N_7105);
and U9331 (N_9331,N_7989,N_6319);
xor U9332 (N_9332,N_7856,N_6656);
or U9333 (N_9333,N_7979,N_6818);
or U9334 (N_9334,N_7612,N_6674);
nand U9335 (N_9335,N_6336,N_7150);
or U9336 (N_9336,N_6988,N_7118);
or U9337 (N_9337,N_6938,N_6324);
xor U9338 (N_9338,N_7175,N_6209);
nand U9339 (N_9339,N_7942,N_7140);
or U9340 (N_9340,N_6012,N_7485);
or U9341 (N_9341,N_6992,N_7836);
or U9342 (N_9342,N_7447,N_7847);
xor U9343 (N_9343,N_6300,N_7705);
or U9344 (N_9344,N_7550,N_6233);
and U9345 (N_9345,N_6873,N_6137);
or U9346 (N_9346,N_7801,N_6350);
and U9347 (N_9347,N_6807,N_6408);
or U9348 (N_9348,N_7459,N_6293);
or U9349 (N_9349,N_7700,N_6816);
xor U9350 (N_9350,N_7582,N_6722);
nand U9351 (N_9351,N_7931,N_6578);
nor U9352 (N_9352,N_7614,N_7111);
nand U9353 (N_9353,N_7975,N_7314);
and U9354 (N_9354,N_6439,N_6854);
xor U9355 (N_9355,N_7302,N_7582);
nand U9356 (N_9356,N_6911,N_7193);
nand U9357 (N_9357,N_6698,N_6644);
nor U9358 (N_9358,N_6106,N_6735);
nand U9359 (N_9359,N_6532,N_6959);
xnor U9360 (N_9360,N_6369,N_6087);
and U9361 (N_9361,N_6562,N_6841);
and U9362 (N_9362,N_7967,N_6975);
and U9363 (N_9363,N_7343,N_7537);
nor U9364 (N_9364,N_6354,N_6072);
or U9365 (N_9365,N_6158,N_7762);
xnor U9366 (N_9366,N_7142,N_7408);
xnor U9367 (N_9367,N_6374,N_7896);
nand U9368 (N_9368,N_7989,N_6018);
nor U9369 (N_9369,N_7701,N_7849);
xnor U9370 (N_9370,N_7949,N_6359);
or U9371 (N_9371,N_6026,N_7828);
or U9372 (N_9372,N_7750,N_7495);
nand U9373 (N_9373,N_7081,N_6297);
nor U9374 (N_9374,N_6428,N_6075);
xor U9375 (N_9375,N_6877,N_6042);
nor U9376 (N_9376,N_7640,N_6550);
nand U9377 (N_9377,N_6412,N_7632);
nor U9378 (N_9378,N_7465,N_7512);
xnor U9379 (N_9379,N_6918,N_7377);
nand U9380 (N_9380,N_6017,N_6317);
and U9381 (N_9381,N_7042,N_7002);
and U9382 (N_9382,N_7840,N_6531);
nand U9383 (N_9383,N_6302,N_6161);
or U9384 (N_9384,N_6128,N_7924);
nor U9385 (N_9385,N_6441,N_7593);
nand U9386 (N_9386,N_6971,N_6870);
nand U9387 (N_9387,N_6659,N_7239);
and U9388 (N_9388,N_6052,N_6922);
and U9389 (N_9389,N_6361,N_6014);
or U9390 (N_9390,N_6583,N_6149);
and U9391 (N_9391,N_6436,N_6940);
nor U9392 (N_9392,N_6140,N_6311);
or U9393 (N_9393,N_7818,N_7397);
or U9394 (N_9394,N_6555,N_7315);
nor U9395 (N_9395,N_7944,N_7420);
nor U9396 (N_9396,N_6783,N_7726);
or U9397 (N_9397,N_6399,N_7320);
and U9398 (N_9398,N_7963,N_6890);
xnor U9399 (N_9399,N_6099,N_6308);
nand U9400 (N_9400,N_7209,N_6771);
or U9401 (N_9401,N_6129,N_6929);
and U9402 (N_9402,N_7980,N_7247);
nor U9403 (N_9403,N_7268,N_7015);
xnor U9404 (N_9404,N_7073,N_6676);
nor U9405 (N_9405,N_6261,N_6901);
nor U9406 (N_9406,N_7522,N_7416);
nand U9407 (N_9407,N_7489,N_6602);
xor U9408 (N_9408,N_6764,N_6044);
nor U9409 (N_9409,N_6204,N_6879);
xnor U9410 (N_9410,N_7160,N_6643);
or U9411 (N_9411,N_7429,N_6664);
nand U9412 (N_9412,N_7615,N_6098);
nand U9413 (N_9413,N_7717,N_7133);
nor U9414 (N_9414,N_7373,N_7633);
nor U9415 (N_9415,N_7306,N_7263);
nor U9416 (N_9416,N_7724,N_7444);
nand U9417 (N_9417,N_6091,N_6671);
or U9418 (N_9418,N_6588,N_6988);
and U9419 (N_9419,N_6636,N_7286);
nand U9420 (N_9420,N_7869,N_6677);
nor U9421 (N_9421,N_6367,N_7214);
xor U9422 (N_9422,N_6429,N_6150);
nor U9423 (N_9423,N_7767,N_7869);
and U9424 (N_9424,N_6041,N_7304);
or U9425 (N_9425,N_7688,N_6122);
or U9426 (N_9426,N_6799,N_6801);
and U9427 (N_9427,N_7201,N_7774);
xnor U9428 (N_9428,N_7835,N_7240);
nand U9429 (N_9429,N_7903,N_7214);
nor U9430 (N_9430,N_7208,N_6381);
nand U9431 (N_9431,N_7360,N_6218);
or U9432 (N_9432,N_7210,N_7542);
or U9433 (N_9433,N_6453,N_7448);
or U9434 (N_9434,N_7117,N_6353);
nand U9435 (N_9435,N_7419,N_7498);
and U9436 (N_9436,N_7700,N_6418);
xor U9437 (N_9437,N_6260,N_6968);
and U9438 (N_9438,N_7432,N_6728);
nand U9439 (N_9439,N_6639,N_6701);
and U9440 (N_9440,N_6064,N_6667);
or U9441 (N_9441,N_6027,N_6492);
nand U9442 (N_9442,N_7179,N_7145);
or U9443 (N_9443,N_6323,N_6077);
xor U9444 (N_9444,N_7526,N_7449);
xor U9445 (N_9445,N_6903,N_7263);
or U9446 (N_9446,N_7220,N_6602);
nor U9447 (N_9447,N_6834,N_6941);
nand U9448 (N_9448,N_6450,N_7649);
and U9449 (N_9449,N_7298,N_6083);
nor U9450 (N_9450,N_6969,N_7244);
nand U9451 (N_9451,N_7170,N_6910);
or U9452 (N_9452,N_7285,N_7833);
and U9453 (N_9453,N_7881,N_7981);
or U9454 (N_9454,N_6158,N_6871);
nor U9455 (N_9455,N_7164,N_7143);
or U9456 (N_9456,N_6798,N_6341);
or U9457 (N_9457,N_7652,N_7851);
nand U9458 (N_9458,N_6666,N_7601);
nor U9459 (N_9459,N_6101,N_7892);
nor U9460 (N_9460,N_6528,N_6465);
or U9461 (N_9461,N_7553,N_7279);
nand U9462 (N_9462,N_7918,N_6797);
or U9463 (N_9463,N_6207,N_6974);
nand U9464 (N_9464,N_6032,N_7604);
nor U9465 (N_9465,N_7936,N_6756);
or U9466 (N_9466,N_7363,N_7913);
nor U9467 (N_9467,N_7984,N_6391);
nor U9468 (N_9468,N_6607,N_7984);
and U9469 (N_9469,N_7675,N_6345);
nor U9470 (N_9470,N_7878,N_6171);
or U9471 (N_9471,N_7014,N_6460);
or U9472 (N_9472,N_6128,N_6139);
and U9473 (N_9473,N_7847,N_6888);
or U9474 (N_9474,N_7949,N_7147);
or U9475 (N_9475,N_7681,N_7288);
nand U9476 (N_9476,N_7400,N_7522);
and U9477 (N_9477,N_7485,N_7927);
or U9478 (N_9478,N_6469,N_6294);
xnor U9479 (N_9479,N_7004,N_6388);
or U9480 (N_9480,N_7413,N_6844);
nand U9481 (N_9481,N_6713,N_6767);
and U9482 (N_9482,N_6226,N_6252);
or U9483 (N_9483,N_6815,N_7723);
and U9484 (N_9484,N_6685,N_6828);
nor U9485 (N_9485,N_7206,N_6188);
and U9486 (N_9486,N_6915,N_7604);
or U9487 (N_9487,N_7356,N_7816);
nand U9488 (N_9488,N_6113,N_6983);
nand U9489 (N_9489,N_7850,N_7111);
nor U9490 (N_9490,N_7085,N_6959);
nand U9491 (N_9491,N_6009,N_6773);
nand U9492 (N_9492,N_6365,N_7669);
nor U9493 (N_9493,N_6599,N_7522);
nand U9494 (N_9494,N_6003,N_7378);
and U9495 (N_9495,N_6626,N_7125);
or U9496 (N_9496,N_7764,N_7441);
or U9497 (N_9497,N_7099,N_7990);
nand U9498 (N_9498,N_6520,N_7809);
nor U9499 (N_9499,N_7306,N_7232);
nor U9500 (N_9500,N_6911,N_7372);
or U9501 (N_9501,N_6704,N_7937);
nand U9502 (N_9502,N_6129,N_7018);
and U9503 (N_9503,N_7595,N_6391);
and U9504 (N_9504,N_7177,N_7636);
or U9505 (N_9505,N_6615,N_6322);
and U9506 (N_9506,N_7757,N_7267);
nand U9507 (N_9507,N_7454,N_6395);
or U9508 (N_9508,N_6823,N_6901);
xnor U9509 (N_9509,N_7267,N_7627);
xnor U9510 (N_9510,N_6338,N_6392);
nand U9511 (N_9511,N_7923,N_7777);
nor U9512 (N_9512,N_7482,N_6171);
nand U9513 (N_9513,N_7550,N_7897);
or U9514 (N_9514,N_7288,N_7870);
nand U9515 (N_9515,N_7874,N_6491);
or U9516 (N_9516,N_6143,N_6121);
nor U9517 (N_9517,N_6511,N_6090);
and U9518 (N_9518,N_7670,N_6427);
xor U9519 (N_9519,N_6800,N_6235);
and U9520 (N_9520,N_6419,N_6028);
xnor U9521 (N_9521,N_6061,N_6677);
nor U9522 (N_9522,N_6959,N_6396);
and U9523 (N_9523,N_7118,N_7823);
or U9524 (N_9524,N_6440,N_7135);
or U9525 (N_9525,N_7586,N_7430);
xor U9526 (N_9526,N_7799,N_7487);
nand U9527 (N_9527,N_7780,N_7491);
or U9528 (N_9528,N_6874,N_6841);
nand U9529 (N_9529,N_6157,N_6302);
or U9530 (N_9530,N_6739,N_7263);
and U9531 (N_9531,N_6157,N_7244);
xnor U9532 (N_9532,N_7797,N_7966);
nor U9533 (N_9533,N_7140,N_6896);
and U9534 (N_9534,N_6685,N_6764);
nor U9535 (N_9535,N_6773,N_7791);
nand U9536 (N_9536,N_7286,N_7886);
or U9537 (N_9537,N_7779,N_7458);
nor U9538 (N_9538,N_7249,N_6369);
or U9539 (N_9539,N_6893,N_7579);
nor U9540 (N_9540,N_6685,N_6128);
nand U9541 (N_9541,N_7382,N_6366);
nor U9542 (N_9542,N_7639,N_7853);
or U9543 (N_9543,N_6155,N_7615);
and U9544 (N_9544,N_6394,N_7161);
nor U9545 (N_9545,N_7485,N_7343);
and U9546 (N_9546,N_7594,N_7216);
nand U9547 (N_9547,N_6100,N_6361);
nand U9548 (N_9548,N_6557,N_7987);
nand U9549 (N_9549,N_7894,N_7634);
or U9550 (N_9550,N_7450,N_6824);
xnor U9551 (N_9551,N_6250,N_7713);
or U9552 (N_9552,N_6211,N_7656);
and U9553 (N_9553,N_7356,N_6172);
nand U9554 (N_9554,N_7225,N_7481);
or U9555 (N_9555,N_7022,N_7592);
or U9556 (N_9556,N_6804,N_7732);
or U9557 (N_9557,N_7002,N_7122);
nand U9558 (N_9558,N_6284,N_7999);
nand U9559 (N_9559,N_7663,N_7088);
or U9560 (N_9560,N_6760,N_7711);
nor U9561 (N_9561,N_7393,N_6862);
or U9562 (N_9562,N_7102,N_6923);
nor U9563 (N_9563,N_6241,N_6497);
and U9564 (N_9564,N_7115,N_7843);
or U9565 (N_9565,N_7162,N_6469);
and U9566 (N_9566,N_6759,N_7200);
or U9567 (N_9567,N_6325,N_7271);
nand U9568 (N_9568,N_7052,N_7765);
and U9569 (N_9569,N_6881,N_6342);
or U9570 (N_9570,N_7938,N_7181);
or U9571 (N_9571,N_6381,N_6678);
nor U9572 (N_9572,N_6562,N_6713);
or U9573 (N_9573,N_7044,N_6741);
nand U9574 (N_9574,N_6498,N_6559);
and U9575 (N_9575,N_7065,N_6883);
nand U9576 (N_9576,N_7371,N_7585);
xnor U9577 (N_9577,N_7511,N_6985);
xnor U9578 (N_9578,N_7564,N_7096);
xnor U9579 (N_9579,N_6809,N_6167);
nor U9580 (N_9580,N_7736,N_6806);
or U9581 (N_9581,N_6748,N_7123);
or U9582 (N_9582,N_7251,N_6427);
and U9583 (N_9583,N_6518,N_7160);
and U9584 (N_9584,N_7138,N_7083);
and U9585 (N_9585,N_7782,N_6960);
and U9586 (N_9586,N_6213,N_7683);
nor U9587 (N_9587,N_6044,N_7487);
or U9588 (N_9588,N_6222,N_6762);
xnor U9589 (N_9589,N_6630,N_7005);
and U9590 (N_9590,N_6959,N_7132);
and U9591 (N_9591,N_6077,N_6752);
or U9592 (N_9592,N_7115,N_7956);
nor U9593 (N_9593,N_7128,N_6932);
nor U9594 (N_9594,N_6568,N_6877);
or U9595 (N_9595,N_6578,N_6869);
and U9596 (N_9596,N_6154,N_7386);
nand U9597 (N_9597,N_7620,N_7125);
xnor U9598 (N_9598,N_7785,N_7244);
xnor U9599 (N_9599,N_7565,N_6143);
nor U9600 (N_9600,N_7737,N_6489);
xnor U9601 (N_9601,N_6127,N_7575);
nor U9602 (N_9602,N_6197,N_7049);
nor U9603 (N_9603,N_6613,N_7197);
nor U9604 (N_9604,N_7298,N_6480);
nand U9605 (N_9605,N_6219,N_7508);
and U9606 (N_9606,N_7467,N_6833);
or U9607 (N_9607,N_6514,N_7956);
nand U9608 (N_9608,N_6860,N_6335);
nand U9609 (N_9609,N_6989,N_7165);
nor U9610 (N_9610,N_7846,N_7747);
nand U9611 (N_9611,N_6153,N_6799);
and U9612 (N_9612,N_6085,N_6862);
xor U9613 (N_9613,N_7415,N_6392);
and U9614 (N_9614,N_6536,N_7042);
xor U9615 (N_9615,N_7741,N_6792);
or U9616 (N_9616,N_6968,N_6181);
xnor U9617 (N_9617,N_6733,N_6803);
or U9618 (N_9618,N_6383,N_7508);
nand U9619 (N_9619,N_7456,N_7617);
nor U9620 (N_9620,N_6185,N_7766);
and U9621 (N_9621,N_7363,N_6815);
nand U9622 (N_9622,N_7875,N_7111);
and U9623 (N_9623,N_7296,N_7865);
or U9624 (N_9624,N_6613,N_7773);
and U9625 (N_9625,N_6879,N_6794);
nor U9626 (N_9626,N_7557,N_6974);
nor U9627 (N_9627,N_7071,N_7072);
xnor U9628 (N_9628,N_7700,N_6880);
nand U9629 (N_9629,N_7952,N_7692);
nor U9630 (N_9630,N_7632,N_7185);
and U9631 (N_9631,N_7714,N_6573);
and U9632 (N_9632,N_7560,N_7689);
and U9633 (N_9633,N_7525,N_6270);
xnor U9634 (N_9634,N_7775,N_7221);
nand U9635 (N_9635,N_6459,N_7276);
and U9636 (N_9636,N_7609,N_7894);
and U9637 (N_9637,N_7388,N_7520);
and U9638 (N_9638,N_7795,N_6481);
nor U9639 (N_9639,N_6899,N_7376);
and U9640 (N_9640,N_7016,N_6508);
and U9641 (N_9641,N_6105,N_6693);
or U9642 (N_9642,N_7357,N_7526);
and U9643 (N_9643,N_7103,N_6275);
xor U9644 (N_9644,N_7971,N_6872);
nor U9645 (N_9645,N_6134,N_6888);
nor U9646 (N_9646,N_6689,N_6220);
and U9647 (N_9647,N_6370,N_6203);
xor U9648 (N_9648,N_7590,N_7461);
nand U9649 (N_9649,N_6790,N_7462);
xnor U9650 (N_9650,N_6037,N_7131);
or U9651 (N_9651,N_7617,N_7335);
nor U9652 (N_9652,N_6207,N_7173);
xnor U9653 (N_9653,N_6559,N_7361);
nand U9654 (N_9654,N_7521,N_6712);
xnor U9655 (N_9655,N_7978,N_7471);
nor U9656 (N_9656,N_7687,N_6502);
nand U9657 (N_9657,N_6122,N_7767);
and U9658 (N_9658,N_7135,N_7378);
nand U9659 (N_9659,N_7085,N_7256);
xor U9660 (N_9660,N_6779,N_6564);
or U9661 (N_9661,N_7958,N_6803);
and U9662 (N_9662,N_6685,N_6881);
or U9663 (N_9663,N_6198,N_6994);
nor U9664 (N_9664,N_6903,N_6541);
xor U9665 (N_9665,N_7938,N_7821);
or U9666 (N_9666,N_6115,N_7010);
nand U9667 (N_9667,N_7911,N_7700);
or U9668 (N_9668,N_6960,N_7106);
or U9669 (N_9669,N_6512,N_6511);
or U9670 (N_9670,N_7020,N_6662);
and U9671 (N_9671,N_6377,N_6653);
and U9672 (N_9672,N_7779,N_7531);
and U9673 (N_9673,N_6919,N_7024);
and U9674 (N_9674,N_7537,N_6773);
and U9675 (N_9675,N_7647,N_6229);
nand U9676 (N_9676,N_7164,N_6168);
or U9677 (N_9677,N_6879,N_7870);
or U9678 (N_9678,N_7031,N_7648);
and U9679 (N_9679,N_7768,N_7003);
and U9680 (N_9680,N_7764,N_6567);
or U9681 (N_9681,N_7345,N_6257);
and U9682 (N_9682,N_7065,N_6811);
nand U9683 (N_9683,N_7772,N_6211);
nand U9684 (N_9684,N_6001,N_6899);
nand U9685 (N_9685,N_6613,N_7866);
nand U9686 (N_9686,N_7964,N_7377);
xor U9687 (N_9687,N_7684,N_6413);
or U9688 (N_9688,N_6646,N_7469);
or U9689 (N_9689,N_6935,N_7215);
or U9690 (N_9690,N_7256,N_6077);
nor U9691 (N_9691,N_7313,N_6161);
and U9692 (N_9692,N_7771,N_7661);
and U9693 (N_9693,N_6199,N_6975);
or U9694 (N_9694,N_7232,N_6770);
nand U9695 (N_9695,N_7819,N_6465);
nor U9696 (N_9696,N_7026,N_6430);
or U9697 (N_9697,N_7309,N_6239);
and U9698 (N_9698,N_7734,N_6239);
nor U9699 (N_9699,N_6452,N_7485);
nor U9700 (N_9700,N_7905,N_7820);
nor U9701 (N_9701,N_6340,N_6814);
and U9702 (N_9702,N_6925,N_7599);
xnor U9703 (N_9703,N_7376,N_7714);
nand U9704 (N_9704,N_6653,N_7723);
and U9705 (N_9705,N_7704,N_7851);
and U9706 (N_9706,N_6276,N_6763);
and U9707 (N_9707,N_6347,N_6399);
nand U9708 (N_9708,N_6124,N_6944);
nand U9709 (N_9709,N_7274,N_6255);
or U9710 (N_9710,N_7107,N_7031);
and U9711 (N_9711,N_7291,N_6367);
nand U9712 (N_9712,N_7157,N_6662);
nand U9713 (N_9713,N_7133,N_7407);
nor U9714 (N_9714,N_6704,N_6259);
nand U9715 (N_9715,N_6995,N_7870);
nor U9716 (N_9716,N_6071,N_7593);
and U9717 (N_9717,N_7921,N_6225);
xnor U9718 (N_9718,N_7078,N_7323);
nand U9719 (N_9719,N_7702,N_7505);
nor U9720 (N_9720,N_7970,N_6133);
nand U9721 (N_9721,N_6205,N_7440);
nand U9722 (N_9722,N_6835,N_7268);
nand U9723 (N_9723,N_6062,N_6162);
and U9724 (N_9724,N_7680,N_7546);
nor U9725 (N_9725,N_7517,N_6644);
nand U9726 (N_9726,N_6932,N_6625);
nand U9727 (N_9727,N_6958,N_6009);
and U9728 (N_9728,N_7606,N_6606);
or U9729 (N_9729,N_6563,N_7206);
or U9730 (N_9730,N_6304,N_6992);
or U9731 (N_9731,N_6827,N_6840);
or U9732 (N_9732,N_7034,N_6416);
nor U9733 (N_9733,N_7726,N_6950);
nor U9734 (N_9734,N_7728,N_7718);
and U9735 (N_9735,N_6072,N_6405);
or U9736 (N_9736,N_7421,N_6576);
and U9737 (N_9737,N_6876,N_7016);
nor U9738 (N_9738,N_6152,N_7876);
and U9739 (N_9739,N_7996,N_7084);
nand U9740 (N_9740,N_7433,N_7905);
or U9741 (N_9741,N_6137,N_7251);
or U9742 (N_9742,N_7710,N_6798);
nor U9743 (N_9743,N_6103,N_6312);
or U9744 (N_9744,N_7497,N_6117);
and U9745 (N_9745,N_7086,N_6045);
or U9746 (N_9746,N_7577,N_6676);
and U9747 (N_9747,N_7287,N_6190);
nor U9748 (N_9748,N_7621,N_7506);
and U9749 (N_9749,N_6819,N_7852);
and U9750 (N_9750,N_7773,N_7632);
or U9751 (N_9751,N_6610,N_6818);
nand U9752 (N_9752,N_6773,N_7007);
nor U9753 (N_9753,N_6862,N_6586);
xor U9754 (N_9754,N_6609,N_7172);
nand U9755 (N_9755,N_6272,N_7273);
nor U9756 (N_9756,N_7814,N_6091);
and U9757 (N_9757,N_6551,N_7643);
xor U9758 (N_9758,N_7992,N_6393);
or U9759 (N_9759,N_7120,N_6035);
nand U9760 (N_9760,N_7249,N_6992);
and U9761 (N_9761,N_7531,N_7663);
nor U9762 (N_9762,N_7914,N_7309);
xor U9763 (N_9763,N_6020,N_6841);
or U9764 (N_9764,N_7718,N_6735);
nand U9765 (N_9765,N_6526,N_6457);
or U9766 (N_9766,N_6833,N_7244);
nor U9767 (N_9767,N_7110,N_7243);
and U9768 (N_9768,N_6824,N_6343);
and U9769 (N_9769,N_6989,N_7877);
xor U9770 (N_9770,N_7108,N_7240);
or U9771 (N_9771,N_6843,N_6786);
xnor U9772 (N_9772,N_7845,N_6949);
nor U9773 (N_9773,N_7038,N_7087);
and U9774 (N_9774,N_7263,N_6669);
or U9775 (N_9775,N_6885,N_6279);
or U9776 (N_9776,N_6260,N_6072);
and U9777 (N_9777,N_6940,N_7165);
xor U9778 (N_9778,N_6060,N_7629);
or U9779 (N_9779,N_6836,N_6212);
nand U9780 (N_9780,N_7306,N_6991);
or U9781 (N_9781,N_7479,N_6499);
nor U9782 (N_9782,N_7932,N_7907);
nand U9783 (N_9783,N_6686,N_7818);
nand U9784 (N_9784,N_7709,N_6934);
nor U9785 (N_9785,N_7646,N_7297);
or U9786 (N_9786,N_6971,N_6495);
xnor U9787 (N_9787,N_6965,N_6165);
nor U9788 (N_9788,N_7115,N_6636);
xor U9789 (N_9789,N_7258,N_7393);
nor U9790 (N_9790,N_7001,N_7141);
or U9791 (N_9791,N_7565,N_6582);
nor U9792 (N_9792,N_7110,N_7009);
and U9793 (N_9793,N_6276,N_6563);
xnor U9794 (N_9794,N_6604,N_6732);
or U9795 (N_9795,N_6332,N_6203);
and U9796 (N_9796,N_7489,N_7483);
or U9797 (N_9797,N_6272,N_7192);
or U9798 (N_9798,N_7284,N_7455);
or U9799 (N_9799,N_7579,N_7066);
and U9800 (N_9800,N_7721,N_7099);
nand U9801 (N_9801,N_7328,N_6895);
nand U9802 (N_9802,N_6852,N_7884);
nand U9803 (N_9803,N_7619,N_6236);
nand U9804 (N_9804,N_6734,N_7574);
and U9805 (N_9805,N_7685,N_7928);
nor U9806 (N_9806,N_7247,N_7553);
xnor U9807 (N_9807,N_7070,N_6978);
and U9808 (N_9808,N_7449,N_6630);
nand U9809 (N_9809,N_6847,N_7985);
nand U9810 (N_9810,N_7931,N_7177);
and U9811 (N_9811,N_7348,N_6185);
nand U9812 (N_9812,N_6280,N_6095);
xnor U9813 (N_9813,N_7760,N_7904);
and U9814 (N_9814,N_7338,N_7457);
or U9815 (N_9815,N_7681,N_6550);
xnor U9816 (N_9816,N_6220,N_6945);
or U9817 (N_9817,N_7621,N_7018);
or U9818 (N_9818,N_7028,N_7543);
xnor U9819 (N_9819,N_7169,N_7075);
nand U9820 (N_9820,N_6404,N_6874);
nand U9821 (N_9821,N_6568,N_6192);
or U9822 (N_9822,N_6440,N_6807);
or U9823 (N_9823,N_6506,N_7158);
xor U9824 (N_9824,N_7453,N_6111);
and U9825 (N_9825,N_7347,N_6611);
xor U9826 (N_9826,N_7686,N_6455);
or U9827 (N_9827,N_6322,N_6965);
nand U9828 (N_9828,N_6900,N_6668);
nor U9829 (N_9829,N_7676,N_6144);
nor U9830 (N_9830,N_7893,N_6539);
nor U9831 (N_9831,N_6678,N_6357);
nor U9832 (N_9832,N_6072,N_6527);
nand U9833 (N_9833,N_7683,N_7524);
and U9834 (N_9834,N_7784,N_6414);
or U9835 (N_9835,N_6561,N_7686);
nor U9836 (N_9836,N_7733,N_6640);
nor U9837 (N_9837,N_7176,N_6536);
nor U9838 (N_9838,N_6089,N_6705);
or U9839 (N_9839,N_7108,N_6970);
xor U9840 (N_9840,N_6798,N_6326);
nor U9841 (N_9841,N_7957,N_6625);
and U9842 (N_9842,N_6622,N_7638);
nand U9843 (N_9843,N_7352,N_7458);
nor U9844 (N_9844,N_7959,N_6592);
or U9845 (N_9845,N_7601,N_7573);
nand U9846 (N_9846,N_6755,N_7925);
or U9847 (N_9847,N_6449,N_6945);
nand U9848 (N_9848,N_6572,N_7524);
nor U9849 (N_9849,N_6098,N_7511);
or U9850 (N_9850,N_7278,N_6504);
nand U9851 (N_9851,N_6879,N_6706);
and U9852 (N_9852,N_7905,N_6033);
and U9853 (N_9853,N_7569,N_7676);
or U9854 (N_9854,N_6329,N_6125);
nand U9855 (N_9855,N_6699,N_7145);
nand U9856 (N_9856,N_6222,N_7012);
nor U9857 (N_9857,N_7126,N_7477);
nand U9858 (N_9858,N_7696,N_6337);
and U9859 (N_9859,N_7128,N_6262);
xnor U9860 (N_9860,N_6959,N_7638);
nor U9861 (N_9861,N_7589,N_6388);
or U9862 (N_9862,N_6361,N_7610);
or U9863 (N_9863,N_7553,N_6368);
nand U9864 (N_9864,N_6056,N_6531);
nand U9865 (N_9865,N_6070,N_7114);
and U9866 (N_9866,N_7141,N_7789);
and U9867 (N_9867,N_6838,N_6504);
nand U9868 (N_9868,N_7890,N_7916);
or U9869 (N_9869,N_7501,N_7235);
and U9870 (N_9870,N_7182,N_7125);
nor U9871 (N_9871,N_7350,N_7018);
nand U9872 (N_9872,N_6275,N_6668);
nand U9873 (N_9873,N_6832,N_7811);
nor U9874 (N_9874,N_6378,N_7683);
xnor U9875 (N_9875,N_7033,N_6546);
and U9876 (N_9876,N_7880,N_7939);
nor U9877 (N_9877,N_6077,N_6440);
nor U9878 (N_9878,N_6945,N_6995);
and U9879 (N_9879,N_6402,N_7829);
or U9880 (N_9880,N_7360,N_6382);
nor U9881 (N_9881,N_6500,N_6344);
nand U9882 (N_9882,N_6870,N_6758);
nand U9883 (N_9883,N_6107,N_7204);
and U9884 (N_9884,N_6314,N_7735);
and U9885 (N_9885,N_7116,N_7173);
and U9886 (N_9886,N_7462,N_6422);
or U9887 (N_9887,N_6415,N_6921);
nand U9888 (N_9888,N_6637,N_7356);
nor U9889 (N_9889,N_7143,N_6203);
xnor U9890 (N_9890,N_7402,N_7430);
or U9891 (N_9891,N_6047,N_7009);
nand U9892 (N_9892,N_6694,N_7985);
nor U9893 (N_9893,N_6709,N_6360);
and U9894 (N_9894,N_7198,N_6994);
nand U9895 (N_9895,N_6847,N_7359);
nor U9896 (N_9896,N_6345,N_7749);
nor U9897 (N_9897,N_6722,N_7590);
xor U9898 (N_9898,N_6750,N_7387);
nor U9899 (N_9899,N_6224,N_7665);
nor U9900 (N_9900,N_6681,N_6980);
and U9901 (N_9901,N_7519,N_6333);
or U9902 (N_9902,N_6489,N_6388);
or U9903 (N_9903,N_6503,N_7010);
and U9904 (N_9904,N_6089,N_7408);
nor U9905 (N_9905,N_7077,N_7046);
nor U9906 (N_9906,N_7400,N_7625);
nand U9907 (N_9907,N_6187,N_6342);
and U9908 (N_9908,N_6656,N_6038);
and U9909 (N_9909,N_7632,N_7998);
nor U9910 (N_9910,N_7329,N_6490);
nand U9911 (N_9911,N_7150,N_7167);
nand U9912 (N_9912,N_6255,N_6365);
nand U9913 (N_9913,N_6370,N_6067);
and U9914 (N_9914,N_7834,N_6636);
nand U9915 (N_9915,N_6663,N_7735);
and U9916 (N_9916,N_6534,N_7366);
xor U9917 (N_9917,N_6173,N_6949);
or U9918 (N_9918,N_6832,N_6489);
or U9919 (N_9919,N_6886,N_6189);
and U9920 (N_9920,N_6016,N_6013);
or U9921 (N_9921,N_6610,N_6731);
nor U9922 (N_9922,N_7452,N_6757);
nor U9923 (N_9923,N_7335,N_6509);
or U9924 (N_9924,N_7901,N_6427);
nor U9925 (N_9925,N_6424,N_7591);
nand U9926 (N_9926,N_6812,N_6748);
xor U9927 (N_9927,N_7781,N_6145);
and U9928 (N_9928,N_7186,N_7709);
or U9929 (N_9929,N_7167,N_7271);
or U9930 (N_9930,N_6341,N_7598);
xnor U9931 (N_9931,N_6837,N_7597);
nor U9932 (N_9932,N_7725,N_7477);
and U9933 (N_9933,N_7969,N_6103);
and U9934 (N_9934,N_6027,N_6094);
xor U9935 (N_9935,N_6693,N_7918);
and U9936 (N_9936,N_7822,N_7776);
xnor U9937 (N_9937,N_7513,N_7063);
xor U9938 (N_9938,N_7868,N_7997);
nand U9939 (N_9939,N_6501,N_6992);
and U9940 (N_9940,N_6968,N_7372);
or U9941 (N_9941,N_7029,N_7709);
nand U9942 (N_9942,N_7635,N_7382);
and U9943 (N_9943,N_7317,N_7973);
and U9944 (N_9944,N_7519,N_6179);
or U9945 (N_9945,N_6651,N_6156);
and U9946 (N_9946,N_6308,N_7324);
xnor U9947 (N_9947,N_7991,N_7498);
nor U9948 (N_9948,N_7106,N_6618);
or U9949 (N_9949,N_7950,N_7323);
and U9950 (N_9950,N_7007,N_7823);
and U9951 (N_9951,N_7157,N_7277);
nor U9952 (N_9952,N_6593,N_7013);
xor U9953 (N_9953,N_6223,N_7068);
xnor U9954 (N_9954,N_7005,N_7473);
xnor U9955 (N_9955,N_7455,N_7858);
nor U9956 (N_9956,N_6006,N_7678);
and U9957 (N_9957,N_6267,N_6979);
nand U9958 (N_9958,N_7912,N_7063);
or U9959 (N_9959,N_6982,N_6534);
nor U9960 (N_9960,N_7486,N_7034);
nand U9961 (N_9961,N_7212,N_7050);
nor U9962 (N_9962,N_6452,N_6998);
or U9963 (N_9963,N_6157,N_7631);
nor U9964 (N_9964,N_7593,N_6135);
or U9965 (N_9965,N_6162,N_7794);
and U9966 (N_9966,N_7147,N_7209);
nand U9967 (N_9967,N_7021,N_6947);
xor U9968 (N_9968,N_7670,N_7539);
nand U9969 (N_9969,N_6792,N_7712);
or U9970 (N_9970,N_7054,N_7932);
nand U9971 (N_9971,N_7043,N_7966);
nand U9972 (N_9972,N_6576,N_6090);
xnor U9973 (N_9973,N_6840,N_6804);
xor U9974 (N_9974,N_7159,N_7266);
nor U9975 (N_9975,N_7920,N_6733);
xnor U9976 (N_9976,N_7932,N_7350);
or U9977 (N_9977,N_6088,N_6913);
or U9978 (N_9978,N_7475,N_7910);
nand U9979 (N_9979,N_7440,N_7961);
or U9980 (N_9980,N_7865,N_7424);
nand U9981 (N_9981,N_7893,N_7583);
nor U9982 (N_9982,N_7274,N_6513);
and U9983 (N_9983,N_7763,N_6177);
and U9984 (N_9984,N_6706,N_6049);
nand U9985 (N_9985,N_7005,N_6070);
nand U9986 (N_9986,N_7292,N_6922);
nand U9987 (N_9987,N_7835,N_6164);
xnor U9988 (N_9988,N_6748,N_6325);
and U9989 (N_9989,N_7136,N_7833);
and U9990 (N_9990,N_6981,N_6484);
or U9991 (N_9991,N_7113,N_6879);
and U9992 (N_9992,N_6638,N_6978);
nor U9993 (N_9993,N_7978,N_7532);
and U9994 (N_9994,N_6266,N_6789);
or U9995 (N_9995,N_7343,N_7476);
nand U9996 (N_9996,N_7356,N_7657);
xor U9997 (N_9997,N_6309,N_7648);
or U9998 (N_9998,N_6128,N_7061);
nand U9999 (N_9999,N_6789,N_7911);
nor UO_0 (O_0,N_8965,N_9832);
and UO_1 (O_1,N_8746,N_9258);
and UO_2 (O_2,N_9046,N_8667);
or UO_3 (O_3,N_9466,N_9527);
nor UO_4 (O_4,N_9242,N_9789);
nor UO_5 (O_5,N_9146,N_9432);
and UO_6 (O_6,N_9438,N_9373);
or UO_7 (O_7,N_8753,N_9967);
and UO_8 (O_8,N_8702,N_8365);
nor UO_9 (O_9,N_8427,N_8716);
nor UO_10 (O_10,N_9964,N_8744);
nand UO_11 (O_11,N_9433,N_9595);
or UO_12 (O_12,N_9890,N_9625);
nor UO_13 (O_13,N_9954,N_8985);
nand UO_14 (O_14,N_9701,N_8270);
nor UO_15 (O_15,N_9197,N_9104);
xor UO_16 (O_16,N_8456,N_9801);
and UO_17 (O_17,N_9153,N_8310);
nand UO_18 (O_18,N_8881,N_9839);
xor UO_19 (O_19,N_8708,N_8550);
nor UO_20 (O_20,N_9722,N_8722);
nor UO_21 (O_21,N_9194,N_8586);
nor UO_22 (O_22,N_8218,N_9350);
nand UO_23 (O_23,N_9323,N_9655);
nand UO_24 (O_24,N_9451,N_9003);
and UO_25 (O_25,N_9074,N_8866);
or UO_26 (O_26,N_8012,N_8600);
or UO_27 (O_27,N_9248,N_8139);
and UO_28 (O_28,N_9700,N_9647);
or UO_29 (O_29,N_8728,N_8158);
xnor UO_30 (O_30,N_8178,N_9804);
nand UO_31 (O_31,N_9468,N_9576);
nor UO_32 (O_32,N_9271,N_8052);
nand UO_33 (O_33,N_8583,N_8079);
nor UO_34 (O_34,N_9580,N_8418);
or UO_35 (O_35,N_9415,N_8833);
xor UO_36 (O_36,N_8650,N_8645);
or UO_37 (O_37,N_8925,N_9262);
and UO_38 (O_38,N_8268,N_8045);
nand UO_39 (O_39,N_9218,N_9151);
nand UO_40 (O_40,N_9965,N_8393);
and UO_41 (O_41,N_8413,N_8820);
nor UO_42 (O_42,N_8942,N_9283);
or UO_43 (O_43,N_8164,N_9116);
nor UO_44 (O_44,N_8569,N_9037);
nor UO_45 (O_45,N_8118,N_9398);
or UO_46 (O_46,N_9048,N_8755);
nand UO_47 (O_47,N_9481,N_9669);
and UO_48 (O_48,N_8732,N_9640);
nand UO_49 (O_49,N_8077,N_9447);
nand UO_50 (O_50,N_9972,N_8912);
or UO_51 (O_51,N_9548,N_9879);
and UO_52 (O_52,N_8132,N_9476);
nor UO_53 (O_53,N_9875,N_9568);
nand UO_54 (O_54,N_8115,N_8256);
nor UO_55 (O_55,N_8900,N_9742);
or UO_56 (O_56,N_9738,N_9612);
and UO_57 (O_57,N_8756,N_9361);
xnor UO_58 (O_58,N_8599,N_8291);
and UO_59 (O_59,N_9045,N_9933);
nor UO_60 (O_60,N_8053,N_8778);
nor UO_61 (O_61,N_9908,N_9970);
and UO_62 (O_62,N_8395,N_9454);
and UO_63 (O_63,N_8886,N_8069);
nand UO_64 (O_64,N_9621,N_8368);
nor UO_65 (O_65,N_9991,N_8621);
or UO_66 (O_66,N_8305,N_8404);
or UO_67 (O_67,N_8027,N_8709);
and UO_68 (O_68,N_8211,N_9178);
xor UO_69 (O_69,N_8814,N_8008);
nor UO_70 (O_70,N_8594,N_9850);
or UO_71 (O_71,N_8482,N_8514);
nor UO_72 (O_72,N_9786,N_8417);
nor UO_73 (O_73,N_8198,N_8160);
and UO_74 (O_74,N_8521,N_9598);
or UO_75 (O_75,N_9511,N_8124);
nand UO_76 (O_76,N_8440,N_9973);
nor UO_77 (O_77,N_9622,N_9946);
nand UO_78 (O_78,N_8789,N_8672);
or UO_79 (O_79,N_9402,N_9697);
nor UO_80 (O_80,N_9223,N_8745);
nand UO_81 (O_81,N_9668,N_9232);
nor UO_82 (O_82,N_9900,N_9921);
or UO_83 (O_83,N_9799,N_9374);
or UO_84 (O_84,N_9077,N_8014);
nor UO_85 (O_85,N_8379,N_9624);
or UO_86 (O_86,N_8346,N_8739);
and UO_87 (O_87,N_9175,N_9031);
xnor UO_88 (O_88,N_8047,N_8625);
xor UO_89 (O_89,N_8960,N_9211);
or UO_90 (O_90,N_8041,N_8236);
nor UO_91 (O_91,N_9030,N_9174);
and UO_92 (O_92,N_8332,N_8114);
and UO_93 (O_93,N_9711,N_9520);
nand UO_94 (O_94,N_8197,N_8390);
and UO_95 (O_95,N_8473,N_9001);
or UO_96 (O_96,N_8434,N_9446);
nand UO_97 (O_97,N_8363,N_8610);
or UO_98 (O_98,N_8408,N_9133);
and UO_99 (O_99,N_9241,N_9391);
and UO_100 (O_100,N_9676,N_8808);
nor UO_101 (O_101,N_9756,N_9033);
and UO_102 (O_102,N_9524,N_8138);
or UO_103 (O_103,N_8227,N_9382);
nor UO_104 (O_104,N_9322,N_8131);
nor UO_105 (O_105,N_9103,N_9995);
or UO_106 (O_106,N_9845,N_9670);
and UO_107 (O_107,N_8604,N_9618);
nand UO_108 (O_108,N_9543,N_9971);
xor UO_109 (O_109,N_9943,N_8328);
or UO_110 (O_110,N_8264,N_8290);
nor UO_111 (O_111,N_8885,N_9502);
nor UO_112 (O_112,N_9523,N_9583);
nor UO_113 (O_113,N_8319,N_8558);
and UO_114 (O_114,N_8286,N_8590);
nand UO_115 (O_115,N_9805,N_9440);
xnor UO_116 (O_116,N_8964,N_8834);
xnor UO_117 (O_117,N_9975,N_8910);
xnor UO_118 (O_118,N_8535,N_8635);
and UO_119 (O_119,N_9063,N_9210);
or UO_120 (O_120,N_9388,N_9196);
and UO_121 (O_121,N_9245,N_8208);
and UO_122 (O_122,N_8002,N_8001);
nand UO_123 (O_123,N_8096,N_8579);
nand UO_124 (O_124,N_8651,N_9575);
or UO_125 (O_125,N_8009,N_9827);
nor UO_126 (O_126,N_9819,N_9633);
nor UO_127 (O_127,N_9263,N_8216);
xnor UO_128 (O_128,N_8729,N_8593);
xnor UO_129 (O_129,N_9076,N_9560);
nand UO_130 (O_130,N_8415,N_9464);
and UO_131 (O_131,N_8752,N_9824);
nor UO_132 (O_132,N_8509,N_9791);
xor UO_133 (O_133,N_8342,N_9022);
xor UO_134 (O_134,N_9491,N_9088);
nor UO_135 (O_135,N_9120,N_8381);
and UO_136 (O_136,N_9741,N_8090);
nor UO_137 (O_137,N_8828,N_8750);
nand UO_138 (O_138,N_8543,N_9069);
xor UO_139 (O_139,N_8813,N_9254);
and UO_140 (O_140,N_9111,N_8083);
nor UO_141 (O_141,N_8260,N_9316);
nand UO_142 (O_142,N_8282,N_9499);
and UO_143 (O_143,N_9328,N_8458);
or UO_144 (O_144,N_8928,N_9472);
xor UO_145 (O_145,N_8220,N_9760);
and UO_146 (O_146,N_8981,N_8715);
xnor UO_147 (O_147,N_9627,N_8524);
or UO_148 (O_148,N_8996,N_8588);
nor UO_149 (O_149,N_9070,N_8006);
and UO_150 (O_150,N_8633,N_9577);
nand UO_151 (O_151,N_8773,N_9772);
or UO_152 (O_152,N_9299,N_9555);
nor UO_153 (O_153,N_8605,N_8483);
nand UO_154 (O_154,N_8991,N_8309);
nand UO_155 (O_155,N_8140,N_9787);
or UO_156 (O_156,N_9895,N_8816);
and UO_157 (O_157,N_9869,N_9993);
and UO_158 (O_158,N_8082,N_9609);
or UO_159 (O_159,N_9565,N_8724);
or UO_160 (O_160,N_9237,N_9025);
nor UO_161 (O_161,N_9118,N_9778);
nor UO_162 (O_162,N_9749,N_9364);
and UO_163 (O_163,N_8312,N_9279);
nand UO_164 (O_164,N_8177,N_9922);
nand UO_165 (O_165,N_9035,N_9808);
or UO_166 (O_166,N_9657,N_9333);
xnor UO_167 (O_167,N_8909,N_9978);
xor UO_168 (O_168,N_9537,N_9958);
or UO_169 (O_169,N_8684,N_8011);
nor UO_170 (O_170,N_9383,N_9847);
or UO_171 (O_171,N_9286,N_8457);
nand UO_172 (O_172,N_9892,N_9252);
nor UO_173 (O_173,N_8343,N_9157);
nor UO_174 (O_174,N_8696,N_9066);
and UO_175 (O_175,N_8636,N_8430);
nor UO_176 (O_176,N_8399,N_8459);
or UO_177 (O_177,N_8400,N_8125);
or UO_178 (O_178,N_9463,N_9055);
or UO_179 (O_179,N_9251,N_8941);
or UO_180 (O_180,N_8801,N_9654);
nor UO_181 (O_181,N_9369,N_8529);
or UO_182 (O_182,N_8134,N_8876);
nand UO_183 (O_183,N_9550,N_8480);
xor UO_184 (O_184,N_9950,N_9441);
nand UO_185 (O_185,N_9909,N_8210);
and UO_186 (O_186,N_8643,N_8331);
or UO_187 (O_187,N_8683,N_9795);
or UO_188 (O_188,N_8168,N_8940);
xor UO_189 (O_189,N_9848,N_9739);
and UO_190 (O_190,N_8230,N_9390);
or UO_191 (O_191,N_8463,N_8503);
xnor UO_192 (O_192,N_9256,N_8105);
and UO_193 (O_193,N_8235,N_8566);
nand UO_194 (O_194,N_8425,N_9866);
and UO_195 (O_195,N_9616,N_9702);
nor UO_196 (O_196,N_9710,N_9338);
and UO_197 (O_197,N_9835,N_9871);
nor UO_198 (O_198,N_9751,N_8841);
or UO_199 (O_199,N_8967,N_9367);
nor UO_200 (O_200,N_8426,N_8066);
nor UO_201 (O_201,N_8574,N_8288);
nor UO_202 (O_202,N_9275,N_8809);
and UO_203 (O_203,N_9889,N_8918);
nor UO_204 (O_204,N_8511,N_9628);
and UO_205 (O_205,N_9243,N_9893);
xor UO_206 (O_206,N_8762,N_8961);
nor UO_207 (O_207,N_9278,N_9794);
nor UO_208 (O_208,N_8970,N_9149);
nand UO_209 (O_209,N_9525,N_9311);
nand UO_210 (O_210,N_9142,N_9920);
and UO_211 (O_211,N_8545,N_8234);
nor UO_212 (O_212,N_9161,N_9042);
nor UO_213 (O_213,N_9306,N_8063);
xor UO_214 (O_214,N_8439,N_8076);
nor UO_215 (O_215,N_9230,N_8573);
and UO_216 (O_216,N_8436,N_9914);
xor UO_217 (O_217,N_8267,N_8423);
nand UO_218 (O_218,N_8403,N_9665);
nand UO_219 (O_219,N_8973,N_9200);
nor UO_220 (O_220,N_9677,N_9268);
nor UO_221 (O_221,N_8073,N_8420);
nand UO_222 (O_222,N_9138,N_8740);
and UO_223 (O_223,N_8274,N_8100);
and UO_224 (O_224,N_9117,N_8632);
and UO_225 (O_225,N_9663,N_8298);
or UO_226 (O_226,N_8107,N_9354);
nor UO_227 (O_227,N_8741,N_8029);
nand UO_228 (O_228,N_9660,N_9018);
and UO_229 (O_229,N_8450,N_8384);
or UO_230 (O_230,N_8944,N_8712);
and UO_231 (O_231,N_9498,N_9864);
and UO_232 (O_232,N_9957,N_9027);
and UO_233 (O_233,N_8631,N_8028);
or UO_234 (O_234,N_8142,N_9007);
nand UO_235 (O_235,N_8104,N_9596);
nor UO_236 (O_236,N_8717,N_9998);
nor UO_237 (O_237,N_9693,N_9384);
and UO_238 (O_238,N_9317,N_9122);
nand UO_239 (O_239,N_9277,N_8923);
nor UO_240 (O_240,N_9486,N_8491);
or UO_241 (O_241,N_8540,N_8601);
nor UO_242 (O_242,N_8183,N_8850);
and UO_243 (O_243,N_8330,N_9708);
nand UO_244 (O_244,N_8931,N_8795);
xor UO_245 (O_245,N_8287,N_9770);
nor UO_246 (O_246,N_9352,N_9357);
and UO_247 (O_247,N_9290,N_9410);
and UO_248 (O_248,N_9154,N_8502);
or UO_249 (O_249,N_9399,N_8101);
nor UO_250 (O_250,N_8999,N_8464);
and UO_251 (O_251,N_8213,N_8562);
nor UO_252 (O_252,N_8432,N_9844);
and UO_253 (O_253,N_9461,N_8226);
and UO_254 (O_254,N_8054,N_8972);
nor UO_255 (O_255,N_8038,N_9615);
or UO_256 (O_256,N_9877,N_9611);
nand UO_257 (O_257,N_9891,N_8484);
and UO_258 (O_258,N_8322,N_8868);
nor UO_259 (O_259,N_8646,N_8182);
nor UO_260 (O_260,N_9928,N_8340);
nand UO_261 (O_261,N_9917,N_8081);
nand UO_262 (O_262,N_9959,N_8099);
nor UO_263 (O_263,N_8689,N_9132);
or UO_264 (O_264,N_9830,N_8007);
nor UO_265 (O_265,N_8068,N_8825);
nand UO_266 (O_266,N_9436,N_8893);
nor UO_267 (O_267,N_9485,N_8301);
or UO_268 (O_268,N_9409,N_9652);
and UO_269 (O_269,N_9777,N_8532);
or UO_270 (O_270,N_9788,N_8659);
nand UO_271 (O_271,N_9919,N_9029);
and UO_272 (O_272,N_8481,N_8341);
or UO_273 (O_273,N_8154,N_9811);
and UO_274 (O_274,N_8383,N_8751);
nand UO_275 (O_275,N_9293,N_8671);
xnor UO_276 (O_276,N_8576,N_8233);
nand UO_277 (O_277,N_8873,N_9162);
or UO_278 (O_278,N_9996,N_8842);
nor UO_279 (O_279,N_8926,N_8348);
nand UO_280 (O_280,N_8257,N_9515);
or UO_281 (O_281,N_8405,N_9462);
nor UO_282 (O_282,N_9617,N_9189);
nand UO_283 (O_283,N_9765,N_8629);
or UO_284 (O_284,N_8065,N_9825);
nor UO_285 (O_285,N_8162,N_8541);
or UO_286 (O_286,N_8510,N_8582);
or UO_287 (O_287,N_8958,N_9816);
and UO_288 (O_288,N_9868,N_8385);
nor UO_289 (O_289,N_8171,N_9821);
xor UO_290 (O_290,N_9872,N_9156);
nand UO_291 (O_291,N_9865,N_9150);
nor UO_292 (O_292,N_8496,N_9796);
or UO_293 (O_293,N_9692,N_8754);
nand UO_294 (O_294,N_8951,N_8655);
and UO_295 (O_295,N_8623,N_9510);
nand UO_296 (O_296,N_9695,N_8244);
and UO_297 (O_297,N_9563,N_9470);
nor UO_298 (O_298,N_8983,N_8325);
or UO_299 (O_299,N_8731,N_9160);
xor UO_300 (O_300,N_9107,N_8902);
nand UO_301 (O_301,N_8145,N_9956);
or UO_302 (O_302,N_8278,N_8534);
nand UO_303 (O_303,N_8719,N_9509);
nor UO_304 (O_304,N_9098,N_8377);
nor UO_305 (O_305,N_9960,N_8544);
nand UO_306 (O_306,N_9773,N_9925);
and UO_307 (O_307,N_8221,N_9423);
nand UO_308 (O_308,N_8552,N_8777);
or UO_309 (O_309,N_9767,N_9536);
nor UO_310 (O_310,N_9280,N_9818);
xor UO_311 (O_311,N_8567,N_8232);
nor UO_312 (O_312,N_8688,N_8357);
nor UO_313 (O_313,N_8039,N_9184);
or UO_314 (O_314,N_8311,N_8258);
nand UO_315 (O_315,N_8898,N_8506);
and UO_316 (O_316,N_8191,N_8725);
nor UO_317 (O_317,N_8085,N_8438);
nor UO_318 (O_318,N_9375,N_8176);
nand UO_319 (O_319,N_8091,N_9547);
nand UO_320 (O_320,N_9300,N_9664);
or UO_321 (O_321,N_8849,N_8686);
and UO_322 (O_322,N_8224,N_8180);
and UO_323 (O_323,N_8392,N_9473);
nor UO_324 (O_324,N_9812,N_9424);
nand UO_325 (O_325,N_8252,N_9852);
nor UO_326 (O_326,N_8159,N_9253);
nand UO_327 (O_327,N_9477,N_8674);
nand UO_328 (O_328,N_8296,N_9726);
nor UO_329 (O_329,N_8272,N_8949);
nor UO_330 (O_330,N_8818,N_9667);
or UO_331 (O_331,N_9714,N_8877);
nor UO_332 (O_332,N_9204,N_8811);
or UO_333 (O_333,N_9746,N_8067);
nor UO_334 (O_334,N_9556,N_8711);
nor UO_335 (O_335,N_9659,N_8641);
or UO_336 (O_336,N_9949,N_8507);
nand UO_337 (O_337,N_8147,N_8092);
nor UO_338 (O_338,N_9854,N_8229);
and UO_339 (O_339,N_8043,N_8854);
nor UO_340 (O_340,N_8705,N_9331);
or UO_341 (O_341,N_9059,N_9836);
and UO_342 (O_342,N_8995,N_9255);
nor UO_343 (O_343,N_8285,N_8794);
or UO_344 (O_344,N_9097,N_9748);
nor UO_345 (O_345,N_9310,N_9587);
and UO_346 (O_346,N_9078,N_9720);
nand UO_347 (O_347,N_9140,N_8447);
or UO_348 (O_348,N_8767,N_8826);
nor UO_349 (O_349,N_8119,N_9800);
or UO_350 (O_350,N_8021,N_8060);
or UO_351 (O_351,N_8974,N_8157);
or UO_352 (O_352,N_8206,N_9744);
or UO_353 (O_353,N_9356,N_8130);
nand UO_354 (O_354,N_9932,N_9155);
or UO_355 (O_355,N_9238,N_9124);
or UO_356 (O_356,N_9802,N_8707);
and UO_357 (O_357,N_8493,N_8861);
and UO_358 (O_358,N_8865,N_9158);
and UO_359 (O_359,N_8787,N_9371);
or UO_360 (O_360,N_9389,N_9206);
nor UO_361 (O_361,N_8106,N_9119);
xnor UO_362 (O_362,N_9434,N_8397);
or UO_363 (O_363,N_8314,N_9139);
or UO_364 (O_364,N_9503,N_8017);
or UO_365 (O_365,N_9163,N_8649);
nor UO_366 (O_366,N_8986,N_9782);
or UO_367 (O_367,N_9784,N_8468);
or UO_368 (O_368,N_8609,N_9820);
and UO_369 (O_369,N_9480,N_8677);
nand UO_370 (O_370,N_9336,N_8097);
nand UO_371 (O_371,N_8660,N_8113);
or UO_372 (O_372,N_8061,N_9519);
and UO_373 (O_373,N_8003,N_9180);
nand UO_374 (O_374,N_8108,N_8366);
and UO_375 (O_375,N_8945,N_9608);
nand UO_376 (O_376,N_8283,N_9539);
nand UO_377 (O_377,N_8701,N_8966);
or UO_378 (O_378,N_9452,N_8444);
nor UO_379 (O_379,N_8186,N_9913);
and UO_380 (O_380,N_9169,N_9507);
nor UO_381 (O_381,N_8334,N_9420);
and UO_382 (O_382,N_8917,N_8831);
and UO_383 (O_383,N_8652,N_8129);
or UO_384 (O_384,N_9730,N_9863);
and UO_385 (O_385,N_9172,N_9947);
nand UO_386 (O_386,N_8058,N_8783);
xnor UO_387 (O_387,N_8475,N_9396);
nor UO_388 (O_388,N_9689,N_9857);
nand UO_389 (O_389,N_9591,N_8477);
nand UO_390 (O_390,N_8155,N_9792);
nor UO_391 (O_391,N_9842,N_8442);
or UO_392 (O_392,N_9906,N_8152);
xor UO_393 (O_393,N_8293,N_9449);
nor UO_394 (O_394,N_8163,N_9638);
or UO_395 (O_395,N_8676,N_9060);
xnor UO_396 (O_396,N_8919,N_9757);
and UO_397 (O_397,N_9724,N_9532);
nor UO_398 (O_398,N_9675,N_8374);
nand UO_399 (O_399,N_8580,N_9766);
nand UO_400 (O_400,N_8888,N_8915);
nor UO_401 (O_401,N_8143,N_9475);
and UO_402 (O_402,N_9345,N_8315);
or UO_403 (O_403,N_9923,N_8345);
or UO_404 (O_404,N_9101,N_9079);
or UO_405 (O_405,N_8044,N_8832);
and UO_406 (O_406,N_9176,N_9425);
nand UO_407 (O_407,N_9859,N_9980);
nor UO_408 (O_408,N_9363,N_8760);
nor UO_409 (O_409,N_8978,N_8372);
nand UO_410 (O_410,N_8495,N_9907);
nand UO_411 (O_411,N_9224,N_9177);
nor UO_412 (O_412,N_8890,N_9883);
or UO_413 (O_413,N_8513,N_8367);
nand UO_414 (O_414,N_9026,N_9554);
and UO_415 (O_415,N_8019,N_8875);
nand UO_416 (O_416,N_9006,N_8431);
or UO_417 (O_417,N_9584,N_9228);
nand UO_418 (O_418,N_9487,N_9731);
nand UO_419 (O_419,N_8557,N_8467);
or UO_420 (O_420,N_8515,N_8170);
or UO_421 (O_421,N_9202,N_9032);
nand UO_422 (O_422,N_9458,N_9259);
nand UO_423 (O_423,N_8694,N_8589);
and UO_424 (O_424,N_9421,N_9979);
nand UO_425 (O_425,N_8608,N_9335);
nand UO_426 (O_426,N_8804,N_8084);
xnor UO_427 (O_427,N_8214,N_8896);
and UO_428 (O_428,N_9797,N_9745);
or UO_429 (O_429,N_8714,N_8273);
nor UO_430 (O_430,N_8336,N_9337);
or UO_431 (O_431,N_8316,N_9272);
and UO_432 (O_432,N_8523,N_9453);
nand UO_433 (O_433,N_9942,N_8271);
nor UO_434 (O_434,N_9405,N_9108);
and UO_435 (O_435,N_9173,N_8990);
or UO_436 (O_436,N_9517,N_9817);
nor UO_437 (O_437,N_8680,N_9634);
xor UO_438 (O_438,N_8547,N_8169);
xor UO_439 (O_439,N_8144,N_8355);
nor UO_440 (O_440,N_9858,N_9083);
and UO_441 (O_441,N_8056,N_9043);
nand UO_442 (O_442,N_9106,N_8872);
or UO_443 (O_443,N_9841,N_9951);
and UO_444 (O_444,N_9244,N_9953);
and UO_445 (O_445,N_9603,N_9269);
and UO_446 (O_446,N_8812,N_9630);
nor UO_447 (O_447,N_9057,N_8292);
nand UO_448 (O_448,N_9780,N_8173);
and UO_449 (O_449,N_8691,N_8046);
nor UO_450 (O_450,N_8333,N_8614);
or UO_451 (O_451,N_8059,N_8772);
and UO_452 (O_452,N_8611,N_8947);
nor UO_453 (O_453,N_9302,N_8098);
nand UO_454 (O_454,N_9944,N_8644);
and UO_455 (O_455,N_9082,N_8905);
or UO_456 (O_456,N_8735,N_9192);
xor UO_457 (O_457,N_8351,N_8955);
or UO_458 (O_458,N_8613,N_8803);
xor UO_459 (O_459,N_8819,N_8591);
nand UO_460 (O_460,N_8499,N_8770);
nor UO_461 (O_461,N_9684,N_9915);
nor UO_462 (O_462,N_8080,N_8102);
nand UO_463 (O_463,N_9831,N_9886);
and UO_464 (O_464,N_8254,N_9823);
and UO_465 (O_465,N_9179,N_8469);
nor UO_466 (O_466,N_9058,N_9986);
nand UO_467 (O_467,N_9100,N_8031);
xnor UO_468 (O_468,N_8276,N_8259);
and UO_469 (O_469,N_9431,N_9650);
and UO_470 (O_470,N_8761,N_8856);
and UO_471 (O_471,N_9068,N_8690);
nand UO_472 (O_472,N_8202,N_8658);
or UO_473 (O_473,N_9687,N_9732);
and UO_474 (O_474,N_8194,N_9287);
and UO_475 (O_475,N_9743,N_9728);
and UO_476 (O_476,N_8817,N_8209);
xnor UO_477 (O_477,N_8560,N_8454);
nand UO_478 (O_478,N_8713,N_9329);
and UO_479 (O_479,N_9094,N_8335);
nor UO_480 (O_480,N_8556,N_8137);
and UO_481 (O_481,N_9240,N_8013);
or UO_482 (O_482,N_8606,N_8703);
or UO_483 (O_483,N_9793,N_8279);
nand UO_484 (O_484,N_8821,N_9394);
or UO_485 (O_485,N_8771,N_8699);
and UO_486 (O_486,N_8373,N_9977);
nor UO_487 (O_487,N_9324,N_9401);
and UO_488 (O_488,N_8205,N_8022);
and UO_489 (O_489,N_9775,N_8110);
nor UO_490 (O_490,N_8836,N_9614);
and UO_491 (O_491,N_9067,N_8538);
or UO_492 (O_492,N_8241,N_9168);
nor UO_493 (O_493,N_8776,N_8853);
nand UO_494 (O_494,N_9312,N_9571);
and UO_495 (O_495,N_8758,N_9081);
nand UO_496 (O_496,N_8398,N_9181);
and UO_497 (O_497,N_8913,N_8308);
or UO_498 (O_498,N_9867,N_8517);
or UO_499 (O_499,N_8706,N_8838);
nor UO_500 (O_500,N_9235,N_9725);
nor UO_501 (O_501,N_9937,N_8135);
or UO_502 (O_502,N_8975,N_9040);
nand UO_503 (O_503,N_9273,N_8294);
and UO_504 (O_504,N_9626,N_9535);
nor UO_505 (O_505,N_9414,N_8466);
nor UO_506 (O_506,N_8988,N_8412);
and UO_507 (O_507,N_9435,N_9341);
or UO_508 (O_508,N_8738,N_9207);
or UO_509 (O_509,N_9901,N_9916);
nor UO_510 (O_510,N_8883,N_9236);
nor UO_511 (O_511,N_9750,N_8035);
or UO_512 (O_512,N_8791,N_9636);
or UO_513 (O_513,N_8485,N_9504);
nand UO_514 (O_514,N_8807,N_9826);
and UO_515 (O_515,N_9455,N_9216);
or UO_516 (O_516,N_8174,N_8533);
nor UO_517 (O_517,N_9247,N_9274);
and UO_518 (O_518,N_8570,N_8307);
or UO_519 (O_519,N_8492,N_9264);
and UO_520 (O_520,N_8402,N_8572);
or UO_521 (O_521,N_9047,N_9939);
nand UO_522 (O_522,N_8441,N_9736);
nand UO_523 (O_523,N_8269,N_9976);
nand UO_524 (O_524,N_8843,N_9755);
nand UO_525 (O_525,N_9326,N_9512);
nand UO_526 (O_526,N_8536,N_8040);
and UO_527 (O_527,N_8980,N_8984);
and UO_528 (O_528,N_8184,N_9723);
nor UO_529 (O_529,N_8721,N_9833);
nand UO_530 (O_530,N_8927,N_8637);
nand UO_531 (O_531,N_8238,N_9690);
and UO_532 (O_532,N_9763,N_9347);
nand UO_533 (O_533,N_8406,N_8387);
or UO_534 (O_534,N_8020,N_9144);
and UO_535 (O_535,N_9378,N_8192);
xor UO_536 (O_536,N_9945,N_8490);
and UO_537 (O_537,N_8049,N_9605);
and UO_538 (O_538,N_8790,N_8117);
and UO_539 (O_539,N_9205,N_8443);
or UO_540 (O_540,N_8074,N_9589);
nor UO_541 (O_541,N_9131,N_8088);
and UO_542 (O_542,N_9814,N_9860);
xor UO_543 (O_543,N_8461,N_9837);
nand UO_544 (O_544,N_8111,N_9683);
nor UO_545 (O_545,N_8414,N_9559);
nor UO_546 (O_546,N_9769,N_8277);
or UO_547 (O_547,N_8971,N_8736);
or UO_548 (O_548,N_8126,N_8122);
or UO_549 (O_549,N_9360,N_8592);
nor UO_550 (O_550,N_8639,N_9903);
or UO_551 (O_551,N_9073,N_8223);
nand UO_552 (O_552,N_9145,N_9910);
or UO_553 (O_553,N_8640,N_9876);
or UO_554 (O_554,N_9296,N_9222);
or UO_555 (O_555,N_8784,N_9021);
and UO_556 (O_556,N_9696,N_9884);
nor UO_557 (O_557,N_9929,N_9988);
xor UO_558 (O_558,N_9759,N_8798);
or UO_559 (O_559,N_8445,N_8539);
nor UO_560 (O_560,N_8775,N_9494);
xor UO_561 (O_561,N_9721,N_9706);
nor UO_562 (O_562,N_8782,N_8622);
nor UO_563 (O_563,N_9052,N_8033);
and UO_564 (O_564,N_9561,N_9071);
nor UO_565 (O_565,N_9044,N_8284);
and UO_566 (O_566,N_8304,N_8847);
nor UO_567 (O_567,N_9553,N_9147);
xnor UO_568 (O_568,N_9645,N_8086);
or UO_569 (O_569,N_9170,N_8240);
and UO_570 (O_570,N_8032,N_8835);
or UO_571 (O_571,N_9346,N_9102);
and UO_572 (O_572,N_8994,N_8824);
nor UO_573 (O_573,N_9715,N_9653);
nand UO_574 (O_574,N_9191,N_9562);
or UO_575 (O_575,N_9303,N_9888);
nor UO_576 (O_576,N_9704,N_9182);
nor UO_577 (O_577,N_8879,N_8769);
or UO_578 (O_578,N_9962,N_9987);
nand UO_579 (O_579,N_9607,N_9096);
nand UO_580 (O_580,N_8429,N_9469);
xor UO_581 (O_581,N_9050,N_9387);
nor UO_582 (O_582,N_9505,N_9320);
nand UO_583 (O_583,N_8857,N_9266);
or UO_584 (O_584,N_8859,N_8700);
nor UO_585 (O_585,N_8478,N_9450);
or UO_586 (O_586,N_9694,N_8362);
or UO_587 (O_587,N_8196,N_8246);
and UO_588 (O_588,N_8887,N_8347);
and UO_589 (O_589,N_8799,N_9989);
nor UO_590 (O_590,N_8727,N_8253);
nor UO_591 (O_591,N_8977,N_9674);
or UO_592 (O_592,N_9362,N_9209);
or UO_593 (O_593,N_9619,N_8265);
xor UO_594 (O_594,N_8989,N_9112);
xor UO_595 (O_595,N_9557,N_8779);
nor UO_596 (O_596,N_8133,N_8249);
nand UO_597 (O_597,N_9544,N_8815);
and UO_598 (O_598,N_8656,N_8559);
nor UO_599 (O_599,N_8858,N_9092);
nand UO_600 (O_600,N_9002,N_8212);
nor UO_601 (O_601,N_8356,N_8231);
xor UO_602 (O_602,N_9250,N_8370);
nand UO_603 (O_603,N_9691,N_8810);
nor UO_604 (O_604,N_8626,N_8844);
nor UO_605 (O_605,N_8166,N_8939);
and UO_606 (O_606,N_8095,N_9528);
nor UO_607 (O_607,N_8952,N_8146);
nand UO_608 (O_608,N_9846,N_9783);
nor UO_609 (O_609,N_9948,N_9288);
and UO_610 (O_610,N_8979,N_9456);
or UO_611 (O_611,N_9529,N_9315);
and UO_612 (O_612,N_8071,N_9671);
nand UO_613 (O_613,N_8391,N_8969);
xor UO_614 (O_614,N_9459,N_8634);
and UO_615 (O_615,N_9134,N_9109);
and UO_616 (O_616,N_9861,N_8848);
nand UO_617 (O_617,N_9225,N_9406);
or UO_618 (O_618,N_8470,N_8584);
nor UO_619 (O_619,N_9992,N_8508);
or UO_620 (O_620,N_8300,N_8512);
and UO_621 (O_621,N_9128,N_9602);
or UO_622 (O_622,N_9581,N_9558);
and UO_623 (O_623,N_9952,N_9516);
or UO_624 (O_624,N_8565,N_9429);
nor UO_625 (O_625,N_8654,N_9474);
and UO_626 (O_626,N_9080,N_8612);
and UO_627 (O_627,N_9359,N_9567);
nand UO_628 (O_628,N_8852,N_8693);
or UO_629 (O_629,N_8516,N_8822);
or UO_630 (O_630,N_8109,N_8867);
and UO_631 (O_631,N_8638,N_8193);
or UO_632 (O_632,N_9164,N_8666);
nand UO_633 (O_633,N_9351,N_8959);
or UO_634 (O_634,N_8869,N_8668);
or UO_635 (O_635,N_9851,N_8121);
or UO_636 (O_636,N_9377,N_8930);
and UO_637 (O_637,N_8561,N_9193);
or UO_638 (O_638,N_9855,N_9213);
or UO_639 (O_639,N_8042,N_9137);
nand UO_640 (O_640,N_9610,N_8542);
and UO_641 (O_641,N_8723,N_8222);
nor UO_642 (O_642,N_9072,N_8797);
nor UO_643 (O_643,N_8034,N_8036);
nor UO_644 (O_644,N_9905,N_9930);
nand UO_645 (O_645,N_9672,N_8647);
or UO_646 (O_646,N_9428,N_8024);
or UO_647 (O_647,N_9566,N_9217);
or UO_648 (O_648,N_9585,N_8181);
nor UO_649 (O_649,N_8681,N_9764);
and UO_650 (O_650,N_9737,N_9620);
nand UO_651 (O_651,N_8765,N_9327);
xnor UO_652 (O_652,N_9552,N_8189);
and UO_653 (O_653,N_8907,N_9093);
and UO_654 (O_654,N_8749,N_8474);
nor UO_655 (O_655,N_8266,N_8156);
and UO_656 (O_656,N_9017,N_8860);
nor UO_657 (O_657,N_8657,N_9955);
or UO_658 (O_658,N_9500,N_8151);
and UO_659 (O_659,N_8548,N_9488);
nor UO_660 (O_660,N_9935,N_8757);
nor UO_661 (O_661,N_8518,N_9843);
nand UO_662 (O_662,N_9776,N_9203);
and UO_663 (O_663,N_9649,N_9422);
and UO_664 (O_664,N_9599,N_8653);
and UO_665 (O_665,N_8863,N_9894);
xor UO_666 (O_666,N_8748,N_9678);
xnor UO_667 (O_667,N_8823,N_8219);
xor UO_668 (O_668,N_8263,N_8829);
and UO_669 (O_669,N_9444,N_9495);
and UO_670 (O_670,N_8764,N_9829);
nand UO_671 (O_671,N_9099,N_9880);
xor UO_672 (O_672,N_9208,N_9212);
nor UO_673 (O_673,N_9358,N_9729);
nor UO_674 (O_674,N_8382,N_8389);
nor UO_675 (O_675,N_8720,N_9931);
or UO_676 (O_676,N_8884,N_9403);
and UO_677 (O_677,N_8245,N_9231);
and UO_678 (O_678,N_8993,N_9355);
or UO_679 (O_679,N_9090,N_9896);
and UO_680 (O_680,N_9121,N_9679);
and UO_681 (O_681,N_9912,N_9295);
nor UO_682 (O_682,N_9918,N_8698);
nand UO_683 (O_683,N_8120,N_8094);
and UO_684 (O_684,N_8595,N_8768);
or UO_685 (O_685,N_8929,N_8465);
nor UO_686 (O_686,N_8437,N_8954);
nand UO_687 (O_687,N_8175,N_8338);
nor UO_688 (O_688,N_8710,N_9870);
nand UO_689 (O_689,N_9265,N_8525);
or UO_690 (O_690,N_8661,N_8936);
nor UO_691 (O_691,N_8317,N_9400);
or UO_692 (O_692,N_8911,N_8933);
nand UO_693 (O_693,N_8489,N_8839);
nand UO_694 (O_694,N_8871,N_8358);
or UO_695 (O_695,N_9790,N_8837);
and UO_696 (O_696,N_9578,N_8242);
nand UO_697 (O_697,N_9199,N_8840);
nand UO_698 (O_698,N_9629,N_9289);
and UO_699 (O_699,N_9604,N_8766);
xnor UO_700 (O_700,N_9095,N_9221);
nor UO_701 (O_701,N_8215,N_9214);
nor UO_702 (O_702,N_8004,N_8354);
or UO_703 (O_703,N_9019,N_9445);
xnor UO_704 (O_704,N_8505,N_8070);
and UO_705 (O_705,N_9437,N_8275);
or UO_706 (O_706,N_8339,N_9934);
and UO_707 (O_707,N_8759,N_8932);
or UO_708 (O_708,N_8935,N_9443);
or UO_709 (O_709,N_8337,N_8603);
nor UO_710 (O_710,N_8048,N_9779);
or UO_711 (O_711,N_9343,N_9984);
nor UO_712 (O_712,N_8785,N_9342);
or UO_713 (O_713,N_8892,N_9513);
nor UO_714 (O_714,N_9056,N_9887);
nand UO_715 (O_715,N_8281,N_9590);
xnor UO_716 (O_716,N_9261,N_8568);
and UO_717 (O_717,N_9249,N_8624);
nor UO_718 (O_718,N_9015,N_9054);
nor UO_719 (O_719,N_9822,N_8320);
or UO_720 (O_720,N_9064,N_9774);
or UO_721 (O_721,N_8846,N_9735);
xor UO_722 (O_722,N_9166,N_8016);
and UO_723 (O_723,N_8669,N_9856);
and UO_724 (O_724,N_8504,N_8161);
nor UO_725 (O_725,N_8718,N_9061);
xor UO_726 (O_726,N_8862,N_8453);
nor UO_727 (O_727,N_9990,N_8963);
or UO_728 (O_728,N_9999,N_8401);
or UO_729 (O_729,N_9034,N_9276);
or UO_730 (O_730,N_9085,N_8921);
and UO_731 (O_731,N_8904,N_8737);
nand UO_732 (O_732,N_8673,N_8500);
or UO_733 (O_733,N_8497,N_9298);
or UO_734 (O_734,N_9038,N_8239);
or UO_735 (O_735,N_9297,N_8141);
xor UO_736 (O_736,N_9386,N_8627);
nand UO_737 (O_737,N_9187,N_8025);
and UO_738 (O_738,N_9651,N_9281);
and UO_739 (O_739,N_9215,N_9878);
or UO_740 (O_740,N_9573,N_8498);
and UO_741 (O_741,N_8578,N_9457);
nor UO_742 (O_742,N_8010,N_8476);
nand UO_743 (O_743,N_9834,N_9167);
and UO_744 (O_744,N_9219,N_8962);
and UO_745 (O_745,N_8692,N_9304);
and UO_746 (O_746,N_8409,N_8956);
and UO_747 (O_747,N_9798,N_9680);
nand UO_748 (O_748,N_8380,N_9803);
nor UO_749 (O_749,N_9483,N_9041);
xnor UO_750 (O_750,N_9762,N_9368);
or UO_751 (O_751,N_8185,N_8237);
nand UO_752 (O_752,N_9530,N_8897);
nor UO_753 (O_753,N_9688,N_9319);
or UO_754 (O_754,N_9049,N_9188);
nor UO_755 (O_755,N_9564,N_8922);
and UO_756 (O_756,N_9601,N_9969);
or UO_757 (O_757,N_9091,N_8449);
or UO_758 (O_758,N_8424,N_9234);
and UO_759 (O_759,N_8796,N_9353);
nor UO_760 (O_760,N_8250,N_8864);
nand UO_761 (O_761,N_9753,N_9666);
xnor UO_762 (O_762,N_9902,N_9013);
and UO_763 (O_763,N_8078,N_9028);
or UO_764 (O_764,N_8255,N_8148);
nor UO_765 (O_765,N_9257,N_8326);
and UO_766 (O_766,N_9039,N_8306);
nor UO_767 (O_767,N_8786,N_9639);
nand UO_768 (O_768,N_9938,N_8217);
nor UO_769 (O_769,N_8527,N_9592);
or UO_770 (O_770,N_8127,N_9712);
and UO_771 (O_771,N_9911,N_8695);
and UO_772 (O_772,N_9961,N_9994);
xnor UO_773 (O_773,N_9897,N_8128);
and UO_774 (O_774,N_8998,N_9635);
nand UO_775 (O_775,N_9012,N_8916);
nand UO_776 (O_776,N_9632,N_8575);
and UO_777 (O_777,N_9407,N_9974);
nor UO_778 (O_778,N_8563,N_9201);
or UO_779 (O_779,N_9471,N_9717);
nand UO_780 (O_780,N_9141,N_9482);
nand UO_781 (O_781,N_9314,N_8522);
or UO_782 (O_782,N_9682,N_8982);
nor UO_783 (O_783,N_8526,N_9227);
or UO_784 (O_784,N_9718,N_9549);
and UO_785 (O_785,N_8486,N_8103);
nor UO_786 (O_786,N_8630,N_9190);
and UO_787 (O_787,N_8302,N_9086);
or UO_788 (O_788,N_9260,N_9586);
and UO_789 (O_789,N_9853,N_9344);
or UO_790 (O_790,N_8802,N_8344);
nor UO_791 (O_791,N_8199,N_8726);
xnor UO_792 (O_792,N_8243,N_9439);
nor UO_793 (O_793,N_9171,N_8321);
nor UO_794 (O_794,N_9014,N_9198);
nor UO_795 (O_795,N_9658,N_8571);
and UO_796 (O_796,N_8855,N_9533);
nand UO_797 (O_797,N_8149,N_8908);
nor UO_798 (O_798,N_8551,N_9478);
and UO_799 (O_799,N_9004,N_8386);
nand UO_800 (O_800,N_8806,N_9129);
nand UO_801 (O_801,N_9963,N_9501);
and UO_802 (O_802,N_9940,N_9417);
nand UO_803 (O_803,N_8553,N_8329);
or UO_804 (O_804,N_9771,N_9114);
or UO_805 (O_805,N_8388,N_9641);
nor UO_806 (O_806,N_8297,N_9642);
or UO_807 (O_807,N_9397,N_8167);
nor UO_808 (O_808,N_8587,N_8793);
nor UO_809 (O_809,N_9703,N_9024);
and UO_810 (O_810,N_9904,N_8055);
nand UO_811 (O_811,N_8360,N_8228);
nand UO_812 (O_812,N_8747,N_9113);
nor UO_813 (O_813,N_9419,N_8487);
or UO_814 (O_814,N_9165,N_8997);
and UO_815 (O_815,N_9385,N_8188);
nor UO_816 (O_816,N_8585,N_9631);
nor UO_817 (O_817,N_8742,N_8165);
and UO_818 (O_818,N_8037,N_8943);
and UO_819 (O_819,N_9365,N_9152);
and UO_820 (O_820,N_9968,N_8891);
nand UO_821 (O_821,N_9699,N_9882);
nor UO_822 (O_822,N_8899,N_8597);
nor UO_823 (O_823,N_8416,N_8204);
nor UO_824 (O_824,N_8471,N_8153);
nor UO_825 (O_825,N_9643,N_8675);
or UO_826 (O_826,N_9159,N_9125);
or UO_827 (O_827,N_8446,N_8247);
nor UO_828 (O_828,N_9412,N_9418);
xnor UO_829 (O_829,N_8615,N_8448);
nand UO_830 (O_830,N_9579,N_9479);
nor UO_831 (O_831,N_9709,N_9413);
or UO_832 (O_832,N_9467,N_9983);
and UO_833 (O_833,N_8976,N_9183);
nor UO_834 (O_834,N_8678,N_9540);
nand UO_835 (O_835,N_9809,N_9348);
or UO_836 (O_836,N_9569,N_9572);
and UO_837 (O_837,N_8889,N_9489);
nor UO_838 (O_838,N_9233,N_9873);
and UO_839 (O_839,N_9526,N_9810);
nand UO_840 (O_840,N_9815,N_8472);
and UO_841 (O_841,N_8878,N_9226);
nand UO_842 (O_842,N_9325,N_8057);
nand UO_843 (O_843,N_9597,N_9985);
or UO_844 (O_844,N_8598,N_9541);
nor UO_845 (O_845,N_8596,N_8378);
and UO_846 (O_846,N_8350,N_9136);
nor UO_847 (O_847,N_8018,N_9518);
nor UO_848 (O_848,N_8396,N_9705);
or UO_849 (O_849,N_9508,N_8555);
nand UO_850 (O_850,N_8528,N_8375);
or UO_851 (O_851,N_9734,N_8546);
nand UO_852 (O_852,N_9828,N_8501);
and UO_853 (O_853,N_8251,N_9239);
nand UO_854 (O_854,N_8617,N_9514);
and UO_855 (O_855,N_8581,N_8364);
nor UO_856 (O_856,N_8261,N_8679);
nor UO_857 (O_857,N_9448,N_9673);
xnor UO_858 (O_858,N_8662,N_8648);
nor UO_859 (O_859,N_8313,N_8179);
and UO_860 (O_860,N_9332,N_8421);
nor UO_861 (O_861,N_8200,N_8903);
and UO_862 (O_862,N_9105,N_9008);
nand UO_863 (O_863,N_8618,N_8262);
nor UO_864 (O_864,N_8937,N_8946);
xnor UO_865 (O_865,N_9781,N_9941);
nand UO_866 (O_866,N_8299,N_9807);
and UO_867 (O_867,N_9613,N_9656);
and UO_868 (O_868,N_9143,N_9698);
nand UO_869 (O_869,N_8451,N_8950);
xor UO_870 (O_870,N_9570,N_9531);
nand UO_871 (O_871,N_8327,N_8554);
and UO_872 (O_872,N_9686,N_9594);
and UO_873 (O_873,N_9246,N_9648);
nor UO_874 (O_874,N_8150,N_9307);
nor UO_875 (O_875,N_9005,N_9662);
and UO_876 (O_876,N_9785,N_9849);
nand UO_877 (O_877,N_9292,N_8050);
and UO_878 (O_878,N_9600,N_9862);
xnor UO_879 (O_879,N_9924,N_8488);
or UO_880 (O_880,N_9318,N_9606);
nor UO_881 (O_881,N_9305,N_9126);
or UO_882 (O_882,N_9110,N_9981);
xor UO_883 (O_883,N_9546,N_9716);
xnor UO_884 (O_884,N_9885,N_8577);
and UO_885 (O_885,N_9582,N_8920);
and UO_886 (O_886,N_9372,N_9393);
and UO_887 (O_887,N_8934,N_9898);
nand UO_888 (O_888,N_9349,N_9115);
and UO_889 (O_889,N_9496,N_9392);
or UO_890 (O_890,N_8687,N_8394);
nor UO_891 (O_891,N_8323,N_9493);
and UO_892 (O_892,N_8602,N_9465);
or UO_893 (O_893,N_8827,N_9733);
or UO_894 (O_894,N_9340,N_8620);
and UO_895 (O_895,N_8564,N_8520);
xor UO_896 (O_896,N_9813,N_8026);
and UO_897 (O_897,N_9020,N_8000);
nand UO_898 (O_898,N_9339,N_9551);
xor UO_899 (O_899,N_8407,N_9294);
nand UO_900 (O_900,N_8733,N_9334);
and UO_901 (O_901,N_9130,N_9982);
or UO_902 (O_902,N_8452,N_9838);
xnor UO_903 (O_903,N_8410,N_9408);
and UO_904 (O_904,N_9768,N_8968);
nand UO_905 (O_905,N_9661,N_9053);
and UO_906 (O_906,N_8894,N_8015);
and UO_907 (O_907,N_9427,N_9395);
or UO_908 (O_908,N_8830,N_8361);
nand UO_909 (O_909,N_8203,N_9713);
nand UO_910 (O_910,N_9997,N_9538);
nor UO_911 (O_911,N_9681,N_9148);
and UO_912 (O_912,N_9727,N_9011);
and UO_913 (O_913,N_9270,N_9484);
nor UO_914 (O_914,N_8324,N_9899);
or UO_915 (O_915,N_9308,N_8628);
nand UO_916 (O_916,N_9285,N_9065);
or UO_917 (O_917,N_9754,N_9637);
xor UO_918 (O_918,N_9545,N_8187);
xnor UO_919 (O_919,N_9542,N_8136);
or UO_920 (O_920,N_9740,N_9747);
xnor UO_921 (O_921,N_8064,N_8280);
or UO_922 (O_922,N_8870,N_8422);
and UO_923 (O_923,N_9646,N_8607);
nor UO_924 (O_924,N_8616,N_8743);
or UO_925 (O_925,N_9806,N_8318);
nand UO_926 (O_926,N_9460,N_9135);
nand UO_927 (O_927,N_8352,N_9313);
and UO_928 (O_928,N_8428,N_8730);
xor UO_929 (O_929,N_9036,N_8123);
nor UO_930 (O_930,N_8201,N_8530);
nand UO_931 (O_931,N_9521,N_8763);
and UO_932 (O_932,N_8663,N_8419);
and UO_933 (O_933,N_8369,N_9442);
xor UO_934 (O_934,N_8901,N_9010);
and UO_935 (O_935,N_9506,N_8303);
and UO_936 (O_936,N_8697,N_8531);
and UO_937 (O_937,N_8948,N_9380);
or UO_938 (O_938,N_8682,N_8172);
xor UO_939 (O_939,N_9291,N_8880);
or UO_940 (O_940,N_9411,N_9840);
xor UO_941 (O_941,N_8295,N_8116);
nor UO_942 (O_942,N_8087,N_8665);
nand UO_943 (O_943,N_8519,N_9927);
xnor UO_944 (O_944,N_9051,N_9379);
or UO_945 (O_945,N_8093,N_8957);
and UO_946 (O_946,N_9588,N_9229);
xor UO_947 (O_947,N_9644,N_8800);
nor UO_948 (O_948,N_9534,N_8734);
nor UO_949 (O_949,N_8851,N_8195);
xor UO_950 (O_950,N_8248,N_8353);
and UO_951 (O_951,N_9936,N_9376);
nand UO_952 (O_952,N_9127,N_8987);
and UO_953 (O_953,N_8359,N_9881);
nand UO_954 (O_954,N_8953,N_9404);
xnor UO_955 (O_955,N_9926,N_9321);
nor UO_956 (O_956,N_9000,N_8895);
nor UO_957 (O_957,N_8089,N_8112);
nor UO_958 (O_958,N_9330,N_9593);
nor UO_959 (O_959,N_8460,N_9087);
xor UO_960 (O_960,N_8190,N_9758);
nor UO_961 (O_961,N_8023,N_8349);
nand UO_962 (O_962,N_9522,N_8371);
xnor UO_963 (O_963,N_9301,N_8845);
nand UO_964 (O_964,N_8914,N_9719);
nand UO_965 (O_965,N_8479,N_8549);
xnor UO_966 (O_966,N_9416,N_8780);
nand UO_967 (O_967,N_9761,N_9426);
or UO_968 (O_968,N_8062,N_9752);
and UO_969 (O_969,N_8781,N_8462);
or UO_970 (O_970,N_8030,N_8537);
xnor UO_971 (O_971,N_9123,N_8289);
nor UO_972 (O_972,N_8992,N_8051);
or UO_973 (O_973,N_9089,N_9492);
xnor UO_974 (O_974,N_9016,N_9284);
nand UO_975 (O_975,N_8642,N_8788);
nand UO_976 (O_976,N_8005,N_8774);
and UO_977 (O_977,N_9370,N_8670);
nand UO_978 (O_978,N_8411,N_8704);
nor UO_979 (O_979,N_9966,N_8455);
xnor UO_980 (O_980,N_8685,N_9381);
nand UO_981 (O_981,N_8376,N_9009);
or UO_982 (O_982,N_9075,N_8664);
nand UO_983 (O_983,N_9707,N_9623);
or UO_984 (O_984,N_9267,N_8435);
nor UO_985 (O_985,N_8494,N_8805);
xor UO_986 (O_986,N_8207,N_9023);
nor UO_987 (O_987,N_9497,N_8225);
nand UO_988 (O_988,N_9685,N_8874);
nand UO_989 (O_989,N_9186,N_8619);
nand UO_990 (O_990,N_9490,N_8792);
nor UO_991 (O_991,N_9874,N_9195);
nand UO_992 (O_992,N_9282,N_9084);
or UO_993 (O_993,N_9185,N_9366);
or UO_994 (O_994,N_9430,N_8924);
nor UO_995 (O_995,N_9309,N_8906);
or UO_996 (O_996,N_8938,N_8433);
or UO_997 (O_997,N_8072,N_9574);
nand UO_998 (O_998,N_9062,N_8075);
and UO_999 (O_999,N_8882,N_9220);
nand UO_1000 (O_1000,N_9162,N_9935);
and UO_1001 (O_1001,N_8533,N_9920);
nand UO_1002 (O_1002,N_8677,N_8456);
nand UO_1003 (O_1003,N_9514,N_9008);
or UO_1004 (O_1004,N_9884,N_9948);
or UO_1005 (O_1005,N_8731,N_8790);
and UO_1006 (O_1006,N_8640,N_9569);
or UO_1007 (O_1007,N_9905,N_8400);
nand UO_1008 (O_1008,N_8991,N_9325);
and UO_1009 (O_1009,N_8313,N_9664);
or UO_1010 (O_1010,N_8309,N_8822);
nor UO_1011 (O_1011,N_8203,N_9498);
nor UO_1012 (O_1012,N_9072,N_8035);
nand UO_1013 (O_1013,N_9232,N_8715);
and UO_1014 (O_1014,N_9959,N_8665);
or UO_1015 (O_1015,N_9913,N_8873);
nand UO_1016 (O_1016,N_8182,N_8459);
nand UO_1017 (O_1017,N_9179,N_9251);
nand UO_1018 (O_1018,N_9750,N_8600);
and UO_1019 (O_1019,N_9465,N_9421);
and UO_1020 (O_1020,N_9882,N_8071);
nand UO_1021 (O_1021,N_9146,N_9499);
nand UO_1022 (O_1022,N_9619,N_8313);
nor UO_1023 (O_1023,N_9378,N_9020);
nand UO_1024 (O_1024,N_9699,N_9275);
nand UO_1025 (O_1025,N_9340,N_9016);
and UO_1026 (O_1026,N_9558,N_9519);
and UO_1027 (O_1027,N_8803,N_8189);
or UO_1028 (O_1028,N_8203,N_8485);
xnor UO_1029 (O_1029,N_8009,N_9738);
and UO_1030 (O_1030,N_8710,N_9452);
and UO_1031 (O_1031,N_8484,N_8050);
nand UO_1032 (O_1032,N_9605,N_8522);
or UO_1033 (O_1033,N_9879,N_9813);
or UO_1034 (O_1034,N_8600,N_8060);
xor UO_1035 (O_1035,N_9216,N_9445);
nand UO_1036 (O_1036,N_9475,N_9081);
nor UO_1037 (O_1037,N_8486,N_9728);
or UO_1038 (O_1038,N_8393,N_8379);
and UO_1039 (O_1039,N_8286,N_9720);
or UO_1040 (O_1040,N_9733,N_8793);
and UO_1041 (O_1041,N_8391,N_9599);
xnor UO_1042 (O_1042,N_8143,N_8544);
nor UO_1043 (O_1043,N_8484,N_9184);
or UO_1044 (O_1044,N_8495,N_8025);
or UO_1045 (O_1045,N_8453,N_9977);
and UO_1046 (O_1046,N_8988,N_9221);
nor UO_1047 (O_1047,N_8813,N_8368);
nor UO_1048 (O_1048,N_9456,N_9955);
and UO_1049 (O_1049,N_9342,N_8196);
nor UO_1050 (O_1050,N_9110,N_9010);
or UO_1051 (O_1051,N_9821,N_9544);
and UO_1052 (O_1052,N_8554,N_9509);
nor UO_1053 (O_1053,N_9464,N_8515);
and UO_1054 (O_1054,N_9904,N_9185);
xnor UO_1055 (O_1055,N_9531,N_8881);
and UO_1056 (O_1056,N_8723,N_8453);
or UO_1057 (O_1057,N_9148,N_8986);
and UO_1058 (O_1058,N_8138,N_8036);
nor UO_1059 (O_1059,N_9578,N_9635);
nor UO_1060 (O_1060,N_8107,N_9464);
and UO_1061 (O_1061,N_8739,N_8173);
and UO_1062 (O_1062,N_8846,N_9856);
or UO_1063 (O_1063,N_8976,N_9766);
or UO_1064 (O_1064,N_9801,N_8564);
and UO_1065 (O_1065,N_8563,N_9535);
xor UO_1066 (O_1066,N_8711,N_9397);
or UO_1067 (O_1067,N_8401,N_8715);
nor UO_1068 (O_1068,N_8909,N_9992);
xor UO_1069 (O_1069,N_9359,N_9792);
and UO_1070 (O_1070,N_8393,N_9782);
and UO_1071 (O_1071,N_9550,N_9512);
and UO_1072 (O_1072,N_8927,N_8337);
nor UO_1073 (O_1073,N_8704,N_8358);
and UO_1074 (O_1074,N_9457,N_9538);
xnor UO_1075 (O_1075,N_9088,N_8467);
xnor UO_1076 (O_1076,N_8109,N_9203);
and UO_1077 (O_1077,N_9721,N_9112);
nand UO_1078 (O_1078,N_9147,N_8644);
nor UO_1079 (O_1079,N_8509,N_8514);
nand UO_1080 (O_1080,N_8754,N_9599);
and UO_1081 (O_1081,N_8526,N_9685);
nor UO_1082 (O_1082,N_9639,N_8812);
nand UO_1083 (O_1083,N_9471,N_9062);
nor UO_1084 (O_1084,N_9010,N_8712);
nor UO_1085 (O_1085,N_8904,N_9633);
or UO_1086 (O_1086,N_9795,N_9150);
nor UO_1087 (O_1087,N_9755,N_9006);
nor UO_1088 (O_1088,N_9289,N_8955);
and UO_1089 (O_1089,N_8100,N_9910);
nand UO_1090 (O_1090,N_9758,N_9517);
or UO_1091 (O_1091,N_9879,N_9920);
nand UO_1092 (O_1092,N_9067,N_8478);
nand UO_1093 (O_1093,N_8853,N_8112);
or UO_1094 (O_1094,N_8637,N_9521);
nor UO_1095 (O_1095,N_9395,N_9171);
nand UO_1096 (O_1096,N_8367,N_8885);
nand UO_1097 (O_1097,N_8627,N_9558);
and UO_1098 (O_1098,N_8906,N_9097);
nor UO_1099 (O_1099,N_8282,N_9534);
nor UO_1100 (O_1100,N_9733,N_8610);
nand UO_1101 (O_1101,N_8431,N_9741);
nand UO_1102 (O_1102,N_8819,N_9564);
or UO_1103 (O_1103,N_8520,N_8262);
and UO_1104 (O_1104,N_8817,N_8156);
nand UO_1105 (O_1105,N_9777,N_8105);
nor UO_1106 (O_1106,N_9697,N_9072);
and UO_1107 (O_1107,N_9184,N_8481);
nor UO_1108 (O_1108,N_9006,N_8641);
xor UO_1109 (O_1109,N_8108,N_9155);
nand UO_1110 (O_1110,N_8018,N_9300);
nor UO_1111 (O_1111,N_9808,N_9521);
or UO_1112 (O_1112,N_8494,N_8463);
and UO_1113 (O_1113,N_9151,N_9459);
nor UO_1114 (O_1114,N_9639,N_8499);
or UO_1115 (O_1115,N_8342,N_9598);
and UO_1116 (O_1116,N_8198,N_8604);
nand UO_1117 (O_1117,N_8142,N_8000);
or UO_1118 (O_1118,N_8936,N_9777);
and UO_1119 (O_1119,N_9812,N_9361);
or UO_1120 (O_1120,N_8116,N_9576);
or UO_1121 (O_1121,N_9567,N_8173);
nor UO_1122 (O_1122,N_8850,N_9626);
xnor UO_1123 (O_1123,N_8890,N_8146);
xnor UO_1124 (O_1124,N_9087,N_8453);
nor UO_1125 (O_1125,N_9840,N_8780);
nor UO_1126 (O_1126,N_9258,N_9352);
nor UO_1127 (O_1127,N_9851,N_9134);
or UO_1128 (O_1128,N_9872,N_8943);
and UO_1129 (O_1129,N_8498,N_9690);
and UO_1130 (O_1130,N_8580,N_8858);
nand UO_1131 (O_1131,N_9035,N_9925);
nor UO_1132 (O_1132,N_8967,N_9688);
nand UO_1133 (O_1133,N_8984,N_9013);
nand UO_1134 (O_1134,N_9777,N_8278);
nor UO_1135 (O_1135,N_9279,N_9615);
or UO_1136 (O_1136,N_9233,N_8055);
nand UO_1137 (O_1137,N_9753,N_8338);
or UO_1138 (O_1138,N_9286,N_8339);
and UO_1139 (O_1139,N_9680,N_8706);
nand UO_1140 (O_1140,N_9457,N_8381);
xnor UO_1141 (O_1141,N_9917,N_9090);
nor UO_1142 (O_1142,N_8037,N_9737);
or UO_1143 (O_1143,N_8704,N_8736);
and UO_1144 (O_1144,N_9276,N_9965);
or UO_1145 (O_1145,N_8876,N_9104);
and UO_1146 (O_1146,N_8558,N_8457);
and UO_1147 (O_1147,N_8966,N_9103);
xor UO_1148 (O_1148,N_9946,N_9931);
nor UO_1149 (O_1149,N_9421,N_8814);
or UO_1150 (O_1150,N_9217,N_9290);
or UO_1151 (O_1151,N_9376,N_8433);
nand UO_1152 (O_1152,N_8097,N_8980);
nor UO_1153 (O_1153,N_9979,N_8296);
nand UO_1154 (O_1154,N_9362,N_8657);
xor UO_1155 (O_1155,N_9043,N_9774);
or UO_1156 (O_1156,N_8894,N_9050);
and UO_1157 (O_1157,N_8957,N_8629);
nor UO_1158 (O_1158,N_8202,N_8211);
nand UO_1159 (O_1159,N_9019,N_9565);
or UO_1160 (O_1160,N_9209,N_9538);
and UO_1161 (O_1161,N_9901,N_9727);
nand UO_1162 (O_1162,N_9981,N_8141);
nand UO_1163 (O_1163,N_9366,N_8247);
or UO_1164 (O_1164,N_8482,N_8948);
and UO_1165 (O_1165,N_8898,N_9361);
nand UO_1166 (O_1166,N_8309,N_8535);
xnor UO_1167 (O_1167,N_8886,N_9027);
or UO_1168 (O_1168,N_8995,N_8899);
nand UO_1169 (O_1169,N_8252,N_8936);
or UO_1170 (O_1170,N_8036,N_8278);
nor UO_1171 (O_1171,N_8509,N_8450);
or UO_1172 (O_1172,N_8715,N_8106);
nand UO_1173 (O_1173,N_8372,N_9101);
nor UO_1174 (O_1174,N_8248,N_9776);
nor UO_1175 (O_1175,N_8828,N_9141);
and UO_1176 (O_1176,N_9112,N_9415);
nor UO_1177 (O_1177,N_9846,N_8494);
nor UO_1178 (O_1178,N_8580,N_8306);
nor UO_1179 (O_1179,N_8074,N_8807);
nor UO_1180 (O_1180,N_9103,N_9372);
nand UO_1181 (O_1181,N_9697,N_8956);
and UO_1182 (O_1182,N_8919,N_9330);
nor UO_1183 (O_1183,N_9562,N_9566);
or UO_1184 (O_1184,N_9452,N_8946);
and UO_1185 (O_1185,N_9372,N_8513);
nand UO_1186 (O_1186,N_9874,N_9955);
and UO_1187 (O_1187,N_8247,N_9454);
or UO_1188 (O_1188,N_8652,N_9009);
or UO_1189 (O_1189,N_9220,N_8831);
nor UO_1190 (O_1190,N_8715,N_9525);
nand UO_1191 (O_1191,N_9592,N_9229);
and UO_1192 (O_1192,N_9348,N_9872);
xor UO_1193 (O_1193,N_9271,N_8032);
nand UO_1194 (O_1194,N_9670,N_8999);
nand UO_1195 (O_1195,N_9053,N_8482);
nand UO_1196 (O_1196,N_9963,N_8322);
and UO_1197 (O_1197,N_8858,N_9350);
nand UO_1198 (O_1198,N_9096,N_9252);
or UO_1199 (O_1199,N_9028,N_9312);
nand UO_1200 (O_1200,N_8504,N_9397);
nand UO_1201 (O_1201,N_8043,N_9446);
or UO_1202 (O_1202,N_8628,N_9854);
and UO_1203 (O_1203,N_9291,N_9854);
or UO_1204 (O_1204,N_9408,N_9137);
and UO_1205 (O_1205,N_9664,N_8172);
or UO_1206 (O_1206,N_8477,N_9550);
and UO_1207 (O_1207,N_8480,N_9390);
nor UO_1208 (O_1208,N_9633,N_8434);
nand UO_1209 (O_1209,N_9717,N_8018);
and UO_1210 (O_1210,N_8397,N_9477);
nand UO_1211 (O_1211,N_8551,N_9734);
nor UO_1212 (O_1212,N_9899,N_8767);
and UO_1213 (O_1213,N_9161,N_9334);
and UO_1214 (O_1214,N_9554,N_8215);
and UO_1215 (O_1215,N_9918,N_9613);
nor UO_1216 (O_1216,N_9498,N_9272);
and UO_1217 (O_1217,N_9332,N_9463);
and UO_1218 (O_1218,N_8978,N_8761);
nor UO_1219 (O_1219,N_8897,N_9793);
and UO_1220 (O_1220,N_8364,N_8373);
nor UO_1221 (O_1221,N_9409,N_8961);
nor UO_1222 (O_1222,N_8259,N_9440);
and UO_1223 (O_1223,N_8153,N_8916);
and UO_1224 (O_1224,N_9496,N_8051);
xor UO_1225 (O_1225,N_9398,N_8247);
and UO_1226 (O_1226,N_9901,N_9737);
nor UO_1227 (O_1227,N_9405,N_8652);
nand UO_1228 (O_1228,N_9014,N_8085);
nor UO_1229 (O_1229,N_8707,N_8861);
or UO_1230 (O_1230,N_8204,N_9305);
or UO_1231 (O_1231,N_8300,N_8772);
nand UO_1232 (O_1232,N_9934,N_8014);
or UO_1233 (O_1233,N_8564,N_9525);
or UO_1234 (O_1234,N_9995,N_8229);
and UO_1235 (O_1235,N_9219,N_8234);
nor UO_1236 (O_1236,N_8480,N_8889);
nand UO_1237 (O_1237,N_9085,N_9371);
nor UO_1238 (O_1238,N_8972,N_9442);
nor UO_1239 (O_1239,N_9009,N_8622);
or UO_1240 (O_1240,N_9020,N_9643);
xor UO_1241 (O_1241,N_8609,N_8871);
nand UO_1242 (O_1242,N_9585,N_9198);
xor UO_1243 (O_1243,N_8108,N_9831);
nand UO_1244 (O_1244,N_8690,N_8303);
nor UO_1245 (O_1245,N_9661,N_8367);
and UO_1246 (O_1246,N_8578,N_8197);
xnor UO_1247 (O_1247,N_8640,N_8363);
or UO_1248 (O_1248,N_9602,N_8374);
and UO_1249 (O_1249,N_8769,N_8291);
and UO_1250 (O_1250,N_9146,N_9428);
xnor UO_1251 (O_1251,N_8729,N_9949);
or UO_1252 (O_1252,N_8888,N_9655);
xnor UO_1253 (O_1253,N_9219,N_8808);
and UO_1254 (O_1254,N_8268,N_9675);
or UO_1255 (O_1255,N_8806,N_8621);
and UO_1256 (O_1256,N_8352,N_9162);
and UO_1257 (O_1257,N_9694,N_8241);
and UO_1258 (O_1258,N_8466,N_9761);
nor UO_1259 (O_1259,N_9179,N_8936);
nor UO_1260 (O_1260,N_9817,N_8985);
nand UO_1261 (O_1261,N_8215,N_8040);
and UO_1262 (O_1262,N_8631,N_8649);
or UO_1263 (O_1263,N_9258,N_9106);
and UO_1264 (O_1264,N_8510,N_9401);
and UO_1265 (O_1265,N_9008,N_9466);
nor UO_1266 (O_1266,N_8164,N_9022);
nor UO_1267 (O_1267,N_9151,N_8361);
nor UO_1268 (O_1268,N_9871,N_8229);
and UO_1269 (O_1269,N_8226,N_8323);
or UO_1270 (O_1270,N_8641,N_8504);
or UO_1271 (O_1271,N_8236,N_9194);
and UO_1272 (O_1272,N_8032,N_8847);
nor UO_1273 (O_1273,N_8176,N_9479);
nand UO_1274 (O_1274,N_8680,N_8625);
xnor UO_1275 (O_1275,N_8306,N_8635);
nor UO_1276 (O_1276,N_9128,N_8263);
nand UO_1277 (O_1277,N_9738,N_9410);
and UO_1278 (O_1278,N_8138,N_9301);
or UO_1279 (O_1279,N_9358,N_9886);
nand UO_1280 (O_1280,N_8250,N_8567);
nor UO_1281 (O_1281,N_9274,N_8966);
or UO_1282 (O_1282,N_9243,N_8526);
xnor UO_1283 (O_1283,N_8999,N_8263);
and UO_1284 (O_1284,N_9673,N_8763);
nor UO_1285 (O_1285,N_9845,N_9292);
nor UO_1286 (O_1286,N_9960,N_9981);
nor UO_1287 (O_1287,N_9339,N_8890);
nand UO_1288 (O_1288,N_8618,N_8438);
or UO_1289 (O_1289,N_9785,N_9671);
and UO_1290 (O_1290,N_9631,N_9386);
nor UO_1291 (O_1291,N_9337,N_8754);
and UO_1292 (O_1292,N_8606,N_8166);
or UO_1293 (O_1293,N_9778,N_9672);
and UO_1294 (O_1294,N_8348,N_8406);
or UO_1295 (O_1295,N_9074,N_8941);
or UO_1296 (O_1296,N_8803,N_9847);
and UO_1297 (O_1297,N_8594,N_9090);
nand UO_1298 (O_1298,N_8937,N_8773);
xnor UO_1299 (O_1299,N_9620,N_8023);
nor UO_1300 (O_1300,N_9508,N_9527);
nand UO_1301 (O_1301,N_9146,N_8143);
nor UO_1302 (O_1302,N_8331,N_9147);
or UO_1303 (O_1303,N_9240,N_8027);
xor UO_1304 (O_1304,N_9826,N_8372);
nor UO_1305 (O_1305,N_9277,N_9404);
nand UO_1306 (O_1306,N_8471,N_9167);
or UO_1307 (O_1307,N_9857,N_9866);
nand UO_1308 (O_1308,N_9224,N_8388);
xor UO_1309 (O_1309,N_9131,N_9726);
and UO_1310 (O_1310,N_8857,N_9479);
nand UO_1311 (O_1311,N_8853,N_9726);
or UO_1312 (O_1312,N_8485,N_9281);
or UO_1313 (O_1313,N_8044,N_9614);
and UO_1314 (O_1314,N_9380,N_8989);
nand UO_1315 (O_1315,N_9551,N_8016);
xnor UO_1316 (O_1316,N_8456,N_8079);
nor UO_1317 (O_1317,N_8442,N_9139);
xor UO_1318 (O_1318,N_8497,N_9489);
and UO_1319 (O_1319,N_9594,N_8246);
nand UO_1320 (O_1320,N_9300,N_8776);
xor UO_1321 (O_1321,N_9261,N_9697);
nand UO_1322 (O_1322,N_9786,N_9366);
and UO_1323 (O_1323,N_8449,N_8445);
nand UO_1324 (O_1324,N_8216,N_9764);
and UO_1325 (O_1325,N_8159,N_9254);
xor UO_1326 (O_1326,N_8770,N_9147);
xor UO_1327 (O_1327,N_9051,N_8047);
or UO_1328 (O_1328,N_8262,N_8625);
nor UO_1329 (O_1329,N_8922,N_8813);
or UO_1330 (O_1330,N_9387,N_9782);
nor UO_1331 (O_1331,N_9140,N_8884);
and UO_1332 (O_1332,N_9704,N_9539);
and UO_1333 (O_1333,N_9199,N_9391);
or UO_1334 (O_1334,N_8282,N_8381);
nand UO_1335 (O_1335,N_8711,N_9032);
nor UO_1336 (O_1336,N_9572,N_8916);
and UO_1337 (O_1337,N_8086,N_8140);
xor UO_1338 (O_1338,N_8119,N_8238);
and UO_1339 (O_1339,N_8176,N_8066);
nor UO_1340 (O_1340,N_8375,N_9457);
nor UO_1341 (O_1341,N_8259,N_8014);
and UO_1342 (O_1342,N_9651,N_9990);
nand UO_1343 (O_1343,N_8143,N_9982);
or UO_1344 (O_1344,N_8196,N_9551);
nor UO_1345 (O_1345,N_9409,N_8004);
nand UO_1346 (O_1346,N_9398,N_9184);
nand UO_1347 (O_1347,N_8954,N_8096);
xor UO_1348 (O_1348,N_8097,N_9559);
or UO_1349 (O_1349,N_8444,N_9532);
or UO_1350 (O_1350,N_8845,N_9212);
or UO_1351 (O_1351,N_9267,N_9804);
or UO_1352 (O_1352,N_9662,N_9797);
or UO_1353 (O_1353,N_8482,N_8248);
nor UO_1354 (O_1354,N_8668,N_8318);
or UO_1355 (O_1355,N_9215,N_8189);
or UO_1356 (O_1356,N_8232,N_9063);
nor UO_1357 (O_1357,N_9705,N_9487);
or UO_1358 (O_1358,N_9098,N_9902);
and UO_1359 (O_1359,N_9717,N_9490);
nand UO_1360 (O_1360,N_9476,N_9792);
xor UO_1361 (O_1361,N_8445,N_9676);
or UO_1362 (O_1362,N_9578,N_8172);
xor UO_1363 (O_1363,N_9321,N_9788);
and UO_1364 (O_1364,N_9110,N_8853);
nand UO_1365 (O_1365,N_8439,N_9403);
nand UO_1366 (O_1366,N_9207,N_8898);
or UO_1367 (O_1367,N_8185,N_8293);
and UO_1368 (O_1368,N_8465,N_8099);
nor UO_1369 (O_1369,N_9220,N_9650);
or UO_1370 (O_1370,N_9981,N_9651);
and UO_1371 (O_1371,N_8742,N_8754);
xnor UO_1372 (O_1372,N_8519,N_8676);
or UO_1373 (O_1373,N_9371,N_9943);
nand UO_1374 (O_1374,N_9905,N_9045);
nor UO_1375 (O_1375,N_9603,N_9430);
and UO_1376 (O_1376,N_8876,N_9385);
or UO_1377 (O_1377,N_9243,N_9121);
xnor UO_1378 (O_1378,N_9902,N_9716);
and UO_1379 (O_1379,N_9318,N_9226);
or UO_1380 (O_1380,N_9720,N_9366);
nor UO_1381 (O_1381,N_9437,N_9945);
and UO_1382 (O_1382,N_8821,N_8959);
xnor UO_1383 (O_1383,N_8128,N_9338);
xnor UO_1384 (O_1384,N_8245,N_8268);
xor UO_1385 (O_1385,N_8818,N_9024);
and UO_1386 (O_1386,N_8674,N_9994);
nor UO_1387 (O_1387,N_8180,N_8358);
nand UO_1388 (O_1388,N_9084,N_8332);
and UO_1389 (O_1389,N_9780,N_8477);
xor UO_1390 (O_1390,N_8704,N_8799);
nor UO_1391 (O_1391,N_9611,N_8421);
or UO_1392 (O_1392,N_8739,N_9591);
or UO_1393 (O_1393,N_9338,N_8263);
or UO_1394 (O_1394,N_9909,N_8042);
and UO_1395 (O_1395,N_8018,N_9882);
nor UO_1396 (O_1396,N_9307,N_9915);
nor UO_1397 (O_1397,N_9128,N_9536);
nand UO_1398 (O_1398,N_8257,N_8615);
or UO_1399 (O_1399,N_9111,N_9945);
nand UO_1400 (O_1400,N_8562,N_9354);
and UO_1401 (O_1401,N_9769,N_8234);
and UO_1402 (O_1402,N_8241,N_9002);
nand UO_1403 (O_1403,N_8761,N_9621);
and UO_1404 (O_1404,N_9130,N_8813);
xor UO_1405 (O_1405,N_8448,N_9082);
xnor UO_1406 (O_1406,N_9739,N_8369);
nand UO_1407 (O_1407,N_8474,N_8430);
nand UO_1408 (O_1408,N_9093,N_9166);
nand UO_1409 (O_1409,N_8606,N_8020);
nor UO_1410 (O_1410,N_9631,N_9195);
and UO_1411 (O_1411,N_9789,N_9216);
and UO_1412 (O_1412,N_8084,N_9317);
or UO_1413 (O_1413,N_8235,N_8612);
xor UO_1414 (O_1414,N_9563,N_8975);
and UO_1415 (O_1415,N_8469,N_9949);
nor UO_1416 (O_1416,N_9556,N_8002);
or UO_1417 (O_1417,N_8077,N_9279);
nand UO_1418 (O_1418,N_9678,N_8029);
nor UO_1419 (O_1419,N_9085,N_8197);
xor UO_1420 (O_1420,N_9552,N_8361);
nand UO_1421 (O_1421,N_9812,N_8688);
and UO_1422 (O_1422,N_8306,N_9003);
nand UO_1423 (O_1423,N_8554,N_8030);
nor UO_1424 (O_1424,N_8712,N_8975);
nand UO_1425 (O_1425,N_9541,N_9771);
and UO_1426 (O_1426,N_8828,N_9740);
and UO_1427 (O_1427,N_8632,N_9008);
nand UO_1428 (O_1428,N_9260,N_8832);
or UO_1429 (O_1429,N_8082,N_8016);
xor UO_1430 (O_1430,N_8287,N_8554);
or UO_1431 (O_1431,N_9021,N_9166);
or UO_1432 (O_1432,N_8350,N_8931);
nor UO_1433 (O_1433,N_9527,N_9883);
xor UO_1434 (O_1434,N_9599,N_8969);
nor UO_1435 (O_1435,N_9941,N_8192);
or UO_1436 (O_1436,N_8276,N_9482);
and UO_1437 (O_1437,N_8806,N_8812);
nand UO_1438 (O_1438,N_8351,N_8684);
or UO_1439 (O_1439,N_9151,N_8681);
nand UO_1440 (O_1440,N_8774,N_9367);
or UO_1441 (O_1441,N_8477,N_9026);
or UO_1442 (O_1442,N_8128,N_8097);
xor UO_1443 (O_1443,N_9744,N_9111);
nor UO_1444 (O_1444,N_8292,N_8149);
xor UO_1445 (O_1445,N_8420,N_9804);
and UO_1446 (O_1446,N_8816,N_8180);
or UO_1447 (O_1447,N_9474,N_8380);
nor UO_1448 (O_1448,N_8626,N_9300);
and UO_1449 (O_1449,N_8150,N_9217);
or UO_1450 (O_1450,N_9795,N_9459);
nor UO_1451 (O_1451,N_8530,N_9547);
or UO_1452 (O_1452,N_9536,N_9596);
or UO_1453 (O_1453,N_9412,N_9064);
or UO_1454 (O_1454,N_8428,N_8456);
or UO_1455 (O_1455,N_9770,N_9700);
xor UO_1456 (O_1456,N_8027,N_9743);
nand UO_1457 (O_1457,N_9047,N_9728);
nand UO_1458 (O_1458,N_8163,N_8851);
xnor UO_1459 (O_1459,N_9691,N_8508);
or UO_1460 (O_1460,N_8682,N_9459);
nor UO_1461 (O_1461,N_8726,N_8857);
and UO_1462 (O_1462,N_9630,N_8050);
or UO_1463 (O_1463,N_9472,N_9055);
nand UO_1464 (O_1464,N_8033,N_8140);
nand UO_1465 (O_1465,N_9206,N_8485);
nand UO_1466 (O_1466,N_9030,N_9698);
nor UO_1467 (O_1467,N_9168,N_9734);
and UO_1468 (O_1468,N_9868,N_8534);
nand UO_1469 (O_1469,N_8602,N_9434);
xor UO_1470 (O_1470,N_8228,N_9054);
and UO_1471 (O_1471,N_9797,N_9389);
xor UO_1472 (O_1472,N_9587,N_9383);
and UO_1473 (O_1473,N_9715,N_8802);
and UO_1474 (O_1474,N_8422,N_8737);
and UO_1475 (O_1475,N_9987,N_9030);
nand UO_1476 (O_1476,N_8484,N_8235);
nor UO_1477 (O_1477,N_9170,N_8507);
or UO_1478 (O_1478,N_8393,N_8422);
nor UO_1479 (O_1479,N_8889,N_8114);
or UO_1480 (O_1480,N_9848,N_9782);
nand UO_1481 (O_1481,N_8683,N_8121);
or UO_1482 (O_1482,N_8004,N_8881);
and UO_1483 (O_1483,N_8509,N_9887);
nor UO_1484 (O_1484,N_8398,N_8473);
or UO_1485 (O_1485,N_9924,N_8290);
nand UO_1486 (O_1486,N_8826,N_8090);
nand UO_1487 (O_1487,N_9457,N_9655);
or UO_1488 (O_1488,N_8532,N_9420);
and UO_1489 (O_1489,N_8899,N_8887);
nor UO_1490 (O_1490,N_9281,N_8265);
nand UO_1491 (O_1491,N_8677,N_8740);
nor UO_1492 (O_1492,N_8669,N_9951);
nor UO_1493 (O_1493,N_8038,N_8641);
nand UO_1494 (O_1494,N_8836,N_9092);
and UO_1495 (O_1495,N_8948,N_8919);
or UO_1496 (O_1496,N_8716,N_9862);
and UO_1497 (O_1497,N_9387,N_9391);
nor UO_1498 (O_1498,N_9837,N_8897);
and UO_1499 (O_1499,N_9778,N_9355);
endmodule