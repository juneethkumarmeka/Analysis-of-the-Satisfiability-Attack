module basic_2000_20000_2500_10_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_1142,In_537);
nor U1 (N_1,In_370,In_445);
nor U2 (N_2,In_1789,In_940);
nand U3 (N_3,In_1116,In_1562);
nand U4 (N_4,In_76,In_1798);
or U5 (N_5,In_1145,In_1107);
nor U6 (N_6,In_507,In_1729);
nand U7 (N_7,In_184,In_413);
xnor U8 (N_8,In_63,In_1169);
or U9 (N_9,In_1243,In_1673);
nand U10 (N_10,In_22,In_15);
nor U11 (N_11,In_23,In_1576);
nand U12 (N_12,In_577,In_788);
nand U13 (N_13,In_885,In_1981);
nor U14 (N_14,In_828,In_1944);
and U15 (N_15,In_1234,In_648);
or U16 (N_16,In_1248,In_688);
nand U17 (N_17,In_402,In_1830);
nand U18 (N_18,In_1083,In_1856);
nand U19 (N_19,In_1113,In_1996);
or U20 (N_20,In_221,In_1613);
or U21 (N_21,In_1115,In_781);
or U22 (N_22,In_349,In_1974);
and U23 (N_23,In_1217,In_1547);
nand U24 (N_24,In_409,In_837);
or U25 (N_25,In_544,In_1386);
nand U26 (N_26,In_1311,In_1004);
or U27 (N_27,In_567,In_1967);
or U28 (N_28,In_1126,In_549);
nand U29 (N_29,In_1552,In_1690);
nand U30 (N_30,In_1771,In_405);
nand U31 (N_31,In_1134,In_473);
xor U32 (N_32,In_821,In_1708);
nor U33 (N_33,In_794,In_1803);
or U34 (N_34,In_1833,In_469);
nand U35 (N_35,In_1725,In_1574);
and U36 (N_36,In_765,In_1881);
and U37 (N_37,In_1223,In_1170);
or U38 (N_38,In_1760,In_457);
or U39 (N_39,In_386,In_213);
and U40 (N_40,In_241,In_1139);
nor U41 (N_41,In_1808,In_981);
and U42 (N_42,In_1596,In_206);
or U43 (N_43,In_1215,In_1431);
nor U44 (N_44,In_724,In_123);
nor U45 (N_45,In_927,In_466);
and U46 (N_46,In_508,In_107);
or U47 (N_47,In_1817,In_1794);
xor U48 (N_48,In_894,In_1230);
xnor U49 (N_49,In_211,In_246);
or U50 (N_50,In_1173,In_1767);
and U51 (N_51,In_1618,In_879);
or U52 (N_52,In_436,In_1517);
and U53 (N_53,In_1800,In_1988);
nor U54 (N_54,In_515,In_566);
and U55 (N_55,In_564,In_547);
nor U56 (N_56,In_1986,In_275);
xor U57 (N_57,In_1713,In_1327);
and U58 (N_58,In_1128,In_430);
nand U59 (N_59,In_408,In_527);
xor U60 (N_60,In_1138,In_923);
or U61 (N_61,In_570,In_795);
and U62 (N_62,In_1978,In_546);
and U63 (N_63,In_480,In_873);
nor U64 (N_64,In_1249,In_932);
or U65 (N_65,In_1916,In_590);
or U66 (N_66,In_960,In_889);
or U67 (N_67,In_139,In_563);
xnor U68 (N_68,In_956,In_155);
nand U69 (N_69,In_704,In_832);
or U70 (N_70,In_202,In_843);
nand U71 (N_71,In_1163,In_91);
and U72 (N_72,In_49,In_1922);
or U73 (N_73,In_1034,In_1802);
xnor U74 (N_74,In_170,In_360);
nor U75 (N_75,In_805,In_1356);
nor U76 (N_76,In_521,In_1861);
nand U77 (N_77,In_841,In_38);
nand U78 (N_78,In_189,In_809);
or U79 (N_79,In_703,In_630);
or U80 (N_80,In_1518,In_1480);
nand U81 (N_81,In_1899,In_1666);
or U82 (N_82,In_1033,In_1401);
and U83 (N_83,In_1943,In_1603);
or U84 (N_84,In_1396,In_207);
or U85 (N_85,In_1866,In_493);
or U86 (N_86,In_341,In_631);
or U87 (N_87,In_1114,In_1970);
and U88 (N_88,In_1739,In_1393);
xnor U89 (N_89,In_254,In_69);
and U90 (N_90,In_818,In_118);
or U91 (N_91,In_1864,In_893);
and U92 (N_92,In_1041,In_398);
nand U93 (N_93,In_20,In_1872);
and U94 (N_94,In_1687,In_1140);
or U95 (N_95,In_1316,In_1254);
nand U96 (N_96,In_1869,In_133);
nand U97 (N_97,In_1056,In_1620);
nor U98 (N_98,In_1512,In_1601);
and U99 (N_99,In_293,In_0);
or U100 (N_100,In_387,In_1065);
nor U101 (N_101,In_1422,In_1913);
or U102 (N_102,In_611,In_56);
or U103 (N_103,In_1067,In_1928);
nand U104 (N_104,In_231,In_1099);
or U105 (N_105,In_1879,In_1372);
and U106 (N_106,In_150,In_1871);
nor U107 (N_107,In_448,In_1473);
nand U108 (N_108,In_1077,In_1556);
nand U109 (N_109,In_1962,In_1726);
nor U110 (N_110,In_793,In_1595);
xnor U111 (N_111,In_1733,In_1615);
nor U112 (N_112,In_1362,In_1822);
nor U113 (N_113,In_1651,In_1717);
or U114 (N_114,In_756,In_1721);
and U115 (N_115,In_926,In_1037);
and U116 (N_116,In_947,In_532);
and U117 (N_117,In_462,In_997);
and U118 (N_118,In_1886,In_1098);
nor U119 (N_119,In_806,In_778);
and U120 (N_120,In_464,In_1937);
or U121 (N_121,In_220,In_1882);
xnor U122 (N_122,In_509,In_198);
and U123 (N_123,In_830,In_602);
nor U124 (N_124,In_1838,In_1627);
nand U125 (N_125,In_318,In_1488);
xor U126 (N_126,In_10,In_367);
and U127 (N_127,In_256,In_880);
and U128 (N_128,In_1549,In_576);
nand U129 (N_129,In_1617,In_1847);
nand U130 (N_130,In_753,In_1266);
nand U131 (N_131,In_574,In_538);
nor U132 (N_132,In_734,In_375);
xnor U133 (N_133,In_957,In_1848);
and U134 (N_134,In_979,In_768);
nand U135 (N_135,In_1697,In_731);
nor U136 (N_136,In_287,In_657);
or U137 (N_137,In_135,In_366);
xnor U138 (N_138,In_1199,In_776);
or U139 (N_139,In_808,In_1481);
nor U140 (N_140,In_1700,In_862);
or U141 (N_141,In_34,In_1436);
and U142 (N_142,In_1742,In_264);
nor U143 (N_143,In_1049,In_742);
and U144 (N_144,In_1060,In_180);
xor U145 (N_145,In_1971,In_815);
or U146 (N_146,In_1514,In_160);
and U147 (N_147,In_481,In_319);
and U148 (N_148,In_482,In_288);
nand U149 (N_149,In_849,In_1323);
and U150 (N_150,In_1374,In_1949);
nand U151 (N_151,In_686,In_1942);
or U152 (N_152,In_959,In_1588);
or U153 (N_153,In_1398,In_513);
xnor U154 (N_154,In_489,In_1051);
nor U155 (N_155,In_449,In_1806);
xor U156 (N_156,In_892,In_1644);
nand U157 (N_157,In_741,In_1277);
nor U158 (N_158,In_320,In_477);
and U159 (N_159,In_1196,In_1357);
and U160 (N_160,In_1634,In_487);
nor U161 (N_161,In_332,In_311);
and U162 (N_162,In_1855,In_1703);
nand U163 (N_163,In_1082,In_1337);
nand U164 (N_164,In_1095,In_266);
or U165 (N_165,In_260,In_154);
and U166 (N_166,In_1598,In_388);
nor U167 (N_167,In_1453,In_1889);
xnor U168 (N_168,In_1509,In_476);
or U169 (N_169,In_665,In_1179);
and U170 (N_170,In_1508,In_215);
nor U171 (N_171,In_581,In_1397);
or U172 (N_172,In_1332,In_1648);
and U173 (N_173,In_798,In_1288);
and U174 (N_174,In_573,In_333);
nor U175 (N_175,In_569,In_1313);
nand U176 (N_176,In_1043,In_1247);
xnor U177 (N_177,In_970,In_1911);
and U178 (N_178,In_512,In_1446);
or U179 (N_179,In_958,In_1735);
nor U180 (N_180,In_774,In_1710);
nand U181 (N_181,In_1074,In_829);
or U182 (N_182,In_132,In_996);
and U183 (N_183,In_586,In_1171);
and U184 (N_184,In_1207,In_1705);
and U185 (N_185,In_371,In_804);
nor U186 (N_186,In_1,In_352);
nor U187 (N_187,In_823,In_588);
xor U188 (N_188,In_751,In_1786);
nor U189 (N_189,In_1209,In_1555);
or U190 (N_190,In_906,In_346);
nor U191 (N_191,In_1376,In_1801);
nor U192 (N_192,In_802,In_551);
and U193 (N_193,In_441,In_623);
or U194 (N_194,In_1302,In_390);
xnor U195 (N_195,In_622,In_1945);
and U196 (N_196,In_1961,In_1137);
or U197 (N_197,In_975,In_833);
nor U198 (N_198,In_933,In_624);
xor U199 (N_199,In_166,In_1053);
and U200 (N_200,In_1746,In_230);
nand U201 (N_201,In_204,In_236);
nand U202 (N_202,In_1764,In_1857);
nor U203 (N_203,In_1274,In_1289);
nand U204 (N_204,In_603,In_1669);
or U205 (N_205,In_1533,In_1476);
and U206 (N_206,In_1605,In_257);
nand U207 (N_207,In_866,In_1519);
nor U208 (N_208,In_506,In_1842);
and U209 (N_209,In_1185,In_1216);
nand U210 (N_210,In_1989,In_1459);
and U211 (N_211,In_1444,In_278);
and U212 (N_212,In_1371,In_416);
nor U213 (N_213,In_785,In_1271);
nor U214 (N_214,In_99,In_1968);
nand U215 (N_215,In_1600,In_522);
nor U216 (N_216,In_1607,In_791);
or U217 (N_217,In_330,In_758);
nor U218 (N_218,In_867,In_79);
nand U219 (N_219,In_1110,In_877);
and U220 (N_220,In_787,In_819);
nand U221 (N_221,In_1692,In_1888);
or U222 (N_222,In_16,In_813);
or U223 (N_223,In_1977,In_1273);
nor U224 (N_224,In_1366,In_1759);
nand U225 (N_225,In_1660,In_297);
nor U226 (N_226,In_357,In_1959);
nor U227 (N_227,In_18,In_1351);
xnor U228 (N_228,In_1003,In_676);
nand U229 (N_229,In_1305,In_219);
nand U230 (N_230,In_993,In_659);
nor U231 (N_231,In_317,In_1483);
nor U232 (N_232,In_1863,In_424);
nor U233 (N_233,In_1293,In_411);
and U234 (N_234,In_895,In_1360);
nor U235 (N_235,In_1463,In_228);
and U236 (N_236,In_255,In_1284);
or U237 (N_237,In_604,In_1706);
or U238 (N_238,In_391,In_212);
nand U239 (N_239,In_437,In_1883);
nand U240 (N_240,In_498,In_519);
and U241 (N_241,In_1845,In_1427);
or U242 (N_242,In_1958,In_1251);
or U243 (N_243,In_1934,In_1526);
xor U244 (N_244,In_1245,In_1191);
or U245 (N_245,In_775,In_651);
nor U246 (N_246,In_948,In_31);
nand U247 (N_247,In_931,In_1407);
and U248 (N_248,In_682,In_1778);
nor U249 (N_249,In_1220,In_1825);
nand U250 (N_250,In_1720,In_605);
nand U251 (N_251,In_966,In_1162);
xor U252 (N_252,In_347,In_552);
nand U253 (N_253,In_542,In_1870);
and U254 (N_254,In_985,In_848);
xor U255 (N_255,In_510,In_355);
nor U256 (N_256,In_921,In_760);
or U257 (N_257,In_1550,In_772);
and U258 (N_258,In_859,In_524);
nor U259 (N_259,In_1278,In_1581);
xor U260 (N_260,In_1557,In_262);
xnor U261 (N_261,In_1221,In_1619);
nand U262 (N_262,In_746,In_1773);
nor U263 (N_263,In_1670,In_593);
nor U264 (N_264,In_1963,In_1513);
and U265 (N_265,In_92,In_1527);
xor U266 (N_266,In_263,In_650);
nand U267 (N_267,In_301,In_138);
or U268 (N_268,In_1662,In_591);
nor U269 (N_269,In_1008,In_1814);
or U270 (N_270,In_1984,In_1202);
or U271 (N_271,In_1136,In_1242);
nor U272 (N_272,In_426,In_1631);
nand U273 (N_273,In_952,In_125);
and U274 (N_274,In_835,In_223);
nor U275 (N_275,In_7,In_702);
nor U276 (N_276,In_1681,In_846);
nor U277 (N_277,In_51,In_354);
nand U278 (N_278,In_1100,In_1679);
xnor U279 (N_279,In_726,In_656);
and U280 (N_280,In_141,In_857);
nand U281 (N_281,In_1568,In_816);
and U282 (N_282,In_1440,In_73);
nand U283 (N_283,In_639,In_109);
and U284 (N_284,In_1540,In_632);
and U285 (N_285,In_1317,In_66);
nor U286 (N_286,In_192,In_693);
nand U287 (N_287,In_748,In_1496);
nor U288 (N_288,In_851,In_157);
nand U289 (N_289,In_1719,In_766);
nand U290 (N_290,In_1409,In_1792);
or U291 (N_291,In_1754,In_1022);
nor U292 (N_292,In_1902,In_899);
xor U293 (N_293,In_488,In_446);
and U294 (N_294,In_1415,In_1458);
and U295 (N_295,In_345,In_976);
nor U296 (N_296,In_111,In_1707);
and U297 (N_297,In_227,In_978);
and U298 (N_298,In_1728,In_226);
nor U299 (N_299,In_1405,In_1938);
and U300 (N_300,In_484,In_280);
nor U301 (N_301,In_70,In_147);
nor U302 (N_302,In_394,In_727);
and U303 (N_303,In_474,In_61);
or U304 (N_304,In_638,In_1625);
or U305 (N_305,In_801,In_1907);
or U306 (N_306,In_839,In_304);
nand U307 (N_307,In_1059,In_356);
nand U308 (N_308,In_1072,In_1569);
or U309 (N_309,In_1105,In_1960);
or U310 (N_310,In_483,In_78);
nand U311 (N_311,In_729,In_1419);
and U312 (N_312,In_1106,In_516);
nor U313 (N_313,In_875,In_30);
nor U314 (N_314,In_1103,In_1628);
xor U315 (N_315,In_41,In_903);
and U316 (N_316,In_383,In_1516);
or U317 (N_317,In_1029,In_1319);
and U318 (N_318,In_222,In_46);
and U319 (N_319,In_271,In_52);
or U320 (N_320,In_1894,In_181);
or U321 (N_321,In_1127,In_1312);
nor U322 (N_322,In_913,In_1521);
nor U323 (N_323,In_208,In_1553);
or U324 (N_324,In_812,In_607);
or U325 (N_325,In_1616,In_1014);
or U326 (N_326,In_1388,In_1612);
xor U327 (N_327,In_1811,In_919);
nand U328 (N_328,In_585,In_1632);
xnor U329 (N_329,In_533,In_578);
and U330 (N_330,In_444,In_990);
and U331 (N_331,In_967,In_269);
or U332 (N_332,In_615,In_1195);
and U333 (N_333,In_158,In_1040);
nor U334 (N_334,In_410,In_1515);
nor U335 (N_335,In_1111,In_415);
nor U336 (N_336,In_1447,In_856);
nor U337 (N_337,In_1490,In_545);
and U338 (N_338,In_1346,In_238);
nor U339 (N_339,In_869,In_1834);
or U340 (N_340,In_1867,In_824);
xnor U341 (N_341,In_143,In_401);
nor U342 (N_342,In_757,In_438);
nor U343 (N_343,In_1722,In_541);
and U344 (N_344,In_1455,In_1176);
and U345 (N_345,In_479,In_1186);
and U346 (N_346,In_486,In_321);
nand U347 (N_347,In_1239,In_1523);
nand U348 (N_348,In_635,In_1671);
nand U349 (N_349,In_247,In_331);
nand U350 (N_350,In_1123,In_1015);
nor U351 (N_351,In_217,In_1365);
or U352 (N_352,In_1865,In_177);
xor U353 (N_353,In_1751,In_190);
or U354 (N_354,In_348,In_252);
or U355 (N_355,In_1743,In_1203);
nor U356 (N_356,In_1304,In_1437);
nor U357 (N_357,In_1572,In_1953);
nor U358 (N_358,In_420,In_689);
and U359 (N_359,In_322,In_1183);
and U360 (N_360,In_1506,In_472);
nor U361 (N_361,In_200,In_800);
nand U362 (N_362,In_55,In_1164);
nand U363 (N_363,In_1931,In_43);
nor U364 (N_364,In_443,In_531);
nor U365 (N_365,In_1210,In_596);
and U366 (N_366,In_303,In_945);
xnor U367 (N_367,In_1375,In_1255);
nand U368 (N_368,In_467,In_1682);
nor U369 (N_369,In_1484,In_917);
nand U370 (N_370,In_1655,In_675);
and U371 (N_371,In_1414,In_1536);
or U372 (N_372,In_244,In_232);
nor U373 (N_373,In_911,In_674);
and U374 (N_374,In_253,In_1227);
nand U375 (N_375,In_1604,In_397);
or U376 (N_376,In_1844,In_429);
nand U377 (N_377,In_660,In_182);
nor U378 (N_378,In_1235,In_1429);
or U379 (N_379,In_442,In_571);
and U380 (N_380,In_980,In_1500);
or U381 (N_381,In_503,In_172);
nor U382 (N_382,In_1658,In_277);
xnor U383 (N_383,In_1464,In_754);
nand U384 (N_384,In_1683,In_1290);
and U385 (N_385,In_767,In_1636);
nor U386 (N_386,In_1434,In_1920);
nor U387 (N_387,In_684,In_1783);
and U388 (N_388,In_68,In_250);
nor U389 (N_389,In_176,In_962);
nor U390 (N_390,In_619,In_562);
xnor U391 (N_391,In_210,In_86);
nor U392 (N_392,In_1734,In_306);
nor U393 (N_393,In_161,In_421);
nor U394 (N_394,In_381,In_1472);
or U395 (N_395,In_1718,In_1776);
and U396 (N_396,In_1025,In_245);
and U397 (N_397,In_965,In_939);
and U398 (N_398,In_1471,In_1565);
nor U399 (N_399,In_1505,In_1795);
nand U400 (N_400,In_989,In_435);
and U401 (N_401,In_1545,In_1238);
or U402 (N_402,In_1264,In_1309);
xor U403 (N_403,In_81,In_834);
nor U404 (N_404,In_718,In_613);
nand U405 (N_405,In_173,In_1350);
and U406 (N_406,In_716,In_1796);
and U407 (N_407,In_1878,In_1112);
nor U408 (N_408,In_162,In_925);
and U409 (N_409,In_553,In_1924);
and U410 (N_410,In_1478,In_900);
nand U411 (N_411,In_74,In_382);
and U412 (N_412,In_362,In_1686);
nor U413 (N_413,In_706,In_598);
or U414 (N_414,In_1387,In_1339);
nor U415 (N_415,In_852,In_1543);
nand U416 (N_416,In_104,In_550);
nor U417 (N_417,In_1016,In_643);
or U418 (N_418,In_499,In_954);
nor U419 (N_419,In_117,In_1983);
xnor U420 (N_420,In_750,In_1267);
nor U421 (N_421,In_1846,In_1222);
nor U422 (N_422,In_1246,In_1390);
nor U423 (N_423,In_928,In_59);
or U424 (N_424,In_314,In_1840);
nor U425 (N_425,In_1167,In_1900);
xnor U426 (N_426,In_50,In_1813);
and U427 (N_427,In_24,In_1300);
nor U428 (N_428,In_1843,In_1353);
nand U429 (N_429,In_929,In_579);
or U430 (N_430,In_140,In_789);
or U431 (N_431,In_1404,In_1629);
nand U432 (N_432,In_597,In_1301);
nor U433 (N_433,In_1769,In_1129);
and U434 (N_434,In_276,In_1815);
nand U435 (N_435,In_175,In_1999);
nor U436 (N_436,In_407,In_1086);
and U437 (N_437,In_1424,In_174);
nand U438 (N_438,In_1544,In_62);
nand U439 (N_439,In_1919,In_580);
and U440 (N_440,In_1124,In_1837);
nand U441 (N_441,In_243,In_283);
nand U442 (N_442,In_12,In_872);
and U443 (N_443,In_518,In_1542);
or U444 (N_444,In_1590,In_1088);
nor U445 (N_445,In_431,In_1741);
and U446 (N_446,In_973,In_1213);
or U447 (N_447,In_440,In_1154);
or U448 (N_448,In_1499,In_1197);
nand U449 (N_449,In_1336,In_1228);
nor U450 (N_450,In_1768,In_1208);
nand U451 (N_451,In_1297,In_491);
nand U452 (N_452,In_1024,In_1954);
and U453 (N_453,In_1281,In_1320);
or U454 (N_454,In_1812,In_769);
and U455 (N_455,In_621,In_1606);
nand U456 (N_456,In_1036,In_1435);
nand U457 (N_457,In_1699,In_216);
xnor U458 (N_458,In_1250,In_1367);
or U459 (N_459,In_1253,In_1647);
or U460 (N_460,In_1343,In_1380);
nand U461 (N_461,In_1150,In_119);
nor U462 (N_462,In_1344,In_1325);
and U463 (N_463,In_629,In_884);
and U464 (N_464,In_677,In_1985);
nor U465 (N_465,In_137,In_194);
or U466 (N_466,In_455,In_836);
or U467 (N_467,In_1157,In_1640);
and U468 (N_468,In_1394,In_273);
and U469 (N_469,In_136,In_1772);
and U470 (N_470,In_764,In_1042);
xnor U471 (N_471,In_1633,In_972);
or U472 (N_472,In_27,In_738);
nor U473 (N_473,In_1175,In_1130);
xor U474 (N_474,In_425,In_529);
nand U475 (N_475,In_705,In_151);
nand U476 (N_476,In_1045,In_797);
nand U477 (N_477,In_186,In_1448);
nand U478 (N_478,In_35,In_1212);
or U479 (N_479,In_1001,In_1586);
or U480 (N_480,In_1987,In_1205);
or U481 (N_481,In_338,In_1991);
and U482 (N_482,In_1724,In_1198);
nand U483 (N_483,In_1310,In_886);
nand U484 (N_484,In_1694,In_1020);
or U485 (N_485,In_1936,In_1952);
and U486 (N_486,In_1933,In_21);
and U487 (N_487,In_548,In_199);
nor U488 (N_488,In_1915,In_1452);
and U489 (N_489,In_633,In_1068);
or U490 (N_490,In_1652,In_1108);
nand U491 (N_491,In_1119,In_1649);
nor U492 (N_492,In_1094,In_658);
or U493 (N_493,In_1460,In_1416);
xnor U494 (N_494,In_337,In_1432);
nand U495 (N_495,In_359,In_326);
and U496 (N_496,In_1487,In_1237);
or U497 (N_497,In_1836,In_114);
nand U498 (N_498,In_384,In_1408);
and U499 (N_499,In_825,In_53);
or U500 (N_500,In_1240,In_1530);
and U501 (N_501,In_864,In_620);
or U502 (N_502,In_1973,In_1260);
and U503 (N_503,In_908,In_1069);
nand U504 (N_504,In_1348,In_910);
nor U505 (N_505,In_999,In_1592);
xnor U506 (N_506,In_33,In_1835);
nand U507 (N_507,In_1950,In_1093);
xor U508 (N_508,In_1873,In_450);
and U509 (N_509,In_1610,In_1653);
xor U510 (N_510,In_1957,In_1283);
or U511 (N_511,In_1012,In_363);
nor U512 (N_512,In_195,In_1331);
or U513 (N_513,In_930,In_148);
nor U514 (N_514,In_747,In_955);
nand U515 (N_515,In_1685,In_1091);
nor U516 (N_516,In_14,In_646);
and U517 (N_517,In_1090,In_1850);
xnor U518 (N_518,In_1645,In_1622);
and U519 (N_519,In_1926,In_142);
nand U520 (N_520,In_1969,In_1218);
nor U521 (N_521,In_1046,In_419);
or U522 (N_522,In_1770,In_740);
nand U523 (N_523,In_242,In_1972);
nand U524 (N_524,In_286,In_1839);
xor U525 (N_525,In_1927,In_1187);
nor U526 (N_526,In_640,In_1828);
and U527 (N_527,In_1951,In_124);
nor U528 (N_528,In_942,In_1998);
and U529 (N_529,In_423,In_1159);
and U530 (N_530,In_389,In_1745);
or U531 (N_531,In_1280,In_485);
nand U532 (N_532,In_1307,In_1548);
and U533 (N_533,In_1704,In_1038);
xnor U534 (N_534,In_514,In_329);
xnor U535 (N_535,In_1275,In_471);
or U536 (N_536,In_75,In_951);
or U537 (N_537,In_912,In_1165);
or U538 (N_538,In_439,In_248);
xnor U539 (N_539,In_490,In_1906);
nor U540 (N_540,In_1876,In_977);
or U541 (N_541,In_1747,In_568);
nand U542 (N_542,In_1563,In_1827);
xor U543 (N_543,In_504,In_618);
and U544 (N_544,In_625,In_1994);
and U545 (N_545,In_1383,In_90);
or U546 (N_546,In_628,In_302);
nor U547 (N_547,In_1057,In_755);
nand U548 (N_548,In_1062,In_1497);
and U549 (N_549,In_540,In_358);
nor U550 (N_550,In_492,In_600);
or U551 (N_551,In_905,In_372);
xnor U552 (N_552,In_453,In_272);
or U553 (N_553,In_1941,In_1976);
and U554 (N_554,In_871,In_720);
nand U555 (N_555,In_1917,In_984);
nand U556 (N_556,In_696,In_265);
or U557 (N_557,In_898,In_47);
or U558 (N_558,In_1539,In_1832);
and U559 (N_559,In_1912,In_1370);
nor U560 (N_560,In_163,In_698);
and U561 (N_561,In_1143,In_82);
nand U562 (N_562,In_1964,In_1005);
nand U563 (N_563,In_1373,In_992);
nand U564 (N_564,In_460,In_1177);
nand U565 (N_565,In_1898,In_1711);
nor U566 (N_566,In_907,In_1314);
and U567 (N_567,In_669,In_465);
nor U568 (N_568,In_1761,In_103);
nand U569 (N_569,In_205,In_1558);
xnor U570 (N_570,In_1474,In_1829);
or U571 (N_571,In_1443,In_1740);
or U572 (N_572,In_281,In_134);
nand U573 (N_573,In_1184,In_188);
nor U574 (N_574,In_295,In_1048);
or U575 (N_575,In_711,In_1265);
or U576 (N_576,In_3,In_868);
nor U577 (N_577,In_105,In_447);
and U578 (N_578,In_1492,In_1564);
and U579 (N_579,In_1862,In_1858);
nand U580 (N_580,In_102,In_122);
nor U581 (N_581,In_773,In_847);
nand U582 (N_582,In_152,In_652);
xor U583 (N_583,In_1676,In_1790);
or U584 (N_584,In_100,In_1433);
or U585 (N_585,In_32,In_739);
and U586 (N_586,In_1997,In_1623);
and U587 (N_587,In_936,In_1120);
and U588 (N_588,In_1391,In_279);
and U589 (N_589,In_1626,In_77);
nor U590 (N_590,In_1322,In_1677);
and U591 (N_591,In_112,In_1630);
nand U592 (N_592,In_685,In_560);
nand U593 (N_593,In_1507,In_1744);
and U594 (N_594,In_865,In_1279);
nor U595 (N_595,In_239,In_183);
or U596 (N_596,In_1347,In_1342);
nor U597 (N_597,In_803,In_203);
xor U598 (N_598,In_1334,In_1172);
xor U599 (N_599,In_725,In_1193);
xor U600 (N_600,In_1716,In_1571);
nand U601 (N_601,In_1285,In_1381);
or U602 (N_602,In_1392,In_1295);
and U603 (N_603,In_149,In_1738);
nand U604 (N_604,In_916,In_106);
nor U605 (N_605,In_1578,In_666);
or U606 (N_606,In_855,In_1809);
and U607 (N_607,In_1287,In_1665);
nand U608 (N_608,In_369,In_1691);
or U609 (N_609,In_1058,In_1299);
and U610 (N_610,In_458,In_379);
nand U611 (N_611,In_1256,In_282);
and U612 (N_612,In_1097,In_328);
and U613 (N_613,In_1663,In_762);
and U614 (N_614,In_904,In_575);
nor U615 (N_615,In_608,In_1621);
nand U616 (N_616,In_1732,In_572);
or U617 (N_617,In_1750,In_452);
and U618 (N_618,In_393,In_1990);
or U619 (N_619,In_454,In_759);
or U620 (N_620,In_983,In_475);
or U621 (N_621,In_994,In_1063);
xnor U622 (N_622,In_101,In_1897);
and U623 (N_623,In_1583,In_1573);
nor U624 (N_624,In_128,In_1182);
nand U625 (N_625,In_1905,In_418);
nor U626 (N_626,In_683,In_1292);
or U627 (N_627,In_502,In_897);
nor U628 (N_628,In_1748,In_1430);
or U629 (N_629,In_1493,In_191);
or U630 (N_630,In_310,In_644);
or U631 (N_631,In_673,In_1262);
xnor U632 (N_632,In_1580,In_1081);
and U633 (N_633,In_780,In_969);
nand U634 (N_634,In_1233,In_316);
and U635 (N_635,In_1089,In_1007);
nor U636 (N_636,In_350,In_1980);
xnor U637 (N_637,In_918,In_964);
and U638 (N_638,In_58,In_1276);
xnor U639 (N_639,In_1194,In_376);
and U640 (N_640,In_422,In_1155);
nand U641 (N_641,In_1715,In_662);
and U642 (N_642,In_1657,In_1765);
and U643 (N_643,In_922,In_378);
or U644 (N_644,In_324,In_1402);
xnor U645 (N_645,In_1087,In_1465);
nand U646 (N_646,In_159,In_953);
nor U647 (N_647,In_67,In_1667);
nor U648 (N_648,In_730,In_1575);
or U649 (N_649,In_1259,In_505);
and U650 (N_650,In_209,In_783);
nor U651 (N_651,In_1914,In_1698);
and U652 (N_652,In_882,In_1192);
nand U653 (N_653,In_240,In_1675);
and U654 (N_654,In_771,In_1328);
nor U655 (N_655,In_399,In_478);
or U656 (N_656,In_1642,In_1009);
and U657 (N_657,In_126,In_1047);
or U658 (N_658,In_1384,In_661);
and U659 (N_659,In_285,In_97);
or U660 (N_660,In_268,In_810);
or U661 (N_661,In_1799,In_888);
and U662 (N_662,In_1158,In_1469);
xnor U663 (N_663,In_1560,In_763);
nor U664 (N_664,In_156,In_1702);
nor U665 (N_665,In_395,In_1345);
and U666 (N_666,In_299,In_1611);
nand U667 (N_667,In_1537,In_1026);
and U668 (N_668,In_5,In_1252);
nor U669 (N_669,In_1161,In_1076);
or U670 (N_670,In_543,In_1477);
or U671 (N_671,In_1468,In_1650);
and U672 (N_672,In_1286,In_949);
and U673 (N_673,In_377,In_1948);
nor U674 (N_674,In_1055,In_728);
and U675 (N_675,In_1000,In_1204);
nand U676 (N_676,In_334,In_1723);
and U677 (N_677,In_1002,In_305);
and U678 (N_678,In_1896,In_1224);
nand U679 (N_679,In_1805,In_556);
or U680 (N_680,In_1166,In_1554);
or U681 (N_681,In_1294,In_627);
xnor U682 (N_682,In_887,In_1413);
xor U683 (N_683,In_653,In_594);
nand U684 (N_684,In_1714,In_1132);
or U685 (N_685,In_692,In_672);
or U686 (N_686,In_6,In_1661);
nor U687 (N_687,In_790,In_1385);
nand U688 (N_688,In_1885,In_1080);
xor U689 (N_689,In_1831,In_1475);
nor U690 (N_690,In_1895,In_1824);
xor U691 (N_691,In_1947,In_1017);
nor U692 (N_692,In_432,In_1052);
nor U693 (N_693,In_1489,In_1449);
nand U694 (N_694,In_129,In_616);
or U695 (N_695,In_878,In_1774);
or U696 (N_696,In_289,In_1762);
nand U697 (N_697,In_64,In_1466);
nand U698 (N_698,In_365,In_461);
and U699 (N_699,In_792,In_463);
or U700 (N_700,In_844,In_93);
xor U701 (N_701,In_637,In_1073);
and U702 (N_702,In_1780,In_168);
nor U703 (N_703,In_820,In_1775);
nand U704 (N_704,In_249,In_599);
or U705 (N_705,In_1891,In_1382);
or U706 (N_706,In_1538,In_1498);
nor U707 (N_707,In_1643,In_863);
nand U708 (N_708,In_1141,In_595);
nand U709 (N_709,In_339,In_434);
nand U710 (N_710,In_11,In_1330);
or U711 (N_711,In_169,In_1071);
nand U712 (N_712,In_617,In_1229);
or U713 (N_713,In_1785,In_1693);
nand U714 (N_714,In_1303,In_1178);
or U715 (N_715,In_83,In_1363);
nand U716 (N_716,In_1624,In_987);
or U717 (N_717,In_251,In_934);
and U718 (N_718,In_883,In_1324);
nor U719 (N_719,In_1078,In_54);
nand U720 (N_720,In_1638,In_1456);
nor U721 (N_721,In_745,In_327);
nor U722 (N_722,In_668,In_1333);
or U723 (N_723,In_343,In_1504);
xor U724 (N_724,In_699,In_1755);
nand U725 (N_725,In_1349,In_1131);
nor U726 (N_726,In_937,In_1445);
nor U727 (N_727,In_1486,In_1841);
or U728 (N_728,In_1160,In_1757);
or U729 (N_729,In_1758,In_782);
nand U730 (N_730,In_396,In_717);
nor U731 (N_731,In_694,In_1032);
xor U732 (N_732,In_1491,In_526);
nand U733 (N_733,In_144,In_986);
nor U734 (N_734,In_353,In_1122);
and U735 (N_735,In_891,In_995);
nand U736 (N_736,In_941,In_1125);
nor U737 (N_737,In_1591,In_667);
nand U738 (N_738,In_1709,In_1501);
nor U739 (N_739,In_1689,In_1462);
nand U740 (N_740,In_850,In_690);
nor U741 (N_741,In_1935,In_1901);
nor U742 (N_742,In_373,In_1296);
nand U743 (N_743,In_1566,In_645);
and U744 (N_744,In_1656,In_1854);
nor U745 (N_745,In_583,In_946);
or U746 (N_746,In_1411,In_1594);
xnor U747 (N_747,In_874,In_1109);
nand U748 (N_748,In_1599,In_1674);
xor U749 (N_749,In_584,In_193);
or U750 (N_750,In_1884,In_1261);
and U751 (N_751,In_722,In_1511);
or U752 (N_752,In_44,In_695);
nand U753 (N_753,In_1039,In_1368);
xor U754 (N_754,In_414,In_292);
nand U755 (N_755,In_1727,In_225);
or U756 (N_756,In_1975,In_364);
nor U757 (N_757,In_1326,In_909);
nor U758 (N_758,In_1030,In_565);
and U759 (N_759,In_1318,In_914);
or U760 (N_760,In_1932,In_1752);
or U761 (N_761,In_121,In_284);
nor U762 (N_762,In_1144,In_497);
or U763 (N_763,In_308,In_25);
and U764 (N_764,In_636,In_1925);
nand U765 (N_765,In_1439,In_1852);
nand U766 (N_766,In_1420,In_1421);
and U767 (N_767,In_670,In_1940);
nand U768 (N_768,In_146,In_1135);
or U769 (N_769,In_1096,In_323);
nor U770 (N_770,In_1352,In_737);
and U771 (N_771,In_36,In_374);
and U772 (N_772,In_1639,In_920);
nor U773 (N_773,In_42,In_88);
or U774 (N_774,In_968,In_587);
and U775 (N_775,In_96,In_340);
nor U776 (N_776,In_13,In_822);
nor U777 (N_777,In_1567,In_1244);
nand U778 (N_778,In_335,In_626);
and U779 (N_779,In_1979,In_845);
nand U780 (N_780,In_520,In_1641);
nand U781 (N_781,In_1791,In_974);
and U782 (N_782,In_1749,In_368);
and U783 (N_783,In_267,In_57);
and U784 (N_784,In_1225,In_201);
nand U785 (N_785,In_1593,In_433);
and U786 (N_786,In_1956,In_1696);
nor U787 (N_787,In_678,In_164);
nor U788 (N_788,In_1880,In_752);
or U789 (N_789,In_85,In_1156);
and U790 (N_790,In_679,In_1579);
or U791 (N_791,In_511,In_1084);
nand U792 (N_792,In_1369,In_1023);
and U793 (N_793,In_1736,In_1389);
nor U794 (N_794,In_235,In_403);
nor U795 (N_795,In_680,In_1887);
nor U796 (N_796,In_1232,In_1993);
xnor U797 (N_797,In_1546,In_344);
nand U798 (N_798,In_218,In_1399);
and U799 (N_799,In_45,In_902);
and U800 (N_800,In_1438,In_1892);
and U801 (N_801,In_171,In_1903);
or U802 (N_802,In_649,In_558);
nor U803 (N_803,In_296,In_890);
and U804 (N_804,In_259,In_701);
nor U805 (N_805,In_1502,In_1263);
xor U806 (N_806,In_642,In_1495);
and U807 (N_807,In_715,In_1298);
and U808 (N_808,In_1201,In_1646);
nor U809 (N_809,In_1403,In_404);
nand U810 (N_810,In_1226,In_1609);
and U811 (N_811,In_1470,In_1152);
nor U812 (N_812,In_39,In_1359);
nand U813 (N_813,In_1753,In_1664);
nand U814 (N_814,In_1451,In_517);
xor U815 (N_815,In_733,In_1321);
nor U816 (N_816,In_1121,In_1180);
and U817 (N_817,In_307,In_1035);
and U818 (N_818,In_1361,In_108);
and U819 (N_819,In_707,In_400);
or U820 (N_820,In_1788,In_915);
and U821 (N_821,In_1777,In_89);
nor U822 (N_822,In_1019,In_1853);
nand U823 (N_823,In_1766,In_853);
xor U824 (N_824,In_539,In_1146);
and U825 (N_825,In_351,In_807);
nor U826 (N_826,In_1737,In_1955);
xnor U827 (N_827,In_1211,In_1425);
xor U828 (N_828,In_961,In_258);
nand U829 (N_829,In_601,In_315);
nand U830 (N_830,In_1781,In_614);
and U831 (N_831,In_1849,In_153);
xor U832 (N_832,In_1821,In_536);
nor U833 (N_833,In_1485,In_664);
xor U834 (N_834,In_528,In_1890);
and U835 (N_835,In_224,In_291);
and U836 (N_836,In_1148,In_523);
xor U837 (N_837,In_1206,In_1582);
or U838 (N_838,In_736,In_495);
nor U839 (N_839,In_270,In_827);
or U840 (N_840,In_1104,In_1441);
and U841 (N_841,In_1482,In_606);
xnor U842 (N_842,In_131,In_1027);
xor U843 (N_843,In_971,In_525);
xnor U844 (N_844,In_708,In_1939);
or U845 (N_845,In_456,In_557);
nand U846 (N_846,In_1860,In_1561);
nand U847 (N_847,In_1730,In_1188);
xor U848 (N_848,In_1587,In_943);
or U849 (N_849,In_641,In_655);
nor U850 (N_850,In_1329,In_1010);
or U851 (N_851,In_1021,In_838);
or U852 (N_852,In_1904,In_1678);
or U853 (N_853,In_761,In_924);
nand U854 (N_854,In_392,In_1826);
nand U855 (N_855,In_697,In_988);
nand U856 (N_856,In_1355,In_998);
nand U857 (N_857,In_500,In_1461);
or U858 (N_858,In_589,In_1820);
nor U859 (N_859,In_380,In_1412);
nor U860 (N_860,In_609,In_1423);
nand U861 (N_861,In_1153,In_1364);
nor U862 (N_862,In_713,In_1308);
and U863 (N_863,In_1918,In_1102);
xor U864 (N_864,In_1525,In_799);
nor U865 (N_865,In_385,In_26);
or U866 (N_866,In_1011,In_1426);
and U867 (N_867,In_779,In_1241);
xnor U868 (N_868,In_944,In_1529);
xnor U869 (N_869,In_687,In_95);
or U870 (N_870,In_796,In_40);
and U871 (N_871,In_1528,In_127);
nand U872 (N_872,In_1868,In_325);
nor U873 (N_873,In_37,In_860);
xor U874 (N_874,In_417,In_1340);
or U875 (N_875,In_1921,In_1117);
nand U876 (N_876,In_935,In_28);
xnor U877 (N_877,In_1494,In_831);
nand U878 (N_878,In_671,In_361);
nor U879 (N_879,In_17,In_1680);
and U880 (N_880,In_1819,In_950);
or U881 (N_881,In_1965,In_1908);
and U882 (N_882,In_826,In_1189);
and U883 (N_883,In_876,In_1875);
and U884 (N_884,In_1450,In_691);
nand U885 (N_885,In_1797,In_1075);
or U886 (N_886,In_309,In_709);
nor U887 (N_887,In_817,In_1442);
nand U888 (N_888,In_1522,In_786);
or U889 (N_889,In_1577,In_858);
nand U890 (N_890,In_19,In_165);
or U891 (N_891,In_938,In_428);
or U892 (N_892,In_861,In_120);
or U893 (N_893,In_459,In_881);
and U894 (N_894,In_1909,In_1608);
nand U895 (N_895,In_29,In_1395);
nand U896 (N_896,In_1282,In_274);
or U897 (N_897,In_229,In_814);
nand U898 (N_898,In_1804,In_451);
nor U899 (N_899,In_9,In_197);
or U900 (N_900,In_1174,In_1712);
nor U901 (N_901,In_714,In_298);
nand U902 (N_902,In_1923,In_261);
and U903 (N_903,In_1028,In_1354);
and U904 (N_904,In_1779,In_1756);
xor U905 (N_905,In_749,In_1379);
and U906 (N_906,In_1272,In_1066);
nor U907 (N_907,In_1701,In_1101);
nand U908 (N_908,In_1672,In_1085);
and U909 (N_909,In_654,In_610);
or U910 (N_910,In_854,In_412);
and U911 (N_911,In_700,In_561);
and U912 (N_912,In_1637,In_896);
nor U913 (N_913,In_1092,In_1534);
nor U914 (N_914,In_145,In_1535);
nand U915 (N_915,In_1231,In_294);
or U916 (N_916,In_113,In_1874);
and U917 (N_917,In_1457,In_991);
or U918 (N_918,In_1147,In_1654);
nand U919 (N_919,In_98,In_1410);
nand U920 (N_920,In_179,In_1763);
nor U921 (N_921,In_300,In_501);
xor U922 (N_922,In_1214,In_94);
nand U923 (N_923,In_470,In_494);
nor U924 (N_924,In_8,In_901);
and U925 (N_925,In_1269,In_237);
xnor U926 (N_926,In_535,In_1291);
or U927 (N_927,In_1149,In_1064);
and U928 (N_928,In_110,In_1597);
and U929 (N_929,In_65,In_1338);
xor U930 (N_930,In_4,In_80);
nor U931 (N_931,In_1570,In_719);
nor U932 (N_932,In_1044,In_1151);
xor U933 (N_933,In_313,In_982);
or U934 (N_934,In_634,In_592);
and U935 (N_935,In_1695,In_1510);
or U936 (N_936,In_712,In_178);
nand U937 (N_937,In_744,In_1315);
or U938 (N_938,In_681,In_1503);
nor U939 (N_939,In_1454,In_1524);
nor U940 (N_940,In_1782,In_1614);
and U941 (N_941,In_1585,In_1018);
nor U942 (N_942,In_1406,In_721);
or U943 (N_943,In_732,In_842);
and U944 (N_944,In_84,In_1378);
or U945 (N_945,In_1992,In_1910);
nor U946 (N_946,In_1731,In_710);
and U947 (N_947,In_167,In_1930);
and U948 (N_948,In_1181,In_555);
nor U949 (N_949,In_1358,In_647);
xnor U950 (N_950,In_743,In_116);
nand U951 (N_951,In_1417,In_1995);
xor U952 (N_952,In_196,In_1467);
nand U953 (N_953,In_1133,In_1688);
and U954 (N_954,In_1877,In_1541);
and U955 (N_955,In_840,In_1418);
nor U956 (N_956,In_1584,In_1793);
nand U957 (N_957,In_1635,In_1168);
and U958 (N_958,In_870,In_1851);
and U959 (N_959,In_1270,In_233);
and U960 (N_960,In_1659,In_1551);
nor U961 (N_961,In_1070,In_1668);
nand U962 (N_962,In_1946,In_1784);
or U963 (N_963,In_1532,In_1982);
and U964 (N_964,In_777,In_1559);
nor U965 (N_965,In_1816,In_1013);
or U966 (N_966,In_1520,In_87);
and U967 (N_967,In_554,In_1257);
and U968 (N_968,In_187,In_1236);
and U969 (N_969,In_1190,In_1810);
nor U970 (N_970,In_1268,In_1079);
nor U971 (N_971,In_811,In_1823);
nand U972 (N_972,In_1479,In_115);
xor U973 (N_973,In_1929,In_530);
nor U974 (N_974,In_342,In_663);
or U975 (N_975,In_1818,In_1054);
nand U976 (N_976,In_185,In_2);
xnor U977 (N_977,In_1859,In_963);
and U978 (N_978,In_1966,In_1219);
and U979 (N_979,In_130,In_1684);
nand U980 (N_980,In_735,In_1531);
nand U981 (N_981,In_582,In_1341);
nor U982 (N_982,In_1602,In_336);
nor U983 (N_983,In_406,In_214);
and U984 (N_984,In_468,In_71);
nand U985 (N_985,In_784,In_1400);
xnor U986 (N_986,In_723,In_1306);
nor U987 (N_987,In_427,In_60);
nand U988 (N_988,In_48,In_1050);
or U989 (N_989,In_1061,In_559);
nor U990 (N_990,In_534,In_1335);
or U991 (N_991,In_72,In_1428);
or U992 (N_992,In_1031,In_312);
nand U993 (N_993,In_1807,In_1589);
nand U994 (N_994,In_1787,In_612);
and U995 (N_995,In_496,In_1200);
and U996 (N_996,In_290,In_1893);
nand U997 (N_997,In_1377,In_770);
or U998 (N_998,In_234,In_1118);
or U999 (N_999,In_1006,In_1258);
and U1000 (N_1000,In_1037,In_863);
and U1001 (N_1001,In_78,In_1659);
nand U1002 (N_1002,In_1134,In_663);
and U1003 (N_1003,In_690,In_1202);
nand U1004 (N_1004,In_903,In_244);
or U1005 (N_1005,In_460,In_394);
and U1006 (N_1006,In_1164,In_1334);
nand U1007 (N_1007,In_1280,In_987);
nor U1008 (N_1008,In_1554,In_247);
xnor U1009 (N_1009,In_840,In_1358);
nand U1010 (N_1010,In_492,In_143);
nand U1011 (N_1011,In_258,In_1308);
or U1012 (N_1012,In_101,In_1472);
or U1013 (N_1013,In_1428,In_498);
nor U1014 (N_1014,In_227,In_304);
and U1015 (N_1015,In_1767,In_67);
and U1016 (N_1016,In_1827,In_1063);
and U1017 (N_1017,In_77,In_2);
xor U1018 (N_1018,In_187,In_25);
and U1019 (N_1019,In_127,In_794);
nand U1020 (N_1020,In_998,In_1262);
nand U1021 (N_1021,In_1353,In_147);
nand U1022 (N_1022,In_1118,In_1868);
nand U1023 (N_1023,In_1737,In_1319);
nor U1024 (N_1024,In_164,In_1661);
or U1025 (N_1025,In_21,In_1758);
and U1026 (N_1026,In_1153,In_826);
or U1027 (N_1027,In_176,In_125);
xnor U1028 (N_1028,In_1003,In_1149);
nor U1029 (N_1029,In_1600,In_1732);
xnor U1030 (N_1030,In_1024,In_164);
or U1031 (N_1031,In_473,In_494);
or U1032 (N_1032,In_1416,In_1497);
or U1033 (N_1033,In_771,In_500);
or U1034 (N_1034,In_1091,In_585);
nand U1035 (N_1035,In_514,In_1419);
and U1036 (N_1036,In_1374,In_1463);
and U1037 (N_1037,In_15,In_1212);
and U1038 (N_1038,In_341,In_174);
nor U1039 (N_1039,In_1775,In_326);
and U1040 (N_1040,In_786,In_179);
or U1041 (N_1041,In_1408,In_822);
nand U1042 (N_1042,In_1218,In_685);
nor U1043 (N_1043,In_529,In_1267);
and U1044 (N_1044,In_1570,In_1836);
or U1045 (N_1045,In_702,In_984);
or U1046 (N_1046,In_703,In_1375);
or U1047 (N_1047,In_654,In_302);
nor U1048 (N_1048,In_89,In_421);
or U1049 (N_1049,In_948,In_1399);
nor U1050 (N_1050,In_1137,In_1622);
nor U1051 (N_1051,In_1081,In_996);
nor U1052 (N_1052,In_1147,In_1368);
nor U1053 (N_1053,In_694,In_1324);
nand U1054 (N_1054,In_1112,In_80);
and U1055 (N_1055,In_468,In_1233);
nand U1056 (N_1056,In_320,In_1578);
nand U1057 (N_1057,In_1085,In_1117);
and U1058 (N_1058,In_1901,In_265);
nor U1059 (N_1059,In_101,In_678);
or U1060 (N_1060,In_1879,In_4);
nand U1061 (N_1061,In_532,In_1966);
and U1062 (N_1062,In_905,In_672);
or U1063 (N_1063,In_281,In_733);
nand U1064 (N_1064,In_1582,In_357);
nand U1065 (N_1065,In_1809,In_111);
nor U1066 (N_1066,In_458,In_1331);
and U1067 (N_1067,In_169,In_1255);
or U1068 (N_1068,In_793,In_71);
xnor U1069 (N_1069,In_50,In_144);
xor U1070 (N_1070,In_1486,In_1952);
nand U1071 (N_1071,In_1120,In_95);
and U1072 (N_1072,In_1565,In_1086);
and U1073 (N_1073,In_366,In_849);
and U1074 (N_1074,In_1617,In_635);
or U1075 (N_1075,In_1410,In_1917);
nor U1076 (N_1076,In_1891,In_1736);
or U1077 (N_1077,In_182,In_160);
nand U1078 (N_1078,In_1648,In_1409);
and U1079 (N_1079,In_422,In_512);
or U1080 (N_1080,In_284,In_208);
and U1081 (N_1081,In_1245,In_485);
or U1082 (N_1082,In_1001,In_839);
nor U1083 (N_1083,In_737,In_517);
nand U1084 (N_1084,In_1995,In_432);
nor U1085 (N_1085,In_584,In_145);
nor U1086 (N_1086,In_1264,In_845);
xor U1087 (N_1087,In_1528,In_1761);
nor U1088 (N_1088,In_1036,In_1266);
xor U1089 (N_1089,In_1318,In_935);
xor U1090 (N_1090,In_1577,In_1011);
xor U1091 (N_1091,In_1506,In_1673);
xor U1092 (N_1092,In_283,In_1900);
nand U1093 (N_1093,In_1743,In_1867);
and U1094 (N_1094,In_319,In_52);
nand U1095 (N_1095,In_1731,In_673);
nand U1096 (N_1096,In_635,In_575);
and U1097 (N_1097,In_255,In_578);
nor U1098 (N_1098,In_1002,In_802);
and U1099 (N_1099,In_1163,In_329);
nand U1100 (N_1100,In_554,In_1718);
or U1101 (N_1101,In_1514,In_92);
nor U1102 (N_1102,In_659,In_1783);
or U1103 (N_1103,In_468,In_661);
or U1104 (N_1104,In_121,In_1650);
nand U1105 (N_1105,In_829,In_1028);
and U1106 (N_1106,In_144,In_898);
xor U1107 (N_1107,In_511,In_816);
nand U1108 (N_1108,In_263,In_1052);
and U1109 (N_1109,In_323,In_1944);
xnor U1110 (N_1110,In_106,In_47);
nand U1111 (N_1111,In_319,In_1321);
nand U1112 (N_1112,In_92,In_1350);
or U1113 (N_1113,In_1623,In_400);
nor U1114 (N_1114,In_677,In_285);
nand U1115 (N_1115,In_372,In_52);
and U1116 (N_1116,In_778,In_1149);
and U1117 (N_1117,In_145,In_941);
nand U1118 (N_1118,In_640,In_1043);
and U1119 (N_1119,In_1964,In_12);
and U1120 (N_1120,In_292,In_106);
xnor U1121 (N_1121,In_1160,In_1827);
and U1122 (N_1122,In_1455,In_1892);
nand U1123 (N_1123,In_1764,In_1695);
xnor U1124 (N_1124,In_1058,In_1729);
and U1125 (N_1125,In_722,In_338);
and U1126 (N_1126,In_1970,In_614);
and U1127 (N_1127,In_793,In_1182);
nor U1128 (N_1128,In_479,In_1086);
nor U1129 (N_1129,In_1698,In_165);
nor U1130 (N_1130,In_921,In_1919);
nor U1131 (N_1131,In_1006,In_304);
or U1132 (N_1132,In_1316,In_947);
or U1133 (N_1133,In_75,In_384);
nor U1134 (N_1134,In_434,In_879);
nand U1135 (N_1135,In_59,In_1308);
nand U1136 (N_1136,In_516,In_537);
nand U1137 (N_1137,In_1920,In_303);
nand U1138 (N_1138,In_1608,In_120);
or U1139 (N_1139,In_1539,In_1394);
nand U1140 (N_1140,In_184,In_1493);
nand U1141 (N_1141,In_1436,In_807);
and U1142 (N_1142,In_182,In_1958);
nor U1143 (N_1143,In_692,In_173);
or U1144 (N_1144,In_635,In_66);
nor U1145 (N_1145,In_1728,In_189);
nor U1146 (N_1146,In_565,In_1964);
nor U1147 (N_1147,In_364,In_1615);
or U1148 (N_1148,In_1114,In_1890);
xnor U1149 (N_1149,In_345,In_1284);
nand U1150 (N_1150,In_1191,In_1404);
xor U1151 (N_1151,In_842,In_468);
nor U1152 (N_1152,In_136,In_1420);
nor U1153 (N_1153,In_153,In_1974);
nand U1154 (N_1154,In_1568,In_1099);
nor U1155 (N_1155,In_546,In_1834);
nor U1156 (N_1156,In_368,In_1855);
nor U1157 (N_1157,In_334,In_66);
or U1158 (N_1158,In_342,In_141);
or U1159 (N_1159,In_61,In_1437);
nor U1160 (N_1160,In_1909,In_223);
or U1161 (N_1161,In_1526,In_855);
nand U1162 (N_1162,In_1528,In_1827);
nor U1163 (N_1163,In_1442,In_1588);
nand U1164 (N_1164,In_1379,In_1245);
and U1165 (N_1165,In_238,In_1192);
and U1166 (N_1166,In_463,In_242);
nor U1167 (N_1167,In_474,In_534);
and U1168 (N_1168,In_1570,In_936);
nand U1169 (N_1169,In_1411,In_1972);
and U1170 (N_1170,In_336,In_295);
and U1171 (N_1171,In_604,In_212);
or U1172 (N_1172,In_1782,In_1376);
or U1173 (N_1173,In_116,In_779);
nor U1174 (N_1174,In_1225,In_1744);
nand U1175 (N_1175,In_595,In_1296);
or U1176 (N_1176,In_261,In_586);
nand U1177 (N_1177,In_1110,In_1157);
nor U1178 (N_1178,In_583,In_1922);
xnor U1179 (N_1179,In_1757,In_701);
and U1180 (N_1180,In_457,In_751);
or U1181 (N_1181,In_1648,In_1507);
or U1182 (N_1182,In_1935,In_1790);
or U1183 (N_1183,In_1510,In_1219);
or U1184 (N_1184,In_313,In_1343);
nor U1185 (N_1185,In_1833,In_1121);
nor U1186 (N_1186,In_321,In_596);
nand U1187 (N_1187,In_1192,In_915);
or U1188 (N_1188,In_831,In_136);
nand U1189 (N_1189,In_836,In_565);
and U1190 (N_1190,In_1565,In_360);
and U1191 (N_1191,In_1855,In_974);
and U1192 (N_1192,In_801,In_382);
and U1193 (N_1193,In_1541,In_994);
or U1194 (N_1194,In_1915,In_1801);
nand U1195 (N_1195,In_1219,In_391);
or U1196 (N_1196,In_1694,In_1124);
or U1197 (N_1197,In_57,In_889);
and U1198 (N_1198,In_1418,In_1602);
or U1199 (N_1199,In_1295,In_248);
and U1200 (N_1200,In_927,In_1304);
and U1201 (N_1201,In_969,In_1485);
nand U1202 (N_1202,In_437,In_1281);
and U1203 (N_1203,In_679,In_53);
nor U1204 (N_1204,In_1533,In_174);
or U1205 (N_1205,In_1196,In_1277);
or U1206 (N_1206,In_1314,In_537);
nand U1207 (N_1207,In_1436,In_1965);
xnor U1208 (N_1208,In_1915,In_620);
and U1209 (N_1209,In_92,In_1513);
and U1210 (N_1210,In_485,In_226);
nor U1211 (N_1211,In_125,In_264);
or U1212 (N_1212,In_1754,In_538);
nor U1213 (N_1213,In_650,In_1622);
nor U1214 (N_1214,In_1266,In_1466);
nor U1215 (N_1215,In_1331,In_172);
nor U1216 (N_1216,In_1636,In_375);
or U1217 (N_1217,In_1106,In_1283);
or U1218 (N_1218,In_658,In_42);
or U1219 (N_1219,In_606,In_16);
and U1220 (N_1220,In_316,In_1291);
xor U1221 (N_1221,In_1216,In_713);
nand U1222 (N_1222,In_465,In_1757);
and U1223 (N_1223,In_745,In_1456);
or U1224 (N_1224,In_1593,In_1095);
or U1225 (N_1225,In_811,In_1710);
nor U1226 (N_1226,In_627,In_292);
and U1227 (N_1227,In_475,In_224);
or U1228 (N_1228,In_1864,In_1848);
or U1229 (N_1229,In_505,In_664);
nor U1230 (N_1230,In_1713,In_1770);
nor U1231 (N_1231,In_1337,In_357);
nand U1232 (N_1232,In_1330,In_606);
and U1233 (N_1233,In_1556,In_1051);
nor U1234 (N_1234,In_413,In_1589);
and U1235 (N_1235,In_1805,In_630);
nand U1236 (N_1236,In_1185,In_917);
xor U1237 (N_1237,In_1275,In_1109);
or U1238 (N_1238,In_1994,In_142);
or U1239 (N_1239,In_524,In_1032);
and U1240 (N_1240,In_1755,In_534);
nor U1241 (N_1241,In_923,In_1833);
nand U1242 (N_1242,In_469,In_1736);
or U1243 (N_1243,In_1779,In_1672);
or U1244 (N_1244,In_1893,In_1264);
or U1245 (N_1245,In_347,In_50);
nor U1246 (N_1246,In_344,In_678);
or U1247 (N_1247,In_1866,In_1755);
or U1248 (N_1248,In_73,In_1628);
nor U1249 (N_1249,In_710,In_298);
nand U1250 (N_1250,In_858,In_1750);
nor U1251 (N_1251,In_293,In_382);
and U1252 (N_1252,In_1154,In_1311);
xnor U1253 (N_1253,In_1894,In_1058);
and U1254 (N_1254,In_1722,In_1495);
or U1255 (N_1255,In_1090,In_77);
nor U1256 (N_1256,In_340,In_876);
or U1257 (N_1257,In_1318,In_1918);
and U1258 (N_1258,In_1683,In_861);
or U1259 (N_1259,In_1492,In_465);
or U1260 (N_1260,In_1552,In_812);
xnor U1261 (N_1261,In_1398,In_1901);
nor U1262 (N_1262,In_907,In_1174);
and U1263 (N_1263,In_647,In_1899);
nand U1264 (N_1264,In_1568,In_143);
xnor U1265 (N_1265,In_588,In_407);
or U1266 (N_1266,In_1894,In_723);
nor U1267 (N_1267,In_910,In_22);
or U1268 (N_1268,In_1610,In_378);
and U1269 (N_1269,In_34,In_1193);
nor U1270 (N_1270,In_1637,In_613);
nor U1271 (N_1271,In_1062,In_644);
nand U1272 (N_1272,In_1849,In_105);
and U1273 (N_1273,In_70,In_1407);
or U1274 (N_1274,In_123,In_1703);
or U1275 (N_1275,In_931,In_1582);
and U1276 (N_1276,In_664,In_606);
or U1277 (N_1277,In_749,In_1988);
and U1278 (N_1278,In_822,In_811);
nand U1279 (N_1279,In_1023,In_98);
and U1280 (N_1280,In_1113,In_1471);
or U1281 (N_1281,In_721,In_596);
nand U1282 (N_1282,In_31,In_1660);
nor U1283 (N_1283,In_1699,In_1744);
xor U1284 (N_1284,In_107,In_1030);
or U1285 (N_1285,In_1927,In_491);
or U1286 (N_1286,In_451,In_1895);
nor U1287 (N_1287,In_1529,In_1869);
and U1288 (N_1288,In_361,In_486);
nor U1289 (N_1289,In_1255,In_1981);
nand U1290 (N_1290,In_1969,In_1614);
or U1291 (N_1291,In_1405,In_421);
and U1292 (N_1292,In_1215,In_1644);
nor U1293 (N_1293,In_1421,In_647);
nor U1294 (N_1294,In_1861,In_1208);
and U1295 (N_1295,In_1378,In_1401);
and U1296 (N_1296,In_840,In_357);
nor U1297 (N_1297,In_1962,In_330);
nor U1298 (N_1298,In_1872,In_370);
nor U1299 (N_1299,In_580,In_750);
nor U1300 (N_1300,In_176,In_1431);
and U1301 (N_1301,In_433,In_1231);
or U1302 (N_1302,In_1684,In_428);
xor U1303 (N_1303,In_187,In_808);
and U1304 (N_1304,In_225,In_50);
nor U1305 (N_1305,In_1000,In_374);
nand U1306 (N_1306,In_998,In_547);
and U1307 (N_1307,In_1991,In_1451);
nand U1308 (N_1308,In_680,In_1677);
or U1309 (N_1309,In_1524,In_859);
xor U1310 (N_1310,In_1868,In_59);
nand U1311 (N_1311,In_1832,In_499);
nand U1312 (N_1312,In_761,In_444);
nor U1313 (N_1313,In_318,In_564);
or U1314 (N_1314,In_1830,In_1489);
or U1315 (N_1315,In_1297,In_88);
nand U1316 (N_1316,In_851,In_318);
or U1317 (N_1317,In_758,In_1931);
and U1318 (N_1318,In_1002,In_157);
nor U1319 (N_1319,In_798,In_267);
and U1320 (N_1320,In_255,In_1623);
and U1321 (N_1321,In_1484,In_650);
nand U1322 (N_1322,In_920,In_783);
nand U1323 (N_1323,In_1624,In_1991);
nor U1324 (N_1324,In_1672,In_1632);
nand U1325 (N_1325,In_1725,In_1768);
nor U1326 (N_1326,In_431,In_323);
nand U1327 (N_1327,In_283,In_335);
nand U1328 (N_1328,In_1382,In_916);
or U1329 (N_1329,In_1666,In_662);
xnor U1330 (N_1330,In_1040,In_1270);
and U1331 (N_1331,In_1450,In_1093);
or U1332 (N_1332,In_1708,In_81);
or U1333 (N_1333,In_1341,In_1143);
nand U1334 (N_1334,In_511,In_1727);
nor U1335 (N_1335,In_1422,In_1424);
and U1336 (N_1336,In_1290,In_722);
or U1337 (N_1337,In_1960,In_1953);
nor U1338 (N_1338,In_1489,In_127);
xor U1339 (N_1339,In_2,In_1949);
or U1340 (N_1340,In_517,In_47);
nor U1341 (N_1341,In_479,In_1171);
or U1342 (N_1342,In_1351,In_1741);
nand U1343 (N_1343,In_894,In_811);
and U1344 (N_1344,In_1355,In_1167);
or U1345 (N_1345,In_818,In_1223);
nor U1346 (N_1346,In_2,In_1286);
and U1347 (N_1347,In_658,In_1493);
nor U1348 (N_1348,In_793,In_695);
and U1349 (N_1349,In_1534,In_1532);
nor U1350 (N_1350,In_934,In_326);
nor U1351 (N_1351,In_406,In_924);
nand U1352 (N_1352,In_45,In_1343);
nor U1353 (N_1353,In_1911,In_263);
nor U1354 (N_1354,In_266,In_1395);
and U1355 (N_1355,In_700,In_14);
or U1356 (N_1356,In_1031,In_1664);
or U1357 (N_1357,In_850,In_1878);
nand U1358 (N_1358,In_1243,In_946);
nor U1359 (N_1359,In_364,In_1916);
or U1360 (N_1360,In_1883,In_1509);
nor U1361 (N_1361,In_1257,In_1440);
nand U1362 (N_1362,In_1245,In_73);
and U1363 (N_1363,In_1738,In_699);
nand U1364 (N_1364,In_1622,In_1709);
nand U1365 (N_1365,In_1029,In_1229);
nand U1366 (N_1366,In_638,In_737);
and U1367 (N_1367,In_41,In_1295);
nand U1368 (N_1368,In_1481,In_904);
nor U1369 (N_1369,In_1642,In_1679);
and U1370 (N_1370,In_1412,In_1142);
and U1371 (N_1371,In_1261,In_1167);
nor U1372 (N_1372,In_403,In_1224);
nand U1373 (N_1373,In_1037,In_1999);
or U1374 (N_1374,In_802,In_422);
nand U1375 (N_1375,In_1877,In_1179);
nand U1376 (N_1376,In_173,In_647);
nand U1377 (N_1377,In_117,In_91);
or U1378 (N_1378,In_1566,In_967);
and U1379 (N_1379,In_1681,In_477);
and U1380 (N_1380,In_1456,In_812);
or U1381 (N_1381,In_1104,In_1333);
nor U1382 (N_1382,In_753,In_1174);
nand U1383 (N_1383,In_1252,In_1063);
nand U1384 (N_1384,In_189,In_1161);
or U1385 (N_1385,In_1401,In_366);
nor U1386 (N_1386,In_303,In_127);
and U1387 (N_1387,In_738,In_664);
nand U1388 (N_1388,In_1976,In_1583);
or U1389 (N_1389,In_1991,In_1129);
xor U1390 (N_1390,In_909,In_1070);
nor U1391 (N_1391,In_615,In_92);
or U1392 (N_1392,In_1421,In_178);
nor U1393 (N_1393,In_689,In_1075);
or U1394 (N_1394,In_1934,In_924);
nand U1395 (N_1395,In_1459,In_1998);
and U1396 (N_1396,In_887,In_760);
and U1397 (N_1397,In_1716,In_400);
nor U1398 (N_1398,In_506,In_898);
or U1399 (N_1399,In_411,In_1413);
and U1400 (N_1400,In_1831,In_203);
nor U1401 (N_1401,In_1479,In_326);
nand U1402 (N_1402,In_495,In_1819);
and U1403 (N_1403,In_1552,In_1255);
xnor U1404 (N_1404,In_257,In_880);
and U1405 (N_1405,In_1833,In_393);
nor U1406 (N_1406,In_1691,In_80);
and U1407 (N_1407,In_872,In_1104);
and U1408 (N_1408,In_1920,In_1985);
nor U1409 (N_1409,In_271,In_968);
or U1410 (N_1410,In_1351,In_1657);
nand U1411 (N_1411,In_1133,In_990);
and U1412 (N_1412,In_1664,In_1161);
or U1413 (N_1413,In_1406,In_1205);
or U1414 (N_1414,In_126,In_1694);
nand U1415 (N_1415,In_230,In_209);
nand U1416 (N_1416,In_680,In_704);
nand U1417 (N_1417,In_1244,In_1142);
and U1418 (N_1418,In_655,In_807);
and U1419 (N_1419,In_261,In_894);
or U1420 (N_1420,In_975,In_973);
and U1421 (N_1421,In_906,In_1495);
or U1422 (N_1422,In_1549,In_925);
or U1423 (N_1423,In_347,In_1143);
xor U1424 (N_1424,In_979,In_510);
and U1425 (N_1425,In_1072,In_1488);
or U1426 (N_1426,In_1976,In_26);
nand U1427 (N_1427,In_1427,In_31);
and U1428 (N_1428,In_632,In_448);
or U1429 (N_1429,In_181,In_509);
nand U1430 (N_1430,In_1086,In_1067);
nand U1431 (N_1431,In_1273,In_596);
and U1432 (N_1432,In_1116,In_144);
and U1433 (N_1433,In_1440,In_655);
and U1434 (N_1434,In_34,In_524);
and U1435 (N_1435,In_740,In_1257);
or U1436 (N_1436,In_515,In_252);
nand U1437 (N_1437,In_274,In_230);
and U1438 (N_1438,In_246,In_1769);
and U1439 (N_1439,In_1063,In_1524);
nor U1440 (N_1440,In_173,In_1019);
or U1441 (N_1441,In_1275,In_333);
nor U1442 (N_1442,In_1552,In_350);
and U1443 (N_1443,In_1555,In_805);
nor U1444 (N_1444,In_373,In_1339);
nand U1445 (N_1445,In_307,In_858);
nand U1446 (N_1446,In_1135,In_324);
nor U1447 (N_1447,In_1728,In_862);
and U1448 (N_1448,In_1622,In_157);
or U1449 (N_1449,In_269,In_1619);
or U1450 (N_1450,In_713,In_471);
and U1451 (N_1451,In_1988,In_1273);
nand U1452 (N_1452,In_1528,In_1610);
and U1453 (N_1453,In_1097,In_1562);
and U1454 (N_1454,In_1887,In_14);
xor U1455 (N_1455,In_1962,In_1184);
or U1456 (N_1456,In_1509,In_501);
nor U1457 (N_1457,In_1872,In_17);
xor U1458 (N_1458,In_678,In_1297);
and U1459 (N_1459,In_1938,In_1220);
nor U1460 (N_1460,In_1314,In_1381);
or U1461 (N_1461,In_412,In_1286);
or U1462 (N_1462,In_912,In_1967);
nand U1463 (N_1463,In_1002,In_1441);
xnor U1464 (N_1464,In_401,In_1158);
nor U1465 (N_1465,In_1187,In_1579);
nor U1466 (N_1466,In_1529,In_1913);
and U1467 (N_1467,In_65,In_1107);
and U1468 (N_1468,In_136,In_392);
nor U1469 (N_1469,In_158,In_1411);
nor U1470 (N_1470,In_732,In_1444);
xor U1471 (N_1471,In_1891,In_848);
nor U1472 (N_1472,In_1865,In_1588);
and U1473 (N_1473,In_1397,In_704);
nand U1474 (N_1474,In_625,In_1775);
or U1475 (N_1475,In_1229,In_986);
nor U1476 (N_1476,In_1475,In_1443);
or U1477 (N_1477,In_282,In_1099);
and U1478 (N_1478,In_595,In_461);
nand U1479 (N_1479,In_1464,In_1835);
or U1480 (N_1480,In_928,In_1341);
nand U1481 (N_1481,In_1512,In_1057);
xor U1482 (N_1482,In_1122,In_965);
and U1483 (N_1483,In_112,In_811);
or U1484 (N_1484,In_650,In_596);
nand U1485 (N_1485,In_1390,In_472);
xor U1486 (N_1486,In_33,In_658);
nor U1487 (N_1487,In_1485,In_1134);
nand U1488 (N_1488,In_683,In_1937);
and U1489 (N_1489,In_1272,In_1677);
nand U1490 (N_1490,In_458,In_922);
nand U1491 (N_1491,In_1855,In_719);
nor U1492 (N_1492,In_1821,In_769);
nand U1493 (N_1493,In_1967,In_1295);
nand U1494 (N_1494,In_1476,In_1491);
nor U1495 (N_1495,In_1109,In_1033);
nor U1496 (N_1496,In_1188,In_1329);
or U1497 (N_1497,In_786,In_1016);
and U1498 (N_1498,In_1095,In_1637);
nor U1499 (N_1499,In_841,In_1457);
and U1500 (N_1500,In_1244,In_35);
xor U1501 (N_1501,In_216,In_1374);
nand U1502 (N_1502,In_1514,In_1857);
and U1503 (N_1503,In_216,In_798);
nand U1504 (N_1504,In_1429,In_373);
nor U1505 (N_1505,In_697,In_1193);
or U1506 (N_1506,In_700,In_400);
or U1507 (N_1507,In_1228,In_1430);
nand U1508 (N_1508,In_1776,In_1390);
nand U1509 (N_1509,In_242,In_364);
nor U1510 (N_1510,In_488,In_555);
nand U1511 (N_1511,In_1222,In_657);
nand U1512 (N_1512,In_1313,In_1572);
nand U1513 (N_1513,In_1588,In_1597);
and U1514 (N_1514,In_57,In_1241);
and U1515 (N_1515,In_783,In_1039);
nand U1516 (N_1516,In_23,In_1913);
nor U1517 (N_1517,In_868,In_163);
and U1518 (N_1518,In_1063,In_739);
nand U1519 (N_1519,In_371,In_299);
or U1520 (N_1520,In_1206,In_983);
or U1521 (N_1521,In_1678,In_669);
or U1522 (N_1522,In_1459,In_1820);
nor U1523 (N_1523,In_201,In_110);
and U1524 (N_1524,In_1682,In_1353);
or U1525 (N_1525,In_569,In_836);
nor U1526 (N_1526,In_1196,In_1623);
nor U1527 (N_1527,In_305,In_163);
and U1528 (N_1528,In_1657,In_342);
and U1529 (N_1529,In_1421,In_704);
nor U1530 (N_1530,In_171,In_1333);
or U1531 (N_1531,In_1010,In_389);
and U1532 (N_1532,In_479,In_1861);
and U1533 (N_1533,In_1491,In_1083);
nand U1534 (N_1534,In_672,In_199);
or U1535 (N_1535,In_1144,In_42);
or U1536 (N_1536,In_420,In_387);
and U1537 (N_1537,In_141,In_730);
nor U1538 (N_1538,In_1826,In_1257);
or U1539 (N_1539,In_172,In_932);
nor U1540 (N_1540,In_323,In_370);
xnor U1541 (N_1541,In_1982,In_146);
and U1542 (N_1542,In_1736,In_281);
nand U1543 (N_1543,In_1480,In_1332);
and U1544 (N_1544,In_327,In_302);
nand U1545 (N_1545,In_30,In_124);
nand U1546 (N_1546,In_1821,In_454);
or U1547 (N_1547,In_202,In_1532);
nand U1548 (N_1548,In_1887,In_1081);
nor U1549 (N_1549,In_830,In_618);
nor U1550 (N_1550,In_254,In_1599);
or U1551 (N_1551,In_1896,In_238);
nand U1552 (N_1552,In_1134,In_157);
nor U1553 (N_1553,In_1994,In_345);
nand U1554 (N_1554,In_869,In_110);
nand U1555 (N_1555,In_50,In_963);
nand U1556 (N_1556,In_167,In_1577);
or U1557 (N_1557,In_573,In_852);
nand U1558 (N_1558,In_378,In_141);
nand U1559 (N_1559,In_1151,In_1239);
and U1560 (N_1560,In_1436,In_318);
and U1561 (N_1561,In_1256,In_474);
or U1562 (N_1562,In_1343,In_1211);
xor U1563 (N_1563,In_1575,In_144);
nor U1564 (N_1564,In_730,In_1574);
nand U1565 (N_1565,In_1079,In_1340);
nand U1566 (N_1566,In_1049,In_840);
nor U1567 (N_1567,In_762,In_371);
and U1568 (N_1568,In_405,In_1380);
nand U1569 (N_1569,In_483,In_762);
nand U1570 (N_1570,In_1501,In_459);
nand U1571 (N_1571,In_1175,In_1146);
and U1572 (N_1572,In_179,In_221);
and U1573 (N_1573,In_1839,In_1612);
and U1574 (N_1574,In_1144,In_620);
and U1575 (N_1575,In_859,In_1996);
or U1576 (N_1576,In_23,In_253);
nor U1577 (N_1577,In_1738,In_1035);
or U1578 (N_1578,In_1663,In_937);
nand U1579 (N_1579,In_1910,In_544);
and U1580 (N_1580,In_1457,In_1180);
and U1581 (N_1581,In_1384,In_376);
nand U1582 (N_1582,In_1370,In_1022);
and U1583 (N_1583,In_1261,In_667);
or U1584 (N_1584,In_202,In_636);
nand U1585 (N_1585,In_949,In_1646);
xnor U1586 (N_1586,In_99,In_1319);
nand U1587 (N_1587,In_1277,In_702);
and U1588 (N_1588,In_563,In_68);
and U1589 (N_1589,In_1636,In_1926);
and U1590 (N_1590,In_722,In_866);
xor U1591 (N_1591,In_1284,In_1270);
nand U1592 (N_1592,In_434,In_1654);
or U1593 (N_1593,In_1914,In_703);
nor U1594 (N_1594,In_1322,In_1580);
or U1595 (N_1595,In_1465,In_96);
nor U1596 (N_1596,In_90,In_1845);
nand U1597 (N_1597,In_1655,In_1640);
nand U1598 (N_1598,In_1356,In_297);
nor U1599 (N_1599,In_1783,In_201);
or U1600 (N_1600,In_1174,In_761);
xor U1601 (N_1601,In_908,In_1415);
and U1602 (N_1602,In_1610,In_1177);
nand U1603 (N_1603,In_233,In_1827);
and U1604 (N_1604,In_1023,In_646);
nand U1605 (N_1605,In_665,In_826);
and U1606 (N_1606,In_1864,In_1862);
or U1607 (N_1607,In_1997,In_199);
and U1608 (N_1608,In_498,In_800);
or U1609 (N_1609,In_1906,In_1735);
xnor U1610 (N_1610,In_1223,In_1764);
nor U1611 (N_1611,In_1780,In_1079);
nand U1612 (N_1612,In_1852,In_407);
and U1613 (N_1613,In_1672,In_957);
or U1614 (N_1614,In_1069,In_1595);
or U1615 (N_1615,In_467,In_1198);
or U1616 (N_1616,In_42,In_1703);
and U1617 (N_1617,In_1782,In_1247);
and U1618 (N_1618,In_1548,In_960);
xnor U1619 (N_1619,In_386,In_1258);
nand U1620 (N_1620,In_828,In_1587);
or U1621 (N_1621,In_1331,In_1551);
xor U1622 (N_1622,In_1243,In_329);
or U1623 (N_1623,In_107,In_926);
or U1624 (N_1624,In_1934,In_1180);
or U1625 (N_1625,In_15,In_495);
xor U1626 (N_1626,In_113,In_1392);
xor U1627 (N_1627,In_1635,In_281);
xnor U1628 (N_1628,In_524,In_47);
nor U1629 (N_1629,In_261,In_107);
and U1630 (N_1630,In_1645,In_1840);
nand U1631 (N_1631,In_343,In_1758);
nor U1632 (N_1632,In_385,In_1856);
nor U1633 (N_1633,In_99,In_105);
or U1634 (N_1634,In_402,In_1952);
and U1635 (N_1635,In_1262,In_1967);
nor U1636 (N_1636,In_734,In_1300);
nand U1637 (N_1637,In_68,In_1132);
and U1638 (N_1638,In_609,In_856);
or U1639 (N_1639,In_1235,In_888);
and U1640 (N_1640,In_1947,In_1067);
and U1641 (N_1641,In_906,In_131);
or U1642 (N_1642,In_1401,In_738);
nor U1643 (N_1643,In_487,In_626);
xor U1644 (N_1644,In_1384,In_1397);
nor U1645 (N_1645,In_788,In_1018);
and U1646 (N_1646,In_180,In_1350);
nand U1647 (N_1647,In_1224,In_454);
nand U1648 (N_1648,In_1067,In_91);
or U1649 (N_1649,In_1157,In_214);
nand U1650 (N_1650,In_360,In_1696);
xor U1651 (N_1651,In_585,In_1167);
or U1652 (N_1652,In_856,In_198);
nor U1653 (N_1653,In_78,In_861);
or U1654 (N_1654,In_1296,In_613);
nand U1655 (N_1655,In_1613,In_1386);
and U1656 (N_1656,In_92,In_1413);
or U1657 (N_1657,In_1861,In_472);
nand U1658 (N_1658,In_564,In_1992);
and U1659 (N_1659,In_1406,In_310);
nand U1660 (N_1660,In_1709,In_26);
and U1661 (N_1661,In_1245,In_1840);
or U1662 (N_1662,In_29,In_582);
nor U1663 (N_1663,In_1821,In_1979);
nand U1664 (N_1664,In_656,In_14);
nand U1665 (N_1665,In_1800,In_1008);
and U1666 (N_1666,In_600,In_572);
and U1667 (N_1667,In_844,In_1881);
xnor U1668 (N_1668,In_990,In_464);
nor U1669 (N_1669,In_1918,In_114);
nor U1670 (N_1670,In_605,In_1149);
and U1671 (N_1671,In_890,In_1584);
or U1672 (N_1672,In_1821,In_263);
nor U1673 (N_1673,In_111,In_811);
nor U1674 (N_1674,In_815,In_1022);
or U1675 (N_1675,In_879,In_1332);
xor U1676 (N_1676,In_905,In_1961);
or U1677 (N_1677,In_848,In_1608);
nor U1678 (N_1678,In_384,In_1461);
xnor U1679 (N_1679,In_442,In_972);
nand U1680 (N_1680,In_776,In_1959);
xnor U1681 (N_1681,In_1069,In_118);
and U1682 (N_1682,In_1166,In_1170);
and U1683 (N_1683,In_1862,In_1952);
nand U1684 (N_1684,In_1275,In_319);
nor U1685 (N_1685,In_1938,In_366);
nand U1686 (N_1686,In_402,In_239);
nand U1687 (N_1687,In_1630,In_1836);
nor U1688 (N_1688,In_651,In_527);
nor U1689 (N_1689,In_1062,In_1721);
nor U1690 (N_1690,In_894,In_1288);
and U1691 (N_1691,In_131,In_1337);
xor U1692 (N_1692,In_1917,In_493);
or U1693 (N_1693,In_1732,In_1655);
and U1694 (N_1694,In_1655,In_1380);
or U1695 (N_1695,In_615,In_319);
or U1696 (N_1696,In_172,In_392);
or U1697 (N_1697,In_1650,In_1020);
and U1698 (N_1698,In_892,In_220);
nor U1699 (N_1699,In_459,In_1751);
nand U1700 (N_1700,In_812,In_1271);
or U1701 (N_1701,In_32,In_665);
nand U1702 (N_1702,In_845,In_1192);
nor U1703 (N_1703,In_1661,In_1139);
nand U1704 (N_1704,In_1428,In_809);
nand U1705 (N_1705,In_1596,In_514);
nor U1706 (N_1706,In_700,In_730);
or U1707 (N_1707,In_1844,In_446);
nor U1708 (N_1708,In_607,In_68);
or U1709 (N_1709,In_1389,In_1730);
nand U1710 (N_1710,In_1256,In_208);
nand U1711 (N_1711,In_602,In_1979);
nand U1712 (N_1712,In_783,In_1368);
and U1713 (N_1713,In_1710,In_1825);
or U1714 (N_1714,In_608,In_637);
or U1715 (N_1715,In_1834,In_1058);
and U1716 (N_1716,In_969,In_1738);
nor U1717 (N_1717,In_821,In_1029);
nand U1718 (N_1718,In_1066,In_1581);
nor U1719 (N_1719,In_1540,In_1054);
nand U1720 (N_1720,In_1604,In_298);
nand U1721 (N_1721,In_949,In_613);
or U1722 (N_1722,In_1542,In_1319);
nor U1723 (N_1723,In_1622,In_467);
xor U1724 (N_1724,In_1019,In_471);
and U1725 (N_1725,In_162,In_1492);
xor U1726 (N_1726,In_897,In_1822);
nand U1727 (N_1727,In_845,In_1252);
and U1728 (N_1728,In_186,In_1279);
and U1729 (N_1729,In_736,In_197);
xnor U1730 (N_1730,In_949,In_518);
nor U1731 (N_1731,In_1144,In_965);
nor U1732 (N_1732,In_1237,In_1076);
nor U1733 (N_1733,In_1046,In_836);
nand U1734 (N_1734,In_1244,In_1989);
and U1735 (N_1735,In_1180,In_759);
and U1736 (N_1736,In_1560,In_1400);
nor U1737 (N_1737,In_1382,In_39);
nor U1738 (N_1738,In_310,In_1094);
nor U1739 (N_1739,In_1524,In_548);
nor U1740 (N_1740,In_1146,In_1241);
nand U1741 (N_1741,In_624,In_1889);
and U1742 (N_1742,In_985,In_1910);
nor U1743 (N_1743,In_1963,In_1031);
nor U1744 (N_1744,In_58,In_1800);
and U1745 (N_1745,In_1952,In_1600);
and U1746 (N_1746,In_1066,In_1173);
nor U1747 (N_1747,In_1130,In_1587);
and U1748 (N_1748,In_811,In_1721);
nor U1749 (N_1749,In_978,In_1708);
and U1750 (N_1750,In_12,In_433);
nor U1751 (N_1751,In_718,In_1224);
or U1752 (N_1752,In_1807,In_430);
or U1753 (N_1753,In_871,In_442);
or U1754 (N_1754,In_1132,In_198);
nand U1755 (N_1755,In_1477,In_948);
or U1756 (N_1756,In_679,In_1715);
nand U1757 (N_1757,In_149,In_1142);
nand U1758 (N_1758,In_71,In_457);
xnor U1759 (N_1759,In_1904,In_1898);
or U1760 (N_1760,In_50,In_1807);
or U1761 (N_1761,In_304,In_136);
xor U1762 (N_1762,In_450,In_850);
nor U1763 (N_1763,In_713,In_1206);
nand U1764 (N_1764,In_1194,In_1475);
nand U1765 (N_1765,In_735,In_1498);
nor U1766 (N_1766,In_1407,In_1664);
and U1767 (N_1767,In_565,In_177);
xnor U1768 (N_1768,In_1715,In_291);
and U1769 (N_1769,In_1734,In_1336);
nand U1770 (N_1770,In_913,In_1237);
or U1771 (N_1771,In_1726,In_1954);
and U1772 (N_1772,In_1088,In_191);
nor U1773 (N_1773,In_246,In_40);
nor U1774 (N_1774,In_107,In_299);
xnor U1775 (N_1775,In_1822,In_1699);
nand U1776 (N_1776,In_199,In_79);
nor U1777 (N_1777,In_167,In_1547);
nor U1778 (N_1778,In_471,In_1220);
nand U1779 (N_1779,In_305,In_165);
or U1780 (N_1780,In_1599,In_989);
or U1781 (N_1781,In_157,In_454);
and U1782 (N_1782,In_41,In_91);
nand U1783 (N_1783,In_1767,In_507);
or U1784 (N_1784,In_700,In_1966);
or U1785 (N_1785,In_514,In_211);
nand U1786 (N_1786,In_968,In_1181);
or U1787 (N_1787,In_101,In_1769);
or U1788 (N_1788,In_546,In_718);
nand U1789 (N_1789,In_947,In_1655);
nand U1790 (N_1790,In_596,In_745);
nor U1791 (N_1791,In_1899,In_886);
xor U1792 (N_1792,In_1547,In_898);
nand U1793 (N_1793,In_722,In_1559);
nor U1794 (N_1794,In_39,In_772);
nand U1795 (N_1795,In_597,In_1548);
nor U1796 (N_1796,In_1717,In_1230);
nor U1797 (N_1797,In_1192,In_818);
or U1798 (N_1798,In_1322,In_254);
nand U1799 (N_1799,In_1576,In_1351);
nor U1800 (N_1800,In_1189,In_1907);
nor U1801 (N_1801,In_376,In_1319);
nand U1802 (N_1802,In_1785,In_1475);
nor U1803 (N_1803,In_21,In_382);
or U1804 (N_1804,In_779,In_675);
or U1805 (N_1805,In_195,In_976);
and U1806 (N_1806,In_1001,In_1141);
nor U1807 (N_1807,In_1534,In_621);
and U1808 (N_1808,In_869,In_1405);
nor U1809 (N_1809,In_1877,In_230);
xor U1810 (N_1810,In_519,In_1737);
nor U1811 (N_1811,In_438,In_1132);
xor U1812 (N_1812,In_537,In_205);
nand U1813 (N_1813,In_1726,In_139);
or U1814 (N_1814,In_1623,In_147);
and U1815 (N_1815,In_419,In_580);
or U1816 (N_1816,In_1132,In_1089);
nand U1817 (N_1817,In_321,In_1041);
nand U1818 (N_1818,In_1451,In_301);
or U1819 (N_1819,In_51,In_793);
and U1820 (N_1820,In_286,In_1719);
nor U1821 (N_1821,In_1316,In_974);
nor U1822 (N_1822,In_1069,In_1354);
or U1823 (N_1823,In_1260,In_405);
or U1824 (N_1824,In_1891,In_572);
and U1825 (N_1825,In_345,In_0);
or U1826 (N_1826,In_1211,In_376);
or U1827 (N_1827,In_1751,In_1327);
nand U1828 (N_1828,In_221,In_1057);
nor U1829 (N_1829,In_526,In_1169);
nand U1830 (N_1830,In_893,In_930);
or U1831 (N_1831,In_1949,In_523);
xor U1832 (N_1832,In_943,In_1920);
xor U1833 (N_1833,In_400,In_492);
and U1834 (N_1834,In_731,In_818);
and U1835 (N_1835,In_1179,In_626);
nor U1836 (N_1836,In_745,In_1836);
and U1837 (N_1837,In_1495,In_773);
and U1838 (N_1838,In_1801,In_860);
nor U1839 (N_1839,In_271,In_470);
xor U1840 (N_1840,In_308,In_1106);
xnor U1841 (N_1841,In_1397,In_1554);
or U1842 (N_1842,In_904,In_661);
and U1843 (N_1843,In_1326,In_1775);
nand U1844 (N_1844,In_1308,In_917);
nand U1845 (N_1845,In_1032,In_1262);
or U1846 (N_1846,In_1527,In_468);
or U1847 (N_1847,In_472,In_1863);
nand U1848 (N_1848,In_591,In_116);
nor U1849 (N_1849,In_785,In_538);
or U1850 (N_1850,In_1788,In_88);
or U1851 (N_1851,In_31,In_42);
nor U1852 (N_1852,In_262,In_502);
or U1853 (N_1853,In_1542,In_588);
xor U1854 (N_1854,In_1715,In_1828);
nor U1855 (N_1855,In_90,In_900);
or U1856 (N_1856,In_1414,In_1018);
nand U1857 (N_1857,In_1498,In_68);
or U1858 (N_1858,In_1268,In_120);
xor U1859 (N_1859,In_642,In_1857);
nor U1860 (N_1860,In_1010,In_1465);
nor U1861 (N_1861,In_1663,In_556);
and U1862 (N_1862,In_138,In_1138);
or U1863 (N_1863,In_243,In_388);
nand U1864 (N_1864,In_494,In_1730);
nand U1865 (N_1865,In_1500,In_451);
or U1866 (N_1866,In_1527,In_1888);
or U1867 (N_1867,In_426,In_710);
nor U1868 (N_1868,In_1129,In_780);
or U1869 (N_1869,In_1296,In_738);
nor U1870 (N_1870,In_1474,In_521);
nor U1871 (N_1871,In_485,In_1423);
xnor U1872 (N_1872,In_125,In_669);
nor U1873 (N_1873,In_1348,In_75);
nor U1874 (N_1874,In_1376,In_1473);
nor U1875 (N_1875,In_987,In_291);
xor U1876 (N_1876,In_1985,In_1202);
xnor U1877 (N_1877,In_1628,In_61);
nand U1878 (N_1878,In_279,In_1613);
and U1879 (N_1879,In_408,In_1381);
or U1880 (N_1880,In_288,In_73);
nand U1881 (N_1881,In_1374,In_1832);
or U1882 (N_1882,In_311,In_125);
or U1883 (N_1883,In_798,In_1089);
nand U1884 (N_1884,In_1004,In_43);
xor U1885 (N_1885,In_292,In_560);
and U1886 (N_1886,In_754,In_272);
and U1887 (N_1887,In_1612,In_1452);
xnor U1888 (N_1888,In_1901,In_1124);
xor U1889 (N_1889,In_174,In_88);
and U1890 (N_1890,In_1626,In_1625);
nor U1891 (N_1891,In_755,In_783);
xor U1892 (N_1892,In_796,In_1652);
or U1893 (N_1893,In_264,In_56);
nand U1894 (N_1894,In_840,In_1946);
nand U1895 (N_1895,In_1450,In_828);
nor U1896 (N_1896,In_370,In_750);
nor U1897 (N_1897,In_1420,In_465);
and U1898 (N_1898,In_81,In_114);
and U1899 (N_1899,In_1836,In_1502);
nand U1900 (N_1900,In_829,In_735);
nor U1901 (N_1901,In_1151,In_1633);
nand U1902 (N_1902,In_1929,In_153);
xnor U1903 (N_1903,In_14,In_673);
nor U1904 (N_1904,In_1360,In_1113);
nand U1905 (N_1905,In_660,In_642);
and U1906 (N_1906,In_1780,In_125);
nand U1907 (N_1907,In_782,In_723);
xor U1908 (N_1908,In_1432,In_1054);
nand U1909 (N_1909,In_1358,In_480);
and U1910 (N_1910,In_600,In_316);
and U1911 (N_1911,In_1929,In_483);
nor U1912 (N_1912,In_345,In_140);
nand U1913 (N_1913,In_18,In_1893);
and U1914 (N_1914,In_534,In_1270);
and U1915 (N_1915,In_273,In_1571);
nand U1916 (N_1916,In_1610,In_674);
nor U1917 (N_1917,In_263,In_1979);
or U1918 (N_1918,In_1659,In_375);
or U1919 (N_1919,In_309,In_934);
and U1920 (N_1920,In_1267,In_808);
nand U1921 (N_1921,In_318,In_218);
nor U1922 (N_1922,In_65,In_697);
nand U1923 (N_1923,In_597,In_873);
nor U1924 (N_1924,In_781,In_162);
or U1925 (N_1925,In_619,In_1205);
nor U1926 (N_1926,In_97,In_1777);
nand U1927 (N_1927,In_1383,In_17);
nand U1928 (N_1928,In_458,In_1894);
nand U1929 (N_1929,In_825,In_343);
nor U1930 (N_1930,In_667,In_554);
nor U1931 (N_1931,In_1685,In_717);
nor U1932 (N_1932,In_393,In_914);
and U1933 (N_1933,In_457,In_870);
nand U1934 (N_1934,In_1868,In_1812);
nor U1935 (N_1935,In_1717,In_1475);
and U1936 (N_1936,In_283,In_383);
or U1937 (N_1937,In_1148,In_358);
xnor U1938 (N_1938,In_1205,In_871);
nand U1939 (N_1939,In_815,In_1417);
or U1940 (N_1940,In_1010,In_1714);
and U1941 (N_1941,In_1904,In_238);
or U1942 (N_1942,In_369,In_217);
or U1943 (N_1943,In_1624,In_1348);
or U1944 (N_1944,In_305,In_284);
or U1945 (N_1945,In_1302,In_8);
or U1946 (N_1946,In_331,In_1242);
nand U1947 (N_1947,In_336,In_1163);
nand U1948 (N_1948,In_1580,In_1514);
nand U1949 (N_1949,In_1178,In_1137);
xor U1950 (N_1950,In_900,In_1766);
nor U1951 (N_1951,In_433,In_1079);
xor U1952 (N_1952,In_1178,In_1332);
nor U1953 (N_1953,In_296,In_1452);
nor U1954 (N_1954,In_1149,In_1106);
nor U1955 (N_1955,In_1300,In_534);
and U1956 (N_1956,In_14,In_1423);
nor U1957 (N_1957,In_1615,In_907);
and U1958 (N_1958,In_788,In_1974);
or U1959 (N_1959,In_1653,In_439);
or U1960 (N_1960,In_1291,In_1601);
and U1961 (N_1961,In_416,In_317);
nor U1962 (N_1962,In_1750,In_735);
nor U1963 (N_1963,In_1616,In_933);
nor U1964 (N_1964,In_1076,In_1700);
nand U1965 (N_1965,In_1587,In_1302);
and U1966 (N_1966,In_681,In_187);
xor U1967 (N_1967,In_536,In_464);
or U1968 (N_1968,In_531,In_1689);
and U1969 (N_1969,In_1308,In_1357);
nor U1970 (N_1970,In_1992,In_351);
and U1971 (N_1971,In_202,In_972);
and U1972 (N_1972,In_216,In_1793);
xnor U1973 (N_1973,In_62,In_592);
nand U1974 (N_1974,In_1800,In_156);
nor U1975 (N_1975,In_1519,In_1566);
nand U1976 (N_1976,In_1917,In_1968);
nor U1977 (N_1977,In_1483,In_235);
nand U1978 (N_1978,In_845,In_324);
and U1979 (N_1979,In_1783,In_1969);
xnor U1980 (N_1980,In_1691,In_1286);
or U1981 (N_1981,In_311,In_1664);
nand U1982 (N_1982,In_615,In_1261);
xnor U1983 (N_1983,In_1573,In_235);
nor U1984 (N_1984,In_1763,In_1537);
and U1985 (N_1985,In_1475,In_594);
and U1986 (N_1986,In_1164,In_1485);
nand U1987 (N_1987,In_1189,In_1454);
and U1988 (N_1988,In_234,In_1321);
and U1989 (N_1989,In_335,In_1470);
and U1990 (N_1990,In_1062,In_1860);
nand U1991 (N_1991,In_884,In_1479);
nor U1992 (N_1992,In_592,In_1934);
and U1993 (N_1993,In_0,In_1949);
nor U1994 (N_1994,In_1567,In_1387);
xor U1995 (N_1995,In_783,In_1092);
and U1996 (N_1996,In_263,In_1271);
nor U1997 (N_1997,In_1282,In_1384);
and U1998 (N_1998,In_420,In_481);
or U1999 (N_1999,In_211,In_186);
and U2000 (N_2000,N_328,N_937);
nor U2001 (N_2001,N_688,N_701);
nor U2002 (N_2002,N_528,N_1801);
and U2003 (N_2003,N_1233,N_660);
and U2004 (N_2004,N_1009,N_1845);
or U2005 (N_2005,N_767,N_1237);
nand U2006 (N_2006,N_943,N_1004);
and U2007 (N_2007,N_1920,N_224);
nand U2008 (N_2008,N_1527,N_1789);
or U2009 (N_2009,N_468,N_1977);
nand U2010 (N_2010,N_1909,N_1366);
nor U2011 (N_2011,N_823,N_187);
or U2012 (N_2012,N_1903,N_49);
or U2013 (N_2013,N_42,N_65);
nor U2014 (N_2014,N_419,N_1324);
and U2015 (N_2015,N_4,N_1255);
nand U2016 (N_2016,N_1769,N_1250);
and U2017 (N_2017,N_731,N_146);
nand U2018 (N_2018,N_891,N_1905);
nand U2019 (N_2019,N_538,N_542);
or U2020 (N_2020,N_782,N_1260);
and U2021 (N_2021,N_703,N_1330);
and U2022 (N_2022,N_352,N_1022);
nor U2023 (N_2023,N_652,N_579);
or U2024 (N_2024,N_1877,N_1174);
nand U2025 (N_2025,N_137,N_1532);
nor U2026 (N_2026,N_322,N_788);
or U2027 (N_2027,N_321,N_1713);
nor U2028 (N_2028,N_1721,N_127);
nand U2029 (N_2029,N_774,N_1358);
nor U2030 (N_2030,N_470,N_118);
xor U2031 (N_2031,N_1427,N_534);
nor U2032 (N_2032,N_120,N_371);
nand U2033 (N_2033,N_1073,N_320);
and U2034 (N_2034,N_1616,N_790);
nor U2035 (N_2035,N_1817,N_346);
nand U2036 (N_2036,N_807,N_170);
nand U2037 (N_2037,N_12,N_682);
nand U2038 (N_2038,N_131,N_584);
or U2039 (N_2039,N_388,N_1630);
or U2040 (N_2040,N_1134,N_1377);
or U2041 (N_2041,N_429,N_112);
nor U2042 (N_2042,N_1695,N_1960);
nor U2043 (N_2043,N_1037,N_217);
nand U2044 (N_2044,N_1390,N_80);
nand U2045 (N_2045,N_953,N_1701);
or U2046 (N_2046,N_1947,N_1720);
nor U2047 (N_2047,N_1809,N_237);
nor U2048 (N_2048,N_1618,N_1738);
xnor U2049 (N_2049,N_1953,N_256);
nand U2050 (N_2050,N_1434,N_1168);
xnor U2051 (N_2051,N_72,N_990);
or U2052 (N_2052,N_272,N_1003);
nor U2053 (N_2053,N_1418,N_1808);
or U2054 (N_2054,N_940,N_420);
nand U2055 (N_2055,N_1535,N_527);
and U2056 (N_2056,N_1724,N_927);
and U2057 (N_2057,N_274,N_110);
and U2058 (N_2058,N_496,N_951);
nor U2059 (N_2059,N_276,N_1405);
and U2060 (N_2060,N_897,N_1671);
and U2061 (N_2061,N_1472,N_1286);
nand U2062 (N_2062,N_464,N_354);
or U2063 (N_2063,N_1144,N_1934);
and U2064 (N_2064,N_1991,N_758);
nor U2065 (N_2065,N_330,N_949);
or U2066 (N_2066,N_1088,N_559);
nor U2067 (N_2067,N_275,N_1807);
and U2068 (N_2068,N_1786,N_625);
nor U2069 (N_2069,N_442,N_934);
xor U2070 (N_2070,N_1647,N_1717);
nand U2071 (N_2071,N_1984,N_1445);
nor U2072 (N_2072,N_1475,N_134);
and U2073 (N_2073,N_373,N_786);
nand U2074 (N_2074,N_1213,N_608);
nand U2075 (N_2075,N_947,N_1800);
or U2076 (N_2076,N_655,N_1774);
nand U2077 (N_2077,N_1644,N_478);
nand U2078 (N_2078,N_163,N_1244);
or U2079 (N_2079,N_1439,N_1958);
nand U2080 (N_2080,N_234,N_1219);
xnor U2081 (N_2081,N_283,N_440);
and U2082 (N_2082,N_878,N_1457);
nand U2083 (N_2083,N_776,N_1334);
or U2084 (N_2084,N_1685,N_200);
nor U2085 (N_2085,N_1452,N_1007);
and U2086 (N_2086,N_610,N_1666);
nand U2087 (N_2087,N_178,N_653);
nor U2088 (N_2088,N_1495,N_1236);
nor U2089 (N_2089,N_1842,N_597);
or U2090 (N_2090,N_1454,N_1185);
xor U2091 (N_2091,N_115,N_1385);
nor U2092 (N_2092,N_545,N_1669);
nor U2093 (N_2093,N_991,N_474);
nand U2094 (N_2094,N_1468,N_693);
xnor U2095 (N_2095,N_1614,N_143);
or U2096 (N_2096,N_1910,N_142);
or U2097 (N_2097,N_1938,N_377);
nand U2098 (N_2098,N_312,N_1230);
nand U2099 (N_2099,N_748,N_1830);
and U2100 (N_2100,N_229,N_454);
or U2101 (N_2101,N_324,N_1756);
nand U2102 (N_2102,N_1613,N_1442);
and U2103 (N_2103,N_211,N_1222);
nand U2104 (N_2104,N_1231,N_1252);
and U2105 (N_2105,N_1187,N_1263);
nor U2106 (N_2106,N_1560,N_1523);
nand U2107 (N_2107,N_1719,N_390);
or U2108 (N_2108,N_325,N_1590);
nand U2109 (N_2109,N_995,N_1224);
nand U2110 (N_2110,N_1032,N_1804);
nand U2111 (N_2111,N_640,N_259);
nand U2112 (N_2112,N_326,N_1478);
or U2113 (N_2113,N_763,N_207);
nor U2114 (N_2114,N_485,N_252);
nor U2115 (N_2115,N_206,N_945);
or U2116 (N_2116,N_1112,N_1396);
xnor U2117 (N_2117,N_1728,N_753);
nand U2118 (N_2118,N_732,N_1421);
or U2119 (N_2119,N_1601,N_1915);
nand U2120 (N_2120,N_457,N_482);
nand U2121 (N_2121,N_556,N_1269);
nand U2122 (N_2122,N_125,N_600);
or U2123 (N_2123,N_1534,N_1514);
and U2124 (N_2124,N_1576,N_755);
and U2125 (N_2125,N_1592,N_1572);
and U2126 (N_2126,N_946,N_1172);
nor U2127 (N_2127,N_1974,N_1785);
and U2128 (N_2128,N_1218,N_973);
nor U2129 (N_2129,N_1556,N_85);
nor U2130 (N_2130,N_216,N_1981);
nor U2131 (N_2131,N_300,N_1023);
or U2132 (N_2132,N_1928,N_220);
nand U2133 (N_2133,N_15,N_382);
xor U2134 (N_2134,N_1841,N_1876);
or U2135 (N_2135,N_530,N_1759);
nand U2136 (N_2136,N_1379,N_1988);
nand U2137 (N_2137,N_109,N_1443);
nand U2138 (N_2138,N_737,N_1425);
and U2139 (N_2139,N_235,N_896);
and U2140 (N_2140,N_1661,N_1684);
or U2141 (N_2141,N_1622,N_155);
or U2142 (N_2142,N_409,N_1776);
and U2143 (N_2143,N_1598,N_1363);
xor U2144 (N_2144,N_396,N_1650);
nor U2145 (N_2145,N_1798,N_1050);
nor U2146 (N_2146,N_1961,N_261);
nand U2147 (N_2147,N_489,N_1325);
and U2148 (N_2148,N_1680,N_179);
and U2149 (N_2149,N_1152,N_884);
xor U2150 (N_2150,N_1065,N_344);
or U2151 (N_2151,N_1931,N_90);
and U2152 (N_2152,N_508,N_1524);
nor U2153 (N_2153,N_1249,N_893);
nand U2154 (N_2154,N_1059,N_315);
nand U2155 (N_2155,N_1536,N_680);
nor U2156 (N_2156,N_1151,N_1742);
and U2157 (N_2157,N_1683,N_1398);
and U2158 (N_2158,N_1469,N_1640);
nand U2159 (N_2159,N_1796,N_509);
nor U2160 (N_2160,N_1966,N_1580);
or U2161 (N_2161,N_647,N_974);
nand U2162 (N_2162,N_1555,N_1788);
nor U2163 (N_2163,N_1892,N_1773);
nor U2164 (N_2164,N_826,N_1304);
and U2165 (N_2165,N_709,N_1027);
and U2166 (N_2166,N_309,N_602);
or U2167 (N_2167,N_1150,N_1948);
nor U2168 (N_2168,N_385,N_867);
nor U2169 (N_2169,N_512,N_749);
nand U2170 (N_2170,N_733,N_540);
and U2171 (N_2171,N_739,N_103);
nand U2172 (N_2172,N_1133,N_191);
nor U2173 (N_2173,N_765,N_1856);
nand U2174 (N_2174,N_1649,N_1307);
and U2175 (N_2175,N_1485,N_1643);
and U2176 (N_2176,N_1462,N_1287);
nand U2177 (N_2177,N_1281,N_1161);
xnor U2178 (N_2178,N_395,N_977);
nor U2179 (N_2179,N_1351,N_184);
nor U2180 (N_2180,N_1766,N_1968);
nand U2181 (N_2181,N_1784,N_720);
nand U2182 (N_2182,N_1013,N_122);
and U2183 (N_2183,N_1939,N_1054);
and U2184 (N_2184,N_975,N_1030);
or U2185 (N_2185,N_1814,N_1705);
nor U2186 (N_2186,N_1567,N_243);
and U2187 (N_2187,N_1171,N_1783);
and U2188 (N_2188,N_333,N_626);
or U2189 (N_2189,N_1285,N_238);
nor U2190 (N_2190,N_1284,N_1319);
and U2191 (N_2191,N_687,N_1078);
or U2192 (N_2192,N_188,N_726);
nor U2193 (N_2193,N_161,N_832);
xnor U2194 (N_2194,N_886,N_1725);
nor U2195 (N_2195,N_1300,N_1505);
or U2196 (N_2196,N_1262,N_711);
or U2197 (N_2197,N_1173,N_1428);
or U2198 (N_2198,N_1952,N_1912);
nor U2199 (N_2199,N_1183,N_879);
and U2200 (N_2200,N_824,N_306);
and U2201 (N_2201,N_648,N_651);
nor U2202 (N_2202,N_1745,N_932);
nor U2203 (N_2203,N_1031,N_1041);
nand U2204 (N_2204,N_1641,N_1143);
xor U2205 (N_2205,N_1615,N_446);
or U2206 (N_2206,N_1651,N_985);
and U2207 (N_2207,N_1645,N_1209);
nor U2208 (N_2208,N_794,N_1875);
nor U2209 (N_2209,N_828,N_1781);
nor U2210 (N_2210,N_705,N_1554);
nor U2211 (N_2211,N_443,N_1289);
nand U2212 (N_2212,N_901,N_54);
or U2213 (N_2213,N_960,N_836);
or U2214 (N_2214,N_598,N_1341);
nor U2215 (N_2215,N_1757,N_1731);
nand U2216 (N_2216,N_1077,N_412);
and U2217 (N_2217,N_784,N_1111);
and U2218 (N_2218,N_1676,N_903);
nand U2219 (N_2219,N_1706,N_26);
xor U2220 (N_2220,N_0,N_455);
and U2221 (N_2221,N_831,N_872);
xnor U2222 (N_2222,N_180,N_1466);
or U2223 (N_2223,N_119,N_278);
and U2224 (N_2224,N_560,N_471);
nor U2225 (N_2225,N_145,N_875);
nor U2226 (N_2226,N_1432,N_89);
or U2227 (N_2227,N_404,N_1137);
and U2228 (N_2228,N_9,N_1955);
nor U2229 (N_2229,N_1058,N_59);
xor U2230 (N_2230,N_1194,N_591);
and U2231 (N_2231,N_1893,N_169);
nor U2232 (N_2232,N_1162,N_1001);
and U2233 (N_2233,N_154,N_24);
or U2234 (N_2234,N_1464,N_1400);
xnor U2235 (N_2235,N_1113,N_1811);
nand U2236 (N_2236,N_91,N_497);
nor U2237 (N_2237,N_1566,N_327);
or U2238 (N_2238,N_323,N_1607);
nor U2239 (N_2239,N_1326,N_132);
and U2240 (N_2240,N_815,N_1930);
or U2241 (N_2241,N_287,N_1299);
or U2242 (N_2242,N_1402,N_1820);
or U2243 (N_2243,N_1247,N_398);
or U2244 (N_2244,N_362,N_37);
xor U2245 (N_2245,N_1487,N_1937);
nor U2246 (N_2246,N_1574,N_19);
nand U2247 (N_2247,N_772,N_1594);
nor U2248 (N_2248,N_307,N_380);
nor U2249 (N_2249,N_644,N_1117);
or U2250 (N_2250,N_1246,N_98);
xnor U2251 (N_2251,N_31,N_363);
or U2252 (N_2252,N_10,N_204);
or U2253 (N_2253,N_596,N_1838);
nor U2254 (N_2254,N_1655,N_1206);
nand U2255 (N_2255,N_86,N_1051);
or U2256 (N_2256,N_288,N_1642);
nand U2257 (N_2257,N_1029,N_1849);
nand U2258 (N_2258,N_339,N_1321);
nand U2259 (N_2259,N_628,N_1829);
nor U2260 (N_2260,N_1093,N_1361);
or U2261 (N_2261,N_821,N_1812);
xnor U2262 (N_2262,N_1703,N_1831);
xor U2263 (N_2263,N_1207,N_1164);
xnor U2264 (N_2264,N_806,N_1921);
nor U2265 (N_2265,N_1987,N_899);
and U2266 (N_2266,N_1416,N_292);
and U2267 (N_2267,N_1220,N_197);
or U2268 (N_2268,N_165,N_96);
and U2269 (N_2269,N_248,N_353);
nor U2270 (N_2270,N_718,N_422);
and U2271 (N_2271,N_631,N_1426);
nand U2272 (N_2272,N_1401,N_885);
nand U2273 (N_2273,N_433,N_1364);
and U2274 (N_2274,N_1256,N_279);
nor U2275 (N_2275,N_1438,N_194);
nor U2276 (N_2276,N_1978,N_51);
nor U2277 (N_2277,N_1226,N_1611);
or U2278 (N_2278,N_1971,N_22);
nand U2279 (N_2279,N_1107,N_515);
or U2280 (N_2280,N_1055,N_1879);
xnor U2281 (N_2281,N_1712,N_76);
nand U2282 (N_2282,N_874,N_695);
nand U2283 (N_2283,N_1081,N_1251);
or U2284 (N_2284,N_182,N_1744);
xnor U2285 (N_2285,N_88,N_1165);
or U2286 (N_2286,N_1242,N_285);
xnor U2287 (N_2287,N_1373,N_1834);
nor U2288 (N_2288,N_657,N_920);
or U2289 (N_2289,N_1391,N_174);
nor U2290 (N_2290,N_221,N_656);
nor U2291 (N_2291,N_1386,N_1780);
or U2292 (N_2292,N_225,N_761);
and U2293 (N_2293,N_1316,N_1866);
nand U2294 (N_2294,N_964,N_1913);
nand U2295 (N_2295,N_1046,N_1253);
xor U2296 (N_2296,N_5,N_1317);
nand U2297 (N_2297,N_980,N_337);
and U2298 (N_2298,N_318,N_77);
and U2299 (N_2299,N_1533,N_510);
nor U2300 (N_2300,N_402,N_1103);
or U2301 (N_2301,N_494,N_506);
nor U2302 (N_2302,N_1129,N_1596);
and U2303 (N_2303,N_183,N_1632);
or U2304 (N_2304,N_595,N_1839);
nor U2305 (N_2305,N_1074,N_1080);
nor U2306 (N_2306,N_157,N_1827);
nor U2307 (N_2307,N_630,N_919);
nor U2308 (N_2308,N_1345,N_375);
nand U2309 (N_2309,N_604,N_1044);
nand U2310 (N_2310,N_838,N_1927);
nor U2311 (N_2311,N_777,N_1751);
and U2312 (N_2312,N_415,N_1696);
nor U2313 (N_2313,N_851,N_1754);
nand U2314 (N_2314,N_391,N_1750);
or U2315 (N_2315,N_1790,N_264);
and U2316 (N_2316,N_1736,N_1499);
or U2317 (N_2317,N_1670,N_490);
nor U2318 (N_2318,N_1895,N_1201);
nor U2319 (N_2319,N_1092,N_588);
nand U2320 (N_2320,N_332,N_1889);
and U2321 (N_2321,N_924,N_302);
nand U2322 (N_2322,N_619,N_744);
or U2323 (N_2323,N_1539,N_1996);
nor U2324 (N_2324,N_107,N_425);
and U2325 (N_2325,N_1232,N_574);
and U2326 (N_2326,N_1393,N_46);
or U2327 (N_2327,N_1094,N_1982);
nand U2328 (N_2328,N_1625,N_1298);
nor U2329 (N_2329,N_1901,N_1943);
or U2330 (N_2330,N_785,N_1558);
or U2331 (N_2331,N_230,N_336);
nand U2332 (N_2332,N_1675,N_1409);
nand U2333 (N_2333,N_63,N_1980);
xnor U2334 (N_2334,N_1118,N_992);
or U2335 (N_2335,N_94,N_411);
or U2336 (N_2336,N_448,N_1639);
nand U2337 (N_2337,N_811,N_764);
nor U2338 (N_2338,N_1371,N_958);
nor U2339 (N_2339,N_314,N_1528);
nand U2340 (N_2340,N_1605,N_799);
or U2341 (N_2341,N_231,N_311);
and U2342 (N_2342,N_1585,N_1564);
nor U2343 (N_2343,N_1312,N_1019);
xor U2344 (N_2344,N_370,N_1709);
xnor U2345 (N_2345,N_724,N_1586);
or U2346 (N_2346,N_1149,N_582);
xnor U2347 (N_2347,N_1707,N_293);
nor U2348 (N_2348,N_193,N_1687);
nand U2349 (N_2349,N_1896,N_1049);
nand U2350 (N_2350,N_580,N_1637);
or U2351 (N_2351,N_846,N_1565);
or U2352 (N_2352,N_847,N_1581);
nor U2353 (N_2353,N_833,N_472);
and U2354 (N_2354,N_281,N_1689);
nor U2355 (N_2355,N_58,N_864);
or U2356 (N_2356,N_912,N_1819);
or U2357 (N_2357,N_1293,N_775);
xor U2358 (N_2358,N_1767,N_1746);
xor U2359 (N_2359,N_1924,N_113);
or U2360 (N_2360,N_599,N_48);
and U2361 (N_2361,N_1169,N_1557);
and U2362 (N_2362,N_849,N_1297);
nand U2363 (N_2363,N_1690,N_1933);
nor U2364 (N_2364,N_684,N_548);
nor U2365 (N_2365,N_809,N_21);
or U2366 (N_2366,N_1571,N_223);
or U2367 (N_2367,N_636,N_1413);
nand U2368 (N_2368,N_814,N_1764);
xnor U2369 (N_2369,N_417,N_441);
or U2370 (N_2370,N_1972,N_715);
and U2371 (N_2371,N_1932,N_926);
and U2372 (N_2372,N_1537,N_1120);
nor U2373 (N_2373,N_1292,N_418);
nor U2374 (N_2374,N_918,N_605);
and U2375 (N_2375,N_71,N_683);
or U2376 (N_2376,N_1857,N_603);
nor U2377 (N_2377,N_414,N_1272);
xor U2378 (N_2378,N_646,N_613);
or U2379 (N_2379,N_389,N_1608);
nor U2380 (N_2380,N_1403,N_1084);
nor U2381 (N_2381,N_1917,N_1257);
nor U2382 (N_2382,N_1470,N_1399);
and U2383 (N_2383,N_825,N_453);
and U2384 (N_2384,N_1089,N_343);
and U2385 (N_2385,N_1825,N_56);
xnor U2386 (N_2386,N_171,N_1423);
or U2387 (N_2387,N_1531,N_305);
or U2388 (N_2388,N_1337,N_623);
nand U2389 (N_2389,N_1483,N_1018);
nand U2390 (N_2390,N_156,N_713);
nor U2391 (N_2391,N_1045,N_1146);
or U2392 (N_2392,N_1148,N_55);
or U2393 (N_2393,N_1192,N_1540);
nor U2394 (N_2394,N_1429,N_568);
or U2395 (N_2395,N_319,N_368);
nor U2396 (N_2396,N_676,N_1052);
nand U2397 (N_2397,N_923,N_246);
nor U2398 (N_2398,N_1225,N_936);
nor U2399 (N_2399,N_1600,N_1593);
nor U2400 (N_2400,N_558,N_1406);
xor U2401 (N_2401,N_1741,N_1347);
and U2402 (N_2402,N_41,N_689);
and U2403 (N_2403,N_812,N_844);
nor U2404 (N_2404,N_962,N_1544);
and U2405 (N_2405,N_994,N_257);
and U2406 (N_2406,N_280,N_1114);
and U2407 (N_2407,N_845,N_1805);
nand U2408 (N_2408,N_1623,N_712);
nor U2409 (N_2409,N_1346,N_808);
xor U2410 (N_2410,N_181,N_578);
xor U2411 (N_2411,N_983,N_752);
and U2412 (N_2412,N_939,N_1739);
or U2413 (N_2413,N_241,N_1359);
xnor U2414 (N_2414,N_1518,N_1479);
nand U2415 (N_2415,N_892,N_933);
nand U2416 (N_2416,N_998,N_524);
and U2417 (N_2417,N_1863,N_813);
nand U2418 (N_2418,N_1633,N_1761);
nor U2419 (N_2419,N_1976,N_451);
nor U2420 (N_2420,N_895,N_999);
and U2421 (N_2421,N_1267,N_650);
nand U2422 (N_2422,N_1458,N_531);
nand U2423 (N_2423,N_913,N_1513);
or U2424 (N_2424,N_296,N_162);
nor U2425 (N_2425,N_1835,N_632);
and U2426 (N_2426,N_942,N_950);
nand U2427 (N_2427,N_1087,N_114);
or U2428 (N_2428,N_1448,N_1659);
xnor U2429 (N_2429,N_164,N_3);
nand U2430 (N_2430,N_716,N_686);
xor U2431 (N_2431,N_253,N_750);
and U2432 (N_2432,N_1323,N_78);
nor U2433 (N_2433,N_817,N_1755);
or U2434 (N_2434,N_1864,N_1283);
and U2435 (N_2435,N_436,N_1275);
and U2436 (N_2436,N_969,N_1266);
nor U2437 (N_2437,N_1090,N_575);
nand U2438 (N_2438,N_1699,N_620);
nor U2439 (N_2439,N_1735,N_639);
and U2440 (N_2440,N_1430,N_1753);
or U2441 (N_2441,N_1521,N_295);
nor U2442 (N_2442,N_1779,N_768);
and U2443 (N_2443,N_1609,N_766);
nor U2444 (N_2444,N_592,N_853);
or U2445 (N_2445,N_381,N_1887);
and U2446 (N_2446,N_34,N_467);
and U2447 (N_2447,N_694,N_459);
nor U2448 (N_2448,N_1388,N_1258);
nand U2449 (N_2449,N_1214,N_1138);
nand U2450 (N_2450,N_1404,N_298);
and U2451 (N_2451,N_1843,N_1453);
and U2452 (N_2452,N_1763,N_1700);
or U2453 (N_2453,N_1119,N_1328);
xnor U2454 (N_2454,N_166,N_294);
and U2455 (N_2455,N_730,N_1204);
nand U2456 (N_2456,N_1714,N_1855);
nand U2457 (N_2457,N_1575,N_1079);
xnor U2458 (N_2458,N_47,N_1579);
or U2459 (N_2459,N_1140,N_1832);
nor U2460 (N_2460,N_1511,N_397);
or U2461 (N_2461,N_929,N_1395);
xor U2462 (N_2462,N_857,N_1407);
or U2463 (N_2463,N_1408,N_1858);
and U2464 (N_2464,N_1840,N_803);
nand U2465 (N_2465,N_1314,N_729);
nand U2466 (N_2466,N_1449,N_1894);
and U2467 (N_2467,N_507,N_14);
nand U2468 (N_2468,N_66,N_8);
xor U2469 (N_2469,N_1014,N_1417);
and U2470 (N_2470,N_1110,N_979);
nor U2471 (N_2471,N_289,N_1749);
nand U2472 (N_2472,N_424,N_1595);
or U2473 (N_2473,N_616,N_553);
nand U2474 (N_2474,N_1387,N_1526);
nor U2475 (N_2475,N_1424,N_151);
or U2476 (N_2476,N_1950,N_1303);
xnor U2477 (N_2477,N_1748,N_444);
and U2478 (N_2478,N_1136,N_781);
nor U2479 (N_2479,N_1854,N_1568);
and U2480 (N_2480,N_1890,N_366);
or U2481 (N_2481,N_1792,N_798);
or U2482 (N_2482,N_1983,N_1447);
xnor U2483 (N_2483,N_555,N_1672);
and U2484 (N_2484,N_317,N_1965);
and U2485 (N_2485,N_228,N_1778);
and U2486 (N_2486,N_1273,N_379);
and U2487 (N_2487,N_740,N_1541);
nor U2488 (N_2488,N_1916,N_247);
and U2489 (N_2489,N_1010,N_1498);
or U2490 (N_2490,N_462,N_593);
nor U2491 (N_2491,N_1178,N_746);
nand U2492 (N_2492,N_1861,N_116);
or U2493 (N_2493,N_890,N_1768);
and U2494 (N_2494,N_430,N_1064);
nand U2495 (N_2495,N_643,N_32);
nor U2496 (N_2496,N_1061,N_1437);
and U2497 (N_2497,N_1504,N_176);
xnor U2498 (N_2498,N_1723,N_434);
nor U2499 (N_2499,N_1654,N_1941);
nor U2500 (N_2500,N_905,N_819);
or U2501 (N_2501,N_190,N_830);
or U2502 (N_2502,N_1477,N_1336);
and U2503 (N_2503,N_1548,N_1125);
nor U2504 (N_2504,N_1322,N_1489);
nand U2505 (N_2505,N_99,N_40);
nor U2506 (N_2506,N_484,N_1951);
and U2507 (N_2507,N_43,N_1195);
nand U2508 (N_2508,N_565,N_818);
nor U2509 (N_2509,N_862,N_473);
xor U2510 (N_2510,N_1553,N_1878);
and U2511 (N_2511,N_1737,N_1296);
and U2512 (N_2512,N_925,N_1166);
nor U2513 (N_2513,N_423,N_1100);
or U2514 (N_2514,N_944,N_27);
nor U2515 (N_2515,N_659,N_1491);
xnor U2516 (N_2516,N_406,N_865);
and U2517 (N_2517,N_1681,N_1847);
or U2518 (N_2518,N_360,N_1115);
and U2519 (N_2519,N_547,N_866);
xor U2520 (N_2520,N_172,N_1874);
nor U2521 (N_2521,N_1197,N_1869);
nand U2522 (N_2522,N_544,N_1508);
or U2523 (N_2523,N_1710,N_661);
and U2524 (N_2524,N_1109,N_1335);
nor U2525 (N_2525,N_1139,N_1196);
nor U2526 (N_2526,N_1038,N_168);
and U2527 (N_2527,N_1543,N_201);
and U2528 (N_2528,N_769,N_1902);
or U2529 (N_2529,N_426,N_374);
nand U2530 (N_2530,N_1493,N_1837);
and U2531 (N_2531,N_299,N_612);
or U2532 (N_2532,N_268,N_1306);
nand U2533 (N_2533,N_1791,N_681);
xnor U2534 (N_2534,N_1069,N_1141);
or U2535 (N_2535,N_263,N_1945);
or U2536 (N_2536,N_1025,N_251);
or U2537 (N_2537,N_1964,N_226);
nor U2538 (N_2538,N_955,N_148);
and U2539 (N_2539,N_1588,N_697);
nand U2540 (N_2540,N_669,N_308);
nor U2541 (N_2541,N_1657,N_1015);
nor U2542 (N_2542,N_1922,N_1584);
or U2543 (N_2543,N_1012,N_771);
xnor U2544 (N_2544,N_736,N_1175);
nor U2545 (N_2545,N_546,N_889);
nor U2546 (N_2546,N_1677,N_1473);
nand U2547 (N_2547,N_1826,N_1787);
or U2548 (N_2548,N_577,N_1476);
xnor U2549 (N_2549,N_930,N_663);
or U2550 (N_2550,N_369,N_710);
or U2551 (N_2551,N_583,N_1066);
or U2552 (N_2552,N_1582,N_439);
and U2553 (N_2553,N_1128,N_780);
nor U2554 (N_2554,N_677,N_1509);
nor U2555 (N_2555,N_1899,N_1510);
nor U2556 (N_2556,N_1130,N_286);
and U2557 (N_2557,N_1075,N_97);
or U2558 (N_2558,N_938,N_1121);
nor U2559 (N_2559,N_1241,N_1357);
or U2560 (N_2560,N_36,N_1963);
nor U2561 (N_2561,N_460,N_340);
nor U2562 (N_2562,N_988,N_270);
and U2563 (N_2563,N_67,N_1621);
and U2564 (N_2564,N_614,N_868);
and U2565 (N_2565,N_100,N_760);
xnor U2566 (N_2566,N_1688,N_1583);
and U2567 (N_2567,N_1760,N_23);
xor U2568 (N_2568,N_1048,N_1648);
nor U2569 (N_2569,N_835,N_1240);
or U2570 (N_2570,N_70,N_1663);
or U2571 (N_2571,N_797,N_1356);
and U2572 (N_2572,N_850,N_1708);
and U2573 (N_2573,N_759,N_719);
or U2574 (N_2574,N_1436,N_881);
and U2575 (N_2575,N_1461,N_1368);
nand U2576 (N_2576,N_1160,N_1142);
or U2577 (N_2577,N_271,N_504);
and U2578 (N_2578,N_997,N_563);
nor U2579 (N_2579,N_1957,N_1154);
or U2580 (N_2580,N_101,N_349);
and U2581 (N_2581,N_1308,N_1280);
nor U2582 (N_2582,N_952,N_1320);
or U2583 (N_2583,N_1309,N_1212);
or U2584 (N_2584,N_260,N_1852);
and U2585 (N_2585,N_1740,N_331);
nor U2586 (N_2586,N_1656,N_522);
nor U2587 (N_2587,N_1372,N_1603);
nor U2588 (N_2588,N_1327,N_1552);
and U2589 (N_2589,N_822,N_126);
nand U2590 (N_2590,N_149,N_348);
nor U2591 (N_2591,N_576,N_1732);
nand U2592 (N_2592,N_236,N_1211);
nor U2593 (N_2593,N_1057,N_987);
and U2594 (N_2594,N_487,N_1216);
nor U2595 (N_2595,N_1072,N_1956);
nor U2596 (N_2596,N_297,N_483);
or U2597 (N_2597,N_129,N_1163);
nand U2598 (N_2598,N_770,N_1122);
and U2599 (N_2599,N_536,N_466);
xnor U2600 (N_2600,N_1718,N_1597);
and U2601 (N_2601,N_242,N_1248);
nand U2602 (N_2602,N_873,N_428);
xnor U2603 (N_2603,N_981,N_62);
or U2604 (N_2604,N_971,N_852);
and U2605 (N_2605,N_1772,N_1463);
or U2606 (N_2606,N_376,N_1098);
or U2607 (N_2607,N_1652,N_791);
xnor U2608 (N_2608,N_606,N_800);
and U2609 (N_2609,N_1747,N_35);
nand U2610 (N_2610,N_1002,N_1188);
nor U2611 (N_2611,N_203,N_961);
or U2612 (N_2612,N_521,N_123);
nor U2613 (N_2613,N_1765,N_1332);
or U2614 (N_2614,N_361,N_1969);
xnor U2615 (N_2615,N_898,N_906);
nor U2616 (N_2616,N_1880,N_1850);
nand U2617 (N_2617,N_787,N_1170);
and U2618 (N_2618,N_1868,N_1668);
or U2619 (N_2619,N_316,N_52);
nor U2620 (N_2620,N_590,N_452);
and U2621 (N_2621,N_1392,N_1135);
or U2622 (N_2622,N_513,N_848);
xor U2623 (N_2623,N_189,N_1083);
and U2624 (N_2624,N_87,N_535);
or U2625 (N_2625,N_877,N_7);
nor U2626 (N_2626,N_691,N_1067);
and U2627 (N_2627,N_909,N_1919);
xor U2628 (N_2628,N_1885,N_670);
or U2629 (N_2629,N_447,N_723);
nand U2630 (N_2630,N_1047,N_674);
xor U2631 (N_2631,N_1276,N_1517);
nand U2632 (N_2632,N_491,N_81);
xor U2633 (N_2633,N_1156,N_75);
nor U2634 (N_2634,N_665,N_1245);
nor U2635 (N_2635,N_882,N_1612);
and U2636 (N_2636,N_202,N_108);
and U2637 (N_2637,N_1848,N_1159);
nand U2638 (N_2638,N_1157,N_1806);
or U2639 (N_2639,N_1456,N_1733);
nand U2640 (N_2640,N_104,N_615);
or U2641 (N_2641,N_1867,N_664);
nor U2642 (N_2642,N_1506,N_329);
or U2643 (N_2643,N_1617,N_668);
nand U2644 (N_2644,N_28,N_461);
nor U2645 (N_2645,N_957,N_1516);
and U2646 (N_2646,N_387,N_1318);
and U2647 (N_2647,N_986,N_1102);
nor U2648 (N_2648,N_1678,N_1907);
nand U2649 (N_2649,N_39,N_93);
xor U2650 (N_2650,N_410,N_1606);
nor U2651 (N_2651,N_1179,N_1865);
nand U2652 (N_2652,N_1906,N_1028);
or U2653 (N_2653,N_721,N_1435);
nor U2654 (N_2654,N_1891,N_1397);
nor U2655 (N_2655,N_1016,N_1006);
nor U2656 (N_2656,N_1823,N_1946);
nand U2657 (N_2657,N_1923,N_1711);
or U2658 (N_2658,N_227,N_445);
nor U2659 (N_2659,N_141,N_1682);
xor U2660 (N_2660,N_792,N_1349);
nand U2661 (N_2661,N_493,N_1131);
nand U2662 (N_2662,N_1589,N_1264);
and U2663 (N_2663,N_1602,N_1570);
nand U2664 (N_2664,N_519,N_523);
or U2665 (N_2665,N_1693,N_543);
xor U2666 (N_2666,N_160,N_1198);
nor U2667 (N_2667,N_561,N_827);
xor U2668 (N_2668,N_303,N_1354);
and U2669 (N_2669,N_372,N_1591);
nor U2670 (N_2670,N_356,N_175);
xor U2671 (N_2671,N_700,N_1180);
and U2672 (N_2672,N_1715,N_641);
or U2673 (N_2673,N_1729,N_1944);
or U2674 (N_2674,N_1882,N_1846);
nand U2675 (N_2675,N_350,N_117);
and U2676 (N_2676,N_820,N_1344);
xor U2677 (N_2677,N_1886,N_267);
nand U2678 (N_2678,N_1099,N_1520);
nand U2679 (N_2679,N_880,N_1635);
nand U2680 (N_2680,N_133,N_477);
or U2681 (N_2681,N_1302,N_1271);
nor U2682 (N_2682,N_128,N_1106);
or U2683 (N_2683,N_1071,N_345);
or U2684 (N_2684,N_159,N_532);
xnor U2685 (N_2685,N_1496,N_1795);
or U2686 (N_2686,N_959,N_1631);
xnor U2687 (N_2687,N_1492,N_581);
nor U2688 (N_2688,N_212,N_401);
xnor U2689 (N_2689,N_282,N_18);
xnor U2690 (N_2690,N_469,N_45);
nor U2691 (N_2691,N_1929,N_481);
xnor U2692 (N_2692,N_239,N_1008);
or U2693 (N_2693,N_20,N_102);
nand U2694 (N_2694,N_982,N_153);
nand U2695 (N_2695,N_1182,N_1343);
or U2696 (N_2696,N_888,N_458);
nand U2697 (N_2697,N_1551,N_533);
or U2698 (N_2698,N_840,N_1897);
or U2699 (N_2699,N_1153,N_1333);
xor U2700 (N_2700,N_1062,N_1762);
or U2701 (N_2701,N_698,N_573);
nor U2702 (N_2702,N_1450,N_1431);
nand U2703 (N_2703,N_1017,N_334);
or U2704 (N_2704,N_635,N_135);
or U2705 (N_2705,N_1782,N_64);
and U2706 (N_2706,N_1722,N_793);
or U2707 (N_2707,N_667,N_1726);
nand U2708 (N_2708,N_922,N_916);
or U2709 (N_2709,N_265,N_585);
nand U2710 (N_2710,N_1021,N_738);
or U2711 (N_2711,N_1949,N_517);
and U2712 (N_2712,N_1305,N_1465);
and U2713 (N_2713,N_399,N_405);
xnor U2714 (N_2714,N_198,N_1127);
nand U2715 (N_2715,N_82,N_1147);
or U2716 (N_2716,N_843,N_638);
xor U2717 (N_2717,N_607,N_642);
and U2718 (N_2718,N_1813,N_416);
nand U2719 (N_2719,N_456,N_1664);
nand U2720 (N_2720,N_1940,N_917);
and U2721 (N_2721,N_1636,N_570);
and U2722 (N_2722,N_106,N_1967);
or U2723 (N_2723,N_1460,N_611);
nand U2724 (N_2724,N_972,N_618);
xor U2725 (N_2725,N_1628,N_1301);
nand U2726 (N_2726,N_1410,N_1752);
xor U2727 (N_2727,N_1519,N_53);
nand U2728 (N_2728,N_779,N_1176);
or U2729 (N_2729,N_702,N_1542);
nand U2730 (N_2730,N_1235,N_1034);
or U2731 (N_2731,N_1375,N_754);
or U2732 (N_2732,N_1734,N_1277);
nand U2733 (N_2733,N_1167,N_1338);
and U2734 (N_2734,N_1559,N_1348);
and U2735 (N_2735,N_887,N_11);
nand U2736 (N_2736,N_1155,N_1068);
or U2737 (N_2737,N_1500,N_25);
or U2738 (N_2738,N_427,N_1362);
nor U2739 (N_2739,N_914,N_124);
and U2740 (N_2740,N_525,N_976);
and U2741 (N_2741,N_304,N_498);
nor U2742 (N_2742,N_150,N_855);
and U2743 (N_2743,N_571,N_1036);
nor U2744 (N_2744,N_1914,N_1279);
or U2745 (N_2745,N_1313,N_662);
nor U2746 (N_2746,N_1295,N_1382);
and U2747 (N_2747,N_796,N_1290);
nand U2748 (N_2748,N_624,N_756);
or U2749 (N_2749,N_900,N_1973);
nand U2750 (N_2750,N_209,N_860);
nor U2751 (N_2751,N_1507,N_1975);
nor U2752 (N_2752,N_1985,N_1873);
and U2753 (N_2753,N_449,N_1350);
xor U2754 (N_2754,N_1384,N_1020);
xor U2755 (N_2755,N_130,N_1270);
nor U2756 (N_2756,N_233,N_1208);
nand U2757 (N_2757,N_707,N_73);
or U2758 (N_2758,N_1758,N_1494);
nor U2759 (N_2759,N_210,N_57);
nor U2760 (N_2760,N_1011,N_968);
nor U2761 (N_2761,N_139,N_480);
and U2762 (N_2762,N_1227,N_254);
nor U2763 (N_2763,N_1451,N_989);
nor U2764 (N_2764,N_751,N_529);
or U2765 (N_2765,N_1501,N_1884);
xor U2766 (N_2766,N_13,N_465);
nor U2767 (N_2767,N_1515,N_105);
or U2768 (N_2768,N_876,N_1638);
or U2769 (N_2769,N_1771,N_863);
xor U2770 (N_2770,N_400,N_1215);
nand U2771 (N_2771,N_68,N_1522);
or U2772 (N_2772,N_1691,N_564);
nor U2773 (N_2773,N_1353,N_810);
xnor U2774 (N_2774,N_192,N_1797);
xor U2775 (N_2775,N_1803,N_1799);
xnor U2776 (N_2776,N_1223,N_1474);
and U2777 (N_2777,N_1578,N_500);
nand U2778 (N_2778,N_1577,N_666);
or U2779 (N_2779,N_413,N_725);
nor U2780 (N_2780,N_699,N_1239);
xor U2781 (N_2781,N_1471,N_1997);
nor U2782 (N_2782,N_1883,N_1383);
or U2783 (N_2783,N_92,N_649);
nand U2784 (N_2784,N_586,N_74);
nor U2785 (N_2785,N_541,N_1274);
nor U2786 (N_2786,N_562,N_358);
or U2787 (N_2787,N_1822,N_6);
and U2788 (N_2788,N_839,N_503);
nor U2789 (N_2789,N_1026,N_38);
xnor U2790 (N_2790,N_1872,N_634);
and U2791 (N_2791,N_1374,N_834);
and U2792 (N_2792,N_935,N_1836);
or U2793 (N_2793,N_692,N_177);
or U2794 (N_2794,N_1853,N_1482);
nor U2795 (N_2795,N_1994,N_1538);
nand U2796 (N_2796,N_1900,N_1340);
xor U2797 (N_2797,N_1097,N_1365);
and U2798 (N_2798,N_1770,N_1459);
and U2799 (N_2799,N_1989,N_1942);
nor U2800 (N_2800,N_258,N_1132);
or U2801 (N_2801,N_883,N_144);
nand U2802 (N_2802,N_138,N_941);
and U2803 (N_2803,N_1042,N_1229);
and U2804 (N_2804,N_904,N_147);
or U2805 (N_2805,N_1743,N_1818);
and U2806 (N_2806,N_948,N_1411);
or U2807 (N_2807,N_690,N_232);
or U2808 (N_2808,N_861,N_383);
and U2809 (N_2809,N_762,N_1076);
nand U2810 (N_2810,N_1992,N_1999);
nor U2811 (N_2811,N_335,N_1056);
nand U2812 (N_2812,N_621,N_1870);
nand U2813 (N_2813,N_1860,N_1624);
nor U2814 (N_2814,N_111,N_622);
nor U2815 (N_2815,N_1995,N_1727);
nor U2816 (N_2816,N_95,N_386);
nor U2817 (N_2817,N_967,N_435);
xnor U2818 (N_2818,N_367,N_1105);
xor U2819 (N_2819,N_1794,N_30);
nand U2820 (N_2820,N_842,N_1070);
xor U2821 (N_2821,N_1108,N_871);
and U2822 (N_2822,N_1694,N_1851);
nand U2823 (N_2823,N_1039,N_1412);
nor U2824 (N_2824,N_1202,N_1673);
xor U2825 (N_2825,N_136,N_1441);
or U2826 (N_2826,N_567,N_240);
nor U2827 (N_2827,N_1315,N_152);
or U2828 (N_2828,N_1415,N_706);
nor U2829 (N_2829,N_514,N_1116);
nand U2830 (N_2830,N_1954,N_1329);
nand U2831 (N_2831,N_516,N_437);
nand U2832 (N_2832,N_1486,N_1833);
nor U2833 (N_2833,N_1440,N_1862);
nand U2834 (N_2834,N_801,N_1191);
and U2835 (N_2835,N_185,N_966);
nand U2836 (N_2836,N_502,N_1189);
nand U2837 (N_2837,N_837,N_1381);
or U2838 (N_2838,N_908,N_262);
xnor U2839 (N_2839,N_1444,N_1497);
nand U2840 (N_2840,N_1024,N_341);
and U2841 (N_2841,N_1573,N_1634);
nand U2842 (N_2842,N_475,N_1935);
nor U2843 (N_2843,N_273,N_1881);
or U2844 (N_2844,N_1360,N_1433);
and U2845 (N_2845,N_1380,N_778);
and U2846 (N_2846,N_854,N_1355);
or U2847 (N_2847,N_394,N_1828);
or U2848 (N_2848,N_520,N_215);
and U2849 (N_2849,N_219,N_505);
nor U2850 (N_2850,N_722,N_609);
xor U2851 (N_2851,N_1053,N_1035);
nand U2852 (N_2852,N_1455,N_728);
or U2853 (N_2853,N_551,N_566);
and U2854 (N_2854,N_1040,N_1265);
and U2855 (N_2855,N_158,N_1802);
nor U2856 (N_2856,N_1619,N_658);
nor U2857 (N_2857,N_678,N_1033);
nand U2858 (N_2858,N_431,N_526);
or U2859 (N_2859,N_1261,N_69);
or U2860 (N_2860,N_617,N_1177);
or U2861 (N_2861,N_408,N_1627);
and U2862 (N_2862,N_488,N_539);
and U2863 (N_2863,N_518,N_1331);
xor U2864 (N_2864,N_747,N_284);
and U2865 (N_2865,N_290,N_1278);
nor U2866 (N_2866,N_213,N_1550);
or U2867 (N_2867,N_393,N_805);
or U2868 (N_2868,N_392,N_1549);
nor U2869 (N_2869,N_587,N_931);
nor U2870 (N_2870,N_196,N_1667);
nor U2871 (N_2871,N_1095,N_1660);
and U2872 (N_2872,N_1490,N_708);
and U2873 (N_2873,N_673,N_1200);
and U2874 (N_2874,N_907,N_1352);
or U2875 (N_2875,N_1376,N_167);
or U2876 (N_2876,N_978,N_1502);
nor U2877 (N_2877,N_629,N_1810);
nand U2878 (N_2878,N_1063,N_1911);
nor U2879 (N_2879,N_359,N_1414);
nand U2880 (N_2880,N_338,N_1815);
nor U2881 (N_2881,N_421,N_501);
nor U2882 (N_2882,N_841,N_1679);
or U2883 (N_2883,N_1367,N_1563);
nand U2884 (N_2884,N_1674,N_486);
nor U2885 (N_2885,N_1546,N_915);
nand U2886 (N_2886,N_1060,N_1793);
nand U2887 (N_2887,N_1254,N_499);
nor U2888 (N_2888,N_858,N_277);
xor U2889 (N_2889,N_205,N_476);
or U2890 (N_2890,N_511,N_1104);
nand U2891 (N_2891,N_633,N_1716);
and U2892 (N_2892,N_269,N_61);
nor U2893 (N_2893,N_1339,N_208);
or U2894 (N_2894,N_250,N_1993);
nand U2895 (N_2895,N_601,N_1124);
nand U2896 (N_2896,N_310,N_789);
or U2897 (N_2897,N_1342,N_1697);
nor U2898 (N_2898,N_1821,N_714);
and U2899 (N_2899,N_218,N_222);
nor U2900 (N_2900,N_1043,N_50);
nand U2901 (N_2901,N_140,N_357);
nand U2902 (N_2902,N_1205,N_963);
and U2903 (N_2903,N_742,N_1918);
xnor U2904 (N_2904,N_696,N_1086);
nor U2905 (N_2905,N_1420,N_1844);
nor U2906 (N_2906,N_1238,N_195);
nor U2907 (N_2907,N_1525,N_557);
nand U2908 (N_2908,N_1193,N_1101);
nor U2909 (N_2909,N_1936,N_1545);
or U2910 (N_2910,N_1998,N_1824);
and U2911 (N_2911,N_378,N_1389);
xor U2912 (N_2912,N_654,N_1199);
nand U2913 (N_2913,N_1702,N_1369);
nand U2914 (N_2914,N_594,N_1658);
and U2915 (N_2915,N_1091,N_783);
nor U2916 (N_2916,N_1986,N_1082);
nand U2917 (N_2917,N_1085,N_1217);
nand U2918 (N_2918,N_1599,N_902);
and U2919 (N_2919,N_313,N_1562);
nand U2920 (N_2920,N_1488,N_741);
xor U2921 (N_2921,N_734,N_121);
or U2922 (N_2922,N_859,N_984);
nand U2923 (N_2923,N_1096,N_301);
and U2924 (N_2924,N_717,N_1629);
or U2925 (N_2925,N_1310,N_589);
nand U2926 (N_2926,N_645,N_727);
and U2927 (N_2927,N_1268,N_1908);
nor U2928 (N_2928,N_1480,N_1481);
or U2929 (N_2929,N_1587,N_1990);
nand U2930 (N_2930,N_1228,N_1419);
nor U2931 (N_2931,N_675,N_743);
xnor U2932 (N_2932,N_1959,N_679);
or U2933 (N_2933,N_1000,N_996);
nand U2934 (N_2934,N_993,N_1282);
or U2935 (N_2935,N_1467,N_1394);
and U2936 (N_2936,N_970,N_1871);
nor U2937 (N_2937,N_1126,N_1610);
and U2938 (N_2938,N_829,N_928);
and U2939 (N_2939,N_214,N_816);
nor U2940 (N_2940,N_403,N_704);
nand U2941 (N_2941,N_1926,N_1311);
and U2942 (N_2942,N_1662,N_16);
or U2943 (N_2943,N_804,N_1210);
or U2944 (N_2944,N_745,N_1484);
nor U2945 (N_2945,N_735,N_199);
nand U2946 (N_2946,N_79,N_1859);
nor U2947 (N_2947,N_255,N_450);
nor U2948 (N_2948,N_347,N_266);
and U2949 (N_2949,N_1184,N_495);
nand U2950 (N_2950,N_33,N_1653);
nand U2951 (N_2951,N_173,N_365);
nor U2952 (N_2952,N_1181,N_1777);
nand U2953 (N_2953,N_921,N_1234);
xor U2954 (N_2954,N_1561,N_83);
or U2955 (N_2955,N_569,N_1190);
or U2956 (N_2956,N_342,N_479);
or U2957 (N_2957,N_1446,N_351);
nand U2958 (N_2958,N_869,N_1503);
nor U2959 (N_2959,N_672,N_549);
or U2960 (N_2960,N_1123,N_1604);
nor U2961 (N_2961,N_1422,N_1370);
nand U2962 (N_2962,N_291,N_965);
nor U2963 (N_2963,N_552,N_1962);
nand U2964 (N_2964,N_894,N_554);
nor U2965 (N_2965,N_1620,N_1686);
nor U2966 (N_2966,N_17,N_244);
or U2967 (N_2967,N_1005,N_1243);
nor U2968 (N_2968,N_60,N_463);
nand U2969 (N_2969,N_1,N_432);
nand U2970 (N_2970,N_249,N_1665);
and U2971 (N_2971,N_671,N_956);
nor U2972 (N_2972,N_1529,N_1145);
xor U2973 (N_2973,N_1704,N_1569);
and U2974 (N_2974,N_550,N_1626);
nor U2975 (N_2975,N_1692,N_1203);
nand U2976 (N_2976,N_1888,N_685);
and U2977 (N_2977,N_911,N_1547);
and U2978 (N_2978,N_84,N_856);
nor U2979 (N_2979,N_1221,N_954);
nand U2980 (N_2980,N_438,N_802);
xnor U2981 (N_2981,N_1925,N_2);
nor U2982 (N_2982,N_795,N_1186);
nand U2983 (N_2983,N_773,N_1378);
nor U2984 (N_2984,N_1646,N_1904);
nor U2985 (N_2985,N_757,N_44);
and U2986 (N_2986,N_1730,N_1158);
nor U2987 (N_2987,N_537,N_1898);
nor U2988 (N_2988,N_1970,N_627);
or U2989 (N_2989,N_1259,N_29);
and U2990 (N_2990,N_910,N_1291);
nor U2991 (N_2991,N_637,N_355);
or U2992 (N_2992,N_245,N_1979);
and U2993 (N_2993,N_1288,N_870);
or U2994 (N_2994,N_1294,N_1816);
and U2995 (N_2995,N_407,N_1698);
xnor U2996 (N_2996,N_492,N_1530);
nand U2997 (N_2997,N_572,N_1775);
or U2998 (N_2998,N_1512,N_384);
and U2999 (N_2999,N_364,N_186);
nand U3000 (N_3000,N_714,N_1750);
xnor U3001 (N_3001,N_99,N_1415);
nor U3002 (N_3002,N_1070,N_862);
and U3003 (N_3003,N_1410,N_683);
nor U3004 (N_3004,N_1694,N_54);
nor U3005 (N_3005,N_1534,N_964);
and U3006 (N_3006,N_672,N_399);
nand U3007 (N_3007,N_1686,N_1576);
nand U3008 (N_3008,N_1344,N_1699);
nor U3009 (N_3009,N_675,N_1060);
or U3010 (N_3010,N_1107,N_71);
and U3011 (N_3011,N_804,N_1135);
or U3012 (N_3012,N_1890,N_1442);
nand U3013 (N_3013,N_1897,N_190);
and U3014 (N_3014,N_570,N_305);
nand U3015 (N_3015,N_965,N_200);
nand U3016 (N_3016,N_1806,N_577);
xnor U3017 (N_3017,N_507,N_940);
and U3018 (N_3018,N_1362,N_127);
xor U3019 (N_3019,N_1239,N_1730);
and U3020 (N_3020,N_1922,N_1799);
and U3021 (N_3021,N_148,N_1682);
xnor U3022 (N_3022,N_1909,N_1545);
or U3023 (N_3023,N_258,N_1133);
or U3024 (N_3024,N_1076,N_1321);
nand U3025 (N_3025,N_744,N_976);
and U3026 (N_3026,N_1781,N_1022);
and U3027 (N_3027,N_403,N_1654);
nor U3028 (N_3028,N_54,N_1241);
and U3029 (N_3029,N_1711,N_462);
and U3030 (N_3030,N_838,N_448);
xnor U3031 (N_3031,N_969,N_856);
nand U3032 (N_3032,N_918,N_382);
and U3033 (N_3033,N_183,N_146);
nand U3034 (N_3034,N_1771,N_545);
nand U3035 (N_3035,N_1865,N_322);
nand U3036 (N_3036,N_110,N_59);
nand U3037 (N_3037,N_299,N_925);
nand U3038 (N_3038,N_1615,N_1992);
and U3039 (N_3039,N_667,N_688);
or U3040 (N_3040,N_743,N_893);
or U3041 (N_3041,N_1068,N_1872);
and U3042 (N_3042,N_1644,N_1853);
and U3043 (N_3043,N_342,N_1917);
or U3044 (N_3044,N_1228,N_315);
or U3045 (N_3045,N_1772,N_87);
nor U3046 (N_3046,N_1758,N_1098);
and U3047 (N_3047,N_332,N_275);
xor U3048 (N_3048,N_585,N_1732);
nor U3049 (N_3049,N_618,N_1979);
nand U3050 (N_3050,N_105,N_502);
xor U3051 (N_3051,N_1909,N_876);
nor U3052 (N_3052,N_1734,N_490);
nand U3053 (N_3053,N_195,N_924);
nor U3054 (N_3054,N_1814,N_977);
and U3055 (N_3055,N_1936,N_126);
xor U3056 (N_3056,N_3,N_1100);
or U3057 (N_3057,N_461,N_1662);
nor U3058 (N_3058,N_1091,N_823);
xnor U3059 (N_3059,N_584,N_346);
xnor U3060 (N_3060,N_1611,N_1361);
nor U3061 (N_3061,N_738,N_941);
xnor U3062 (N_3062,N_1923,N_1435);
and U3063 (N_3063,N_5,N_1733);
nand U3064 (N_3064,N_573,N_389);
or U3065 (N_3065,N_446,N_58);
nor U3066 (N_3066,N_1635,N_1003);
nor U3067 (N_3067,N_153,N_1826);
nor U3068 (N_3068,N_1928,N_297);
nand U3069 (N_3069,N_1424,N_12);
and U3070 (N_3070,N_357,N_229);
and U3071 (N_3071,N_609,N_1323);
and U3072 (N_3072,N_329,N_1657);
nor U3073 (N_3073,N_1829,N_20);
and U3074 (N_3074,N_1027,N_1672);
or U3075 (N_3075,N_469,N_145);
xnor U3076 (N_3076,N_530,N_1769);
or U3077 (N_3077,N_1583,N_1316);
nor U3078 (N_3078,N_354,N_1358);
nand U3079 (N_3079,N_415,N_1491);
nand U3080 (N_3080,N_899,N_1563);
xnor U3081 (N_3081,N_17,N_1517);
nand U3082 (N_3082,N_1549,N_1179);
or U3083 (N_3083,N_1639,N_1591);
and U3084 (N_3084,N_1348,N_1433);
nand U3085 (N_3085,N_1073,N_132);
nor U3086 (N_3086,N_1617,N_1988);
nor U3087 (N_3087,N_1632,N_422);
or U3088 (N_3088,N_1859,N_649);
or U3089 (N_3089,N_1177,N_189);
and U3090 (N_3090,N_1277,N_670);
nor U3091 (N_3091,N_1882,N_577);
or U3092 (N_3092,N_1835,N_1200);
or U3093 (N_3093,N_1642,N_933);
nand U3094 (N_3094,N_1282,N_1198);
nand U3095 (N_3095,N_996,N_976);
and U3096 (N_3096,N_1245,N_1602);
nor U3097 (N_3097,N_1085,N_88);
and U3098 (N_3098,N_300,N_890);
and U3099 (N_3099,N_252,N_1068);
nor U3100 (N_3100,N_377,N_500);
nor U3101 (N_3101,N_1519,N_587);
xnor U3102 (N_3102,N_621,N_1648);
nand U3103 (N_3103,N_183,N_277);
nor U3104 (N_3104,N_176,N_1313);
xnor U3105 (N_3105,N_1164,N_4);
xor U3106 (N_3106,N_1938,N_145);
nor U3107 (N_3107,N_804,N_1044);
or U3108 (N_3108,N_92,N_1492);
and U3109 (N_3109,N_39,N_753);
nor U3110 (N_3110,N_1874,N_1372);
nor U3111 (N_3111,N_927,N_390);
nor U3112 (N_3112,N_161,N_1538);
xor U3113 (N_3113,N_1838,N_289);
and U3114 (N_3114,N_814,N_1761);
xnor U3115 (N_3115,N_668,N_571);
xnor U3116 (N_3116,N_1771,N_404);
xnor U3117 (N_3117,N_745,N_239);
and U3118 (N_3118,N_832,N_1655);
nand U3119 (N_3119,N_1151,N_417);
and U3120 (N_3120,N_1631,N_1521);
and U3121 (N_3121,N_41,N_978);
nor U3122 (N_3122,N_718,N_717);
nor U3123 (N_3123,N_484,N_731);
nand U3124 (N_3124,N_1899,N_912);
and U3125 (N_3125,N_413,N_883);
or U3126 (N_3126,N_1199,N_260);
and U3127 (N_3127,N_1366,N_246);
nand U3128 (N_3128,N_540,N_765);
nand U3129 (N_3129,N_985,N_821);
nand U3130 (N_3130,N_796,N_299);
or U3131 (N_3131,N_729,N_124);
nor U3132 (N_3132,N_670,N_1751);
and U3133 (N_3133,N_490,N_644);
or U3134 (N_3134,N_801,N_250);
and U3135 (N_3135,N_1597,N_82);
nor U3136 (N_3136,N_1407,N_1989);
nor U3137 (N_3137,N_1532,N_1919);
nand U3138 (N_3138,N_1404,N_623);
nor U3139 (N_3139,N_1161,N_1682);
nor U3140 (N_3140,N_733,N_1054);
nor U3141 (N_3141,N_611,N_1499);
or U3142 (N_3142,N_243,N_1189);
nand U3143 (N_3143,N_1745,N_1496);
nand U3144 (N_3144,N_1133,N_996);
nor U3145 (N_3145,N_157,N_1785);
and U3146 (N_3146,N_1336,N_1120);
and U3147 (N_3147,N_340,N_367);
nor U3148 (N_3148,N_513,N_431);
and U3149 (N_3149,N_852,N_637);
xor U3150 (N_3150,N_1038,N_1851);
nand U3151 (N_3151,N_1571,N_1124);
and U3152 (N_3152,N_1521,N_761);
or U3153 (N_3153,N_301,N_1743);
or U3154 (N_3154,N_923,N_197);
nand U3155 (N_3155,N_333,N_12);
nor U3156 (N_3156,N_365,N_1021);
and U3157 (N_3157,N_1004,N_1241);
nor U3158 (N_3158,N_189,N_516);
nor U3159 (N_3159,N_1436,N_275);
nor U3160 (N_3160,N_204,N_730);
nor U3161 (N_3161,N_1010,N_639);
xor U3162 (N_3162,N_1273,N_1387);
and U3163 (N_3163,N_805,N_1502);
nand U3164 (N_3164,N_200,N_1815);
xnor U3165 (N_3165,N_1502,N_491);
and U3166 (N_3166,N_1992,N_1755);
and U3167 (N_3167,N_918,N_1180);
nor U3168 (N_3168,N_163,N_611);
and U3169 (N_3169,N_702,N_1649);
and U3170 (N_3170,N_1851,N_656);
nand U3171 (N_3171,N_666,N_1724);
and U3172 (N_3172,N_1993,N_1888);
nor U3173 (N_3173,N_1615,N_1947);
nor U3174 (N_3174,N_1888,N_1518);
nor U3175 (N_3175,N_166,N_1259);
and U3176 (N_3176,N_559,N_669);
nand U3177 (N_3177,N_421,N_1625);
nor U3178 (N_3178,N_1180,N_403);
or U3179 (N_3179,N_976,N_1025);
nor U3180 (N_3180,N_1558,N_341);
nor U3181 (N_3181,N_1895,N_1128);
nor U3182 (N_3182,N_1195,N_611);
or U3183 (N_3183,N_1167,N_1501);
nand U3184 (N_3184,N_1598,N_1799);
and U3185 (N_3185,N_1137,N_635);
xor U3186 (N_3186,N_236,N_1877);
and U3187 (N_3187,N_930,N_842);
or U3188 (N_3188,N_1647,N_1363);
nand U3189 (N_3189,N_1049,N_1830);
nor U3190 (N_3190,N_1125,N_1179);
or U3191 (N_3191,N_303,N_1054);
and U3192 (N_3192,N_1758,N_1545);
or U3193 (N_3193,N_1121,N_886);
nand U3194 (N_3194,N_1606,N_844);
nor U3195 (N_3195,N_943,N_463);
or U3196 (N_3196,N_1826,N_577);
nor U3197 (N_3197,N_1713,N_713);
or U3198 (N_3198,N_196,N_1371);
nor U3199 (N_3199,N_804,N_1586);
nand U3200 (N_3200,N_278,N_678);
nor U3201 (N_3201,N_1132,N_187);
nand U3202 (N_3202,N_1988,N_934);
nor U3203 (N_3203,N_1043,N_437);
nand U3204 (N_3204,N_1424,N_1583);
and U3205 (N_3205,N_1310,N_1857);
nor U3206 (N_3206,N_1575,N_979);
nand U3207 (N_3207,N_1227,N_1429);
xnor U3208 (N_3208,N_859,N_391);
xnor U3209 (N_3209,N_1680,N_1429);
xor U3210 (N_3210,N_733,N_1260);
nand U3211 (N_3211,N_1809,N_1968);
xor U3212 (N_3212,N_425,N_621);
and U3213 (N_3213,N_728,N_226);
or U3214 (N_3214,N_687,N_669);
xnor U3215 (N_3215,N_1364,N_197);
nor U3216 (N_3216,N_364,N_1227);
and U3217 (N_3217,N_1380,N_1791);
nand U3218 (N_3218,N_1408,N_810);
nor U3219 (N_3219,N_338,N_290);
xor U3220 (N_3220,N_348,N_1183);
and U3221 (N_3221,N_894,N_365);
nor U3222 (N_3222,N_557,N_237);
nor U3223 (N_3223,N_691,N_1985);
and U3224 (N_3224,N_1946,N_819);
xor U3225 (N_3225,N_854,N_247);
and U3226 (N_3226,N_1086,N_532);
xor U3227 (N_3227,N_268,N_1397);
and U3228 (N_3228,N_106,N_988);
and U3229 (N_3229,N_505,N_1060);
nand U3230 (N_3230,N_23,N_1601);
and U3231 (N_3231,N_236,N_805);
or U3232 (N_3232,N_31,N_1083);
nand U3233 (N_3233,N_1600,N_816);
nand U3234 (N_3234,N_1726,N_1367);
nand U3235 (N_3235,N_1624,N_1229);
and U3236 (N_3236,N_802,N_1902);
xor U3237 (N_3237,N_293,N_1164);
or U3238 (N_3238,N_998,N_482);
or U3239 (N_3239,N_1995,N_768);
nor U3240 (N_3240,N_1813,N_414);
nor U3241 (N_3241,N_1432,N_63);
nand U3242 (N_3242,N_1049,N_1286);
nand U3243 (N_3243,N_705,N_840);
nand U3244 (N_3244,N_1235,N_1821);
nand U3245 (N_3245,N_602,N_66);
xor U3246 (N_3246,N_1014,N_1658);
or U3247 (N_3247,N_1532,N_1109);
nand U3248 (N_3248,N_633,N_26);
nor U3249 (N_3249,N_567,N_1164);
and U3250 (N_3250,N_796,N_1617);
and U3251 (N_3251,N_1727,N_422);
nand U3252 (N_3252,N_1592,N_901);
nand U3253 (N_3253,N_929,N_1753);
nand U3254 (N_3254,N_515,N_970);
or U3255 (N_3255,N_1097,N_1427);
and U3256 (N_3256,N_116,N_785);
or U3257 (N_3257,N_1368,N_1962);
and U3258 (N_3258,N_1629,N_293);
or U3259 (N_3259,N_515,N_1229);
nor U3260 (N_3260,N_1973,N_1708);
nand U3261 (N_3261,N_1484,N_847);
nor U3262 (N_3262,N_851,N_208);
nor U3263 (N_3263,N_221,N_362);
and U3264 (N_3264,N_13,N_1137);
xnor U3265 (N_3265,N_1656,N_1446);
and U3266 (N_3266,N_936,N_1545);
or U3267 (N_3267,N_1513,N_1281);
nand U3268 (N_3268,N_169,N_1954);
nand U3269 (N_3269,N_1294,N_1477);
nor U3270 (N_3270,N_65,N_170);
nor U3271 (N_3271,N_566,N_707);
nor U3272 (N_3272,N_328,N_1519);
and U3273 (N_3273,N_1043,N_1800);
and U3274 (N_3274,N_1160,N_564);
and U3275 (N_3275,N_1762,N_1429);
nand U3276 (N_3276,N_1153,N_471);
or U3277 (N_3277,N_305,N_1691);
nor U3278 (N_3278,N_1413,N_442);
and U3279 (N_3279,N_459,N_1595);
nor U3280 (N_3280,N_1988,N_966);
or U3281 (N_3281,N_179,N_1615);
and U3282 (N_3282,N_1581,N_1658);
nand U3283 (N_3283,N_1623,N_1387);
or U3284 (N_3284,N_1454,N_1301);
nand U3285 (N_3285,N_1794,N_1809);
and U3286 (N_3286,N_1429,N_190);
nand U3287 (N_3287,N_1637,N_323);
or U3288 (N_3288,N_510,N_894);
or U3289 (N_3289,N_227,N_314);
nor U3290 (N_3290,N_1111,N_1356);
or U3291 (N_3291,N_1169,N_1150);
or U3292 (N_3292,N_1200,N_1161);
nor U3293 (N_3293,N_703,N_1882);
and U3294 (N_3294,N_1351,N_451);
or U3295 (N_3295,N_1061,N_978);
and U3296 (N_3296,N_416,N_898);
nor U3297 (N_3297,N_432,N_333);
and U3298 (N_3298,N_145,N_370);
xor U3299 (N_3299,N_1860,N_604);
and U3300 (N_3300,N_1771,N_241);
nor U3301 (N_3301,N_236,N_1130);
and U3302 (N_3302,N_1912,N_1852);
and U3303 (N_3303,N_700,N_1165);
or U3304 (N_3304,N_1091,N_1337);
and U3305 (N_3305,N_543,N_778);
nor U3306 (N_3306,N_1199,N_1539);
nand U3307 (N_3307,N_1684,N_632);
nand U3308 (N_3308,N_804,N_694);
nor U3309 (N_3309,N_873,N_1797);
xnor U3310 (N_3310,N_972,N_1070);
xor U3311 (N_3311,N_208,N_1279);
nor U3312 (N_3312,N_1846,N_753);
nor U3313 (N_3313,N_1607,N_1268);
nor U3314 (N_3314,N_1044,N_1261);
nor U3315 (N_3315,N_151,N_1873);
nand U3316 (N_3316,N_449,N_808);
or U3317 (N_3317,N_1428,N_1756);
nand U3318 (N_3318,N_1619,N_102);
nor U3319 (N_3319,N_1663,N_766);
and U3320 (N_3320,N_771,N_1251);
nand U3321 (N_3321,N_528,N_1435);
or U3322 (N_3322,N_1086,N_1423);
nor U3323 (N_3323,N_1700,N_878);
or U3324 (N_3324,N_54,N_1963);
and U3325 (N_3325,N_1264,N_78);
xnor U3326 (N_3326,N_1561,N_285);
and U3327 (N_3327,N_1664,N_232);
nand U3328 (N_3328,N_350,N_1794);
and U3329 (N_3329,N_1792,N_1677);
nand U3330 (N_3330,N_1770,N_238);
xor U3331 (N_3331,N_917,N_730);
nand U3332 (N_3332,N_271,N_1544);
and U3333 (N_3333,N_1261,N_121);
nor U3334 (N_3334,N_951,N_1079);
and U3335 (N_3335,N_633,N_308);
and U3336 (N_3336,N_61,N_1129);
nor U3337 (N_3337,N_1247,N_856);
nor U3338 (N_3338,N_1256,N_1869);
xnor U3339 (N_3339,N_377,N_1739);
and U3340 (N_3340,N_1140,N_1551);
or U3341 (N_3341,N_1623,N_1734);
or U3342 (N_3342,N_1885,N_1902);
and U3343 (N_3343,N_15,N_1108);
nand U3344 (N_3344,N_1485,N_1015);
or U3345 (N_3345,N_638,N_1722);
and U3346 (N_3346,N_1513,N_1309);
or U3347 (N_3347,N_1573,N_138);
or U3348 (N_3348,N_1458,N_1605);
nor U3349 (N_3349,N_1801,N_1338);
nor U3350 (N_3350,N_1056,N_582);
nand U3351 (N_3351,N_31,N_788);
xor U3352 (N_3352,N_1574,N_930);
nor U3353 (N_3353,N_1395,N_1824);
or U3354 (N_3354,N_1035,N_14);
nand U3355 (N_3355,N_10,N_652);
nand U3356 (N_3356,N_429,N_803);
and U3357 (N_3357,N_1429,N_210);
and U3358 (N_3358,N_1028,N_375);
nand U3359 (N_3359,N_1654,N_1042);
or U3360 (N_3360,N_280,N_691);
xnor U3361 (N_3361,N_151,N_1847);
nor U3362 (N_3362,N_825,N_1888);
nand U3363 (N_3363,N_1375,N_631);
xor U3364 (N_3364,N_416,N_1724);
nor U3365 (N_3365,N_675,N_699);
and U3366 (N_3366,N_0,N_1936);
or U3367 (N_3367,N_420,N_159);
nor U3368 (N_3368,N_1767,N_319);
nand U3369 (N_3369,N_1955,N_180);
nand U3370 (N_3370,N_179,N_466);
nor U3371 (N_3371,N_927,N_366);
or U3372 (N_3372,N_1037,N_661);
nand U3373 (N_3373,N_46,N_369);
or U3374 (N_3374,N_523,N_771);
xor U3375 (N_3375,N_1721,N_475);
nand U3376 (N_3376,N_171,N_640);
nor U3377 (N_3377,N_1573,N_512);
and U3378 (N_3378,N_1801,N_159);
nor U3379 (N_3379,N_1430,N_1096);
or U3380 (N_3380,N_755,N_1230);
nor U3381 (N_3381,N_1786,N_1376);
and U3382 (N_3382,N_200,N_1312);
nand U3383 (N_3383,N_802,N_1133);
and U3384 (N_3384,N_1570,N_1920);
nor U3385 (N_3385,N_155,N_412);
nand U3386 (N_3386,N_1675,N_1589);
or U3387 (N_3387,N_1073,N_379);
and U3388 (N_3388,N_852,N_1109);
xnor U3389 (N_3389,N_1944,N_1097);
nand U3390 (N_3390,N_342,N_1118);
nor U3391 (N_3391,N_1431,N_816);
nor U3392 (N_3392,N_735,N_597);
xor U3393 (N_3393,N_1424,N_148);
xnor U3394 (N_3394,N_1956,N_535);
nand U3395 (N_3395,N_67,N_545);
and U3396 (N_3396,N_1162,N_406);
xnor U3397 (N_3397,N_1792,N_945);
nand U3398 (N_3398,N_867,N_676);
nand U3399 (N_3399,N_1650,N_452);
nand U3400 (N_3400,N_726,N_1214);
or U3401 (N_3401,N_968,N_1269);
and U3402 (N_3402,N_1594,N_1252);
nand U3403 (N_3403,N_1276,N_852);
or U3404 (N_3404,N_795,N_1172);
xor U3405 (N_3405,N_425,N_1148);
nand U3406 (N_3406,N_1732,N_671);
nand U3407 (N_3407,N_1545,N_1942);
nor U3408 (N_3408,N_1412,N_47);
and U3409 (N_3409,N_1353,N_395);
and U3410 (N_3410,N_529,N_1918);
nor U3411 (N_3411,N_1488,N_965);
nor U3412 (N_3412,N_1741,N_751);
nor U3413 (N_3413,N_1482,N_1625);
nor U3414 (N_3414,N_461,N_112);
or U3415 (N_3415,N_785,N_31);
or U3416 (N_3416,N_683,N_1824);
nor U3417 (N_3417,N_1857,N_546);
or U3418 (N_3418,N_1934,N_881);
or U3419 (N_3419,N_484,N_964);
nor U3420 (N_3420,N_318,N_1135);
nor U3421 (N_3421,N_1200,N_1682);
xor U3422 (N_3422,N_1882,N_206);
nor U3423 (N_3423,N_1897,N_1331);
nor U3424 (N_3424,N_429,N_762);
or U3425 (N_3425,N_1456,N_674);
and U3426 (N_3426,N_518,N_1885);
or U3427 (N_3427,N_178,N_1700);
nand U3428 (N_3428,N_1909,N_331);
xnor U3429 (N_3429,N_268,N_593);
nor U3430 (N_3430,N_312,N_1265);
nand U3431 (N_3431,N_815,N_979);
xor U3432 (N_3432,N_151,N_1465);
or U3433 (N_3433,N_1532,N_1869);
nor U3434 (N_3434,N_737,N_1687);
nor U3435 (N_3435,N_736,N_523);
or U3436 (N_3436,N_1260,N_286);
xnor U3437 (N_3437,N_410,N_1910);
nand U3438 (N_3438,N_1142,N_1954);
and U3439 (N_3439,N_421,N_365);
or U3440 (N_3440,N_1260,N_1025);
nand U3441 (N_3441,N_410,N_1520);
and U3442 (N_3442,N_673,N_1714);
or U3443 (N_3443,N_1122,N_1820);
and U3444 (N_3444,N_924,N_1535);
and U3445 (N_3445,N_869,N_572);
nand U3446 (N_3446,N_1021,N_1487);
xnor U3447 (N_3447,N_1999,N_228);
nand U3448 (N_3448,N_235,N_1401);
or U3449 (N_3449,N_1796,N_529);
xnor U3450 (N_3450,N_1091,N_1968);
or U3451 (N_3451,N_58,N_1745);
and U3452 (N_3452,N_1416,N_1731);
and U3453 (N_3453,N_54,N_1804);
nor U3454 (N_3454,N_1793,N_1018);
nor U3455 (N_3455,N_126,N_1432);
and U3456 (N_3456,N_694,N_658);
or U3457 (N_3457,N_1408,N_984);
nand U3458 (N_3458,N_1674,N_1025);
or U3459 (N_3459,N_580,N_990);
or U3460 (N_3460,N_607,N_1238);
nand U3461 (N_3461,N_1121,N_181);
xnor U3462 (N_3462,N_902,N_685);
nand U3463 (N_3463,N_784,N_746);
and U3464 (N_3464,N_512,N_7);
xor U3465 (N_3465,N_1949,N_1619);
nor U3466 (N_3466,N_1002,N_342);
nand U3467 (N_3467,N_1566,N_1582);
nand U3468 (N_3468,N_1675,N_1479);
nand U3469 (N_3469,N_1093,N_1961);
nand U3470 (N_3470,N_1058,N_1772);
and U3471 (N_3471,N_18,N_447);
and U3472 (N_3472,N_1313,N_373);
nor U3473 (N_3473,N_181,N_1710);
and U3474 (N_3474,N_851,N_684);
nor U3475 (N_3475,N_1553,N_1092);
nand U3476 (N_3476,N_958,N_402);
nand U3477 (N_3477,N_132,N_26);
nor U3478 (N_3478,N_1881,N_859);
nand U3479 (N_3479,N_1229,N_131);
nand U3480 (N_3480,N_1593,N_865);
nand U3481 (N_3481,N_722,N_0);
or U3482 (N_3482,N_469,N_1401);
xor U3483 (N_3483,N_1893,N_1871);
and U3484 (N_3484,N_1435,N_1540);
or U3485 (N_3485,N_1084,N_1857);
nand U3486 (N_3486,N_893,N_1088);
xnor U3487 (N_3487,N_1031,N_1163);
nand U3488 (N_3488,N_691,N_457);
and U3489 (N_3489,N_1103,N_1920);
or U3490 (N_3490,N_1350,N_897);
nor U3491 (N_3491,N_1163,N_1817);
or U3492 (N_3492,N_996,N_1452);
nand U3493 (N_3493,N_608,N_1772);
xnor U3494 (N_3494,N_963,N_1131);
or U3495 (N_3495,N_211,N_1082);
and U3496 (N_3496,N_261,N_1945);
nor U3497 (N_3497,N_1775,N_19);
nand U3498 (N_3498,N_249,N_153);
xor U3499 (N_3499,N_1412,N_1269);
nor U3500 (N_3500,N_1235,N_588);
and U3501 (N_3501,N_1677,N_376);
nand U3502 (N_3502,N_1147,N_1631);
and U3503 (N_3503,N_1374,N_1701);
and U3504 (N_3504,N_1793,N_280);
nor U3505 (N_3505,N_1446,N_1607);
or U3506 (N_3506,N_138,N_106);
nor U3507 (N_3507,N_1940,N_1133);
or U3508 (N_3508,N_1385,N_1020);
or U3509 (N_3509,N_1495,N_1040);
nor U3510 (N_3510,N_740,N_1865);
nor U3511 (N_3511,N_1417,N_301);
xnor U3512 (N_3512,N_868,N_1389);
nand U3513 (N_3513,N_1247,N_1510);
xnor U3514 (N_3514,N_583,N_1511);
nor U3515 (N_3515,N_1400,N_810);
nor U3516 (N_3516,N_378,N_1928);
and U3517 (N_3517,N_1607,N_1547);
nand U3518 (N_3518,N_107,N_1208);
or U3519 (N_3519,N_1833,N_22);
or U3520 (N_3520,N_1841,N_153);
and U3521 (N_3521,N_1288,N_1514);
nor U3522 (N_3522,N_374,N_1896);
nand U3523 (N_3523,N_1221,N_231);
or U3524 (N_3524,N_1404,N_1847);
and U3525 (N_3525,N_1332,N_608);
nor U3526 (N_3526,N_1882,N_1658);
nor U3527 (N_3527,N_861,N_1746);
and U3528 (N_3528,N_236,N_1572);
and U3529 (N_3529,N_1970,N_328);
nor U3530 (N_3530,N_1196,N_11);
and U3531 (N_3531,N_1664,N_1846);
and U3532 (N_3532,N_1290,N_472);
nor U3533 (N_3533,N_882,N_1338);
nor U3534 (N_3534,N_850,N_1426);
nor U3535 (N_3535,N_1715,N_1909);
nand U3536 (N_3536,N_1386,N_1815);
xnor U3537 (N_3537,N_814,N_134);
nor U3538 (N_3538,N_906,N_482);
xor U3539 (N_3539,N_1479,N_1689);
nor U3540 (N_3540,N_178,N_1429);
or U3541 (N_3541,N_111,N_1835);
xnor U3542 (N_3542,N_579,N_1912);
xnor U3543 (N_3543,N_1434,N_1574);
nand U3544 (N_3544,N_143,N_580);
xor U3545 (N_3545,N_846,N_1996);
and U3546 (N_3546,N_815,N_1700);
and U3547 (N_3547,N_75,N_523);
nor U3548 (N_3548,N_1765,N_1185);
or U3549 (N_3549,N_1004,N_1505);
nand U3550 (N_3550,N_1531,N_738);
or U3551 (N_3551,N_398,N_1758);
and U3552 (N_3552,N_14,N_522);
xor U3553 (N_3553,N_711,N_75);
and U3554 (N_3554,N_946,N_1731);
nand U3555 (N_3555,N_1501,N_588);
xnor U3556 (N_3556,N_1174,N_672);
nand U3557 (N_3557,N_1758,N_39);
and U3558 (N_3558,N_373,N_1098);
xor U3559 (N_3559,N_477,N_945);
and U3560 (N_3560,N_987,N_159);
nand U3561 (N_3561,N_1292,N_1863);
and U3562 (N_3562,N_610,N_701);
nand U3563 (N_3563,N_57,N_686);
nand U3564 (N_3564,N_1178,N_470);
or U3565 (N_3565,N_227,N_611);
xor U3566 (N_3566,N_1685,N_1922);
nand U3567 (N_3567,N_423,N_28);
nand U3568 (N_3568,N_391,N_776);
or U3569 (N_3569,N_833,N_385);
nand U3570 (N_3570,N_1169,N_435);
nand U3571 (N_3571,N_1555,N_1401);
nor U3572 (N_3572,N_1548,N_1764);
nor U3573 (N_3573,N_1,N_1969);
nand U3574 (N_3574,N_816,N_1404);
or U3575 (N_3575,N_1769,N_1010);
xnor U3576 (N_3576,N_184,N_1552);
and U3577 (N_3577,N_1519,N_706);
nand U3578 (N_3578,N_1956,N_989);
nand U3579 (N_3579,N_1034,N_1888);
nor U3580 (N_3580,N_1730,N_1393);
nor U3581 (N_3581,N_1249,N_285);
or U3582 (N_3582,N_180,N_1244);
nand U3583 (N_3583,N_927,N_22);
nand U3584 (N_3584,N_1106,N_1034);
or U3585 (N_3585,N_74,N_1822);
or U3586 (N_3586,N_1079,N_508);
nand U3587 (N_3587,N_1475,N_753);
nand U3588 (N_3588,N_1835,N_1134);
and U3589 (N_3589,N_21,N_1505);
nor U3590 (N_3590,N_1076,N_290);
nor U3591 (N_3591,N_962,N_1419);
nor U3592 (N_3592,N_1893,N_1526);
or U3593 (N_3593,N_1072,N_446);
nand U3594 (N_3594,N_1524,N_1791);
nor U3595 (N_3595,N_1660,N_1595);
nor U3596 (N_3596,N_534,N_9);
nor U3597 (N_3597,N_1487,N_1684);
or U3598 (N_3598,N_849,N_1000);
and U3599 (N_3599,N_425,N_1781);
nor U3600 (N_3600,N_285,N_363);
and U3601 (N_3601,N_1722,N_1264);
or U3602 (N_3602,N_260,N_885);
or U3603 (N_3603,N_1339,N_1854);
or U3604 (N_3604,N_1612,N_48);
nor U3605 (N_3605,N_106,N_1216);
nor U3606 (N_3606,N_1904,N_851);
nor U3607 (N_3607,N_1225,N_308);
and U3608 (N_3608,N_1397,N_1999);
and U3609 (N_3609,N_1962,N_962);
or U3610 (N_3610,N_1829,N_638);
or U3611 (N_3611,N_1505,N_1412);
nand U3612 (N_3612,N_609,N_1567);
nor U3613 (N_3613,N_876,N_163);
or U3614 (N_3614,N_569,N_905);
xor U3615 (N_3615,N_979,N_405);
or U3616 (N_3616,N_435,N_1269);
nor U3617 (N_3617,N_104,N_1091);
nand U3618 (N_3618,N_1908,N_175);
and U3619 (N_3619,N_943,N_1677);
and U3620 (N_3620,N_1757,N_1256);
and U3621 (N_3621,N_1075,N_780);
nor U3622 (N_3622,N_659,N_1441);
nor U3623 (N_3623,N_785,N_1457);
or U3624 (N_3624,N_499,N_1726);
and U3625 (N_3625,N_1373,N_1574);
xnor U3626 (N_3626,N_1007,N_1532);
nor U3627 (N_3627,N_1570,N_552);
xor U3628 (N_3628,N_634,N_287);
and U3629 (N_3629,N_919,N_1368);
and U3630 (N_3630,N_862,N_581);
nand U3631 (N_3631,N_1385,N_601);
and U3632 (N_3632,N_1146,N_1574);
and U3633 (N_3633,N_1056,N_1164);
xor U3634 (N_3634,N_1425,N_1641);
and U3635 (N_3635,N_648,N_1891);
or U3636 (N_3636,N_42,N_754);
nand U3637 (N_3637,N_1122,N_116);
and U3638 (N_3638,N_1831,N_1796);
and U3639 (N_3639,N_1376,N_1866);
and U3640 (N_3640,N_1986,N_1903);
nand U3641 (N_3641,N_1270,N_845);
nor U3642 (N_3642,N_28,N_1415);
or U3643 (N_3643,N_1233,N_319);
and U3644 (N_3644,N_581,N_1898);
nor U3645 (N_3645,N_1928,N_1105);
xor U3646 (N_3646,N_369,N_1846);
or U3647 (N_3647,N_646,N_85);
or U3648 (N_3648,N_1093,N_1543);
xor U3649 (N_3649,N_1855,N_57);
or U3650 (N_3650,N_1610,N_474);
nor U3651 (N_3651,N_494,N_1764);
nor U3652 (N_3652,N_1956,N_351);
or U3653 (N_3653,N_1925,N_1358);
and U3654 (N_3654,N_966,N_1102);
and U3655 (N_3655,N_722,N_1628);
nand U3656 (N_3656,N_378,N_264);
or U3657 (N_3657,N_1457,N_293);
xnor U3658 (N_3658,N_1714,N_598);
or U3659 (N_3659,N_919,N_1453);
nor U3660 (N_3660,N_1066,N_1850);
or U3661 (N_3661,N_1837,N_953);
nor U3662 (N_3662,N_268,N_1186);
nor U3663 (N_3663,N_1935,N_1553);
nor U3664 (N_3664,N_1830,N_302);
nor U3665 (N_3665,N_476,N_579);
or U3666 (N_3666,N_1278,N_190);
nor U3667 (N_3667,N_342,N_1312);
and U3668 (N_3668,N_1825,N_370);
nor U3669 (N_3669,N_925,N_1143);
nand U3670 (N_3670,N_1891,N_1126);
nor U3671 (N_3671,N_293,N_546);
nor U3672 (N_3672,N_692,N_1856);
nor U3673 (N_3673,N_1667,N_1746);
and U3674 (N_3674,N_538,N_1620);
or U3675 (N_3675,N_1072,N_1046);
and U3676 (N_3676,N_1306,N_1348);
and U3677 (N_3677,N_1752,N_1181);
nor U3678 (N_3678,N_1438,N_618);
nor U3679 (N_3679,N_1949,N_1104);
or U3680 (N_3680,N_1792,N_1538);
nand U3681 (N_3681,N_1009,N_1315);
nand U3682 (N_3682,N_457,N_1816);
nor U3683 (N_3683,N_1287,N_1078);
and U3684 (N_3684,N_1726,N_1525);
nor U3685 (N_3685,N_1449,N_1057);
and U3686 (N_3686,N_1870,N_249);
nand U3687 (N_3687,N_1894,N_1031);
nand U3688 (N_3688,N_475,N_310);
nand U3689 (N_3689,N_1699,N_1230);
and U3690 (N_3690,N_1967,N_639);
xnor U3691 (N_3691,N_336,N_467);
nand U3692 (N_3692,N_1327,N_1309);
nand U3693 (N_3693,N_1069,N_407);
or U3694 (N_3694,N_381,N_1598);
and U3695 (N_3695,N_1019,N_1242);
and U3696 (N_3696,N_960,N_133);
or U3697 (N_3697,N_821,N_399);
nand U3698 (N_3698,N_1589,N_895);
nor U3699 (N_3699,N_1535,N_183);
or U3700 (N_3700,N_682,N_1733);
and U3701 (N_3701,N_1453,N_640);
and U3702 (N_3702,N_1465,N_506);
and U3703 (N_3703,N_1381,N_615);
and U3704 (N_3704,N_967,N_133);
or U3705 (N_3705,N_1267,N_1797);
nand U3706 (N_3706,N_1269,N_1769);
and U3707 (N_3707,N_160,N_459);
nand U3708 (N_3708,N_951,N_240);
nor U3709 (N_3709,N_1257,N_1983);
nor U3710 (N_3710,N_1601,N_1149);
nor U3711 (N_3711,N_450,N_781);
xnor U3712 (N_3712,N_299,N_328);
nor U3713 (N_3713,N_589,N_919);
nand U3714 (N_3714,N_762,N_111);
nor U3715 (N_3715,N_664,N_1908);
and U3716 (N_3716,N_1855,N_1313);
nand U3717 (N_3717,N_352,N_1616);
or U3718 (N_3718,N_545,N_148);
xor U3719 (N_3719,N_709,N_796);
and U3720 (N_3720,N_360,N_951);
or U3721 (N_3721,N_247,N_995);
or U3722 (N_3722,N_327,N_439);
or U3723 (N_3723,N_545,N_1729);
or U3724 (N_3724,N_1325,N_1987);
and U3725 (N_3725,N_1540,N_1419);
nor U3726 (N_3726,N_396,N_1657);
nor U3727 (N_3727,N_1565,N_1592);
and U3728 (N_3728,N_1408,N_823);
nand U3729 (N_3729,N_190,N_1382);
or U3730 (N_3730,N_465,N_624);
nand U3731 (N_3731,N_1608,N_263);
xnor U3732 (N_3732,N_1974,N_1652);
or U3733 (N_3733,N_226,N_1671);
and U3734 (N_3734,N_61,N_1032);
nand U3735 (N_3735,N_1820,N_1477);
or U3736 (N_3736,N_1083,N_1830);
and U3737 (N_3737,N_101,N_707);
or U3738 (N_3738,N_1345,N_1002);
and U3739 (N_3739,N_1732,N_1011);
xnor U3740 (N_3740,N_232,N_1503);
and U3741 (N_3741,N_1236,N_823);
or U3742 (N_3742,N_962,N_1558);
and U3743 (N_3743,N_302,N_1371);
and U3744 (N_3744,N_1079,N_1798);
or U3745 (N_3745,N_156,N_747);
xnor U3746 (N_3746,N_873,N_1460);
or U3747 (N_3747,N_25,N_578);
nand U3748 (N_3748,N_1092,N_806);
nor U3749 (N_3749,N_631,N_1551);
nand U3750 (N_3750,N_1091,N_1829);
or U3751 (N_3751,N_370,N_244);
nand U3752 (N_3752,N_551,N_1013);
and U3753 (N_3753,N_1355,N_1178);
nor U3754 (N_3754,N_353,N_133);
nand U3755 (N_3755,N_1827,N_1251);
and U3756 (N_3756,N_1796,N_1541);
and U3757 (N_3757,N_1699,N_274);
nor U3758 (N_3758,N_393,N_836);
or U3759 (N_3759,N_1283,N_718);
nand U3760 (N_3760,N_1143,N_587);
or U3761 (N_3761,N_1523,N_83);
nor U3762 (N_3762,N_1294,N_1860);
xnor U3763 (N_3763,N_1618,N_1221);
and U3764 (N_3764,N_751,N_1161);
nor U3765 (N_3765,N_404,N_918);
nand U3766 (N_3766,N_20,N_1512);
nand U3767 (N_3767,N_1884,N_639);
xnor U3768 (N_3768,N_1498,N_1746);
nand U3769 (N_3769,N_1740,N_1725);
nand U3770 (N_3770,N_1950,N_1160);
xnor U3771 (N_3771,N_1757,N_1129);
nand U3772 (N_3772,N_919,N_763);
and U3773 (N_3773,N_457,N_1261);
or U3774 (N_3774,N_1614,N_451);
and U3775 (N_3775,N_1479,N_60);
and U3776 (N_3776,N_1781,N_1376);
or U3777 (N_3777,N_1109,N_1611);
nand U3778 (N_3778,N_794,N_674);
xor U3779 (N_3779,N_887,N_988);
xor U3780 (N_3780,N_898,N_1339);
nand U3781 (N_3781,N_45,N_1464);
and U3782 (N_3782,N_1969,N_725);
nor U3783 (N_3783,N_1285,N_751);
nand U3784 (N_3784,N_1363,N_321);
nand U3785 (N_3785,N_137,N_320);
and U3786 (N_3786,N_588,N_1880);
or U3787 (N_3787,N_937,N_1234);
or U3788 (N_3788,N_127,N_532);
xnor U3789 (N_3789,N_710,N_322);
and U3790 (N_3790,N_1567,N_229);
and U3791 (N_3791,N_21,N_1917);
xnor U3792 (N_3792,N_379,N_595);
xor U3793 (N_3793,N_1696,N_1538);
nand U3794 (N_3794,N_1531,N_456);
nand U3795 (N_3795,N_564,N_668);
and U3796 (N_3796,N_1048,N_922);
and U3797 (N_3797,N_1374,N_1002);
and U3798 (N_3798,N_410,N_922);
nor U3799 (N_3799,N_1231,N_821);
nor U3800 (N_3800,N_958,N_160);
nor U3801 (N_3801,N_1882,N_1140);
nand U3802 (N_3802,N_756,N_1232);
nor U3803 (N_3803,N_1308,N_1057);
nand U3804 (N_3804,N_1858,N_881);
or U3805 (N_3805,N_1752,N_1264);
and U3806 (N_3806,N_1743,N_1471);
nand U3807 (N_3807,N_1605,N_80);
and U3808 (N_3808,N_1381,N_1536);
and U3809 (N_3809,N_909,N_632);
nand U3810 (N_3810,N_768,N_662);
or U3811 (N_3811,N_301,N_1864);
or U3812 (N_3812,N_324,N_1424);
xor U3813 (N_3813,N_1697,N_1951);
nand U3814 (N_3814,N_1710,N_401);
nor U3815 (N_3815,N_382,N_916);
and U3816 (N_3816,N_1227,N_924);
nor U3817 (N_3817,N_1520,N_417);
and U3818 (N_3818,N_1591,N_874);
or U3819 (N_3819,N_823,N_898);
and U3820 (N_3820,N_171,N_949);
and U3821 (N_3821,N_883,N_157);
or U3822 (N_3822,N_871,N_1274);
nor U3823 (N_3823,N_1689,N_866);
and U3824 (N_3824,N_1849,N_1035);
or U3825 (N_3825,N_1570,N_887);
nand U3826 (N_3826,N_520,N_897);
nand U3827 (N_3827,N_883,N_224);
nand U3828 (N_3828,N_1177,N_1452);
nand U3829 (N_3829,N_1380,N_1672);
nand U3830 (N_3830,N_729,N_660);
and U3831 (N_3831,N_38,N_434);
nor U3832 (N_3832,N_434,N_477);
or U3833 (N_3833,N_857,N_408);
xnor U3834 (N_3834,N_611,N_930);
and U3835 (N_3835,N_1636,N_1048);
and U3836 (N_3836,N_1633,N_1365);
nand U3837 (N_3837,N_1493,N_1330);
or U3838 (N_3838,N_275,N_825);
nand U3839 (N_3839,N_711,N_340);
and U3840 (N_3840,N_390,N_1231);
nor U3841 (N_3841,N_1659,N_1077);
nor U3842 (N_3842,N_916,N_308);
nor U3843 (N_3843,N_807,N_202);
or U3844 (N_3844,N_684,N_201);
nand U3845 (N_3845,N_862,N_917);
nand U3846 (N_3846,N_1275,N_1057);
xnor U3847 (N_3847,N_621,N_833);
nor U3848 (N_3848,N_796,N_68);
nand U3849 (N_3849,N_1110,N_138);
or U3850 (N_3850,N_1279,N_879);
nand U3851 (N_3851,N_1915,N_795);
or U3852 (N_3852,N_908,N_1151);
nand U3853 (N_3853,N_137,N_409);
or U3854 (N_3854,N_283,N_1142);
nand U3855 (N_3855,N_1978,N_981);
nand U3856 (N_3856,N_1960,N_579);
and U3857 (N_3857,N_1390,N_1834);
nand U3858 (N_3858,N_1980,N_1865);
and U3859 (N_3859,N_529,N_1583);
nor U3860 (N_3860,N_1610,N_369);
and U3861 (N_3861,N_980,N_57);
or U3862 (N_3862,N_1461,N_1452);
nor U3863 (N_3863,N_1087,N_436);
nand U3864 (N_3864,N_437,N_629);
or U3865 (N_3865,N_504,N_593);
and U3866 (N_3866,N_1593,N_1164);
or U3867 (N_3867,N_1358,N_1104);
nor U3868 (N_3868,N_1441,N_1107);
nand U3869 (N_3869,N_1113,N_1490);
and U3870 (N_3870,N_233,N_1845);
nand U3871 (N_3871,N_168,N_301);
nand U3872 (N_3872,N_510,N_767);
nand U3873 (N_3873,N_1680,N_1414);
or U3874 (N_3874,N_1900,N_1719);
nor U3875 (N_3875,N_380,N_1739);
or U3876 (N_3876,N_24,N_1553);
and U3877 (N_3877,N_984,N_1755);
nor U3878 (N_3878,N_829,N_1555);
nor U3879 (N_3879,N_268,N_489);
or U3880 (N_3880,N_1558,N_1659);
nand U3881 (N_3881,N_848,N_1156);
nor U3882 (N_3882,N_1921,N_133);
xnor U3883 (N_3883,N_899,N_1518);
xnor U3884 (N_3884,N_150,N_1499);
nand U3885 (N_3885,N_393,N_775);
nand U3886 (N_3886,N_1121,N_1514);
nand U3887 (N_3887,N_559,N_1597);
nor U3888 (N_3888,N_1958,N_1797);
nand U3889 (N_3889,N_761,N_1957);
nor U3890 (N_3890,N_394,N_1592);
xnor U3891 (N_3891,N_121,N_842);
nor U3892 (N_3892,N_390,N_1048);
xnor U3893 (N_3893,N_398,N_1304);
or U3894 (N_3894,N_1529,N_1908);
or U3895 (N_3895,N_1683,N_1876);
nor U3896 (N_3896,N_1717,N_922);
or U3897 (N_3897,N_850,N_80);
and U3898 (N_3898,N_987,N_670);
nand U3899 (N_3899,N_541,N_1926);
or U3900 (N_3900,N_1971,N_1601);
nand U3901 (N_3901,N_1018,N_29);
nand U3902 (N_3902,N_1769,N_561);
or U3903 (N_3903,N_1013,N_1908);
nor U3904 (N_3904,N_1183,N_290);
nand U3905 (N_3905,N_958,N_1413);
or U3906 (N_3906,N_484,N_1102);
nand U3907 (N_3907,N_1862,N_902);
and U3908 (N_3908,N_1813,N_1027);
nand U3909 (N_3909,N_1159,N_199);
or U3910 (N_3910,N_60,N_1595);
nor U3911 (N_3911,N_822,N_1676);
nand U3912 (N_3912,N_1265,N_556);
nand U3913 (N_3913,N_72,N_1297);
or U3914 (N_3914,N_814,N_169);
xnor U3915 (N_3915,N_1456,N_1852);
or U3916 (N_3916,N_141,N_1575);
or U3917 (N_3917,N_1385,N_619);
xnor U3918 (N_3918,N_1055,N_1383);
nor U3919 (N_3919,N_297,N_1165);
and U3920 (N_3920,N_1785,N_1074);
and U3921 (N_3921,N_1404,N_499);
or U3922 (N_3922,N_167,N_830);
xnor U3923 (N_3923,N_1525,N_1832);
xnor U3924 (N_3924,N_730,N_418);
and U3925 (N_3925,N_1423,N_189);
nand U3926 (N_3926,N_714,N_567);
and U3927 (N_3927,N_666,N_908);
nand U3928 (N_3928,N_800,N_1888);
xnor U3929 (N_3929,N_1134,N_1423);
xor U3930 (N_3930,N_1543,N_615);
or U3931 (N_3931,N_1629,N_420);
nor U3932 (N_3932,N_793,N_205);
or U3933 (N_3933,N_880,N_953);
nor U3934 (N_3934,N_1181,N_520);
xnor U3935 (N_3935,N_840,N_1721);
nand U3936 (N_3936,N_1645,N_1100);
and U3937 (N_3937,N_1405,N_924);
nor U3938 (N_3938,N_1448,N_837);
and U3939 (N_3939,N_93,N_857);
nand U3940 (N_3940,N_95,N_674);
nand U3941 (N_3941,N_1183,N_543);
or U3942 (N_3942,N_1627,N_987);
nand U3943 (N_3943,N_284,N_163);
xnor U3944 (N_3944,N_1737,N_1870);
or U3945 (N_3945,N_1800,N_783);
and U3946 (N_3946,N_1675,N_1232);
or U3947 (N_3947,N_991,N_660);
nor U3948 (N_3948,N_855,N_1162);
nand U3949 (N_3949,N_1313,N_1217);
or U3950 (N_3950,N_503,N_11);
xnor U3951 (N_3951,N_47,N_1052);
nand U3952 (N_3952,N_695,N_1309);
nor U3953 (N_3953,N_1847,N_1352);
xor U3954 (N_3954,N_60,N_1618);
nand U3955 (N_3955,N_1477,N_389);
or U3956 (N_3956,N_978,N_864);
xnor U3957 (N_3957,N_1019,N_1521);
or U3958 (N_3958,N_773,N_324);
nand U3959 (N_3959,N_755,N_332);
nor U3960 (N_3960,N_1161,N_1899);
nand U3961 (N_3961,N_648,N_105);
or U3962 (N_3962,N_1693,N_730);
and U3963 (N_3963,N_468,N_1961);
and U3964 (N_3964,N_121,N_1109);
nor U3965 (N_3965,N_1410,N_1457);
nand U3966 (N_3966,N_1862,N_779);
and U3967 (N_3967,N_576,N_1485);
and U3968 (N_3968,N_374,N_1481);
nor U3969 (N_3969,N_1229,N_579);
and U3970 (N_3970,N_506,N_1603);
and U3971 (N_3971,N_1812,N_1234);
nor U3972 (N_3972,N_971,N_730);
nand U3973 (N_3973,N_1236,N_1755);
nand U3974 (N_3974,N_728,N_1276);
or U3975 (N_3975,N_987,N_369);
and U3976 (N_3976,N_5,N_137);
xor U3977 (N_3977,N_1003,N_890);
or U3978 (N_3978,N_20,N_19);
and U3979 (N_3979,N_1895,N_1254);
and U3980 (N_3980,N_1870,N_27);
xor U3981 (N_3981,N_902,N_1566);
nand U3982 (N_3982,N_1204,N_972);
nor U3983 (N_3983,N_160,N_1583);
or U3984 (N_3984,N_1744,N_1765);
xor U3985 (N_3985,N_664,N_1303);
and U3986 (N_3986,N_1804,N_654);
nor U3987 (N_3987,N_1484,N_277);
nand U3988 (N_3988,N_1907,N_295);
nor U3989 (N_3989,N_1311,N_249);
or U3990 (N_3990,N_461,N_1016);
or U3991 (N_3991,N_284,N_1017);
nor U3992 (N_3992,N_1225,N_1247);
and U3993 (N_3993,N_478,N_1850);
or U3994 (N_3994,N_164,N_576);
nand U3995 (N_3995,N_62,N_1884);
nor U3996 (N_3996,N_160,N_791);
or U3997 (N_3997,N_1962,N_1776);
nor U3998 (N_3998,N_1676,N_1578);
nand U3999 (N_3999,N_1852,N_427);
nand U4000 (N_4000,N_3265,N_3390);
xor U4001 (N_4001,N_3917,N_2330);
and U4002 (N_4002,N_3904,N_3964);
or U4003 (N_4003,N_2667,N_2722);
nor U4004 (N_4004,N_2303,N_3594);
and U4005 (N_4005,N_2275,N_2370);
nand U4006 (N_4006,N_3667,N_3123);
and U4007 (N_4007,N_3277,N_2659);
and U4008 (N_4008,N_2091,N_3120);
or U4009 (N_4009,N_3126,N_2719);
xor U4010 (N_4010,N_3600,N_2577);
nor U4011 (N_4011,N_3525,N_2891);
and U4012 (N_4012,N_2819,N_2098);
or U4013 (N_4013,N_2400,N_3151);
and U4014 (N_4014,N_2916,N_2249);
xor U4015 (N_4015,N_2403,N_2900);
nor U4016 (N_4016,N_3872,N_3546);
nand U4017 (N_4017,N_3376,N_3293);
nor U4018 (N_4018,N_2467,N_2849);
and U4019 (N_4019,N_2110,N_3219);
and U4020 (N_4020,N_2525,N_2935);
nand U4021 (N_4021,N_2449,N_2382);
xnor U4022 (N_4022,N_2247,N_3560);
nand U4023 (N_4023,N_3564,N_2172);
and U4024 (N_4024,N_3436,N_3065);
and U4025 (N_4025,N_3645,N_3588);
nor U4026 (N_4026,N_2643,N_3441);
and U4027 (N_4027,N_2123,N_2688);
and U4028 (N_4028,N_3721,N_2493);
and U4029 (N_4029,N_3761,N_3678);
nor U4030 (N_4030,N_3996,N_3179);
and U4031 (N_4031,N_3599,N_2919);
nor U4032 (N_4032,N_3103,N_3924);
nor U4033 (N_4033,N_2011,N_3337);
or U4034 (N_4034,N_2317,N_2202);
or U4035 (N_4035,N_3576,N_3346);
or U4036 (N_4036,N_3838,N_3325);
or U4037 (N_4037,N_3938,N_2628);
nor U4038 (N_4038,N_3510,N_2352);
nor U4039 (N_4039,N_2936,N_2072);
and U4040 (N_4040,N_3225,N_2047);
nor U4041 (N_4041,N_3314,N_3134);
nor U4042 (N_4042,N_2333,N_2086);
nand U4043 (N_4043,N_2534,N_2353);
or U4044 (N_4044,N_2677,N_3983);
or U4045 (N_4045,N_2351,N_2608);
nor U4046 (N_4046,N_3654,N_3979);
or U4047 (N_4047,N_2093,N_3211);
nor U4048 (N_4048,N_3319,N_2166);
nand U4049 (N_4049,N_2368,N_2298);
nor U4050 (N_4050,N_3919,N_3534);
and U4051 (N_4051,N_2447,N_3117);
nand U4052 (N_4052,N_3821,N_3460);
and U4053 (N_4053,N_3128,N_2282);
nand U4054 (N_4054,N_2068,N_3063);
nand U4055 (N_4055,N_3552,N_3495);
xor U4056 (N_4056,N_2700,N_3630);
or U4057 (N_4057,N_2035,N_3439);
nand U4058 (N_4058,N_2087,N_3596);
nand U4059 (N_4059,N_2452,N_2004);
and U4060 (N_4060,N_2552,N_3612);
and U4061 (N_4061,N_3090,N_3703);
and U4062 (N_4062,N_3429,N_3110);
and U4063 (N_4063,N_3885,N_3694);
nand U4064 (N_4064,N_3250,N_3816);
or U4065 (N_4065,N_2531,N_3178);
and U4066 (N_4066,N_3953,N_2567);
nand U4067 (N_4067,N_2080,N_2085);
nor U4068 (N_4068,N_3352,N_2626);
and U4069 (N_4069,N_3805,N_3054);
xnor U4070 (N_4070,N_3375,N_2242);
and U4071 (N_4071,N_2599,N_2825);
nand U4072 (N_4072,N_3545,N_2863);
and U4073 (N_4073,N_2171,N_3882);
and U4074 (N_4074,N_2573,N_2704);
nand U4075 (N_4075,N_3172,N_2446);
nor U4076 (N_4076,N_2651,N_3501);
nor U4077 (N_4077,N_2150,N_3527);
nor U4078 (N_4078,N_2977,N_3034);
nand U4079 (N_4079,N_2218,N_3454);
and U4080 (N_4080,N_3614,N_3832);
nor U4081 (N_4081,N_2813,N_2789);
and U4082 (N_4082,N_3758,N_3089);
nand U4083 (N_4083,N_3310,N_3666);
or U4084 (N_4084,N_3773,N_2990);
or U4085 (N_4085,N_2926,N_3253);
nor U4086 (N_4086,N_3543,N_2945);
xnor U4087 (N_4087,N_2685,N_3001);
nand U4088 (N_4088,N_2959,N_3131);
or U4089 (N_4089,N_3458,N_3580);
nor U4090 (N_4090,N_2886,N_3391);
nor U4091 (N_4091,N_3493,N_3108);
nor U4092 (N_4092,N_2019,N_3003);
xor U4093 (N_4093,N_3792,N_2769);
nor U4094 (N_4094,N_3035,N_3130);
and U4095 (N_4095,N_3323,N_2551);
or U4096 (N_4096,N_2804,N_3831);
nor U4097 (N_4097,N_2345,N_3149);
xor U4098 (N_4098,N_2025,N_3371);
or U4099 (N_4099,N_3412,N_3058);
and U4100 (N_4100,N_3107,N_3733);
nand U4101 (N_4101,N_2103,N_3189);
or U4102 (N_4102,N_2031,N_2294);
nor U4103 (N_4103,N_3651,N_2033);
and U4104 (N_4104,N_3389,N_2720);
nor U4105 (N_4105,N_2770,N_3574);
nor U4106 (N_4106,N_3186,N_3064);
or U4107 (N_4107,N_2005,N_3680);
and U4108 (N_4108,N_2416,N_2799);
nor U4109 (N_4109,N_2864,N_2523);
and U4110 (N_4110,N_3096,N_2854);
nand U4111 (N_4111,N_3074,N_3078);
nor U4112 (N_4112,N_2413,N_2794);
nor U4113 (N_4113,N_3213,N_2765);
nand U4114 (N_4114,N_2844,N_3039);
nor U4115 (N_4115,N_2852,N_2417);
nand U4116 (N_4116,N_3586,N_2342);
nor U4117 (N_4117,N_3359,N_2028);
or U4118 (N_4118,N_3749,N_2873);
nand U4119 (N_4119,N_2461,N_3767);
nor U4120 (N_4120,N_2848,N_3555);
nor U4121 (N_4121,N_2939,N_3809);
or U4122 (N_4122,N_2940,N_3762);
nor U4123 (N_4123,N_2271,N_2327);
nor U4124 (N_4124,N_2728,N_2645);
xor U4125 (N_4125,N_2159,N_3868);
nor U4126 (N_4126,N_2843,N_2419);
and U4127 (N_4127,N_2438,N_2829);
nor U4128 (N_4128,N_2509,N_3852);
and U4129 (N_4129,N_2000,N_3930);
nor U4130 (N_4130,N_2961,N_3264);
nand U4131 (N_4131,N_3661,N_3619);
and U4132 (N_4132,N_2678,N_3918);
and U4133 (N_4133,N_2928,N_2931);
or U4134 (N_4134,N_3989,N_2772);
and U4135 (N_4135,N_2308,N_3477);
nor U4136 (N_4136,N_2328,N_3158);
nor U4137 (N_4137,N_3633,N_2563);
nand U4138 (N_4138,N_3320,N_2823);
and U4139 (N_4139,N_2008,N_3598);
nand U4140 (N_4140,N_3780,N_2780);
and U4141 (N_4141,N_2623,N_2927);
nor U4142 (N_4142,N_3027,N_3981);
or U4143 (N_4143,N_2557,N_3741);
nand U4144 (N_4144,N_2660,N_2715);
and U4145 (N_4145,N_2965,N_2251);
or U4146 (N_4146,N_3424,N_2032);
xnor U4147 (N_4147,N_3940,N_2228);
or U4148 (N_4148,N_3331,N_2395);
or U4149 (N_4149,N_2290,N_3632);
xor U4150 (N_4150,N_3031,N_3044);
nand U4151 (N_4151,N_3242,N_3068);
and U4152 (N_4152,N_3797,N_2445);
nand U4153 (N_4153,N_3479,N_3071);
and U4154 (N_4154,N_2361,N_2778);
or U4155 (N_4155,N_3509,N_3687);
nor U4156 (N_4156,N_3112,N_2260);
xor U4157 (N_4157,N_3911,N_3283);
nand U4158 (N_4158,N_2473,N_2040);
xnor U4159 (N_4159,N_2605,N_2458);
nor U4160 (N_4160,N_3897,N_2853);
or U4161 (N_4161,N_2401,N_3245);
nand U4162 (N_4162,N_3905,N_2606);
xor U4163 (N_4163,N_2572,N_2138);
nand U4164 (N_4164,N_3629,N_2244);
and U4165 (N_4165,N_3269,N_3069);
nand U4166 (N_4166,N_3469,N_2077);
or U4167 (N_4167,N_3512,N_2276);
and U4168 (N_4168,N_3162,N_2556);
or U4169 (N_4169,N_2329,N_2131);
xor U4170 (N_4170,N_2256,N_2578);
and U4171 (N_4171,N_2991,N_2430);
nor U4172 (N_4172,N_3018,N_3430);
nor U4173 (N_4173,N_3975,N_3876);
xnor U4174 (N_4174,N_3674,N_3354);
nand U4175 (N_4175,N_2281,N_2670);
xor U4176 (N_4176,N_3308,N_2186);
and U4177 (N_4177,N_2518,N_3461);
nor U4178 (N_4178,N_3582,N_2754);
or U4179 (N_4179,N_2966,N_2462);
nor U4180 (N_4180,N_2513,N_2671);
and U4181 (N_4181,N_3384,N_2946);
nor U4182 (N_4182,N_2061,N_3340);
and U4183 (N_4183,N_3717,N_3038);
xor U4184 (N_4184,N_2869,N_2027);
and U4185 (N_4185,N_2768,N_3829);
and U4186 (N_4186,N_2358,N_2614);
nand U4187 (N_4187,N_3474,N_3305);
or U4188 (N_4188,N_2117,N_2998);
nor U4189 (N_4189,N_2151,N_2127);
nand U4190 (N_4190,N_3641,N_2341);
xnor U4191 (N_4191,N_3272,N_3777);
xnor U4192 (N_4192,N_2297,N_3148);
xnor U4193 (N_4193,N_3693,N_2526);
nand U4194 (N_4194,N_3326,N_2976);
or U4195 (N_4195,N_2725,N_3966);
xnor U4196 (N_4196,N_2665,N_2586);
xnor U4197 (N_4197,N_3855,N_3754);
nor U4198 (N_4198,N_3382,N_2129);
xor U4199 (N_4199,N_3794,N_3472);
and U4200 (N_4200,N_2496,N_2189);
or U4201 (N_4201,N_3046,N_3800);
nor U4202 (N_4202,N_2953,N_3714);
or U4203 (N_4203,N_3528,N_2646);
xnor U4204 (N_4204,N_2310,N_3113);
nor U4205 (N_4205,N_2639,N_3526);
and U4206 (N_4206,N_3462,N_2135);
and U4207 (N_4207,N_2376,N_2755);
xor U4208 (N_4208,N_3150,N_2680);
nand U4209 (N_4209,N_2870,N_2633);
nor U4210 (N_4210,N_2668,N_3570);
or U4211 (N_4211,N_2817,N_3812);
nand U4212 (N_4212,N_2740,N_2437);
or U4213 (N_4213,N_2954,N_2672);
nand U4214 (N_4214,N_2681,N_3788);
or U4215 (N_4215,N_3124,N_2459);
xor U4216 (N_4216,N_2958,N_3779);
nand U4217 (N_4217,N_3569,N_2283);
and U4218 (N_4218,N_2266,N_2206);
or U4219 (N_4219,N_3668,N_2180);
nor U4220 (N_4220,N_3273,N_3763);
nor U4221 (N_4221,N_2409,N_2357);
and U4222 (N_4222,N_3553,N_2197);
nor U4223 (N_4223,N_3377,N_3486);
nand U4224 (N_4224,N_3214,N_2280);
nand U4225 (N_4225,N_3874,N_2974);
nand U4226 (N_4226,N_2058,N_3239);
nand U4227 (N_4227,N_2391,N_3077);
nand U4228 (N_4228,N_2257,N_3009);
nor U4229 (N_4229,N_2487,N_3615);
nor U4230 (N_4230,N_2508,N_2495);
or U4231 (N_4231,N_3042,N_3862);
and U4232 (N_4232,N_2846,N_2845);
nor U4233 (N_4233,N_3037,N_2264);
nand U4234 (N_4234,N_2405,N_2827);
or U4235 (N_4235,N_2293,N_3175);
or U4236 (N_4236,N_3743,N_2250);
and U4237 (N_4237,N_2914,N_2761);
or U4238 (N_4238,N_3254,N_3476);
and U4239 (N_4239,N_2512,N_2017);
nor U4240 (N_4240,N_2270,N_2111);
and U4241 (N_4241,N_2460,N_3008);
or U4242 (N_4242,N_2893,N_3663);
or U4243 (N_4243,N_2192,N_2491);
xor U4244 (N_4244,N_2820,N_3490);
xnor U4245 (N_4245,N_3715,N_3274);
nand U4246 (N_4246,N_2584,N_3991);
nand U4247 (N_4247,N_3365,N_2217);
nand U4248 (N_4248,N_3497,N_3830);
and U4249 (N_4249,N_3066,N_2985);
or U4250 (N_4250,N_2909,N_2607);
or U4251 (N_4251,N_3861,N_3297);
nor U4252 (N_4252,N_3099,N_2568);
and U4253 (N_4253,N_2737,N_2099);
nand U4254 (N_4254,N_3907,N_3723);
nor U4255 (N_4255,N_3402,N_2949);
nor U4256 (N_4256,N_2950,N_3785);
and U4257 (N_4257,N_3052,N_2007);
nor U4258 (N_4258,N_3114,N_3783);
nand U4259 (N_4259,N_3505,N_2790);
nand U4260 (N_4260,N_3238,N_3154);
nor U4261 (N_4261,N_2598,N_2002);
nand U4262 (N_4262,N_2215,N_3900);
or U4263 (N_4263,N_2885,N_3180);
nand U4264 (N_4264,N_3828,N_2362);
nand U4265 (N_4265,N_2288,N_2065);
nor U4266 (N_4266,N_3648,N_2423);
or U4267 (N_4267,N_3771,N_3482);
nor U4268 (N_4268,N_2588,N_2212);
xor U4269 (N_4269,N_2999,N_3351);
xor U4270 (N_4270,N_2147,N_3191);
nor U4271 (N_4271,N_2980,N_2906);
or U4272 (N_4272,N_2630,N_2880);
nor U4273 (N_4273,N_2913,N_3276);
and U4274 (N_4274,N_3928,N_2996);
nand U4275 (N_4275,N_3432,N_2359);
and U4276 (N_4276,N_3252,N_3210);
xnor U4277 (N_4277,N_2624,N_3636);
nor U4278 (N_4278,N_2580,N_3984);
xor U4279 (N_4279,N_2161,N_3237);
xnor U4280 (N_4280,N_2937,N_2805);
nor U4281 (N_4281,N_3736,N_2992);
or U4282 (N_4282,N_2629,N_3270);
and U4283 (N_4283,N_3621,N_3062);
nor U4284 (N_4284,N_3522,N_3220);
nor U4285 (N_4285,N_3691,N_3899);
and U4286 (N_4286,N_2533,N_3379);
nand U4287 (N_4287,N_2543,N_2049);
nor U4288 (N_4288,N_3914,N_3129);
xor U4289 (N_4289,N_2708,N_2082);
nand U4290 (N_4290,N_2687,N_3562);
xnor U4291 (N_4291,N_2402,N_3311);
and U4292 (N_4292,N_2311,N_3994);
nand U4293 (N_4293,N_3132,N_3248);
nand U4294 (N_4294,N_3475,N_3013);
and U4295 (N_4295,N_3335,N_3824);
nor U4296 (N_4296,N_2775,N_2354);
or U4297 (N_4297,N_2904,N_3577);
nand U4298 (N_4298,N_2272,N_2081);
and U4299 (N_4299,N_3022,N_2995);
and U4300 (N_4300,N_3769,N_2113);
or U4301 (N_4301,N_2248,N_3451);
nand U4302 (N_4302,N_2070,N_2383);
or U4303 (N_4303,N_2868,N_3637);
and U4304 (N_4304,N_2056,N_2570);
nor U4305 (N_4305,N_3877,N_3121);
xnor U4306 (N_4306,N_3716,N_3866);
nand U4307 (N_4307,N_3083,N_2750);
and U4308 (N_4308,N_3165,N_2721);
and U4309 (N_4309,N_2315,N_3755);
or U4310 (N_4310,N_3169,N_3879);
nand U4311 (N_4311,N_3665,N_2812);
nor U4312 (N_4312,N_2652,N_3115);
nor U4313 (N_4313,N_2676,N_2743);
nor U4314 (N_4314,N_3437,N_3550);
nand U4315 (N_4315,N_3959,N_3086);
and U4316 (N_4316,N_3152,N_2300);
and U4317 (N_4317,N_3367,N_3125);
or U4318 (N_4318,N_2975,N_2798);
xor U4319 (N_4319,N_3339,N_2170);
or U4320 (N_4320,N_2398,N_2903);
nand U4321 (N_4321,N_3492,N_2637);
or U4322 (N_4322,N_3355,N_3652);
nand U4323 (N_4323,N_2902,N_3000);
nor U4324 (N_4324,N_3662,N_2674);
or U4325 (N_4325,N_2105,N_2596);
and U4326 (N_4326,N_3499,N_2238);
nor U4327 (N_4327,N_3847,N_2422);
nand U4328 (N_4328,N_2696,N_2023);
or U4329 (N_4329,N_2339,N_2468);
nor U4330 (N_4330,N_3153,N_2892);
and U4331 (N_4331,N_2384,N_2371);
nand U4332 (N_4332,N_2894,N_2124);
nand U4333 (N_4333,N_2647,N_3963);
and U4334 (N_4334,N_2693,N_3489);
xnor U4335 (N_4335,N_3881,N_3909);
nor U4336 (N_4336,N_2529,N_2621);
nand U4337 (N_4337,N_3296,N_2911);
and U4338 (N_4338,N_3161,N_3005);
nand U4339 (N_4339,N_3167,N_3313);
nand U4340 (N_4340,N_3646,N_3587);
nand U4341 (N_4341,N_2648,N_2134);
or U4342 (N_4342,N_2781,N_3190);
or U4343 (N_4343,N_3332,N_2947);
nor U4344 (N_4344,N_3978,N_2695);
nor U4345 (N_4345,N_2851,N_3768);
nand U4346 (N_4346,N_3511,N_2520);
and U4347 (N_4347,N_2654,N_2627);
xnor U4348 (N_4348,N_2455,N_2269);
nor U4349 (N_4349,N_2766,N_2622);
nand U4350 (N_4350,N_3572,N_2746);
and U4351 (N_4351,N_2592,N_3057);
nor U4352 (N_4352,N_3608,N_2528);
or U4353 (N_4353,N_3922,N_3221);
xnor U4354 (N_4354,N_2717,N_3752);
xor U4355 (N_4355,N_3168,N_3413);
or U4356 (N_4356,N_2655,N_3625);
nor U4357 (N_4357,N_2232,N_2279);
or U4358 (N_4358,N_3240,N_2479);
or U4359 (N_4359,N_3804,N_3094);
and U4360 (N_4360,N_3342,N_3109);
nand U4361 (N_4361,N_2874,N_2565);
nand U4362 (N_4362,N_3408,N_3607);
nor U4363 (N_4363,N_2295,N_2649);
xor U4364 (N_4364,N_2686,N_2641);
and U4365 (N_4365,N_3706,N_2378);
and U4366 (N_4366,N_3181,N_3374);
xnor U4367 (N_4367,N_3873,N_3593);
or U4368 (N_4368,N_2336,N_3176);
nand U4369 (N_4369,N_2234,N_3333);
or U4370 (N_4370,N_3993,N_3443);
nor U4371 (N_4371,N_2751,N_3669);
nand U4372 (N_4372,N_2972,N_3775);
nand U4373 (N_4373,N_3781,N_2429);
and U4374 (N_4374,N_3259,N_3690);
and U4375 (N_4375,N_2394,N_3015);
or U4376 (N_4376,N_3048,N_3456);
xor U4377 (N_4377,N_2807,N_3846);
and U4378 (N_4378,N_3540,N_3854);
nand U4379 (N_4379,N_3676,N_3471);
nand U4380 (N_4380,N_3547,N_2967);
nand U4381 (N_4381,N_2532,N_2360);
or U4382 (N_4382,N_2611,N_3503);
xnor U4383 (N_4383,N_3657,N_3362);
and U4384 (N_4384,N_3935,N_2857);
nand U4385 (N_4385,N_3695,N_2296);
nand U4386 (N_4386,N_2284,N_2600);
nand U4387 (N_4387,N_2287,N_2822);
and U4388 (N_4388,N_2285,N_2233);
and U4389 (N_4389,N_2003,N_3815);
and U4390 (N_4390,N_2752,N_2942);
nor U4391 (N_4391,N_3467,N_3921);
or U4392 (N_4392,N_3556,N_3122);
nor U4393 (N_4393,N_3184,N_3278);
nor U4394 (N_4394,N_2877,N_2177);
and U4395 (N_4395,N_2955,N_2542);
nor U4396 (N_4396,N_3581,N_2026);
nor U4397 (N_4397,N_2841,N_2055);
and U4398 (N_4398,N_2970,N_2101);
nor U4399 (N_4399,N_3892,N_3685);
or U4400 (N_4400,N_3740,N_3072);
or U4401 (N_4401,N_3014,N_2433);
xor U4402 (N_4402,N_3638,N_3183);
nor U4403 (N_4403,N_3853,N_2306);
or U4404 (N_4404,N_3656,N_2771);
nor U4405 (N_4405,N_3823,N_3887);
nor U4406 (N_4406,N_2243,N_2956);
nand U4407 (N_4407,N_3751,N_2213);
and U4408 (N_4408,N_2036,N_3087);
and U4409 (N_4409,N_2392,N_3660);
nand U4410 (N_4410,N_3949,N_3481);
or U4411 (N_4411,N_2118,N_3447);
and U4412 (N_4412,N_3584,N_2540);
and U4413 (N_4413,N_3520,N_2921);
nand U4414 (N_4414,N_2348,N_2830);
or U4415 (N_4415,N_2457,N_3383);
nor U4416 (N_4416,N_2505,N_3291);
and U4417 (N_4417,N_3356,N_2236);
and U4418 (N_4418,N_3399,N_2223);
or U4419 (N_4419,N_2088,N_3067);
nand U4420 (N_4420,N_2516,N_2252);
and U4421 (N_4421,N_3207,N_3886);
nor U4422 (N_4422,N_2175,N_2486);
and U4423 (N_4423,N_2268,N_2095);
nand U4424 (N_4424,N_2120,N_2130);
or U4425 (N_4425,N_3127,N_2635);
nand U4426 (N_4426,N_3536,N_3093);
nor U4427 (N_4427,N_2037,N_2699);
nand U4428 (N_4428,N_3971,N_3947);
nand U4429 (N_4429,N_2106,N_2561);
nand U4430 (N_4430,N_2261,N_3026);
nand U4431 (N_4431,N_3400,N_2211);
or U4432 (N_4432,N_2145,N_2176);
or U4433 (N_4433,N_2941,N_3284);
or U4434 (N_4434,N_3271,N_3765);
xnor U4435 (N_4435,N_2158,N_3060);
or U4436 (N_4436,N_2744,N_2163);
nand U4437 (N_4437,N_3146,N_2774);
and U4438 (N_4438,N_2193,N_2421);
nor U4439 (N_4439,N_3982,N_2432);
nor U4440 (N_4440,N_3890,N_3842);
nor U4441 (N_4441,N_2554,N_2375);
nand U4442 (N_4442,N_3147,N_2385);
nor U4443 (N_4443,N_3418,N_2682);
and U4444 (N_4444,N_2571,N_3732);
or U4445 (N_4445,N_3610,N_3193);
nand U4446 (N_4446,N_3756,N_2834);
or U4447 (N_4447,N_3627,N_2675);
and U4448 (N_4448,N_3537,N_2666);
or U4449 (N_4449,N_2816,N_2139);
and U4450 (N_4450,N_2811,N_2489);
and U4451 (N_4451,N_2334,N_2638);
or U4452 (N_4452,N_3519,N_3302);
and U4453 (N_4453,N_2060,N_2051);
or U4454 (N_4454,N_2604,N_3863);
and U4455 (N_4455,N_3050,N_2809);
or U4456 (N_4456,N_2500,N_3195);
or U4457 (N_4457,N_2764,N_2610);
or U4458 (N_4458,N_3182,N_2184);
nand U4459 (N_4459,N_2918,N_2558);
or U4460 (N_4460,N_2689,N_2842);
nor U4461 (N_4461,N_2390,N_3507);
nor U4462 (N_4462,N_3187,N_2404);
and U4463 (N_4463,N_2444,N_2644);
nor U4464 (N_4464,N_3944,N_2439);
and U4465 (N_4465,N_2803,N_2968);
nor U4466 (N_4466,N_2861,N_3972);
nand U4467 (N_4467,N_3415,N_2690);
nor U4468 (N_4468,N_2364,N_3934);
nor U4469 (N_4469,N_2199,N_2912);
xor U4470 (N_4470,N_3188,N_2701);
and U4471 (N_4471,N_2915,N_3603);
nand U4472 (N_4472,N_3609,N_3565);
xnor U4473 (N_4473,N_3144,N_2289);
nand U4474 (N_4474,N_3300,N_3840);
or U4475 (N_4475,N_2934,N_2788);
nand U4476 (N_4476,N_2393,N_2149);
xnor U4477 (N_4477,N_2480,N_3453);
xnor U4478 (N_4478,N_3488,N_2258);
nor U4479 (N_4479,N_3388,N_3757);
and U4480 (N_4480,N_3450,N_2125);
or U4481 (N_4481,N_2152,N_3101);
xor U4482 (N_4482,N_3517,N_3640);
nand U4483 (N_4483,N_3306,N_3137);
and U4484 (N_4484,N_2792,N_3702);
and U4485 (N_4485,N_3813,N_3538);
nor U4486 (N_4486,N_2663,N_3502);
and U4487 (N_4487,N_2219,N_3055);
nand U4488 (N_4488,N_3226,N_2408);
or U4489 (N_4489,N_3200,N_2691);
and U4490 (N_4490,N_2302,N_2399);
or U4491 (N_4491,N_3712,N_2856);
xor U4492 (N_4492,N_2828,N_3960);
nand U4493 (N_4493,N_2366,N_2800);
and U4494 (N_4494,N_3315,N_2274);
nor U4495 (N_4495,N_3604,N_3024);
xor U4496 (N_4496,N_3197,N_2569);
nor U4497 (N_4497,N_2389,N_3464);
and U4498 (N_4498,N_2664,N_3438);
and U4499 (N_4499,N_3864,N_3231);
xnor U4500 (N_4500,N_3244,N_2550);
nor U4501 (N_4501,N_3051,N_3222);
and U4502 (N_4502,N_2875,N_3076);
nor U4503 (N_4503,N_2661,N_3737);
nor U4504 (N_4504,N_3626,N_2262);
nand U4505 (N_4505,N_2016,N_3021);
and U4506 (N_4506,N_2022,N_3251);
nor U4507 (N_4507,N_2114,N_3860);
or U4508 (N_4508,N_3243,N_3778);
or U4509 (N_4509,N_3896,N_2443);
nand U4510 (N_4510,N_2920,N_3770);
nor U4511 (N_4511,N_3990,N_3309);
xnor U4512 (N_4512,N_2356,N_3616);
or U4513 (N_4513,N_3631,N_2136);
nor U4514 (N_4514,N_2756,N_2168);
nand U4515 (N_4515,N_3185,N_2507);
and U4516 (N_4516,N_3324,N_3422);
or U4517 (N_4517,N_2733,N_3233);
and U4518 (N_4518,N_2410,N_3260);
nand U4519 (N_4519,N_2710,N_3257);
and U4520 (N_4520,N_3827,N_2786);
or U4521 (N_4521,N_2724,N_2010);
or U4522 (N_4522,N_3521,N_3875);
xor U4523 (N_4523,N_3016,N_3140);
nand U4524 (N_4524,N_3931,N_2165);
nor U4525 (N_4525,N_2732,N_3833);
nor U4526 (N_4526,N_2562,N_2555);
nor U4527 (N_4527,N_3987,N_2191);
nor U4528 (N_4528,N_2535,N_2254);
and U4529 (N_4529,N_2818,N_2198);
nor U4530 (N_4530,N_2971,N_3997);
nand U4531 (N_4531,N_3601,N_3677);
or U4532 (N_4532,N_3295,N_3196);
nor U4533 (N_4533,N_2636,N_2943);
or U4534 (N_4534,N_3826,N_3498);
and U4535 (N_4535,N_2878,N_3174);
nand U4536 (N_4536,N_3470,N_2386);
and U4537 (N_4537,N_3419,N_3417);
nor U4538 (N_4538,N_3045,N_3156);
or U4539 (N_4539,N_2374,N_2471);
nand U4540 (N_4540,N_3561,N_3976);
and U4541 (N_4541,N_3901,N_2239);
or U4542 (N_4542,N_3957,N_3739);
nand U4543 (N_4543,N_3795,N_2866);
nor U4544 (N_4544,N_3844,N_3177);
nand U4545 (N_4545,N_3655,N_3675);
and U4546 (N_4546,N_2484,N_2018);
nor U4547 (N_4547,N_3485,N_3301);
xnor U4548 (N_4548,N_2539,N_3895);
or U4549 (N_4549,N_3910,N_2453);
and U4550 (N_4550,N_3246,N_3611);
and U4551 (N_4551,N_2204,N_3925);
or U4552 (N_4552,N_3133,N_3164);
or U4553 (N_4553,N_3010,N_3092);
xor U4554 (N_4554,N_3407,N_2498);
and U4555 (N_4555,N_3682,N_3330);
xor U4556 (N_4556,N_3004,N_2221);
and U4557 (N_4557,N_2897,N_2052);
or U4558 (N_4558,N_2146,N_3411);
and U4559 (N_4559,N_2576,N_3258);
nand U4560 (N_4560,N_3684,N_3670);
or U4561 (N_4561,N_3760,N_3508);
or U4562 (N_4562,N_3163,N_3241);
nand U4563 (N_4563,N_3649,N_3793);
and U4564 (N_4564,N_2320,N_3870);
nand U4565 (N_4565,N_2041,N_2631);
and U4566 (N_4566,N_3557,N_2890);
and U4567 (N_4567,N_3988,N_2442);
and U4568 (N_4568,N_3906,N_2178);
nor U4569 (N_4569,N_3290,N_2933);
and U4570 (N_4570,N_3791,N_2938);
or U4571 (N_4571,N_2397,N_3835);
and U4572 (N_4572,N_2420,N_3328);
and U4573 (N_4573,N_3920,N_2632);
and U4574 (N_4574,N_3618,N_3956);
nor U4575 (N_4575,N_2898,N_2142);
or U4576 (N_4576,N_2387,N_3261);
or U4577 (N_4577,N_3532,N_2859);
and U4578 (N_4578,N_2963,N_3205);
xor U4579 (N_4579,N_2133,N_2729);
or U4580 (N_4580,N_3401,N_3951);
xnor U4581 (N_4581,N_2983,N_2723);
nor U4582 (N_4582,N_2226,N_3445);
nor U4583 (N_4583,N_3798,N_3030);
nand U4584 (N_4584,N_3859,N_3579);
nor U4585 (N_4585,N_2006,N_2726);
nand U4586 (N_4586,N_2048,N_2575);
and U4587 (N_4587,N_3945,N_3227);
nand U4588 (N_4588,N_2824,N_2548);
nor U4589 (N_4589,N_3494,N_3533);
nor U4590 (N_4590,N_3554,N_2777);
and U4591 (N_4591,N_3228,N_2029);
nor U4592 (N_4592,N_2119,N_3635);
or U4593 (N_4593,N_2053,N_3724);
or U4594 (N_4594,N_3985,N_2148);
nand U4595 (N_4595,N_3002,N_2640);
nand U4596 (N_4596,N_2169,N_3343);
and U4597 (N_4597,N_2650,N_3466);
nand U4598 (N_4598,N_2589,N_3082);
and U4599 (N_4599,N_3336,N_2634);
nor U4600 (N_4600,N_3398,N_3403);
nor U4601 (N_4601,N_3387,N_3880);
and U4602 (N_4602,N_2951,N_3224);
and U4603 (N_4603,N_2100,N_2205);
nand U4604 (N_4604,N_2494,N_2616);
or U4605 (N_4605,N_3145,N_3698);
nand U4606 (N_4606,N_2521,N_2618);
xnor U4607 (N_4607,N_3420,N_3776);
nand U4608 (N_4608,N_3806,N_3653);
and U4609 (N_4609,N_3166,N_2735);
nand U4610 (N_4610,N_2519,N_2319);
xor U4611 (N_4611,N_2259,N_2984);
and U4612 (N_4612,N_2365,N_2503);
or U4613 (N_4613,N_2112,N_2988);
and U4614 (N_4614,N_3266,N_2888);
nand U4615 (N_4615,N_3856,N_2741);
xnor U4616 (N_4616,N_3697,N_3433);
nand U4617 (N_4617,N_2895,N_2739);
or U4618 (N_4618,N_2501,N_3954);
and U4619 (N_4619,N_3427,N_3267);
or U4620 (N_4620,N_2511,N_3747);
nand U4621 (N_4621,N_3605,N_3696);
or U4622 (N_4622,N_2090,N_3595);
nand U4623 (N_4623,N_2126,N_3159);
xor U4624 (N_4624,N_2075,N_2964);
and U4625 (N_4625,N_2952,N_2325);
xnor U4626 (N_4626,N_3995,N_3468);
nor U4627 (N_4627,N_3484,N_2910);
or U4628 (N_4628,N_3617,N_2711);
or U4629 (N_4629,N_2063,N_3170);
or U4630 (N_4630,N_3759,N_3992);
nand U4631 (N_4631,N_2414,N_3692);
nand U4632 (N_4632,N_2698,N_3566);
nor U4633 (N_4633,N_3659,N_2174);
or U4634 (N_4634,N_2791,N_3097);
or U4635 (N_4635,N_3622,N_3431);
xor U4636 (N_4636,N_3748,N_2309);
and U4637 (N_4637,N_2742,N_2316);
and U4638 (N_4638,N_3102,N_2340);
or U4639 (N_4639,N_3592,N_3967);
and U4640 (N_4640,N_2860,N_2190);
and U4641 (N_4641,N_3961,N_2020);
or U4642 (N_4642,N_3738,N_3893);
nand U4643 (N_4643,N_2579,N_2128);
nand U4644 (N_4644,N_3491,N_3380);
nor U4645 (N_4645,N_2896,N_3465);
nor U4646 (N_4646,N_3782,N_2312);
or U4647 (N_4647,N_2102,N_3571);
or U4648 (N_4648,N_2763,N_2759);
nor U4649 (N_4649,N_3444,N_3926);
and U4650 (N_4650,N_3891,N_2730);
nor U4651 (N_4651,N_3529,N_3119);
and U4652 (N_4652,N_2154,N_2046);
nand U4653 (N_4653,N_3155,N_3745);
nand U4654 (N_4654,N_2814,N_3817);
and U4655 (N_4655,N_3658,N_3007);
and U4656 (N_4656,N_2406,N_2923);
or U4657 (N_4657,N_3299,N_2832);
xor U4658 (N_4658,N_3317,N_2784);
and U4659 (N_4659,N_2987,N_2425);
and U4660 (N_4660,N_3361,N_2590);
xnor U4661 (N_4661,N_2712,N_2839);
nand U4662 (N_4662,N_3404,N_2044);
nand U4663 (N_4663,N_2989,N_2143);
and U4664 (N_4664,N_3708,N_3671);
or U4665 (N_4665,N_3686,N_2475);
xnor U4666 (N_4666,N_2506,N_3268);
or U4667 (N_4667,N_2510,N_3851);
and U4668 (N_4668,N_3933,N_3329);
nand U4669 (N_4669,N_2476,N_3192);
and U4670 (N_4670,N_2188,N_2908);
and U4671 (N_4671,N_2173,N_2703);
nor U4672 (N_4672,N_2587,N_2195);
nand U4673 (N_4673,N_3888,N_3334);
and U4674 (N_4674,N_3962,N_3459);
nor U4675 (N_4675,N_3116,N_3327);
nand U4676 (N_4676,N_3234,N_2709);
and U4677 (N_4677,N_3304,N_3915);
or U4678 (N_4678,N_3878,N_3849);
nand U4679 (N_4679,N_2349,N_3100);
nand U4680 (N_4680,N_2203,N_3968);
nor U4681 (N_4681,N_3378,N_3364);
xor U4682 (N_4682,N_3941,N_3764);
and U4683 (N_4683,N_2167,N_2847);
or U4684 (N_4684,N_3043,N_2986);
and U4685 (N_4685,N_2253,N_3903);
or U4686 (N_4686,N_3672,N_2882);
nand U4687 (N_4687,N_3558,N_3366);
and U4688 (N_4688,N_3814,N_2653);
nor U4689 (N_4689,N_3539,N_2246);
or U4690 (N_4690,N_2483,N_3292);
or U4691 (N_4691,N_2625,N_2054);
nand U4692 (N_4692,N_2917,N_2922);
or U4693 (N_4693,N_3679,N_2067);
nand U4694 (N_4694,N_3799,N_3029);
nor U4695 (N_4695,N_2076,N_3111);
nand U4696 (N_4696,N_2064,N_2305);
and U4697 (N_4697,N_3728,N_3118);
or U4698 (N_4698,N_3081,N_3913);
nand U4699 (N_4699,N_3338,N_2094);
and U4700 (N_4700,N_2960,N_2981);
xor U4701 (N_4701,N_2706,N_2108);
nor U4702 (N_4702,N_2597,N_3735);
and U4703 (N_4703,N_3372,N_3699);
nor U4704 (N_4704,N_3634,N_3710);
and U4705 (N_4705,N_3711,N_2994);
nor U4706 (N_4706,N_2731,N_3496);
or U4707 (N_4707,N_3784,N_2039);
or U4708 (N_4708,N_3139,N_2009);
and U4709 (N_4709,N_2015,N_3084);
nand U4710 (N_4710,N_2545,N_2734);
and U4711 (N_4711,N_3726,N_3157);
or U4712 (N_4712,N_2840,N_2440);
and U4713 (N_4713,N_3948,N_2767);
and U4714 (N_4714,N_3544,N_3986);
nand U4715 (N_4715,N_3056,N_3255);
and U4716 (N_4716,N_2380,N_2074);
and U4717 (N_4717,N_2831,N_2948);
and U4718 (N_4718,N_3514,N_2216);
xnor U4719 (N_4719,N_2235,N_3559);
nand U4720 (N_4720,N_3229,N_3344);
or U4721 (N_4721,N_2071,N_2299);
xor U4722 (N_4722,N_2214,N_3312);
nand U4723 (N_4723,N_2872,N_3789);
or U4724 (N_4724,N_2337,N_2515);
and U4725 (N_4725,N_2121,N_2338);
or U4726 (N_4726,N_2448,N_3473);
and U4727 (N_4727,N_2372,N_3578);
xor U4728 (N_4728,N_2601,N_3628);
nor U4729 (N_4729,N_2657,N_2424);
xor U4730 (N_4730,N_3288,N_2482);
and U4731 (N_4731,N_3041,N_3980);
nand U4732 (N_4732,N_2718,N_2713);
nand U4733 (N_4733,N_2012,N_3575);
nor U4734 (N_4734,N_2369,N_3819);
or U4735 (N_4735,N_3019,N_2773);
and U4736 (N_4736,N_3262,N_3567);
nand U4737 (N_4737,N_2220,N_3020);
and U4738 (N_4738,N_3406,N_2969);
and U4739 (N_4739,N_2692,N_3958);
nor U4740 (N_4740,N_3442,N_3916);
nand U4741 (N_4741,N_3867,N_2183);
or U4742 (N_4742,N_2162,N_3073);
xnor U4743 (N_4743,N_3047,N_3845);
nand U4744 (N_4744,N_2407,N_2619);
nor U4745 (N_4745,N_3282,N_2749);
and U4746 (N_4746,N_2583,N_2412);
nor U4747 (N_4747,N_2787,N_3837);
nand U4748 (N_4748,N_2209,N_3718);
nand U4749 (N_4749,N_3613,N_3036);
nand U4750 (N_4750,N_3753,N_3973);
or U4751 (N_4751,N_2472,N_3198);
nor U4752 (N_4752,N_2115,N_2669);
or U4753 (N_4753,N_2530,N_2517);
and U4754 (N_4754,N_3644,N_3590);
and U4755 (N_4755,N_3766,N_3235);
nor U4756 (N_4756,N_3869,N_3583);
xnor U4757 (N_4757,N_3104,N_2497);
nor U4758 (N_4758,N_2156,N_2021);
nand U4759 (N_4759,N_3709,N_3848);
xor U4760 (N_4760,N_3871,N_3884);
nand U4761 (N_4761,N_3095,N_2779);
and U4762 (N_4762,N_2544,N_2901);
and U4763 (N_4763,N_3746,N_2255);
nand U4764 (N_4764,N_3321,N_2292);
and U4765 (N_4765,N_2179,N_2314);
and U4766 (N_4766,N_3006,N_2566);
or U4767 (N_4767,N_2714,N_3850);
or U4768 (N_4768,N_2182,N_2388);
and U4769 (N_4769,N_2835,N_2208);
nand U4770 (N_4770,N_2153,N_3394);
nand U4771 (N_4771,N_2602,N_2796);
nand U4772 (N_4772,N_2683,N_3435);
or U4773 (N_4773,N_2263,N_2431);
and U4774 (N_4774,N_2466,N_2957);
and U4775 (N_4775,N_2907,N_3075);
nor U4776 (N_4776,N_3688,N_3858);
or U4777 (N_4777,N_3079,N_3236);
and U4778 (N_4778,N_2194,N_3171);
nor U4779 (N_4779,N_2050,N_2524);
or U4780 (N_4780,N_3970,N_3825);
and U4781 (N_4781,N_2925,N_2083);
nor U4782 (N_4782,N_3088,N_2267);
nor U4783 (N_4783,N_2694,N_2474);
and U4784 (N_4784,N_3209,N_2838);
nor U4785 (N_4785,N_2595,N_2073);
xor U4786 (N_4786,N_3203,N_2585);
nor U4787 (N_4787,N_3053,N_3025);
and U4788 (N_4788,N_3303,N_2346);
and U4789 (N_4789,N_2335,N_3028);
xor U4790 (N_4790,N_2454,N_2062);
nand U4791 (N_4791,N_3275,N_2140);
and U4792 (N_4792,N_3307,N_2485);
and U4793 (N_4793,N_3513,N_2428);
nor U4794 (N_4794,N_2808,N_3345);
and U4795 (N_4795,N_3942,N_2785);
xnor U4796 (N_4796,N_2104,N_2286);
nor U4797 (N_4797,N_3409,N_2096);
and U4798 (N_4798,N_2207,N_3810);
xnor U4799 (N_4799,N_2549,N_2240);
nand U4800 (N_4800,N_2884,N_2795);
or U4801 (N_4801,N_3011,N_3836);
or U4802 (N_4802,N_3952,N_2229);
or U4803 (N_4803,N_2225,N_3531);
nor U4804 (N_4804,N_3396,N_2642);
xor U4805 (N_4805,N_3230,N_3950);
or U4806 (N_4806,N_2492,N_3085);
and U4807 (N_4807,N_3523,N_3518);
nand U4808 (N_4808,N_2982,N_3136);
xnor U4809 (N_4809,N_3263,N_2702);
or U4810 (N_4810,N_3286,N_2450);
nand U4811 (N_4811,N_3386,N_2553);
or U4812 (N_4812,N_3455,N_3423);
nand U4813 (N_4813,N_3357,N_2200);
or U4814 (N_4814,N_3719,N_2536);
nor U4815 (N_4815,N_3373,N_2546);
or U4816 (N_4816,N_3889,N_3705);
or U4817 (N_4817,N_3839,N_2753);
or U4818 (N_4818,N_3393,N_2245);
or U4819 (N_4819,N_2181,N_3368);
xnor U4820 (N_4820,N_3943,N_3426);
nand U4821 (N_4821,N_3202,N_2451);
nand U4822 (N_4822,N_2490,N_3232);
nand U4823 (N_4823,N_3923,N_3218);
or U4824 (N_4824,N_3902,N_2679);
or U4825 (N_4825,N_3012,N_3385);
xnor U4826 (N_4826,N_2883,N_3434);
nor U4827 (N_4827,N_3786,N_2089);
xnor U4828 (N_4828,N_3217,N_3541);
nand U4829 (N_4829,N_2821,N_2973);
nor U4830 (N_4830,N_3929,N_2736);
or U4831 (N_4831,N_2887,N_2344);
nor U4832 (N_4832,N_3440,N_3597);
nand U4833 (N_4833,N_2801,N_2069);
xor U4834 (N_4834,N_3969,N_2463);
or U4835 (N_4835,N_3381,N_2826);
xnor U4836 (N_4836,N_2836,N_2196);
xnor U4837 (N_4837,N_3247,N_2673);
nand U4838 (N_4838,N_3535,N_2324);
and U4839 (N_4839,N_2355,N_2656);
xor U4840 (N_4840,N_2612,N_2465);
or U4841 (N_4841,N_2343,N_2322);
nand U4842 (N_4842,N_3392,N_2132);
and U4843 (N_4843,N_2547,N_3713);
nor U4844 (N_4844,N_2930,N_3563);
or U4845 (N_4845,N_2855,N_3865);
nor U4846 (N_4846,N_3965,N_2613);
nor U4847 (N_4847,N_3927,N_3730);
and U4848 (N_4848,N_3585,N_3744);
nand U4849 (N_4849,N_3322,N_3841);
nand U4850 (N_4850,N_2273,N_3700);
xor U4851 (N_4851,N_3568,N_2783);
nor U4852 (N_4852,N_3206,N_3936);
nand U4853 (N_4853,N_2157,N_2867);
nor U4854 (N_4854,N_3353,N_2560);
nand U4855 (N_4855,N_2059,N_3201);
nor U4856 (N_4856,N_3141,N_2707);
and U4857 (N_4857,N_2837,N_3289);
xor U4858 (N_4858,N_3212,N_3360);
nor U4859 (N_4859,N_3542,N_2373);
nor U4860 (N_4860,N_3138,N_2504);
or U4861 (N_4861,N_2377,N_3080);
and U4862 (N_4862,N_2541,N_2684);
nand U4863 (N_4863,N_3549,N_2265);
or U4864 (N_4864,N_2747,N_3017);
or U4865 (N_4865,N_2231,N_3955);
and U4866 (N_4866,N_2929,N_2030);
or U4867 (N_4867,N_2237,N_3256);
xor U4868 (N_4868,N_3281,N_2582);
nand U4869 (N_4869,N_2488,N_3642);
xnor U4870 (N_4870,N_2603,N_3912);
or U4871 (N_4871,N_3316,N_3811);
nand U4872 (N_4872,N_3516,N_2304);
nor U4873 (N_4873,N_3463,N_2107);
and U4874 (N_4874,N_2499,N_3725);
nor U4875 (N_4875,N_3215,N_3551);
nand U4876 (N_4876,N_2326,N_3298);
and U4877 (N_4877,N_2426,N_2321);
nand U4878 (N_4878,N_3683,N_3937);
nand U4879 (N_4879,N_3142,N_2084);
or U4880 (N_4880,N_3673,N_2066);
nor U4881 (N_4881,N_3704,N_3946);
nand U4882 (N_4882,N_3318,N_3524);
or U4883 (N_4883,N_2155,N_2318);
nand U4884 (N_4884,N_3742,N_3405);
and U4885 (N_4885,N_3070,N_2806);
and U4886 (N_4886,N_3287,N_2122);
xor U4887 (N_4887,N_3894,N_3620);
xor U4888 (N_4888,N_2464,N_2277);
nor U4889 (N_4889,N_2537,N_3410);
nand U4890 (N_4890,N_3425,N_3999);
and U4891 (N_4891,N_3932,N_2411);
and U4892 (N_4892,N_3883,N_2230);
nand U4893 (N_4893,N_3091,N_2738);
and U4894 (N_4894,N_2109,N_3370);
xor U4895 (N_4895,N_2758,N_2396);
nand U4896 (N_4896,N_2662,N_3349);
xnor U4897 (N_4897,N_2932,N_2620);
nand U4898 (N_4898,N_3216,N_2137);
nand U4899 (N_4899,N_3796,N_2144);
and U4900 (N_4900,N_3294,N_3105);
or U4901 (N_4901,N_3395,N_2227);
nor U4902 (N_4902,N_2862,N_2993);
nor U4903 (N_4903,N_2815,N_2418);
and U4904 (N_4904,N_2379,N_3602);
or U4905 (N_4905,N_2160,N_2858);
and U4906 (N_4906,N_2810,N_3032);
nand U4907 (N_4907,N_3194,N_2456);
nand U4908 (N_4908,N_2797,N_3643);
and U4909 (N_4909,N_2415,N_2313);
xnor U4910 (N_4910,N_2079,N_2833);
nand U4911 (N_4911,N_3358,N_3208);
xnor U4912 (N_4912,N_3843,N_2962);
nand U4913 (N_4913,N_3803,N_2307);
xor U4914 (N_4914,N_3573,N_3998);
nor U4915 (N_4915,N_3414,N_3591);
or U4916 (N_4916,N_3647,N_3023);
nand U4917 (N_4917,N_3787,N_3049);
and U4918 (N_4918,N_2187,N_2865);
nor U4919 (N_4919,N_3750,N_2441);
nor U4920 (N_4920,N_2802,N_2697);
or U4921 (N_4921,N_2850,N_3199);
nand U4922 (N_4922,N_3160,N_2332);
or U4923 (N_4923,N_2658,N_2889);
and U4924 (N_4924,N_2705,N_3772);
nor U4925 (N_4925,N_2538,N_2347);
and U4926 (N_4926,N_2881,N_2793);
xnor U4927 (N_4927,N_2185,N_3774);
nor U4928 (N_4928,N_2481,N_3681);
nor U4929 (N_4929,N_2210,N_3448);
xor U4930 (N_4930,N_2024,N_3446);
xor U4931 (N_4931,N_2978,N_3478);
nand U4932 (N_4932,N_2042,N_3457);
and U4933 (N_4933,N_2776,N_3347);
nand U4934 (N_4934,N_3421,N_2617);
and U4935 (N_4935,N_3729,N_3106);
and U4936 (N_4936,N_2367,N_3807);
or U4937 (N_4937,N_2879,N_2522);
or U4938 (N_4938,N_2899,N_2038);
nand U4939 (N_4939,N_2564,N_3249);
xor U4940 (N_4940,N_3974,N_3707);
nor U4941 (N_4941,N_2434,N_2514);
nor U4942 (N_4942,N_3808,N_2291);
or U4943 (N_4943,N_3606,N_2222);
and U4944 (N_4944,N_3898,N_2092);
and U4945 (N_4945,N_2057,N_2436);
and U4946 (N_4946,N_3204,N_2470);
xnor U4947 (N_4947,N_3452,N_3480);
or U4948 (N_4948,N_2164,N_3589);
nand U4949 (N_4949,N_2871,N_3802);
or U4950 (N_4950,N_3734,N_2045);
nor U4951 (N_4951,N_3348,N_3801);
and U4952 (N_4952,N_3280,N_2278);
and U4953 (N_4953,N_3818,N_3143);
nor U4954 (N_4954,N_2469,N_2979);
xor U4955 (N_4955,N_2924,N_2748);
xnor U4956 (N_4956,N_3487,N_2301);
nand U4957 (N_4957,N_2435,N_2876);
xnor U4958 (N_4958,N_2097,N_2760);
nand U4959 (N_4959,N_3820,N_2594);
xor U4960 (N_4960,N_2116,N_3722);
nand U4961 (N_4961,N_3223,N_3834);
nor U4962 (N_4962,N_2141,N_2001);
xnor U4963 (N_4963,N_2078,N_2224);
nor U4964 (N_4964,N_3483,N_3285);
and U4965 (N_4965,N_2013,N_3341);
and U4966 (N_4966,N_3548,N_2527);
nor U4967 (N_4967,N_2593,N_3664);
xnor U4968 (N_4968,N_2609,N_2478);
xnor U4969 (N_4969,N_2591,N_3428);
nand U4970 (N_4970,N_2727,N_2350);
nor U4971 (N_4971,N_3363,N_3731);
or U4972 (N_4972,N_2762,N_2043);
or U4973 (N_4973,N_2034,N_2014);
or U4974 (N_4974,N_3530,N_3623);
nand U4975 (N_4975,N_2905,N_2782);
or U4976 (N_4976,N_3500,N_3061);
nand U4977 (N_4977,N_2745,N_2716);
nor U4978 (N_4978,N_2757,N_3701);
nor U4979 (N_4979,N_3689,N_3397);
nor U4980 (N_4980,N_3033,N_2363);
and U4981 (N_4981,N_3506,N_2201);
nor U4982 (N_4982,N_3639,N_3908);
or U4983 (N_4983,N_3040,N_2581);
nor U4984 (N_4984,N_3059,N_3939);
or U4985 (N_4985,N_2574,N_3977);
nor U4986 (N_4986,N_3173,N_2559);
and U4987 (N_4987,N_3515,N_3624);
or U4988 (N_4988,N_2615,N_2944);
nand U4989 (N_4989,N_3416,N_3727);
and U4990 (N_4990,N_3350,N_2427);
or U4991 (N_4991,N_3135,N_2241);
nor U4992 (N_4992,N_2477,N_3822);
and U4993 (N_4993,N_2331,N_2502);
nand U4994 (N_4994,N_3857,N_3098);
nand U4995 (N_4995,N_3720,N_3650);
nor U4996 (N_4996,N_2323,N_3790);
or U4997 (N_4997,N_2997,N_3504);
nand U4998 (N_4998,N_3449,N_3279);
or U4999 (N_4999,N_2381,N_3369);
nand U5000 (N_5000,N_2642,N_3175);
nor U5001 (N_5001,N_2617,N_3879);
and U5002 (N_5002,N_2152,N_2412);
and U5003 (N_5003,N_3349,N_3454);
xnor U5004 (N_5004,N_2492,N_3289);
and U5005 (N_5005,N_3370,N_3992);
and U5006 (N_5006,N_2984,N_3715);
nand U5007 (N_5007,N_2303,N_3831);
nor U5008 (N_5008,N_2043,N_3854);
and U5009 (N_5009,N_3811,N_2738);
or U5010 (N_5010,N_3905,N_3279);
and U5011 (N_5011,N_3722,N_3918);
nand U5012 (N_5012,N_2991,N_3798);
xor U5013 (N_5013,N_3877,N_3180);
or U5014 (N_5014,N_3086,N_3393);
nand U5015 (N_5015,N_3661,N_3381);
xnor U5016 (N_5016,N_2178,N_3257);
and U5017 (N_5017,N_2302,N_3295);
or U5018 (N_5018,N_3109,N_2821);
or U5019 (N_5019,N_3019,N_3947);
or U5020 (N_5020,N_2715,N_2896);
nor U5021 (N_5021,N_3453,N_2033);
or U5022 (N_5022,N_2595,N_2331);
nand U5023 (N_5023,N_2108,N_2057);
nand U5024 (N_5024,N_2432,N_2743);
nand U5025 (N_5025,N_2266,N_3201);
xor U5026 (N_5026,N_3053,N_2429);
and U5027 (N_5027,N_3219,N_3421);
and U5028 (N_5028,N_3825,N_3947);
nor U5029 (N_5029,N_3954,N_2315);
or U5030 (N_5030,N_2129,N_2573);
and U5031 (N_5031,N_3040,N_3697);
nor U5032 (N_5032,N_2597,N_2546);
nor U5033 (N_5033,N_2364,N_2699);
nor U5034 (N_5034,N_3372,N_2160);
xnor U5035 (N_5035,N_3130,N_3936);
nand U5036 (N_5036,N_3052,N_2153);
or U5037 (N_5037,N_3833,N_2850);
and U5038 (N_5038,N_2429,N_2572);
or U5039 (N_5039,N_2586,N_2723);
and U5040 (N_5040,N_3815,N_2371);
and U5041 (N_5041,N_3163,N_3362);
nand U5042 (N_5042,N_3221,N_3722);
nor U5043 (N_5043,N_2909,N_3443);
xnor U5044 (N_5044,N_3322,N_3604);
nor U5045 (N_5045,N_3895,N_2607);
xnor U5046 (N_5046,N_3875,N_2187);
or U5047 (N_5047,N_3255,N_3351);
and U5048 (N_5048,N_2482,N_2632);
xnor U5049 (N_5049,N_3011,N_3169);
xnor U5050 (N_5050,N_3688,N_2481);
nand U5051 (N_5051,N_2455,N_2524);
xnor U5052 (N_5052,N_2649,N_3900);
or U5053 (N_5053,N_3162,N_3515);
nor U5054 (N_5054,N_3404,N_2401);
and U5055 (N_5055,N_2924,N_3595);
nor U5056 (N_5056,N_2611,N_2146);
and U5057 (N_5057,N_3026,N_3993);
and U5058 (N_5058,N_2760,N_3567);
or U5059 (N_5059,N_2127,N_3251);
nand U5060 (N_5060,N_3463,N_3980);
or U5061 (N_5061,N_2758,N_2825);
or U5062 (N_5062,N_3369,N_2437);
or U5063 (N_5063,N_2831,N_3907);
nand U5064 (N_5064,N_2291,N_2189);
or U5065 (N_5065,N_3699,N_2945);
nand U5066 (N_5066,N_3867,N_2667);
nand U5067 (N_5067,N_2531,N_2397);
and U5068 (N_5068,N_3990,N_2158);
nor U5069 (N_5069,N_3476,N_3059);
nand U5070 (N_5070,N_2079,N_2925);
and U5071 (N_5071,N_2191,N_2142);
nand U5072 (N_5072,N_3992,N_2288);
nor U5073 (N_5073,N_3263,N_2342);
nor U5074 (N_5074,N_3162,N_3003);
nand U5075 (N_5075,N_3315,N_3649);
nor U5076 (N_5076,N_3962,N_2019);
or U5077 (N_5077,N_2646,N_3218);
or U5078 (N_5078,N_3647,N_2339);
xor U5079 (N_5079,N_3376,N_3207);
nor U5080 (N_5080,N_3014,N_2867);
nor U5081 (N_5081,N_3334,N_2230);
nand U5082 (N_5082,N_3630,N_2441);
nand U5083 (N_5083,N_3730,N_3357);
nor U5084 (N_5084,N_3058,N_3572);
or U5085 (N_5085,N_3159,N_2365);
or U5086 (N_5086,N_2645,N_2339);
xor U5087 (N_5087,N_2682,N_3176);
nand U5088 (N_5088,N_2709,N_2460);
nor U5089 (N_5089,N_2039,N_3008);
nand U5090 (N_5090,N_3270,N_2011);
or U5091 (N_5091,N_3757,N_3977);
nand U5092 (N_5092,N_2696,N_3196);
and U5093 (N_5093,N_3312,N_2638);
nand U5094 (N_5094,N_2908,N_2324);
nand U5095 (N_5095,N_2076,N_2275);
nor U5096 (N_5096,N_3102,N_2295);
and U5097 (N_5097,N_3029,N_2599);
and U5098 (N_5098,N_3852,N_3832);
and U5099 (N_5099,N_3117,N_3302);
xor U5100 (N_5100,N_3336,N_2330);
xnor U5101 (N_5101,N_3791,N_2478);
xnor U5102 (N_5102,N_3640,N_3716);
or U5103 (N_5103,N_2790,N_2499);
xor U5104 (N_5104,N_2861,N_2712);
nor U5105 (N_5105,N_3993,N_2988);
and U5106 (N_5106,N_3166,N_3160);
or U5107 (N_5107,N_2127,N_2712);
and U5108 (N_5108,N_3041,N_2814);
and U5109 (N_5109,N_3126,N_2456);
or U5110 (N_5110,N_2359,N_2374);
and U5111 (N_5111,N_2188,N_3741);
xor U5112 (N_5112,N_2437,N_2007);
nor U5113 (N_5113,N_3230,N_3134);
nor U5114 (N_5114,N_3440,N_2231);
nand U5115 (N_5115,N_3768,N_2985);
and U5116 (N_5116,N_2767,N_3922);
nor U5117 (N_5117,N_2823,N_3861);
or U5118 (N_5118,N_3482,N_3076);
or U5119 (N_5119,N_3792,N_3312);
nand U5120 (N_5120,N_2699,N_2379);
and U5121 (N_5121,N_3792,N_3988);
nor U5122 (N_5122,N_2065,N_3425);
and U5123 (N_5123,N_2407,N_3784);
nor U5124 (N_5124,N_2234,N_3026);
nand U5125 (N_5125,N_3119,N_2705);
or U5126 (N_5126,N_2165,N_2394);
and U5127 (N_5127,N_2522,N_2082);
and U5128 (N_5128,N_3514,N_2050);
or U5129 (N_5129,N_2491,N_3257);
and U5130 (N_5130,N_3529,N_2278);
or U5131 (N_5131,N_3541,N_2930);
nand U5132 (N_5132,N_2359,N_3313);
nand U5133 (N_5133,N_2394,N_2405);
or U5134 (N_5134,N_3094,N_3421);
nor U5135 (N_5135,N_2501,N_3536);
or U5136 (N_5136,N_2334,N_3100);
and U5137 (N_5137,N_3390,N_2996);
nand U5138 (N_5138,N_3280,N_3104);
and U5139 (N_5139,N_3172,N_2128);
xor U5140 (N_5140,N_2341,N_3391);
xnor U5141 (N_5141,N_2012,N_3947);
xnor U5142 (N_5142,N_2566,N_2821);
and U5143 (N_5143,N_2076,N_3269);
nor U5144 (N_5144,N_3354,N_2239);
nand U5145 (N_5145,N_3002,N_3961);
nor U5146 (N_5146,N_3567,N_2442);
nor U5147 (N_5147,N_3773,N_2530);
and U5148 (N_5148,N_2685,N_2043);
or U5149 (N_5149,N_3862,N_3359);
or U5150 (N_5150,N_3765,N_3772);
and U5151 (N_5151,N_2962,N_3497);
nor U5152 (N_5152,N_2981,N_3843);
xnor U5153 (N_5153,N_2104,N_3668);
and U5154 (N_5154,N_3269,N_3366);
xor U5155 (N_5155,N_2526,N_3660);
xnor U5156 (N_5156,N_3106,N_3735);
or U5157 (N_5157,N_2372,N_2502);
nand U5158 (N_5158,N_2708,N_3929);
nand U5159 (N_5159,N_3814,N_2162);
or U5160 (N_5160,N_3597,N_3575);
and U5161 (N_5161,N_3080,N_3757);
nand U5162 (N_5162,N_3845,N_2893);
nand U5163 (N_5163,N_2978,N_2744);
and U5164 (N_5164,N_3367,N_3845);
or U5165 (N_5165,N_3374,N_2775);
or U5166 (N_5166,N_3915,N_3467);
nor U5167 (N_5167,N_3102,N_3600);
xor U5168 (N_5168,N_2478,N_3553);
and U5169 (N_5169,N_2306,N_2621);
nand U5170 (N_5170,N_2216,N_2142);
nor U5171 (N_5171,N_3466,N_3519);
and U5172 (N_5172,N_2905,N_3883);
or U5173 (N_5173,N_3892,N_2340);
or U5174 (N_5174,N_3004,N_2002);
and U5175 (N_5175,N_3671,N_2722);
or U5176 (N_5176,N_2663,N_3015);
and U5177 (N_5177,N_2532,N_2001);
and U5178 (N_5178,N_3127,N_3051);
nor U5179 (N_5179,N_2346,N_2440);
xor U5180 (N_5180,N_2302,N_2068);
nor U5181 (N_5181,N_2302,N_2297);
nor U5182 (N_5182,N_2192,N_2831);
nand U5183 (N_5183,N_3680,N_2878);
nand U5184 (N_5184,N_2732,N_3055);
or U5185 (N_5185,N_3522,N_2489);
or U5186 (N_5186,N_2839,N_3868);
nor U5187 (N_5187,N_3244,N_3280);
nand U5188 (N_5188,N_3949,N_3312);
nand U5189 (N_5189,N_3066,N_2646);
nand U5190 (N_5190,N_3928,N_2293);
nor U5191 (N_5191,N_3829,N_2120);
and U5192 (N_5192,N_3945,N_3430);
or U5193 (N_5193,N_2899,N_3275);
and U5194 (N_5194,N_3245,N_3455);
nand U5195 (N_5195,N_3074,N_3951);
and U5196 (N_5196,N_3787,N_3409);
and U5197 (N_5197,N_3547,N_3465);
or U5198 (N_5198,N_3372,N_3000);
xor U5199 (N_5199,N_3763,N_3051);
nand U5200 (N_5200,N_2788,N_3496);
nand U5201 (N_5201,N_2597,N_3897);
nand U5202 (N_5202,N_3865,N_2495);
nand U5203 (N_5203,N_3489,N_3427);
nor U5204 (N_5204,N_3304,N_3736);
or U5205 (N_5205,N_2487,N_3066);
nor U5206 (N_5206,N_2622,N_3882);
nand U5207 (N_5207,N_2302,N_3327);
nor U5208 (N_5208,N_3881,N_2138);
nor U5209 (N_5209,N_2839,N_2894);
xnor U5210 (N_5210,N_3294,N_3184);
nand U5211 (N_5211,N_2853,N_2054);
nand U5212 (N_5212,N_3131,N_2527);
nand U5213 (N_5213,N_3600,N_3722);
xor U5214 (N_5214,N_2561,N_3573);
nand U5215 (N_5215,N_2069,N_3885);
or U5216 (N_5216,N_2519,N_2342);
nor U5217 (N_5217,N_3718,N_2043);
xor U5218 (N_5218,N_3822,N_3667);
nor U5219 (N_5219,N_3825,N_2621);
and U5220 (N_5220,N_3433,N_2551);
nand U5221 (N_5221,N_3878,N_2172);
or U5222 (N_5222,N_2777,N_3946);
or U5223 (N_5223,N_2730,N_3312);
or U5224 (N_5224,N_3839,N_2103);
nor U5225 (N_5225,N_2403,N_2523);
or U5226 (N_5226,N_3642,N_3347);
nor U5227 (N_5227,N_2167,N_2935);
xor U5228 (N_5228,N_3750,N_3073);
nor U5229 (N_5229,N_3151,N_2277);
or U5230 (N_5230,N_2376,N_3017);
and U5231 (N_5231,N_2918,N_3878);
or U5232 (N_5232,N_3504,N_2847);
and U5233 (N_5233,N_2371,N_2550);
nand U5234 (N_5234,N_2609,N_2445);
or U5235 (N_5235,N_2556,N_2187);
nor U5236 (N_5236,N_3587,N_2310);
and U5237 (N_5237,N_2012,N_2311);
nor U5238 (N_5238,N_2799,N_2904);
nand U5239 (N_5239,N_3552,N_3367);
nor U5240 (N_5240,N_3276,N_3418);
and U5241 (N_5241,N_2523,N_3446);
xor U5242 (N_5242,N_2113,N_3258);
or U5243 (N_5243,N_3287,N_2528);
nor U5244 (N_5244,N_3768,N_3236);
or U5245 (N_5245,N_3861,N_2479);
and U5246 (N_5246,N_3415,N_3042);
nor U5247 (N_5247,N_3821,N_2054);
xnor U5248 (N_5248,N_3988,N_2173);
nand U5249 (N_5249,N_3672,N_2352);
nor U5250 (N_5250,N_3850,N_2156);
or U5251 (N_5251,N_2968,N_3568);
xor U5252 (N_5252,N_2110,N_3050);
nand U5253 (N_5253,N_3800,N_2422);
or U5254 (N_5254,N_2860,N_2372);
nand U5255 (N_5255,N_2847,N_2113);
and U5256 (N_5256,N_2352,N_2538);
or U5257 (N_5257,N_3556,N_2161);
nor U5258 (N_5258,N_3570,N_2639);
nor U5259 (N_5259,N_3319,N_2743);
nand U5260 (N_5260,N_3197,N_2411);
and U5261 (N_5261,N_2562,N_2795);
nor U5262 (N_5262,N_3247,N_2071);
or U5263 (N_5263,N_3656,N_3716);
nand U5264 (N_5264,N_2688,N_2019);
and U5265 (N_5265,N_2709,N_2925);
and U5266 (N_5266,N_2848,N_3991);
nand U5267 (N_5267,N_2340,N_2254);
nor U5268 (N_5268,N_2752,N_2508);
xnor U5269 (N_5269,N_3759,N_2737);
or U5270 (N_5270,N_2276,N_2280);
and U5271 (N_5271,N_3116,N_3615);
and U5272 (N_5272,N_2809,N_3164);
nand U5273 (N_5273,N_3719,N_3333);
nor U5274 (N_5274,N_3277,N_3329);
and U5275 (N_5275,N_2550,N_3374);
and U5276 (N_5276,N_2621,N_3432);
and U5277 (N_5277,N_2675,N_2971);
or U5278 (N_5278,N_3846,N_3763);
nor U5279 (N_5279,N_2986,N_3029);
and U5280 (N_5280,N_3358,N_3652);
nor U5281 (N_5281,N_2596,N_2878);
xor U5282 (N_5282,N_3099,N_3487);
nor U5283 (N_5283,N_3110,N_2411);
nand U5284 (N_5284,N_3194,N_3670);
or U5285 (N_5285,N_2307,N_3571);
nor U5286 (N_5286,N_2503,N_3486);
and U5287 (N_5287,N_3760,N_3571);
and U5288 (N_5288,N_3060,N_3557);
nor U5289 (N_5289,N_2525,N_3838);
nand U5290 (N_5290,N_3795,N_2125);
nand U5291 (N_5291,N_2677,N_3895);
or U5292 (N_5292,N_3326,N_2375);
or U5293 (N_5293,N_3243,N_3751);
nand U5294 (N_5294,N_2482,N_3999);
or U5295 (N_5295,N_3352,N_3214);
and U5296 (N_5296,N_2055,N_3403);
nor U5297 (N_5297,N_3153,N_3756);
nor U5298 (N_5298,N_3056,N_3444);
and U5299 (N_5299,N_3546,N_2924);
nand U5300 (N_5300,N_2589,N_3284);
nand U5301 (N_5301,N_3426,N_2197);
or U5302 (N_5302,N_3182,N_2396);
nand U5303 (N_5303,N_2144,N_3531);
nor U5304 (N_5304,N_3912,N_3450);
nor U5305 (N_5305,N_3700,N_3235);
nand U5306 (N_5306,N_2615,N_2313);
nand U5307 (N_5307,N_3117,N_3940);
nor U5308 (N_5308,N_3388,N_3545);
nand U5309 (N_5309,N_3946,N_3208);
xor U5310 (N_5310,N_2114,N_3922);
nor U5311 (N_5311,N_3610,N_2188);
nand U5312 (N_5312,N_3421,N_2142);
xnor U5313 (N_5313,N_3287,N_2885);
nor U5314 (N_5314,N_3112,N_2254);
or U5315 (N_5315,N_3586,N_2824);
and U5316 (N_5316,N_3144,N_2521);
nand U5317 (N_5317,N_3014,N_2071);
or U5318 (N_5318,N_3881,N_2605);
and U5319 (N_5319,N_2006,N_2600);
nor U5320 (N_5320,N_2120,N_3019);
nor U5321 (N_5321,N_3133,N_2708);
and U5322 (N_5322,N_3154,N_2822);
nor U5323 (N_5323,N_3168,N_2227);
xnor U5324 (N_5324,N_2757,N_2356);
xnor U5325 (N_5325,N_3829,N_3655);
xor U5326 (N_5326,N_2511,N_2393);
or U5327 (N_5327,N_2960,N_3906);
nor U5328 (N_5328,N_2176,N_3244);
nand U5329 (N_5329,N_2505,N_3016);
nand U5330 (N_5330,N_2416,N_2370);
and U5331 (N_5331,N_3921,N_3196);
and U5332 (N_5332,N_2970,N_3501);
and U5333 (N_5333,N_3396,N_2047);
or U5334 (N_5334,N_2392,N_2875);
nand U5335 (N_5335,N_3621,N_2786);
or U5336 (N_5336,N_2312,N_2251);
or U5337 (N_5337,N_2053,N_3448);
and U5338 (N_5338,N_3652,N_3030);
and U5339 (N_5339,N_3628,N_2441);
xnor U5340 (N_5340,N_3096,N_3905);
nand U5341 (N_5341,N_2739,N_3538);
and U5342 (N_5342,N_3600,N_2075);
nor U5343 (N_5343,N_3070,N_3962);
or U5344 (N_5344,N_2220,N_3120);
and U5345 (N_5345,N_3509,N_2422);
nor U5346 (N_5346,N_3965,N_3341);
nor U5347 (N_5347,N_2787,N_2598);
nand U5348 (N_5348,N_3800,N_2128);
xnor U5349 (N_5349,N_2434,N_2964);
and U5350 (N_5350,N_2622,N_3382);
nor U5351 (N_5351,N_3582,N_2443);
or U5352 (N_5352,N_3722,N_3964);
nor U5353 (N_5353,N_2995,N_3341);
or U5354 (N_5354,N_2387,N_2185);
nand U5355 (N_5355,N_2472,N_3543);
or U5356 (N_5356,N_3403,N_2234);
and U5357 (N_5357,N_3628,N_3057);
nor U5358 (N_5358,N_3109,N_3997);
nor U5359 (N_5359,N_3140,N_3351);
nand U5360 (N_5360,N_2333,N_3697);
or U5361 (N_5361,N_2580,N_2114);
xnor U5362 (N_5362,N_2169,N_2503);
and U5363 (N_5363,N_2404,N_2913);
nand U5364 (N_5364,N_3088,N_2989);
nand U5365 (N_5365,N_2888,N_3214);
nor U5366 (N_5366,N_3764,N_3427);
or U5367 (N_5367,N_2233,N_3831);
or U5368 (N_5368,N_3333,N_2117);
or U5369 (N_5369,N_3975,N_2648);
nand U5370 (N_5370,N_2545,N_3543);
or U5371 (N_5371,N_2699,N_2215);
nand U5372 (N_5372,N_3802,N_2243);
xor U5373 (N_5373,N_2400,N_2875);
nor U5374 (N_5374,N_2384,N_3826);
nand U5375 (N_5375,N_2230,N_2723);
and U5376 (N_5376,N_3017,N_3752);
and U5377 (N_5377,N_3383,N_3610);
nor U5378 (N_5378,N_3470,N_2218);
or U5379 (N_5379,N_2866,N_2363);
or U5380 (N_5380,N_3760,N_2552);
nand U5381 (N_5381,N_3889,N_2820);
and U5382 (N_5382,N_3558,N_2722);
nor U5383 (N_5383,N_2031,N_2593);
nor U5384 (N_5384,N_2995,N_2329);
nand U5385 (N_5385,N_2323,N_2469);
xor U5386 (N_5386,N_2618,N_2843);
nand U5387 (N_5387,N_2735,N_3758);
or U5388 (N_5388,N_3339,N_3698);
nand U5389 (N_5389,N_2419,N_2695);
or U5390 (N_5390,N_3708,N_2040);
and U5391 (N_5391,N_3638,N_2602);
nor U5392 (N_5392,N_3115,N_3554);
nand U5393 (N_5393,N_3805,N_2890);
or U5394 (N_5394,N_2678,N_2097);
and U5395 (N_5395,N_2848,N_3921);
nand U5396 (N_5396,N_2891,N_3649);
and U5397 (N_5397,N_2949,N_2154);
and U5398 (N_5398,N_3337,N_2470);
nor U5399 (N_5399,N_2159,N_2886);
and U5400 (N_5400,N_2730,N_3873);
xor U5401 (N_5401,N_3390,N_3163);
and U5402 (N_5402,N_2950,N_2403);
and U5403 (N_5403,N_2820,N_3202);
nor U5404 (N_5404,N_2757,N_3344);
or U5405 (N_5405,N_2466,N_2923);
and U5406 (N_5406,N_2965,N_3933);
xnor U5407 (N_5407,N_3116,N_2420);
nand U5408 (N_5408,N_3834,N_3320);
nand U5409 (N_5409,N_3604,N_2636);
or U5410 (N_5410,N_3272,N_2299);
and U5411 (N_5411,N_2019,N_2687);
or U5412 (N_5412,N_2924,N_3663);
and U5413 (N_5413,N_2423,N_3492);
nor U5414 (N_5414,N_3160,N_3890);
nand U5415 (N_5415,N_3498,N_3612);
nand U5416 (N_5416,N_2123,N_3601);
or U5417 (N_5417,N_2884,N_2412);
nor U5418 (N_5418,N_3498,N_3122);
nor U5419 (N_5419,N_2967,N_2101);
nand U5420 (N_5420,N_2403,N_2429);
and U5421 (N_5421,N_2291,N_2848);
and U5422 (N_5422,N_2274,N_3805);
nand U5423 (N_5423,N_2128,N_3970);
nand U5424 (N_5424,N_2256,N_3984);
or U5425 (N_5425,N_3590,N_3683);
and U5426 (N_5426,N_2489,N_2141);
and U5427 (N_5427,N_3901,N_2725);
and U5428 (N_5428,N_3688,N_2012);
or U5429 (N_5429,N_2325,N_3747);
nor U5430 (N_5430,N_3130,N_3526);
nor U5431 (N_5431,N_3381,N_3413);
or U5432 (N_5432,N_2572,N_3817);
or U5433 (N_5433,N_2955,N_3461);
nor U5434 (N_5434,N_2323,N_3340);
nor U5435 (N_5435,N_3356,N_3418);
or U5436 (N_5436,N_2317,N_2907);
or U5437 (N_5437,N_3759,N_3803);
nand U5438 (N_5438,N_3586,N_3298);
xor U5439 (N_5439,N_2232,N_3393);
or U5440 (N_5440,N_3587,N_3876);
or U5441 (N_5441,N_2506,N_3980);
nand U5442 (N_5442,N_2637,N_3637);
and U5443 (N_5443,N_2849,N_2103);
xor U5444 (N_5444,N_3213,N_3698);
nand U5445 (N_5445,N_3790,N_3322);
nor U5446 (N_5446,N_2861,N_3379);
nand U5447 (N_5447,N_2612,N_2970);
nor U5448 (N_5448,N_3537,N_2918);
nand U5449 (N_5449,N_3261,N_2918);
nand U5450 (N_5450,N_3499,N_2941);
nand U5451 (N_5451,N_3841,N_2817);
and U5452 (N_5452,N_2586,N_2169);
nand U5453 (N_5453,N_2188,N_3488);
or U5454 (N_5454,N_3264,N_2356);
nand U5455 (N_5455,N_2385,N_2032);
and U5456 (N_5456,N_3427,N_2172);
nor U5457 (N_5457,N_2775,N_3879);
and U5458 (N_5458,N_3105,N_2933);
nand U5459 (N_5459,N_3715,N_2436);
and U5460 (N_5460,N_2391,N_3857);
or U5461 (N_5461,N_3538,N_2134);
nor U5462 (N_5462,N_2579,N_3139);
nor U5463 (N_5463,N_3582,N_3912);
xnor U5464 (N_5464,N_3049,N_3201);
nor U5465 (N_5465,N_2627,N_2382);
and U5466 (N_5466,N_3537,N_3746);
and U5467 (N_5467,N_2919,N_2728);
or U5468 (N_5468,N_2312,N_3584);
nand U5469 (N_5469,N_3804,N_3038);
nor U5470 (N_5470,N_3623,N_2459);
nor U5471 (N_5471,N_3211,N_3145);
nand U5472 (N_5472,N_2777,N_2376);
and U5473 (N_5473,N_3862,N_3987);
and U5474 (N_5474,N_3844,N_2909);
xor U5475 (N_5475,N_3293,N_3977);
and U5476 (N_5476,N_3677,N_3624);
nor U5477 (N_5477,N_3651,N_2876);
or U5478 (N_5478,N_2779,N_3310);
nor U5479 (N_5479,N_3585,N_3162);
nand U5480 (N_5480,N_3232,N_2871);
or U5481 (N_5481,N_3698,N_3082);
or U5482 (N_5482,N_3147,N_3742);
nor U5483 (N_5483,N_3064,N_2712);
nor U5484 (N_5484,N_3100,N_2330);
nand U5485 (N_5485,N_3388,N_3558);
nor U5486 (N_5486,N_3949,N_2144);
nor U5487 (N_5487,N_3997,N_3691);
or U5488 (N_5488,N_2005,N_2246);
nor U5489 (N_5489,N_3876,N_3147);
and U5490 (N_5490,N_2507,N_2255);
or U5491 (N_5491,N_2785,N_2760);
or U5492 (N_5492,N_2175,N_2333);
nand U5493 (N_5493,N_2344,N_2457);
nand U5494 (N_5494,N_3583,N_3761);
or U5495 (N_5495,N_3325,N_2002);
nand U5496 (N_5496,N_2412,N_2960);
and U5497 (N_5497,N_2527,N_3865);
or U5498 (N_5498,N_3758,N_2487);
xor U5499 (N_5499,N_2961,N_2862);
and U5500 (N_5500,N_2076,N_3771);
nor U5501 (N_5501,N_3049,N_3084);
and U5502 (N_5502,N_3693,N_2133);
and U5503 (N_5503,N_2129,N_3409);
and U5504 (N_5504,N_2529,N_2292);
and U5505 (N_5505,N_3030,N_3995);
nor U5506 (N_5506,N_2723,N_3109);
or U5507 (N_5507,N_3507,N_3841);
nand U5508 (N_5508,N_2902,N_2427);
nor U5509 (N_5509,N_3319,N_3672);
nand U5510 (N_5510,N_2165,N_3664);
or U5511 (N_5511,N_2286,N_2076);
and U5512 (N_5512,N_3577,N_3094);
or U5513 (N_5513,N_3628,N_3511);
nand U5514 (N_5514,N_2765,N_3709);
nand U5515 (N_5515,N_2382,N_3536);
nand U5516 (N_5516,N_2065,N_2444);
and U5517 (N_5517,N_2979,N_3854);
nand U5518 (N_5518,N_2059,N_3719);
nor U5519 (N_5519,N_2130,N_3568);
or U5520 (N_5520,N_2360,N_2608);
nand U5521 (N_5521,N_3422,N_2598);
or U5522 (N_5522,N_3808,N_3684);
or U5523 (N_5523,N_3323,N_2757);
nor U5524 (N_5524,N_3028,N_3994);
or U5525 (N_5525,N_2716,N_2185);
and U5526 (N_5526,N_2797,N_3843);
and U5527 (N_5527,N_2507,N_2031);
and U5528 (N_5528,N_3965,N_2554);
xnor U5529 (N_5529,N_2236,N_3406);
nand U5530 (N_5530,N_2714,N_2176);
or U5531 (N_5531,N_3844,N_2581);
or U5532 (N_5532,N_2823,N_3715);
or U5533 (N_5533,N_2080,N_2641);
or U5534 (N_5534,N_2501,N_3740);
xor U5535 (N_5535,N_2801,N_2118);
nand U5536 (N_5536,N_3987,N_2793);
xnor U5537 (N_5537,N_3366,N_3011);
or U5538 (N_5538,N_3426,N_3247);
or U5539 (N_5539,N_3456,N_3017);
and U5540 (N_5540,N_3928,N_2047);
nand U5541 (N_5541,N_2841,N_2501);
xor U5542 (N_5542,N_2806,N_3417);
nor U5543 (N_5543,N_3722,N_3330);
nor U5544 (N_5544,N_2124,N_2289);
and U5545 (N_5545,N_2292,N_3119);
nor U5546 (N_5546,N_2001,N_2161);
nand U5547 (N_5547,N_2589,N_3144);
or U5548 (N_5548,N_3313,N_3874);
or U5549 (N_5549,N_3862,N_3062);
and U5550 (N_5550,N_2514,N_3313);
nand U5551 (N_5551,N_3383,N_2271);
and U5552 (N_5552,N_2823,N_2621);
and U5553 (N_5553,N_2535,N_2929);
nor U5554 (N_5554,N_2669,N_2063);
or U5555 (N_5555,N_3943,N_2122);
and U5556 (N_5556,N_3087,N_3194);
nor U5557 (N_5557,N_3982,N_3166);
or U5558 (N_5558,N_2462,N_2224);
nand U5559 (N_5559,N_2560,N_2069);
xor U5560 (N_5560,N_3255,N_2306);
or U5561 (N_5561,N_3842,N_2203);
xor U5562 (N_5562,N_2941,N_2554);
nand U5563 (N_5563,N_2751,N_3561);
nor U5564 (N_5564,N_3695,N_2693);
and U5565 (N_5565,N_3534,N_3926);
or U5566 (N_5566,N_2919,N_3391);
nand U5567 (N_5567,N_3951,N_2709);
and U5568 (N_5568,N_3229,N_3795);
nor U5569 (N_5569,N_3345,N_2761);
nand U5570 (N_5570,N_2437,N_2250);
or U5571 (N_5571,N_2579,N_2541);
xnor U5572 (N_5572,N_2330,N_3740);
nor U5573 (N_5573,N_3814,N_2797);
nor U5574 (N_5574,N_3459,N_2239);
nand U5575 (N_5575,N_3120,N_3113);
or U5576 (N_5576,N_2881,N_3336);
nand U5577 (N_5577,N_2921,N_3330);
nand U5578 (N_5578,N_3773,N_3957);
nor U5579 (N_5579,N_3271,N_2921);
and U5580 (N_5580,N_3056,N_2011);
nor U5581 (N_5581,N_3112,N_2368);
xor U5582 (N_5582,N_2516,N_2456);
and U5583 (N_5583,N_2894,N_2258);
xor U5584 (N_5584,N_3666,N_2356);
or U5585 (N_5585,N_2716,N_2020);
and U5586 (N_5586,N_2888,N_3367);
nand U5587 (N_5587,N_3705,N_3212);
nor U5588 (N_5588,N_2383,N_2454);
nand U5589 (N_5589,N_3499,N_3541);
nor U5590 (N_5590,N_2119,N_2743);
nand U5591 (N_5591,N_2181,N_3586);
nand U5592 (N_5592,N_3392,N_3610);
or U5593 (N_5593,N_2767,N_2948);
and U5594 (N_5594,N_3455,N_2116);
or U5595 (N_5595,N_3372,N_3003);
nor U5596 (N_5596,N_3574,N_3391);
nor U5597 (N_5597,N_3832,N_2993);
or U5598 (N_5598,N_2919,N_3432);
nand U5599 (N_5599,N_3535,N_2513);
and U5600 (N_5600,N_2515,N_3568);
or U5601 (N_5601,N_3911,N_3883);
nor U5602 (N_5602,N_3369,N_3307);
or U5603 (N_5603,N_3343,N_2638);
nand U5604 (N_5604,N_3102,N_3046);
nor U5605 (N_5605,N_2442,N_2211);
nor U5606 (N_5606,N_3583,N_2614);
nand U5607 (N_5607,N_3219,N_3217);
or U5608 (N_5608,N_2982,N_2422);
or U5609 (N_5609,N_3970,N_3686);
or U5610 (N_5610,N_3917,N_3102);
nand U5611 (N_5611,N_2734,N_3885);
xnor U5612 (N_5612,N_3718,N_3021);
nor U5613 (N_5613,N_3546,N_2587);
and U5614 (N_5614,N_2750,N_3323);
and U5615 (N_5615,N_2589,N_2086);
nand U5616 (N_5616,N_3481,N_2853);
nand U5617 (N_5617,N_3323,N_2812);
or U5618 (N_5618,N_2076,N_2333);
or U5619 (N_5619,N_2875,N_3271);
nor U5620 (N_5620,N_3709,N_2777);
or U5621 (N_5621,N_3659,N_2289);
and U5622 (N_5622,N_3257,N_2764);
nand U5623 (N_5623,N_3802,N_3443);
and U5624 (N_5624,N_2341,N_3151);
or U5625 (N_5625,N_3122,N_2332);
xor U5626 (N_5626,N_3012,N_3630);
nor U5627 (N_5627,N_3154,N_2842);
or U5628 (N_5628,N_2239,N_3454);
nor U5629 (N_5629,N_2649,N_3363);
and U5630 (N_5630,N_3645,N_3491);
and U5631 (N_5631,N_3511,N_3142);
or U5632 (N_5632,N_3165,N_2266);
and U5633 (N_5633,N_3181,N_3332);
nand U5634 (N_5634,N_2247,N_2500);
nand U5635 (N_5635,N_2925,N_3446);
or U5636 (N_5636,N_3796,N_3928);
and U5637 (N_5637,N_2626,N_3017);
and U5638 (N_5638,N_3143,N_3806);
nor U5639 (N_5639,N_3035,N_2576);
nand U5640 (N_5640,N_2353,N_3629);
nand U5641 (N_5641,N_3198,N_2386);
nand U5642 (N_5642,N_3830,N_2355);
and U5643 (N_5643,N_2062,N_3882);
nand U5644 (N_5644,N_3062,N_3752);
and U5645 (N_5645,N_3132,N_3928);
or U5646 (N_5646,N_3473,N_2814);
or U5647 (N_5647,N_2428,N_3363);
nand U5648 (N_5648,N_2419,N_3210);
nand U5649 (N_5649,N_3607,N_2648);
nand U5650 (N_5650,N_3358,N_3127);
or U5651 (N_5651,N_2307,N_2260);
nand U5652 (N_5652,N_3763,N_2109);
nand U5653 (N_5653,N_2625,N_3395);
xnor U5654 (N_5654,N_2567,N_2764);
nand U5655 (N_5655,N_3346,N_3924);
or U5656 (N_5656,N_2005,N_2806);
nor U5657 (N_5657,N_2730,N_2439);
nand U5658 (N_5658,N_3125,N_2450);
or U5659 (N_5659,N_3475,N_3341);
or U5660 (N_5660,N_2727,N_3904);
nand U5661 (N_5661,N_3178,N_3170);
nor U5662 (N_5662,N_3097,N_3365);
nor U5663 (N_5663,N_3766,N_3289);
nor U5664 (N_5664,N_2292,N_3230);
nand U5665 (N_5665,N_2418,N_3049);
and U5666 (N_5666,N_3652,N_2785);
nor U5667 (N_5667,N_3565,N_2128);
nor U5668 (N_5668,N_2339,N_2817);
or U5669 (N_5669,N_2428,N_3129);
xor U5670 (N_5670,N_2175,N_3074);
nor U5671 (N_5671,N_2002,N_2263);
or U5672 (N_5672,N_3517,N_3804);
or U5673 (N_5673,N_2153,N_2038);
xnor U5674 (N_5674,N_3572,N_3186);
or U5675 (N_5675,N_3330,N_3402);
xnor U5676 (N_5676,N_3533,N_2395);
xnor U5677 (N_5677,N_3387,N_2681);
nor U5678 (N_5678,N_3851,N_2120);
nand U5679 (N_5679,N_3054,N_3302);
nor U5680 (N_5680,N_2873,N_2172);
or U5681 (N_5681,N_3973,N_3443);
xnor U5682 (N_5682,N_2703,N_2815);
nand U5683 (N_5683,N_3843,N_3832);
nand U5684 (N_5684,N_2706,N_2934);
nand U5685 (N_5685,N_2644,N_3419);
nand U5686 (N_5686,N_3648,N_3634);
nand U5687 (N_5687,N_3431,N_2279);
and U5688 (N_5688,N_3131,N_3327);
or U5689 (N_5689,N_2858,N_3332);
and U5690 (N_5690,N_3192,N_2803);
nor U5691 (N_5691,N_2173,N_3762);
nor U5692 (N_5692,N_2963,N_3919);
and U5693 (N_5693,N_3239,N_2651);
nor U5694 (N_5694,N_3820,N_3680);
nor U5695 (N_5695,N_3825,N_3289);
or U5696 (N_5696,N_3773,N_3977);
nand U5697 (N_5697,N_2198,N_3837);
xnor U5698 (N_5698,N_3413,N_2746);
or U5699 (N_5699,N_2337,N_3954);
xnor U5700 (N_5700,N_3027,N_3384);
and U5701 (N_5701,N_3170,N_3519);
nand U5702 (N_5702,N_2517,N_3193);
nor U5703 (N_5703,N_2636,N_2523);
or U5704 (N_5704,N_2104,N_3461);
or U5705 (N_5705,N_2178,N_2520);
or U5706 (N_5706,N_3269,N_3805);
or U5707 (N_5707,N_2636,N_3705);
nor U5708 (N_5708,N_2272,N_3576);
nor U5709 (N_5709,N_3477,N_2139);
nand U5710 (N_5710,N_2592,N_3004);
nor U5711 (N_5711,N_3290,N_2753);
nand U5712 (N_5712,N_2814,N_3281);
and U5713 (N_5713,N_3628,N_3936);
nand U5714 (N_5714,N_3743,N_3723);
xnor U5715 (N_5715,N_3875,N_3793);
nand U5716 (N_5716,N_3452,N_2112);
nor U5717 (N_5717,N_2589,N_2327);
xnor U5718 (N_5718,N_3904,N_2448);
xnor U5719 (N_5719,N_3125,N_3894);
xor U5720 (N_5720,N_3662,N_3344);
nand U5721 (N_5721,N_2714,N_2530);
nand U5722 (N_5722,N_3156,N_3545);
or U5723 (N_5723,N_2615,N_3847);
and U5724 (N_5724,N_2861,N_2100);
nor U5725 (N_5725,N_3884,N_2684);
or U5726 (N_5726,N_3880,N_2573);
nor U5727 (N_5727,N_2446,N_3462);
and U5728 (N_5728,N_3081,N_3942);
or U5729 (N_5729,N_3698,N_3767);
and U5730 (N_5730,N_3426,N_3604);
nor U5731 (N_5731,N_3434,N_2524);
nor U5732 (N_5732,N_3427,N_2948);
xor U5733 (N_5733,N_2015,N_2191);
or U5734 (N_5734,N_2759,N_3744);
nor U5735 (N_5735,N_3214,N_3907);
and U5736 (N_5736,N_3944,N_2617);
nand U5737 (N_5737,N_2762,N_3352);
and U5738 (N_5738,N_3952,N_3903);
nand U5739 (N_5739,N_2047,N_3997);
and U5740 (N_5740,N_3301,N_2699);
nand U5741 (N_5741,N_3921,N_3675);
or U5742 (N_5742,N_2403,N_3651);
nand U5743 (N_5743,N_3852,N_2802);
nand U5744 (N_5744,N_2233,N_3789);
and U5745 (N_5745,N_2790,N_3141);
and U5746 (N_5746,N_3819,N_3912);
nor U5747 (N_5747,N_2327,N_3860);
and U5748 (N_5748,N_2650,N_3819);
nor U5749 (N_5749,N_3743,N_3396);
nand U5750 (N_5750,N_3280,N_2367);
and U5751 (N_5751,N_3646,N_2902);
or U5752 (N_5752,N_3697,N_3547);
nand U5753 (N_5753,N_3065,N_2246);
nand U5754 (N_5754,N_2135,N_3709);
nand U5755 (N_5755,N_2153,N_2742);
or U5756 (N_5756,N_2117,N_3100);
or U5757 (N_5757,N_2141,N_2171);
nor U5758 (N_5758,N_2472,N_3323);
nand U5759 (N_5759,N_3430,N_2797);
and U5760 (N_5760,N_2577,N_3019);
nor U5761 (N_5761,N_2462,N_2906);
and U5762 (N_5762,N_2925,N_3682);
and U5763 (N_5763,N_3313,N_2672);
nand U5764 (N_5764,N_2534,N_2739);
and U5765 (N_5765,N_2142,N_2407);
nor U5766 (N_5766,N_3168,N_3421);
nor U5767 (N_5767,N_3120,N_2908);
or U5768 (N_5768,N_3731,N_2226);
and U5769 (N_5769,N_2045,N_3432);
xnor U5770 (N_5770,N_2045,N_2860);
nor U5771 (N_5771,N_3290,N_2527);
or U5772 (N_5772,N_3773,N_3691);
or U5773 (N_5773,N_2917,N_3788);
and U5774 (N_5774,N_2839,N_2814);
nor U5775 (N_5775,N_2760,N_3829);
or U5776 (N_5776,N_3692,N_2420);
or U5777 (N_5777,N_2106,N_3583);
nor U5778 (N_5778,N_3588,N_3501);
and U5779 (N_5779,N_2915,N_3763);
nand U5780 (N_5780,N_3779,N_2942);
nand U5781 (N_5781,N_2543,N_2565);
and U5782 (N_5782,N_3834,N_2605);
nor U5783 (N_5783,N_3684,N_3200);
or U5784 (N_5784,N_3366,N_3564);
nand U5785 (N_5785,N_3890,N_3046);
nand U5786 (N_5786,N_2315,N_2846);
nor U5787 (N_5787,N_3704,N_2900);
nor U5788 (N_5788,N_2029,N_3504);
or U5789 (N_5789,N_3685,N_3540);
and U5790 (N_5790,N_3819,N_2981);
or U5791 (N_5791,N_3303,N_2366);
xnor U5792 (N_5792,N_3778,N_3936);
nand U5793 (N_5793,N_2894,N_2049);
or U5794 (N_5794,N_2954,N_2283);
or U5795 (N_5795,N_3962,N_2894);
and U5796 (N_5796,N_3957,N_2912);
and U5797 (N_5797,N_2269,N_3353);
or U5798 (N_5798,N_2173,N_2632);
nor U5799 (N_5799,N_2689,N_2882);
and U5800 (N_5800,N_3746,N_2688);
or U5801 (N_5801,N_3951,N_3527);
xor U5802 (N_5802,N_2737,N_2266);
and U5803 (N_5803,N_3462,N_3492);
xor U5804 (N_5804,N_2645,N_3696);
xnor U5805 (N_5805,N_3212,N_3308);
nor U5806 (N_5806,N_3988,N_2118);
nand U5807 (N_5807,N_3909,N_3768);
nor U5808 (N_5808,N_3341,N_3950);
or U5809 (N_5809,N_2219,N_3540);
nor U5810 (N_5810,N_3446,N_2550);
or U5811 (N_5811,N_2449,N_3704);
xnor U5812 (N_5812,N_2713,N_3467);
or U5813 (N_5813,N_2945,N_2971);
xnor U5814 (N_5814,N_3654,N_2929);
nor U5815 (N_5815,N_3773,N_2360);
nand U5816 (N_5816,N_3632,N_2261);
and U5817 (N_5817,N_2084,N_3048);
nor U5818 (N_5818,N_3841,N_3667);
or U5819 (N_5819,N_3668,N_2080);
or U5820 (N_5820,N_2850,N_2555);
and U5821 (N_5821,N_2417,N_2312);
or U5822 (N_5822,N_2443,N_3598);
nor U5823 (N_5823,N_3127,N_3132);
nor U5824 (N_5824,N_3492,N_3990);
or U5825 (N_5825,N_2900,N_2437);
or U5826 (N_5826,N_3254,N_2919);
nor U5827 (N_5827,N_3252,N_3672);
xor U5828 (N_5828,N_2634,N_2880);
nand U5829 (N_5829,N_3128,N_3396);
nand U5830 (N_5830,N_2558,N_2554);
nor U5831 (N_5831,N_3018,N_3110);
xor U5832 (N_5832,N_2207,N_2288);
nor U5833 (N_5833,N_3304,N_2688);
and U5834 (N_5834,N_2932,N_3717);
xor U5835 (N_5835,N_2732,N_2117);
nand U5836 (N_5836,N_2703,N_3054);
nand U5837 (N_5837,N_2592,N_2668);
nor U5838 (N_5838,N_3859,N_2070);
or U5839 (N_5839,N_3029,N_2407);
or U5840 (N_5840,N_3886,N_2366);
nor U5841 (N_5841,N_2576,N_2622);
and U5842 (N_5842,N_2906,N_2089);
and U5843 (N_5843,N_3274,N_3622);
and U5844 (N_5844,N_2551,N_3388);
nor U5845 (N_5845,N_3575,N_3195);
or U5846 (N_5846,N_3463,N_2223);
or U5847 (N_5847,N_3119,N_2378);
or U5848 (N_5848,N_3695,N_3342);
xnor U5849 (N_5849,N_2738,N_2373);
nand U5850 (N_5850,N_2169,N_2132);
nand U5851 (N_5851,N_3381,N_3625);
nand U5852 (N_5852,N_2183,N_2694);
nand U5853 (N_5853,N_2939,N_2647);
and U5854 (N_5854,N_3640,N_2733);
and U5855 (N_5855,N_3436,N_3874);
or U5856 (N_5856,N_3326,N_2734);
and U5857 (N_5857,N_3173,N_3993);
nor U5858 (N_5858,N_2011,N_2097);
xnor U5859 (N_5859,N_2680,N_3223);
nor U5860 (N_5860,N_3950,N_2689);
and U5861 (N_5861,N_3800,N_2840);
nand U5862 (N_5862,N_2698,N_2873);
nand U5863 (N_5863,N_2985,N_2086);
nand U5864 (N_5864,N_3500,N_2030);
and U5865 (N_5865,N_2922,N_3350);
nor U5866 (N_5866,N_2660,N_3250);
and U5867 (N_5867,N_3982,N_3869);
and U5868 (N_5868,N_3573,N_3821);
or U5869 (N_5869,N_2331,N_3534);
and U5870 (N_5870,N_3736,N_2581);
xor U5871 (N_5871,N_2820,N_2116);
xnor U5872 (N_5872,N_2748,N_2765);
nor U5873 (N_5873,N_2573,N_2319);
or U5874 (N_5874,N_3047,N_2753);
or U5875 (N_5875,N_3518,N_2851);
or U5876 (N_5876,N_2553,N_2744);
nand U5877 (N_5877,N_2824,N_3447);
nand U5878 (N_5878,N_2027,N_2186);
nor U5879 (N_5879,N_2712,N_2407);
nand U5880 (N_5880,N_3569,N_3239);
nand U5881 (N_5881,N_3903,N_3495);
or U5882 (N_5882,N_2853,N_2813);
and U5883 (N_5883,N_2901,N_2448);
nor U5884 (N_5884,N_3915,N_2686);
and U5885 (N_5885,N_2528,N_2275);
nand U5886 (N_5886,N_2584,N_3671);
nor U5887 (N_5887,N_3412,N_3468);
nor U5888 (N_5888,N_3667,N_3844);
and U5889 (N_5889,N_2393,N_2020);
nor U5890 (N_5890,N_2964,N_3863);
and U5891 (N_5891,N_2862,N_3659);
nor U5892 (N_5892,N_2237,N_2417);
xnor U5893 (N_5893,N_3715,N_3381);
or U5894 (N_5894,N_2036,N_2518);
nor U5895 (N_5895,N_2515,N_2743);
nor U5896 (N_5896,N_2083,N_3777);
and U5897 (N_5897,N_2584,N_2804);
nand U5898 (N_5898,N_2162,N_3023);
nor U5899 (N_5899,N_2119,N_3713);
nor U5900 (N_5900,N_3458,N_2362);
or U5901 (N_5901,N_3039,N_2861);
nor U5902 (N_5902,N_2992,N_3024);
nor U5903 (N_5903,N_3075,N_3735);
nand U5904 (N_5904,N_2084,N_3651);
or U5905 (N_5905,N_3229,N_2488);
or U5906 (N_5906,N_3327,N_3169);
and U5907 (N_5907,N_2752,N_2565);
or U5908 (N_5908,N_2877,N_2655);
and U5909 (N_5909,N_2964,N_2844);
or U5910 (N_5910,N_3827,N_2143);
nor U5911 (N_5911,N_2443,N_2284);
nand U5912 (N_5912,N_2133,N_3289);
or U5913 (N_5913,N_3032,N_3732);
or U5914 (N_5914,N_2495,N_3863);
nand U5915 (N_5915,N_3366,N_3013);
and U5916 (N_5916,N_2757,N_2060);
or U5917 (N_5917,N_3672,N_2962);
nand U5918 (N_5918,N_2573,N_3220);
and U5919 (N_5919,N_3718,N_2468);
or U5920 (N_5920,N_3029,N_3476);
or U5921 (N_5921,N_2006,N_2522);
or U5922 (N_5922,N_2023,N_2772);
and U5923 (N_5923,N_3636,N_2725);
and U5924 (N_5924,N_3056,N_3203);
or U5925 (N_5925,N_3084,N_3774);
and U5926 (N_5926,N_3490,N_2512);
xor U5927 (N_5927,N_2495,N_2281);
nor U5928 (N_5928,N_3487,N_2894);
or U5929 (N_5929,N_2571,N_3300);
nor U5930 (N_5930,N_2752,N_3275);
nand U5931 (N_5931,N_2331,N_2044);
nand U5932 (N_5932,N_2204,N_2561);
nor U5933 (N_5933,N_2892,N_2540);
nor U5934 (N_5934,N_2584,N_2456);
or U5935 (N_5935,N_3464,N_3455);
nor U5936 (N_5936,N_2405,N_2461);
and U5937 (N_5937,N_3258,N_2501);
or U5938 (N_5938,N_2251,N_2801);
xnor U5939 (N_5939,N_2122,N_3932);
or U5940 (N_5940,N_3680,N_3345);
nand U5941 (N_5941,N_3776,N_2452);
nor U5942 (N_5942,N_2563,N_2423);
nand U5943 (N_5943,N_3492,N_2947);
nor U5944 (N_5944,N_2488,N_3978);
nand U5945 (N_5945,N_3701,N_3277);
or U5946 (N_5946,N_3372,N_2869);
and U5947 (N_5947,N_2923,N_3391);
or U5948 (N_5948,N_2685,N_3639);
nor U5949 (N_5949,N_3990,N_2156);
nand U5950 (N_5950,N_2224,N_3809);
xor U5951 (N_5951,N_3897,N_3753);
nand U5952 (N_5952,N_3264,N_3824);
xor U5953 (N_5953,N_2854,N_3053);
nor U5954 (N_5954,N_2805,N_3010);
or U5955 (N_5955,N_2952,N_3423);
and U5956 (N_5956,N_3167,N_2511);
nand U5957 (N_5957,N_3270,N_2221);
or U5958 (N_5958,N_2434,N_2938);
xor U5959 (N_5959,N_2556,N_2514);
nand U5960 (N_5960,N_3974,N_2531);
and U5961 (N_5961,N_2746,N_3571);
and U5962 (N_5962,N_2452,N_3107);
or U5963 (N_5963,N_2113,N_2046);
nor U5964 (N_5964,N_2733,N_3820);
xor U5965 (N_5965,N_2436,N_2946);
xor U5966 (N_5966,N_2682,N_3855);
and U5967 (N_5967,N_2287,N_3027);
and U5968 (N_5968,N_3602,N_3267);
or U5969 (N_5969,N_2197,N_3263);
nor U5970 (N_5970,N_3105,N_3729);
nor U5971 (N_5971,N_3155,N_3375);
nor U5972 (N_5972,N_2846,N_2343);
nor U5973 (N_5973,N_3396,N_2686);
nor U5974 (N_5974,N_2743,N_3219);
or U5975 (N_5975,N_3427,N_2543);
nand U5976 (N_5976,N_3871,N_3005);
or U5977 (N_5977,N_3911,N_3574);
nor U5978 (N_5978,N_3338,N_2352);
and U5979 (N_5979,N_2932,N_2615);
xnor U5980 (N_5980,N_3327,N_3059);
and U5981 (N_5981,N_3216,N_2852);
and U5982 (N_5982,N_3476,N_3101);
and U5983 (N_5983,N_3526,N_2512);
nand U5984 (N_5984,N_2160,N_2315);
nand U5985 (N_5985,N_3335,N_3168);
xnor U5986 (N_5986,N_3229,N_2337);
nand U5987 (N_5987,N_3059,N_2003);
nor U5988 (N_5988,N_3405,N_2480);
nor U5989 (N_5989,N_2077,N_2083);
nand U5990 (N_5990,N_3276,N_2464);
and U5991 (N_5991,N_2934,N_2793);
nor U5992 (N_5992,N_3103,N_2685);
and U5993 (N_5993,N_3714,N_3995);
nor U5994 (N_5994,N_2394,N_3924);
nor U5995 (N_5995,N_3624,N_2076);
or U5996 (N_5996,N_2880,N_3362);
nor U5997 (N_5997,N_2095,N_3871);
or U5998 (N_5998,N_2045,N_3203);
nor U5999 (N_5999,N_2484,N_2344);
nand U6000 (N_6000,N_4723,N_5043);
or U6001 (N_6001,N_4103,N_4364);
or U6002 (N_6002,N_4847,N_5791);
and U6003 (N_6003,N_4708,N_5998);
xnor U6004 (N_6004,N_4016,N_4309);
nand U6005 (N_6005,N_4340,N_5696);
or U6006 (N_6006,N_4948,N_4085);
or U6007 (N_6007,N_5124,N_4277);
or U6008 (N_6008,N_4183,N_4589);
nor U6009 (N_6009,N_4453,N_4147);
or U6010 (N_6010,N_5955,N_4933);
nor U6011 (N_6011,N_5214,N_5751);
nand U6012 (N_6012,N_5721,N_4499);
xnor U6013 (N_6013,N_5767,N_4189);
nand U6014 (N_6014,N_4638,N_4654);
nand U6015 (N_6015,N_5636,N_5780);
nand U6016 (N_6016,N_4730,N_4455);
nor U6017 (N_6017,N_4547,N_5677);
nand U6018 (N_6018,N_5291,N_5611);
and U6019 (N_6019,N_4439,N_5670);
and U6020 (N_6020,N_5096,N_5429);
nand U6021 (N_6021,N_5774,N_4172);
nand U6022 (N_6022,N_4432,N_5699);
or U6023 (N_6023,N_4395,N_5901);
nor U6024 (N_6024,N_5257,N_4670);
nand U6025 (N_6025,N_5606,N_5837);
xnor U6026 (N_6026,N_4668,N_5757);
nand U6027 (N_6027,N_4086,N_4662);
or U6028 (N_6028,N_4351,N_4625);
and U6029 (N_6029,N_4749,N_4816);
and U6030 (N_6030,N_5603,N_5404);
nand U6031 (N_6031,N_4032,N_4304);
nand U6032 (N_6032,N_4377,N_5815);
and U6033 (N_6033,N_5111,N_4078);
and U6034 (N_6034,N_4812,N_5331);
and U6035 (N_6035,N_4899,N_4821);
nand U6036 (N_6036,N_5804,N_5294);
nand U6037 (N_6037,N_5547,N_4554);
nor U6038 (N_6038,N_4953,N_5682);
and U6039 (N_6039,N_5763,N_4817);
nand U6040 (N_6040,N_5741,N_4731);
or U6041 (N_6041,N_5252,N_4229);
xor U6042 (N_6042,N_5969,N_5660);
nand U6043 (N_6043,N_4409,N_5044);
nand U6044 (N_6044,N_5614,N_5458);
or U6045 (N_6045,N_5217,N_4041);
and U6046 (N_6046,N_5383,N_5920);
or U6047 (N_6047,N_5876,N_4047);
nand U6048 (N_6048,N_5673,N_4891);
and U6049 (N_6049,N_5539,N_4145);
or U6050 (N_6050,N_5373,N_5959);
nor U6051 (N_6051,N_5307,N_4746);
or U6052 (N_6052,N_5720,N_5716);
and U6053 (N_6053,N_5196,N_4838);
and U6054 (N_6054,N_5836,N_4688);
or U6055 (N_6055,N_4140,N_5719);
nor U6056 (N_6056,N_5874,N_4242);
or U6057 (N_6057,N_5320,N_4563);
and U6058 (N_6058,N_4516,N_5066);
nand U6059 (N_6059,N_5266,N_5330);
nor U6060 (N_6060,N_5916,N_5678);
or U6061 (N_6061,N_5830,N_4157);
or U6062 (N_6062,N_5370,N_4408);
and U6063 (N_6063,N_4760,N_5665);
nor U6064 (N_6064,N_5563,N_4162);
and U6065 (N_6065,N_5122,N_5050);
nand U6066 (N_6066,N_5733,N_5166);
nor U6067 (N_6067,N_5645,N_4387);
nor U6068 (N_6068,N_4384,N_4988);
nor U6069 (N_6069,N_5988,N_5604);
or U6070 (N_6070,N_5597,N_5258);
and U6071 (N_6071,N_5642,N_4813);
or U6072 (N_6072,N_5332,N_4835);
nand U6073 (N_6073,N_4378,N_5193);
and U6074 (N_6074,N_4431,N_4217);
xor U6075 (N_6075,N_4867,N_5149);
nor U6076 (N_6076,N_5263,N_5361);
nor U6077 (N_6077,N_5034,N_5686);
nand U6078 (N_6078,N_4941,N_4770);
xnor U6079 (N_6079,N_4976,N_5036);
or U6080 (N_6080,N_4262,N_4514);
nor U6081 (N_6081,N_4295,N_4343);
nor U6082 (N_6082,N_5651,N_5760);
nor U6083 (N_6083,N_5662,N_5843);
nand U6084 (N_6084,N_4287,N_5299);
or U6085 (N_6085,N_4366,N_5004);
xnor U6086 (N_6086,N_4596,N_5706);
xor U6087 (N_6087,N_5045,N_4942);
nand U6088 (N_6088,N_4112,N_5703);
or U6089 (N_6089,N_5411,N_4567);
or U6090 (N_6090,N_4440,N_4703);
or U6091 (N_6091,N_5279,N_5346);
nand U6092 (N_6092,N_4080,N_5438);
and U6093 (N_6093,N_5672,N_5977);
and U6094 (N_6094,N_4744,N_5701);
or U6095 (N_6095,N_4270,N_4187);
or U6096 (N_6096,N_5226,N_5020);
nand U6097 (N_6097,N_4535,N_5726);
nand U6098 (N_6098,N_5349,N_5579);
nor U6099 (N_6099,N_5509,N_5165);
and U6100 (N_6100,N_5067,N_5156);
or U6101 (N_6101,N_4268,N_5758);
nand U6102 (N_6102,N_4360,N_5061);
or U6103 (N_6103,N_4079,N_4743);
and U6104 (N_6104,N_4370,N_4115);
nor U6105 (N_6105,N_5181,N_4274);
nor U6106 (N_6106,N_4578,N_5211);
nand U6107 (N_6107,N_5759,N_5355);
nand U6108 (N_6108,N_4796,N_4206);
xor U6109 (N_6109,N_4982,N_5039);
xor U6110 (N_6110,N_4222,N_4125);
nand U6111 (N_6111,N_5494,N_4237);
nand U6112 (N_6112,N_4250,N_4128);
nand U6113 (N_6113,N_4960,N_5556);
or U6114 (N_6114,N_5419,N_5956);
and U6115 (N_6115,N_5182,N_4335);
nor U6116 (N_6116,N_5881,N_4594);
nor U6117 (N_6117,N_5629,N_4861);
or U6118 (N_6118,N_4799,N_4834);
and U6119 (N_6119,N_4163,N_5054);
xor U6120 (N_6120,N_5350,N_5930);
nor U6121 (N_6121,N_5794,N_4342);
xnor U6122 (N_6122,N_5431,N_5126);
or U6123 (N_6123,N_5971,N_5272);
and U6124 (N_6124,N_4735,N_5778);
or U6125 (N_6125,N_4236,N_4068);
and U6126 (N_6126,N_4918,N_5869);
or U6127 (N_6127,N_5492,N_4152);
nor U6128 (N_6128,N_4191,N_4987);
nand U6129 (N_6129,N_5308,N_4774);
or U6130 (N_6130,N_4042,N_4221);
or U6131 (N_6131,N_4204,N_4561);
and U6132 (N_6132,N_5255,N_4102);
and U6133 (N_6133,N_5100,N_4122);
nand U6134 (N_6134,N_5136,N_4859);
nand U6135 (N_6135,N_5797,N_5380);
and U6136 (N_6136,N_5293,N_4996);
nor U6137 (N_6137,N_4716,N_5410);
nand U6138 (N_6138,N_4851,N_5533);
nor U6139 (N_6139,N_4488,N_5209);
or U6140 (N_6140,N_5465,N_4509);
nand U6141 (N_6141,N_5644,N_5418);
nand U6142 (N_6142,N_5074,N_4846);
or U6143 (N_6143,N_5188,N_4321);
nand U6144 (N_6144,N_5773,N_5345);
nor U6145 (N_6145,N_5273,N_5110);
nand U6146 (N_6146,N_4031,N_4572);
and U6147 (N_6147,N_5484,N_4069);
and U6148 (N_6148,N_4092,N_5530);
nor U6149 (N_6149,N_5745,N_4510);
and U6150 (N_6150,N_5982,N_5595);
nand U6151 (N_6151,N_4880,N_5184);
or U6152 (N_6152,N_4995,N_4185);
nand U6153 (N_6153,N_5864,N_4350);
nor U6154 (N_6154,N_4361,N_4544);
nand U6155 (N_6155,N_5551,N_5992);
or U6156 (N_6156,N_4886,N_4029);
and U6157 (N_6157,N_4738,N_4628);
and U6158 (N_6158,N_4761,N_5063);
xor U6159 (N_6159,N_5498,N_4952);
xor U6160 (N_6160,N_5659,N_4494);
nor U6161 (N_6161,N_4758,N_4515);
or U6162 (N_6162,N_5860,N_4144);
xnor U6163 (N_6163,N_5285,N_5236);
and U6164 (N_6164,N_5878,N_5402);
nor U6165 (N_6165,N_5582,N_5933);
nor U6166 (N_6166,N_4419,N_4975);
and U6167 (N_6167,N_4444,N_5886);
nand U6168 (N_6168,N_4930,N_4986);
and U6169 (N_6169,N_5693,N_4026);
and U6170 (N_6170,N_4734,N_5295);
and U6171 (N_6171,N_5967,N_4365);
or U6172 (N_6172,N_4403,N_5416);
nand U6173 (N_6173,N_4393,N_5189);
nor U6174 (N_6174,N_5812,N_4776);
and U6175 (N_6175,N_4061,N_4265);
nor U6176 (N_6176,N_4246,N_5123);
nor U6177 (N_6177,N_4566,N_4665);
and U6178 (N_6178,N_5506,N_5489);
or U6179 (N_6179,N_4329,N_5347);
or U6180 (N_6180,N_5839,N_4917);
and U6181 (N_6181,N_4754,N_4777);
nor U6182 (N_6182,N_5769,N_4195);
nor U6183 (N_6183,N_4482,N_5367);
or U6184 (N_6184,N_5951,N_5101);
and U6185 (N_6185,N_4955,N_5808);
nand U6186 (N_6186,N_4306,N_5022);
nor U6187 (N_6187,N_4194,N_5552);
and U6188 (N_6188,N_5796,N_4402);
nand U6189 (N_6189,N_4282,N_5499);
nor U6190 (N_6190,N_5602,N_5208);
or U6191 (N_6191,N_5568,N_5042);
nor U6192 (N_6192,N_5392,N_5212);
or U6193 (N_6193,N_4339,N_4223);
or U6194 (N_6194,N_5927,N_4491);
nand U6195 (N_6195,N_4755,N_5639);
nand U6196 (N_6196,N_4705,N_4921);
and U6197 (N_6197,N_4788,N_5608);
xor U6198 (N_6198,N_5816,N_5577);
nand U6199 (N_6199,N_4373,N_4814);
nand U6200 (N_6200,N_4700,N_5931);
and U6201 (N_6201,N_4720,N_4564);
or U6202 (N_6202,N_5961,N_4245);
and U6203 (N_6203,N_4584,N_4363);
or U6204 (N_6204,N_5792,N_5174);
nor U6205 (N_6205,N_5278,N_4990);
or U6206 (N_6206,N_4833,N_4965);
and U6207 (N_6207,N_5460,N_5439);
and U6208 (N_6208,N_4649,N_4279);
or U6209 (N_6209,N_5232,N_5264);
nand U6210 (N_6210,N_5766,N_4780);
xor U6211 (N_6211,N_4998,N_4215);
and U6212 (N_6212,N_4934,N_5496);
or U6213 (N_6213,N_4374,N_5996);
or U6214 (N_6214,N_4548,N_4712);
or U6215 (N_6215,N_4117,N_5409);
or U6216 (N_6216,N_5432,N_5650);
or U6217 (N_6217,N_5870,N_4619);
or U6218 (N_6218,N_5875,N_5964);
nor U6219 (N_6219,N_4660,N_5146);
nand U6220 (N_6220,N_5178,N_4003);
and U6221 (N_6221,N_4493,N_5323);
or U6222 (N_6222,N_5075,N_5296);
or U6223 (N_6223,N_4093,N_4354);
and U6224 (N_6224,N_4475,N_5055);
and U6225 (N_6225,N_4655,N_5443);
and U6226 (N_6226,N_4260,N_4071);
xor U6227 (N_6227,N_5403,N_4303);
and U6228 (N_6228,N_5097,N_5134);
or U6229 (N_6229,N_4517,N_5938);
xnor U6230 (N_6230,N_5633,N_4599);
and U6231 (N_6231,N_4938,N_5789);
and U6232 (N_6232,N_4511,N_5274);
nand U6233 (N_6233,N_5301,N_5396);
or U6234 (N_6234,N_4994,N_5398);
xor U6235 (N_6235,N_4503,N_4525);
and U6236 (N_6236,N_4243,N_5049);
nor U6237 (N_6237,N_5840,N_5793);
and U6238 (N_6238,N_5851,N_4894);
nand U6239 (N_6239,N_5343,N_4296);
nand U6240 (N_6240,N_4099,N_4508);
nor U6241 (N_6241,N_4862,N_4434);
nand U6242 (N_6242,N_4970,N_4849);
xor U6243 (N_6243,N_5973,N_5480);
nand U6244 (N_6244,N_5080,N_5685);
nor U6245 (N_6245,N_4985,N_4005);
and U6246 (N_6246,N_4549,N_5401);
and U6247 (N_6247,N_4954,N_4090);
nor U6248 (N_6248,N_4436,N_4878);
or U6249 (N_6249,N_4631,N_4136);
or U6250 (N_6250,N_4214,N_4196);
xor U6251 (N_6251,N_5456,N_5923);
nand U6252 (N_6252,N_5717,N_4701);
nor U6253 (N_6253,N_5817,N_4368);
or U6254 (N_6254,N_5708,N_5203);
nand U6255 (N_6255,N_5434,N_4044);
or U6256 (N_6256,N_5655,N_5483);
nand U6257 (N_6257,N_5736,N_4652);
nand U6258 (N_6258,N_4010,N_5085);
or U6259 (N_6259,N_4745,N_5880);
nor U6260 (N_6260,N_5035,N_4696);
or U6261 (N_6261,N_4231,N_5377);
nand U6262 (N_6262,N_4801,N_4359);
nor U6263 (N_6263,N_5822,N_4661);
nor U6264 (N_6264,N_5150,N_4273);
nor U6265 (N_6265,N_5374,N_5504);
nand U6266 (N_6266,N_5479,N_5463);
and U6267 (N_6267,N_4528,N_5848);
nand U6268 (N_6268,N_5186,N_5737);
or U6269 (N_6269,N_4672,N_4857);
or U6270 (N_6270,N_4272,N_4523);
or U6271 (N_6271,N_5173,N_4981);
nor U6272 (N_6272,N_5247,N_5368);
or U6273 (N_6273,N_4173,N_5095);
xor U6274 (N_6274,N_5753,N_4487);
nand U6275 (N_6275,N_5536,N_5302);
and U6276 (N_6276,N_5240,N_4627);
and U6277 (N_6277,N_4490,N_5040);
nor U6278 (N_6278,N_4641,N_5872);
and U6279 (N_6279,N_5909,N_4910);
nand U6280 (N_6280,N_5306,N_5338);
xnor U6281 (N_6281,N_4219,N_4445);
nor U6282 (N_6282,N_4967,N_5527);
nand U6283 (N_6283,N_4133,N_5810);
xnor U6284 (N_6284,N_5157,N_4526);
or U6285 (N_6285,N_4401,N_4969);
nand U6286 (N_6286,N_4858,N_4827);
xnor U6287 (N_6287,N_5104,N_4682);
nor U6288 (N_6288,N_5185,N_5477);
nor U6289 (N_6289,N_5092,N_4275);
or U6290 (N_6290,N_5995,N_4602);
and U6291 (N_6291,N_5929,N_5038);
and U6292 (N_6292,N_4873,N_5855);
or U6293 (N_6293,N_4116,N_4956);
xor U6294 (N_6294,N_5129,N_5994);
or U6295 (N_6295,N_4227,N_4964);
nor U6296 (N_6296,N_5567,N_4959);
nand U6297 (N_6297,N_5592,N_4288);
nand U6298 (N_6298,N_4650,N_4038);
nand U6299 (N_6299,N_4860,N_4966);
nand U6300 (N_6300,N_4771,N_5856);
and U6301 (N_6301,N_5356,N_5534);
nor U6302 (N_6302,N_5825,N_4310);
or U6303 (N_6303,N_5687,N_5697);
nand U6304 (N_6304,N_5554,N_4576);
and U6305 (N_6305,N_4454,N_5105);
and U6306 (N_6306,N_5116,N_5674);
nor U6307 (N_6307,N_5109,N_4841);
xnor U6308 (N_6308,N_4480,N_4100);
nor U6309 (N_6309,N_5298,N_5421);
or U6310 (N_6310,N_4946,N_4485);
or U6311 (N_6311,N_5382,N_5254);
or U6312 (N_6312,N_5544,N_4664);
or U6313 (N_6313,N_4890,N_5029);
and U6314 (N_6314,N_4466,N_5190);
nor U6315 (N_6315,N_4551,N_5915);
nand U6316 (N_6316,N_4875,N_4083);
and U6317 (N_6317,N_5788,N_5102);
and U6318 (N_6318,N_4175,N_5500);
nor U6319 (N_6319,N_5106,N_4823);
or U6320 (N_6320,N_4114,N_5897);
and U6321 (N_6321,N_4865,N_4600);
and U6322 (N_6322,N_5495,N_5657);
or U6323 (N_6323,N_4106,N_4369);
and U6324 (N_6324,N_5844,N_5318);
or U6325 (N_6325,N_5724,N_4607);
xor U6326 (N_6326,N_4477,N_5680);
and U6327 (N_6327,N_5654,N_4063);
nor U6328 (N_6328,N_4714,N_4597);
nor U6329 (N_6329,N_5922,N_4824);
nand U6330 (N_6330,N_5470,N_5940);
or U6331 (N_6331,N_5945,N_5569);
xnor U6332 (N_6332,N_4543,N_4165);
xor U6333 (N_6333,N_5112,N_4685);
nor U6334 (N_6334,N_4529,N_4601);
nand U6335 (N_6335,N_5099,N_4422);
nand U6336 (N_6336,N_4385,N_5128);
and U6337 (N_6337,N_4129,N_5221);
and U6338 (N_6338,N_5161,N_5454);
xnor U6339 (N_6339,N_5053,N_4291);
and U6340 (N_6340,N_4240,N_4922);
nand U6341 (N_6341,N_4271,N_5289);
and U6342 (N_6342,N_5183,N_5947);
or U6343 (N_6343,N_4171,N_5535);
nand U6344 (N_6344,N_4328,N_5518);
nand U6345 (N_6345,N_4898,N_4552);
nand U6346 (N_6346,N_5246,N_4647);
or U6347 (N_6347,N_5032,N_4610);
nand U6348 (N_6348,N_4747,N_4235);
and U6349 (N_6349,N_4149,N_4141);
or U6350 (N_6350,N_5118,N_4009);
nor U6351 (N_6351,N_5525,N_4980);
nor U6352 (N_6352,N_4629,N_4201);
nor U6353 (N_6353,N_4298,N_4239);
xor U6354 (N_6354,N_5847,N_5227);
nor U6355 (N_6355,N_4389,N_5200);
or U6356 (N_6356,N_4159,N_4341);
or U6357 (N_6357,N_4143,N_5414);
nand U6358 (N_6358,N_5026,N_4430);
nand U6359 (N_6359,N_4199,N_5508);
nor U6360 (N_6360,N_5877,N_5607);
and U6361 (N_6361,N_4810,N_5671);
and U6362 (N_6362,N_5406,N_4333);
nand U6363 (N_6363,N_5459,N_5485);
nand U6364 (N_6364,N_5175,N_5892);
nor U6365 (N_6365,N_4459,N_5060);
xnor U6366 (N_6366,N_5317,N_5906);
nor U6367 (N_6367,N_4974,N_4392);
or U6368 (N_6368,N_4615,N_5167);
nand U6369 (N_6369,N_5290,N_4557);
and U6370 (N_6370,N_4766,N_4656);
and U6371 (N_6371,N_5658,N_4104);
xnor U6372 (N_6372,N_5714,N_4920);
or U6373 (N_6373,N_4166,N_4943);
and U6374 (N_6374,N_4391,N_5222);
nand U6375 (N_6375,N_4507,N_4313);
and U6376 (N_6376,N_4586,N_4055);
nor U6377 (N_6377,N_5805,N_4822);
nor U6378 (N_6378,N_4299,N_4151);
or U6379 (N_6379,N_4539,N_5133);
nand U6380 (N_6380,N_5315,N_4740);
and U6381 (N_6381,N_5850,N_5566);
nor U6382 (N_6382,N_5936,N_5275);
and U6383 (N_6383,N_5984,N_5863);
nand U6384 (N_6384,N_5632,N_5545);
and U6385 (N_6385,N_4840,N_5683);
nand U6386 (N_6386,N_4075,N_4283);
or U6387 (N_6387,N_4565,N_4793);
or U6388 (N_6388,N_4230,N_4791);
or U6389 (N_6389,N_4807,N_4786);
nor U6390 (N_6390,N_4863,N_5113);
nand U6391 (N_6391,N_5831,N_5276);
nor U6392 (N_6392,N_4019,N_4238);
nand U6393 (N_6393,N_4698,N_4376);
xnor U6394 (N_6394,N_5871,N_5366);
nand U6395 (N_6395,N_4438,N_5046);
nor U6396 (N_6396,N_5239,N_5268);
or U6397 (N_6397,N_5466,N_4137);
xor U6398 (N_6398,N_4164,N_4218);
or U6399 (N_6399,N_5625,N_5488);
nand U6400 (N_6400,N_4018,N_4887);
nand U6401 (N_6401,N_4778,N_5070);
and U6402 (N_6402,N_4498,N_5250);
or U6403 (N_6403,N_5084,N_4689);
and U6404 (N_6404,N_4150,N_5088);
and U6405 (N_6405,N_5337,N_4739);
nor U6406 (N_6406,N_5647,N_4254);
or U6407 (N_6407,N_4465,N_5051);
nor U6408 (N_6408,N_5441,N_5482);
or U6409 (N_6409,N_4205,N_4410);
nor U6410 (N_6410,N_4530,N_4521);
xor U6411 (N_6411,N_5888,N_4330);
nor U6412 (N_6412,N_4721,N_5771);
nand U6413 (N_6413,N_5169,N_5283);
and U6414 (N_6414,N_5444,N_4573);
and U6415 (N_6415,N_4736,N_4914);
nand U6416 (N_6416,N_4322,N_5761);
nor U6417 (N_6417,N_5896,N_4879);
xor U6418 (N_6418,N_4289,N_5605);
nand U6419 (N_6419,N_4435,N_4612);
and U6420 (N_6420,N_5435,N_4888);
nand U6421 (N_6421,N_4800,N_4297);
nor U6422 (N_6422,N_4462,N_5882);
and U6423 (N_6423,N_5790,N_4624);
or U6424 (N_6424,N_5231,N_4470);
nor U6425 (N_6425,N_4179,N_4923);
nand U6426 (N_6426,N_4947,N_4028);
and U6427 (N_6427,N_5823,N_5388);
nor U6428 (N_6428,N_4932,N_5198);
and U6429 (N_6429,N_5442,N_5939);
xnor U6430 (N_6430,N_4259,N_4502);
nor U6431 (N_6431,N_4913,N_5225);
and U6432 (N_6432,N_4476,N_4193);
and U6433 (N_6433,N_5164,N_4866);
xor U6434 (N_6434,N_4854,N_5369);
or U6435 (N_6435,N_5142,N_4611);
nand U6436 (N_6436,N_4371,N_5835);
and U6437 (N_6437,N_5244,N_5627);
nor U6438 (N_6438,N_5024,N_5065);
nor U6439 (N_6439,N_4234,N_5970);
or U6440 (N_6440,N_5584,N_4675);
nand U6441 (N_6441,N_5091,N_5433);
nor U6442 (N_6442,N_5979,N_5912);
nor U6443 (N_6443,N_5462,N_5626);
or U6444 (N_6444,N_4101,N_5224);
and U6445 (N_6445,N_5172,N_5571);
or U6446 (N_6446,N_4541,N_4323);
nand U6447 (N_6447,N_4950,N_5314);
and U6448 (N_6448,N_5461,N_4856);
or U6449 (N_6449,N_5017,N_4842);
or U6450 (N_6450,N_4447,N_4790);
or U6451 (N_6451,N_4496,N_5081);
and U6452 (N_6452,N_5891,N_5827);
and U6453 (N_6453,N_5452,N_4292);
or U6454 (N_6454,N_5505,N_5137);
or U6455 (N_6455,N_5451,N_4519);
and U6456 (N_6456,N_4072,N_4651);
nor U6457 (N_6457,N_5574,N_5430);
nand U6458 (N_6458,N_5309,N_5140);
or U6459 (N_6459,N_4935,N_5709);
nand U6460 (N_6460,N_5474,N_5715);
nor U6461 (N_6461,N_4811,N_4278);
nor U6462 (N_6462,N_5132,N_5313);
and U6463 (N_6463,N_5422,N_4285);
and U6464 (N_6464,N_4836,N_5623);
or U6465 (N_6465,N_4358,N_4848);
nand U6466 (N_6466,N_5842,N_4871);
nor U6467 (N_6467,N_5027,N_4706);
nand U6468 (N_6468,N_4691,N_5179);
or U6469 (N_6469,N_4460,N_4011);
or U6470 (N_6470,N_5408,N_4677);
or U6471 (N_6471,N_4829,N_4451);
or U6472 (N_6472,N_5256,N_5321);
xor U6473 (N_6473,N_5130,N_5640);
or U6474 (N_6474,N_5555,N_4481);
and U6475 (N_6475,N_5204,N_5637);
nand U6476 (N_6476,N_5513,N_5354);
nor U6477 (N_6477,N_4639,N_5233);
and U6478 (N_6478,N_4684,N_5609);
nand U6479 (N_6479,N_5006,N_5543);
or U6480 (N_6480,N_5748,N_5712);
or U6481 (N_6481,N_4052,N_4489);
xor U6482 (N_6482,N_4412,N_4174);
nor U6483 (N_6483,N_5980,N_4725);
nand U6484 (N_6484,N_5905,N_5335);
xnor U6485 (N_6485,N_5286,N_4659);
or U6486 (N_6486,N_4002,N_5756);
nor U6487 (N_6487,N_4520,N_5229);
nand U6488 (N_6488,N_5676,N_5824);
or U6489 (N_6489,N_5903,N_5010);
nand U6490 (N_6490,N_5553,N_5372);
or U6491 (N_6491,N_5491,N_5087);
and U6492 (N_6492,N_4901,N_4006);
and U6493 (N_6493,N_5652,N_5007);
nor U6494 (N_6494,N_4819,N_5012);
nor U6495 (N_6495,N_5427,N_4414);
and U6496 (N_6496,N_4156,N_4686);
or U6497 (N_6497,N_4896,N_4906);
and U6498 (N_6498,N_5379,N_4417);
nor U6499 (N_6499,N_5516,N_4756);
nand U6500 (N_6500,N_4357,N_5475);
or U6501 (N_6501,N_5919,N_4198);
or U6502 (N_6502,N_4545,N_5587);
or U6503 (N_6503,N_4828,N_5859);
or U6504 (N_6504,N_5524,N_5037);
xor U6505 (N_6505,N_4021,N_4580);
and U6506 (N_6506,N_4560,N_4537);
nor U6507 (N_6507,N_4184,N_4603);
or U6508 (N_6508,N_5910,N_5103);
or U6509 (N_6509,N_5585,N_4792);
and U6510 (N_6510,N_5962,N_4690);
nor U6511 (N_6511,N_4642,N_5834);
nor U6512 (N_6512,N_4484,N_5245);
nor U6513 (N_6513,N_4023,N_4407);
nor U6514 (N_6514,N_5885,N_4046);
or U6515 (N_6515,N_5618,N_4673);
nor U6516 (N_6516,N_5785,N_5924);
nor U6517 (N_6517,N_5052,N_5328);
and U6518 (N_6518,N_5925,N_4495);
and U6519 (N_6519,N_5394,N_4999);
and U6520 (N_6520,N_5503,N_5216);
or U6521 (N_6521,N_4207,N_5478);
or U6522 (N_6522,N_5643,N_5968);
and U6523 (N_6523,N_5127,N_4614);
and U6524 (N_6524,N_5818,N_5391);
or U6525 (N_6525,N_4895,N_5420);
nor U6526 (N_6526,N_5481,N_5739);
nor U6527 (N_6527,N_4033,N_4681);
or U6528 (N_6528,N_4795,N_5852);
or U6529 (N_6529,N_4066,N_5151);
nand U6530 (N_6530,N_5900,N_4680);
nand U6531 (N_6531,N_5238,N_5201);
xor U6532 (N_6532,N_4804,N_4711);
or U6533 (N_6533,N_4893,N_5206);
and U6534 (N_6534,N_5453,N_5357);
nand U6535 (N_6535,N_5600,N_4362);
nand U6536 (N_6536,N_4697,N_5235);
nor U6537 (N_6537,N_5363,N_4931);
or U6538 (N_6538,N_4424,N_4057);
or U6539 (N_6539,N_4413,N_5730);
or U6540 (N_6540,N_5734,N_5879);
and U6541 (N_6541,N_5983,N_4785);
or U6542 (N_6542,N_4160,N_4989);
or U6543 (N_6543,N_5468,N_4324);
or U6544 (N_6544,N_5768,N_4794);
and U6545 (N_6545,N_4513,N_4135);
and U6546 (N_6546,N_5809,N_4098);
and U6547 (N_6547,N_5918,N_5664);
or U6548 (N_6548,N_4067,N_5476);
nor U6549 (N_6549,N_4750,N_4581);
xor U6550 (N_6550,N_4280,N_5634);
or U6551 (N_6551,N_4618,N_4443);
nor U6552 (N_6552,N_4782,N_5661);
or U6553 (N_6553,N_4437,N_4375);
xnor U6554 (N_6554,N_5727,N_5192);
nand U6555 (N_6555,N_4134,N_4830);
nand U6556 (N_6556,N_4609,N_5400);
and U6557 (N_6557,N_5436,N_4345);
nor U6558 (N_6558,N_5141,N_4383);
or U6559 (N_6559,N_5329,N_4138);
nor U6560 (N_6560,N_4399,N_5125);
nor U6561 (N_6561,N_4924,N_4263);
xnor U6562 (N_6562,N_4765,N_4852);
nand U6563 (N_6563,N_5570,N_5344);
and U6564 (N_6564,N_5679,N_4884);
xnor U6565 (N_6565,N_5288,N_5941);
nand U6566 (N_6566,N_5580,N_4261);
or U6567 (N_6567,N_5009,N_4188);
and U6568 (N_6568,N_4082,N_4468);
and U6569 (N_6569,N_4062,N_5324);
nor U6570 (N_6570,N_5467,N_5943);
and U6571 (N_6571,N_4595,N_5270);
or U6572 (N_6572,N_5068,N_4077);
or U6573 (N_6573,N_5950,N_4326);
or U6574 (N_6574,N_5334,N_4110);
nand U6575 (N_6575,N_5949,N_4772);
xor U6576 (N_6576,N_4043,N_5907);
nor U6577 (N_6577,N_5393,N_4962);
and U6578 (N_6578,N_5199,N_5079);
nor U6579 (N_6579,N_5194,N_4497);
or U6580 (N_6580,N_4971,N_4168);
xor U6581 (N_6581,N_5493,N_4949);
or U6582 (N_6582,N_4623,N_5445);
or U6583 (N_6583,N_4864,N_4719);
nor U6584 (N_6584,N_5280,N_5407);
and U6585 (N_6585,N_5803,N_5972);
or U6586 (N_6586,N_4534,N_4542);
nor U6587 (N_6587,N_4267,N_5153);
or U6588 (N_6588,N_5913,N_4787);
or U6589 (N_6589,N_5845,N_5312);
and U6590 (N_6590,N_5887,N_5548);
or U6591 (N_6591,N_5935,N_5364);
nor U6592 (N_6592,N_5071,N_5292);
and U6593 (N_6593,N_4524,N_5001);
nor U6594 (N_6594,N_5147,N_5205);
nor U6595 (N_6595,N_4726,N_4676);
and U6596 (N_6596,N_4233,N_5028);
or U6597 (N_6597,N_4958,N_4784);
or U6598 (N_6598,N_5740,N_5832);
nor U6599 (N_6599,N_4056,N_5025);
nand U6600 (N_6600,N_5779,N_5596);
or U6601 (N_6601,N_4640,N_5180);
nand U6602 (N_6602,N_4094,N_5378);
or U6603 (N_6603,N_4569,N_4732);
nand U6604 (N_6604,N_5326,N_4308);
and U6605 (N_6605,N_4874,N_5615);
or U6606 (N_6606,N_5828,N_5381);
nor U6607 (N_6607,N_5772,N_5707);
and U6608 (N_6608,N_5914,N_4433);
or U6609 (N_6609,N_4653,N_5041);
nand U6610 (N_6610,N_5646,N_4646);
and U6611 (N_6611,N_5215,N_5237);
xnor U6612 (N_6612,N_4728,N_4553);
and U6613 (N_6613,N_5365,N_5705);
nor U6614 (N_6614,N_5019,N_5520);
nor U6615 (N_6615,N_5348,N_5561);
or U6616 (N_6616,N_5207,N_4479);
nor U6617 (N_6617,N_5359,N_5993);
nand U6618 (N_6618,N_4161,N_5656);
or U6619 (N_6619,N_4096,N_4605);
or U6620 (N_6620,N_4251,N_5135);
xnor U6621 (N_6621,N_5762,N_4928);
and U6622 (N_6622,N_5210,N_5976);
and U6623 (N_6623,N_5523,N_5853);
and U6624 (N_6624,N_4753,N_4826);
xor U6625 (N_6625,N_5163,N_5144);
nand U6626 (N_6626,N_5575,N_4346);
nor U6627 (N_6627,N_5251,N_4571);
and U6628 (N_6628,N_4327,N_5883);
and U6629 (N_6629,N_5729,N_4153);
xnor U6630 (N_6630,N_5528,N_5937);
nor U6631 (N_6631,N_4390,N_4416);
xnor U6632 (N_6632,N_5058,N_5814);
and U6633 (N_6633,N_4314,N_5997);
nor U6634 (N_6634,N_5387,N_5322);
nand U6635 (N_6635,N_5742,N_5316);
and U6636 (N_6636,N_5838,N_4773);
and U6637 (N_6637,N_4064,N_4504);
nor U6638 (N_6638,N_4636,N_5073);
nand U6639 (N_6639,N_4818,N_4825);
or U6640 (N_6640,N_4767,N_5541);
or U6641 (N_6641,N_5395,N_4939);
or U6642 (N_6642,N_5090,N_4317);
or U6643 (N_6643,N_4900,N_5351);
nor U6644 (N_6644,N_4048,N_4978);
and U6645 (N_6645,N_5963,N_5002);
xor U6646 (N_6646,N_5865,N_4319);
and U6647 (N_6647,N_4775,N_5710);
and U6648 (N_6648,N_4170,N_4718);
and U6649 (N_6649,N_5559,N_5704);
xor U6650 (N_6650,N_4577,N_4574);
and U6651 (N_6651,N_5800,N_5787);
or U6652 (N_6652,N_5958,N_5108);
or U6653 (N_6653,N_4717,N_4051);
nor U6654 (N_6654,N_5743,N_4216);
nand U6655 (N_6655,N_4501,N_4590);
and U6656 (N_6656,N_4281,N_4902);
or U6657 (N_6657,N_4815,N_5271);
nand U6658 (N_6658,N_4853,N_5265);
nand U6659 (N_6659,N_4058,N_4182);
and U6660 (N_6660,N_4457,N_4926);
or U6661 (N_6661,N_4148,N_5069);
nand U6662 (N_6662,N_5668,N_5911);
and U6663 (N_6663,N_4752,N_5904);
or U6664 (N_6664,N_4474,N_5449);
nand U6665 (N_6665,N_4617,N_5841);
or U6666 (N_6666,N_5448,N_4264);
xor U6667 (N_6667,N_4331,N_5613);
or U6668 (N_6668,N_5098,N_5486);
nor U6669 (N_6669,N_5187,N_4616);
or U6670 (N_6670,N_5228,N_4500);
and U6671 (N_6671,N_4225,N_4429);
and U6672 (N_6672,N_5738,N_4907);
and U6673 (N_6673,N_5138,N_4256);
nor U6674 (N_6674,N_4748,N_5287);
xor U6675 (N_6675,N_5728,N_5532);
and U6676 (N_6676,N_4411,N_5564);
nand U6677 (N_6677,N_4126,N_4940);
or U6678 (N_6678,N_4559,N_5953);
nor U6679 (N_6679,N_5056,N_5281);
and U6680 (N_6680,N_4017,N_5806);
and U6681 (N_6681,N_5735,N_5114);
nor U6682 (N_6682,N_4737,N_5638);
nor U6683 (N_6683,N_4155,N_4876);
or U6684 (N_6684,N_5786,N_4423);
nand U6685 (N_6685,N_4769,N_4583);
nand U6686 (N_6686,N_5170,N_5519);
and U6687 (N_6687,N_5243,N_5089);
or U6688 (N_6688,N_5415,N_4972);
and U6689 (N_6689,N_5107,N_5784);
nor U6690 (N_6690,N_4763,N_5159);
or U6691 (N_6691,N_4178,N_5340);
or U6692 (N_6692,N_5957,N_4355);
nand U6693 (N_6693,N_5457,N_4845);
or U6694 (N_6694,N_5512,N_5003);
nor U6695 (N_6695,N_5471,N_5873);
or U6696 (N_6696,N_4425,N_4802);
xnor U6697 (N_6697,N_5898,N_5277);
xor U6698 (N_6698,N_5667,N_4709);
and U6699 (N_6699,N_5581,N_4040);
and U6700 (N_6700,N_5576,N_5731);
or U6701 (N_6701,N_4911,N_4582);
nand U6702 (N_6702,N_4013,N_4789);
or U6703 (N_6703,N_4404,N_4905);
nand U6704 (N_6704,N_4266,N_4305);
nor U6705 (N_6705,N_4892,N_5781);
or U6706 (N_6706,N_5948,N_4742);
and U6707 (N_6707,N_5782,N_4593);
nor U6708 (N_6708,N_4088,N_5586);
nor U6709 (N_6709,N_4883,N_5752);
nand U6710 (N_6710,N_4693,N_5148);
or U6711 (N_6711,N_5426,N_5325);
nand U6712 (N_6712,N_4108,N_4154);
nor U6713 (N_6713,N_5725,N_5588);
nor U6714 (N_6714,N_5540,N_4951);
nor U6715 (N_6715,N_5487,N_5016);
nand U6716 (N_6716,N_4585,N_5399);
and U6717 (N_6717,N_5511,N_4473);
and U6718 (N_6718,N_4398,N_4645);
or U6719 (N_6719,N_4027,N_5261);
or U6720 (N_6720,N_4555,N_5849);
nand U6721 (N_6721,N_4556,N_4606);
nand U6722 (N_6722,N_5692,N_4197);
nor U6723 (N_6723,N_5526,N_5249);
and U6724 (N_6724,N_5560,N_4348);
or U6725 (N_6725,N_4707,N_4715);
and U6726 (N_6726,N_5057,N_4741);
and U6727 (N_6727,N_4505,N_4123);
nand U6728 (N_6728,N_4200,N_4781);
nand U6729 (N_6729,N_4284,N_5424);
nor U6730 (N_6730,N_4868,N_5744);
or U6731 (N_6731,N_4307,N_4118);
nor U6732 (N_6732,N_5455,N_5619);
nand U6733 (N_6733,N_5700,N_4400);
and U6734 (N_6734,N_4927,N_5946);
and U6735 (N_6735,N_5267,N_5902);
nand U6736 (N_6736,N_4427,N_4025);
or U6737 (N_6737,N_4226,N_4192);
nand U6738 (N_6738,N_4426,N_5008);
and U6739 (N_6739,N_5549,N_5213);
nor U6740 (N_6740,N_5620,N_5801);
nand U6741 (N_6741,N_4805,N_4255);
xnor U6742 (N_6742,N_5158,N_5558);
or U6743 (N_6743,N_4084,N_4783);
and U6744 (N_6744,N_4146,N_5353);
or U6745 (N_6745,N_4727,N_4211);
nand U6746 (N_6746,N_4300,N_5064);
nor U6747 (N_6747,N_5732,N_5775);
and U6748 (N_6748,N_4983,N_4167);
nand U6749 (N_6749,N_4059,N_4558);
nor U6750 (N_6750,N_5573,N_4562);
nand U6751 (N_6751,N_5746,N_5684);
or U6752 (N_6752,N_4591,N_5405);
nand U6753 (N_6753,N_5230,N_5154);
xnor U6754 (N_6754,N_4347,N_4344);
and U6755 (N_6755,N_4997,N_4367);
or U6756 (N_6756,N_4420,N_5932);
nor U6757 (N_6757,N_4657,N_5305);
or U6758 (N_6758,N_5799,N_5965);
and U6759 (N_6759,N_4957,N_4352);
nand U6760 (N_6760,N_4020,N_4109);
and U6761 (N_6761,N_4729,N_5152);
xnor U6762 (N_6762,N_4014,N_4724);
and U6763 (N_6763,N_5327,N_5867);
nand U6764 (N_6764,N_5833,N_5770);
nand U6765 (N_6765,N_5975,N_5718);
and U6766 (N_6766,N_4269,N_4850);
and U6767 (N_6767,N_5985,N_4442);
nor U6768 (N_6768,N_5986,N_4658);
and U6769 (N_6769,N_5021,N_5723);
and U6770 (N_6770,N_5764,N_4337);
nor U6771 (N_6771,N_5776,N_5546);
xnor U6772 (N_6772,N_4472,N_4483);
nor U6773 (N_6773,N_5145,N_4081);
nor U6774 (N_6774,N_5310,N_4695);
nand U6775 (N_6775,N_4963,N_4353);
and U6776 (N_6776,N_4637,N_4000);
and U6777 (N_6777,N_5005,N_5688);
nor U6778 (N_6778,N_5282,N_4702);
nor U6779 (N_6779,N_5829,N_5162);
or U6780 (N_6780,N_4806,N_5062);
nor U6781 (N_6781,N_4415,N_5333);
nor U6782 (N_6782,N_4916,N_4049);
nand U6783 (N_6783,N_4325,N_4318);
and U6784 (N_6784,N_4276,N_4808);
and U6785 (N_6785,N_4379,N_4798);
or U6786 (N_6786,N_4486,N_5059);
nand U6787 (N_6787,N_5926,N_4803);
and U6788 (N_6788,N_5978,N_5990);
xor U6789 (N_6789,N_4441,N_4598);
nand U6790 (N_6790,N_5339,N_5622);
nand U6791 (N_6791,N_4091,N_4113);
and U6792 (N_6792,N_4293,N_4004);
nand U6793 (N_6793,N_4540,N_5413);
xnor U6794 (N_6794,N_5531,N_5358);
nor U6795 (N_6795,N_4111,N_4692);
or U6796 (N_6796,N_4396,N_4478);
nand U6797 (N_6797,N_5537,N_5412);
nor U6798 (N_6798,N_4944,N_4158);
nand U6799 (N_6799,N_5259,N_5669);
or U6800 (N_6800,N_4448,N_4620);
xor U6801 (N_6801,N_4679,N_4608);
nor U6802 (N_6802,N_4418,N_4666);
nor U6803 (N_6803,N_5031,N_5663);
nor U6804 (N_6804,N_5497,N_5397);
and U6805 (N_6805,N_5242,N_4461);
xnor U6806 (N_6806,N_4381,N_4034);
nand U6807 (N_6807,N_4797,N_4388);
nor U6808 (N_6808,N_4522,N_5417);
and U6809 (N_6809,N_5934,N_4039);
nand U6810 (N_6810,N_5423,N_5078);
xnor U6811 (N_6811,N_4877,N_5854);
and U6812 (N_6812,N_4973,N_4855);
nor U6813 (N_6813,N_5675,N_4604);
nand U6814 (N_6814,N_4904,N_4587);
and U6815 (N_6815,N_5813,N_5428);
nor U6816 (N_6816,N_4181,N_4132);
xor U6817 (N_6817,N_5262,N_5820);
nand U6818 (N_6818,N_4394,N_5018);
nor U6819 (N_6819,N_5681,N_5641);
xor U6820 (N_6820,N_5472,N_4915);
and U6821 (N_6821,N_5030,N_4382);
and U6822 (N_6822,N_4632,N_5572);
nand U6823 (N_6823,N_5908,N_4015);
or U6824 (N_6824,N_5304,N_4671);
nand U6825 (N_6825,N_5297,N_5015);
or U6826 (N_6826,N_5371,N_5115);
nor U6827 (N_6827,N_4065,N_4286);
and U6828 (N_6828,N_4630,N_4213);
and U6829 (N_6829,N_4037,N_5218);
nor U6830 (N_6830,N_5033,N_5469);
nor U6831 (N_6831,N_5749,N_5522);
nor U6832 (N_6832,N_4456,N_4130);
nor U6833 (N_6833,N_5966,N_5866);
nor U6834 (N_6834,N_4993,N_5464);
or U6835 (N_6835,N_4209,N_4127);
or U6836 (N_6836,N_4142,N_4180);
nand U6837 (N_6837,N_4315,N_5944);
or U6838 (N_6838,N_5093,N_5047);
or U6839 (N_6839,N_4648,N_4527);
xnor U6840 (N_6840,N_5889,N_5599);
nand U6841 (N_6841,N_4882,N_5450);
xnor U6842 (N_6842,N_5750,N_4053);
and U6843 (N_6843,N_5284,N_5589);
and U6844 (N_6844,N_4699,N_4839);
nor U6845 (N_6845,N_5076,N_5648);
and U6846 (N_6846,N_4030,N_4449);
and U6847 (N_6847,N_4634,N_4012);
xnor U6848 (N_6848,N_4311,N_5593);
nor U6849 (N_6849,N_4302,N_5514);
and U6850 (N_6850,N_4991,N_5253);
nor U6851 (N_6851,N_4506,N_5942);
or U6852 (N_6852,N_5385,N_4228);
nand U6853 (N_6853,N_4249,N_4809);
nand U6854 (N_6854,N_5974,N_4356);
xor U6855 (N_6855,N_5260,N_5755);
xnor U6856 (N_6856,N_4463,N_4757);
nor U6857 (N_6857,N_4961,N_4626);
nand U6858 (N_6858,N_4458,N_5077);
or U6859 (N_6859,N_4169,N_5538);
or U6860 (N_6860,N_5689,N_4687);
xnor U6861 (N_6861,N_5117,N_5072);
nor U6862 (N_6862,N_5311,N_4332);
nand U6863 (N_6863,N_5894,N_4570);
nor U6864 (N_6864,N_4945,N_5783);
nor U6865 (N_6865,N_5248,N_4467);
nor U6866 (N_6866,N_4397,N_4622);
xnor U6867 (N_6867,N_4452,N_4220);
and U6868 (N_6868,N_4405,N_5811);
nor U6869 (N_6869,N_4937,N_5219);
nor U6870 (N_6870,N_5868,N_4050);
or U6871 (N_6871,N_5490,N_4843);
nor U6872 (N_6872,N_4471,N_5846);
or U6873 (N_6873,N_4320,N_5501);
nand U6874 (N_6874,N_5360,N_5515);
nand U6875 (N_6875,N_5542,N_4203);
xnor U6876 (N_6876,N_4713,N_4536);
or U6877 (N_6877,N_4968,N_4889);
nor U6878 (N_6878,N_5352,N_5691);
nor U6879 (N_6879,N_4253,N_5698);
nor U6880 (N_6880,N_4621,N_4837);
nor U6881 (N_6881,N_4120,N_4241);
and U6882 (N_6882,N_5121,N_4669);
xnor U6883 (N_6883,N_5502,N_5425);
and U6884 (N_6884,N_4258,N_5594);
and U6885 (N_6885,N_5507,N_5139);
nor U6886 (N_6886,N_4119,N_4428);
nor U6887 (N_6887,N_5921,N_4678);
xnor U6888 (N_6888,N_4633,N_4912);
or U6889 (N_6889,N_5991,N_4095);
and U6890 (N_6890,N_4704,N_5191);
and U6891 (N_6891,N_5119,N_4045);
or U6892 (N_6892,N_5168,N_4532);
or U6893 (N_6893,N_4464,N_5389);
nor U6894 (N_6894,N_5362,N_5695);
or U6895 (N_6895,N_5048,N_4512);
xor U6896 (N_6896,N_5550,N_5384);
nor U6897 (N_6897,N_5754,N_5666);
or U6898 (N_6898,N_5083,N_5336);
or U6899 (N_6899,N_5023,N_5616);
and U6900 (N_6900,N_5375,N_5631);
nand U6901 (N_6901,N_5928,N_5234);
xor U6902 (N_6902,N_4208,N_4294);
and U6903 (N_6903,N_4244,N_4831);
xor U6904 (N_6904,N_5143,N_4232);
nor U6905 (N_6905,N_4349,N_4105);
nor U6906 (N_6906,N_4768,N_5447);
nand U6907 (N_6907,N_4764,N_5826);
nand U6908 (N_6908,N_4186,N_5694);
nor U6909 (N_6909,N_4024,N_4076);
nand U6910 (N_6910,N_5861,N_4733);
and U6911 (N_6911,N_5437,N_4533);
or U6912 (N_6912,N_5160,N_5510);
or U6913 (N_6913,N_4881,N_5899);
or U6914 (N_6914,N_5711,N_5197);
nand U6915 (N_6915,N_5202,N_5591);
nor U6916 (N_6916,N_5120,N_4176);
nor U6917 (N_6917,N_4872,N_4121);
xnor U6918 (N_6918,N_4210,N_4008);
or U6919 (N_6919,N_4252,N_4546);
or U6920 (N_6920,N_4469,N_4762);
nor U6921 (N_6921,N_4869,N_5517);
nand U6922 (N_6922,N_4592,N_4885);
nor U6923 (N_6923,N_5300,N_4759);
nand U6924 (N_6924,N_4290,N_5917);
or U6925 (N_6925,N_4124,N_4635);
xnor U6926 (N_6926,N_4054,N_4386);
and U6927 (N_6927,N_4036,N_5220);
and U6928 (N_6928,N_4257,N_4492);
nand U6929 (N_6929,N_4722,N_5981);
nor U6930 (N_6930,N_4316,N_4074);
xor U6931 (N_6931,N_5617,N_4060);
or U6932 (N_6932,N_4372,N_4674);
nor U6933 (N_6933,N_4202,N_5171);
xnor U6934 (N_6934,N_5557,N_4247);
xor U6935 (N_6935,N_5341,N_4936);
nor U6936 (N_6936,N_5960,N_5440);
nand U6937 (N_6937,N_5890,N_5082);
or U6938 (N_6938,N_5802,N_4683);
and U6939 (N_6939,N_5303,N_5086);
nand U6940 (N_6940,N_5386,N_5529);
xnor U6941 (N_6941,N_5195,N_5521);
xor U6942 (N_6942,N_5765,N_5562);
and U6943 (N_6943,N_4001,N_4925);
or U6944 (N_6944,N_5893,N_4550);
and U6945 (N_6945,N_4312,N_5747);
nand U6946 (N_6946,N_5999,N_5989);
or U6947 (N_6947,N_5653,N_5952);
xor U6948 (N_6948,N_4844,N_5342);
xor U6949 (N_6949,N_5954,N_5013);
and U6950 (N_6950,N_4575,N_5628);
and U6951 (N_6951,N_5690,N_4568);
or U6952 (N_6952,N_4336,N_5319);
nor U6953 (N_6953,N_5590,N_5884);
nor U6954 (N_6954,N_4977,N_4984);
or U6955 (N_6955,N_5777,N_5612);
or U6956 (N_6956,N_4089,N_5821);
or U6957 (N_6957,N_4643,N_4694);
nor U6958 (N_6958,N_5713,N_5446);
nand U6959 (N_6959,N_5987,N_4538);
nor U6960 (N_6960,N_5241,N_5895);
nand U6961 (N_6961,N_4908,N_4107);
nand U6962 (N_6962,N_5621,N_4779);
and U6963 (N_6963,N_5624,N_4903);
nor U6964 (N_6964,N_4909,N_4421);
and U6965 (N_6965,N_5390,N_4820);
or U6966 (N_6966,N_4644,N_5862);
nand U6967 (N_6967,N_4450,N_5094);
or U6968 (N_6968,N_5376,N_5630);
nor U6969 (N_6969,N_4212,N_5177);
nor U6970 (N_6970,N_4531,N_4832);
nand U6971 (N_6971,N_5000,N_5795);
nor U6972 (N_6972,N_5798,N_4667);
nand U6973 (N_6973,N_4406,N_4097);
xnor U6974 (N_6974,N_4301,N_5807);
nor U6975 (N_6975,N_5722,N_5565);
nor U6976 (N_6976,N_4518,N_4131);
or U6977 (N_6977,N_4929,N_5610);
and U6978 (N_6978,N_5601,N_5011);
or U6979 (N_6979,N_5858,N_5857);
and U6980 (N_6980,N_5223,N_4919);
and U6981 (N_6981,N_4248,N_4579);
nor U6982 (N_6982,N_5131,N_5583);
nand U6983 (N_6983,N_4446,N_4070);
and U6984 (N_6984,N_5702,N_4710);
or U6985 (N_6985,N_4139,N_5269);
and U6986 (N_6986,N_5014,N_5819);
and U6987 (N_6987,N_4022,N_4087);
and U6988 (N_6988,N_4073,N_5176);
and U6989 (N_6989,N_5635,N_5649);
and U6990 (N_6990,N_4224,N_4979);
or U6991 (N_6991,N_4338,N_4751);
nor U6992 (N_6992,N_4190,N_4870);
or U6993 (N_6993,N_4663,N_5155);
nand U6994 (N_6994,N_4380,N_5473);
or U6995 (N_6995,N_5578,N_4035);
xor U6996 (N_6996,N_4613,N_4897);
or U6997 (N_6997,N_4334,N_4992);
and U6998 (N_6998,N_4007,N_4177);
or U6999 (N_6999,N_5598,N_4588);
and U7000 (N_7000,N_5543,N_5257);
nand U7001 (N_7001,N_5010,N_5557);
or U7002 (N_7002,N_4314,N_5790);
nand U7003 (N_7003,N_5975,N_5526);
nand U7004 (N_7004,N_5173,N_5670);
xor U7005 (N_7005,N_4722,N_4996);
or U7006 (N_7006,N_4964,N_5370);
or U7007 (N_7007,N_4911,N_5741);
nand U7008 (N_7008,N_4909,N_4028);
and U7009 (N_7009,N_4051,N_4024);
and U7010 (N_7010,N_5234,N_5752);
nor U7011 (N_7011,N_5209,N_5133);
or U7012 (N_7012,N_4930,N_4504);
or U7013 (N_7013,N_4480,N_5996);
and U7014 (N_7014,N_4894,N_4956);
nand U7015 (N_7015,N_5903,N_5708);
nor U7016 (N_7016,N_5386,N_4436);
or U7017 (N_7017,N_5596,N_4394);
and U7018 (N_7018,N_4722,N_4071);
xor U7019 (N_7019,N_5097,N_4160);
and U7020 (N_7020,N_5820,N_5298);
or U7021 (N_7021,N_5255,N_5573);
and U7022 (N_7022,N_4665,N_4140);
or U7023 (N_7023,N_5551,N_4664);
nor U7024 (N_7024,N_5793,N_4232);
or U7025 (N_7025,N_5769,N_4519);
nand U7026 (N_7026,N_4319,N_4574);
nand U7027 (N_7027,N_4333,N_4885);
nor U7028 (N_7028,N_5006,N_5807);
or U7029 (N_7029,N_4119,N_5141);
or U7030 (N_7030,N_5714,N_4085);
nor U7031 (N_7031,N_4566,N_4015);
nor U7032 (N_7032,N_4501,N_5938);
nor U7033 (N_7033,N_4612,N_4829);
nand U7034 (N_7034,N_5135,N_5430);
nor U7035 (N_7035,N_4479,N_5926);
nor U7036 (N_7036,N_5604,N_4194);
nor U7037 (N_7037,N_4278,N_4063);
or U7038 (N_7038,N_4084,N_4215);
and U7039 (N_7039,N_5704,N_5012);
nor U7040 (N_7040,N_4533,N_4871);
and U7041 (N_7041,N_4986,N_4718);
or U7042 (N_7042,N_4120,N_5270);
nor U7043 (N_7043,N_4773,N_4014);
and U7044 (N_7044,N_4815,N_4205);
nand U7045 (N_7045,N_4554,N_5174);
nand U7046 (N_7046,N_5815,N_5113);
nand U7047 (N_7047,N_5757,N_5394);
or U7048 (N_7048,N_5892,N_5402);
and U7049 (N_7049,N_4930,N_5339);
nand U7050 (N_7050,N_5860,N_4234);
nor U7051 (N_7051,N_4640,N_5611);
nand U7052 (N_7052,N_5425,N_5047);
nor U7053 (N_7053,N_4244,N_5386);
xor U7054 (N_7054,N_5665,N_4183);
nand U7055 (N_7055,N_5940,N_4530);
or U7056 (N_7056,N_4592,N_4488);
nor U7057 (N_7057,N_4039,N_5043);
and U7058 (N_7058,N_5134,N_4475);
or U7059 (N_7059,N_4012,N_4927);
nor U7060 (N_7060,N_4801,N_5140);
nand U7061 (N_7061,N_5620,N_4927);
xnor U7062 (N_7062,N_5130,N_5625);
nor U7063 (N_7063,N_4978,N_5883);
and U7064 (N_7064,N_5138,N_5525);
or U7065 (N_7065,N_5422,N_5103);
nand U7066 (N_7066,N_4760,N_4478);
nand U7067 (N_7067,N_5734,N_4556);
nand U7068 (N_7068,N_4264,N_4123);
and U7069 (N_7069,N_4401,N_5917);
or U7070 (N_7070,N_5341,N_4812);
nor U7071 (N_7071,N_4479,N_5708);
nor U7072 (N_7072,N_5945,N_4286);
nand U7073 (N_7073,N_5317,N_4698);
nor U7074 (N_7074,N_5689,N_5884);
nor U7075 (N_7075,N_4750,N_4718);
or U7076 (N_7076,N_5427,N_4840);
xor U7077 (N_7077,N_5657,N_4274);
or U7078 (N_7078,N_4351,N_4137);
and U7079 (N_7079,N_4805,N_5104);
nand U7080 (N_7080,N_4002,N_5738);
or U7081 (N_7081,N_5426,N_4759);
or U7082 (N_7082,N_5297,N_5390);
and U7083 (N_7083,N_5833,N_4877);
nand U7084 (N_7084,N_4357,N_5908);
and U7085 (N_7085,N_5111,N_4864);
nor U7086 (N_7086,N_5036,N_5171);
or U7087 (N_7087,N_5149,N_4916);
xnor U7088 (N_7088,N_4779,N_5409);
nor U7089 (N_7089,N_5109,N_4386);
nor U7090 (N_7090,N_4210,N_5224);
nor U7091 (N_7091,N_4210,N_5642);
nand U7092 (N_7092,N_5137,N_4936);
nand U7093 (N_7093,N_4496,N_5164);
and U7094 (N_7094,N_5308,N_5878);
and U7095 (N_7095,N_5233,N_5438);
or U7096 (N_7096,N_4063,N_5299);
nand U7097 (N_7097,N_4456,N_5195);
or U7098 (N_7098,N_4033,N_5709);
nand U7099 (N_7099,N_5127,N_5860);
nand U7100 (N_7100,N_5060,N_5648);
or U7101 (N_7101,N_4766,N_5358);
and U7102 (N_7102,N_5963,N_5478);
and U7103 (N_7103,N_4974,N_5104);
and U7104 (N_7104,N_4164,N_4562);
nor U7105 (N_7105,N_4756,N_4506);
nor U7106 (N_7106,N_4338,N_5133);
nand U7107 (N_7107,N_5581,N_5125);
and U7108 (N_7108,N_4557,N_4048);
nand U7109 (N_7109,N_4005,N_5677);
xor U7110 (N_7110,N_5847,N_4836);
or U7111 (N_7111,N_4826,N_5275);
xnor U7112 (N_7112,N_5381,N_4925);
nand U7113 (N_7113,N_5394,N_5957);
nand U7114 (N_7114,N_4505,N_4981);
xnor U7115 (N_7115,N_4007,N_5002);
and U7116 (N_7116,N_5644,N_5834);
xor U7117 (N_7117,N_4209,N_5267);
or U7118 (N_7118,N_5027,N_5347);
or U7119 (N_7119,N_4472,N_5381);
nor U7120 (N_7120,N_4006,N_4406);
or U7121 (N_7121,N_5361,N_4107);
nor U7122 (N_7122,N_5040,N_5351);
nor U7123 (N_7123,N_4246,N_4348);
or U7124 (N_7124,N_4513,N_5905);
xor U7125 (N_7125,N_4377,N_4980);
and U7126 (N_7126,N_4384,N_5124);
nor U7127 (N_7127,N_4032,N_5221);
nand U7128 (N_7128,N_4851,N_4429);
or U7129 (N_7129,N_4099,N_4167);
nor U7130 (N_7130,N_5717,N_5969);
and U7131 (N_7131,N_5758,N_4663);
or U7132 (N_7132,N_5461,N_5460);
nor U7133 (N_7133,N_4351,N_5055);
and U7134 (N_7134,N_5755,N_4054);
nor U7135 (N_7135,N_5643,N_5215);
nand U7136 (N_7136,N_4625,N_5443);
and U7137 (N_7137,N_4621,N_5027);
nor U7138 (N_7138,N_5284,N_5315);
and U7139 (N_7139,N_5627,N_5539);
xnor U7140 (N_7140,N_4082,N_5299);
nand U7141 (N_7141,N_4647,N_5339);
or U7142 (N_7142,N_5685,N_4834);
and U7143 (N_7143,N_5939,N_5980);
nor U7144 (N_7144,N_4823,N_4043);
nand U7145 (N_7145,N_5233,N_5638);
or U7146 (N_7146,N_4769,N_5550);
nor U7147 (N_7147,N_4430,N_4553);
and U7148 (N_7148,N_4751,N_5041);
or U7149 (N_7149,N_4648,N_5364);
and U7150 (N_7150,N_5593,N_5058);
nor U7151 (N_7151,N_5058,N_4455);
and U7152 (N_7152,N_5749,N_4903);
or U7153 (N_7153,N_4695,N_5389);
and U7154 (N_7154,N_5657,N_5176);
and U7155 (N_7155,N_4052,N_5828);
nand U7156 (N_7156,N_5102,N_5539);
and U7157 (N_7157,N_4003,N_4593);
or U7158 (N_7158,N_4382,N_5674);
nor U7159 (N_7159,N_5797,N_4929);
or U7160 (N_7160,N_5312,N_5884);
nor U7161 (N_7161,N_5048,N_5728);
nor U7162 (N_7162,N_5509,N_5866);
xor U7163 (N_7163,N_4073,N_4595);
nand U7164 (N_7164,N_5762,N_4261);
and U7165 (N_7165,N_5148,N_5905);
nand U7166 (N_7166,N_5575,N_5341);
and U7167 (N_7167,N_5610,N_5023);
xor U7168 (N_7168,N_4655,N_5537);
nand U7169 (N_7169,N_5408,N_4989);
or U7170 (N_7170,N_4657,N_4945);
and U7171 (N_7171,N_5810,N_5717);
nor U7172 (N_7172,N_4900,N_5334);
nor U7173 (N_7173,N_4264,N_4626);
nor U7174 (N_7174,N_5577,N_5723);
or U7175 (N_7175,N_5371,N_4109);
nor U7176 (N_7176,N_5592,N_5174);
or U7177 (N_7177,N_4598,N_4147);
nor U7178 (N_7178,N_5176,N_5474);
or U7179 (N_7179,N_4062,N_5654);
nand U7180 (N_7180,N_4314,N_5587);
nor U7181 (N_7181,N_4368,N_5548);
and U7182 (N_7182,N_5284,N_5506);
and U7183 (N_7183,N_5457,N_4753);
xor U7184 (N_7184,N_5868,N_4763);
or U7185 (N_7185,N_5979,N_4974);
and U7186 (N_7186,N_4381,N_4554);
nor U7187 (N_7187,N_5417,N_4324);
or U7188 (N_7188,N_5743,N_4900);
nand U7189 (N_7189,N_4991,N_5798);
or U7190 (N_7190,N_5227,N_4049);
nor U7191 (N_7191,N_5850,N_5480);
and U7192 (N_7192,N_5653,N_4734);
nand U7193 (N_7193,N_5870,N_4758);
nor U7194 (N_7194,N_4124,N_5733);
or U7195 (N_7195,N_5370,N_5690);
nand U7196 (N_7196,N_5405,N_5021);
or U7197 (N_7197,N_5408,N_5142);
and U7198 (N_7198,N_5059,N_4277);
xnor U7199 (N_7199,N_4295,N_4225);
and U7200 (N_7200,N_4516,N_5670);
or U7201 (N_7201,N_5432,N_4374);
and U7202 (N_7202,N_4069,N_5984);
nand U7203 (N_7203,N_5718,N_4326);
or U7204 (N_7204,N_5721,N_5213);
and U7205 (N_7205,N_4594,N_5507);
or U7206 (N_7206,N_5490,N_4183);
nor U7207 (N_7207,N_4557,N_5186);
nor U7208 (N_7208,N_5026,N_4696);
nand U7209 (N_7209,N_5424,N_4352);
and U7210 (N_7210,N_5380,N_5291);
or U7211 (N_7211,N_4105,N_4311);
or U7212 (N_7212,N_5344,N_4737);
nor U7213 (N_7213,N_4113,N_5093);
and U7214 (N_7214,N_4071,N_4488);
xnor U7215 (N_7215,N_5227,N_4593);
and U7216 (N_7216,N_4395,N_4204);
nor U7217 (N_7217,N_5995,N_4849);
nand U7218 (N_7218,N_4971,N_5745);
nand U7219 (N_7219,N_4568,N_5705);
nor U7220 (N_7220,N_4757,N_5957);
and U7221 (N_7221,N_5696,N_4871);
nor U7222 (N_7222,N_4098,N_5115);
nand U7223 (N_7223,N_4193,N_4523);
nor U7224 (N_7224,N_5773,N_4815);
nand U7225 (N_7225,N_5817,N_4327);
nand U7226 (N_7226,N_5958,N_4561);
nand U7227 (N_7227,N_5198,N_4666);
xnor U7228 (N_7228,N_4070,N_4549);
and U7229 (N_7229,N_5149,N_5446);
and U7230 (N_7230,N_5001,N_5395);
xnor U7231 (N_7231,N_4741,N_4026);
and U7232 (N_7232,N_5453,N_4039);
or U7233 (N_7233,N_4237,N_5564);
nand U7234 (N_7234,N_4874,N_5265);
xor U7235 (N_7235,N_5355,N_5994);
and U7236 (N_7236,N_4740,N_4576);
and U7237 (N_7237,N_5803,N_4131);
and U7238 (N_7238,N_4588,N_4920);
or U7239 (N_7239,N_5969,N_4870);
or U7240 (N_7240,N_5007,N_4159);
or U7241 (N_7241,N_5112,N_4568);
nand U7242 (N_7242,N_4521,N_4485);
nor U7243 (N_7243,N_5732,N_4692);
and U7244 (N_7244,N_4136,N_5970);
and U7245 (N_7245,N_5443,N_4500);
and U7246 (N_7246,N_5699,N_4395);
nor U7247 (N_7247,N_4100,N_4711);
nor U7248 (N_7248,N_4486,N_4026);
and U7249 (N_7249,N_5126,N_5685);
nand U7250 (N_7250,N_4614,N_4428);
and U7251 (N_7251,N_5885,N_5856);
nor U7252 (N_7252,N_5980,N_5199);
nor U7253 (N_7253,N_5592,N_4210);
xor U7254 (N_7254,N_4976,N_5898);
xor U7255 (N_7255,N_4609,N_4856);
xor U7256 (N_7256,N_4031,N_5558);
and U7257 (N_7257,N_4871,N_5858);
nand U7258 (N_7258,N_4479,N_4681);
nor U7259 (N_7259,N_5964,N_5141);
xor U7260 (N_7260,N_5331,N_4999);
and U7261 (N_7261,N_4156,N_5844);
or U7262 (N_7262,N_5127,N_4700);
nand U7263 (N_7263,N_5658,N_5626);
nand U7264 (N_7264,N_4978,N_4281);
and U7265 (N_7265,N_4209,N_4490);
xor U7266 (N_7266,N_4860,N_4035);
and U7267 (N_7267,N_5651,N_4049);
nand U7268 (N_7268,N_5092,N_4990);
and U7269 (N_7269,N_5514,N_4217);
nor U7270 (N_7270,N_5724,N_4581);
and U7271 (N_7271,N_4476,N_4577);
nor U7272 (N_7272,N_4867,N_5717);
nor U7273 (N_7273,N_5461,N_5214);
nor U7274 (N_7274,N_5965,N_4938);
and U7275 (N_7275,N_4230,N_5530);
nand U7276 (N_7276,N_5220,N_5247);
xnor U7277 (N_7277,N_4085,N_4049);
or U7278 (N_7278,N_4398,N_4808);
nand U7279 (N_7279,N_5820,N_4605);
xnor U7280 (N_7280,N_5573,N_5250);
and U7281 (N_7281,N_4107,N_5072);
or U7282 (N_7282,N_5572,N_4376);
and U7283 (N_7283,N_4519,N_5160);
nand U7284 (N_7284,N_5994,N_4507);
or U7285 (N_7285,N_5053,N_4911);
nand U7286 (N_7286,N_5060,N_5569);
nor U7287 (N_7287,N_5457,N_4386);
nand U7288 (N_7288,N_4051,N_5650);
nand U7289 (N_7289,N_4550,N_4721);
and U7290 (N_7290,N_4543,N_5513);
or U7291 (N_7291,N_5287,N_5671);
or U7292 (N_7292,N_5525,N_4114);
xor U7293 (N_7293,N_5676,N_5834);
xor U7294 (N_7294,N_5429,N_5044);
nor U7295 (N_7295,N_5914,N_4215);
and U7296 (N_7296,N_5449,N_5649);
nor U7297 (N_7297,N_5903,N_5880);
nand U7298 (N_7298,N_5711,N_4099);
nor U7299 (N_7299,N_4645,N_4512);
nand U7300 (N_7300,N_5779,N_4722);
and U7301 (N_7301,N_4979,N_5882);
nand U7302 (N_7302,N_4975,N_5995);
and U7303 (N_7303,N_4070,N_5302);
nand U7304 (N_7304,N_5506,N_5680);
and U7305 (N_7305,N_4024,N_4595);
or U7306 (N_7306,N_4986,N_4491);
xnor U7307 (N_7307,N_5508,N_5851);
or U7308 (N_7308,N_4510,N_5436);
nor U7309 (N_7309,N_4110,N_4009);
and U7310 (N_7310,N_4165,N_4131);
nand U7311 (N_7311,N_4275,N_4887);
or U7312 (N_7312,N_5339,N_5320);
and U7313 (N_7313,N_5509,N_5600);
or U7314 (N_7314,N_5872,N_4818);
xnor U7315 (N_7315,N_4793,N_4600);
nand U7316 (N_7316,N_4795,N_5084);
or U7317 (N_7317,N_4522,N_4875);
xor U7318 (N_7318,N_5364,N_5009);
nor U7319 (N_7319,N_5405,N_5801);
and U7320 (N_7320,N_4025,N_5921);
nand U7321 (N_7321,N_5424,N_4627);
and U7322 (N_7322,N_5672,N_4033);
or U7323 (N_7323,N_5931,N_5504);
nor U7324 (N_7324,N_5890,N_4624);
nand U7325 (N_7325,N_5782,N_4794);
nor U7326 (N_7326,N_5491,N_5584);
nand U7327 (N_7327,N_4126,N_5505);
or U7328 (N_7328,N_5401,N_5077);
nor U7329 (N_7329,N_5085,N_4043);
and U7330 (N_7330,N_4563,N_4218);
or U7331 (N_7331,N_4459,N_5955);
and U7332 (N_7332,N_5689,N_5249);
and U7333 (N_7333,N_5790,N_4656);
xnor U7334 (N_7334,N_5349,N_4943);
or U7335 (N_7335,N_5959,N_4876);
or U7336 (N_7336,N_4518,N_4648);
and U7337 (N_7337,N_5072,N_5525);
and U7338 (N_7338,N_5774,N_4960);
nand U7339 (N_7339,N_4565,N_4361);
and U7340 (N_7340,N_5064,N_5951);
nor U7341 (N_7341,N_4922,N_5115);
or U7342 (N_7342,N_5215,N_5784);
nand U7343 (N_7343,N_5797,N_4040);
and U7344 (N_7344,N_5600,N_5744);
or U7345 (N_7345,N_4951,N_4782);
nand U7346 (N_7346,N_5057,N_4148);
nand U7347 (N_7347,N_4369,N_5751);
xnor U7348 (N_7348,N_4513,N_4014);
or U7349 (N_7349,N_5454,N_4485);
or U7350 (N_7350,N_4378,N_5133);
nor U7351 (N_7351,N_5910,N_4465);
xor U7352 (N_7352,N_4995,N_4981);
nand U7353 (N_7353,N_5413,N_4615);
or U7354 (N_7354,N_5294,N_5716);
nor U7355 (N_7355,N_5982,N_5372);
nand U7356 (N_7356,N_5036,N_4498);
and U7357 (N_7357,N_4663,N_4770);
nor U7358 (N_7358,N_5082,N_4453);
or U7359 (N_7359,N_4455,N_4536);
and U7360 (N_7360,N_5944,N_5169);
nand U7361 (N_7361,N_4678,N_5950);
nor U7362 (N_7362,N_4325,N_5637);
nor U7363 (N_7363,N_5973,N_4906);
nand U7364 (N_7364,N_4887,N_4642);
and U7365 (N_7365,N_4683,N_5860);
and U7366 (N_7366,N_4695,N_4441);
and U7367 (N_7367,N_5620,N_5384);
xnor U7368 (N_7368,N_4134,N_4385);
or U7369 (N_7369,N_5900,N_5793);
nand U7370 (N_7370,N_4619,N_4070);
and U7371 (N_7371,N_5826,N_5688);
xnor U7372 (N_7372,N_4489,N_5681);
and U7373 (N_7373,N_4569,N_5888);
xor U7374 (N_7374,N_5967,N_5996);
xor U7375 (N_7375,N_4595,N_4366);
nand U7376 (N_7376,N_4961,N_5693);
nor U7377 (N_7377,N_5742,N_4044);
and U7378 (N_7378,N_4941,N_5652);
nor U7379 (N_7379,N_5508,N_4266);
nor U7380 (N_7380,N_4498,N_5711);
or U7381 (N_7381,N_5105,N_5631);
and U7382 (N_7382,N_4458,N_4779);
nor U7383 (N_7383,N_4963,N_5796);
and U7384 (N_7384,N_4804,N_4842);
nor U7385 (N_7385,N_5600,N_5004);
and U7386 (N_7386,N_5135,N_4077);
nor U7387 (N_7387,N_4725,N_4351);
nor U7388 (N_7388,N_4242,N_4126);
nor U7389 (N_7389,N_4393,N_5038);
or U7390 (N_7390,N_4167,N_4951);
or U7391 (N_7391,N_4722,N_4097);
and U7392 (N_7392,N_5505,N_4182);
nand U7393 (N_7393,N_4181,N_5949);
and U7394 (N_7394,N_4239,N_4595);
and U7395 (N_7395,N_4706,N_4211);
or U7396 (N_7396,N_5760,N_5719);
or U7397 (N_7397,N_4827,N_4386);
xor U7398 (N_7398,N_5567,N_5980);
or U7399 (N_7399,N_4427,N_5530);
or U7400 (N_7400,N_4244,N_4158);
nand U7401 (N_7401,N_4475,N_5146);
nand U7402 (N_7402,N_4018,N_5768);
nor U7403 (N_7403,N_4369,N_4037);
and U7404 (N_7404,N_4671,N_4391);
xnor U7405 (N_7405,N_4696,N_4195);
nor U7406 (N_7406,N_5205,N_4556);
and U7407 (N_7407,N_5940,N_5977);
or U7408 (N_7408,N_4383,N_4361);
nand U7409 (N_7409,N_5043,N_5970);
xnor U7410 (N_7410,N_4036,N_5053);
nand U7411 (N_7411,N_5916,N_5059);
nor U7412 (N_7412,N_5697,N_5416);
and U7413 (N_7413,N_4736,N_5744);
nand U7414 (N_7414,N_5924,N_5164);
or U7415 (N_7415,N_4948,N_4839);
and U7416 (N_7416,N_5171,N_4562);
or U7417 (N_7417,N_4600,N_4980);
nand U7418 (N_7418,N_4041,N_4312);
nor U7419 (N_7419,N_5583,N_5069);
nand U7420 (N_7420,N_5637,N_5758);
nor U7421 (N_7421,N_5489,N_4611);
and U7422 (N_7422,N_4254,N_5777);
nor U7423 (N_7423,N_4628,N_4645);
and U7424 (N_7424,N_4179,N_4385);
or U7425 (N_7425,N_5444,N_5047);
and U7426 (N_7426,N_4414,N_4567);
nor U7427 (N_7427,N_4998,N_4288);
nor U7428 (N_7428,N_5613,N_4305);
nand U7429 (N_7429,N_5081,N_4611);
nand U7430 (N_7430,N_4839,N_4652);
and U7431 (N_7431,N_4046,N_4018);
nand U7432 (N_7432,N_5525,N_5337);
xnor U7433 (N_7433,N_5851,N_4548);
or U7434 (N_7434,N_4275,N_5945);
nand U7435 (N_7435,N_5780,N_5539);
nor U7436 (N_7436,N_4098,N_5410);
or U7437 (N_7437,N_5626,N_4788);
nor U7438 (N_7438,N_4164,N_5972);
xnor U7439 (N_7439,N_4760,N_4049);
nand U7440 (N_7440,N_4947,N_5268);
nor U7441 (N_7441,N_5217,N_4197);
xnor U7442 (N_7442,N_5945,N_5506);
nor U7443 (N_7443,N_4033,N_5365);
xnor U7444 (N_7444,N_5105,N_5150);
and U7445 (N_7445,N_4597,N_4758);
nor U7446 (N_7446,N_5686,N_5719);
or U7447 (N_7447,N_4242,N_4912);
nor U7448 (N_7448,N_4777,N_5872);
and U7449 (N_7449,N_5792,N_4308);
and U7450 (N_7450,N_5709,N_4542);
and U7451 (N_7451,N_5255,N_4819);
xor U7452 (N_7452,N_4098,N_5731);
nor U7453 (N_7453,N_4231,N_4047);
xor U7454 (N_7454,N_4067,N_4694);
nor U7455 (N_7455,N_4375,N_4668);
xor U7456 (N_7456,N_4285,N_4797);
nand U7457 (N_7457,N_5286,N_4007);
xor U7458 (N_7458,N_4176,N_5234);
xnor U7459 (N_7459,N_5568,N_4144);
or U7460 (N_7460,N_5632,N_4164);
nor U7461 (N_7461,N_5381,N_4392);
nor U7462 (N_7462,N_4646,N_5856);
xor U7463 (N_7463,N_4052,N_4131);
and U7464 (N_7464,N_5395,N_4845);
or U7465 (N_7465,N_5431,N_5334);
and U7466 (N_7466,N_4253,N_4916);
nor U7467 (N_7467,N_4763,N_5112);
xor U7468 (N_7468,N_5586,N_4576);
or U7469 (N_7469,N_5260,N_4255);
nand U7470 (N_7470,N_5891,N_4062);
nor U7471 (N_7471,N_5693,N_5053);
nor U7472 (N_7472,N_4460,N_5149);
xor U7473 (N_7473,N_4546,N_5530);
xnor U7474 (N_7474,N_5828,N_5020);
nand U7475 (N_7475,N_5050,N_5407);
and U7476 (N_7476,N_5066,N_4762);
and U7477 (N_7477,N_4556,N_5047);
and U7478 (N_7478,N_4425,N_5652);
nand U7479 (N_7479,N_5519,N_4806);
nand U7480 (N_7480,N_5224,N_4322);
and U7481 (N_7481,N_4019,N_5945);
nor U7482 (N_7482,N_5435,N_5772);
or U7483 (N_7483,N_4405,N_5552);
nor U7484 (N_7484,N_5611,N_5013);
nor U7485 (N_7485,N_5421,N_4676);
and U7486 (N_7486,N_5994,N_4756);
nor U7487 (N_7487,N_4984,N_5777);
nand U7488 (N_7488,N_5866,N_5827);
or U7489 (N_7489,N_4405,N_5146);
or U7490 (N_7490,N_4907,N_4770);
and U7491 (N_7491,N_4193,N_5409);
xnor U7492 (N_7492,N_5023,N_4602);
nor U7493 (N_7493,N_5830,N_4631);
and U7494 (N_7494,N_5620,N_4240);
nor U7495 (N_7495,N_4792,N_4205);
and U7496 (N_7496,N_4241,N_5419);
nor U7497 (N_7497,N_5988,N_5764);
xnor U7498 (N_7498,N_5253,N_5462);
nor U7499 (N_7499,N_5180,N_5657);
and U7500 (N_7500,N_5277,N_5370);
and U7501 (N_7501,N_5560,N_4701);
xnor U7502 (N_7502,N_4132,N_5088);
or U7503 (N_7503,N_5990,N_4358);
nor U7504 (N_7504,N_4865,N_5367);
or U7505 (N_7505,N_4452,N_4897);
xnor U7506 (N_7506,N_4411,N_5916);
nand U7507 (N_7507,N_4429,N_4100);
nor U7508 (N_7508,N_5736,N_4350);
and U7509 (N_7509,N_5690,N_4762);
xor U7510 (N_7510,N_5412,N_4409);
or U7511 (N_7511,N_4135,N_5094);
and U7512 (N_7512,N_5352,N_4583);
xor U7513 (N_7513,N_5767,N_4689);
or U7514 (N_7514,N_5085,N_4879);
nand U7515 (N_7515,N_5921,N_4465);
or U7516 (N_7516,N_4425,N_4730);
and U7517 (N_7517,N_5643,N_4408);
or U7518 (N_7518,N_5197,N_5578);
nor U7519 (N_7519,N_4753,N_5173);
nand U7520 (N_7520,N_5736,N_4311);
or U7521 (N_7521,N_5498,N_5320);
nand U7522 (N_7522,N_4515,N_4264);
nor U7523 (N_7523,N_5946,N_5795);
nand U7524 (N_7524,N_5882,N_4763);
and U7525 (N_7525,N_4433,N_5272);
nor U7526 (N_7526,N_4723,N_4182);
xnor U7527 (N_7527,N_4863,N_4225);
and U7528 (N_7528,N_5823,N_5221);
nand U7529 (N_7529,N_4543,N_4699);
xnor U7530 (N_7530,N_4219,N_5224);
xnor U7531 (N_7531,N_5352,N_4399);
and U7532 (N_7532,N_5098,N_4107);
and U7533 (N_7533,N_5949,N_5374);
or U7534 (N_7534,N_5084,N_4052);
nor U7535 (N_7535,N_5260,N_4221);
nand U7536 (N_7536,N_4763,N_5505);
or U7537 (N_7537,N_5801,N_4608);
nand U7538 (N_7538,N_5883,N_4018);
xnor U7539 (N_7539,N_5900,N_4355);
or U7540 (N_7540,N_4391,N_5255);
or U7541 (N_7541,N_4793,N_5140);
or U7542 (N_7542,N_4678,N_5352);
and U7543 (N_7543,N_5347,N_5327);
and U7544 (N_7544,N_5177,N_4898);
and U7545 (N_7545,N_5455,N_4046);
or U7546 (N_7546,N_5580,N_5130);
nand U7547 (N_7547,N_4745,N_4375);
xor U7548 (N_7548,N_5758,N_5461);
nand U7549 (N_7549,N_4664,N_4412);
nand U7550 (N_7550,N_4889,N_5968);
and U7551 (N_7551,N_4519,N_4193);
xnor U7552 (N_7552,N_4324,N_4230);
or U7553 (N_7553,N_4362,N_5573);
and U7554 (N_7554,N_5044,N_5035);
nand U7555 (N_7555,N_5485,N_4258);
nand U7556 (N_7556,N_4779,N_4407);
or U7557 (N_7557,N_4448,N_4951);
nor U7558 (N_7558,N_5889,N_5499);
and U7559 (N_7559,N_4851,N_5186);
or U7560 (N_7560,N_5702,N_5808);
and U7561 (N_7561,N_5770,N_5394);
or U7562 (N_7562,N_4832,N_5929);
or U7563 (N_7563,N_4184,N_4613);
nor U7564 (N_7564,N_4333,N_5396);
or U7565 (N_7565,N_5295,N_5159);
and U7566 (N_7566,N_4898,N_4678);
and U7567 (N_7567,N_4469,N_5825);
nor U7568 (N_7568,N_5398,N_5325);
nor U7569 (N_7569,N_5122,N_5833);
or U7570 (N_7570,N_5767,N_4856);
and U7571 (N_7571,N_5271,N_5865);
and U7572 (N_7572,N_5950,N_5078);
or U7573 (N_7573,N_5677,N_4043);
and U7574 (N_7574,N_4468,N_4867);
or U7575 (N_7575,N_4794,N_5988);
nand U7576 (N_7576,N_5769,N_5115);
xor U7577 (N_7577,N_4428,N_4582);
nand U7578 (N_7578,N_4093,N_4854);
xor U7579 (N_7579,N_5689,N_4727);
and U7580 (N_7580,N_5089,N_4064);
nor U7581 (N_7581,N_4542,N_5260);
nor U7582 (N_7582,N_5032,N_4467);
and U7583 (N_7583,N_4596,N_5121);
nor U7584 (N_7584,N_5228,N_4816);
nand U7585 (N_7585,N_4333,N_4604);
nor U7586 (N_7586,N_5137,N_4624);
nand U7587 (N_7587,N_5144,N_4668);
nor U7588 (N_7588,N_5037,N_5347);
nor U7589 (N_7589,N_4563,N_4350);
or U7590 (N_7590,N_4602,N_4307);
or U7591 (N_7591,N_5502,N_4645);
xor U7592 (N_7592,N_5131,N_5156);
nor U7593 (N_7593,N_4370,N_4920);
and U7594 (N_7594,N_5940,N_4948);
nor U7595 (N_7595,N_4100,N_5715);
and U7596 (N_7596,N_5570,N_5108);
or U7597 (N_7597,N_4148,N_4802);
and U7598 (N_7598,N_5835,N_4227);
and U7599 (N_7599,N_4131,N_4807);
nand U7600 (N_7600,N_4311,N_4542);
nand U7601 (N_7601,N_4500,N_5689);
or U7602 (N_7602,N_4915,N_5583);
nand U7603 (N_7603,N_4958,N_5294);
nand U7604 (N_7604,N_5063,N_5772);
and U7605 (N_7605,N_4504,N_5204);
and U7606 (N_7606,N_4047,N_5125);
nor U7607 (N_7607,N_5836,N_4824);
nor U7608 (N_7608,N_5489,N_5186);
nand U7609 (N_7609,N_4786,N_4348);
and U7610 (N_7610,N_4174,N_5153);
xnor U7611 (N_7611,N_4035,N_5621);
nand U7612 (N_7612,N_4521,N_4692);
and U7613 (N_7613,N_4134,N_4086);
and U7614 (N_7614,N_5917,N_4552);
and U7615 (N_7615,N_4885,N_5875);
or U7616 (N_7616,N_4210,N_5629);
xnor U7617 (N_7617,N_5229,N_4169);
nand U7618 (N_7618,N_5042,N_5007);
or U7619 (N_7619,N_4368,N_5957);
nand U7620 (N_7620,N_4391,N_5331);
or U7621 (N_7621,N_5177,N_5521);
nand U7622 (N_7622,N_4659,N_5228);
nor U7623 (N_7623,N_4727,N_4085);
and U7624 (N_7624,N_4190,N_5008);
nand U7625 (N_7625,N_4019,N_4486);
and U7626 (N_7626,N_4993,N_5654);
and U7627 (N_7627,N_4928,N_5429);
and U7628 (N_7628,N_4298,N_5579);
and U7629 (N_7629,N_5082,N_5781);
nand U7630 (N_7630,N_5117,N_5937);
xor U7631 (N_7631,N_4095,N_5271);
nand U7632 (N_7632,N_4064,N_4776);
and U7633 (N_7633,N_4147,N_4806);
nor U7634 (N_7634,N_5474,N_5017);
nand U7635 (N_7635,N_4807,N_4198);
or U7636 (N_7636,N_4988,N_5337);
nor U7637 (N_7637,N_4217,N_4125);
nand U7638 (N_7638,N_4678,N_5839);
nand U7639 (N_7639,N_5905,N_5784);
nor U7640 (N_7640,N_5849,N_5260);
nor U7641 (N_7641,N_5684,N_4469);
nor U7642 (N_7642,N_5114,N_5080);
nor U7643 (N_7643,N_4178,N_5757);
or U7644 (N_7644,N_4517,N_4918);
and U7645 (N_7645,N_4984,N_4265);
nor U7646 (N_7646,N_4827,N_5058);
nor U7647 (N_7647,N_5545,N_4383);
nand U7648 (N_7648,N_5726,N_4748);
and U7649 (N_7649,N_4838,N_4281);
nand U7650 (N_7650,N_4866,N_5617);
nor U7651 (N_7651,N_4753,N_5448);
or U7652 (N_7652,N_5546,N_5959);
nor U7653 (N_7653,N_5487,N_5993);
nor U7654 (N_7654,N_4236,N_4511);
xnor U7655 (N_7655,N_5452,N_4662);
nor U7656 (N_7656,N_4302,N_4769);
and U7657 (N_7657,N_4643,N_4144);
xor U7658 (N_7658,N_5078,N_4987);
and U7659 (N_7659,N_4023,N_4503);
nor U7660 (N_7660,N_4896,N_5292);
nor U7661 (N_7661,N_4006,N_5965);
and U7662 (N_7662,N_4278,N_4990);
nand U7663 (N_7663,N_5888,N_5654);
and U7664 (N_7664,N_4020,N_5371);
or U7665 (N_7665,N_5684,N_5450);
nor U7666 (N_7666,N_4560,N_5367);
nor U7667 (N_7667,N_5930,N_5210);
nand U7668 (N_7668,N_4507,N_4440);
or U7669 (N_7669,N_5233,N_4579);
nor U7670 (N_7670,N_5542,N_5303);
or U7671 (N_7671,N_5596,N_5273);
nor U7672 (N_7672,N_5410,N_5944);
or U7673 (N_7673,N_4294,N_5762);
and U7674 (N_7674,N_4456,N_5716);
xnor U7675 (N_7675,N_4185,N_5535);
and U7676 (N_7676,N_5868,N_5674);
xnor U7677 (N_7677,N_4382,N_4753);
xor U7678 (N_7678,N_5081,N_5257);
or U7679 (N_7679,N_5819,N_4121);
nor U7680 (N_7680,N_4463,N_5369);
nand U7681 (N_7681,N_5260,N_5693);
nor U7682 (N_7682,N_5600,N_4457);
xor U7683 (N_7683,N_5329,N_4407);
nor U7684 (N_7684,N_4033,N_5522);
and U7685 (N_7685,N_5914,N_5342);
or U7686 (N_7686,N_4192,N_4391);
nand U7687 (N_7687,N_4026,N_4202);
nand U7688 (N_7688,N_4469,N_5215);
or U7689 (N_7689,N_4752,N_5462);
xor U7690 (N_7690,N_4399,N_5675);
nor U7691 (N_7691,N_5633,N_4283);
or U7692 (N_7692,N_5213,N_4513);
or U7693 (N_7693,N_4921,N_5560);
or U7694 (N_7694,N_5083,N_4526);
nand U7695 (N_7695,N_5606,N_4244);
xor U7696 (N_7696,N_5646,N_5534);
and U7697 (N_7697,N_4754,N_5743);
and U7698 (N_7698,N_5826,N_5630);
xor U7699 (N_7699,N_5058,N_5801);
and U7700 (N_7700,N_4191,N_5408);
and U7701 (N_7701,N_5414,N_5450);
nand U7702 (N_7702,N_5979,N_5053);
nor U7703 (N_7703,N_5614,N_4030);
or U7704 (N_7704,N_4462,N_5976);
nor U7705 (N_7705,N_5279,N_4384);
nand U7706 (N_7706,N_5297,N_4297);
and U7707 (N_7707,N_5809,N_4501);
xor U7708 (N_7708,N_4889,N_4918);
and U7709 (N_7709,N_5661,N_5816);
or U7710 (N_7710,N_5045,N_4904);
nand U7711 (N_7711,N_5303,N_5608);
or U7712 (N_7712,N_5731,N_5251);
nor U7713 (N_7713,N_4713,N_5396);
or U7714 (N_7714,N_4706,N_4312);
xnor U7715 (N_7715,N_4124,N_4976);
nor U7716 (N_7716,N_5951,N_5777);
nand U7717 (N_7717,N_5666,N_5237);
nor U7718 (N_7718,N_4028,N_4459);
xnor U7719 (N_7719,N_5887,N_5133);
or U7720 (N_7720,N_4043,N_4775);
and U7721 (N_7721,N_4907,N_4332);
nand U7722 (N_7722,N_5145,N_5551);
nand U7723 (N_7723,N_4225,N_4999);
nand U7724 (N_7724,N_4749,N_4278);
or U7725 (N_7725,N_5468,N_4318);
nor U7726 (N_7726,N_4430,N_5266);
or U7727 (N_7727,N_5645,N_4315);
nand U7728 (N_7728,N_5388,N_5423);
nand U7729 (N_7729,N_5442,N_4360);
or U7730 (N_7730,N_4080,N_5366);
and U7731 (N_7731,N_4243,N_4575);
nand U7732 (N_7732,N_4964,N_4294);
nand U7733 (N_7733,N_5572,N_5247);
or U7734 (N_7734,N_4541,N_5287);
nand U7735 (N_7735,N_4273,N_5818);
nand U7736 (N_7736,N_5162,N_4114);
nand U7737 (N_7737,N_5400,N_5984);
and U7738 (N_7738,N_4543,N_5319);
nand U7739 (N_7739,N_4231,N_5910);
and U7740 (N_7740,N_4760,N_4370);
nand U7741 (N_7741,N_4548,N_4759);
and U7742 (N_7742,N_5555,N_5918);
nand U7743 (N_7743,N_4377,N_5379);
and U7744 (N_7744,N_5882,N_5686);
and U7745 (N_7745,N_5521,N_5142);
nor U7746 (N_7746,N_5555,N_5173);
nor U7747 (N_7747,N_4275,N_5963);
and U7748 (N_7748,N_5416,N_5289);
nor U7749 (N_7749,N_4218,N_5229);
nor U7750 (N_7750,N_5615,N_4844);
nor U7751 (N_7751,N_4741,N_5995);
xor U7752 (N_7752,N_4107,N_5502);
nand U7753 (N_7753,N_4771,N_5389);
xnor U7754 (N_7754,N_5228,N_5386);
nand U7755 (N_7755,N_4844,N_5362);
nand U7756 (N_7756,N_5575,N_5433);
or U7757 (N_7757,N_5817,N_5400);
nor U7758 (N_7758,N_5914,N_4804);
nand U7759 (N_7759,N_5637,N_5622);
nor U7760 (N_7760,N_5005,N_5195);
and U7761 (N_7761,N_4363,N_5124);
nor U7762 (N_7762,N_5626,N_4644);
nor U7763 (N_7763,N_5499,N_4281);
nand U7764 (N_7764,N_5093,N_4526);
nor U7765 (N_7765,N_5509,N_4229);
and U7766 (N_7766,N_4178,N_4744);
nor U7767 (N_7767,N_5280,N_5744);
or U7768 (N_7768,N_5868,N_4750);
and U7769 (N_7769,N_5346,N_5240);
and U7770 (N_7770,N_5103,N_5220);
nand U7771 (N_7771,N_4638,N_5611);
nor U7772 (N_7772,N_4405,N_4307);
nor U7773 (N_7773,N_4330,N_4556);
nor U7774 (N_7774,N_5636,N_4779);
and U7775 (N_7775,N_4821,N_4992);
xor U7776 (N_7776,N_5279,N_5693);
and U7777 (N_7777,N_4693,N_5285);
and U7778 (N_7778,N_4728,N_4651);
or U7779 (N_7779,N_4014,N_4030);
and U7780 (N_7780,N_5454,N_4024);
or U7781 (N_7781,N_4174,N_4999);
and U7782 (N_7782,N_5459,N_5244);
and U7783 (N_7783,N_5268,N_4373);
nand U7784 (N_7784,N_5009,N_4591);
or U7785 (N_7785,N_5962,N_5805);
nand U7786 (N_7786,N_5165,N_4185);
nor U7787 (N_7787,N_5841,N_4990);
and U7788 (N_7788,N_4771,N_5171);
or U7789 (N_7789,N_5979,N_4720);
or U7790 (N_7790,N_4257,N_5511);
nor U7791 (N_7791,N_4929,N_5184);
or U7792 (N_7792,N_4318,N_5906);
nand U7793 (N_7793,N_5553,N_4063);
nand U7794 (N_7794,N_5799,N_4015);
xnor U7795 (N_7795,N_4656,N_4552);
nand U7796 (N_7796,N_5590,N_4619);
nor U7797 (N_7797,N_4024,N_5333);
and U7798 (N_7798,N_5301,N_4664);
or U7799 (N_7799,N_4020,N_4692);
or U7800 (N_7800,N_5146,N_4232);
nand U7801 (N_7801,N_5940,N_5064);
or U7802 (N_7802,N_4580,N_5006);
or U7803 (N_7803,N_5736,N_4675);
nand U7804 (N_7804,N_5538,N_5257);
nand U7805 (N_7805,N_4157,N_5520);
and U7806 (N_7806,N_4337,N_4214);
xnor U7807 (N_7807,N_4993,N_5087);
nor U7808 (N_7808,N_4136,N_4886);
or U7809 (N_7809,N_5572,N_5974);
nor U7810 (N_7810,N_5783,N_5355);
nor U7811 (N_7811,N_5002,N_4570);
or U7812 (N_7812,N_4356,N_4419);
nand U7813 (N_7813,N_4177,N_4801);
xor U7814 (N_7814,N_5937,N_5582);
nand U7815 (N_7815,N_4981,N_5807);
xnor U7816 (N_7816,N_4051,N_4023);
or U7817 (N_7817,N_5050,N_4811);
or U7818 (N_7818,N_4611,N_4252);
and U7819 (N_7819,N_5096,N_5840);
nand U7820 (N_7820,N_4016,N_4559);
nor U7821 (N_7821,N_4505,N_5695);
and U7822 (N_7822,N_5483,N_5437);
nand U7823 (N_7823,N_4514,N_4449);
and U7824 (N_7824,N_5008,N_4215);
nor U7825 (N_7825,N_4136,N_5693);
nand U7826 (N_7826,N_5218,N_5262);
and U7827 (N_7827,N_5581,N_4711);
nor U7828 (N_7828,N_4058,N_4367);
and U7829 (N_7829,N_5442,N_4896);
nand U7830 (N_7830,N_5595,N_5243);
xor U7831 (N_7831,N_5426,N_5552);
and U7832 (N_7832,N_5824,N_4736);
or U7833 (N_7833,N_5030,N_4495);
and U7834 (N_7834,N_4406,N_5704);
xnor U7835 (N_7835,N_4739,N_4401);
nor U7836 (N_7836,N_4831,N_5220);
and U7837 (N_7837,N_4360,N_5928);
xnor U7838 (N_7838,N_5231,N_5192);
nand U7839 (N_7839,N_4636,N_4887);
nor U7840 (N_7840,N_4388,N_4334);
nand U7841 (N_7841,N_5710,N_4833);
nand U7842 (N_7842,N_4970,N_4572);
nand U7843 (N_7843,N_5053,N_4503);
xnor U7844 (N_7844,N_4170,N_4177);
nand U7845 (N_7845,N_5167,N_5017);
xor U7846 (N_7846,N_5197,N_4532);
or U7847 (N_7847,N_4769,N_4394);
or U7848 (N_7848,N_4476,N_5317);
or U7849 (N_7849,N_5577,N_5319);
xnor U7850 (N_7850,N_5329,N_4862);
or U7851 (N_7851,N_4006,N_4323);
or U7852 (N_7852,N_4553,N_5056);
xor U7853 (N_7853,N_4768,N_5916);
nor U7854 (N_7854,N_4311,N_5309);
and U7855 (N_7855,N_5688,N_4537);
xor U7856 (N_7856,N_4357,N_4974);
nor U7857 (N_7857,N_5258,N_5741);
and U7858 (N_7858,N_5248,N_5571);
nor U7859 (N_7859,N_5108,N_5957);
nand U7860 (N_7860,N_5032,N_4257);
nand U7861 (N_7861,N_4723,N_5621);
or U7862 (N_7862,N_4241,N_4292);
and U7863 (N_7863,N_4122,N_4441);
or U7864 (N_7864,N_5151,N_4411);
nand U7865 (N_7865,N_4015,N_4421);
nand U7866 (N_7866,N_4498,N_4118);
xnor U7867 (N_7867,N_5914,N_5074);
nand U7868 (N_7868,N_4873,N_4043);
or U7869 (N_7869,N_4652,N_5751);
and U7870 (N_7870,N_5478,N_4800);
or U7871 (N_7871,N_5782,N_5275);
and U7872 (N_7872,N_5172,N_5446);
xor U7873 (N_7873,N_4888,N_5978);
nor U7874 (N_7874,N_4790,N_4612);
nand U7875 (N_7875,N_4101,N_5047);
nor U7876 (N_7876,N_5965,N_4913);
nand U7877 (N_7877,N_4245,N_4731);
xor U7878 (N_7878,N_5430,N_5049);
nand U7879 (N_7879,N_5237,N_4523);
nor U7880 (N_7880,N_5491,N_5483);
nor U7881 (N_7881,N_5571,N_4210);
or U7882 (N_7882,N_5705,N_5210);
and U7883 (N_7883,N_5217,N_4562);
nor U7884 (N_7884,N_4632,N_4317);
nor U7885 (N_7885,N_4294,N_5591);
and U7886 (N_7886,N_5513,N_5611);
or U7887 (N_7887,N_4678,N_5063);
or U7888 (N_7888,N_5770,N_4161);
nand U7889 (N_7889,N_4896,N_4862);
or U7890 (N_7890,N_5530,N_4780);
nor U7891 (N_7891,N_4171,N_5886);
nand U7892 (N_7892,N_4728,N_4319);
nor U7893 (N_7893,N_5912,N_5419);
nand U7894 (N_7894,N_4754,N_5991);
nand U7895 (N_7895,N_4181,N_5605);
nand U7896 (N_7896,N_4187,N_5751);
or U7897 (N_7897,N_4616,N_4338);
or U7898 (N_7898,N_5148,N_4358);
nand U7899 (N_7899,N_5419,N_4963);
nor U7900 (N_7900,N_4699,N_5227);
and U7901 (N_7901,N_4491,N_5150);
nor U7902 (N_7902,N_4973,N_5153);
and U7903 (N_7903,N_4641,N_5720);
or U7904 (N_7904,N_5607,N_4075);
and U7905 (N_7905,N_5708,N_4279);
or U7906 (N_7906,N_4620,N_5386);
nand U7907 (N_7907,N_5056,N_5823);
and U7908 (N_7908,N_5578,N_5832);
nor U7909 (N_7909,N_4994,N_4980);
or U7910 (N_7910,N_5130,N_4019);
nand U7911 (N_7911,N_5967,N_5909);
xnor U7912 (N_7912,N_4341,N_5911);
nor U7913 (N_7913,N_5238,N_5442);
or U7914 (N_7914,N_5367,N_4687);
and U7915 (N_7915,N_5735,N_4592);
and U7916 (N_7916,N_4440,N_5616);
or U7917 (N_7917,N_5869,N_4723);
or U7918 (N_7918,N_4413,N_4431);
or U7919 (N_7919,N_5660,N_4015);
nand U7920 (N_7920,N_5125,N_5576);
or U7921 (N_7921,N_4111,N_4198);
xor U7922 (N_7922,N_5480,N_4943);
nand U7923 (N_7923,N_5744,N_5424);
and U7924 (N_7924,N_4141,N_5824);
nor U7925 (N_7925,N_4012,N_5630);
nand U7926 (N_7926,N_4258,N_4262);
or U7927 (N_7927,N_4602,N_4440);
or U7928 (N_7928,N_5217,N_4343);
or U7929 (N_7929,N_5225,N_4093);
nor U7930 (N_7930,N_4844,N_5655);
nor U7931 (N_7931,N_4324,N_4458);
or U7932 (N_7932,N_5826,N_4083);
nor U7933 (N_7933,N_4111,N_5264);
or U7934 (N_7934,N_4413,N_4601);
nor U7935 (N_7935,N_4968,N_5845);
and U7936 (N_7936,N_4721,N_5103);
nand U7937 (N_7937,N_5731,N_4465);
nand U7938 (N_7938,N_4487,N_5411);
nor U7939 (N_7939,N_5957,N_4663);
nand U7940 (N_7940,N_5633,N_4440);
nand U7941 (N_7941,N_4125,N_5273);
nor U7942 (N_7942,N_5932,N_4268);
or U7943 (N_7943,N_5157,N_5365);
or U7944 (N_7944,N_5816,N_4171);
nand U7945 (N_7945,N_5719,N_4023);
and U7946 (N_7946,N_5639,N_5846);
or U7947 (N_7947,N_5924,N_4909);
nor U7948 (N_7948,N_5697,N_5584);
and U7949 (N_7949,N_5702,N_4527);
and U7950 (N_7950,N_4499,N_4736);
nand U7951 (N_7951,N_4682,N_4203);
or U7952 (N_7952,N_5354,N_5193);
nor U7953 (N_7953,N_5928,N_5222);
nand U7954 (N_7954,N_5966,N_5999);
nor U7955 (N_7955,N_5972,N_5797);
nor U7956 (N_7956,N_4412,N_5410);
and U7957 (N_7957,N_5175,N_5426);
nand U7958 (N_7958,N_4102,N_4945);
and U7959 (N_7959,N_5137,N_5060);
or U7960 (N_7960,N_5561,N_5786);
and U7961 (N_7961,N_5665,N_4620);
or U7962 (N_7962,N_4037,N_5111);
or U7963 (N_7963,N_5934,N_4768);
and U7964 (N_7964,N_4097,N_5148);
nor U7965 (N_7965,N_4284,N_5101);
nor U7966 (N_7966,N_4226,N_5852);
nor U7967 (N_7967,N_5183,N_5345);
and U7968 (N_7968,N_4650,N_4150);
or U7969 (N_7969,N_4866,N_4567);
xnor U7970 (N_7970,N_5899,N_5526);
nand U7971 (N_7971,N_4828,N_4054);
nor U7972 (N_7972,N_4544,N_4211);
nor U7973 (N_7973,N_4960,N_5669);
or U7974 (N_7974,N_5358,N_5627);
or U7975 (N_7975,N_5503,N_5378);
nor U7976 (N_7976,N_4857,N_5121);
nand U7977 (N_7977,N_5696,N_4009);
xor U7978 (N_7978,N_4237,N_4378);
nand U7979 (N_7979,N_4167,N_5251);
nor U7980 (N_7980,N_5478,N_5066);
and U7981 (N_7981,N_4651,N_4993);
or U7982 (N_7982,N_4955,N_4822);
nand U7983 (N_7983,N_4157,N_5411);
and U7984 (N_7984,N_5154,N_5714);
xnor U7985 (N_7985,N_4146,N_4516);
and U7986 (N_7986,N_4379,N_4562);
nand U7987 (N_7987,N_5736,N_4599);
nand U7988 (N_7988,N_5699,N_4146);
and U7989 (N_7989,N_4279,N_5062);
and U7990 (N_7990,N_5733,N_4690);
xor U7991 (N_7991,N_4563,N_4032);
and U7992 (N_7992,N_4441,N_5761);
xnor U7993 (N_7993,N_5568,N_5992);
and U7994 (N_7994,N_5861,N_4436);
or U7995 (N_7995,N_4518,N_5091);
nand U7996 (N_7996,N_5372,N_4282);
xor U7997 (N_7997,N_4493,N_4460);
nand U7998 (N_7998,N_4561,N_4705);
nor U7999 (N_7999,N_4487,N_4908);
nand U8000 (N_8000,N_6643,N_7554);
or U8001 (N_8001,N_6330,N_6768);
xor U8002 (N_8002,N_6020,N_6389);
xor U8003 (N_8003,N_6195,N_6023);
and U8004 (N_8004,N_6361,N_6858);
and U8005 (N_8005,N_6052,N_7084);
nor U8006 (N_8006,N_6497,N_6337);
or U8007 (N_8007,N_6840,N_7990);
and U8008 (N_8008,N_6019,N_7630);
nor U8009 (N_8009,N_6568,N_7137);
and U8010 (N_8010,N_6945,N_6825);
or U8011 (N_8011,N_7668,N_6594);
nor U8012 (N_8012,N_7740,N_7949);
nor U8013 (N_8013,N_6249,N_7984);
or U8014 (N_8014,N_7366,N_7970);
xnor U8015 (N_8015,N_7000,N_6327);
or U8016 (N_8016,N_7491,N_6662);
nor U8017 (N_8017,N_6095,N_7169);
nor U8018 (N_8018,N_7284,N_6364);
or U8019 (N_8019,N_7188,N_7475);
and U8020 (N_8020,N_7149,N_6414);
nor U8021 (N_8021,N_7427,N_6002);
and U8022 (N_8022,N_7125,N_6494);
nor U8023 (N_8023,N_7869,N_7547);
or U8024 (N_8024,N_7297,N_6715);
xor U8025 (N_8025,N_7868,N_6388);
or U8026 (N_8026,N_6678,N_7627);
nand U8027 (N_8027,N_6233,N_7150);
nand U8028 (N_8028,N_7811,N_6882);
and U8029 (N_8029,N_7660,N_6823);
nand U8030 (N_8030,N_6991,N_7457);
nor U8031 (N_8031,N_7005,N_6055);
xnor U8032 (N_8032,N_7294,N_6036);
nand U8033 (N_8033,N_7160,N_6001);
and U8034 (N_8034,N_7363,N_6629);
nor U8035 (N_8035,N_7670,N_7336);
xor U8036 (N_8036,N_7575,N_6656);
nand U8037 (N_8037,N_7099,N_6919);
or U8038 (N_8038,N_6419,N_7656);
and U8039 (N_8039,N_7742,N_6783);
or U8040 (N_8040,N_6852,N_7770);
or U8041 (N_8041,N_7771,N_7796);
nor U8042 (N_8042,N_6903,N_6582);
or U8043 (N_8043,N_6863,N_6659);
nand U8044 (N_8044,N_7092,N_6561);
or U8045 (N_8045,N_7305,N_6123);
nor U8046 (N_8046,N_6965,N_7584);
and U8047 (N_8047,N_7975,N_7790);
and U8048 (N_8048,N_6299,N_7748);
and U8049 (N_8049,N_7763,N_6218);
xnor U8050 (N_8050,N_6304,N_6203);
and U8051 (N_8051,N_7911,N_7227);
and U8052 (N_8052,N_7918,N_6705);
or U8053 (N_8053,N_6560,N_6745);
nor U8054 (N_8054,N_7064,N_6131);
xnor U8055 (N_8055,N_7808,N_7541);
and U8056 (N_8056,N_6596,N_6246);
xnor U8057 (N_8057,N_6722,N_7538);
and U8058 (N_8058,N_6275,N_7794);
nand U8059 (N_8059,N_7906,N_6577);
nand U8060 (N_8060,N_7060,N_6378);
nand U8061 (N_8061,N_6365,N_6737);
xnor U8062 (N_8062,N_6581,N_7513);
and U8063 (N_8063,N_6828,N_6819);
nor U8064 (N_8064,N_6812,N_7940);
xnor U8065 (N_8065,N_7304,N_7420);
and U8066 (N_8066,N_6326,N_6433);
and U8067 (N_8067,N_6752,N_6790);
or U8068 (N_8068,N_7819,N_6871);
nand U8069 (N_8069,N_6704,N_7737);
or U8070 (N_8070,N_7610,N_7686);
nor U8071 (N_8071,N_6401,N_6422);
and U8072 (N_8072,N_6210,N_7499);
and U8073 (N_8073,N_7874,N_7919);
nor U8074 (N_8074,N_6073,N_7365);
or U8075 (N_8075,N_7553,N_7082);
or U8076 (N_8076,N_6572,N_6487);
or U8077 (N_8077,N_6022,N_6830);
or U8078 (N_8078,N_6845,N_7027);
nor U8079 (N_8079,N_7521,N_7494);
nand U8080 (N_8080,N_7841,N_7502);
and U8081 (N_8081,N_6405,N_6846);
nand U8082 (N_8082,N_6839,N_6350);
and U8083 (N_8083,N_7145,N_6847);
nand U8084 (N_8084,N_7981,N_7661);
nor U8085 (N_8085,N_7389,N_6804);
or U8086 (N_8086,N_7102,N_6503);
or U8087 (N_8087,N_6007,N_7489);
nand U8088 (N_8088,N_6089,N_6535);
or U8089 (N_8089,N_7681,N_6385);
and U8090 (N_8090,N_6734,N_7194);
nor U8091 (N_8091,N_7865,N_6394);
or U8092 (N_8092,N_7533,N_6966);
and U8093 (N_8093,N_6543,N_6941);
nor U8094 (N_8094,N_6802,N_7016);
or U8095 (N_8095,N_6763,N_6976);
or U8096 (N_8096,N_6532,N_7514);
nand U8097 (N_8097,N_7658,N_6094);
nor U8098 (N_8098,N_7409,N_6933);
xor U8099 (N_8099,N_6910,N_7382);
or U8100 (N_8100,N_6428,N_6829);
nor U8101 (N_8101,N_7311,N_6256);
or U8102 (N_8102,N_6066,N_6436);
nor U8103 (N_8103,N_6196,N_7707);
nand U8104 (N_8104,N_6603,N_7685);
and U8105 (N_8105,N_7912,N_7876);
and U8106 (N_8106,N_6669,N_7801);
and U8107 (N_8107,N_6794,N_7348);
and U8108 (N_8108,N_7379,N_7065);
nand U8109 (N_8109,N_7856,N_6619);
nand U8110 (N_8110,N_6542,N_7993);
xnor U8111 (N_8111,N_7959,N_7019);
and U8112 (N_8112,N_7262,N_7378);
nor U8113 (N_8113,N_7580,N_7086);
nand U8114 (N_8114,N_7684,N_6167);
nand U8115 (N_8115,N_7530,N_7044);
nor U8116 (N_8116,N_6390,N_6711);
and U8117 (N_8117,N_6041,N_6979);
or U8118 (N_8118,N_6479,N_7370);
nand U8119 (N_8119,N_7059,N_7923);
and U8120 (N_8120,N_6575,N_6174);
and U8121 (N_8121,N_7645,N_6043);
nor U8122 (N_8122,N_6311,N_7051);
nand U8123 (N_8123,N_6569,N_7980);
xor U8124 (N_8124,N_7511,N_6694);
nand U8125 (N_8125,N_6455,N_6145);
and U8126 (N_8126,N_6538,N_7750);
xnor U8127 (N_8127,N_7663,N_7280);
nand U8128 (N_8128,N_7814,N_6730);
or U8129 (N_8129,N_7377,N_7972);
xor U8130 (N_8130,N_7723,N_6680);
nor U8131 (N_8131,N_7098,N_7447);
xnor U8132 (N_8132,N_6254,N_7076);
nand U8133 (N_8133,N_6975,N_7560);
and U8134 (N_8134,N_6972,N_7900);
nand U8135 (N_8135,N_7053,N_7855);
nand U8136 (N_8136,N_7877,N_7013);
nand U8137 (N_8137,N_6236,N_7916);
nor U8138 (N_8138,N_7588,N_6736);
or U8139 (N_8139,N_6039,N_7569);
or U8140 (N_8140,N_6584,N_6376);
nand U8141 (N_8141,N_7667,N_7581);
xnor U8142 (N_8142,N_7958,N_6449);
nor U8143 (N_8143,N_6929,N_6398);
nor U8144 (N_8144,N_7821,N_7628);
nand U8145 (N_8145,N_6521,N_6059);
or U8146 (N_8146,N_7552,N_6166);
nand U8147 (N_8147,N_7589,N_7515);
xnor U8148 (N_8148,N_7831,N_7122);
and U8149 (N_8149,N_7785,N_7844);
nand U8150 (N_8150,N_6585,N_6461);
and U8151 (N_8151,N_7709,N_6178);
nand U8152 (N_8152,N_7110,N_7342);
nand U8153 (N_8153,N_7741,N_7134);
or U8154 (N_8154,N_6237,N_7969);
nor U8155 (N_8155,N_7903,N_7593);
and U8156 (N_8156,N_7410,N_7647);
nor U8157 (N_8157,N_6641,N_7526);
nor U8158 (N_8158,N_7724,N_6772);
nand U8159 (N_8159,N_7252,N_6402);
nand U8160 (N_8160,N_7505,N_6344);
nor U8161 (N_8161,N_6587,N_6363);
and U8162 (N_8162,N_7755,N_6064);
or U8163 (N_8163,N_6030,N_7894);
nor U8164 (N_8164,N_7132,N_7600);
nor U8165 (N_8165,N_6320,N_7784);
nand U8166 (N_8166,N_6093,N_6848);
or U8167 (N_8167,N_6477,N_7226);
nand U8168 (N_8168,N_6668,N_7299);
and U8169 (N_8169,N_6129,N_6435);
and U8170 (N_8170,N_6597,N_7185);
and U8171 (N_8171,N_7253,N_7343);
nor U8172 (N_8172,N_7640,N_6396);
nor U8173 (N_8173,N_6690,N_7007);
and U8174 (N_8174,N_7333,N_7786);
and U8175 (N_8175,N_6683,N_7107);
and U8176 (N_8176,N_6645,N_7706);
and U8177 (N_8177,N_7069,N_6761);
nand U8178 (N_8178,N_7196,N_7544);
nor U8179 (N_8179,N_7921,N_6011);
and U8180 (N_8180,N_6334,N_7485);
or U8181 (N_8181,N_6138,N_6489);
nand U8182 (N_8182,N_6673,N_7144);
and U8183 (N_8183,N_7701,N_6159);
and U8184 (N_8184,N_7947,N_6609);
nor U8185 (N_8185,N_6938,N_6540);
nor U8186 (N_8186,N_6434,N_7096);
or U8187 (N_8187,N_6693,N_7536);
and U8188 (N_8188,N_6671,N_6931);
nand U8189 (N_8189,N_7840,N_6546);
and U8190 (N_8190,N_7837,N_6054);
and U8191 (N_8191,N_6885,N_6674);
nand U8192 (N_8192,N_7392,N_7967);
or U8193 (N_8193,N_6120,N_7331);
and U8194 (N_8194,N_7133,N_6226);
or U8195 (N_8195,N_6689,N_6756);
or U8196 (N_8196,N_6815,N_7866);
xnor U8197 (N_8197,N_7384,N_6317);
nand U8198 (N_8198,N_7130,N_6646);
nor U8199 (N_8199,N_7435,N_7142);
xnor U8200 (N_8200,N_7999,N_6040);
nor U8201 (N_8201,N_7985,N_6035);
or U8202 (N_8202,N_7117,N_7173);
nand U8203 (N_8203,N_6420,N_7424);
xor U8204 (N_8204,N_7079,N_6295);
nor U8205 (N_8205,N_7849,N_6124);
nor U8206 (N_8206,N_6670,N_7622);
nor U8207 (N_8207,N_7804,N_7633);
nor U8208 (N_8208,N_7049,N_6085);
or U8209 (N_8209,N_7001,N_7345);
nor U8210 (N_8210,N_6198,N_6925);
nor U8211 (N_8211,N_6250,N_6961);
and U8212 (N_8212,N_7792,N_7854);
or U8213 (N_8213,N_6024,N_7250);
nor U8214 (N_8214,N_7915,N_7004);
nand U8215 (N_8215,N_6352,N_6343);
nand U8216 (N_8216,N_6312,N_7545);
and U8217 (N_8217,N_7634,N_6453);
and U8218 (N_8218,N_7863,N_7994);
xnor U8219 (N_8219,N_7644,N_6551);
or U8220 (N_8220,N_7490,N_7308);
and U8221 (N_8221,N_7467,N_6215);
nor U8222 (N_8222,N_7401,N_6512);
nor U8223 (N_8223,N_6700,N_6285);
nor U8224 (N_8224,N_7022,N_7797);
nand U8225 (N_8225,N_7291,N_6962);
nand U8226 (N_8226,N_7687,N_6245);
nor U8227 (N_8227,N_7057,N_7592);
or U8228 (N_8228,N_7042,N_7503);
and U8229 (N_8229,N_7517,N_6744);
or U8230 (N_8230,N_7765,N_7455);
or U8231 (N_8231,N_7432,N_6316);
nor U8232 (N_8232,N_7310,N_7599);
and U8233 (N_8233,N_7011,N_7577);
nor U8234 (N_8234,N_6213,N_7812);
nand U8235 (N_8235,N_6781,N_6757);
nand U8236 (N_8236,N_6786,N_7974);
nor U8237 (N_8237,N_7285,N_6563);
nand U8238 (N_8238,N_7810,N_6545);
nand U8239 (N_8239,N_7193,N_6881);
and U8240 (N_8240,N_7359,N_7951);
nand U8241 (N_8241,N_6163,N_6305);
and U8242 (N_8242,N_7871,N_7408);
nand U8243 (N_8243,N_6319,N_6746);
or U8244 (N_8244,N_7167,N_6873);
nor U8245 (N_8245,N_6411,N_7726);
and U8246 (N_8246,N_6475,N_6292);
nor U8247 (N_8247,N_6519,N_6194);
nor U8248 (N_8248,N_6654,N_7809);
or U8249 (N_8249,N_6142,N_6854);
xor U8250 (N_8250,N_7071,N_6676);
nand U8251 (N_8251,N_6286,N_7988);
nor U8252 (N_8252,N_7946,N_7442);
and U8253 (N_8253,N_6620,N_7418);
xor U8254 (N_8254,N_7463,N_6336);
nor U8255 (N_8255,N_6549,N_6894);
xor U8256 (N_8256,N_7220,N_6952);
xor U8257 (N_8257,N_6905,N_6706);
and U8258 (N_8258,N_6958,N_7452);
nand U8259 (N_8259,N_7830,N_6895);
nor U8260 (N_8260,N_7971,N_7507);
nand U8261 (N_8261,N_6306,N_6119);
nor U8262 (N_8262,N_7230,N_6807);
nor U8263 (N_8263,N_7965,N_7884);
nand U8264 (N_8264,N_6809,N_6907);
and U8265 (N_8265,N_6998,N_7459);
nor U8266 (N_8266,N_7638,N_6004);
or U8267 (N_8267,N_7651,N_7269);
nand U8268 (N_8268,N_6014,N_7183);
xnor U8269 (N_8269,N_7825,N_7932);
or U8270 (N_8270,N_6239,N_7757);
nor U8271 (N_8271,N_7391,N_7646);
xor U8272 (N_8272,N_6988,N_7035);
xor U8273 (N_8273,N_7032,N_6273);
xor U8274 (N_8274,N_7629,N_6835);
nor U8275 (N_8275,N_6759,N_6155);
nor U8276 (N_8276,N_7565,N_6633);
xnor U8277 (N_8277,N_6499,N_6180);
and U8278 (N_8278,N_7497,N_7721);
nor U8279 (N_8279,N_6114,N_7428);
nor U8280 (N_8280,N_7157,N_7556);
or U8281 (N_8281,N_7104,N_7669);
or U8282 (N_8282,N_7211,N_7327);
xnor U8283 (N_8283,N_7174,N_7488);
and U8284 (N_8284,N_6484,N_6622);
nor U8285 (N_8285,N_6156,N_7606);
and U8286 (N_8286,N_7023,N_7649);
or U8287 (N_8287,N_7760,N_6010);
and U8288 (N_8288,N_7931,N_6170);
or U8289 (N_8289,N_7303,N_7690);
nor U8290 (N_8290,N_7052,N_7198);
nand U8291 (N_8291,N_7067,N_6780);
nor U8292 (N_8292,N_6764,N_6520);
or U8293 (N_8293,N_6212,N_6501);
nor U8294 (N_8294,N_7689,N_6602);
and U8295 (N_8295,N_6369,N_6686);
and U8296 (N_8296,N_6732,N_6099);
and U8297 (N_8297,N_7776,N_7465);
and U8298 (N_8298,N_7462,N_6778);
and U8299 (N_8299,N_6314,N_7140);
nand U8300 (N_8300,N_7539,N_7436);
nand U8301 (N_8301,N_6407,N_6758);
and U8302 (N_8302,N_7329,N_6109);
nand U8303 (N_8303,N_6032,N_6787);
or U8304 (N_8304,N_6438,N_6088);
nand U8305 (N_8305,N_7917,N_7268);
nor U8306 (N_8306,N_6935,N_7857);
and U8307 (N_8307,N_6760,N_7882);
or U8308 (N_8308,N_7914,N_7908);
and U8309 (N_8309,N_7500,N_7322);
or U8310 (N_8310,N_6855,N_6348);
nor U8311 (N_8311,N_6749,N_7012);
or U8312 (N_8312,N_6221,N_6324);
nand U8313 (N_8313,N_7131,N_6162);
or U8314 (N_8314,N_6614,N_6898);
nor U8315 (N_8315,N_7480,N_7003);
nor U8316 (N_8316,N_6849,N_7901);
and U8317 (N_8317,N_7422,N_6644);
and U8318 (N_8318,N_6607,N_6647);
and U8319 (N_8319,N_6943,N_7800);
nand U8320 (N_8320,N_6315,N_7278);
nor U8321 (N_8321,N_7529,N_6591);
nor U8322 (N_8322,N_6726,N_6775);
nand U8323 (N_8323,N_6627,N_7263);
nand U8324 (N_8324,N_7264,N_7828);
or U8325 (N_8325,N_6151,N_7184);
nand U8326 (N_8326,N_6813,N_6038);
and U8327 (N_8327,N_7506,N_7778);
or U8328 (N_8328,N_6130,N_7653);
or U8329 (N_8329,N_7910,N_7703);
or U8330 (N_8330,N_7314,N_7761);
nand U8331 (N_8331,N_6485,N_7405);
and U8332 (N_8332,N_7880,N_6467);
nand U8333 (N_8333,N_6949,N_6168);
nor U8334 (N_8334,N_7292,N_7139);
xor U8335 (N_8335,N_7558,N_6608);
nand U8336 (N_8336,N_7473,N_7213);
nor U8337 (N_8337,N_7254,N_7164);
or U8338 (N_8338,N_7026,N_7306);
or U8339 (N_8339,N_6228,N_6510);
xor U8340 (N_8340,N_7361,N_6559);
nand U8341 (N_8341,N_6974,N_6403);
or U8342 (N_8342,N_6912,N_6639);
nand U8343 (N_8343,N_6526,N_6631);
nand U8344 (N_8344,N_7017,N_6103);
nor U8345 (N_8345,N_6824,N_6444);
and U8346 (N_8346,N_7534,N_6611);
or U8347 (N_8347,N_6956,N_7241);
or U8348 (N_8348,N_6567,N_7815);
or U8349 (N_8349,N_6719,N_6838);
nor U8350 (N_8350,N_6000,N_7037);
nand U8351 (N_8351,N_7381,N_7735);
nor U8352 (N_8352,N_6527,N_6735);
or U8353 (N_8353,N_7477,N_6899);
nand U8354 (N_8354,N_6748,N_7624);
and U8355 (N_8355,N_6459,N_6031);
and U8356 (N_8356,N_7199,N_7460);
nor U8357 (N_8357,N_6214,N_7380);
or U8358 (N_8358,N_6413,N_6183);
nor U8359 (N_8359,N_6377,N_7347);
and U8360 (N_8360,N_7504,N_7586);
nor U8361 (N_8361,N_6235,N_7952);
and U8362 (N_8362,N_7591,N_7728);
nor U8363 (N_8363,N_6294,N_7862);
xor U8364 (N_8364,N_6950,N_6939);
xor U8365 (N_8365,N_7267,N_7070);
nor U8366 (N_8366,N_7838,N_7597);
nand U8367 (N_8367,N_6983,N_6296);
nand U8368 (N_8368,N_6963,N_7151);
nor U8369 (N_8369,N_6500,N_7373);
xor U8370 (N_8370,N_7764,N_7434);
or U8371 (N_8371,N_6147,N_6200);
xnor U8372 (N_8372,N_6960,N_7714);
or U8373 (N_8373,N_7478,N_6297);
and U8374 (N_8374,N_6465,N_7368);
and U8375 (N_8375,N_7788,N_7056);
nor U8376 (N_8376,N_7858,N_7813);
nand U8377 (N_8377,N_6859,N_7271);
and U8378 (N_8378,N_6716,N_6134);
and U8379 (N_8379,N_6383,N_6086);
nor U8380 (N_8380,N_7889,N_7482);
or U8381 (N_8381,N_6204,N_7341);
and U8382 (N_8382,N_7124,N_6776);
nand U8383 (N_8383,N_6853,N_7043);
and U8384 (N_8384,N_7989,N_7907);
and U8385 (N_8385,N_7870,N_6518);
and U8386 (N_8386,N_6707,N_7009);
and U8387 (N_8387,N_6102,N_6217);
nor U8388 (N_8388,N_6851,N_7734);
nand U8389 (N_8389,N_7977,N_7176);
nand U8390 (N_8390,N_6068,N_7697);
or U8391 (N_8391,N_6069,N_7416);
nor U8392 (N_8392,N_7228,N_7672);
or U8393 (N_8393,N_7054,N_6968);
or U8394 (N_8394,N_6954,N_6137);
and U8395 (N_8395,N_6588,N_7369);
and U8396 (N_8396,N_7316,N_6999);
nor U8397 (N_8397,N_6892,N_7062);
or U8398 (N_8398,N_7073,N_7829);
or U8399 (N_8399,N_7845,N_7641);
and U8400 (N_8400,N_6058,N_7326);
or U8401 (N_8401,N_7571,N_6626);
and U8402 (N_8402,N_6349,N_6112);
nor U8403 (N_8403,N_6589,N_6917);
nand U8404 (N_8404,N_7986,N_7626);
and U8405 (N_8405,N_7398,N_7887);
nand U8406 (N_8406,N_7093,N_6682);
nor U8407 (N_8407,N_7293,N_7146);
or U8408 (N_8408,N_6471,N_6874);
and U8409 (N_8409,N_6747,N_7564);
nor U8410 (N_8410,N_7758,N_6883);
and U8411 (N_8411,N_7312,N_6578);
or U8412 (N_8412,N_6583,N_6805);
or U8413 (N_8413,N_6490,N_7330);
nor U8414 (N_8414,N_6878,N_6082);
or U8415 (N_8415,N_6439,N_7864);
xnor U8416 (N_8416,N_7242,N_7962);
and U8417 (N_8417,N_6667,N_7791);
nor U8418 (N_8418,N_6720,N_7083);
nor U8419 (N_8419,N_6046,N_6995);
nor U8420 (N_8420,N_7002,N_6291);
nand U8421 (N_8421,N_6247,N_7590);
xor U8422 (N_8422,N_6021,N_6118);
or U8423 (N_8423,N_7578,N_7927);
and U8424 (N_8424,N_6071,N_6908);
nor U8425 (N_8425,N_6739,N_7153);
xnor U8426 (N_8426,N_7454,N_6751);
nor U8427 (N_8427,N_6712,N_7354);
or U8428 (N_8428,N_7444,N_6049);
and U8429 (N_8429,N_6785,N_7818);
nand U8430 (N_8430,N_7030,N_6552);
nand U8431 (N_8431,N_7563,N_6081);
xnor U8432 (N_8432,N_6857,N_7978);
nand U8433 (N_8433,N_6901,N_6460);
nor U8434 (N_8434,N_7387,N_7729);
nor U8435 (N_8435,N_6301,N_6817);
nand U8436 (N_8436,N_6981,N_7938);
or U8437 (N_8437,N_6013,N_6604);
nand U8438 (N_8438,N_6679,N_6865);
and U8439 (N_8439,N_7548,N_7441);
or U8440 (N_8440,N_7835,N_6877);
nor U8441 (N_8441,N_7966,N_6491);
nor U8442 (N_8442,N_6753,N_6157);
xnor U8443 (N_8443,N_7650,N_7913);
nand U8444 (N_8444,N_6985,N_6224);
nand U8445 (N_8445,N_6573,N_7437);
and U8446 (N_8446,N_6870,N_6179);
or U8447 (N_8447,N_7014,N_6920);
and U8448 (N_8448,N_6153,N_7234);
nand U8449 (N_8449,N_7820,N_7525);
or U8450 (N_8450,N_7702,N_6922);
nor U8451 (N_8451,N_6408,N_7483);
xor U8452 (N_8452,N_7806,N_6474);
nand U8453 (N_8453,N_7450,N_7487);
nor U8454 (N_8454,N_7246,N_7161);
nor U8455 (N_8455,N_7983,N_6406);
or U8456 (N_8456,N_6713,N_6132);
nor U8457 (N_8457,N_6996,N_6658);
xor U8458 (N_8458,N_7128,N_6393);
or U8459 (N_8459,N_6513,N_6127);
nand U8460 (N_8460,N_7859,N_6087);
and U8461 (N_8461,N_7944,N_6160);
and U8462 (N_8462,N_6025,N_6033);
and U8463 (N_8463,N_6612,N_6598);
xor U8464 (N_8464,N_7301,N_7614);
nand U8465 (N_8465,N_6106,N_6053);
and U8466 (N_8466,N_6121,N_7925);
and U8467 (N_8467,N_7190,N_6992);
or U8468 (N_8468,N_6135,N_7295);
xor U8469 (N_8469,N_7135,N_7147);
or U8470 (N_8470,N_7982,N_7411);
and U8471 (N_8471,N_7699,N_7848);
nand U8472 (N_8472,N_6799,N_6869);
xor U8473 (N_8473,N_7555,N_7061);
nor U8474 (N_8474,N_6618,N_6300);
or U8475 (N_8475,N_7888,N_7675);
and U8476 (N_8476,N_6889,N_7106);
xnor U8477 (N_8477,N_6593,N_7446);
nand U8478 (N_8478,N_7933,N_7274);
or U8479 (N_8479,N_6698,N_6012);
xor U8480 (N_8480,N_6826,N_7964);
nand U8481 (N_8481,N_6986,N_7891);
xor U8482 (N_8482,N_7777,N_7632);
and U8483 (N_8483,N_6592,N_6321);
or U8484 (N_8484,N_6897,N_6386);
and U8485 (N_8485,N_6769,N_7393);
or U8486 (N_8486,N_6205,N_7710);
and U8487 (N_8487,N_6806,N_7332);
or U8488 (N_8488,N_6926,N_7334);
nor U8489 (N_8489,N_6478,N_7739);
nand U8490 (N_8490,N_7942,N_6307);
or U8491 (N_8491,N_6367,N_7895);
or U8492 (N_8492,N_7458,N_7561);
and U8493 (N_8493,N_6505,N_7574);
nand U8494 (N_8494,N_6843,N_7579);
or U8495 (N_8495,N_6496,N_6189);
or U8496 (N_8496,N_6721,N_7961);
nand U8497 (N_8497,N_6784,N_7088);
or U8498 (N_8498,N_7839,N_7175);
nor U8499 (N_8499,N_7323,N_7535);
nor U8500 (N_8500,N_7182,N_6636);
or U8501 (N_8501,N_6558,N_6727);
nand U8502 (N_8502,N_6842,N_7671);
and U8503 (N_8503,N_6789,N_7399);
and U8504 (N_8504,N_6113,N_7367);
or U8505 (N_8505,N_6531,N_6380);
nand U8506 (N_8506,N_6564,N_6672);
nor U8507 (N_8507,N_6282,N_7168);
nand U8508 (N_8508,N_6472,N_6397);
xnor U8509 (N_8509,N_7136,N_7249);
nand U8510 (N_8510,N_6357,N_7941);
and U8511 (N_8511,N_6313,N_6891);
nand U8512 (N_8512,N_6557,N_7782);
nor U8513 (N_8513,N_7817,N_7025);
and U8514 (N_8514,N_7423,N_6801);
nand U8515 (N_8515,N_7356,N_6860);
or U8516 (N_8516,N_6323,N_7691);
or U8517 (N_8517,N_6523,N_6067);
or U8518 (N_8518,N_6628,N_7404);
nand U8519 (N_8519,N_7383,N_6424);
xor U8520 (N_8520,N_6429,N_6879);
or U8521 (N_8521,N_7733,N_6231);
and U8522 (N_8522,N_6648,N_7237);
nand U8523 (N_8523,N_7619,N_7214);
and U8524 (N_8524,N_6267,N_7943);
nand U8525 (N_8525,N_7024,N_7486);
and U8526 (N_8526,N_7566,N_6649);
nand U8527 (N_8527,N_7126,N_6340);
nand U8528 (N_8528,N_7781,N_7479);
or U8529 (N_8529,N_7772,N_6447);
or U8530 (N_8530,N_7221,N_6006);
nor U8531 (N_8531,N_7537,N_6921);
nand U8532 (N_8532,N_7138,N_7616);
or U8533 (N_8533,N_7476,N_7767);
or U8534 (N_8534,N_6164,N_6773);
or U8535 (N_8535,N_7805,N_7224);
nor U8536 (N_8536,N_7461,N_7509);
nor U8537 (N_8537,N_7717,N_6506);
and U8538 (N_8538,N_6900,N_7358);
nand U8539 (N_8539,N_6084,N_6225);
or U8540 (N_8540,N_6257,N_7688);
or U8541 (N_8541,N_7081,N_7256);
and U8542 (N_8542,N_7716,N_7072);
nand U8543 (N_8543,N_7605,N_7842);
and U8544 (N_8544,N_6770,N_6325);
or U8545 (N_8545,N_7779,N_6452);
nand U8546 (N_8546,N_7860,N_6158);
nor U8547 (N_8547,N_6268,N_6834);
and U8548 (N_8548,N_6867,N_7235);
and U8549 (N_8549,N_6930,N_7210);
nand U8550 (N_8550,N_7773,N_7209);
or U8551 (N_8551,N_6695,N_7350);
nor U8552 (N_8552,N_7105,N_6570);
nor U8553 (N_8553,N_6417,N_6795);
or U8554 (N_8554,N_7058,N_7015);
nand U8555 (N_8555,N_7374,N_6029);
or U8556 (N_8556,N_7623,N_7385);
xnor U8557 (N_8557,N_7960,N_7187);
nor U8558 (N_8558,N_7991,N_6997);
nand U8559 (N_8559,N_7928,N_6370);
nand U8560 (N_8560,N_6440,N_7587);
and U8561 (N_8561,N_7747,N_7708);
xor U8562 (N_8562,N_6009,N_6358);
nand U8563 (N_8563,N_7443,N_6057);
nand U8564 (N_8564,N_6192,N_7313);
or U8565 (N_8565,N_7127,N_7364);
and U8566 (N_8566,N_6182,N_6473);
and U8567 (N_8567,N_6850,N_6309);
nor U8568 (N_8568,N_7273,N_7236);
and U8569 (N_8569,N_6973,N_7594);
xor U8570 (N_8570,N_6928,N_7119);
nand U8571 (N_8571,N_7836,N_6616);
xor U8572 (N_8572,N_7415,N_6516);
xor U8573 (N_8573,N_6601,N_6463);
nand U8574 (N_8574,N_6276,N_6169);
or U8575 (N_8575,N_6811,N_6096);
nor U8576 (N_8576,N_6951,N_6483);
and U8577 (N_8577,N_7732,N_6274);
xnor U8578 (N_8578,N_6371,N_6234);
or U8579 (N_8579,N_7010,N_6171);
or U8580 (N_8580,N_6181,N_7827);
and U8581 (N_8581,N_7047,N_7319);
and U8582 (N_8582,N_7317,N_7998);
nand U8583 (N_8583,N_6008,N_6277);
nor U8584 (N_8584,N_7935,N_7033);
nor U8585 (N_8585,N_7087,N_6107);
and U8586 (N_8586,N_7039,N_7222);
nand U8587 (N_8587,N_6379,N_6175);
nor U8588 (N_8588,N_7238,N_6728);
nor U8589 (N_8589,N_6524,N_6777);
nand U8590 (N_8590,N_7074,N_6681);
nor U8591 (N_8591,N_6946,N_6421);
or U8592 (N_8592,N_7172,N_7789);
nand U8593 (N_8593,N_7693,N_7259);
or U8594 (N_8594,N_7754,N_7020);
nand U8595 (N_8595,N_7700,N_6443);
xnor U8596 (N_8596,N_7956,N_7756);
and U8597 (N_8597,N_7639,N_7665);
nor U8598 (N_8598,N_7795,N_6016);
and U8599 (N_8599,N_7112,N_7006);
nor U8600 (N_8600,N_7396,N_7611);
or U8601 (N_8601,N_7178,N_7567);
nand U8602 (N_8602,N_6493,N_6079);
nand U8603 (N_8603,N_7232,N_7725);
nand U8604 (N_8604,N_7909,N_6116);
xor U8605 (N_8605,N_7852,N_6936);
or U8606 (N_8606,N_7068,N_6423);
and U8607 (N_8607,N_6115,N_7636);
xor U8608 (N_8608,N_7286,N_7683);
or U8609 (N_8609,N_6685,N_7583);
or U8610 (N_8610,N_7601,N_7055);
or U8611 (N_8611,N_7682,N_7893);
nor U8612 (N_8612,N_7166,N_7595);
or U8613 (N_8613,N_6525,N_7674);
nor U8614 (N_8614,N_6562,N_6372);
or U8615 (N_8615,N_6074,N_7421);
xnor U8616 (N_8616,N_7582,N_6798);
nor U8617 (N_8617,N_6482,N_7585);
nor U8618 (N_8618,N_7170,N_7621);
or U8619 (N_8619,N_7559,N_6515);
nand U8620 (N_8620,N_7596,N_7243);
or U8621 (N_8621,N_7109,N_6193);
or U8622 (N_8622,N_7445,N_6464);
or U8623 (N_8623,N_7987,N_7315);
or U8624 (N_8624,N_7108,N_6269);
or U8625 (N_8625,N_6456,N_6149);
xnor U8626 (N_8626,N_6451,N_6003);
and U8627 (N_8627,N_6065,N_6792);
and U8628 (N_8628,N_7743,N_7853);
nand U8629 (N_8629,N_7186,N_6005);
nand U8630 (N_8630,N_6640,N_7531);
nand U8631 (N_8631,N_7937,N_7802);
nor U8632 (N_8632,N_6266,N_6740);
nor U8633 (N_8633,N_6832,N_6122);
and U8634 (N_8634,N_6632,N_7618);
nand U8635 (N_8635,N_7696,N_6856);
nor U8636 (N_8636,N_6384,N_7655);
nor U8637 (N_8637,N_7205,N_6876);
or U8638 (N_8638,N_6660,N_6216);
and U8639 (N_8639,N_6392,N_7247);
and U8640 (N_8640,N_6702,N_6037);
or U8641 (N_8641,N_7008,N_6290);
and U8642 (N_8642,N_6270,N_7371);
or U8643 (N_8643,N_7562,N_6289);
or U8644 (N_8644,N_6599,N_7426);
nand U8645 (N_8645,N_7094,N_6544);
nand U8646 (N_8646,N_7867,N_7715);
nor U8647 (N_8647,N_7775,N_6425);
xnor U8648 (N_8648,N_7824,N_6880);
nor U8649 (N_8649,N_7846,N_7216);
nor U8650 (N_8650,N_7413,N_7300);
and U8651 (N_8651,N_7851,N_7648);
or U8652 (N_8652,N_7826,N_7077);
nand U8653 (N_8653,N_7787,N_7279);
nor U8654 (N_8654,N_7386,N_6947);
or U8655 (N_8655,N_7449,N_6141);
nor U8656 (N_8656,N_6555,N_7276);
or U8657 (N_8657,N_6415,N_7929);
xor U8658 (N_8658,N_7116,N_6675);
and U8659 (N_8659,N_7570,N_7111);
nand U8660 (N_8660,N_6310,N_6703);
nor U8661 (N_8661,N_6190,N_6481);
nor U8662 (N_8662,N_6373,N_7883);
xnor U8663 (N_8663,N_6186,N_6993);
and U8664 (N_8664,N_7158,N_6400);
nor U8665 (N_8665,N_6430,N_7090);
nand U8666 (N_8666,N_6161,N_6051);
and U8667 (N_8667,N_7484,N_6508);
xnor U8668 (N_8668,N_7200,N_6362);
xor U8669 (N_8669,N_7288,N_6665);
and U8670 (N_8670,N_6957,N_6666);
nor U8671 (N_8671,N_7968,N_6729);
or U8672 (N_8672,N_7180,N_7519);
or U8673 (N_8673,N_7328,N_7120);
xor U8674 (N_8674,N_7752,N_6070);
nand U8675 (N_8675,N_6916,N_7352);
nand U8676 (N_8676,N_6617,N_7046);
and U8677 (N_8677,N_7948,N_6927);
xnor U8678 (N_8678,N_7040,N_6076);
nand U8679 (N_8679,N_6446,N_7793);
and U8680 (N_8680,N_6201,N_7419);
nand U8681 (N_8681,N_7177,N_6944);
xor U8682 (N_8682,N_7950,N_6571);
and U8683 (N_8683,N_6111,N_7197);
nor U8684 (N_8684,N_6866,N_7934);
and U8685 (N_8685,N_7730,N_6539);
nor U8686 (N_8686,N_7832,N_6977);
nand U8687 (N_8687,N_6034,N_6308);
and U8688 (N_8688,N_6092,N_7400);
nor U8689 (N_8689,N_6255,N_7448);
and U8690 (N_8690,N_6381,N_6511);
nand U8691 (N_8691,N_7097,N_6800);
or U8692 (N_8692,N_6075,N_6605);
nand U8693 (N_8693,N_6243,N_7861);
nand U8694 (N_8694,N_7890,N_6953);
nor U8695 (N_8695,N_6661,N_6822);
nand U8696 (N_8696,N_6056,N_6437);
nand U8697 (N_8697,N_6634,N_7353);
nand U8698 (N_8698,N_6779,N_7118);
nor U8699 (N_8699,N_6624,N_7281);
and U8700 (N_8700,N_7550,N_6288);
or U8701 (N_8701,N_7162,N_7397);
nand U8702 (N_8702,N_7736,N_6279);
and U8703 (N_8703,N_7272,N_7320);
or U8704 (N_8704,N_7464,N_7976);
nor U8705 (N_8705,N_6782,N_7524);
nor U8706 (N_8706,N_7215,N_7666);
nand U8707 (N_8707,N_7936,N_7206);
nor U8708 (N_8708,N_6574,N_7664);
nor U8709 (N_8709,N_7471,N_7335);
nor U8710 (N_8710,N_6896,N_6143);
or U8711 (N_8711,N_7021,N_7637);
or U8712 (N_8712,N_6630,N_6104);
or U8713 (N_8713,N_7568,N_6502);
or U8714 (N_8714,N_7129,N_7834);
or U8715 (N_8715,N_6466,N_6514);
or U8716 (N_8716,N_6165,N_7225);
xor U8717 (N_8717,N_7201,N_7275);
nand U8718 (N_8718,N_7066,N_6152);
xor U8719 (N_8719,N_7018,N_6476);
or U8720 (N_8720,N_7692,N_7362);
nand U8721 (N_8721,N_7338,N_6328);
nor U8722 (N_8722,N_6657,N_7659);
nand U8723 (N_8723,N_7346,N_6875);
nand U8724 (N_8724,N_7528,N_7540);
or U8725 (N_8725,N_6909,N_6252);
and U8726 (N_8726,N_6360,N_7896);
nor U8727 (N_8727,N_6227,N_6664);
nand U8728 (N_8728,N_7673,N_6223);
or U8729 (N_8729,N_6837,N_6959);
and U8730 (N_8730,N_7508,N_6253);
or U8731 (N_8731,N_6207,N_6374);
and U8732 (N_8732,N_7496,N_7745);
and U8733 (N_8733,N_7270,N_6934);
and U8734 (N_8734,N_7351,N_7878);
and U8735 (N_8735,N_6366,N_6126);
and U8736 (N_8736,N_7239,N_6530);
or U8737 (N_8737,N_6796,N_7095);
nor U8738 (N_8738,N_7159,N_7337);
nor U8739 (N_8739,N_7114,N_6967);
or U8740 (N_8740,N_7296,N_6548);
nand U8741 (N_8741,N_7165,N_6206);
nor U8742 (N_8742,N_7433,N_7694);
and U8743 (N_8743,N_7631,N_7695);
or U8744 (N_8744,N_6154,N_7607);
xnor U8745 (N_8745,N_7657,N_7608);
and U8746 (N_8746,N_6133,N_7282);
or U8747 (N_8747,N_7712,N_6441);
nor U8748 (N_8748,N_6606,N_6655);
and U8749 (N_8749,N_6725,N_6710);
xor U8750 (N_8750,N_7872,N_7979);
and U8751 (N_8751,N_6042,N_6409);
nor U8752 (N_8752,N_7542,N_7417);
and U8753 (N_8753,N_6188,N_7470);
or U8754 (N_8754,N_6293,N_6942);
or U8755 (N_8755,N_7261,N_7780);
and U8756 (N_8756,N_7498,N_6743);
and U8757 (N_8757,N_6045,N_7897);
or U8758 (N_8758,N_7751,N_7875);
nor U8759 (N_8759,N_7881,N_6553);
nor U8760 (N_8760,N_6184,N_6861);
nor U8761 (N_8761,N_7604,N_6391);
and U8762 (N_8762,N_6814,N_7642);
and U8763 (N_8763,N_6427,N_7203);
or U8764 (N_8764,N_7546,N_6416);
xor U8765 (N_8765,N_7028,N_7302);
nand U8766 (N_8766,N_6911,N_7898);
nand U8767 (N_8767,N_7718,N_7248);
or U8768 (N_8768,N_7233,N_6990);
nor U8769 (N_8769,N_7152,N_6767);
xor U8770 (N_8770,N_7089,N_6063);
and U8771 (N_8771,N_7953,N_7635);
and U8772 (N_8772,N_6495,N_7822);
or U8773 (N_8773,N_6090,N_6128);
or U8774 (N_8774,N_6888,N_7543);
or U8775 (N_8775,N_6048,N_7431);
and U8776 (N_8776,N_7244,N_6462);
nand U8777 (N_8777,N_6015,N_6342);
nor U8778 (N_8778,N_7727,N_6651);
and U8779 (N_8779,N_7048,N_7148);
or U8780 (N_8780,N_6872,N_7501);
nand U8781 (N_8781,N_7945,N_7101);
nand U8782 (N_8782,N_6788,N_6955);
nor U8783 (N_8783,N_7698,N_6808);
nand U8784 (N_8784,N_6259,N_6220);
xor U8785 (N_8785,N_7034,N_6172);
nand U8786 (N_8786,N_6890,N_7481);
xnor U8787 (N_8787,N_6356,N_7290);
and U8788 (N_8788,N_6027,N_6187);
nor U8789 (N_8789,N_7847,N_7523);
or U8790 (N_8790,N_7711,N_6028);
nor U8791 (N_8791,N_7613,N_6265);
nor U8792 (N_8792,N_6354,N_7930);
or U8793 (N_8793,N_7223,N_6723);
and U8794 (N_8794,N_6600,N_7080);
nor U8795 (N_8795,N_6541,N_7085);
or U8796 (N_8796,N_6091,N_6529);
or U8797 (N_8797,N_7402,N_7609);
or U8798 (N_8798,N_7036,N_6263);
nand U8799 (N_8799,N_6346,N_7171);
xnor U8800 (N_8800,N_7766,N_7372);
nand U8801 (N_8801,N_6375,N_7922);
nor U8802 (N_8802,N_7654,N_6399);
nor U8803 (N_8803,N_7924,N_7439);
nor U8804 (N_8804,N_6791,N_6771);
nor U8805 (N_8805,N_6528,N_6199);
nand U8806 (N_8806,N_6923,N_7265);
and U8807 (N_8807,N_7746,N_7260);
xnor U8808 (N_8808,N_7154,N_7617);
or U8809 (N_8809,N_6688,N_7643);
nor U8810 (N_8810,N_7318,N_6445);
or U8811 (N_8811,N_6717,N_7375);
or U8812 (N_8812,N_7557,N_6576);
nor U8813 (N_8813,N_6448,N_7440);
or U8814 (N_8814,N_6442,N_6208);
and U8815 (N_8815,N_6222,N_6733);
and U8816 (N_8816,N_7212,N_6741);
or U8817 (N_8817,N_6595,N_6841);
and U8818 (N_8818,N_7939,N_7955);
and U8819 (N_8819,N_6339,N_6623);
xnor U8820 (N_8820,N_6969,N_6219);
and U8821 (N_8821,N_7340,N_6230);
and U8822 (N_8822,N_7307,N_6893);
nor U8823 (N_8823,N_7192,N_7902);
xnor U8824 (N_8824,N_7527,N_6504);
nor U8825 (N_8825,N_6827,N_6264);
nor U8826 (N_8826,N_7078,N_7807);
nor U8827 (N_8827,N_7722,N_6971);
and U8828 (N_8828,N_6699,N_7407);
xnor U8829 (N_8829,N_7430,N_6762);
or U8830 (N_8830,N_6271,N_6060);
or U8831 (N_8831,N_6318,N_7029);
or U8832 (N_8832,N_6816,N_7451);
or U8833 (N_8833,N_7258,N_7905);
nor U8834 (N_8834,N_6565,N_6426);
or U8835 (N_8835,N_6332,N_6191);
nand U8836 (N_8836,N_6844,N_6238);
nand U8837 (N_8837,N_6062,N_6836);
xor U8838 (N_8838,N_6283,N_6098);
nand U8839 (N_8839,N_7704,N_7749);
nand U8840 (N_8840,N_6754,N_7753);
nor U8841 (N_8841,N_7045,N_6353);
nand U8842 (N_8842,N_7532,N_7816);
nand U8843 (N_8843,N_6244,N_7572);
nand U8844 (N_8844,N_6450,N_6258);
or U8845 (N_8845,N_7231,N_6904);
nor U8846 (N_8846,N_6708,N_6793);
xnor U8847 (N_8847,N_7257,N_7395);
and U8848 (N_8848,N_6047,N_7251);
nand U8849 (N_8849,N_6486,N_7769);
nand U8850 (N_8850,N_6902,N_6831);
or U8851 (N_8851,N_7873,N_7973);
or U8852 (N_8852,N_6387,N_7360);
nor U8853 (N_8853,N_6653,N_6136);
and U8854 (N_8854,N_6637,N_7189);
nor U8855 (N_8855,N_6287,N_6468);
or U8856 (N_8856,N_7744,N_6989);
and U8857 (N_8857,N_7996,N_7195);
nor U8858 (N_8858,N_6536,N_7388);
nand U8859 (N_8859,N_6948,N_7041);
or U8860 (N_8860,N_7625,N_6101);
xnor U8861 (N_8861,N_7926,N_6556);
xnor U8862 (N_8862,N_6303,N_6061);
xnor U8863 (N_8863,N_7602,N_7652);
or U8864 (N_8864,N_6026,N_6044);
and U8865 (N_8865,N_7298,N_7163);
nand U8866 (N_8866,N_6579,N_7615);
and U8867 (N_8867,N_6821,N_6642);
and U8868 (N_8868,N_6978,N_7963);
or U8869 (N_8869,N_7549,N_6211);
and U8870 (N_8870,N_7493,N_6110);
nor U8871 (N_8871,N_7339,N_6322);
or U8872 (N_8872,N_7957,N_6229);
nor U8873 (N_8873,N_6868,N_7255);
nand U8874 (N_8874,N_7678,N_6140);
and U8875 (N_8875,N_7266,N_6980);
nand U8876 (N_8876,N_6331,N_6338);
nand U8877 (N_8877,N_7414,N_6148);
and U8878 (N_8878,N_6260,N_6507);
and U8879 (N_8879,N_6625,N_6833);
or U8880 (N_8880,N_7208,N_6984);
xor U8881 (N_8881,N_6547,N_7576);
nand U8882 (N_8882,N_6580,N_6418);
nor U8883 (N_8883,N_6696,N_6517);
and U8884 (N_8884,N_6347,N_6994);
and U8885 (N_8885,N_7217,N_7850);
and U8886 (N_8886,N_6248,N_7843);
or U8887 (N_8887,N_7719,N_7103);
and U8888 (N_8888,N_6083,N_6820);
and U8889 (N_8889,N_6146,N_6077);
or U8890 (N_8890,N_6906,N_6684);
xor U8891 (N_8891,N_6335,N_6108);
nor U8892 (N_8892,N_6862,N_6610);
or U8893 (N_8893,N_6554,N_7229);
nand U8894 (N_8894,N_6395,N_6197);
nor U8895 (N_8895,N_6469,N_7344);
or U8896 (N_8896,N_6522,N_6886);
or U8897 (N_8897,N_7179,N_6333);
or U8898 (N_8898,N_7063,N_7219);
xnor U8899 (N_8899,N_6691,N_7412);
and U8900 (N_8900,N_6431,N_6537);
nor U8901 (N_8901,N_6638,N_7123);
nor U8902 (N_8902,N_6492,N_6750);
and U8903 (N_8903,N_7823,N_6765);
or U8904 (N_8904,N_7156,N_6272);
nand U8905 (N_8905,N_7798,N_7992);
or U8906 (N_8906,N_6755,N_7245);
and U8907 (N_8907,N_7522,N_7612);
and U8908 (N_8908,N_7141,N_7181);
nand U8909 (N_8909,N_7768,N_6454);
nor U8910 (N_8910,N_7355,N_6714);
nor U8911 (N_8911,N_7321,N_7050);
and U8912 (N_8912,N_7287,N_6080);
nor U8913 (N_8913,N_6509,N_7677);
nand U8914 (N_8914,N_7324,N_6887);
or U8915 (N_8915,N_7031,N_7466);
and U8916 (N_8916,N_6488,N_7349);
or U8917 (N_8917,N_7390,N_6150);
nor U8918 (N_8918,N_6533,N_6177);
nor U8919 (N_8919,N_6176,N_7731);
or U8920 (N_8920,N_7762,N_7155);
or U8921 (N_8921,N_7603,N_6280);
nor U8922 (N_8922,N_7357,N_6202);
or U8923 (N_8923,N_7204,N_6351);
nor U8924 (N_8924,N_6818,N_7075);
nand U8925 (N_8925,N_6884,N_7191);
and U8926 (N_8926,N_7472,N_6018);
nand U8927 (N_8927,N_7680,N_6534);
nor U8928 (N_8928,N_6410,N_6404);
or U8929 (N_8929,N_6241,N_7676);
or U8930 (N_8930,N_6742,N_6382);
nand U8931 (N_8931,N_7394,N_7309);
or U8932 (N_8932,N_7510,N_6278);
and U8933 (N_8933,N_7892,N_6621);
nand U8934 (N_8934,N_6173,N_7038);
nand U8935 (N_8935,N_6412,N_6209);
or U8936 (N_8936,N_6613,N_7518);
nand U8937 (N_8937,N_7429,N_7376);
or U8938 (N_8938,N_6078,N_6937);
and U8939 (N_8939,N_6117,N_7833);
nand U8940 (N_8940,N_7954,N_6663);
or U8941 (N_8941,N_7516,N_6932);
xor U8942 (N_8942,N_6924,N_6298);
and U8943 (N_8943,N_6987,N_6692);
or U8944 (N_8944,N_7325,N_6232);
or U8945 (N_8945,N_6914,N_7899);
nor U8946 (N_8946,N_7207,N_7403);
or U8947 (N_8947,N_6709,N_7438);
nand U8948 (N_8948,N_7679,N_6432);
and U8949 (N_8949,N_7277,N_7453);
nand U8950 (N_8950,N_7406,N_6261);
nor U8951 (N_8951,N_6864,N_6810);
nor U8952 (N_8952,N_6586,N_7100);
nand U8953 (N_8953,N_6970,N_7520);
or U8954 (N_8954,N_6797,N_7759);
nand U8955 (N_8955,N_7202,N_6687);
xnor U8956 (N_8956,N_6139,N_6590);
or U8957 (N_8957,N_6281,N_6766);
nand U8958 (N_8958,N_7879,N_7113);
and U8959 (N_8959,N_6615,N_6724);
or U8960 (N_8960,N_7425,N_6498);
and U8961 (N_8961,N_7705,N_7799);
nor U8962 (N_8962,N_7468,N_6329);
nand U8963 (N_8963,N_6918,N_7240);
xor U8964 (N_8964,N_7091,N_7115);
xnor U8965 (N_8965,N_6302,N_7662);
and U8966 (N_8966,N_6635,N_7289);
and U8967 (N_8967,N_6368,N_6345);
nand U8968 (N_8968,N_7885,N_7620);
and U8969 (N_8969,N_7904,N_6457);
or U8970 (N_8970,N_7283,N_7783);
or U8971 (N_8971,N_7469,N_6072);
and U8972 (N_8972,N_6677,N_6550);
nand U8973 (N_8973,N_7495,N_6915);
nor U8974 (N_8974,N_6650,N_7713);
nor U8975 (N_8975,N_7920,N_6566);
nand U8976 (N_8976,N_6964,N_6982);
nor U8977 (N_8977,N_6470,N_7456);
and U8978 (N_8978,N_6803,N_7218);
and U8979 (N_8979,N_6017,N_6359);
and U8980 (N_8980,N_6738,N_7803);
nand U8981 (N_8981,N_7512,N_7598);
or U8982 (N_8982,N_6262,N_7143);
and U8983 (N_8983,N_6774,N_7738);
or U8984 (N_8984,N_6144,N_6251);
nor U8985 (N_8985,N_6242,N_7121);
and U8986 (N_8986,N_7474,N_6731);
and U8987 (N_8987,N_6458,N_6341);
xnor U8988 (N_8988,N_6185,N_7997);
nand U8989 (N_8989,N_7720,N_6718);
nor U8990 (N_8990,N_6105,N_7573);
or U8991 (N_8991,N_6355,N_6697);
nor U8992 (N_8992,N_6284,N_6913);
or U8993 (N_8993,N_6701,N_6652);
or U8994 (N_8994,N_6480,N_7886);
nor U8995 (N_8995,N_7995,N_6940);
nand U8996 (N_8996,N_7774,N_6100);
or U8997 (N_8997,N_6050,N_7492);
or U8998 (N_8998,N_6240,N_6125);
nor U8999 (N_8999,N_6097,N_7551);
nor U9000 (N_9000,N_6291,N_7043);
nand U9001 (N_9001,N_6969,N_7353);
nor U9002 (N_9002,N_7884,N_7306);
or U9003 (N_9003,N_7385,N_6105);
and U9004 (N_9004,N_6990,N_7245);
xor U9005 (N_9005,N_7475,N_7769);
nand U9006 (N_9006,N_7979,N_7818);
nand U9007 (N_9007,N_7714,N_6495);
or U9008 (N_9008,N_6940,N_7313);
or U9009 (N_9009,N_6796,N_7292);
xor U9010 (N_9010,N_7987,N_7790);
or U9011 (N_9011,N_6364,N_6756);
nor U9012 (N_9012,N_7160,N_6454);
and U9013 (N_9013,N_6312,N_7449);
nor U9014 (N_9014,N_7730,N_7555);
nand U9015 (N_9015,N_7890,N_7401);
nor U9016 (N_9016,N_7445,N_7993);
nor U9017 (N_9017,N_7746,N_6931);
nand U9018 (N_9018,N_7244,N_6047);
xnor U9019 (N_9019,N_6793,N_6989);
nand U9020 (N_9020,N_7300,N_6039);
or U9021 (N_9021,N_7342,N_7224);
or U9022 (N_9022,N_7735,N_7859);
nand U9023 (N_9023,N_6007,N_7158);
nor U9024 (N_9024,N_7949,N_6661);
xor U9025 (N_9025,N_7024,N_7015);
or U9026 (N_9026,N_7255,N_7921);
nor U9027 (N_9027,N_7886,N_7987);
nand U9028 (N_9028,N_6147,N_7109);
nor U9029 (N_9029,N_7928,N_6563);
xor U9030 (N_9030,N_7646,N_7151);
nor U9031 (N_9031,N_6669,N_6609);
nand U9032 (N_9032,N_6759,N_7680);
and U9033 (N_9033,N_7554,N_6753);
nor U9034 (N_9034,N_7055,N_7923);
xor U9035 (N_9035,N_6522,N_7376);
xor U9036 (N_9036,N_6057,N_6826);
nor U9037 (N_9037,N_7892,N_6460);
nand U9038 (N_9038,N_7997,N_7140);
xor U9039 (N_9039,N_6289,N_6162);
nand U9040 (N_9040,N_6148,N_7062);
or U9041 (N_9041,N_7712,N_6398);
and U9042 (N_9042,N_6997,N_7661);
and U9043 (N_9043,N_7782,N_6305);
nand U9044 (N_9044,N_6840,N_6038);
and U9045 (N_9045,N_7032,N_6526);
nand U9046 (N_9046,N_6978,N_7274);
nor U9047 (N_9047,N_7988,N_6425);
nor U9048 (N_9048,N_7449,N_7805);
and U9049 (N_9049,N_7123,N_6172);
nand U9050 (N_9050,N_6912,N_6508);
or U9051 (N_9051,N_7622,N_6738);
and U9052 (N_9052,N_6312,N_6630);
and U9053 (N_9053,N_6773,N_6714);
nor U9054 (N_9054,N_6631,N_6138);
xor U9055 (N_9055,N_6195,N_7592);
nor U9056 (N_9056,N_7633,N_7725);
and U9057 (N_9057,N_7637,N_6887);
nand U9058 (N_9058,N_7054,N_6328);
nor U9059 (N_9059,N_7914,N_7144);
and U9060 (N_9060,N_7814,N_7835);
nand U9061 (N_9061,N_6654,N_7592);
nor U9062 (N_9062,N_7089,N_6703);
nor U9063 (N_9063,N_7628,N_6995);
nand U9064 (N_9064,N_6916,N_6518);
xnor U9065 (N_9065,N_6584,N_7099);
nand U9066 (N_9066,N_7152,N_7411);
and U9067 (N_9067,N_6682,N_7620);
or U9068 (N_9068,N_6055,N_6186);
and U9069 (N_9069,N_7235,N_6525);
nand U9070 (N_9070,N_6667,N_6051);
or U9071 (N_9071,N_6027,N_6288);
and U9072 (N_9072,N_7069,N_7995);
nor U9073 (N_9073,N_6767,N_6092);
and U9074 (N_9074,N_7375,N_7391);
nand U9075 (N_9075,N_7036,N_7606);
nor U9076 (N_9076,N_7777,N_6936);
nand U9077 (N_9077,N_7067,N_7282);
and U9078 (N_9078,N_7021,N_6445);
and U9079 (N_9079,N_6285,N_6119);
nand U9080 (N_9080,N_6737,N_6839);
nand U9081 (N_9081,N_7079,N_7840);
nor U9082 (N_9082,N_7351,N_7165);
nor U9083 (N_9083,N_7540,N_7373);
nor U9084 (N_9084,N_7690,N_6074);
or U9085 (N_9085,N_6661,N_6763);
and U9086 (N_9086,N_7535,N_6605);
or U9087 (N_9087,N_6356,N_6778);
or U9088 (N_9088,N_6955,N_7904);
and U9089 (N_9089,N_7763,N_6538);
nand U9090 (N_9090,N_7305,N_6190);
and U9091 (N_9091,N_7276,N_7575);
nand U9092 (N_9092,N_7133,N_7333);
or U9093 (N_9093,N_7582,N_6315);
nand U9094 (N_9094,N_7999,N_7391);
nand U9095 (N_9095,N_6839,N_6916);
or U9096 (N_9096,N_6897,N_7321);
nor U9097 (N_9097,N_6396,N_6650);
nor U9098 (N_9098,N_7017,N_6135);
xnor U9099 (N_9099,N_7238,N_6513);
or U9100 (N_9100,N_6663,N_6393);
nand U9101 (N_9101,N_7787,N_7973);
and U9102 (N_9102,N_7456,N_6439);
nor U9103 (N_9103,N_7939,N_7851);
and U9104 (N_9104,N_6290,N_6186);
or U9105 (N_9105,N_7530,N_7954);
nand U9106 (N_9106,N_6848,N_6434);
nor U9107 (N_9107,N_6632,N_7210);
and U9108 (N_9108,N_7017,N_6505);
or U9109 (N_9109,N_7710,N_6948);
nand U9110 (N_9110,N_6109,N_6995);
nand U9111 (N_9111,N_6045,N_6770);
nand U9112 (N_9112,N_7072,N_7882);
and U9113 (N_9113,N_6871,N_6235);
nand U9114 (N_9114,N_7624,N_7470);
nand U9115 (N_9115,N_6398,N_6023);
nor U9116 (N_9116,N_6140,N_7995);
and U9117 (N_9117,N_7475,N_6710);
nand U9118 (N_9118,N_7683,N_7651);
nand U9119 (N_9119,N_7087,N_7744);
and U9120 (N_9120,N_6932,N_6976);
and U9121 (N_9121,N_7832,N_7857);
and U9122 (N_9122,N_7264,N_7627);
nor U9123 (N_9123,N_7907,N_7717);
or U9124 (N_9124,N_6456,N_7719);
nand U9125 (N_9125,N_6272,N_6280);
nand U9126 (N_9126,N_6673,N_7778);
nand U9127 (N_9127,N_6339,N_7439);
nand U9128 (N_9128,N_6588,N_6785);
or U9129 (N_9129,N_7956,N_7365);
and U9130 (N_9130,N_7049,N_6240);
nor U9131 (N_9131,N_6325,N_6623);
and U9132 (N_9132,N_7730,N_6094);
and U9133 (N_9133,N_6933,N_7717);
nor U9134 (N_9134,N_6565,N_6222);
nor U9135 (N_9135,N_6862,N_6177);
and U9136 (N_9136,N_7440,N_6636);
and U9137 (N_9137,N_7856,N_7688);
nand U9138 (N_9138,N_6528,N_6769);
nor U9139 (N_9139,N_6889,N_6024);
and U9140 (N_9140,N_6354,N_6843);
nor U9141 (N_9141,N_6984,N_7124);
or U9142 (N_9142,N_6105,N_6959);
or U9143 (N_9143,N_6913,N_6426);
xor U9144 (N_9144,N_7775,N_6717);
and U9145 (N_9145,N_7620,N_7061);
or U9146 (N_9146,N_7412,N_6793);
xnor U9147 (N_9147,N_7055,N_6784);
xor U9148 (N_9148,N_6149,N_7265);
nand U9149 (N_9149,N_6924,N_7076);
and U9150 (N_9150,N_6875,N_7400);
and U9151 (N_9151,N_6837,N_7028);
nor U9152 (N_9152,N_7143,N_7180);
and U9153 (N_9153,N_7095,N_7235);
and U9154 (N_9154,N_6284,N_6728);
or U9155 (N_9155,N_7899,N_7396);
nand U9156 (N_9156,N_7978,N_7429);
nand U9157 (N_9157,N_7708,N_7546);
nor U9158 (N_9158,N_7231,N_6300);
nand U9159 (N_9159,N_6053,N_6252);
xnor U9160 (N_9160,N_7368,N_7793);
and U9161 (N_9161,N_6437,N_7462);
and U9162 (N_9162,N_7308,N_7379);
nor U9163 (N_9163,N_6351,N_7936);
or U9164 (N_9164,N_7555,N_7207);
and U9165 (N_9165,N_6680,N_7063);
nor U9166 (N_9166,N_6431,N_6873);
and U9167 (N_9167,N_6489,N_6194);
nand U9168 (N_9168,N_7758,N_6752);
xor U9169 (N_9169,N_6794,N_7332);
or U9170 (N_9170,N_7861,N_7432);
nand U9171 (N_9171,N_7075,N_7197);
or U9172 (N_9172,N_6978,N_6922);
nor U9173 (N_9173,N_7330,N_6852);
nor U9174 (N_9174,N_6385,N_7037);
or U9175 (N_9175,N_7610,N_6882);
nor U9176 (N_9176,N_6758,N_6017);
nand U9177 (N_9177,N_6172,N_7903);
and U9178 (N_9178,N_6458,N_7199);
nand U9179 (N_9179,N_6762,N_6858);
nand U9180 (N_9180,N_6325,N_7285);
and U9181 (N_9181,N_7902,N_6315);
nor U9182 (N_9182,N_7814,N_7010);
nand U9183 (N_9183,N_7729,N_7186);
xor U9184 (N_9184,N_6255,N_6406);
nor U9185 (N_9185,N_7792,N_7028);
xnor U9186 (N_9186,N_6404,N_7983);
nand U9187 (N_9187,N_7532,N_7659);
nor U9188 (N_9188,N_6089,N_6565);
xor U9189 (N_9189,N_7067,N_7207);
nand U9190 (N_9190,N_7439,N_7178);
nand U9191 (N_9191,N_7493,N_7130);
or U9192 (N_9192,N_7391,N_6075);
nor U9193 (N_9193,N_6022,N_7779);
nor U9194 (N_9194,N_7321,N_6927);
nor U9195 (N_9195,N_7254,N_7498);
or U9196 (N_9196,N_6288,N_7190);
nor U9197 (N_9197,N_6659,N_6730);
or U9198 (N_9198,N_6055,N_6610);
or U9199 (N_9199,N_6710,N_6975);
nor U9200 (N_9200,N_6430,N_7524);
xor U9201 (N_9201,N_7350,N_6342);
and U9202 (N_9202,N_6861,N_6319);
or U9203 (N_9203,N_6295,N_7663);
nor U9204 (N_9204,N_6110,N_7479);
or U9205 (N_9205,N_6070,N_7820);
nor U9206 (N_9206,N_6393,N_6020);
xnor U9207 (N_9207,N_7877,N_6284);
xnor U9208 (N_9208,N_7126,N_7433);
and U9209 (N_9209,N_7211,N_6829);
xor U9210 (N_9210,N_7930,N_7087);
and U9211 (N_9211,N_6504,N_6388);
nor U9212 (N_9212,N_7780,N_7402);
nand U9213 (N_9213,N_6441,N_6596);
nor U9214 (N_9214,N_7425,N_6625);
nand U9215 (N_9215,N_7556,N_6819);
nand U9216 (N_9216,N_6179,N_7907);
or U9217 (N_9217,N_6231,N_6525);
nand U9218 (N_9218,N_7556,N_7489);
nand U9219 (N_9219,N_6309,N_6553);
or U9220 (N_9220,N_6832,N_6411);
and U9221 (N_9221,N_7189,N_7559);
or U9222 (N_9222,N_6530,N_6481);
nand U9223 (N_9223,N_7525,N_7876);
nand U9224 (N_9224,N_6572,N_6721);
or U9225 (N_9225,N_7027,N_7209);
or U9226 (N_9226,N_6631,N_7958);
and U9227 (N_9227,N_7920,N_6487);
nor U9228 (N_9228,N_7579,N_6228);
or U9229 (N_9229,N_7234,N_7456);
nor U9230 (N_9230,N_6593,N_6295);
nand U9231 (N_9231,N_7441,N_6367);
or U9232 (N_9232,N_6439,N_6836);
nor U9233 (N_9233,N_7274,N_6127);
nor U9234 (N_9234,N_6567,N_7866);
nand U9235 (N_9235,N_7102,N_6641);
or U9236 (N_9236,N_7741,N_6220);
and U9237 (N_9237,N_7563,N_6409);
nor U9238 (N_9238,N_7771,N_6641);
nor U9239 (N_9239,N_6283,N_7176);
or U9240 (N_9240,N_6004,N_6527);
xnor U9241 (N_9241,N_7890,N_7856);
or U9242 (N_9242,N_7314,N_7145);
or U9243 (N_9243,N_7358,N_6636);
nor U9244 (N_9244,N_7516,N_6681);
and U9245 (N_9245,N_6115,N_7360);
nor U9246 (N_9246,N_7248,N_7862);
nand U9247 (N_9247,N_7914,N_6182);
or U9248 (N_9248,N_6907,N_7132);
or U9249 (N_9249,N_6677,N_6915);
or U9250 (N_9250,N_7363,N_7633);
or U9251 (N_9251,N_7245,N_6491);
or U9252 (N_9252,N_7623,N_6319);
and U9253 (N_9253,N_6866,N_6099);
and U9254 (N_9254,N_7283,N_6107);
nor U9255 (N_9255,N_7721,N_7557);
nand U9256 (N_9256,N_6418,N_6190);
and U9257 (N_9257,N_7963,N_6392);
nand U9258 (N_9258,N_6531,N_7323);
and U9259 (N_9259,N_6098,N_7469);
and U9260 (N_9260,N_7257,N_6193);
xor U9261 (N_9261,N_7592,N_7623);
and U9262 (N_9262,N_7422,N_6013);
or U9263 (N_9263,N_6949,N_7203);
or U9264 (N_9264,N_7868,N_6606);
nor U9265 (N_9265,N_7984,N_7286);
and U9266 (N_9266,N_7099,N_7091);
and U9267 (N_9267,N_6323,N_6388);
and U9268 (N_9268,N_7858,N_6364);
and U9269 (N_9269,N_7100,N_7409);
nand U9270 (N_9270,N_7434,N_7725);
or U9271 (N_9271,N_7395,N_7346);
and U9272 (N_9272,N_6776,N_7948);
nand U9273 (N_9273,N_6819,N_6491);
or U9274 (N_9274,N_7533,N_6953);
nor U9275 (N_9275,N_6921,N_7701);
or U9276 (N_9276,N_7935,N_6299);
and U9277 (N_9277,N_6638,N_7249);
xnor U9278 (N_9278,N_6868,N_6517);
nand U9279 (N_9279,N_7690,N_6929);
and U9280 (N_9280,N_7400,N_7816);
and U9281 (N_9281,N_6200,N_7241);
or U9282 (N_9282,N_7206,N_6339);
and U9283 (N_9283,N_6072,N_6456);
nand U9284 (N_9284,N_7894,N_7746);
nor U9285 (N_9285,N_7117,N_6656);
and U9286 (N_9286,N_6772,N_7943);
nor U9287 (N_9287,N_6440,N_6376);
or U9288 (N_9288,N_7415,N_6232);
and U9289 (N_9289,N_7677,N_6306);
nand U9290 (N_9290,N_6380,N_6373);
xnor U9291 (N_9291,N_7328,N_6848);
and U9292 (N_9292,N_6422,N_7546);
nor U9293 (N_9293,N_6175,N_6251);
and U9294 (N_9294,N_7882,N_6905);
nor U9295 (N_9295,N_6672,N_6355);
xor U9296 (N_9296,N_7027,N_7127);
and U9297 (N_9297,N_6401,N_6891);
and U9298 (N_9298,N_7230,N_7065);
xnor U9299 (N_9299,N_7510,N_7714);
nand U9300 (N_9300,N_6629,N_7146);
xor U9301 (N_9301,N_7136,N_7219);
xnor U9302 (N_9302,N_6640,N_7484);
and U9303 (N_9303,N_7649,N_7417);
and U9304 (N_9304,N_7394,N_6561);
and U9305 (N_9305,N_6846,N_6380);
and U9306 (N_9306,N_6001,N_6568);
nand U9307 (N_9307,N_7143,N_7182);
nor U9308 (N_9308,N_7171,N_6517);
or U9309 (N_9309,N_6407,N_7399);
nand U9310 (N_9310,N_6234,N_7278);
nor U9311 (N_9311,N_6173,N_7562);
or U9312 (N_9312,N_7676,N_7932);
nand U9313 (N_9313,N_6717,N_6804);
or U9314 (N_9314,N_7874,N_7361);
xor U9315 (N_9315,N_6778,N_7158);
nand U9316 (N_9316,N_6720,N_6004);
and U9317 (N_9317,N_7611,N_7767);
nand U9318 (N_9318,N_7509,N_6383);
or U9319 (N_9319,N_6589,N_7337);
nor U9320 (N_9320,N_7747,N_6988);
and U9321 (N_9321,N_6148,N_6129);
nor U9322 (N_9322,N_7554,N_6099);
or U9323 (N_9323,N_6772,N_6607);
and U9324 (N_9324,N_6357,N_7563);
or U9325 (N_9325,N_7295,N_6957);
or U9326 (N_9326,N_7825,N_7726);
or U9327 (N_9327,N_6280,N_7569);
nand U9328 (N_9328,N_6630,N_7206);
nor U9329 (N_9329,N_7807,N_7431);
nand U9330 (N_9330,N_7544,N_6273);
or U9331 (N_9331,N_7704,N_6464);
or U9332 (N_9332,N_7147,N_6667);
nor U9333 (N_9333,N_7572,N_7420);
or U9334 (N_9334,N_7136,N_7475);
or U9335 (N_9335,N_7712,N_7166);
nand U9336 (N_9336,N_7549,N_6059);
nor U9337 (N_9337,N_7989,N_7232);
or U9338 (N_9338,N_6216,N_7570);
nand U9339 (N_9339,N_6918,N_7566);
or U9340 (N_9340,N_6671,N_7715);
xnor U9341 (N_9341,N_6538,N_7153);
and U9342 (N_9342,N_6494,N_6307);
and U9343 (N_9343,N_7185,N_7743);
or U9344 (N_9344,N_7635,N_7594);
or U9345 (N_9345,N_6118,N_7553);
and U9346 (N_9346,N_6733,N_7729);
nor U9347 (N_9347,N_6533,N_7477);
xor U9348 (N_9348,N_6535,N_6945);
and U9349 (N_9349,N_6761,N_7552);
nand U9350 (N_9350,N_7200,N_6383);
nand U9351 (N_9351,N_7395,N_6699);
or U9352 (N_9352,N_7439,N_7177);
nand U9353 (N_9353,N_7106,N_7815);
and U9354 (N_9354,N_6086,N_6455);
and U9355 (N_9355,N_7123,N_6397);
nand U9356 (N_9356,N_7455,N_7203);
xor U9357 (N_9357,N_7546,N_7737);
and U9358 (N_9358,N_7758,N_6585);
nor U9359 (N_9359,N_6664,N_7997);
nand U9360 (N_9360,N_7689,N_7792);
nor U9361 (N_9361,N_7814,N_7099);
nor U9362 (N_9362,N_7987,N_6074);
nand U9363 (N_9363,N_7473,N_6649);
and U9364 (N_9364,N_7080,N_7000);
nand U9365 (N_9365,N_6966,N_7506);
nor U9366 (N_9366,N_7183,N_7606);
nor U9367 (N_9367,N_7158,N_6450);
nand U9368 (N_9368,N_7614,N_6480);
nor U9369 (N_9369,N_7551,N_7510);
nor U9370 (N_9370,N_6913,N_7388);
nand U9371 (N_9371,N_6589,N_6458);
xor U9372 (N_9372,N_6120,N_6013);
and U9373 (N_9373,N_6496,N_6886);
and U9374 (N_9374,N_7260,N_7816);
and U9375 (N_9375,N_6538,N_7485);
nor U9376 (N_9376,N_6898,N_7235);
nand U9377 (N_9377,N_7234,N_7498);
and U9378 (N_9378,N_7807,N_6716);
nor U9379 (N_9379,N_6277,N_6446);
or U9380 (N_9380,N_7855,N_6011);
xor U9381 (N_9381,N_6255,N_7231);
nor U9382 (N_9382,N_7969,N_7485);
nor U9383 (N_9383,N_7853,N_7829);
nand U9384 (N_9384,N_6600,N_6531);
nand U9385 (N_9385,N_6570,N_7167);
and U9386 (N_9386,N_7778,N_6773);
and U9387 (N_9387,N_7194,N_7968);
nor U9388 (N_9388,N_7610,N_6923);
or U9389 (N_9389,N_6559,N_7466);
or U9390 (N_9390,N_7726,N_7520);
xor U9391 (N_9391,N_7745,N_6497);
nor U9392 (N_9392,N_6483,N_6311);
nand U9393 (N_9393,N_6586,N_6538);
nand U9394 (N_9394,N_6029,N_7119);
and U9395 (N_9395,N_6087,N_6035);
and U9396 (N_9396,N_6569,N_6337);
or U9397 (N_9397,N_6515,N_6081);
nor U9398 (N_9398,N_7713,N_6982);
nand U9399 (N_9399,N_7422,N_7880);
and U9400 (N_9400,N_7304,N_7341);
nand U9401 (N_9401,N_6325,N_7440);
and U9402 (N_9402,N_7019,N_7501);
xor U9403 (N_9403,N_7732,N_7247);
or U9404 (N_9404,N_7664,N_6752);
and U9405 (N_9405,N_6727,N_7081);
and U9406 (N_9406,N_7875,N_7865);
nand U9407 (N_9407,N_6287,N_7418);
nand U9408 (N_9408,N_7071,N_6905);
and U9409 (N_9409,N_7798,N_7877);
nand U9410 (N_9410,N_6729,N_7586);
or U9411 (N_9411,N_7585,N_6049);
and U9412 (N_9412,N_7596,N_6787);
or U9413 (N_9413,N_7093,N_6790);
and U9414 (N_9414,N_6134,N_6140);
and U9415 (N_9415,N_7593,N_6899);
or U9416 (N_9416,N_7325,N_6819);
or U9417 (N_9417,N_6984,N_6761);
and U9418 (N_9418,N_7056,N_6462);
and U9419 (N_9419,N_6253,N_7992);
and U9420 (N_9420,N_7993,N_6439);
or U9421 (N_9421,N_6485,N_7176);
nor U9422 (N_9422,N_7459,N_6879);
xnor U9423 (N_9423,N_6520,N_6347);
or U9424 (N_9424,N_7835,N_6091);
or U9425 (N_9425,N_7455,N_6616);
nor U9426 (N_9426,N_6511,N_7545);
nor U9427 (N_9427,N_6238,N_7866);
nand U9428 (N_9428,N_7932,N_7176);
nor U9429 (N_9429,N_6597,N_7744);
and U9430 (N_9430,N_7952,N_6585);
xnor U9431 (N_9431,N_6813,N_6066);
nand U9432 (N_9432,N_6946,N_7167);
nand U9433 (N_9433,N_7648,N_7261);
and U9434 (N_9434,N_7889,N_7923);
nor U9435 (N_9435,N_7612,N_7379);
xnor U9436 (N_9436,N_7997,N_7502);
and U9437 (N_9437,N_7197,N_7125);
and U9438 (N_9438,N_7245,N_6953);
nor U9439 (N_9439,N_6719,N_7870);
or U9440 (N_9440,N_7022,N_6386);
nor U9441 (N_9441,N_6400,N_6129);
xor U9442 (N_9442,N_6138,N_6470);
nand U9443 (N_9443,N_6857,N_7462);
or U9444 (N_9444,N_6436,N_7444);
nand U9445 (N_9445,N_7344,N_6569);
or U9446 (N_9446,N_6753,N_6492);
nor U9447 (N_9447,N_6408,N_7212);
nor U9448 (N_9448,N_7266,N_6045);
nand U9449 (N_9449,N_7392,N_7634);
nor U9450 (N_9450,N_7430,N_7721);
or U9451 (N_9451,N_7222,N_6478);
and U9452 (N_9452,N_6814,N_6076);
or U9453 (N_9453,N_6789,N_6585);
nand U9454 (N_9454,N_6871,N_6439);
nor U9455 (N_9455,N_6149,N_6223);
or U9456 (N_9456,N_7457,N_7039);
and U9457 (N_9457,N_6555,N_6597);
nor U9458 (N_9458,N_6555,N_7679);
and U9459 (N_9459,N_7671,N_7223);
and U9460 (N_9460,N_7638,N_6051);
nand U9461 (N_9461,N_7418,N_6600);
and U9462 (N_9462,N_7103,N_6730);
xor U9463 (N_9463,N_6932,N_6234);
nor U9464 (N_9464,N_7770,N_7523);
nand U9465 (N_9465,N_6222,N_7196);
xnor U9466 (N_9466,N_7678,N_7598);
and U9467 (N_9467,N_7694,N_7757);
xnor U9468 (N_9468,N_6939,N_6301);
nor U9469 (N_9469,N_6288,N_6794);
and U9470 (N_9470,N_7054,N_7513);
nor U9471 (N_9471,N_7194,N_6280);
or U9472 (N_9472,N_6925,N_6131);
nand U9473 (N_9473,N_7567,N_7543);
and U9474 (N_9474,N_7137,N_6991);
nor U9475 (N_9475,N_6105,N_7595);
and U9476 (N_9476,N_6947,N_6291);
or U9477 (N_9477,N_6005,N_7647);
nand U9478 (N_9478,N_7008,N_7258);
and U9479 (N_9479,N_6387,N_7845);
or U9480 (N_9480,N_6952,N_6475);
xor U9481 (N_9481,N_6295,N_7278);
xnor U9482 (N_9482,N_7096,N_6014);
or U9483 (N_9483,N_6359,N_7120);
or U9484 (N_9484,N_7209,N_6507);
xnor U9485 (N_9485,N_7879,N_7246);
or U9486 (N_9486,N_7581,N_7766);
xor U9487 (N_9487,N_7193,N_6842);
or U9488 (N_9488,N_6965,N_7378);
xnor U9489 (N_9489,N_6133,N_7575);
nor U9490 (N_9490,N_6468,N_7305);
nand U9491 (N_9491,N_6359,N_6687);
nor U9492 (N_9492,N_6475,N_6336);
nand U9493 (N_9493,N_6950,N_7939);
and U9494 (N_9494,N_7722,N_6970);
or U9495 (N_9495,N_6352,N_7138);
nand U9496 (N_9496,N_6008,N_7918);
nand U9497 (N_9497,N_6302,N_6030);
nand U9498 (N_9498,N_6524,N_6243);
and U9499 (N_9499,N_6717,N_6803);
nor U9500 (N_9500,N_6521,N_7639);
nand U9501 (N_9501,N_7639,N_7794);
and U9502 (N_9502,N_7086,N_7544);
or U9503 (N_9503,N_7801,N_6359);
or U9504 (N_9504,N_7962,N_6955);
or U9505 (N_9505,N_7292,N_6654);
nor U9506 (N_9506,N_6419,N_7089);
xor U9507 (N_9507,N_7450,N_7137);
xnor U9508 (N_9508,N_6240,N_7980);
nor U9509 (N_9509,N_7550,N_7243);
and U9510 (N_9510,N_7282,N_7183);
or U9511 (N_9511,N_6910,N_7504);
and U9512 (N_9512,N_6569,N_7580);
xnor U9513 (N_9513,N_7735,N_7530);
nand U9514 (N_9514,N_7465,N_6579);
nor U9515 (N_9515,N_7807,N_7561);
nand U9516 (N_9516,N_6409,N_6737);
or U9517 (N_9517,N_7812,N_7890);
nor U9518 (N_9518,N_7425,N_7338);
xnor U9519 (N_9519,N_6430,N_7838);
or U9520 (N_9520,N_6041,N_7377);
nand U9521 (N_9521,N_6049,N_7997);
xnor U9522 (N_9522,N_7561,N_6831);
and U9523 (N_9523,N_7430,N_7192);
nor U9524 (N_9524,N_7124,N_6556);
nor U9525 (N_9525,N_6067,N_6196);
nand U9526 (N_9526,N_7812,N_7933);
nand U9527 (N_9527,N_7338,N_7497);
or U9528 (N_9528,N_6667,N_7890);
and U9529 (N_9529,N_7320,N_7139);
or U9530 (N_9530,N_7411,N_7062);
or U9531 (N_9531,N_7018,N_7566);
and U9532 (N_9532,N_6376,N_6262);
nor U9533 (N_9533,N_7737,N_6442);
nor U9534 (N_9534,N_7258,N_7404);
or U9535 (N_9535,N_6236,N_7016);
nand U9536 (N_9536,N_7100,N_7344);
and U9537 (N_9537,N_6182,N_7984);
and U9538 (N_9538,N_6688,N_6744);
xnor U9539 (N_9539,N_6130,N_6306);
nand U9540 (N_9540,N_6889,N_7051);
nor U9541 (N_9541,N_6306,N_6962);
and U9542 (N_9542,N_7947,N_7705);
nor U9543 (N_9543,N_7156,N_6248);
or U9544 (N_9544,N_6590,N_6709);
nand U9545 (N_9545,N_7378,N_7299);
nor U9546 (N_9546,N_6407,N_7961);
and U9547 (N_9547,N_7706,N_7242);
nand U9548 (N_9548,N_6408,N_7671);
nor U9549 (N_9549,N_7108,N_7549);
nand U9550 (N_9550,N_6439,N_6924);
and U9551 (N_9551,N_7628,N_6255);
nor U9552 (N_9552,N_6072,N_7262);
and U9553 (N_9553,N_7489,N_6743);
nand U9554 (N_9554,N_7179,N_7290);
nand U9555 (N_9555,N_7666,N_7730);
or U9556 (N_9556,N_7110,N_7483);
nor U9557 (N_9557,N_7621,N_6457);
and U9558 (N_9558,N_7634,N_7317);
nor U9559 (N_9559,N_7203,N_6857);
nand U9560 (N_9560,N_7840,N_6694);
and U9561 (N_9561,N_6485,N_7541);
nand U9562 (N_9562,N_7670,N_7947);
nor U9563 (N_9563,N_6850,N_6297);
and U9564 (N_9564,N_7587,N_7426);
nand U9565 (N_9565,N_7014,N_7846);
nor U9566 (N_9566,N_7185,N_6953);
nand U9567 (N_9567,N_7983,N_7177);
nor U9568 (N_9568,N_7743,N_6298);
and U9569 (N_9569,N_6772,N_6246);
or U9570 (N_9570,N_7694,N_7645);
and U9571 (N_9571,N_6431,N_6998);
nor U9572 (N_9572,N_6664,N_7725);
or U9573 (N_9573,N_7454,N_6812);
nor U9574 (N_9574,N_6093,N_7631);
nor U9575 (N_9575,N_6463,N_7375);
or U9576 (N_9576,N_6600,N_7107);
or U9577 (N_9577,N_6886,N_7070);
nand U9578 (N_9578,N_7729,N_7872);
or U9579 (N_9579,N_7279,N_6195);
nand U9580 (N_9580,N_6477,N_7062);
nor U9581 (N_9581,N_7198,N_6345);
nand U9582 (N_9582,N_6470,N_7886);
nor U9583 (N_9583,N_6006,N_6727);
nor U9584 (N_9584,N_7187,N_6258);
or U9585 (N_9585,N_7449,N_6361);
nand U9586 (N_9586,N_6163,N_6530);
nor U9587 (N_9587,N_6589,N_7065);
and U9588 (N_9588,N_6325,N_7205);
nor U9589 (N_9589,N_6472,N_6312);
and U9590 (N_9590,N_7081,N_7799);
nor U9591 (N_9591,N_6847,N_7999);
or U9592 (N_9592,N_6373,N_6334);
nor U9593 (N_9593,N_6061,N_7944);
and U9594 (N_9594,N_6790,N_7536);
nor U9595 (N_9595,N_6919,N_7681);
nor U9596 (N_9596,N_6701,N_7632);
nor U9597 (N_9597,N_7294,N_6115);
nand U9598 (N_9598,N_6674,N_7537);
nand U9599 (N_9599,N_7715,N_6002);
xnor U9600 (N_9600,N_7834,N_7592);
or U9601 (N_9601,N_7028,N_7670);
nor U9602 (N_9602,N_7895,N_7181);
nand U9603 (N_9603,N_7694,N_6490);
and U9604 (N_9604,N_6179,N_7389);
nand U9605 (N_9605,N_6396,N_6182);
nor U9606 (N_9606,N_7159,N_6102);
nand U9607 (N_9607,N_6328,N_7168);
and U9608 (N_9608,N_7521,N_6225);
nand U9609 (N_9609,N_6753,N_6979);
xor U9610 (N_9610,N_6506,N_6626);
nor U9611 (N_9611,N_7669,N_6826);
nand U9612 (N_9612,N_6171,N_7031);
nand U9613 (N_9613,N_6217,N_7216);
nand U9614 (N_9614,N_6117,N_7017);
or U9615 (N_9615,N_6574,N_6103);
and U9616 (N_9616,N_6248,N_7476);
and U9617 (N_9617,N_6996,N_6868);
or U9618 (N_9618,N_6062,N_7942);
and U9619 (N_9619,N_6202,N_7858);
or U9620 (N_9620,N_7408,N_6254);
or U9621 (N_9621,N_7307,N_6465);
nor U9622 (N_9622,N_7236,N_7102);
and U9623 (N_9623,N_7755,N_7024);
nor U9624 (N_9624,N_7727,N_7895);
nand U9625 (N_9625,N_7870,N_6439);
nand U9626 (N_9626,N_7238,N_6842);
nand U9627 (N_9627,N_7031,N_7518);
and U9628 (N_9628,N_7311,N_6122);
or U9629 (N_9629,N_7813,N_7910);
nand U9630 (N_9630,N_6069,N_6565);
and U9631 (N_9631,N_7836,N_6345);
or U9632 (N_9632,N_6868,N_6789);
nor U9633 (N_9633,N_7694,N_6092);
or U9634 (N_9634,N_6132,N_7937);
xor U9635 (N_9635,N_6239,N_7644);
nand U9636 (N_9636,N_6849,N_6077);
xor U9637 (N_9637,N_6451,N_6024);
nor U9638 (N_9638,N_7277,N_7739);
nand U9639 (N_9639,N_6873,N_7709);
and U9640 (N_9640,N_7692,N_6348);
nand U9641 (N_9641,N_6803,N_7065);
or U9642 (N_9642,N_6741,N_6156);
nand U9643 (N_9643,N_6207,N_7863);
nand U9644 (N_9644,N_6658,N_7535);
xor U9645 (N_9645,N_7661,N_7497);
nand U9646 (N_9646,N_7570,N_6037);
xnor U9647 (N_9647,N_6390,N_7680);
nor U9648 (N_9648,N_7301,N_6317);
and U9649 (N_9649,N_7580,N_7504);
nor U9650 (N_9650,N_6056,N_7312);
nand U9651 (N_9651,N_7702,N_6092);
and U9652 (N_9652,N_6716,N_7444);
nand U9653 (N_9653,N_7488,N_6856);
or U9654 (N_9654,N_7062,N_6893);
and U9655 (N_9655,N_6700,N_7812);
or U9656 (N_9656,N_7847,N_7875);
nand U9657 (N_9657,N_7037,N_7150);
or U9658 (N_9658,N_7214,N_7485);
xor U9659 (N_9659,N_7791,N_7129);
nor U9660 (N_9660,N_7841,N_7401);
and U9661 (N_9661,N_7508,N_7655);
and U9662 (N_9662,N_7257,N_6906);
and U9663 (N_9663,N_6797,N_7941);
and U9664 (N_9664,N_7678,N_7548);
and U9665 (N_9665,N_7349,N_6887);
and U9666 (N_9666,N_7739,N_7655);
nor U9667 (N_9667,N_6000,N_7107);
and U9668 (N_9668,N_6417,N_6198);
or U9669 (N_9669,N_6162,N_6732);
nand U9670 (N_9670,N_7116,N_6456);
nor U9671 (N_9671,N_6127,N_6711);
and U9672 (N_9672,N_7281,N_7302);
nand U9673 (N_9673,N_6970,N_6282);
nand U9674 (N_9674,N_6902,N_6514);
and U9675 (N_9675,N_7696,N_7916);
nor U9676 (N_9676,N_6093,N_7395);
or U9677 (N_9677,N_7311,N_6808);
and U9678 (N_9678,N_6283,N_7378);
xnor U9679 (N_9679,N_6518,N_6636);
nand U9680 (N_9680,N_6946,N_6505);
and U9681 (N_9681,N_6697,N_6091);
or U9682 (N_9682,N_7376,N_7522);
nor U9683 (N_9683,N_6038,N_7248);
nor U9684 (N_9684,N_6669,N_7496);
xor U9685 (N_9685,N_7139,N_6423);
xnor U9686 (N_9686,N_6328,N_7929);
and U9687 (N_9687,N_6229,N_6279);
nand U9688 (N_9688,N_7963,N_6087);
and U9689 (N_9689,N_7605,N_6333);
or U9690 (N_9690,N_6039,N_7814);
and U9691 (N_9691,N_6922,N_7212);
and U9692 (N_9692,N_7886,N_6845);
nand U9693 (N_9693,N_6547,N_7327);
nand U9694 (N_9694,N_6649,N_6939);
xnor U9695 (N_9695,N_7040,N_7311);
nor U9696 (N_9696,N_7525,N_6033);
or U9697 (N_9697,N_6446,N_6889);
nand U9698 (N_9698,N_7572,N_6135);
nor U9699 (N_9699,N_7631,N_6944);
nor U9700 (N_9700,N_7624,N_6468);
nand U9701 (N_9701,N_6318,N_7613);
and U9702 (N_9702,N_6641,N_6663);
or U9703 (N_9703,N_7063,N_7654);
or U9704 (N_9704,N_7691,N_7044);
and U9705 (N_9705,N_6915,N_6855);
or U9706 (N_9706,N_7377,N_6168);
and U9707 (N_9707,N_7919,N_6235);
nor U9708 (N_9708,N_6463,N_7040);
nand U9709 (N_9709,N_7631,N_7868);
and U9710 (N_9710,N_7341,N_7080);
nand U9711 (N_9711,N_6708,N_7122);
nor U9712 (N_9712,N_6347,N_6900);
nor U9713 (N_9713,N_7669,N_7763);
and U9714 (N_9714,N_6518,N_6970);
nor U9715 (N_9715,N_7535,N_6541);
or U9716 (N_9716,N_6056,N_7313);
nand U9717 (N_9717,N_6637,N_7992);
and U9718 (N_9718,N_6590,N_7212);
nand U9719 (N_9719,N_7380,N_6009);
or U9720 (N_9720,N_7941,N_6111);
nand U9721 (N_9721,N_6337,N_6755);
xnor U9722 (N_9722,N_7580,N_7417);
nor U9723 (N_9723,N_7545,N_7222);
and U9724 (N_9724,N_7643,N_7541);
nand U9725 (N_9725,N_6978,N_6301);
nor U9726 (N_9726,N_6991,N_7518);
nand U9727 (N_9727,N_7219,N_7795);
or U9728 (N_9728,N_6380,N_7204);
nor U9729 (N_9729,N_7585,N_7124);
and U9730 (N_9730,N_6567,N_7024);
or U9731 (N_9731,N_6887,N_7563);
or U9732 (N_9732,N_6137,N_6042);
nand U9733 (N_9733,N_7913,N_6442);
nand U9734 (N_9734,N_7133,N_6140);
or U9735 (N_9735,N_7641,N_7224);
nand U9736 (N_9736,N_6659,N_6082);
nor U9737 (N_9737,N_7308,N_7466);
nand U9738 (N_9738,N_6383,N_6399);
nor U9739 (N_9739,N_7671,N_6927);
xor U9740 (N_9740,N_6205,N_7770);
or U9741 (N_9741,N_6154,N_7526);
nor U9742 (N_9742,N_7658,N_7813);
and U9743 (N_9743,N_7144,N_6015);
nor U9744 (N_9744,N_6900,N_6910);
and U9745 (N_9745,N_6297,N_7445);
or U9746 (N_9746,N_6543,N_7928);
and U9747 (N_9747,N_7002,N_7371);
and U9748 (N_9748,N_6682,N_7352);
nor U9749 (N_9749,N_7522,N_7059);
nor U9750 (N_9750,N_7317,N_7222);
xnor U9751 (N_9751,N_6985,N_7349);
nand U9752 (N_9752,N_7914,N_6455);
xnor U9753 (N_9753,N_7327,N_6205);
and U9754 (N_9754,N_6992,N_6604);
xor U9755 (N_9755,N_7130,N_7647);
and U9756 (N_9756,N_7361,N_7430);
and U9757 (N_9757,N_7228,N_6184);
nor U9758 (N_9758,N_7953,N_6570);
or U9759 (N_9759,N_7964,N_6375);
nor U9760 (N_9760,N_7451,N_6150);
or U9761 (N_9761,N_7444,N_7579);
and U9762 (N_9762,N_7893,N_6272);
or U9763 (N_9763,N_6382,N_6325);
and U9764 (N_9764,N_7930,N_6839);
xnor U9765 (N_9765,N_6230,N_7518);
and U9766 (N_9766,N_6778,N_6488);
or U9767 (N_9767,N_6506,N_7104);
or U9768 (N_9768,N_7852,N_6361);
or U9769 (N_9769,N_7859,N_7648);
nor U9770 (N_9770,N_6116,N_7338);
nor U9771 (N_9771,N_6725,N_6871);
and U9772 (N_9772,N_6929,N_6042);
and U9773 (N_9773,N_7932,N_6393);
and U9774 (N_9774,N_7857,N_7493);
nand U9775 (N_9775,N_6019,N_7333);
or U9776 (N_9776,N_7952,N_7010);
nand U9777 (N_9777,N_6560,N_6071);
nor U9778 (N_9778,N_6299,N_7064);
nor U9779 (N_9779,N_6398,N_7354);
or U9780 (N_9780,N_6039,N_6560);
nand U9781 (N_9781,N_7420,N_7465);
nor U9782 (N_9782,N_7083,N_6669);
nor U9783 (N_9783,N_6674,N_7802);
and U9784 (N_9784,N_7181,N_7883);
or U9785 (N_9785,N_6415,N_6981);
and U9786 (N_9786,N_7215,N_6476);
xor U9787 (N_9787,N_7604,N_7448);
and U9788 (N_9788,N_6177,N_7158);
nor U9789 (N_9789,N_6284,N_7020);
nor U9790 (N_9790,N_6645,N_7583);
and U9791 (N_9791,N_6032,N_7932);
or U9792 (N_9792,N_7455,N_7107);
and U9793 (N_9793,N_6937,N_7270);
nand U9794 (N_9794,N_7880,N_6212);
and U9795 (N_9795,N_6342,N_6660);
nand U9796 (N_9796,N_7869,N_6280);
nor U9797 (N_9797,N_6138,N_6368);
nor U9798 (N_9798,N_7362,N_7258);
and U9799 (N_9799,N_7879,N_7747);
nor U9800 (N_9800,N_6562,N_6220);
or U9801 (N_9801,N_7812,N_6077);
nand U9802 (N_9802,N_7566,N_7157);
nor U9803 (N_9803,N_6273,N_6950);
and U9804 (N_9804,N_6571,N_7286);
nor U9805 (N_9805,N_7992,N_6143);
nand U9806 (N_9806,N_7650,N_7248);
and U9807 (N_9807,N_7931,N_6331);
or U9808 (N_9808,N_6009,N_7750);
nand U9809 (N_9809,N_6356,N_7870);
xor U9810 (N_9810,N_7390,N_7687);
or U9811 (N_9811,N_7477,N_7303);
or U9812 (N_9812,N_6837,N_7219);
nor U9813 (N_9813,N_6538,N_7142);
or U9814 (N_9814,N_6645,N_6814);
or U9815 (N_9815,N_7768,N_7824);
or U9816 (N_9816,N_7695,N_6956);
nand U9817 (N_9817,N_6828,N_7150);
or U9818 (N_9818,N_6000,N_6404);
nor U9819 (N_9819,N_7735,N_7131);
nand U9820 (N_9820,N_7941,N_7142);
nand U9821 (N_9821,N_7942,N_7852);
or U9822 (N_9822,N_7340,N_7989);
nor U9823 (N_9823,N_6757,N_6366);
and U9824 (N_9824,N_7003,N_6558);
and U9825 (N_9825,N_6552,N_6340);
nand U9826 (N_9826,N_6401,N_7026);
nand U9827 (N_9827,N_7517,N_7197);
nand U9828 (N_9828,N_6261,N_7565);
or U9829 (N_9829,N_7596,N_7540);
or U9830 (N_9830,N_7764,N_6722);
nor U9831 (N_9831,N_7602,N_6294);
or U9832 (N_9832,N_7758,N_6052);
or U9833 (N_9833,N_7583,N_7813);
nand U9834 (N_9834,N_7224,N_6489);
nand U9835 (N_9835,N_7982,N_6649);
or U9836 (N_9836,N_6488,N_6436);
nand U9837 (N_9837,N_7519,N_6122);
nand U9838 (N_9838,N_7955,N_7494);
xor U9839 (N_9839,N_7677,N_6891);
nand U9840 (N_9840,N_6623,N_6461);
and U9841 (N_9841,N_6795,N_6410);
or U9842 (N_9842,N_7103,N_7841);
nand U9843 (N_9843,N_6258,N_6084);
nor U9844 (N_9844,N_6667,N_6162);
nor U9845 (N_9845,N_6853,N_7228);
or U9846 (N_9846,N_7734,N_7353);
or U9847 (N_9847,N_7560,N_6661);
nor U9848 (N_9848,N_7878,N_7233);
or U9849 (N_9849,N_6138,N_7237);
nand U9850 (N_9850,N_6873,N_7426);
or U9851 (N_9851,N_7827,N_6543);
or U9852 (N_9852,N_6200,N_6463);
xnor U9853 (N_9853,N_7807,N_6268);
xor U9854 (N_9854,N_7274,N_6417);
or U9855 (N_9855,N_7849,N_6172);
nand U9856 (N_9856,N_6941,N_6899);
nor U9857 (N_9857,N_7804,N_6659);
or U9858 (N_9858,N_7110,N_6085);
and U9859 (N_9859,N_7849,N_7804);
nand U9860 (N_9860,N_6700,N_7074);
nor U9861 (N_9861,N_6707,N_6160);
or U9862 (N_9862,N_7360,N_7111);
nand U9863 (N_9863,N_7086,N_6618);
or U9864 (N_9864,N_6258,N_6210);
nor U9865 (N_9865,N_7989,N_6799);
nor U9866 (N_9866,N_6014,N_6490);
and U9867 (N_9867,N_6400,N_7025);
or U9868 (N_9868,N_7214,N_6824);
or U9869 (N_9869,N_7598,N_7226);
xnor U9870 (N_9870,N_7935,N_6348);
nand U9871 (N_9871,N_6943,N_7164);
xor U9872 (N_9872,N_6490,N_7595);
nor U9873 (N_9873,N_6107,N_7457);
xor U9874 (N_9874,N_6330,N_7303);
nor U9875 (N_9875,N_7520,N_6474);
and U9876 (N_9876,N_7024,N_6704);
and U9877 (N_9877,N_7424,N_6585);
and U9878 (N_9878,N_6740,N_6863);
or U9879 (N_9879,N_7459,N_6374);
and U9880 (N_9880,N_6184,N_6762);
nand U9881 (N_9881,N_7115,N_6243);
nor U9882 (N_9882,N_7173,N_7135);
nor U9883 (N_9883,N_7999,N_7067);
nand U9884 (N_9884,N_7218,N_6265);
nor U9885 (N_9885,N_6516,N_7730);
and U9886 (N_9886,N_6953,N_6416);
or U9887 (N_9887,N_6294,N_7746);
or U9888 (N_9888,N_6028,N_7418);
and U9889 (N_9889,N_6462,N_7218);
nand U9890 (N_9890,N_6179,N_7386);
and U9891 (N_9891,N_6521,N_7575);
xor U9892 (N_9892,N_6195,N_6553);
and U9893 (N_9893,N_6500,N_7794);
nor U9894 (N_9894,N_6796,N_7644);
or U9895 (N_9895,N_6587,N_6220);
and U9896 (N_9896,N_7359,N_7285);
and U9897 (N_9897,N_7222,N_7743);
nand U9898 (N_9898,N_6212,N_7906);
nand U9899 (N_9899,N_6922,N_7740);
and U9900 (N_9900,N_7077,N_6117);
xnor U9901 (N_9901,N_7904,N_7206);
or U9902 (N_9902,N_7940,N_7177);
nor U9903 (N_9903,N_6626,N_7096);
or U9904 (N_9904,N_7729,N_6645);
nand U9905 (N_9905,N_7637,N_7587);
nand U9906 (N_9906,N_7395,N_6679);
nand U9907 (N_9907,N_7300,N_7776);
nor U9908 (N_9908,N_7038,N_7228);
nor U9909 (N_9909,N_7114,N_6271);
nor U9910 (N_9910,N_6325,N_7923);
and U9911 (N_9911,N_7790,N_7671);
and U9912 (N_9912,N_7424,N_7775);
nor U9913 (N_9913,N_7463,N_7555);
and U9914 (N_9914,N_6447,N_6849);
or U9915 (N_9915,N_6340,N_6229);
and U9916 (N_9916,N_7944,N_7778);
nor U9917 (N_9917,N_6929,N_6972);
or U9918 (N_9918,N_7651,N_6797);
nor U9919 (N_9919,N_6466,N_7269);
or U9920 (N_9920,N_7950,N_6197);
or U9921 (N_9921,N_7397,N_6948);
or U9922 (N_9922,N_7187,N_6116);
nor U9923 (N_9923,N_6052,N_6653);
xnor U9924 (N_9924,N_7297,N_6126);
and U9925 (N_9925,N_7932,N_6273);
or U9926 (N_9926,N_6173,N_7622);
or U9927 (N_9927,N_6384,N_6666);
xnor U9928 (N_9928,N_6796,N_6938);
nand U9929 (N_9929,N_6068,N_7969);
xnor U9930 (N_9930,N_7485,N_6425);
or U9931 (N_9931,N_7017,N_6406);
and U9932 (N_9932,N_7048,N_6201);
xor U9933 (N_9933,N_6188,N_6369);
or U9934 (N_9934,N_7840,N_6184);
nor U9935 (N_9935,N_7436,N_6941);
nand U9936 (N_9936,N_7940,N_7049);
nor U9937 (N_9937,N_7176,N_7085);
nand U9938 (N_9938,N_7723,N_6139);
and U9939 (N_9939,N_7859,N_7091);
nor U9940 (N_9940,N_7822,N_6844);
nand U9941 (N_9941,N_6549,N_7235);
nor U9942 (N_9942,N_6107,N_7759);
and U9943 (N_9943,N_7090,N_6763);
and U9944 (N_9944,N_7467,N_7607);
nor U9945 (N_9945,N_7822,N_7693);
and U9946 (N_9946,N_6271,N_6911);
or U9947 (N_9947,N_7213,N_7233);
nand U9948 (N_9948,N_6651,N_7457);
nand U9949 (N_9949,N_7474,N_6516);
and U9950 (N_9950,N_6747,N_7847);
xnor U9951 (N_9951,N_6708,N_7036);
nor U9952 (N_9952,N_6513,N_6484);
or U9953 (N_9953,N_6667,N_7336);
nor U9954 (N_9954,N_7061,N_7709);
nand U9955 (N_9955,N_7366,N_7618);
and U9956 (N_9956,N_6114,N_6746);
nor U9957 (N_9957,N_7163,N_7190);
or U9958 (N_9958,N_7937,N_6170);
or U9959 (N_9959,N_7245,N_6334);
nor U9960 (N_9960,N_7077,N_6930);
xor U9961 (N_9961,N_7301,N_7914);
or U9962 (N_9962,N_7279,N_7499);
xor U9963 (N_9963,N_7036,N_7210);
or U9964 (N_9964,N_7268,N_7668);
nor U9965 (N_9965,N_6506,N_7468);
nand U9966 (N_9966,N_6558,N_6600);
nand U9967 (N_9967,N_6297,N_7220);
nor U9968 (N_9968,N_7319,N_6163);
xor U9969 (N_9969,N_6126,N_7160);
and U9970 (N_9970,N_6729,N_6711);
nor U9971 (N_9971,N_7381,N_7314);
or U9972 (N_9972,N_7656,N_7447);
or U9973 (N_9973,N_6856,N_6662);
xor U9974 (N_9974,N_6100,N_7486);
nand U9975 (N_9975,N_6922,N_6092);
or U9976 (N_9976,N_7987,N_7640);
nand U9977 (N_9977,N_7583,N_6982);
nand U9978 (N_9978,N_7442,N_7615);
nor U9979 (N_9979,N_6056,N_6523);
nor U9980 (N_9980,N_7886,N_7366);
nor U9981 (N_9981,N_6863,N_6744);
xnor U9982 (N_9982,N_6724,N_6822);
and U9983 (N_9983,N_7142,N_6125);
xor U9984 (N_9984,N_7315,N_6833);
nor U9985 (N_9985,N_7239,N_7624);
nand U9986 (N_9986,N_6034,N_6143);
xor U9987 (N_9987,N_7721,N_7738);
or U9988 (N_9988,N_6065,N_6181);
or U9989 (N_9989,N_7731,N_6439);
and U9990 (N_9990,N_7723,N_7654);
and U9991 (N_9991,N_6950,N_6436);
and U9992 (N_9992,N_7653,N_7674);
xnor U9993 (N_9993,N_6349,N_7434);
or U9994 (N_9994,N_6258,N_7070);
or U9995 (N_9995,N_7132,N_6130);
nor U9996 (N_9996,N_6051,N_6198);
nand U9997 (N_9997,N_6406,N_6730);
nand U9998 (N_9998,N_6897,N_7797);
and U9999 (N_9999,N_6339,N_6166);
xnor U10000 (N_10000,N_9232,N_8073);
xnor U10001 (N_10001,N_8079,N_9551);
and U10002 (N_10002,N_8166,N_8267);
and U10003 (N_10003,N_9577,N_9279);
nor U10004 (N_10004,N_9800,N_8493);
nor U10005 (N_10005,N_8984,N_8829);
nand U10006 (N_10006,N_9376,N_8476);
xnor U10007 (N_10007,N_8193,N_8531);
nand U10008 (N_10008,N_9737,N_9256);
xnor U10009 (N_10009,N_8860,N_8249);
or U10010 (N_10010,N_9280,N_9424);
nand U10011 (N_10011,N_9168,N_9674);
and U10012 (N_10012,N_8097,N_8845);
nor U10013 (N_10013,N_9982,N_9564);
and U10014 (N_10014,N_8184,N_8220);
and U10015 (N_10015,N_9409,N_8540);
or U10016 (N_10016,N_8530,N_9334);
and U10017 (N_10017,N_8289,N_8551);
or U10018 (N_10018,N_8924,N_9683);
nor U10019 (N_10019,N_8115,N_8585);
nor U10020 (N_10020,N_9178,N_9948);
or U10021 (N_10021,N_9174,N_9297);
and U10022 (N_10022,N_9228,N_8396);
and U10023 (N_10023,N_8251,N_9151);
and U10024 (N_10024,N_9557,N_9816);
nand U10025 (N_10025,N_9937,N_8228);
xor U10026 (N_10026,N_8576,N_8254);
nand U10027 (N_10027,N_8809,N_8794);
and U10028 (N_10028,N_9540,N_9497);
and U10029 (N_10029,N_8415,N_8666);
xnor U10030 (N_10030,N_9131,N_8606);
or U10031 (N_10031,N_9111,N_9341);
nor U10032 (N_10032,N_9701,N_8838);
nand U10033 (N_10033,N_9296,N_8726);
nor U10034 (N_10034,N_8188,N_8769);
and U10035 (N_10035,N_8474,N_9020);
and U10036 (N_10036,N_8933,N_8496);
nand U10037 (N_10037,N_8930,N_9299);
and U10038 (N_10038,N_8620,N_8003);
xor U10039 (N_10039,N_8385,N_9668);
or U10040 (N_10040,N_8944,N_9696);
or U10041 (N_10041,N_9861,N_8679);
or U10042 (N_10042,N_8376,N_8755);
and U10043 (N_10043,N_9226,N_8298);
nand U10044 (N_10044,N_8871,N_9153);
or U10045 (N_10045,N_9294,N_8028);
nand U10046 (N_10046,N_9543,N_8525);
or U10047 (N_10047,N_8767,N_9118);
and U10048 (N_10048,N_8813,N_9849);
nand U10049 (N_10049,N_8368,N_8138);
nor U10050 (N_10050,N_8872,N_8114);
nand U10051 (N_10051,N_9927,N_8418);
nand U10052 (N_10052,N_8405,N_9378);
xnor U10053 (N_10053,N_9621,N_9330);
nor U10054 (N_10054,N_9824,N_9912);
xor U10055 (N_10055,N_8817,N_8909);
xor U10056 (N_10056,N_8294,N_8102);
nor U10057 (N_10057,N_9063,N_9522);
and U10058 (N_10058,N_9004,N_8070);
and U10059 (N_10059,N_9440,N_9198);
nor U10060 (N_10060,N_8692,N_8482);
and U10061 (N_10061,N_8049,N_8314);
nor U10062 (N_10062,N_8043,N_9900);
nand U10063 (N_10063,N_8619,N_9850);
nand U10064 (N_10064,N_8963,N_8194);
and U10065 (N_10065,N_9333,N_9976);
nor U10066 (N_10066,N_8002,N_8554);
nor U10067 (N_10067,N_9753,N_8222);
nand U10068 (N_10068,N_8532,N_8015);
or U10069 (N_10069,N_9902,N_9887);
or U10070 (N_10070,N_8216,N_9726);
nand U10071 (N_10071,N_9391,N_8051);
and U10072 (N_10072,N_9840,N_9618);
and U10073 (N_10073,N_9767,N_8107);
nand U10074 (N_10074,N_9157,N_9066);
xnor U10075 (N_10075,N_8357,N_8912);
nand U10076 (N_10076,N_9782,N_8489);
xnor U10077 (N_10077,N_8142,N_8446);
nor U10078 (N_10078,N_9370,N_9936);
or U10079 (N_10079,N_8127,N_9244);
or U10080 (N_10080,N_8130,N_8853);
nor U10081 (N_10081,N_9970,N_8006);
and U10082 (N_10082,N_9284,N_9605);
or U10083 (N_10083,N_9471,N_8318);
and U10084 (N_10084,N_8290,N_9302);
or U10085 (N_10085,N_9991,N_9710);
nor U10086 (N_10086,N_8875,N_9636);
nand U10087 (N_10087,N_9094,N_8940);
and U10088 (N_10088,N_8161,N_8306);
and U10089 (N_10089,N_8144,N_9494);
and U10090 (N_10090,N_9595,N_8371);
and U10091 (N_10091,N_9435,N_9030);
nor U10092 (N_10092,N_8750,N_8126);
and U10093 (N_10093,N_8334,N_9882);
and U10094 (N_10094,N_9629,N_9007);
xor U10095 (N_10095,N_8310,N_8305);
nand U10096 (N_10096,N_8041,N_8517);
nand U10097 (N_10097,N_8694,N_8480);
nand U10098 (N_10098,N_9730,N_9940);
nor U10099 (N_10099,N_8000,N_8046);
nor U10100 (N_10100,N_9672,N_8091);
nand U10101 (N_10101,N_9310,N_8100);
nor U10102 (N_10102,N_9291,N_9585);
and U10103 (N_10103,N_9687,N_9868);
or U10104 (N_10104,N_8815,N_9445);
nand U10105 (N_10105,N_8658,N_8843);
nand U10106 (N_10106,N_9798,N_9345);
and U10107 (N_10107,N_9758,N_8200);
nand U10108 (N_10108,N_9775,N_9285);
and U10109 (N_10109,N_8240,N_9653);
and U10110 (N_10110,N_8259,N_8779);
xor U10111 (N_10111,N_8004,N_9537);
and U10112 (N_10112,N_8141,N_8708);
xor U10113 (N_10113,N_9593,N_8934);
nor U10114 (N_10114,N_8938,N_9448);
xor U10115 (N_10115,N_8967,N_9073);
and U10116 (N_10116,N_8656,N_8491);
or U10117 (N_10117,N_9721,N_9200);
nand U10118 (N_10118,N_9490,N_8822);
nand U10119 (N_10119,N_8348,N_8646);
xnor U10120 (N_10120,N_9881,N_8430);
and U10121 (N_10121,N_9960,N_9132);
and U10122 (N_10122,N_9432,N_8440);
nand U10123 (N_10123,N_8659,N_9259);
nor U10124 (N_10124,N_9112,N_8602);
xor U10125 (N_10125,N_9086,N_8987);
and U10126 (N_10126,N_8980,N_9312);
and U10127 (N_10127,N_8673,N_8895);
and U10128 (N_10128,N_8660,N_9565);
or U10129 (N_10129,N_8899,N_8283);
nor U10130 (N_10130,N_8927,N_8326);
nand U10131 (N_10131,N_9590,N_8614);
and U10132 (N_10132,N_8235,N_8607);
and U10133 (N_10133,N_9155,N_9804);
and U10134 (N_10134,N_8529,N_9688);
nor U10135 (N_10135,N_8390,N_9139);
or U10136 (N_10136,N_8771,N_9644);
nand U10137 (N_10137,N_9757,N_8150);
nor U10138 (N_10138,N_9603,N_8324);
nor U10139 (N_10139,N_8723,N_8662);
xnor U10140 (N_10140,N_8377,N_9371);
and U10141 (N_10141,N_9029,N_8502);
or U10142 (N_10142,N_8080,N_9837);
or U10143 (N_10143,N_8902,N_9984);
and U10144 (N_10144,N_9365,N_8883);
or U10145 (N_10145,N_8147,N_9171);
and U10146 (N_10146,N_8103,N_8788);
nor U10147 (N_10147,N_9179,N_8175);
and U10148 (N_10148,N_9495,N_9344);
or U10149 (N_10149,N_9260,N_9649);
and U10150 (N_10150,N_9985,N_9517);
and U10151 (N_10151,N_8083,N_8626);
nand U10152 (N_10152,N_9486,N_8499);
nand U10153 (N_10153,N_9449,N_8317);
and U10154 (N_10154,N_9229,N_9324);
nor U10155 (N_10155,N_8510,N_9931);
or U10156 (N_10156,N_8219,N_8189);
and U10157 (N_10157,N_9361,N_8885);
and U10158 (N_10158,N_9170,N_9119);
nor U10159 (N_10159,N_8805,N_9212);
nor U10160 (N_10160,N_8842,N_9165);
and U10161 (N_10161,N_9305,N_9160);
xnor U10162 (N_10162,N_9142,N_8935);
nand U10163 (N_10163,N_9476,N_9813);
xnor U10164 (N_10164,N_8279,N_9508);
or U10165 (N_10165,N_9182,N_8155);
nor U10166 (N_10166,N_9113,N_9193);
nand U10167 (N_10167,N_8492,N_8281);
nand U10168 (N_10168,N_8498,N_8803);
xor U10169 (N_10169,N_9809,N_8878);
xor U10170 (N_10170,N_8774,N_8678);
nor U10171 (N_10171,N_8461,N_9999);
or U10172 (N_10172,N_8449,N_8854);
nand U10173 (N_10173,N_8687,N_9414);
and U10174 (N_10174,N_9582,N_8722);
nand U10175 (N_10175,N_8071,N_8037);
nand U10176 (N_10176,N_8896,N_9971);
nand U10177 (N_10177,N_8343,N_8426);
or U10178 (N_10178,N_8158,N_9068);
nand U10179 (N_10179,N_9675,N_8462);
and U10180 (N_10180,N_9574,N_9834);
nor U10181 (N_10181,N_8411,N_8918);
and U10182 (N_10182,N_9320,N_8686);
and U10183 (N_10183,N_8017,N_8557);
and U10184 (N_10184,N_9853,N_9203);
nand U10185 (N_10185,N_9908,N_9944);
nand U10186 (N_10186,N_9829,N_8255);
and U10187 (N_10187,N_9434,N_9657);
and U10188 (N_10188,N_8680,N_8555);
nand U10189 (N_10189,N_9921,N_9247);
or U10190 (N_10190,N_8024,N_8572);
nand U10191 (N_10191,N_8773,N_8455);
and U10192 (N_10192,N_9958,N_9705);
and U10193 (N_10193,N_9707,N_9941);
nor U10194 (N_10194,N_9403,N_9552);
xor U10195 (N_10195,N_9271,N_9390);
xnor U10196 (N_10196,N_8316,N_9006);
xor U10197 (N_10197,N_9472,N_8976);
and U10198 (N_10198,N_8647,N_8431);
and U10199 (N_10199,N_9520,N_9389);
and U10200 (N_10200,N_9453,N_8231);
and U10201 (N_10201,N_9755,N_9116);
and U10202 (N_10202,N_8218,N_8888);
or U10203 (N_10203,N_8820,N_9347);
nand U10204 (N_10204,N_8970,N_9231);
nand U10205 (N_10205,N_9901,N_8047);
nor U10206 (N_10206,N_8981,N_8772);
xor U10207 (N_10207,N_8151,N_8284);
and U10208 (N_10208,N_8579,N_9515);
nor U10209 (N_10209,N_8033,N_9114);
and U10210 (N_10210,N_9134,N_9161);
or U10211 (N_10211,N_8471,N_9778);
and U10212 (N_10212,N_9790,N_9196);
xor U10213 (N_10213,N_8761,N_9567);
nor U10214 (N_10214,N_8969,N_8404);
xnor U10215 (N_10215,N_9092,N_8867);
nand U10216 (N_10216,N_9780,N_9919);
and U10217 (N_10217,N_8459,N_9872);
and U10218 (N_10218,N_9062,N_9120);
nand U10219 (N_10219,N_8746,N_9052);
and U10220 (N_10220,N_8238,N_8401);
nor U10221 (N_10221,N_8470,N_8710);
nor U10222 (N_10222,N_9933,N_9017);
xor U10223 (N_10223,N_9623,N_8355);
nand U10224 (N_10224,N_9925,N_8148);
and U10225 (N_10225,N_8855,N_9768);
or U10226 (N_10226,N_9355,N_8389);
or U10227 (N_10227,N_8263,N_8738);
nor U10228 (N_10228,N_9444,N_8353);
and U10229 (N_10229,N_9709,N_9127);
and U10230 (N_10230,N_9541,N_8745);
and U10231 (N_10231,N_9394,N_8162);
or U10232 (N_10232,N_8973,N_9663);
nand U10233 (N_10233,N_8029,N_9144);
or U10234 (N_10234,N_8668,N_9000);
nor U10235 (N_10235,N_9963,N_8342);
xor U10236 (N_10236,N_9906,N_8835);
or U10237 (N_10237,N_9743,N_8986);
or U10238 (N_10238,N_9505,N_9398);
or U10239 (N_10239,N_8756,N_8565);
nor U10240 (N_10240,N_9993,N_9034);
or U10241 (N_10241,N_9996,N_8580);
or U10242 (N_10242,N_8562,N_8018);
nor U10243 (N_10243,N_8699,N_9686);
nor U10244 (N_10244,N_9863,N_9162);
and U10245 (N_10245,N_8582,N_8282);
and U10246 (N_10246,N_8475,N_8950);
or U10247 (N_10247,N_9599,N_8567);
or U10248 (N_10248,N_8055,N_9479);
or U10249 (N_10249,N_9379,N_9706);
nand U10250 (N_10250,N_8995,N_9124);
nor U10251 (N_10251,N_9640,N_9402);
nor U10252 (N_10252,N_9465,N_8358);
and U10253 (N_10253,N_8329,N_8864);
or U10254 (N_10254,N_9416,N_8721);
nor U10255 (N_10255,N_8250,N_8672);
or U10256 (N_10256,N_9968,N_8543);
and U10257 (N_10257,N_9581,N_9817);
nand U10258 (N_10258,N_8208,N_9292);
or U10259 (N_10259,N_8395,N_9147);
nand U10260 (N_10260,N_9136,N_9087);
nor U10261 (N_10261,N_8074,N_8793);
and U10262 (N_10262,N_9833,N_9723);
nand U10263 (N_10263,N_8364,N_8365);
or U10264 (N_10264,N_9374,N_8372);
nor U10265 (N_10265,N_8583,N_9571);
and U10266 (N_10266,N_8876,N_9869);
or U10267 (N_10267,N_8889,N_9239);
or U10268 (N_10268,N_9533,N_8192);
nand U10269 (N_10269,N_8067,N_8236);
or U10270 (N_10270,N_8176,N_9454);
nor U10271 (N_10271,N_9372,N_8122);
xor U10272 (N_10272,N_9519,N_9346);
and U10273 (N_10273,N_8439,N_8032);
nor U10274 (N_10274,N_8123,N_9255);
nor U10275 (N_10275,N_8728,N_8108);
and U10276 (N_10276,N_8951,N_8782);
nor U10277 (N_10277,N_9488,N_8592);
nor U10278 (N_10278,N_9484,N_9481);
nand U10279 (N_10279,N_9439,N_8088);
and U10280 (N_10280,N_8713,N_9351);
nor U10281 (N_10281,N_8961,N_9547);
xor U10282 (N_10282,N_8752,N_8907);
nor U10283 (N_10283,N_9612,N_8052);
nand U10284 (N_10284,N_8790,N_8514);
and U10285 (N_10285,N_9295,N_9306);
nor U10286 (N_10286,N_9048,N_8383);
or U10287 (N_10287,N_9878,N_9895);
nand U10288 (N_10288,N_9288,N_9383);
or U10289 (N_10289,N_9679,N_9332);
and U10290 (N_10290,N_9792,N_8800);
nand U10291 (N_10291,N_8109,N_9652);
or U10292 (N_10292,N_8847,N_8941);
nand U10293 (N_10293,N_9915,N_9822);
and U10294 (N_10294,N_9635,N_9560);
nand U10295 (N_10295,N_9219,N_8998);
or U10296 (N_10296,N_8783,N_8558);
nand U10297 (N_10297,N_8273,N_9880);
and U10298 (N_10298,N_8915,N_9032);
and U10299 (N_10299,N_8214,N_9385);
or U10300 (N_10300,N_9965,N_8164);
or U10301 (N_10301,N_8432,N_9138);
and U10302 (N_10302,N_8437,N_9380);
nor U10303 (N_10303,N_8541,N_9311);
and U10304 (N_10304,N_8393,N_8098);
or U10305 (N_10305,N_8863,N_8163);
and U10306 (N_10306,N_8749,N_8295);
or U10307 (N_10307,N_8609,N_9797);
nand U10308 (N_10308,N_9217,N_8747);
or U10309 (N_10309,N_9410,N_8865);
xor U10310 (N_10310,N_8293,N_9399);
or U10311 (N_10311,N_9015,N_9716);
and U10312 (N_10312,N_8419,N_9067);
or U10313 (N_10313,N_9734,N_9423);
nor U10314 (N_10314,N_8438,N_9317);
or U10315 (N_10315,N_8586,N_8792);
and U10316 (N_10316,N_9069,N_8488);
and U10317 (N_10317,N_9518,N_9002);
and U10318 (N_10318,N_9761,N_8827);
xor U10319 (N_10319,N_9521,N_8374);
and U10320 (N_10320,N_8160,N_8593);
or U10321 (N_10321,N_8485,N_8204);
nor U10322 (N_10322,N_9724,N_8511);
nor U10323 (N_10323,N_8441,N_9406);
or U10324 (N_10324,N_9387,N_9617);
nand U10325 (N_10325,N_8178,N_8223);
or U10326 (N_10326,N_8801,N_8149);
or U10327 (N_10327,N_8191,N_8691);
nor U10328 (N_10328,N_9988,N_9854);
xor U10329 (N_10329,N_8020,N_9149);
and U10330 (N_10330,N_8784,N_8139);
xnor U10331 (N_10331,N_9916,N_9877);
and U10332 (N_10332,N_8920,N_8552);
nand U10333 (N_10333,N_8023,N_8806);
nor U10334 (N_10334,N_9690,N_8739);
xor U10335 (N_10335,N_8914,N_9539);
nand U10336 (N_10336,N_9923,N_9172);
or U10337 (N_10337,N_9081,N_9749);
nand U10338 (N_10338,N_8605,N_9667);
and U10339 (N_10339,N_8137,N_8604);
or U10340 (N_10340,N_9265,N_9751);
nand U10341 (N_10341,N_9846,N_9729);
nand U10342 (N_10342,N_8524,N_9273);
nand U10343 (N_10343,N_9818,N_8380);
or U10344 (N_10344,N_9430,N_9061);
and U10345 (N_10345,N_9754,N_9562);
nor U10346 (N_10346,N_8265,N_8416);
and U10347 (N_10347,N_8113,N_8087);
nor U10348 (N_10348,N_9401,N_9866);
or U10349 (N_10349,N_8090,N_8447);
nor U10350 (N_10350,N_9354,N_9856);
and U10351 (N_10351,N_9358,N_8320);
or U10352 (N_10352,N_8891,N_9240);
and U10353 (N_10353,N_9209,N_9110);
nor U10354 (N_10354,N_9233,N_9152);
nand U10355 (N_10355,N_9932,N_9050);
nor U10356 (N_10356,N_9436,N_9466);
and U10357 (N_10357,N_8302,N_9181);
or U10358 (N_10358,N_8642,N_9899);
nand U10359 (N_10359,N_8928,N_9022);
xnor U10360 (N_10360,N_8338,N_8717);
or U10361 (N_10361,N_9702,N_9404);
nor U10362 (N_10362,N_9133,N_9507);
nand U10363 (N_10363,N_9648,N_8735);
nand U10364 (N_10364,N_9082,N_8387);
xnor U10365 (N_10365,N_8180,N_9720);
or U10366 (N_10366,N_8198,N_8766);
nand U10367 (N_10367,N_8421,N_9106);
nor U10368 (N_10368,N_9553,N_9415);
nand U10369 (N_10369,N_8807,N_9375);
or U10370 (N_10370,N_8424,N_8195);
or U10371 (N_10371,N_9215,N_8154);
nor U10372 (N_10372,N_8005,N_8811);
and U10373 (N_10373,N_9051,N_8065);
and U10374 (N_10374,N_8635,N_9531);
nand U10375 (N_10375,N_9691,N_9504);
nor U10376 (N_10376,N_8247,N_9037);
nand U10377 (N_10377,N_8732,N_8436);
and U10378 (N_10378,N_9643,N_8117);
nand U10379 (N_10379,N_9366,N_9628);
nor U10380 (N_10380,N_9819,N_9717);
or U10381 (N_10381,N_8985,N_9858);
nand U10382 (N_10382,N_8442,N_8862);
and U10383 (N_10383,N_9386,N_9090);
and U10384 (N_10384,N_9759,N_9884);
and U10385 (N_10385,N_8850,N_8725);
nand U10386 (N_10386,N_9159,N_8651);
nand U10387 (N_10387,N_8135,N_8744);
xnor U10388 (N_10388,N_8197,N_8594);
nand U10389 (N_10389,N_8288,N_8633);
or U10390 (N_10390,N_8654,N_9121);
and U10391 (N_10391,N_8076,N_8584);
or U10392 (N_10392,N_9930,N_9805);
nand U10393 (N_10393,N_8360,N_9570);
nand U10394 (N_10394,N_9188,N_9852);
and U10395 (N_10395,N_8095,N_9634);
nand U10396 (N_10396,N_9787,N_9130);
xnor U10397 (N_10397,N_9216,N_8134);
and U10398 (N_10398,N_8187,N_8274);
xor U10399 (N_10399,N_8061,N_9031);
and U10400 (N_10400,N_9980,N_8520);
nor U10401 (N_10401,N_9100,N_9665);
xnor U10402 (N_10402,N_8156,N_8542);
nor U10403 (N_10403,N_9493,N_9502);
or U10404 (N_10404,N_8403,N_9283);
nor U10405 (N_10405,N_9123,N_9827);
nor U10406 (N_10406,N_8768,N_9516);
and U10407 (N_10407,N_9154,N_9461);
nor U10408 (N_10408,N_8169,N_8569);
or U10409 (N_10409,N_9975,N_9619);
and U10410 (N_10410,N_8291,N_8237);
xnor U10411 (N_10411,N_8057,N_9747);
and U10412 (N_10412,N_8174,N_8199);
and U10413 (N_10413,N_8202,N_8574);
or U10414 (N_10414,N_8780,N_8466);
nor U10415 (N_10415,N_9396,N_9146);
or U10416 (N_10416,N_8544,N_8042);
nor U10417 (N_10417,N_9862,N_9711);
nor U10418 (N_10418,N_8587,N_9926);
and U10419 (N_10419,N_8053,N_8227);
and U10420 (N_10420,N_9810,N_9400);
or U10421 (N_10421,N_8483,N_8962);
nand U10422 (N_10422,N_9876,N_8671);
nor U10423 (N_10423,N_8589,N_8545);
nor U10424 (N_10424,N_9530,N_9339);
nor U10425 (N_10425,N_8253,N_9983);
or U10426 (N_10426,N_9194,N_9616);
nor U10427 (N_10427,N_8509,N_8534);
or U10428 (N_10428,N_8106,N_8762);
nand U10429 (N_10429,N_8257,N_9776);
nand U10430 (N_10430,N_8906,N_9433);
nor U10431 (N_10431,N_8707,N_8408);
or U10432 (N_10432,N_8937,N_8521);
and U10433 (N_10433,N_9814,N_8693);
nor U10434 (N_10434,N_8111,N_9857);
or U10435 (N_10435,N_9316,N_9214);
or U10436 (N_10436,N_8315,N_9314);
and U10437 (N_10437,N_8637,N_9645);
or U10438 (N_10438,N_9677,N_8869);
and U10439 (N_10439,N_8753,N_9268);
or U10440 (N_10440,N_9442,N_8495);
nand U10441 (N_10441,N_9555,N_8308);
nand U10442 (N_10442,N_8965,N_8705);
and U10443 (N_10443,N_9252,N_9609);
or U10444 (N_10444,N_9093,N_8982);
nand U10445 (N_10445,N_8760,N_8645);
nand U10446 (N_10446,N_8210,N_9859);
nand U10447 (N_10447,N_9452,N_9506);
xnor U10448 (N_10448,N_9586,N_8622);
nor U10449 (N_10449,N_8956,N_8297);
or U10450 (N_10450,N_8269,N_8069);
nand U10451 (N_10451,N_9742,N_9913);
or U10452 (N_10452,N_8131,N_8681);
or U10453 (N_10453,N_8868,N_9627);
nor U10454 (N_10454,N_9041,N_8643);
and U10455 (N_10455,N_9836,N_8190);
and U10456 (N_10456,N_9276,N_9903);
nand U10457 (N_10457,N_8954,N_8797);
nand U10458 (N_10458,N_8591,N_8712);
and U10459 (N_10459,N_8292,N_8309);
and U10460 (N_10460,N_8303,N_8212);
nand U10461 (N_10461,N_9765,N_9978);
and U10462 (N_10462,N_8140,N_9825);
xor U10463 (N_10463,N_8341,N_9013);
nand U10464 (N_10464,N_9290,N_8370);
nand U10465 (N_10465,N_8022,N_8570);
and U10466 (N_10466,N_8373,N_8698);
nand U10467 (N_10467,N_8019,N_8778);
and U10468 (N_10468,N_9084,N_8423);
and U10469 (N_10469,N_8571,N_9096);
and U10470 (N_10470,N_8038,N_9725);
nor U10471 (N_10471,N_9319,N_8270);
nor U10472 (N_10472,N_9584,N_8851);
nand U10473 (N_10473,N_8665,N_9070);
xor U10474 (N_10474,N_9422,N_9485);
nand U10475 (N_10475,N_8913,N_8812);
or U10476 (N_10476,N_9098,N_9591);
and U10477 (N_10477,N_9548,N_8230);
and U10478 (N_10478,N_8628,N_9956);
nor U10479 (N_10479,N_8547,N_8464);
or U10480 (N_10480,N_9350,N_8777);
or U10481 (N_10481,N_8852,N_9680);
nor U10482 (N_10482,N_9289,N_8296);
nor U10483 (N_10483,N_8988,N_9898);
nor U10484 (N_10484,N_9467,N_8903);
and U10485 (N_10485,N_9213,N_8990);
or U10486 (N_10486,N_8677,N_8099);
xor U10487 (N_10487,N_9647,N_9045);
xnor U10488 (N_10488,N_8966,N_8388);
nor U10489 (N_10489,N_8733,N_9596);
and U10490 (N_10490,N_9736,N_8946);
and U10491 (N_10491,N_8764,N_9468);
nor U10492 (N_10492,N_9997,N_9021);
nand U10493 (N_10493,N_8500,N_8639);
nand U10494 (N_10494,N_8206,N_8339);
or U10495 (N_10495,N_8039,N_8560);
nor U10496 (N_10496,N_8392,N_8012);
or U10497 (N_10497,N_9536,N_9164);
and U10498 (N_10498,N_9177,N_8661);
nand U10499 (N_10499,N_9060,N_8215);
or U10500 (N_10500,N_8406,N_9924);
nand U10501 (N_10501,N_9771,N_8078);
or U10502 (N_10502,N_8056,N_8248);
nand U10503 (N_10503,N_8670,N_9821);
or U10504 (N_10504,N_9267,N_9241);
nor U10505 (N_10505,N_9807,N_8751);
xnor U10506 (N_10506,N_8849,N_9626);
nand U10507 (N_10507,N_8233,N_8636);
nor U10508 (N_10508,N_8960,N_8615);
nand U10509 (N_10509,N_9959,N_9499);
and U10510 (N_10510,N_9301,N_9694);
and U10511 (N_10511,N_8382,N_9277);
or U10512 (N_10512,N_9309,N_9189);
xor U10513 (N_10513,N_8034,N_8487);
nor U10514 (N_10514,N_9230,N_9613);
nor U10515 (N_10515,N_8252,N_9620);
xor U10516 (N_10516,N_8217,N_9949);
nand U10517 (N_10517,N_8714,N_9287);
nand U10518 (N_10518,N_8832,N_9835);
nand U10519 (N_10519,N_9803,N_9914);
or U10520 (N_10520,N_9888,N_8264);
xnor U10521 (N_10521,N_9373,N_8804);
xor U10522 (N_10522,N_8031,N_9732);
nor U10523 (N_10523,N_9338,N_8527);
or U10524 (N_10524,N_8085,N_8481);
nor U10525 (N_10525,N_8634,N_9864);
nand U10526 (N_10526,N_8537,N_9072);
nor U10527 (N_10527,N_9243,N_8834);
and U10528 (N_10528,N_8066,N_8943);
nor U10529 (N_10529,N_8814,N_8839);
nand U10530 (N_10530,N_9546,N_9097);
or U10531 (N_10531,N_8335,N_8971);
or U10532 (N_10532,N_8718,N_9080);
and U10533 (N_10533,N_8063,N_9362);
or U10534 (N_10534,N_8285,N_8837);
or U10535 (N_10535,N_9848,N_8414);
or U10536 (N_10536,N_9421,N_9236);
nand U10537 (N_10537,N_8009,N_8968);
xor U10538 (N_10538,N_9576,N_8612);
or U10539 (N_10539,N_9183,N_9298);
nand U10540 (N_10540,N_9563,N_9197);
and U10541 (N_10541,N_8556,N_8874);
xor U10542 (N_10542,N_8021,N_9731);
or U10543 (N_10543,N_8719,N_9225);
or U10544 (N_10544,N_8116,N_8690);
and U10545 (N_10545,N_9470,N_9478);
or U10546 (N_10546,N_9055,N_9042);
and U10547 (N_10547,N_8886,N_9079);
or U10548 (N_10548,N_9789,N_9820);
nor U10549 (N_10549,N_9875,N_8327);
and U10550 (N_10550,N_8030,N_9326);
and U10551 (N_10551,N_8831,N_8893);
or U10552 (N_10552,N_8729,N_9117);
nor U10553 (N_10553,N_9263,N_8287);
nand U10554 (N_10554,N_9487,N_9733);
and U10555 (N_10555,N_8494,N_9437);
or U10556 (N_10556,N_9166,N_8538);
or U10557 (N_10557,N_8460,N_8948);
and U10558 (N_10558,N_9969,N_9431);
nor U10559 (N_10559,N_8445,N_9573);
and U10560 (N_10560,N_8081,N_9143);
nor U10561 (N_10561,N_8452,N_9746);
xor U10562 (N_10562,N_9245,N_8001);
nand U10563 (N_10563,N_9542,N_8911);
or U10564 (N_10564,N_9639,N_8224);
or U10565 (N_10565,N_8840,N_9801);
and U10566 (N_10566,N_8226,N_9740);
nor U10567 (N_10567,N_9981,N_8526);
nor U10568 (N_10568,N_9101,N_9673);
or U10569 (N_10569,N_8068,N_8535);
nand U10570 (N_10570,N_8207,N_8157);
or U10571 (N_10571,N_9033,N_8564);
and U10572 (N_10572,N_8278,N_9772);
nand U10573 (N_10573,N_8624,N_9935);
nor U10574 (N_10574,N_9501,N_8603);
or U10575 (N_10575,N_8861,N_9831);
and U10576 (N_10576,N_9528,N_8121);
nand U10577 (N_10577,N_9322,N_9129);
nor U10578 (N_10578,N_8110,N_9393);
nor U10579 (N_10579,N_9363,N_9242);
and U10580 (N_10580,N_9682,N_9806);
nor U10581 (N_10581,N_9167,N_8798);
nand U10582 (N_10582,N_9943,N_9911);
xnor U10583 (N_10583,N_9514,N_9750);
nand U10584 (N_10584,N_9992,N_9841);
nor U10585 (N_10585,N_9451,N_9126);
and U10586 (N_10586,N_8035,N_8344);
and U10587 (N_10587,N_9357,N_9025);
nor U10588 (N_10588,N_9703,N_8926);
and U10589 (N_10589,N_9766,N_9922);
nor U10590 (N_10590,N_9741,N_9075);
nor U10591 (N_10591,N_9169,N_9426);
or U10592 (N_10592,N_9369,N_8448);
nor U10593 (N_10593,N_8501,N_8333);
nor U10594 (N_10594,N_9974,N_8472);
nor U10595 (N_10595,N_8958,N_8075);
nor U10596 (N_10596,N_8743,N_9275);
nor U10597 (N_10597,N_9340,N_8900);
nor U10598 (N_10598,N_8345,N_8844);
nand U10599 (N_10599,N_8715,N_9947);
or U10600 (N_10600,N_8177,N_8016);
or U10601 (N_10601,N_9028,N_9678);
and U10602 (N_10602,N_9569,N_9083);
nand U10603 (N_10603,N_9659,N_9572);
nor U10604 (N_10604,N_8518,N_8167);
nor U10605 (N_10605,N_8590,N_8549);
xnor U10606 (N_10606,N_9738,N_8599);
nor U10607 (N_10607,N_9860,N_9140);
nand U10608 (N_10608,N_8399,N_8354);
nand U10609 (N_10609,N_9286,N_8757);
or U10610 (N_10610,N_8630,N_9342);
nor U10611 (N_10611,N_8386,N_9427);
xor U10612 (N_10612,N_9141,N_8734);
nand U10613 (N_10613,N_8939,N_8618);
or U10614 (N_10614,N_8833,N_8676);
nand U10615 (N_10615,N_8422,N_8873);
xor U10616 (N_10616,N_8064,N_8351);
or U10617 (N_10617,N_9500,N_8262);
nor U10618 (N_10618,N_9367,N_8165);
or U10619 (N_10619,N_8120,N_9074);
and U10620 (N_10620,N_8910,N_9660);
nand U10621 (N_10621,N_8463,N_8539);
xnor U10622 (N_10622,N_8062,N_8391);
nor U10623 (N_10623,N_9655,N_9250);
nor U10624 (N_10624,N_8092,N_9994);
or U10625 (N_10625,N_9238,N_9477);
nand U10626 (N_10626,N_8763,N_8467);
or U10627 (N_10627,N_8823,N_9509);
or U10628 (N_10628,N_8682,N_8808);
nor U10629 (N_10629,N_9718,N_9575);
nand U10630 (N_10630,N_8945,N_9099);
nor U10631 (N_10631,N_9307,N_8468);
and U10632 (N_10632,N_8588,N_8685);
nand U10633 (N_10633,N_8770,N_8407);
and U10634 (N_10634,N_8011,N_8923);
nand U10635 (N_10635,N_9175,N_8304);
xor U10636 (N_10636,N_9799,N_8992);
nor U10637 (N_10637,N_9795,N_9885);
nor U10638 (N_10638,N_8616,N_8892);
xnor U10639 (N_10639,N_9784,N_8776);
and U10640 (N_10640,N_8925,N_8908);
xor U10641 (N_10641,N_9892,N_9429);
nand U10642 (N_10642,N_9184,N_8887);
nand U10643 (N_10643,N_9313,N_9566);
nor U10644 (N_10644,N_8086,N_8703);
xnor U10645 (N_10645,N_8810,N_9979);
nand U10646 (N_10646,N_8731,N_8947);
or U10647 (N_10647,N_8904,N_8566);
and U10648 (N_10648,N_9463,N_8349);
or U10649 (N_10649,N_9535,N_9638);
or U10650 (N_10650,N_9071,N_8942);
or U10651 (N_10651,N_8124,N_8929);
or U10652 (N_10652,N_8546,N_9204);
and U10653 (N_10653,N_8170,N_8171);
xor U10654 (N_10654,N_9692,N_8008);
nand U10655 (N_10655,N_9918,N_9637);
nand U10656 (N_10656,N_9395,N_9642);
and U10657 (N_10657,N_8978,N_9669);
nand U10658 (N_10658,N_9523,N_8848);
nand U10659 (N_10659,N_8846,N_8347);
nor U10660 (N_10660,N_9600,N_8652);
nand U10661 (N_10661,N_8245,N_8451);
xnor U10662 (N_10662,N_9735,N_9158);
and U10663 (N_10663,N_9480,N_8196);
xor U10664 (N_10664,N_8957,N_9559);
nand U10665 (N_10665,N_8640,N_8112);
and U10666 (N_10666,N_8775,N_8818);
and U10667 (N_10667,N_8601,N_9890);
nand U10668 (N_10668,N_9762,N_9580);
or U10669 (N_10669,N_9770,N_9957);
and U10670 (N_10670,N_9005,N_8741);
nor U10671 (N_10671,N_8882,N_9163);
nor U10672 (N_10672,N_9781,N_8173);
or U10673 (N_10673,N_9102,N_8897);
or U10674 (N_10674,N_9036,N_9987);
nor U10675 (N_10675,N_9195,N_8352);
and U10676 (N_10676,N_8381,N_9335);
and U10677 (N_10677,N_8932,N_8105);
or U10678 (N_10678,N_8994,N_8748);
or U10679 (N_10679,N_9962,N_9843);
nand U10680 (N_10680,N_9293,N_9425);
nand U10681 (N_10681,N_8044,N_9026);
nand U10682 (N_10682,N_8953,N_8655);
nand U10683 (N_10683,N_9253,N_8720);
or U10684 (N_10684,N_8096,N_9039);
and U10685 (N_10685,N_9568,N_8243);
nand U10686 (N_10686,N_8533,N_8610);
and U10687 (N_10687,N_8786,N_8515);
and U10688 (N_10688,N_8397,N_9224);
or U10689 (N_10689,N_8621,N_8201);
and U10690 (N_10690,N_9952,N_8964);
nand U10691 (N_10691,N_9223,N_9331);
and U10692 (N_10692,N_8417,N_8512);
nand U10693 (N_10693,N_9526,N_9328);
or U10694 (N_10694,N_9828,N_8977);
or U10695 (N_10695,N_9343,N_9356);
nor U10696 (N_10696,N_8277,N_9695);
nor U10697 (N_10697,N_9671,N_9764);
nor U10698 (N_10698,N_9794,N_8241);
and U10699 (N_10699,N_9187,N_9558);
or U10700 (N_10700,N_8577,N_8856);
nand U10701 (N_10701,N_8866,N_9190);
nand U10702 (N_10702,N_9783,N_9708);
nor U10703 (N_10703,N_9381,N_9053);
nor U10704 (N_10704,N_9889,N_8146);
nand U10705 (N_10705,N_9085,N_8077);
nand U10706 (N_10706,N_9303,N_9728);
and U10707 (N_10707,N_9474,N_9353);
nand U10708 (N_10708,N_9873,N_8014);
nand U10709 (N_10709,N_9457,N_9826);
and U10710 (N_10710,N_9221,N_9047);
and U10711 (N_10711,N_9946,N_9774);
or U10712 (N_10712,N_8629,N_8328);
and U10713 (N_10713,N_9254,N_9227);
nand U10714 (N_10714,N_9788,N_9839);
xnor U10715 (N_10715,N_9610,N_8050);
nand U10716 (N_10716,N_8684,N_8082);
nor U10717 (N_10717,N_8434,N_9607);
xor U10718 (N_10718,N_8638,N_9666);
and U10719 (N_10719,N_8706,N_8425);
or U10720 (N_10720,N_9046,N_8203);
or U10721 (N_10721,N_8244,N_9745);
and U10722 (N_10722,N_8979,N_9503);
nand U10723 (N_10723,N_9554,N_9418);
nor U10724 (N_10724,N_8575,N_9348);
nand U10725 (N_10725,N_8796,N_9496);
or U10726 (N_10726,N_8894,N_9274);
and U10727 (N_10727,N_8523,N_9939);
xor U10728 (N_10728,N_8975,N_8789);
and U10729 (N_10729,N_9904,N_8125);
nand U10730 (N_10730,N_8740,N_8179);
nand U10731 (N_10731,N_8825,N_8409);
and U10732 (N_10732,N_8410,N_9905);
nand U10733 (N_10733,N_8058,N_8936);
xor U10734 (N_10734,N_9412,N_9137);
nand U10735 (N_10735,N_8013,N_9871);
and U10736 (N_10736,N_9990,N_9583);
or U10737 (N_10737,N_9405,N_9234);
nand U10738 (N_10738,N_8465,N_8669);
nand U10739 (N_10739,N_9109,N_9920);
or U10740 (N_10740,N_9325,N_9808);
or U10741 (N_10741,N_9715,N_9714);
and U10742 (N_10742,N_8870,N_9760);
xnor U10743 (N_10743,N_8275,N_8816);
and U10744 (N_10744,N_9851,N_9336);
or U10745 (N_10745,N_8597,N_9744);
nor U10746 (N_10746,N_8689,N_9364);
nand U10747 (N_10747,N_9482,N_9512);
nor U10748 (N_10748,N_8168,N_9973);
nand U10749 (N_10749,N_9995,N_9823);
nand U10750 (N_10750,N_8675,N_8007);
nand U10751 (N_10751,N_8997,N_8674);
nand U10752 (N_10752,N_9625,N_8428);
nand U10753 (N_10753,N_8683,N_8362);
nand U10754 (N_10754,N_9125,N_8398);
nor U10755 (N_10755,N_9513,N_9419);
and U10756 (N_10756,N_9796,N_8632);
nand U10757 (N_10757,N_8600,N_9459);
nand U10758 (N_10758,N_9698,N_9360);
xnor U10759 (N_10759,N_9498,N_8272);
and U10760 (N_10760,N_8504,N_9611);
xnor U10761 (N_10761,N_8898,N_9689);
and U10762 (N_10762,N_9597,N_8754);
or U10763 (N_10763,N_8641,N_9608);
and U10764 (N_10764,N_8143,N_9700);
nor U10765 (N_10765,N_9934,N_8486);
or U10766 (N_10766,N_9786,N_9812);
xnor U10767 (N_10767,N_9262,N_8477);
nand U10768 (N_10768,N_8089,N_8697);
nand U10769 (N_10769,N_8513,N_9281);
xor U10770 (N_10770,N_8258,N_9544);
and U10771 (N_10771,N_8369,N_9043);
or U10772 (N_10772,N_8359,N_8657);
or U10773 (N_10773,N_9077,N_9018);
xnor U10774 (N_10774,N_9874,N_9327);
nor U10775 (N_10775,N_9220,N_8094);
xnor U10776 (N_10776,N_8221,N_9847);
nor U10777 (N_10777,N_9078,N_9967);
and U10778 (N_10778,N_8611,N_9879);
or U10779 (N_10779,N_8301,N_9855);
or U10780 (N_10780,N_8182,N_8454);
or U10781 (N_10781,N_9264,N_9368);
nand U10782 (N_10782,N_9460,N_9938);
nand U10783 (N_10783,N_8420,N_8478);
or U10784 (N_10784,N_8759,N_8331);
nor U10785 (N_10785,N_9122,N_8307);
or U10786 (N_10786,N_8993,N_8802);
nand U10787 (N_10787,N_8129,N_9211);
nand U10788 (N_10788,N_9107,N_9237);
nor U10789 (N_10789,N_8356,N_8045);
nor U10790 (N_10790,N_9752,N_9009);
nand U10791 (N_10791,N_8578,N_9630);
and U10792 (N_10792,N_8152,N_9953);
xnor U10793 (N_10793,N_9897,N_8858);
and U10794 (N_10794,N_8025,N_8702);
nand U10795 (N_10795,N_8663,N_9589);
or U10796 (N_10796,N_9972,N_9489);
nand U10797 (N_10797,N_9909,N_8048);
nand U10798 (N_10798,N_8093,N_9719);
and U10799 (N_10799,N_9447,N_9525);
nand U10800 (N_10800,N_8473,N_9891);
or U10801 (N_10801,N_9420,N_9989);
nor U10802 (N_10802,N_8648,N_9945);
and U10803 (N_10803,N_8983,N_8922);
nand U10804 (N_10804,N_9192,N_9763);
and U10805 (N_10805,N_9035,N_9049);
or U10806 (N_10806,N_8040,N_9329);
or U10807 (N_10807,N_8644,N_9699);
and U10808 (N_10808,N_8553,N_9910);
nand U10809 (N_10809,N_8260,N_8522);
nor U10810 (N_10810,N_8559,N_9676);
nor U10811 (N_10811,N_9928,N_9323);
or U10812 (N_10812,N_9779,N_8367);
or U10813 (N_10813,N_8996,N_9704);
nor U10814 (N_10814,N_9894,N_8613);
and U10815 (N_10815,N_9308,N_8952);
and U10816 (N_10816,N_9272,N_9950);
or U10817 (N_10817,N_8625,N_8225);
nand U10818 (N_10818,N_8989,N_9222);
and U10819 (N_10819,N_8132,N_9838);
and U10820 (N_10820,N_9208,N_9384);
nor U10821 (N_10821,N_9210,N_8026);
nor U10822 (N_10822,N_8568,N_8881);
xor U10823 (N_10823,N_8181,N_9511);
and U10824 (N_10824,N_8457,N_8312);
nor U10825 (N_10825,N_8490,N_9661);
xnor U10826 (N_10826,N_8128,N_9441);
nand U10827 (N_10827,N_8664,N_9176);
or U10828 (N_10828,N_9359,N_8709);
nand U10829 (N_10829,N_9527,N_9964);
nor U10830 (N_10830,N_9811,N_8905);
nor U10831 (N_10831,N_8917,N_8581);
nor U10832 (N_10832,N_9670,N_9201);
nand U10833 (N_10833,N_9257,N_8340);
nand U10834 (N_10834,N_8503,N_8649);
nand U10835 (N_10835,N_9469,N_9269);
nand U10836 (N_10836,N_9186,N_9483);
and U10837 (N_10837,N_8266,N_9377);
xor U10838 (N_10838,N_9058,N_9961);
xnor U10839 (N_10839,N_8060,N_9413);
nor U10840 (N_10840,N_8336,N_8186);
nor U10841 (N_10841,N_9739,N_8479);
and U10842 (N_10842,N_9524,N_9664);
and U10843 (N_10843,N_8450,N_9712);
nand U10844 (N_10844,N_9534,N_9830);
nor U10845 (N_10845,N_9088,N_8999);
and U10846 (N_10846,N_9010,N_9594);
nand U10847 (N_10847,N_9662,N_8261);
xnor U10848 (N_10848,N_9842,N_8433);
xnor U10849 (N_10849,N_9756,N_9614);
xnor U10850 (N_10850,N_8239,N_8059);
xnor U10851 (N_10851,N_8608,N_9321);
and U10852 (N_10852,N_9040,N_8737);
and U10853 (N_10853,N_9641,N_9550);
xnor U10854 (N_10854,N_9128,N_8286);
and U10855 (N_10855,N_9337,N_9024);
nand U10856 (N_10856,N_8949,N_9545);
or U10857 (N_10857,N_9199,N_9417);
and U10858 (N_10858,N_8507,N_9561);
or U10859 (N_10859,N_9601,N_8435);
and U10860 (N_10860,N_9473,N_8036);
or U10861 (N_10861,N_9844,N_9057);
or U10862 (N_10862,N_9091,N_8209);
or U10863 (N_10863,N_8830,N_8824);
xnor U10864 (N_10864,N_9491,N_9845);
or U10865 (N_10865,N_8133,N_8653);
xor U10866 (N_10866,N_8346,N_9693);
xor U10867 (N_10867,N_9681,N_8027);
and U10868 (N_10868,N_8828,N_8667);
xnor U10869 (N_10869,N_8299,N_9304);
or U10870 (N_10870,N_8711,N_9727);
or U10871 (N_10871,N_9388,N_9300);
and U10872 (N_10872,N_8563,N_8598);
or U10873 (N_10873,N_9173,N_9235);
and U10874 (N_10874,N_8730,N_9105);
and U10875 (N_10875,N_9011,N_9604);
or U10876 (N_10876,N_8276,N_8322);
xnor U10877 (N_10877,N_9592,N_8506);
nand U10878 (N_10878,N_9135,N_9115);
nand U10879 (N_10879,N_9606,N_9977);
nor U10880 (N_10880,N_9428,N_9893);
nand U10881 (N_10881,N_9202,N_9654);
xor U10882 (N_10882,N_9815,N_9998);
nor U10883 (N_10883,N_9392,N_9438);
nor U10884 (N_10884,N_8271,N_9867);
and U10885 (N_10885,N_8879,N_9108);
xor U10886 (N_10886,N_9352,N_8826);
and U10887 (N_10887,N_8400,N_8366);
or U10888 (N_10888,N_8919,N_8857);
and U10889 (N_10889,N_8330,N_9697);
or U10890 (N_10890,N_9150,N_8561);
and U10891 (N_10891,N_9510,N_9349);
or U10892 (N_10892,N_9556,N_8836);
nand U10893 (N_10893,N_9258,N_9206);
nand U10894 (N_10894,N_9579,N_9095);
and U10895 (N_10895,N_9407,N_8159);
and U10896 (N_10896,N_9769,N_9315);
nand U10897 (N_10897,N_8688,N_9446);
or U10898 (N_10898,N_9777,N_8916);
and U10899 (N_10899,N_9631,N_8516);
and U10900 (N_10900,N_9602,N_8361);
nor U10901 (N_10901,N_9038,N_9261);
nor U10902 (N_10902,N_8444,N_9059);
and U10903 (N_10903,N_9748,N_9598);
and U10904 (N_10904,N_9632,N_8972);
or U10905 (N_10905,N_8791,N_9865);
nor U10906 (N_10906,N_9656,N_9896);
or U10907 (N_10907,N_9870,N_8205);
xor U10908 (N_10908,N_9942,N_9549);
nand U10909 (N_10909,N_9475,N_8890);
nor U10910 (N_10910,N_8627,N_9646);
and U10911 (N_10911,N_8300,N_9529);
nor U10912 (N_10912,N_8736,N_8211);
or U10913 (N_10913,N_8332,N_8054);
or U10914 (N_10914,N_8337,N_8704);
or U10915 (N_10915,N_8695,N_9012);
nor U10916 (N_10916,N_9023,N_9064);
xnor U10917 (N_10917,N_8412,N_8821);
and U10918 (N_10918,N_9065,N_8781);
nor U10919 (N_10919,N_8901,N_8443);
nor U10920 (N_10920,N_8884,N_8350);
nand U10921 (N_10921,N_9658,N_9624);
or U10922 (N_10922,N_8880,N_8268);
nand U10923 (N_10923,N_9615,N_8456);
or U10924 (N_10924,N_8548,N_9722);
and U10925 (N_10925,N_8799,N_9076);
and U10926 (N_10926,N_8118,N_9246);
or U10927 (N_10927,N_9456,N_9492);
nand U10928 (N_10928,N_8375,N_9832);
xnor U10929 (N_10929,N_9791,N_8427);
nor U10930 (N_10930,N_8136,N_9027);
or U10931 (N_10931,N_9443,N_9588);
or U10932 (N_10932,N_8379,N_8010);
and U10933 (N_10933,N_8573,N_8413);
nand U10934 (N_10934,N_8384,N_9270);
or U10935 (N_10935,N_8931,N_8623);
or U10936 (N_10936,N_8716,N_8955);
xor U10937 (N_10937,N_9966,N_9156);
or U10938 (N_10938,N_9793,N_9001);
or U10939 (N_10939,N_9180,N_9411);
and U10940 (N_10940,N_8325,N_9802);
xor U10941 (N_10941,N_9318,N_8727);
or U10942 (N_10942,N_9785,N_8819);
xnor U10943 (N_10943,N_9278,N_8363);
nand U10944 (N_10944,N_8402,N_9019);
nor U10945 (N_10945,N_8724,N_9951);
and U10946 (N_10946,N_8519,N_8700);
and U10947 (N_10947,N_9104,N_9685);
nand U10948 (N_10948,N_8323,N_9185);
nor U10949 (N_10949,N_9650,N_9462);
and U10950 (N_10950,N_8650,N_9578);
and U10951 (N_10951,N_9089,N_9282);
nand U10952 (N_10952,N_8550,N_8795);
nor U10953 (N_10953,N_8394,N_9014);
nand U10954 (N_10954,N_9382,N_9455);
nor U10955 (N_10955,N_8696,N_8229);
nand U10956 (N_10956,N_8246,N_9191);
nor U10957 (N_10957,N_9587,N_9251);
xor U10958 (N_10958,N_9986,N_8841);
xor U10959 (N_10959,N_9538,N_8536);
and U10960 (N_10960,N_8153,N_8877);
nor U10961 (N_10961,N_8280,N_8528);
nor U10962 (N_10962,N_9054,N_9713);
and U10963 (N_10963,N_8921,N_9008);
xnor U10964 (N_10964,N_8484,N_9205);
nor U10965 (N_10965,N_9532,N_9773);
and U10966 (N_10966,N_8742,N_8256);
and U10967 (N_10967,N_9249,N_8596);
and U10968 (N_10968,N_8145,N_9955);
nor U10969 (N_10969,N_8505,N_8242);
nor U10970 (N_10970,N_8617,N_9016);
nand U10971 (N_10971,N_8104,N_9003);
nor U10972 (N_10972,N_8232,N_8313);
xnor U10973 (N_10973,N_9408,N_8758);
nand U10974 (N_10974,N_8213,N_8765);
nor U10975 (N_10975,N_9458,N_9218);
or U10976 (N_10976,N_9103,N_8508);
or U10977 (N_10977,N_9954,N_9397);
nor U10978 (N_10978,N_9145,N_9883);
or U10979 (N_10979,N_8172,N_8378);
nor U10980 (N_10980,N_8701,N_9633);
xnor U10981 (N_10981,N_9684,N_8429);
nor U10982 (N_10982,N_9248,N_8311);
nand U10983 (N_10983,N_9266,N_8974);
nor U10984 (N_10984,N_8785,N_8991);
nor U10985 (N_10985,N_8319,N_8321);
nand U10986 (N_10986,N_9044,N_9886);
nand U10987 (N_10987,N_9056,N_9148);
and U10988 (N_10988,N_9622,N_8959);
xor U10989 (N_10989,N_9929,N_8497);
or U10990 (N_10990,N_8183,N_8234);
nand U10991 (N_10991,N_9207,N_8631);
nor U10992 (N_10992,N_8787,N_9450);
nand U10993 (N_10993,N_8101,N_9907);
or U10994 (N_10994,N_9651,N_8453);
nor U10995 (N_10995,N_9464,N_8072);
xnor U10996 (N_10996,N_8458,N_8469);
nor U10997 (N_10997,N_8084,N_8119);
nand U10998 (N_10998,N_9917,N_8595);
and U10999 (N_10999,N_8185,N_8859);
and U11000 (N_11000,N_8586,N_9244);
xor U11001 (N_11001,N_8578,N_9608);
nor U11002 (N_11002,N_9850,N_8818);
nand U11003 (N_11003,N_8413,N_9648);
or U11004 (N_11004,N_8876,N_8790);
nor U11005 (N_11005,N_8292,N_8694);
and U11006 (N_11006,N_8545,N_8777);
nand U11007 (N_11007,N_8428,N_9048);
nand U11008 (N_11008,N_8280,N_8618);
or U11009 (N_11009,N_9562,N_9462);
and U11010 (N_11010,N_9545,N_8069);
xnor U11011 (N_11011,N_8383,N_9441);
xor U11012 (N_11012,N_9952,N_8065);
and U11013 (N_11013,N_8475,N_9450);
nand U11014 (N_11014,N_9990,N_8970);
nand U11015 (N_11015,N_8091,N_8453);
xnor U11016 (N_11016,N_8460,N_9194);
or U11017 (N_11017,N_8910,N_8611);
or U11018 (N_11018,N_8360,N_8581);
nand U11019 (N_11019,N_9857,N_8437);
and U11020 (N_11020,N_9901,N_9389);
nor U11021 (N_11021,N_8415,N_8617);
nand U11022 (N_11022,N_8613,N_8703);
or U11023 (N_11023,N_9267,N_9418);
nand U11024 (N_11024,N_8011,N_9235);
nor U11025 (N_11025,N_8522,N_9270);
nand U11026 (N_11026,N_9407,N_9257);
nor U11027 (N_11027,N_8265,N_8107);
or U11028 (N_11028,N_8488,N_8471);
nor U11029 (N_11029,N_9946,N_8180);
or U11030 (N_11030,N_8216,N_9001);
nor U11031 (N_11031,N_9350,N_8705);
nor U11032 (N_11032,N_8801,N_8053);
or U11033 (N_11033,N_9505,N_9022);
and U11034 (N_11034,N_8552,N_8518);
nand U11035 (N_11035,N_9973,N_9509);
nor U11036 (N_11036,N_9674,N_9112);
and U11037 (N_11037,N_9095,N_8785);
or U11038 (N_11038,N_8599,N_9267);
nor U11039 (N_11039,N_8320,N_8315);
or U11040 (N_11040,N_9731,N_8417);
and U11041 (N_11041,N_8749,N_9324);
nor U11042 (N_11042,N_8644,N_8355);
nor U11043 (N_11043,N_9121,N_9274);
or U11044 (N_11044,N_9419,N_9009);
or U11045 (N_11045,N_8047,N_8268);
nand U11046 (N_11046,N_9504,N_9215);
and U11047 (N_11047,N_8100,N_9988);
or U11048 (N_11048,N_8193,N_8034);
or U11049 (N_11049,N_9983,N_9772);
nor U11050 (N_11050,N_9833,N_9337);
nor U11051 (N_11051,N_9691,N_9795);
nand U11052 (N_11052,N_8091,N_9852);
nor U11053 (N_11053,N_9855,N_8408);
and U11054 (N_11054,N_9391,N_8008);
and U11055 (N_11055,N_8522,N_8546);
nor U11056 (N_11056,N_9046,N_9712);
nor U11057 (N_11057,N_8605,N_9435);
nor U11058 (N_11058,N_9117,N_9673);
nand U11059 (N_11059,N_8083,N_8327);
and U11060 (N_11060,N_9007,N_8659);
or U11061 (N_11061,N_9276,N_9333);
nor U11062 (N_11062,N_9473,N_8797);
nand U11063 (N_11063,N_9431,N_8345);
or U11064 (N_11064,N_8600,N_9019);
nand U11065 (N_11065,N_9987,N_9031);
and U11066 (N_11066,N_8302,N_8835);
or U11067 (N_11067,N_9295,N_8043);
and U11068 (N_11068,N_9993,N_9793);
or U11069 (N_11069,N_9891,N_9073);
nand U11070 (N_11070,N_8932,N_9683);
or U11071 (N_11071,N_9642,N_8733);
nor U11072 (N_11072,N_9602,N_9813);
nand U11073 (N_11073,N_8122,N_9954);
nand U11074 (N_11074,N_9703,N_8545);
xnor U11075 (N_11075,N_9457,N_9983);
and U11076 (N_11076,N_8683,N_8796);
nor U11077 (N_11077,N_8693,N_9647);
nand U11078 (N_11078,N_8516,N_9840);
nand U11079 (N_11079,N_8356,N_9264);
or U11080 (N_11080,N_8709,N_8310);
nand U11081 (N_11081,N_9701,N_8446);
nand U11082 (N_11082,N_9556,N_9955);
nand U11083 (N_11083,N_9324,N_9514);
and U11084 (N_11084,N_9947,N_9803);
nor U11085 (N_11085,N_8742,N_9701);
and U11086 (N_11086,N_8532,N_8591);
or U11087 (N_11087,N_8078,N_9168);
or U11088 (N_11088,N_9227,N_9239);
and U11089 (N_11089,N_9102,N_8591);
or U11090 (N_11090,N_8502,N_9167);
xnor U11091 (N_11091,N_9891,N_8616);
and U11092 (N_11092,N_8908,N_9552);
nor U11093 (N_11093,N_8606,N_8282);
or U11094 (N_11094,N_8936,N_9835);
xnor U11095 (N_11095,N_8366,N_8268);
and U11096 (N_11096,N_8527,N_8250);
nand U11097 (N_11097,N_8817,N_9667);
xor U11098 (N_11098,N_9602,N_8034);
nor U11099 (N_11099,N_9215,N_8460);
nand U11100 (N_11100,N_9954,N_9904);
nor U11101 (N_11101,N_9316,N_8429);
xor U11102 (N_11102,N_9729,N_8175);
nand U11103 (N_11103,N_8493,N_8788);
nor U11104 (N_11104,N_9927,N_8192);
nand U11105 (N_11105,N_8136,N_8669);
and U11106 (N_11106,N_8527,N_8594);
and U11107 (N_11107,N_8824,N_9071);
and U11108 (N_11108,N_8507,N_8695);
nand U11109 (N_11109,N_9905,N_9733);
nand U11110 (N_11110,N_8065,N_8074);
xnor U11111 (N_11111,N_8532,N_9191);
xor U11112 (N_11112,N_9026,N_8852);
and U11113 (N_11113,N_8679,N_8145);
nand U11114 (N_11114,N_9620,N_9096);
or U11115 (N_11115,N_9776,N_8350);
or U11116 (N_11116,N_9846,N_8383);
or U11117 (N_11117,N_8162,N_9169);
and U11118 (N_11118,N_8717,N_9414);
nand U11119 (N_11119,N_8642,N_9025);
and U11120 (N_11120,N_8329,N_9714);
nand U11121 (N_11121,N_8457,N_9369);
or U11122 (N_11122,N_8781,N_8609);
nor U11123 (N_11123,N_9537,N_9266);
nor U11124 (N_11124,N_8655,N_8842);
or U11125 (N_11125,N_8237,N_9261);
xnor U11126 (N_11126,N_9696,N_9154);
and U11127 (N_11127,N_9744,N_9283);
nand U11128 (N_11128,N_9703,N_8267);
or U11129 (N_11129,N_8896,N_8495);
and U11130 (N_11130,N_9249,N_9359);
nor U11131 (N_11131,N_8444,N_8830);
nor U11132 (N_11132,N_8100,N_8672);
and U11133 (N_11133,N_9500,N_9134);
nand U11134 (N_11134,N_9102,N_8507);
nand U11135 (N_11135,N_9143,N_9341);
or U11136 (N_11136,N_8805,N_8564);
nand U11137 (N_11137,N_8657,N_9228);
nand U11138 (N_11138,N_8625,N_9196);
or U11139 (N_11139,N_9922,N_9534);
nor U11140 (N_11140,N_8931,N_8605);
and U11141 (N_11141,N_9035,N_8935);
nand U11142 (N_11142,N_8892,N_8328);
and U11143 (N_11143,N_9274,N_9267);
and U11144 (N_11144,N_8320,N_8939);
nor U11145 (N_11145,N_8378,N_9196);
nor U11146 (N_11146,N_8343,N_8937);
nand U11147 (N_11147,N_9624,N_8854);
nand U11148 (N_11148,N_9099,N_8656);
and U11149 (N_11149,N_9322,N_8816);
and U11150 (N_11150,N_9998,N_9852);
or U11151 (N_11151,N_9544,N_8370);
nand U11152 (N_11152,N_9039,N_9447);
and U11153 (N_11153,N_9248,N_9659);
nor U11154 (N_11154,N_9574,N_8775);
or U11155 (N_11155,N_8306,N_9981);
or U11156 (N_11156,N_8079,N_9913);
and U11157 (N_11157,N_8324,N_8166);
xor U11158 (N_11158,N_8806,N_8647);
and U11159 (N_11159,N_9032,N_9515);
or U11160 (N_11160,N_9568,N_9466);
or U11161 (N_11161,N_9940,N_8573);
or U11162 (N_11162,N_9441,N_9221);
or U11163 (N_11163,N_9606,N_8964);
nand U11164 (N_11164,N_8981,N_8018);
or U11165 (N_11165,N_8758,N_9742);
nor U11166 (N_11166,N_8610,N_9136);
and U11167 (N_11167,N_9755,N_8562);
nor U11168 (N_11168,N_9855,N_8320);
or U11169 (N_11169,N_8433,N_8204);
and U11170 (N_11170,N_8142,N_9602);
nand U11171 (N_11171,N_8438,N_8929);
nor U11172 (N_11172,N_8155,N_9104);
xnor U11173 (N_11173,N_8492,N_8176);
and U11174 (N_11174,N_9500,N_8631);
nor U11175 (N_11175,N_8318,N_8063);
or U11176 (N_11176,N_9664,N_9765);
nor U11177 (N_11177,N_8874,N_9236);
and U11178 (N_11178,N_8878,N_8821);
nand U11179 (N_11179,N_8467,N_9657);
nor U11180 (N_11180,N_8434,N_9822);
or U11181 (N_11181,N_8092,N_9136);
nand U11182 (N_11182,N_9953,N_9212);
or U11183 (N_11183,N_9021,N_9395);
nand U11184 (N_11184,N_9643,N_9161);
nand U11185 (N_11185,N_9847,N_9119);
and U11186 (N_11186,N_8693,N_9174);
or U11187 (N_11187,N_8709,N_9547);
nand U11188 (N_11188,N_9567,N_9414);
nor U11189 (N_11189,N_9443,N_8214);
or U11190 (N_11190,N_9433,N_8305);
and U11191 (N_11191,N_8125,N_9374);
and U11192 (N_11192,N_9022,N_9738);
xnor U11193 (N_11193,N_8916,N_9868);
nor U11194 (N_11194,N_9012,N_8292);
nand U11195 (N_11195,N_8663,N_9393);
and U11196 (N_11196,N_8389,N_9835);
xnor U11197 (N_11197,N_8587,N_8859);
and U11198 (N_11198,N_8246,N_9464);
and U11199 (N_11199,N_8795,N_9142);
nor U11200 (N_11200,N_9337,N_9766);
or U11201 (N_11201,N_9332,N_8424);
nand U11202 (N_11202,N_9928,N_8049);
and U11203 (N_11203,N_9991,N_9642);
and U11204 (N_11204,N_8601,N_8564);
nand U11205 (N_11205,N_8352,N_9700);
nor U11206 (N_11206,N_8247,N_8673);
xnor U11207 (N_11207,N_9325,N_9451);
or U11208 (N_11208,N_8575,N_8584);
or U11209 (N_11209,N_8198,N_9790);
and U11210 (N_11210,N_9632,N_8204);
or U11211 (N_11211,N_8242,N_9131);
nand U11212 (N_11212,N_8964,N_8515);
and U11213 (N_11213,N_9844,N_9411);
and U11214 (N_11214,N_9744,N_8543);
nand U11215 (N_11215,N_9526,N_9451);
or U11216 (N_11216,N_8883,N_9195);
and U11217 (N_11217,N_9037,N_9936);
nor U11218 (N_11218,N_8637,N_9222);
nor U11219 (N_11219,N_8761,N_9775);
nor U11220 (N_11220,N_8103,N_8816);
and U11221 (N_11221,N_8036,N_9545);
nor U11222 (N_11222,N_8580,N_9108);
nor U11223 (N_11223,N_8070,N_9372);
and U11224 (N_11224,N_9441,N_8483);
nor U11225 (N_11225,N_8360,N_9923);
and U11226 (N_11226,N_8338,N_8455);
nor U11227 (N_11227,N_8520,N_9027);
nor U11228 (N_11228,N_9032,N_8319);
nor U11229 (N_11229,N_8093,N_9866);
nor U11230 (N_11230,N_8647,N_8102);
and U11231 (N_11231,N_8518,N_9105);
nor U11232 (N_11232,N_8500,N_9230);
nand U11233 (N_11233,N_8728,N_8503);
nor U11234 (N_11234,N_9276,N_9487);
nor U11235 (N_11235,N_9471,N_9563);
nor U11236 (N_11236,N_9514,N_8043);
or U11237 (N_11237,N_9759,N_8579);
and U11238 (N_11238,N_8133,N_9003);
xor U11239 (N_11239,N_9095,N_8598);
nor U11240 (N_11240,N_8791,N_8653);
or U11241 (N_11241,N_9655,N_9982);
nor U11242 (N_11242,N_8845,N_9319);
nand U11243 (N_11243,N_9065,N_9893);
and U11244 (N_11244,N_8758,N_8555);
or U11245 (N_11245,N_8016,N_8381);
or U11246 (N_11246,N_8471,N_9561);
nor U11247 (N_11247,N_9904,N_8137);
xor U11248 (N_11248,N_8573,N_9708);
nand U11249 (N_11249,N_8946,N_8227);
and U11250 (N_11250,N_9705,N_9294);
and U11251 (N_11251,N_8675,N_8785);
and U11252 (N_11252,N_9019,N_8653);
nand U11253 (N_11253,N_8918,N_8060);
nor U11254 (N_11254,N_9866,N_8936);
nor U11255 (N_11255,N_8106,N_9249);
and U11256 (N_11256,N_8089,N_9596);
nor U11257 (N_11257,N_9558,N_8530);
nor U11258 (N_11258,N_8866,N_9499);
xor U11259 (N_11259,N_9734,N_9731);
and U11260 (N_11260,N_8294,N_9846);
and U11261 (N_11261,N_8608,N_8512);
nand U11262 (N_11262,N_8399,N_8499);
nand U11263 (N_11263,N_8492,N_9124);
nand U11264 (N_11264,N_9438,N_8325);
nor U11265 (N_11265,N_9320,N_8583);
and U11266 (N_11266,N_8994,N_9243);
and U11267 (N_11267,N_9902,N_9159);
nor U11268 (N_11268,N_9053,N_9127);
nor U11269 (N_11269,N_9051,N_9556);
or U11270 (N_11270,N_9240,N_9775);
or U11271 (N_11271,N_8725,N_8693);
nand U11272 (N_11272,N_8180,N_9437);
nand U11273 (N_11273,N_8679,N_8578);
nand U11274 (N_11274,N_9463,N_9266);
and U11275 (N_11275,N_9294,N_8656);
nand U11276 (N_11276,N_8189,N_8281);
nor U11277 (N_11277,N_9206,N_9465);
or U11278 (N_11278,N_8563,N_8557);
xor U11279 (N_11279,N_9130,N_9911);
and U11280 (N_11280,N_8069,N_9247);
xor U11281 (N_11281,N_9311,N_9892);
or U11282 (N_11282,N_9221,N_9369);
nor U11283 (N_11283,N_8872,N_8307);
nor U11284 (N_11284,N_8217,N_8488);
nand U11285 (N_11285,N_9247,N_8918);
nor U11286 (N_11286,N_8393,N_9803);
nor U11287 (N_11287,N_8159,N_9439);
nor U11288 (N_11288,N_8095,N_8128);
or U11289 (N_11289,N_8831,N_8170);
nor U11290 (N_11290,N_8469,N_9885);
or U11291 (N_11291,N_9086,N_8896);
or U11292 (N_11292,N_8843,N_9586);
nand U11293 (N_11293,N_9064,N_8800);
nor U11294 (N_11294,N_9119,N_9229);
nand U11295 (N_11295,N_8722,N_9552);
or U11296 (N_11296,N_8517,N_9538);
nor U11297 (N_11297,N_8561,N_9616);
or U11298 (N_11298,N_9629,N_9505);
xnor U11299 (N_11299,N_9739,N_9887);
nor U11300 (N_11300,N_8666,N_8992);
or U11301 (N_11301,N_8218,N_8473);
nor U11302 (N_11302,N_8043,N_8404);
nand U11303 (N_11303,N_9884,N_8398);
and U11304 (N_11304,N_8965,N_9870);
or U11305 (N_11305,N_8821,N_9220);
nor U11306 (N_11306,N_9542,N_9264);
nor U11307 (N_11307,N_9210,N_9645);
xor U11308 (N_11308,N_8407,N_9208);
and U11309 (N_11309,N_8833,N_8485);
nor U11310 (N_11310,N_9183,N_9896);
or U11311 (N_11311,N_9472,N_8211);
or U11312 (N_11312,N_9474,N_8671);
or U11313 (N_11313,N_8112,N_9332);
and U11314 (N_11314,N_8908,N_9351);
nand U11315 (N_11315,N_8376,N_8340);
nand U11316 (N_11316,N_8806,N_8182);
nand U11317 (N_11317,N_8375,N_9199);
or U11318 (N_11318,N_8858,N_9520);
nor U11319 (N_11319,N_9488,N_8243);
nor U11320 (N_11320,N_9143,N_8360);
or U11321 (N_11321,N_8961,N_9562);
xnor U11322 (N_11322,N_8165,N_8370);
xor U11323 (N_11323,N_9944,N_8866);
nand U11324 (N_11324,N_9436,N_9173);
nand U11325 (N_11325,N_8675,N_8547);
nand U11326 (N_11326,N_9691,N_8800);
nand U11327 (N_11327,N_8180,N_9876);
or U11328 (N_11328,N_8263,N_8133);
nand U11329 (N_11329,N_8195,N_9465);
xnor U11330 (N_11330,N_9659,N_8459);
nand U11331 (N_11331,N_9417,N_9449);
nand U11332 (N_11332,N_9321,N_8044);
nor U11333 (N_11333,N_9238,N_8847);
and U11334 (N_11334,N_9658,N_8656);
or U11335 (N_11335,N_8930,N_9889);
nor U11336 (N_11336,N_9929,N_9864);
or U11337 (N_11337,N_9305,N_9552);
nor U11338 (N_11338,N_8601,N_8304);
nor U11339 (N_11339,N_8012,N_9632);
or U11340 (N_11340,N_8218,N_9032);
nor U11341 (N_11341,N_8604,N_8051);
nor U11342 (N_11342,N_9667,N_8124);
nor U11343 (N_11343,N_8938,N_8487);
xnor U11344 (N_11344,N_8100,N_8157);
nand U11345 (N_11345,N_8733,N_9623);
or U11346 (N_11346,N_8807,N_9815);
and U11347 (N_11347,N_9157,N_8309);
nor U11348 (N_11348,N_9997,N_9007);
nand U11349 (N_11349,N_9224,N_8261);
nand U11350 (N_11350,N_8608,N_9120);
or U11351 (N_11351,N_9888,N_8623);
and U11352 (N_11352,N_9614,N_9498);
or U11353 (N_11353,N_9259,N_9002);
and U11354 (N_11354,N_9256,N_8185);
and U11355 (N_11355,N_8988,N_9117);
nor U11356 (N_11356,N_9799,N_9329);
xor U11357 (N_11357,N_9078,N_8929);
nand U11358 (N_11358,N_9063,N_8775);
and U11359 (N_11359,N_8111,N_8586);
xor U11360 (N_11360,N_9705,N_8887);
or U11361 (N_11361,N_8233,N_8634);
xor U11362 (N_11362,N_8886,N_8219);
xnor U11363 (N_11363,N_8780,N_8158);
or U11364 (N_11364,N_9725,N_8184);
and U11365 (N_11365,N_9579,N_8407);
nand U11366 (N_11366,N_8967,N_9489);
xor U11367 (N_11367,N_8486,N_9520);
and U11368 (N_11368,N_9691,N_8176);
or U11369 (N_11369,N_8773,N_8513);
or U11370 (N_11370,N_9325,N_8474);
nor U11371 (N_11371,N_8501,N_8619);
nand U11372 (N_11372,N_8766,N_9703);
nand U11373 (N_11373,N_9934,N_9186);
or U11374 (N_11374,N_8189,N_8880);
nand U11375 (N_11375,N_9223,N_9662);
nor U11376 (N_11376,N_8115,N_9408);
xnor U11377 (N_11377,N_8609,N_8474);
and U11378 (N_11378,N_8588,N_9111);
nor U11379 (N_11379,N_9686,N_8428);
xnor U11380 (N_11380,N_8469,N_9719);
or U11381 (N_11381,N_8974,N_8729);
or U11382 (N_11382,N_8605,N_8141);
or U11383 (N_11383,N_9610,N_9472);
or U11384 (N_11384,N_9478,N_9790);
xnor U11385 (N_11385,N_8504,N_8402);
or U11386 (N_11386,N_8522,N_9422);
nand U11387 (N_11387,N_9120,N_9341);
and U11388 (N_11388,N_9365,N_9158);
and U11389 (N_11389,N_8656,N_8296);
xor U11390 (N_11390,N_8566,N_8068);
nand U11391 (N_11391,N_8785,N_9862);
nor U11392 (N_11392,N_8105,N_9138);
and U11393 (N_11393,N_8277,N_9232);
and U11394 (N_11394,N_9554,N_8004);
nand U11395 (N_11395,N_9698,N_9701);
nand U11396 (N_11396,N_9847,N_9702);
nand U11397 (N_11397,N_9486,N_9267);
nand U11398 (N_11398,N_9598,N_8965);
or U11399 (N_11399,N_9391,N_8558);
nand U11400 (N_11400,N_8619,N_9976);
nor U11401 (N_11401,N_8840,N_8217);
nor U11402 (N_11402,N_9764,N_9002);
and U11403 (N_11403,N_8106,N_8416);
or U11404 (N_11404,N_8097,N_8393);
or U11405 (N_11405,N_9850,N_9032);
or U11406 (N_11406,N_9385,N_9425);
nand U11407 (N_11407,N_9858,N_8071);
and U11408 (N_11408,N_9934,N_9174);
or U11409 (N_11409,N_8134,N_8633);
nor U11410 (N_11410,N_9475,N_9508);
or U11411 (N_11411,N_8123,N_9646);
and U11412 (N_11412,N_9923,N_8921);
xor U11413 (N_11413,N_8401,N_9224);
xor U11414 (N_11414,N_9773,N_9180);
nand U11415 (N_11415,N_9784,N_8185);
xor U11416 (N_11416,N_8154,N_9622);
or U11417 (N_11417,N_8598,N_8952);
nor U11418 (N_11418,N_8382,N_8508);
nor U11419 (N_11419,N_9158,N_9169);
nand U11420 (N_11420,N_8285,N_9649);
or U11421 (N_11421,N_9568,N_8709);
nor U11422 (N_11422,N_9621,N_9991);
xor U11423 (N_11423,N_8833,N_9003);
nor U11424 (N_11424,N_8515,N_8317);
xnor U11425 (N_11425,N_9453,N_9172);
xnor U11426 (N_11426,N_8612,N_9837);
and U11427 (N_11427,N_9285,N_8343);
nand U11428 (N_11428,N_9495,N_8164);
nand U11429 (N_11429,N_8806,N_8854);
nand U11430 (N_11430,N_9676,N_9025);
or U11431 (N_11431,N_8489,N_9794);
nand U11432 (N_11432,N_8539,N_8767);
nand U11433 (N_11433,N_9705,N_9884);
or U11434 (N_11434,N_8175,N_8045);
nor U11435 (N_11435,N_9573,N_8629);
nor U11436 (N_11436,N_9572,N_9333);
or U11437 (N_11437,N_8916,N_8155);
or U11438 (N_11438,N_8685,N_9691);
or U11439 (N_11439,N_8813,N_8400);
and U11440 (N_11440,N_8256,N_9351);
nand U11441 (N_11441,N_9839,N_9504);
nor U11442 (N_11442,N_9414,N_8463);
or U11443 (N_11443,N_9431,N_8639);
nor U11444 (N_11444,N_9930,N_9260);
xnor U11445 (N_11445,N_9723,N_8584);
nor U11446 (N_11446,N_9292,N_8439);
nand U11447 (N_11447,N_9780,N_9747);
or U11448 (N_11448,N_8542,N_9854);
nor U11449 (N_11449,N_8197,N_8680);
and U11450 (N_11450,N_8698,N_8818);
nor U11451 (N_11451,N_8745,N_9078);
nand U11452 (N_11452,N_9026,N_9945);
nand U11453 (N_11453,N_9597,N_9792);
or U11454 (N_11454,N_8226,N_9574);
or U11455 (N_11455,N_9887,N_8959);
nor U11456 (N_11456,N_9297,N_9123);
and U11457 (N_11457,N_9606,N_9278);
and U11458 (N_11458,N_8874,N_9726);
and U11459 (N_11459,N_9843,N_9184);
nor U11460 (N_11460,N_8690,N_8163);
nand U11461 (N_11461,N_8705,N_8062);
or U11462 (N_11462,N_9354,N_9084);
or U11463 (N_11463,N_8227,N_9912);
nand U11464 (N_11464,N_8389,N_8273);
nand U11465 (N_11465,N_9141,N_9346);
nand U11466 (N_11466,N_8863,N_8781);
or U11467 (N_11467,N_9430,N_8685);
and U11468 (N_11468,N_8048,N_8384);
and U11469 (N_11469,N_9311,N_8208);
nor U11470 (N_11470,N_8510,N_9929);
nor U11471 (N_11471,N_9445,N_8770);
and U11472 (N_11472,N_9470,N_9165);
xnor U11473 (N_11473,N_9689,N_9478);
or U11474 (N_11474,N_9546,N_9133);
nor U11475 (N_11475,N_8767,N_8213);
and U11476 (N_11476,N_8986,N_9704);
nand U11477 (N_11477,N_8548,N_8946);
or U11478 (N_11478,N_8955,N_9411);
nand U11479 (N_11479,N_8974,N_8404);
or U11480 (N_11480,N_9379,N_8980);
or U11481 (N_11481,N_9544,N_8899);
and U11482 (N_11482,N_8498,N_8435);
or U11483 (N_11483,N_9483,N_8932);
nand U11484 (N_11484,N_8537,N_8232);
and U11485 (N_11485,N_8779,N_9667);
and U11486 (N_11486,N_9708,N_9375);
or U11487 (N_11487,N_9086,N_9876);
and U11488 (N_11488,N_8478,N_8075);
nand U11489 (N_11489,N_9915,N_9905);
xnor U11490 (N_11490,N_9480,N_8479);
and U11491 (N_11491,N_8283,N_9245);
xnor U11492 (N_11492,N_9808,N_8794);
or U11493 (N_11493,N_8887,N_9318);
and U11494 (N_11494,N_9278,N_9192);
or U11495 (N_11495,N_9371,N_8526);
and U11496 (N_11496,N_9794,N_9716);
or U11497 (N_11497,N_8044,N_8654);
and U11498 (N_11498,N_8611,N_9040);
nor U11499 (N_11499,N_8377,N_9638);
xnor U11500 (N_11500,N_9999,N_8029);
and U11501 (N_11501,N_8661,N_8456);
nor U11502 (N_11502,N_9891,N_8330);
nor U11503 (N_11503,N_8312,N_9531);
nor U11504 (N_11504,N_8995,N_9026);
or U11505 (N_11505,N_8187,N_9264);
or U11506 (N_11506,N_9054,N_8073);
xor U11507 (N_11507,N_9357,N_8959);
nand U11508 (N_11508,N_9234,N_8134);
nor U11509 (N_11509,N_9548,N_9251);
or U11510 (N_11510,N_8515,N_9611);
and U11511 (N_11511,N_8330,N_9188);
or U11512 (N_11512,N_8051,N_8657);
or U11513 (N_11513,N_8251,N_8990);
nor U11514 (N_11514,N_8454,N_9250);
or U11515 (N_11515,N_8553,N_9465);
nor U11516 (N_11516,N_9191,N_8966);
nand U11517 (N_11517,N_9821,N_9598);
nand U11518 (N_11518,N_9654,N_9399);
xnor U11519 (N_11519,N_8759,N_9380);
nor U11520 (N_11520,N_9563,N_8007);
and U11521 (N_11521,N_8532,N_8670);
nand U11522 (N_11522,N_9676,N_9122);
or U11523 (N_11523,N_9567,N_8541);
or U11524 (N_11524,N_9202,N_9413);
or U11525 (N_11525,N_8679,N_8592);
nand U11526 (N_11526,N_8366,N_9481);
or U11527 (N_11527,N_8747,N_9863);
and U11528 (N_11528,N_8013,N_8234);
nand U11529 (N_11529,N_8944,N_8549);
nor U11530 (N_11530,N_8661,N_8470);
and U11531 (N_11531,N_9043,N_8662);
and U11532 (N_11532,N_8684,N_9113);
xor U11533 (N_11533,N_9414,N_9544);
and U11534 (N_11534,N_9989,N_8831);
nand U11535 (N_11535,N_8124,N_8810);
and U11536 (N_11536,N_9590,N_9188);
nor U11537 (N_11537,N_9589,N_9265);
or U11538 (N_11538,N_9513,N_9913);
nor U11539 (N_11539,N_8649,N_9910);
nor U11540 (N_11540,N_8849,N_9633);
nand U11541 (N_11541,N_8748,N_9717);
or U11542 (N_11542,N_9149,N_9022);
or U11543 (N_11543,N_8758,N_8908);
xnor U11544 (N_11544,N_9582,N_8221);
nor U11545 (N_11545,N_8854,N_9899);
or U11546 (N_11546,N_8241,N_9063);
or U11547 (N_11547,N_9997,N_9578);
xor U11548 (N_11548,N_8201,N_9776);
nor U11549 (N_11549,N_8086,N_9523);
or U11550 (N_11550,N_9158,N_8853);
nor U11551 (N_11551,N_8408,N_9129);
nor U11552 (N_11552,N_8507,N_9005);
or U11553 (N_11553,N_8133,N_9459);
nand U11554 (N_11554,N_9140,N_8906);
nand U11555 (N_11555,N_9445,N_9178);
and U11556 (N_11556,N_8459,N_9816);
nor U11557 (N_11557,N_8022,N_9475);
nor U11558 (N_11558,N_9352,N_8190);
or U11559 (N_11559,N_8290,N_9927);
and U11560 (N_11560,N_9618,N_8038);
and U11561 (N_11561,N_9112,N_9008);
or U11562 (N_11562,N_9660,N_8737);
and U11563 (N_11563,N_9191,N_9275);
xor U11564 (N_11564,N_9405,N_9595);
or U11565 (N_11565,N_9820,N_8611);
xnor U11566 (N_11566,N_9066,N_8216);
or U11567 (N_11567,N_8632,N_9459);
nand U11568 (N_11568,N_8665,N_9083);
or U11569 (N_11569,N_9512,N_9484);
or U11570 (N_11570,N_9891,N_9196);
or U11571 (N_11571,N_9705,N_8446);
and U11572 (N_11572,N_9901,N_9421);
nor U11573 (N_11573,N_8646,N_9392);
or U11574 (N_11574,N_9455,N_8119);
or U11575 (N_11575,N_8720,N_8204);
and U11576 (N_11576,N_8197,N_8377);
nor U11577 (N_11577,N_9850,N_8875);
and U11578 (N_11578,N_9721,N_8827);
nand U11579 (N_11579,N_8454,N_8234);
nor U11580 (N_11580,N_9962,N_8274);
or U11581 (N_11581,N_8760,N_8966);
nand U11582 (N_11582,N_9440,N_9171);
or U11583 (N_11583,N_9524,N_8506);
nand U11584 (N_11584,N_9902,N_9063);
nand U11585 (N_11585,N_8697,N_8549);
nor U11586 (N_11586,N_9009,N_9731);
and U11587 (N_11587,N_8478,N_9463);
xnor U11588 (N_11588,N_8611,N_9965);
nor U11589 (N_11589,N_9730,N_8031);
or U11590 (N_11590,N_8054,N_8078);
and U11591 (N_11591,N_9433,N_8569);
or U11592 (N_11592,N_9904,N_8252);
or U11593 (N_11593,N_8048,N_9932);
nand U11594 (N_11594,N_8944,N_8877);
nor U11595 (N_11595,N_8304,N_8571);
nor U11596 (N_11596,N_9114,N_9082);
nor U11597 (N_11597,N_8303,N_8669);
xor U11598 (N_11598,N_9435,N_9160);
or U11599 (N_11599,N_9391,N_9091);
or U11600 (N_11600,N_8004,N_8044);
and U11601 (N_11601,N_9299,N_8270);
xor U11602 (N_11602,N_9649,N_9556);
nor U11603 (N_11603,N_8297,N_9625);
xor U11604 (N_11604,N_9469,N_8821);
nand U11605 (N_11605,N_9670,N_9956);
or U11606 (N_11606,N_9758,N_8070);
and U11607 (N_11607,N_9920,N_9838);
and U11608 (N_11608,N_9698,N_9376);
nand U11609 (N_11609,N_9699,N_8668);
xor U11610 (N_11610,N_9106,N_8102);
nor U11611 (N_11611,N_8880,N_8322);
or U11612 (N_11612,N_9142,N_9998);
nor U11613 (N_11613,N_9517,N_8964);
and U11614 (N_11614,N_8585,N_8141);
or U11615 (N_11615,N_8365,N_9224);
or U11616 (N_11616,N_9568,N_9721);
and U11617 (N_11617,N_8211,N_9563);
or U11618 (N_11618,N_8260,N_8905);
and U11619 (N_11619,N_8956,N_8495);
nand U11620 (N_11620,N_9164,N_8089);
and U11621 (N_11621,N_8755,N_8171);
or U11622 (N_11622,N_8984,N_9285);
nand U11623 (N_11623,N_8728,N_9332);
nor U11624 (N_11624,N_8741,N_9029);
nand U11625 (N_11625,N_8276,N_9375);
xor U11626 (N_11626,N_9223,N_8725);
nor U11627 (N_11627,N_8115,N_8346);
or U11628 (N_11628,N_8016,N_8979);
nand U11629 (N_11629,N_9519,N_8396);
xor U11630 (N_11630,N_9181,N_9547);
nand U11631 (N_11631,N_8817,N_8509);
nand U11632 (N_11632,N_9165,N_9887);
and U11633 (N_11633,N_8892,N_9555);
or U11634 (N_11634,N_9230,N_9862);
xor U11635 (N_11635,N_8090,N_8612);
and U11636 (N_11636,N_8244,N_9385);
or U11637 (N_11637,N_9210,N_9960);
and U11638 (N_11638,N_9154,N_9350);
nand U11639 (N_11639,N_8928,N_9654);
and U11640 (N_11640,N_8468,N_9838);
or U11641 (N_11641,N_9922,N_9482);
nand U11642 (N_11642,N_8678,N_8931);
nor U11643 (N_11643,N_8919,N_9002);
or U11644 (N_11644,N_9768,N_9448);
xnor U11645 (N_11645,N_9143,N_9086);
nand U11646 (N_11646,N_8805,N_9987);
nand U11647 (N_11647,N_9134,N_9728);
nand U11648 (N_11648,N_8995,N_8217);
or U11649 (N_11649,N_9596,N_9077);
or U11650 (N_11650,N_9102,N_8319);
nor U11651 (N_11651,N_9772,N_8790);
and U11652 (N_11652,N_8310,N_8384);
nor U11653 (N_11653,N_9115,N_9989);
or U11654 (N_11654,N_8999,N_8125);
or U11655 (N_11655,N_8932,N_9434);
nor U11656 (N_11656,N_9560,N_8336);
nand U11657 (N_11657,N_9210,N_9314);
and U11658 (N_11658,N_8328,N_8871);
nand U11659 (N_11659,N_8919,N_9920);
nand U11660 (N_11660,N_9654,N_8341);
or U11661 (N_11661,N_8962,N_8903);
nand U11662 (N_11662,N_9104,N_9723);
nor U11663 (N_11663,N_9891,N_9916);
and U11664 (N_11664,N_9204,N_9803);
nor U11665 (N_11665,N_9695,N_8555);
nor U11666 (N_11666,N_8684,N_8865);
xnor U11667 (N_11667,N_8917,N_9393);
and U11668 (N_11668,N_9926,N_9435);
and U11669 (N_11669,N_8330,N_9970);
and U11670 (N_11670,N_8532,N_8524);
and U11671 (N_11671,N_8058,N_8899);
nor U11672 (N_11672,N_9807,N_8098);
xor U11673 (N_11673,N_8837,N_9758);
and U11674 (N_11674,N_8123,N_8607);
nor U11675 (N_11675,N_8707,N_9670);
and U11676 (N_11676,N_8064,N_8814);
and U11677 (N_11677,N_9391,N_9133);
nor U11678 (N_11678,N_9868,N_8715);
and U11679 (N_11679,N_8696,N_9797);
or U11680 (N_11680,N_8627,N_9902);
nor U11681 (N_11681,N_8851,N_9677);
or U11682 (N_11682,N_8178,N_8664);
or U11683 (N_11683,N_8649,N_9815);
nand U11684 (N_11684,N_9933,N_9760);
or U11685 (N_11685,N_9780,N_8996);
and U11686 (N_11686,N_9504,N_8755);
or U11687 (N_11687,N_8988,N_9439);
xor U11688 (N_11688,N_9154,N_9998);
xor U11689 (N_11689,N_9239,N_9449);
xor U11690 (N_11690,N_9381,N_8719);
and U11691 (N_11691,N_9842,N_9529);
nand U11692 (N_11692,N_8931,N_8212);
nor U11693 (N_11693,N_9581,N_8080);
xor U11694 (N_11694,N_8307,N_9011);
and U11695 (N_11695,N_9446,N_9375);
xnor U11696 (N_11696,N_9762,N_8042);
or U11697 (N_11697,N_8191,N_8018);
nand U11698 (N_11698,N_9338,N_8158);
and U11699 (N_11699,N_8153,N_9111);
nor U11700 (N_11700,N_9562,N_9740);
nand U11701 (N_11701,N_8788,N_8646);
nand U11702 (N_11702,N_8104,N_8383);
xnor U11703 (N_11703,N_9498,N_9954);
and U11704 (N_11704,N_9604,N_9482);
nand U11705 (N_11705,N_9042,N_8963);
nor U11706 (N_11706,N_9520,N_8592);
or U11707 (N_11707,N_8518,N_8264);
xor U11708 (N_11708,N_8615,N_9204);
or U11709 (N_11709,N_9409,N_9874);
nor U11710 (N_11710,N_8118,N_9626);
xor U11711 (N_11711,N_9099,N_8813);
nand U11712 (N_11712,N_9837,N_8352);
or U11713 (N_11713,N_9681,N_8796);
and U11714 (N_11714,N_8443,N_8120);
or U11715 (N_11715,N_8738,N_9287);
or U11716 (N_11716,N_8683,N_9285);
nor U11717 (N_11717,N_9197,N_8231);
or U11718 (N_11718,N_8074,N_8767);
and U11719 (N_11719,N_9427,N_9066);
nand U11720 (N_11720,N_9925,N_8711);
and U11721 (N_11721,N_8641,N_8781);
or U11722 (N_11722,N_9760,N_8745);
nand U11723 (N_11723,N_9630,N_8471);
or U11724 (N_11724,N_8563,N_9663);
or U11725 (N_11725,N_8048,N_8205);
and U11726 (N_11726,N_8035,N_8456);
or U11727 (N_11727,N_8007,N_9335);
nor U11728 (N_11728,N_8961,N_9499);
xnor U11729 (N_11729,N_9518,N_8622);
xor U11730 (N_11730,N_9058,N_9021);
nand U11731 (N_11731,N_9462,N_9393);
or U11732 (N_11732,N_8099,N_9906);
or U11733 (N_11733,N_8217,N_9495);
and U11734 (N_11734,N_8607,N_8545);
or U11735 (N_11735,N_8412,N_9525);
nor U11736 (N_11736,N_9835,N_8717);
xnor U11737 (N_11737,N_8042,N_8863);
nor U11738 (N_11738,N_8253,N_9343);
or U11739 (N_11739,N_9007,N_8963);
nor U11740 (N_11740,N_9310,N_8670);
or U11741 (N_11741,N_9825,N_8004);
nor U11742 (N_11742,N_9305,N_9812);
nor U11743 (N_11743,N_8332,N_8857);
nor U11744 (N_11744,N_9674,N_9737);
nand U11745 (N_11745,N_9301,N_9536);
nand U11746 (N_11746,N_9981,N_8560);
nand U11747 (N_11747,N_9930,N_9849);
or U11748 (N_11748,N_9624,N_9818);
or U11749 (N_11749,N_8121,N_8774);
or U11750 (N_11750,N_9985,N_8867);
or U11751 (N_11751,N_9794,N_9989);
or U11752 (N_11752,N_9268,N_9552);
nand U11753 (N_11753,N_9166,N_8889);
or U11754 (N_11754,N_8433,N_8032);
and U11755 (N_11755,N_9675,N_8275);
or U11756 (N_11756,N_9500,N_9938);
xor U11757 (N_11757,N_9339,N_9878);
nor U11758 (N_11758,N_8097,N_9069);
nor U11759 (N_11759,N_8336,N_9736);
or U11760 (N_11760,N_9566,N_8388);
nor U11761 (N_11761,N_9034,N_8825);
and U11762 (N_11762,N_9299,N_9860);
nor U11763 (N_11763,N_8691,N_9860);
or U11764 (N_11764,N_9598,N_8543);
xnor U11765 (N_11765,N_8438,N_8762);
or U11766 (N_11766,N_9961,N_8905);
or U11767 (N_11767,N_9783,N_8309);
nand U11768 (N_11768,N_9389,N_8660);
or U11769 (N_11769,N_9077,N_9103);
nor U11770 (N_11770,N_8317,N_9500);
or U11771 (N_11771,N_8404,N_9829);
and U11772 (N_11772,N_8111,N_8294);
and U11773 (N_11773,N_8100,N_8994);
and U11774 (N_11774,N_8062,N_8722);
nand U11775 (N_11775,N_8316,N_9722);
nand U11776 (N_11776,N_8991,N_8689);
xnor U11777 (N_11777,N_9866,N_9273);
nor U11778 (N_11778,N_8511,N_8137);
and U11779 (N_11779,N_8089,N_8302);
nor U11780 (N_11780,N_8157,N_8976);
nor U11781 (N_11781,N_8693,N_8254);
nand U11782 (N_11782,N_9831,N_8316);
nand U11783 (N_11783,N_8379,N_9943);
or U11784 (N_11784,N_8098,N_8993);
nand U11785 (N_11785,N_9389,N_8398);
nor U11786 (N_11786,N_9747,N_9371);
nand U11787 (N_11787,N_8060,N_9186);
xnor U11788 (N_11788,N_8939,N_8602);
xor U11789 (N_11789,N_9536,N_9040);
or U11790 (N_11790,N_8730,N_9912);
and U11791 (N_11791,N_9494,N_9189);
or U11792 (N_11792,N_8746,N_8462);
nand U11793 (N_11793,N_8693,N_8815);
nand U11794 (N_11794,N_9966,N_9212);
or U11795 (N_11795,N_8976,N_8282);
or U11796 (N_11796,N_9453,N_9312);
or U11797 (N_11797,N_8049,N_8693);
or U11798 (N_11798,N_8076,N_8021);
nor U11799 (N_11799,N_8390,N_8818);
nor U11800 (N_11800,N_8437,N_9704);
nand U11801 (N_11801,N_8099,N_8866);
nand U11802 (N_11802,N_9932,N_8891);
or U11803 (N_11803,N_9911,N_9062);
nand U11804 (N_11804,N_8989,N_9494);
and U11805 (N_11805,N_8957,N_8276);
or U11806 (N_11806,N_9572,N_8394);
nand U11807 (N_11807,N_8018,N_8821);
and U11808 (N_11808,N_8361,N_9718);
nor U11809 (N_11809,N_8634,N_8798);
nand U11810 (N_11810,N_8335,N_8798);
nor U11811 (N_11811,N_9260,N_8082);
and U11812 (N_11812,N_8107,N_8971);
nand U11813 (N_11813,N_8491,N_8394);
nor U11814 (N_11814,N_8791,N_8881);
or U11815 (N_11815,N_8291,N_8991);
or U11816 (N_11816,N_9477,N_8770);
nor U11817 (N_11817,N_8143,N_9326);
nor U11818 (N_11818,N_9293,N_9676);
and U11819 (N_11819,N_8178,N_9986);
nor U11820 (N_11820,N_9659,N_9078);
nor U11821 (N_11821,N_8228,N_8388);
or U11822 (N_11822,N_9069,N_9829);
and U11823 (N_11823,N_8931,N_8301);
and U11824 (N_11824,N_9353,N_9290);
or U11825 (N_11825,N_8464,N_8105);
and U11826 (N_11826,N_8703,N_9515);
or U11827 (N_11827,N_8639,N_9678);
xnor U11828 (N_11828,N_9153,N_9882);
xor U11829 (N_11829,N_9489,N_8639);
and U11830 (N_11830,N_9170,N_9330);
or U11831 (N_11831,N_8388,N_8236);
or U11832 (N_11832,N_9161,N_8054);
or U11833 (N_11833,N_8107,N_8780);
xnor U11834 (N_11834,N_8130,N_9373);
and U11835 (N_11835,N_9386,N_9050);
or U11836 (N_11836,N_8050,N_9757);
or U11837 (N_11837,N_9981,N_8716);
xor U11838 (N_11838,N_8672,N_8112);
nand U11839 (N_11839,N_9868,N_9497);
nor U11840 (N_11840,N_8283,N_9277);
nand U11841 (N_11841,N_9373,N_9327);
nand U11842 (N_11842,N_9490,N_9191);
or U11843 (N_11843,N_9428,N_9257);
and U11844 (N_11844,N_9899,N_9060);
or U11845 (N_11845,N_9128,N_8982);
and U11846 (N_11846,N_8103,N_9629);
xnor U11847 (N_11847,N_9400,N_9594);
nor U11848 (N_11848,N_8744,N_9697);
nor U11849 (N_11849,N_9983,N_8789);
and U11850 (N_11850,N_8296,N_9097);
nor U11851 (N_11851,N_8096,N_9896);
nand U11852 (N_11852,N_9568,N_9523);
nand U11853 (N_11853,N_9175,N_9959);
nand U11854 (N_11854,N_8742,N_8952);
xnor U11855 (N_11855,N_8100,N_9160);
and U11856 (N_11856,N_8592,N_8883);
or U11857 (N_11857,N_9806,N_8947);
nand U11858 (N_11858,N_8019,N_9835);
nor U11859 (N_11859,N_9479,N_9303);
or U11860 (N_11860,N_8201,N_9880);
and U11861 (N_11861,N_9711,N_8827);
and U11862 (N_11862,N_9923,N_9179);
or U11863 (N_11863,N_9405,N_9926);
or U11864 (N_11864,N_8067,N_9807);
and U11865 (N_11865,N_9020,N_9054);
nor U11866 (N_11866,N_9098,N_9062);
or U11867 (N_11867,N_9245,N_8537);
and U11868 (N_11868,N_9499,N_9834);
nand U11869 (N_11869,N_8313,N_8445);
and U11870 (N_11870,N_9666,N_8072);
or U11871 (N_11871,N_9654,N_8080);
and U11872 (N_11872,N_9176,N_8647);
nand U11873 (N_11873,N_9964,N_8770);
or U11874 (N_11874,N_9532,N_8815);
xnor U11875 (N_11875,N_9388,N_9818);
or U11876 (N_11876,N_9248,N_9308);
nand U11877 (N_11877,N_9282,N_9710);
nor U11878 (N_11878,N_9773,N_8046);
and U11879 (N_11879,N_8537,N_9823);
or U11880 (N_11880,N_8642,N_9357);
or U11881 (N_11881,N_8120,N_9253);
nand U11882 (N_11882,N_9224,N_9118);
or U11883 (N_11883,N_9720,N_9257);
nand U11884 (N_11884,N_9010,N_8860);
nor U11885 (N_11885,N_9188,N_9212);
and U11886 (N_11886,N_8405,N_9471);
or U11887 (N_11887,N_9074,N_8793);
and U11888 (N_11888,N_8209,N_9333);
nor U11889 (N_11889,N_8534,N_9774);
and U11890 (N_11890,N_8995,N_8127);
nor U11891 (N_11891,N_8639,N_9176);
xor U11892 (N_11892,N_8847,N_9331);
nor U11893 (N_11893,N_9672,N_8729);
or U11894 (N_11894,N_8766,N_8165);
or U11895 (N_11895,N_8877,N_9066);
and U11896 (N_11896,N_9026,N_8429);
xnor U11897 (N_11897,N_9098,N_9746);
nand U11898 (N_11898,N_8740,N_9844);
and U11899 (N_11899,N_8560,N_9740);
and U11900 (N_11900,N_8896,N_9278);
nor U11901 (N_11901,N_9742,N_9120);
or U11902 (N_11902,N_9196,N_9694);
or U11903 (N_11903,N_8466,N_8082);
and U11904 (N_11904,N_8673,N_9594);
xnor U11905 (N_11905,N_9607,N_9687);
xnor U11906 (N_11906,N_9312,N_9825);
nor U11907 (N_11907,N_8633,N_8333);
nor U11908 (N_11908,N_8811,N_9569);
and U11909 (N_11909,N_9347,N_9791);
nand U11910 (N_11910,N_8438,N_8901);
nand U11911 (N_11911,N_9276,N_8085);
nor U11912 (N_11912,N_9572,N_9282);
xor U11913 (N_11913,N_9729,N_8194);
xor U11914 (N_11914,N_9612,N_8317);
nand U11915 (N_11915,N_9694,N_9284);
nor U11916 (N_11916,N_9467,N_8201);
nand U11917 (N_11917,N_8736,N_8275);
nand U11918 (N_11918,N_9379,N_9681);
nand U11919 (N_11919,N_8701,N_9444);
nor U11920 (N_11920,N_9064,N_9495);
nand U11921 (N_11921,N_8672,N_9377);
nand U11922 (N_11922,N_8034,N_9570);
or U11923 (N_11923,N_8678,N_9331);
or U11924 (N_11924,N_9129,N_8399);
or U11925 (N_11925,N_9692,N_8218);
nand U11926 (N_11926,N_9398,N_8107);
and U11927 (N_11927,N_9396,N_8692);
nor U11928 (N_11928,N_9474,N_9445);
or U11929 (N_11929,N_9541,N_8546);
or U11930 (N_11930,N_9183,N_9046);
nand U11931 (N_11931,N_9618,N_9144);
or U11932 (N_11932,N_9403,N_8011);
and U11933 (N_11933,N_8382,N_9493);
or U11934 (N_11934,N_8641,N_9005);
or U11935 (N_11935,N_8045,N_9570);
nor U11936 (N_11936,N_8991,N_9213);
nand U11937 (N_11937,N_9187,N_8058);
xnor U11938 (N_11938,N_8027,N_9850);
nor U11939 (N_11939,N_9564,N_8630);
nand U11940 (N_11940,N_8705,N_9200);
nand U11941 (N_11941,N_8782,N_9907);
and U11942 (N_11942,N_8575,N_9991);
and U11943 (N_11943,N_8282,N_8771);
nand U11944 (N_11944,N_9360,N_9341);
xor U11945 (N_11945,N_9979,N_9628);
nor U11946 (N_11946,N_8296,N_9082);
or U11947 (N_11947,N_9988,N_8058);
nor U11948 (N_11948,N_9481,N_8894);
or U11949 (N_11949,N_8068,N_8953);
or U11950 (N_11950,N_9052,N_8084);
nor U11951 (N_11951,N_9825,N_8836);
nor U11952 (N_11952,N_8020,N_8606);
and U11953 (N_11953,N_8478,N_8421);
and U11954 (N_11954,N_8346,N_9241);
nand U11955 (N_11955,N_9456,N_8405);
nor U11956 (N_11956,N_8197,N_8618);
or U11957 (N_11957,N_8370,N_9600);
nand U11958 (N_11958,N_8160,N_9166);
or U11959 (N_11959,N_8366,N_9830);
nor U11960 (N_11960,N_9153,N_8579);
or U11961 (N_11961,N_8013,N_8266);
or U11962 (N_11962,N_9475,N_9207);
nand U11963 (N_11963,N_9106,N_9157);
or U11964 (N_11964,N_8532,N_8700);
and U11965 (N_11965,N_9495,N_9301);
nor U11966 (N_11966,N_9771,N_9512);
nor U11967 (N_11967,N_8716,N_8447);
or U11968 (N_11968,N_9595,N_8737);
nand U11969 (N_11969,N_9312,N_9205);
xnor U11970 (N_11970,N_8201,N_8755);
and U11971 (N_11971,N_8696,N_8986);
nor U11972 (N_11972,N_9693,N_9740);
nand U11973 (N_11973,N_8171,N_8929);
and U11974 (N_11974,N_8802,N_9318);
and U11975 (N_11975,N_8726,N_9005);
or U11976 (N_11976,N_8343,N_9043);
nor U11977 (N_11977,N_9667,N_9919);
and U11978 (N_11978,N_8011,N_8883);
nand U11979 (N_11979,N_9076,N_8720);
nor U11980 (N_11980,N_8953,N_8518);
and U11981 (N_11981,N_9710,N_8223);
nand U11982 (N_11982,N_8311,N_8675);
and U11983 (N_11983,N_8149,N_9649);
or U11984 (N_11984,N_8442,N_9241);
or U11985 (N_11985,N_9080,N_8663);
nand U11986 (N_11986,N_8495,N_9231);
nor U11987 (N_11987,N_8334,N_9538);
or U11988 (N_11988,N_8480,N_9363);
and U11989 (N_11989,N_9857,N_9423);
nor U11990 (N_11990,N_8294,N_9063);
and U11991 (N_11991,N_8519,N_8701);
or U11992 (N_11992,N_8829,N_8876);
or U11993 (N_11993,N_8979,N_8645);
nand U11994 (N_11994,N_8031,N_9907);
nand U11995 (N_11995,N_9585,N_9199);
nor U11996 (N_11996,N_9007,N_8688);
nand U11997 (N_11997,N_9850,N_8650);
nor U11998 (N_11998,N_9319,N_8001);
xnor U11999 (N_11999,N_9811,N_8011);
or U12000 (N_12000,N_11074,N_10684);
or U12001 (N_12001,N_11217,N_11053);
nor U12002 (N_12002,N_10976,N_10756);
and U12003 (N_12003,N_11834,N_11429);
and U12004 (N_12004,N_10545,N_11489);
xor U12005 (N_12005,N_11818,N_11430);
or U12006 (N_12006,N_10941,N_10900);
nor U12007 (N_12007,N_10642,N_11092);
and U12008 (N_12008,N_10554,N_11690);
or U12009 (N_12009,N_11778,N_10062);
or U12010 (N_12010,N_11722,N_11970);
or U12011 (N_12011,N_10481,N_11601);
xor U12012 (N_12012,N_10455,N_11120);
and U12013 (N_12013,N_11898,N_11290);
and U12014 (N_12014,N_10166,N_11638);
and U12015 (N_12015,N_11569,N_10274);
or U12016 (N_12016,N_10237,N_10435);
and U12017 (N_12017,N_11617,N_10712);
and U12018 (N_12018,N_10946,N_10624);
or U12019 (N_12019,N_11312,N_10602);
and U12020 (N_12020,N_10326,N_10551);
nor U12021 (N_12021,N_10560,N_10557);
or U12022 (N_12022,N_11226,N_11990);
nor U12023 (N_12023,N_10936,N_10484);
nor U12024 (N_12024,N_11713,N_10760);
nand U12025 (N_12025,N_11014,N_11697);
or U12026 (N_12026,N_10812,N_11067);
nor U12027 (N_12027,N_11519,N_11740);
nor U12028 (N_12028,N_11339,N_10650);
and U12029 (N_12029,N_11329,N_11321);
nor U12030 (N_12030,N_10857,N_11622);
and U12031 (N_12031,N_11841,N_10352);
or U12032 (N_12032,N_10988,N_11694);
or U12033 (N_12033,N_11300,N_11018);
and U12034 (N_12034,N_11753,N_11931);
or U12035 (N_12035,N_10828,N_10165);
and U12036 (N_12036,N_10821,N_11106);
and U12037 (N_12037,N_10771,N_10395);
and U12038 (N_12038,N_10945,N_10409);
nand U12039 (N_12039,N_11468,N_11550);
nor U12040 (N_12040,N_10553,N_11806);
xor U12041 (N_12041,N_10788,N_10232);
nor U12042 (N_12042,N_10518,N_11775);
nand U12043 (N_12043,N_10718,N_10790);
and U12044 (N_12044,N_10468,N_10669);
nor U12045 (N_12045,N_10851,N_11835);
or U12046 (N_12046,N_10618,N_11234);
or U12047 (N_12047,N_10499,N_10569);
or U12048 (N_12048,N_11409,N_11153);
xnor U12049 (N_12049,N_11041,N_10065);
xor U12050 (N_12050,N_10411,N_11735);
or U12051 (N_12051,N_10447,N_11207);
nand U12052 (N_12052,N_10928,N_11703);
and U12053 (N_12053,N_11221,N_11439);
nand U12054 (N_12054,N_11431,N_11619);
nor U12055 (N_12055,N_10283,N_11864);
and U12056 (N_12056,N_11802,N_11559);
and U12057 (N_12057,N_11073,N_10391);
nand U12058 (N_12058,N_11228,N_11317);
nor U12059 (N_12059,N_11257,N_10994);
nand U12060 (N_12060,N_11664,N_11170);
nor U12061 (N_12061,N_11936,N_10972);
nor U12062 (N_12062,N_11705,N_11318);
nor U12063 (N_12063,N_11050,N_11309);
nand U12064 (N_12064,N_11680,N_11253);
and U12065 (N_12065,N_11245,N_10182);
nand U12066 (N_12066,N_10498,N_10504);
and U12067 (N_12067,N_10501,N_11404);
or U12068 (N_12068,N_11255,N_10987);
or U12069 (N_12069,N_11260,N_10451);
or U12070 (N_12070,N_10735,N_10933);
nand U12071 (N_12071,N_10920,N_11525);
or U12072 (N_12072,N_11296,N_10862);
xnor U12073 (N_12073,N_10750,N_11032);
nor U12074 (N_12074,N_11646,N_11417);
and U12075 (N_12075,N_11425,N_10815);
nand U12076 (N_12076,N_10161,N_10121);
and U12077 (N_12077,N_10886,N_11536);
and U12078 (N_12078,N_10369,N_10893);
and U12079 (N_12079,N_11797,N_10691);
nor U12080 (N_12080,N_11975,N_11408);
nand U12081 (N_12081,N_11169,N_10172);
xnor U12082 (N_12082,N_10427,N_10915);
nand U12083 (N_12083,N_11395,N_11564);
and U12084 (N_12084,N_10874,N_10983);
or U12085 (N_12085,N_10526,N_10654);
nor U12086 (N_12086,N_11803,N_11514);
or U12087 (N_12087,N_10977,N_11055);
and U12088 (N_12088,N_10826,N_11526);
nand U12089 (N_12089,N_11322,N_10860);
or U12090 (N_12090,N_11668,N_10007);
nor U12091 (N_12091,N_11266,N_11289);
nand U12092 (N_12092,N_10752,N_10548);
nor U12093 (N_12093,N_11866,N_10599);
and U12094 (N_12094,N_10377,N_10998);
and U12095 (N_12095,N_10903,N_10677);
and U12096 (N_12096,N_11469,N_11575);
or U12097 (N_12097,N_11028,N_10861);
xnor U12098 (N_12098,N_10048,N_10025);
xor U12099 (N_12099,N_11412,N_10350);
nor U12100 (N_12100,N_10619,N_10533);
or U12101 (N_12101,N_10895,N_11886);
and U12102 (N_12102,N_10600,N_10187);
and U12103 (N_12103,N_10690,N_11381);
xor U12104 (N_12104,N_11655,N_10367);
xor U12105 (N_12105,N_10939,N_10622);
and U12106 (N_12106,N_11667,N_10434);
nand U12107 (N_12107,N_10576,N_10050);
or U12108 (N_12108,N_10470,N_10797);
nand U12109 (N_12109,N_10613,N_11952);
nor U12110 (N_12110,N_11534,N_11872);
xor U12111 (N_12111,N_11472,N_11214);
xnor U12112 (N_12112,N_10016,N_10316);
and U12113 (N_12113,N_10102,N_11467);
and U12114 (N_12114,N_11024,N_11000);
or U12115 (N_12115,N_11710,N_10767);
and U12116 (N_12116,N_11552,N_10272);
nor U12117 (N_12117,N_10761,N_11611);
and U12118 (N_12118,N_10625,N_10399);
nor U12119 (N_12119,N_11428,N_11083);
nor U12120 (N_12120,N_10734,N_11268);
and U12121 (N_12121,N_11200,N_11861);
or U12122 (N_12122,N_10170,N_10015);
xor U12123 (N_12123,N_11440,N_11167);
nand U12124 (N_12124,N_11019,N_11565);
nor U12125 (N_12125,N_11356,N_10889);
or U12126 (N_12126,N_11093,N_11874);
and U12127 (N_12127,N_10478,N_11549);
nor U12128 (N_12128,N_10355,N_10227);
and U12129 (N_12129,N_10241,N_10985);
or U12130 (N_12130,N_10331,N_11855);
nand U12131 (N_12131,N_11635,N_11567);
nand U12132 (N_12132,N_10702,N_11963);
xor U12133 (N_12133,N_11711,N_10280);
and U12134 (N_12134,N_11695,N_10133);
nand U12135 (N_12135,N_11513,N_11940);
nor U12136 (N_12136,N_10014,N_11971);
nand U12137 (N_12137,N_10595,N_10009);
xor U12138 (N_12138,N_11572,N_11660);
or U12139 (N_12139,N_11117,N_10728);
nand U12140 (N_12140,N_10175,N_11299);
nand U12141 (N_12141,N_11029,N_11726);
and U12142 (N_12142,N_10726,N_11235);
or U12143 (N_12143,N_10151,N_10781);
nand U12144 (N_12144,N_11026,N_10343);
nand U12145 (N_12145,N_10366,N_11754);
nand U12146 (N_12146,N_11605,N_10219);
or U12147 (N_12147,N_11478,N_10229);
or U12148 (N_12148,N_10611,N_10858);
nor U12149 (N_12149,N_11663,N_11085);
nand U12150 (N_12150,N_10466,N_11424);
nor U12151 (N_12151,N_11091,N_10603);
or U12152 (N_12152,N_11807,N_10070);
nand U12153 (N_12153,N_10419,N_10104);
or U12154 (N_12154,N_11479,N_11491);
nor U12155 (N_12155,N_10824,N_11293);
or U12156 (N_12156,N_11282,N_11691);
or U12157 (N_12157,N_11744,N_10829);
and U12158 (N_12158,N_10268,N_10672);
nand U12159 (N_12159,N_11320,N_10615);
or U12160 (N_12160,N_11810,N_11328);
xnor U12161 (N_12161,N_11361,N_10055);
or U12162 (N_12162,N_11910,N_10745);
and U12163 (N_12163,N_11331,N_10944);
nor U12164 (N_12164,N_11865,N_10527);
and U12165 (N_12165,N_11079,N_10281);
xnor U12166 (N_12166,N_10278,N_10666);
or U12167 (N_12167,N_11851,N_11977);
nor U12168 (N_12168,N_10271,N_11881);
or U12169 (N_12169,N_11808,N_10679);
nand U12170 (N_12170,N_10032,N_10086);
nor U12171 (N_12171,N_10778,N_11517);
nor U12172 (N_12172,N_10100,N_11627);
nand U12173 (N_12173,N_10585,N_10688);
and U12174 (N_12174,N_11890,N_11352);
and U12175 (N_12175,N_11259,N_10233);
and U12176 (N_12176,N_10510,N_10968);
and U12177 (N_12177,N_11893,N_10221);
nand U12178 (N_12178,N_10480,N_11887);
nand U12179 (N_12179,N_11162,N_10975);
xnor U12180 (N_12180,N_11670,N_10730);
and U12181 (N_12181,N_11480,N_11750);
nand U12182 (N_12182,N_10795,N_11728);
nand U12183 (N_12183,N_11801,N_11107);
xor U12184 (N_12184,N_11791,N_11347);
or U12185 (N_12185,N_10774,N_11578);
nor U12186 (N_12186,N_11845,N_10040);
and U12187 (N_12187,N_11508,N_11109);
nor U12188 (N_12188,N_11758,N_10899);
nand U12189 (N_12189,N_11626,N_10514);
and U12190 (N_12190,N_11579,N_11943);
and U12191 (N_12191,N_11315,N_10964);
nor U12192 (N_12192,N_10380,N_10635);
and U12193 (N_12193,N_11701,N_11856);
nor U12194 (N_12194,N_11637,N_11860);
nor U12195 (N_12195,N_11685,N_10827);
and U12196 (N_12196,N_11964,N_11606);
nor U12197 (N_12197,N_11100,N_10562);
xor U12198 (N_12198,N_10064,N_10808);
nand U12199 (N_12199,N_11288,N_10888);
nand U12200 (N_12200,N_10246,N_11741);
and U12201 (N_12201,N_10191,N_11270);
nand U12202 (N_12202,N_10969,N_10661);
nor U12203 (N_12203,N_11367,N_11189);
or U12204 (N_12204,N_10436,N_11548);
and U12205 (N_12205,N_10907,N_11190);
nor U12206 (N_12206,N_11607,N_11337);
and U12207 (N_12207,N_11209,N_10142);
nor U12208 (N_12208,N_10565,N_11850);
nor U12209 (N_12209,N_11516,N_10674);
nor U12210 (N_12210,N_11389,N_10739);
nand U12211 (N_12211,N_10646,N_10573);
and U12212 (N_12212,N_10365,N_11244);
or U12213 (N_12213,N_10073,N_11927);
nor U12214 (N_12214,N_10426,N_11166);
or U12215 (N_12215,N_10906,N_11124);
and U12216 (N_12216,N_11644,N_10584);
and U12217 (N_12217,N_11999,N_11144);
nor U12218 (N_12218,N_11277,N_11949);
xnor U12219 (N_12219,N_11651,N_10692);
xor U12220 (N_12220,N_10444,N_10564);
or U12221 (N_12221,N_10962,N_10437);
or U12222 (N_12222,N_10793,N_10115);
nor U12223 (N_12223,N_10189,N_11991);
nand U12224 (N_12224,N_10430,N_10556);
or U12225 (N_12225,N_10494,N_11016);
nand U12226 (N_12226,N_10522,N_11995);
nand U12227 (N_12227,N_10277,N_10623);
and U12228 (N_12228,N_11973,N_10333);
nor U12229 (N_12229,N_11133,N_11362);
nand U12230 (N_12230,N_11507,N_10974);
or U12231 (N_12231,N_11847,N_11836);
nand U12232 (N_12232,N_11043,N_10013);
and U12233 (N_12233,N_11471,N_10817);
and U12234 (N_12234,N_10568,N_11585);
and U12235 (N_12235,N_11199,N_10762);
nand U12236 (N_12236,N_10226,N_10461);
nor U12237 (N_12237,N_11933,N_11267);
nand U12238 (N_12238,N_11707,N_11984);
or U12239 (N_12239,N_11901,N_10413);
and U12240 (N_12240,N_11399,N_10183);
or U12241 (N_12241,N_11979,N_10396);
xnor U12242 (N_12242,N_10604,N_11348);
nor U12243 (N_12243,N_10748,N_11538);
nor U12244 (N_12244,N_11563,N_10741);
nor U12245 (N_12245,N_10483,N_10587);
nand U12246 (N_12246,N_11105,N_10539);
nand U12247 (N_12247,N_11463,N_10495);
xnor U12248 (N_12248,N_10432,N_11415);
and U12249 (N_12249,N_10833,N_11344);
and U12250 (N_12250,N_11139,N_11176);
nor U12251 (N_12251,N_11388,N_11966);
nand U12252 (N_12252,N_11110,N_11600);
nor U12253 (N_12253,N_10317,N_10856);
and U12254 (N_12254,N_10417,N_11980);
nand U12255 (N_12255,N_10534,N_10109);
nor U12256 (N_12256,N_10608,N_10908);
nand U12257 (N_12257,N_10563,N_11152);
or U12258 (N_12258,N_10382,N_10388);
nand U12259 (N_12259,N_11897,N_11291);
or U12260 (N_12260,N_10022,N_10927);
nand U12261 (N_12261,N_11437,N_11863);
nor U12262 (N_12262,N_11269,N_11895);
nand U12263 (N_12263,N_11049,N_10947);
and U12264 (N_12264,N_10125,N_11613);
nand U12265 (N_12265,N_10488,N_11363);
nor U12266 (N_12266,N_11698,N_11342);
nor U12267 (N_12267,N_10717,N_11208);
nor U12268 (N_12268,N_10029,N_10647);
nand U12269 (N_12269,N_11355,N_11066);
nor U12270 (N_12270,N_10953,N_11383);
and U12271 (N_12271,N_11512,N_11725);
nand U12272 (N_12272,N_10415,N_11671);
xnor U12273 (N_12273,N_10414,N_10453);
or U12274 (N_12274,N_11609,N_11378);
and U12275 (N_12275,N_10129,N_11168);
xnor U12276 (N_12276,N_11017,N_11276);
nand U12277 (N_12277,N_10181,N_11988);
and U12278 (N_12278,N_11360,N_10402);
nor U12279 (N_12279,N_10465,N_11661);
or U12280 (N_12280,N_11787,N_10106);
nor U12281 (N_12281,N_10284,N_10578);
nor U12282 (N_12282,N_10176,N_11240);
nor U12283 (N_12283,N_11566,N_11785);
and U12284 (N_12284,N_10044,N_11715);
nor U12285 (N_12285,N_10225,N_11391);
and U12286 (N_12286,N_11242,N_11179);
and U12287 (N_12287,N_10847,N_11098);
and U12288 (N_12288,N_10929,N_10875);
and U12289 (N_12289,N_11821,N_10462);
nand U12290 (N_12290,N_11599,N_10474);
or U12291 (N_12291,N_10911,N_11568);
nor U12292 (N_12292,N_11330,N_10337);
or U12293 (N_12293,N_10250,N_10640);
nor U12294 (N_12294,N_11115,N_11464);
nand U12295 (N_12295,N_11006,N_10269);
and U12296 (N_12296,N_10150,N_11205);
and U12297 (N_12297,N_11792,N_10989);
nand U12298 (N_12298,N_10113,N_11751);
nand U12299 (N_12299,N_10082,N_11776);
and U12300 (N_12300,N_10397,N_11553);
xnor U12301 (N_12301,N_11620,N_11057);
nand U12302 (N_12302,N_11369,N_10982);
nor U12303 (N_12303,N_10429,N_11885);
nand U12304 (N_12304,N_10934,N_11164);
or U12305 (N_12305,N_10297,N_10678);
or U12306 (N_12306,N_10144,N_11768);
nor U12307 (N_12307,N_11958,N_10452);
or U12308 (N_12308,N_11119,N_11156);
nor U12309 (N_12309,N_10368,N_10696);
nand U12310 (N_12310,N_11723,N_10507);
xor U12311 (N_12311,N_11581,N_10547);
xor U12312 (N_12312,N_10194,N_10973);
and U12313 (N_12313,N_10529,N_11216);
and U12314 (N_12314,N_11486,N_11749);
and U12315 (N_12315,N_10279,N_10071);
or U12316 (N_12316,N_10626,N_11700);
xnor U12317 (N_12317,N_11603,N_10047);
nor U12318 (N_12318,N_11545,N_10923);
or U12319 (N_12319,N_10612,N_11647);
and U12320 (N_12320,N_11761,N_10035);
or U12321 (N_12321,N_11560,N_10107);
nor U12322 (N_12322,N_11978,N_11483);
and U12323 (N_12323,N_10863,N_10772);
nand U12324 (N_12324,N_11686,N_11656);
nand U12325 (N_12325,N_10154,N_10063);
nand U12326 (N_12326,N_11002,N_11708);
nand U12327 (N_12327,N_10543,N_11301);
nor U12328 (N_12328,N_10984,N_11184);
nor U12329 (N_12329,N_11923,N_10096);
or U12330 (N_12330,N_11147,N_11784);
and U12331 (N_12331,N_10966,N_10996);
nor U12332 (N_12332,N_11522,N_10214);
or U12333 (N_12333,N_11727,N_10262);
nand U12334 (N_12334,N_10135,N_11136);
nand U12335 (N_12335,N_10777,N_11005);
or U12336 (N_12336,N_10589,N_11307);
or U12337 (N_12337,N_11688,N_10428);
and U12338 (N_12338,N_11684,N_11547);
or U12339 (N_12339,N_11137,N_11892);
nor U12340 (N_12340,N_10017,N_10300);
or U12341 (N_12341,N_10719,N_11672);
nand U12342 (N_12342,N_10511,N_10667);
nand U12343 (N_12343,N_10239,N_11879);
or U12344 (N_12344,N_10869,N_11477);
nand U12345 (N_12345,N_11794,N_10558);
or U12346 (N_12346,N_11633,N_10260);
and U12347 (N_12347,N_11729,N_10303);
nand U12348 (N_12348,N_10766,N_10502);
nand U12349 (N_12349,N_11530,N_11739);
or U12350 (N_12350,N_10655,N_11121);
nand U12351 (N_12351,N_10765,N_10505);
nor U12352 (N_12352,N_10512,N_10342);
nand U12353 (N_12353,N_11774,N_10685);
nand U12354 (N_12354,N_11632,N_10544);
nand U12355 (N_12355,N_11994,N_10160);
nor U12356 (N_12356,N_10835,N_11976);
nand U12357 (N_12357,N_11323,N_10901);
nand U12358 (N_12358,N_11689,N_11747);
nand U12359 (N_12359,N_11956,N_10405);
or U12360 (N_12360,N_11254,N_11937);
and U12361 (N_12361,N_11673,N_10503);
or U12362 (N_12362,N_10320,N_11580);
or U12363 (N_12363,N_11843,N_11122);
or U12364 (N_12364,N_10079,N_11040);
xor U12365 (N_12365,N_10406,N_10311);
or U12366 (N_12366,N_11303,N_10844);
or U12367 (N_12367,N_11842,N_10290);
and U12368 (N_12368,N_11612,N_11762);
and U12369 (N_12369,N_11528,N_10707);
or U12370 (N_12370,N_11570,N_10410);
nand U12371 (N_12371,N_10932,N_11222);
nor U12372 (N_12372,N_10354,N_10392);
and U12373 (N_12373,N_11125,N_10782);
nor U12374 (N_12374,N_11227,N_10114);
and U12375 (N_12375,N_11914,N_11113);
or U12376 (N_12376,N_11418,N_11193);
nand U12377 (N_12377,N_11875,N_10292);
and U12378 (N_12378,N_11237,N_10332);
xor U12379 (N_12379,N_10078,N_11150);
nor U12380 (N_12380,N_10582,N_11476);
nand U12381 (N_12381,N_10457,N_11163);
nand U12382 (N_12382,N_11143,N_10665);
xnor U12383 (N_12383,N_11718,N_11871);
and U12384 (N_12384,N_11906,N_10359);
or U12385 (N_12385,N_10532,N_11334);
xnor U12386 (N_12386,N_10705,N_10081);
nor U12387 (N_12387,N_11196,N_11905);
and U12388 (N_12388,N_10649,N_11343);
and U12389 (N_12389,N_11154,N_11224);
or U12390 (N_12390,N_10819,N_11972);
or U12391 (N_12391,N_11398,N_11406);
nor U12392 (N_12392,N_11285,N_10822);
nor U12393 (N_12393,N_11371,N_11387);
nand U12394 (N_12394,N_10383,N_10266);
or U12395 (N_12395,N_11075,N_11069);
nor U12396 (N_12396,N_10506,N_11062);
nor U12397 (N_12397,N_11252,N_10836);
nand U12398 (N_12398,N_10276,N_10509);
or U12399 (N_12399,N_10912,N_10379);
nand U12400 (N_12400,N_11261,N_11116);
nand U12401 (N_12401,N_10141,N_10149);
or U12402 (N_12402,N_11275,N_10891);
nand U12403 (N_12403,N_11932,N_10754);
xnor U12404 (N_12404,N_11524,N_11445);
xor U12405 (N_12405,N_10019,N_11202);
xnor U12406 (N_12406,N_11145,N_11960);
nand U12407 (N_12407,N_10807,N_11621);
or U12408 (N_12408,N_10683,N_10327);
and U12409 (N_12409,N_11752,N_10491);
and U12410 (N_12410,N_10328,N_11748);
and U12411 (N_12411,N_10949,N_10136);
and U12412 (N_12412,N_11717,N_10287);
nand U12413 (N_12413,N_10559,N_10094);
or U12414 (N_12414,N_10921,N_11392);
nor U12415 (N_12415,N_11681,N_10231);
nand U12416 (N_12416,N_11665,N_11755);
and U12417 (N_12417,N_10991,N_10876);
nor U12418 (N_12418,N_10085,N_11394);
and U12419 (N_12419,N_10885,N_11593);
xnor U12420 (N_12420,N_10404,N_11488);
or U12421 (N_12421,N_11554,N_10763);
or U12422 (N_12422,N_11704,N_10749);
and U12423 (N_12423,N_10843,N_11546);
or U12424 (N_12424,N_11231,N_10403);
and U12425 (N_12425,N_11506,N_11993);
nor U12426 (N_12426,N_11919,N_10792);
nand U12427 (N_12427,N_11658,N_10089);
xnor U12428 (N_12428,N_11078,N_10525);
nand U12429 (N_12429,N_10168,N_11925);
xor U12430 (N_12430,N_11908,N_10882);
nand U12431 (N_12431,N_10143,N_10254);
or U12432 (N_12432,N_10832,N_10185);
nor U12433 (N_12433,N_10999,N_11891);
xor U12434 (N_12434,N_10597,N_11438);
nand U12435 (N_12435,N_11048,N_11087);
and U12436 (N_12436,N_10753,N_11859);
or U12437 (N_12437,N_11108,N_11372);
nor U12438 (N_12438,N_10699,N_10251);
and U12439 (N_12439,N_11416,N_11132);
or U12440 (N_12440,N_11013,N_10803);
or U12441 (N_12441,N_11455,N_10192);
xnor U12442 (N_12442,N_11376,N_10769);
or U12443 (N_12443,N_11587,N_10634);
nand U12444 (N_12444,N_11135,N_10138);
nor U12445 (N_12445,N_11295,N_10463);
and U12446 (N_12446,N_10360,N_10223);
xnor U12447 (N_12447,N_11131,N_10530);
or U12448 (N_12448,N_11675,N_11454);
nor U12449 (N_12449,N_11349,N_11903);
or U12450 (N_12450,N_10839,N_10140);
and U12451 (N_12451,N_10158,N_11765);
nand U12452 (N_12452,N_10258,N_11219);
nand U12453 (N_12453,N_10706,N_10031);
and U12454 (N_12454,N_11610,N_10703);
or U12455 (N_12455,N_10211,N_10145);
nor U12456 (N_12456,N_10605,N_10310);
nand U12457 (N_12457,N_11628,N_11783);
or U12458 (N_12458,N_11888,N_10549);
nor U12459 (N_12459,N_10066,N_11571);
nor U12460 (N_12460,N_10524,N_11173);
and U12461 (N_12461,N_11614,N_11008);
nand U12462 (N_12462,N_11243,N_10348);
nand U12463 (N_12463,N_11870,N_10887);
xnor U12464 (N_12464,N_10080,N_11448);
xnor U12465 (N_12465,N_11089,N_10636);
nor U12466 (N_12466,N_11965,N_11858);
nor U12467 (N_12467,N_11878,N_10288);
and U12468 (N_12468,N_10727,N_10639);
and U12469 (N_12469,N_11782,N_11215);
nor U12470 (N_12470,N_10190,N_10570);
or U12471 (N_12471,N_10157,N_11287);
or U12472 (N_12472,N_10641,N_11421);
and U12473 (N_12473,N_10475,N_11959);
nor U12474 (N_12474,N_10243,N_10442);
and U12475 (N_12475,N_10309,N_10301);
nor U12476 (N_12476,N_11909,N_10775);
nor U12477 (N_12477,N_11099,N_11402);
or U12478 (N_12478,N_10126,N_10660);
nand U12479 (N_12479,N_11781,N_11038);
nor U12480 (N_12480,N_10378,N_10971);
xnor U12481 (N_12481,N_11456,N_10816);
or U12482 (N_12482,N_11583,N_10036);
nand U12483 (N_12483,N_10629,N_10023);
nand U12484 (N_12484,N_11509,N_11780);
or U12485 (N_12485,N_10813,N_11523);
xor U12486 (N_12486,N_10721,N_11541);
or U12487 (N_12487,N_10242,N_11904);
and U12488 (N_12488,N_11944,N_10255);
xnor U12489 (N_12489,N_11081,N_11072);
nor U12490 (N_12490,N_10162,N_11760);
nand U12491 (N_12491,N_11283,N_10476);
nor U12492 (N_12492,N_10147,N_10637);
nand U12493 (N_12493,N_10275,N_11380);
nand U12494 (N_12494,N_11426,N_10628);
and U12495 (N_12495,N_10784,N_10345);
nand U12496 (N_12496,N_10448,N_11687);
or U12497 (N_12497,N_10385,N_11746);
nand U12498 (N_12498,N_11068,N_11178);
or U12499 (N_12499,N_10550,N_10653);
nand U12500 (N_12500,N_11716,N_10643);
nor U12501 (N_12501,N_10845,N_11917);
and U12502 (N_12502,N_11414,N_11157);
nand U12503 (N_12503,N_10386,N_10357);
or U12504 (N_12504,N_11354,N_11313);
nor U12505 (N_12505,N_11759,N_11766);
xnor U12506 (N_12506,N_11432,N_11848);
or U12507 (N_12507,N_11070,N_10093);
xor U12508 (N_12508,N_10601,N_11118);
nor U12509 (N_12509,N_10122,N_10076);
or U12510 (N_12510,N_10644,N_10810);
nor U12511 (N_12511,N_10535,N_10177);
and U12512 (N_12512,N_11840,N_10892);
and U12513 (N_12513,N_10799,N_11191);
or U12514 (N_12514,N_10313,N_11239);
nand U12515 (N_12515,N_10108,N_11770);
and U12516 (N_12516,N_10729,N_10871);
nand U12517 (N_12517,N_10913,N_11839);
and U12518 (N_12518,N_10574,N_10841);
or U12519 (N_12519,N_10212,N_11957);
xor U12520 (N_12520,N_10818,N_11332);
and U12521 (N_12521,N_10068,N_10758);
and U12522 (N_12522,N_10981,N_10713);
or U12523 (N_12523,N_10006,N_11037);
or U12524 (N_12524,N_10460,N_11643);
or U12525 (N_12525,N_11829,N_11111);
nand U12526 (N_12526,N_10257,N_11736);
or U12527 (N_12527,N_11504,N_11811);
and U12528 (N_12528,N_10917,N_10235);
nand U12529 (N_12529,N_10517,N_11447);
nand U12530 (N_12530,N_11877,N_11112);
or U12531 (N_12531,N_10049,N_10441);
and U12532 (N_12532,N_10315,N_10868);
xnor U12533 (N_12533,N_10978,N_10338);
and U12534 (N_12534,N_10184,N_11816);
and U12535 (N_12535,N_11114,N_10349);
nor U12536 (N_12536,N_10412,N_10632);
or U12537 (N_12537,N_10420,N_10467);
nand U12538 (N_12538,N_11065,N_11452);
nor U12539 (N_12539,N_11427,N_11359);
xnor U12540 (N_12540,N_10764,N_10645);
and U12541 (N_12541,N_10823,N_10387);
nor U12542 (N_12542,N_10954,N_10583);
nor U12543 (N_12543,N_11003,N_10633);
and U12544 (N_12544,N_11529,N_11795);
nand U12545 (N_12545,N_10198,N_10222);
or U12546 (N_12546,N_10904,N_11505);
xor U12547 (N_12547,N_10676,N_11997);
or U12548 (N_12548,N_10124,N_11922);
or U12549 (N_12549,N_10027,N_10592);
or U12550 (N_12550,N_11831,N_11433);
and U12551 (N_12551,N_10263,N_11833);
nand U12552 (N_12552,N_10620,N_10700);
nor U12553 (N_12553,N_10445,N_10591);
nor U12554 (N_12554,N_10203,N_10358);
and U12555 (N_12555,N_11586,N_10008);
xnor U12556 (N_12556,N_11368,N_10018);
and U12557 (N_12557,N_10773,N_11813);
nand U12558 (N_12558,N_10722,N_11129);
and U12559 (N_12559,N_11194,N_11533);
xor U12560 (N_12560,N_11442,N_11084);
and U12561 (N_12561,N_10285,N_10831);
nor U12562 (N_12562,N_10439,N_10230);
nand U12563 (N_12563,N_10330,N_11232);
and U12564 (N_12564,N_11058,N_11800);
or U12565 (N_12565,N_11757,N_10489);
or U12566 (N_12566,N_11375,N_11160);
or U12567 (N_12567,N_11732,N_11278);
xnor U12568 (N_12568,N_11798,N_10673);
and U12569 (N_12569,N_11007,N_11720);
nor U12570 (N_12570,N_10866,N_10877);
nand U12571 (N_12571,N_10322,N_11102);
and U12572 (N_12572,N_11054,N_10950);
xor U12573 (N_12573,N_11187,N_10867);
nor U12574 (N_12574,N_10648,N_10312);
xnor U12575 (N_12575,N_11992,N_11955);
nor U12576 (N_12576,N_10010,N_11652);
nor U12577 (N_12577,N_10037,N_10139);
and U12578 (N_12578,N_10873,N_10374);
nor U12579 (N_12579,N_10299,N_11064);
nand U12580 (N_12580,N_10293,N_10054);
and U12581 (N_12581,N_10638,N_11662);
and U12582 (N_12582,N_11212,N_11159);
and U12583 (N_12583,N_11838,N_10725);
nor U12584 (N_12584,N_10249,N_10747);
nand U12585 (N_12585,N_10789,N_10259);
and U12586 (N_12586,N_11047,N_10607);
nor U12587 (N_12587,N_11764,N_11592);
and U12588 (N_12588,N_10356,N_11849);
or U12589 (N_12589,N_10606,N_10811);
nand U12590 (N_12590,N_11076,N_10433);
or U12591 (N_12591,N_10508,N_10252);
nand U12592 (N_12592,N_10755,N_10805);
and U12593 (N_12593,N_11206,N_10208);
or U12594 (N_12594,N_11444,N_10733);
or U12595 (N_12595,N_11385,N_10134);
nor U12596 (N_12596,N_11527,N_11837);
nand U12597 (N_12597,N_11011,N_10407);
xor U12598 (N_12598,N_10870,N_11146);
nor U12599 (N_12599,N_10711,N_11096);
or U12600 (N_12600,N_11351,N_11390);
nand U12601 (N_12601,N_10909,N_10456);
and U12602 (N_12602,N_11262,N_10105);
or U12603 (N_12603,N_10473,N_10794);
or U12604 (N_12604,N_11316,N_11590);
nor U12605 (N_12605,N_10786,N_11071);
or U12606 (N_12606,N_10128,N_10264);
nor U12607 (N_12607,N_10042,N_11001);
nor U12608 (N_12608,N_10091,N_10060);
and U12609 (N_12609,N_11820,N_11407);
xnor U12610 (N_12610,N_10746,N_11574);
or U12611 (N_12611,N_11824,N_10687);
nor U12612 (N_12612,N_10740,N_10205);
nand U12613 (N_12613,N_11256,N_11998);
nand U12614 (N_12614,N_11948,N_11357);
or U12615 (N_12615,N_11281,N_11225);
xor U12616 (N_12616,N_10069,N_11051);
or U12617 (N_12617,N_11487,N_10308);
nor U12618 (N_12618,N_11822,N_11790);
nand U12619 (N_12619,N_10155,N_11987);
and U12620 (N_12620,N_10742,N_11462);
or U12621 (N_12621,N_11101,N_10884);
and U12622 (N_12622,N_11819,N_11518);
and U12623 (N_12623,N_10806,N_11451);
nand U12624 (N_12624,N_11779,N_11738);
and U12625 (N_12625,N_10418,N_11247);
or U12626 (N_12626,N_10872,N_10067);
nand U12627 (N_12627,N_11088,N_11183);
or U12628 (N_12628,N_10970,N_10384);
nor U12629 (N_12629,N_10804,N_10111);
nand U12630 (N_12630,N_11989,N_11771);
or U12631 (N_12631,N_11198,N_10848);
nor U12632 (N_12632,N_10370,N_11763);
nor U12633 (N_12633,N_11982,N_10152);
nand U12634 (N_12634,N_10472,N_11719);
nor U12635 (N_12635,N_10120,N_10234);
or U12636 (N_12636,N_10670,N_10849);
nor U12637 (N_12637,N_10708,N_10853);
and U12638 (N_12638,N_10116,N_11186);
and U12639 (N_12639,N_10694,N_11034);
or U12640 (N_12640,N_10137,N_11284);
or U12641 (N_12641,N_10770,N_10846);
and U12642 (N_12642,N_11138,N_11336);
nor U12643 (N_12643,N_10757,N_11346);
or U12644 (N_12644,N_11500,N_10236);
and U12645 (N_12645,N_10077,N_11297);
nand U12646 (N_12646,N_11434,N_10340);
nor U12647 (N_12647,N_10926,N_10095);
and U12648 (N_12648,N_11010,N_11827);
nand U12649 (N_12649,N_11961,N_10555);
xnor U12650 (N_12650,N_11659,N_11962);
and U12651 (N_12651,N_10714,N_10894);
xnor U12652 (N_12652,N_10119,N_11130);
nand U12653 (N_12653,N_11677,N_10854);
xor U12654 (N_12654,N_11182,N_11185);
nand U12655 (N_12655,N_11172,N_10610);
nand U12656 (N_12656,N_10627,N_10083);
and U12657 (N_12657,N_10521,N_11246);
nand U12658 (N_12658,N_11880,N_10581);
nand U12659 (N_12659,N_10153,N_11618);
xnor U12660 (N_12660,N_10937,N_11229);
and U12661 (N_12661,N_11458,N_11595);
nand U12662 (N_12662,N_10056,N_10652);
and U12663 (N_12663,N_10130,N_10351);
or U12664 (N_12664,N_10098,N_10695);
or U12665 (N_12665,N_10671,N_10318);
nand U12666 (N_12666,N_10215,N_10045);
nand U12667 (N_12667,N_11777,N_11103);
and U12668 (N_12668,N_11678,N_11577);
xor U12669 (N_12669,N_10919,N_10097);
or U12670 (N_12670,N_11304,N_10737);
xor U12671 (N_12671,N_11273,N_11544);
and U12672 (N_12672,N_11310,N_10580);
xnor U12673 (N_12673,N_10980,N_11884);
and U12674 (N_12674,N_10616,N_10270);
nor U12675 (N_12675,N_11031,N_10914);
and U12676 (N_12676,N_10959,N_11712);
or U12677 (N_12677,N_11983,N_10759);
or U12678 (N_12678,N_10362,N_11012);
or U12679 (N_12679,N_10614,N_10003);
or U12680 (N_12680,N_11772,N_10195);
and U12681 (N_12681,N_10881,N_11082);
xnor U12682 (N_12682,N_10979,N_11248);
or U12683 (N_12683,N_11921,N_11556);
nand U12684 (N_12684,N_10058,N_11044);
or U12685 (N_12685,N_11305,N_11805);
nor U12686 (N_12686,N_10286,N_11692);
nand U12687 (N_12687,N_11882,N_10716);
nor U12688 (N_12688,N_11702,N_11589);
xor U12689 (N_12689,N_10572,N_11022);
or U12690 (N_12690,N_11573,N_11280);
or U12691 (N_12691,N_11539,N_10967);
and U12692 (N_12692,N_11080,N_10193);
nand U12693 (N_12693,N_11985,N_11954);
nand U12694 (N_12694,N_10046,N_10896);
or U12695 (N_12695,N_10701,N_11035);
nor U12696 (N_12696,N_10957,N_11341);
nor U12697 (N_12697,N_10486,N_10898);
nand U12698 (N_12698,N_11180,N_10879);
and U12699 (N_12699,N_10958,N_11271);
or U12700 (N_12700,N_11419,N_11649);
nor U12701 (N_12701,N_10865,N_11405);
xor U12702 (N_12702,N_11591,N_11941);
or U12703 (N_12703,N_10295,N_10074);
nand U12704 (N_12704,N_10577,N_10952);
nand U12705 (N_12705,N_11128,N_10566);
nand U12706 (N_12706,N_11602,N_10656);
nor U12707 (N_12707,N_10001,N_10110);
nor U12708 (N_12708,N_11461,N_10704);
xor U12709 (N_12709,N_10438,N_10393);
xnor U12710 (N_12710,N_10092,N_11063);
xnor U12711 (N_12711,N_10791,N_10224);
nor U12712 (N_12712,N_11210,N_11631);
and U12713 (N_12713,N_10840,N_10751);
nor U12714 (N_12714,N_11557,N_10375);
nor U12715 (N_12715,N_10520,N_10021);
nor U12716 (N_12716,N_10609,N_11350);
nor U12717 (N_12717,N_11292,N_11493);
nand U12718 (N_12718,N_10103,N_11423);
nand U12719 (N_12719,N_10940,N_11188);
or U12720 (N_12720,N_10075,N_10743);
nand U12721 (N_12721,N_11411,N_11521);
or U12722 (N_12722,N_11499,N_10248);
and U12723 (N_12723,N_11465,N_10541);
nand U12724 (N_12724,N_11358,N_11666);
and U12725 (N_12725,N_10471,N_10041);
or U12726 (N_12726,N_11862,N_11345);
or U12727 (N_12727,N_11364,N_10088);
xnor U12728 (N_12728,N_10265,N_11857);
nand U12729 (N_12729,N_10961,N_10171);
nand U12730 (N_12730,N_10209,N_10785);
or U12731 (N_12731,N_10202,N_10992);
and U12732 (N_12732,N_11537,N_11902);
or U12733 (N_12733,N_11796,N_11365);
nand U12734 (N_12734,N_10732,N_10099);
nor U12735 (N_12735,N_11742,N_10780);
nor U12736 (N_12736,N_10240,N_10852);
nand U12737 (N_12737,N_10500,N_11492);
nor U12738 (N_12738,N_10493,N_11158);
and U12739 (N_12739,N_11676,N_11241);
xnor U12740 (N_12740,N_11211,N_10796);
and U12741 (N_12741,N_11639,N_11969);
nor U12742 (N_12742,N_11793,N_11481);
and U12743 (N_12743,N_10443,N_11615);
xor U12744 (N_12744,N_10294,N_10188);
or U12745 (N_12745,N_10880,N_11272);
or U12746 (N_12746,N_10731,N_11386);
nor U12747 (N_12747,N_10890,N_11097);
and U12748 (N_12748,N_10421,N_11986);
nand U12749 (N_12749,N_11679,N_11817);
nand U12750 (N_12750,N_11370,N_11756);
nor U12751 (N_12751,N_11400,N_10477);
and U12752 (N_12752,N_10002,N_11636);
nand U12753 (N_12753,N_10663,N_10697);
nand U12754 (N_12754,N_11466,N_11485);
and U12755 (N_12755,N_11218,N_10408);
xor U12756 (N_12756,N_10026,N_11743);
nor U12757 (N_12757,N_10995,N_10878);
or U12758 (N_12758,N_11913,N_11382);
and U12759 (N_12759,N_11374,N_10376);
and U12760 (N_12760,N_11263,N_10101);
or U12761 (N_12761,N_10148,N_11420);
nand U12762 (N_12762,N_10398,N_11625);
nand U12763 (N_12763,N_10538,N_10210);
and U12764 (N_12764,N_10496,N_11974);
nand U12765 (N_12765,N_11642,N_10361);
nand U12766 (N_12766,N_11453,N_11023);
and U12767 (N_12767,N_10118,N_11497);
xnor U12768 (N_12768,N_10682,N_11745);
xor U12769 (N_12769,N_11786,N_10024);
xnor U12770 (N_12770,N_11543,N_10204);
or U12771 (N_12771,N_10373,N_11061);
nand U12772 (N_12772,N_11258,N_11733);
or U12773 (N_12773,N_10072,N_11095);
nor U12774 (N_12774,N_11446,N_11867);
nand U12775 (N_12775,N_10336,N_11942);
and U12776 (N_12776,N_11441,N_10838);
or U12777 (N_12777,N_11555,N_11868);
or U12778 (N_12778,N_11588,N_11192);
nand U12779 (N_12779,N_10540,N_11396);
nand U12780 (N_12780,N_10668,N_11203);
or U12781 (N_12781,N_11490,N_10163);
or U12782 (N_12782,N_11213,N_11302);
or U12783 (N_12783,N_11737,N_11929);
xnor U12784 (N_12784,N_10305,N_11501);
nand U12785 (N_12785,N_11327,N_11654);
and U12786 (N_12786,N_11624,N_10314);
nor U12787 (N_12787,N_11175,N_11470);
nor U12788 (N_12788,N_11630,N_10423);
or U12789 (N_12789,N_10686,N_10321);
and U12790 (N_12790,N_10347,N_10801);
xor U12791 (N_12791,N_11230,N_10542);
nor U12792 (N_12792,N_10346,N_10117);
or U12793 (N_12793,N_10329,N_11475);
nor U12794 (N_12794,N_11379,N_10631);
nand U12795 (N_12795,N_10943,N_10390);
nor U12796 (N_12796,N_10197,N_11502);
nor U12797 (N_12797,N_11924,N_11450);
or U12798 (N_12798,N_10938,N_10052);
and U12799 (N_12799,N_11799,N_11027);
and U12800 (N_12800,N_11773,N_10487);
nor U12801 (N_12801,N_10842,N_10217);
or U12802 (N_12802,N_11604,N_10132);
or U12803 (N_12803,N_10997,N_11562);
nor U12804 (N_12804,N_10993,N_11876);
or U12805 (N_12805,N_10948,N_11495);
and U12806 (N_12806,N_10723,N_10061);
and U12807 (N_12807,N_11056,N_11645);
nand U12808 (N_12808,N_10681,N_10662);
xnor U12809 (N_12809,N_10850,N_10942);
or U12810 (N_12810,N_10302,N_10787);
or U12811 (N_12811,N_11616,N_11788);
or U12812 (N_12812,N_11377,N_10657);
nand U12813 (N_12813,N_11629,N_11482);
and U12814 (N_12814,N_10051,N_10482);
nand U12815 (N_12815,N_10199,N_10736);
nand U12816 (N_12816,N_11197,N_10431);
or U12817 (N_12817,N_10449,N_11950);
nor U12818 (N_12818,N_11457,N_11657);
nand U12819 (N_12819,N_10306,N_11828);
nor U12820 (N_12820,N_10956,N_11046);
or U12821 (N_12821,N_11928,N_11809);
nand U12822 (N_12822,N_10485,N_11515);
nor U12823 (N_12823,N_11025,N_10965);
nand U12824 (N_12824,N_10131,N_10030);
nor U12825 (N_12825,N_11033,N_11410);
and U12826 (N_12826,N_11459,N_10567);
and U12827 (N_12827,N_10693,N_11140);
nor U12828 (N_12828,N_11873,N_10864);
and U12829 (N_12829,N_10372,N_10528);
nor U12830 (N_12830,N_11734,N_10834);
nor U12831 (N_12831,N_11149,N_10479);
and U12832 (N_12832,N_11165,N_11900);
nor U12833 (N_12833,N_10497,N_10990);
and U12834 (N_12834,N_11823,N_10779);
nand U12835 (N_12835,N_10201,N_11832);
xnor U12836 (N_12836,N_10709,N_11598);
nor U12837 (N_12837,N_11134,N_10401);
nor U12838 (N_12838,N_10519,N_10238);
and U12839 (N_12839,N_10173,N_11335);
nor U12840 (N_12840,N_11249,N_10028);
and U12841 (N_12841,N_10207,N_10344);
and U12842 (N_12842,N_11706,N_10307);
and U12843 (N_12843,N_10513,N_10289);
nor U12844 (N_12844,N_11996,N_11889);
and U12845 (N_12845,N_10916,N_10244);
and U12846 (N_12846,N_10245,N_11009);
nor U12847 (N_12847,N_10552,N_10621);
nor U12848 (N_12848,N_10651,N_11319);
nand U12849 (N_12849,N_11951,N_11594);
or U12850 (N_12850,N_11401,N_11883);
or U12851 (N_12851,N_11251,N_10922);
nand U12852 (N_12852,N_11916,N_11077);
nor U12853 (N_12853,N_10127,N_10715);
xor U12854 (N_12854,N_11934,N_11238);
and U12855 (N_12855,N_11939,N_11767);
and U12856 (N_12856,N_10371,N_10087);
nor U12857 (N_12857,N_11947,N_11094);
xnor U12858 (N_12858,N_10925,N_10720);
xnor U12859 (N_12859,N_11696,N_11844);
nand U12860 (N_12860,N_11161,N_10617);
or U12861 (N_12861,N_11052,N_10931);
nand U12862 (N_12862,N_11968,N_10282);
xnor U12863 (N_12863,N_11397,N_10123);
nand U12864 (N_12864,N_11059,N_10335);
nor U12865 (N_12865,N_10178,N_10364);
nor U12866 (N_12866,N_10164,N_10902);
nor U12867 (N_12867,N_11279,N_11946);
nand U12868 (N_12868,N_10825,N_10658);
nand U12869 (N_12869,N_10675,N_11177);
nand U12870 (N_12870,N_10011,N_10897);
and U12871 (N_12871,N_11815,N_11683);
nand U12872 (N_12872,N_11250,N_11030);
or U12873 (N_12873,N_10353,N_11498);
nor U12874 (N_12874,N_10363,N_10038);
or U12875 (N_12875,N_10000,N_10256);
nor U12876 (N_12876,N_11721,N_11503);
nand U12877 (N_12877,N_10963,N_11830);
and U12878 (N_12878,N_11104,N_11938);
nor U12879 (N_12879,N_10220,N_10905);
or U12880 (N_12880,N_11494,N_10588);
nor U12881 (N_12881,N_10830,N_10516);
nor U12882 (N_12882,N_10334,N_11789);
or U12883 (N_12883,N_10090,N_11540);
and U12884 (N_12884,N_11804,N_10536);
or U12885 (N_12885,N_10960,N_10213);
xor U12886 (N_12886,N_11981,N_11561);
or U12887 (N_12887,N_11195,N_11484);
or U12888 (N_12888,N_10598,N_11148);
and U12889 (N_12889,N_11511,N_10416);
nor U12890 (N_12890,N_11912,N_10859);
nand U12891 (N_12891,N_10768,N_11460);
or U12892 (N_12892,N_11582,N_10724);
nand U12893 (N_12893,N_11473,N_10424);
or U12894 (N_12894,N_11576,N_11648);
nor U12895 (N_12895,N_11918,N_10200);
and U12896 (N_12896,N_11123,N_11812);
or U12897 (N_12897,N_10710,N_10454);
and U12898 (N_12898,N_11264,N_10159);
and U12899 (N_12899,N_10798,N_11584);
or U12900 (N_12900,N_10820,N_10698);
and U12901 (N_12901,N_11814,N_10323);
and U12902 (N_12902,N_10935,N_11036);
and U12903 (N_12903,N_10112,N_11907);
nand U12904 (N_12904,N_11474,N_11920);
and U12905 (N_12905,N_11155,N_11020);
and U12906 (N_12906,N_11338,N_11201);
nor U12907 (N_12907,N_10515,N_11608);
nor U12908 (N_12908,N_11181,N_10146);
and U12909 (N_12909,N_10196,N_11435);
nand U12910 (N_12910,N_11325,N_10228);
or U12911 (N_12911,N_11535,N_11674);
nand U12912 (N_12912,N_11265,N_11510);
nor U12913 (N_12913,N_10422,N_10324);
or U12914 (N_12914,N_11945,N_10020);
nor U12915 (N_12915,N_10561,N_11436);
xor U12916 (N_12916,N_11393,N_10186);
or U12917 (N_12917,N_11326,N_11311);
or U12918 (N_12918,N_10594,N_10053);
and U12919 (N_12919,N_11769,N_10575);
and U12920 (N_12920,N_10458,N_10389);
xor U12921 (N_12921,N_11641,N_10034);
nor U12922 (N_12922,N_11640,N_11846);
and U12923 (N_12923,N_11308,N_10339);
nand U12924 (N_12924,N_11353,N_11825);
and U12925 (N_12925,N_10537,N_11558);
xor U12926 (N_12926,N_10680,N_11853);
nand U12927 (N_12927,N_10059,N_10216);
nor U12928 (N_12928,N_11682,N_10800);
or U12929 (N_12929,N_11015,N_11233);
nor U12930 (N_12930,N_10930,N_11042);
nand U12931 (N_12931,N_10596,N_11449);
xnor U12932 (N_12932,N_11911,N_10450);
nor U12933 (N_12933,N_10955,N_11714);
nor U12934 (N_12934,N_11004,N_11693);
or U12935 (N_12935,N_10630,N_10174);
nand U12936 (N_12936,N_11634,N_10446);
nor U12937 (N_12937,N_11403,N_10802);
nor U12938 (N_12938,N_10464,N_10837);
nor U12939 (N_12939,N_11090,N_11967);
nand U12940 (N_12940,N_10253,N_10986);
nor U12941 (N_12941,N_10531,N_11422);
or U12942 (N_12942,N_10492,N_11542);
and U12943 (N_12943,N_10004,N_10738);
nand U12944 (N_12944,N_10169,N_10043);
xor U12945 (N_12945,N_11324,N_11915);
or U12946 (N_12946,N_10039,N_11926);
xnor U12947 (N_12947,N_11596,N_11531);
nand U12948 (N_12948,N_10440,N_11854);
or U12949 (N_12949,N_11220,N_10855);
xor U12950 (N_12950,N_10394,N_10084);
xnor U12951 (N_12951,N_11709,N_11852);
xnor U12952 (N_12952,N_11730,N_10325);
or U12953 (N_12953,N_11141,N_11294);
nand U12954 (N_12954,N_10593,N_10247);
nand U12955 (N_12955,N_11894,N_11731);
nor U12956 (N_12956,N_10179,N_10571);
and U12957 (N_12957,N_11174,N_11039);
or U12958 (N_12958,N_11045,N_10744);
nand U12959 (N_12959,N_11127,N_10005);
or U12960 (N_12960,N_10319,N_11086);
or U12961 (N_12961,N_10664,N_11896);
or U12962 (N_12962,N_10659,N_11223);
nor U12963 (N_12963,N_10033,N_11236);
nand U12964 (N_12964,N_10523,N_11413);
nand U12965 (N_12965,N_11930,N_10206);
nor U12966 (N_12966,N_11899,N_11384);
xnor U12967 (N_12967,N_10057,N_10291);
and U12968 (N_12968,N_11443,N_11496);
nor U12969 (N_12969,N_10267,N_10156);
and U12970 (N_12970,N_11935,N_10167);
and U12971 (N_12971,N_11340,N_11171);
or U12972 (N_12972,N_11126,N_10776);
and U12973 (N_12973,N_11669,N_11366);
and U12974 (N_12974,N_10304,N_10296);
xnor U12975 (N_12975,N_10783,N_10341);
xnor U12976 (N_12976,N_10910,N_10459);
xnor U12977 (N_12977,N_10012,N_11597);
and U12978 (N_12978,N_11274,N_11314);
or U12979 (N_12979,N_10814,N_10951);
or U12980 (N_12980,N_11650,N_11953);
and U12981 (N_12981,N_11869,N_11373);
nand U12982 (N_12982,N_11333,N_11298);
nor U12983 (N_12983,N_11021,N_10400);
nand U12984 (N_12984,N_10425,N_11826);
or U12985 (N_12985,N_10273,N_10809);
or U12986 (N_12986,N_10218,N_10261);
and U12987 (N_12987,N_10883,N_10579);
or U12988 (N_12988,N_10180,N_11286);
and U12989 (N_12989,N_11532,N_10918);
xor U12990 (N_12990,N_10381,N_10924);
or U12991 (N_12991,N_11623,N_10586);
nand U12992 (N_12992,N_11151,N_11724);
or U12993 (N_12993,N_11306,N_10546);
nand U12994 (N_12994,N_11060,N_11520);
nand U12995 (N_12995,N_10689,N_10490);
nand U12996 (N_12996,N_11204,N_11699);
nor U12997 (N_12997,N_10590,N_10469);
nand U12998 (N_12998,N_11142,N_10298);
nor U12999 (N_12999,N_11551,N_11653);
and U13000 (N_13000,N_10472,N_11250);
xnor U13001 (N_13001,N_10798,N_10713);
nand U13002 (N_13002,N_11714,N_11843);
nand U13003 (N_13003,N_10893,N_11896);
nor U13004 (N_13004,N_11872,N_10140);
and U13005 (N_13005,N_10066,N_10077);
nor U13006 (N_13006,N_10515,N_11452);
and U13007 (N_13007,N_11527,N_10769);
or U13008 (N_13008,N_10857,N_10208);
nand U13009 (N_13009,N_11199,N_11389);
nor U13010 (N_13010,N_11602,N_10447);
nor U13011 (N_13011,N_11449,N_11439);
and U13012 (N_13012,N_10931,N_11322);
xor U13013 (N_13013,N_11773,N_10803);
or U13014 (N_13014,N_11679,N_10583);
or U13015 (N_13015,N_10925,N_10082);
nor U13016 (N_13016,N_11182,N_10429);
nor U13017 (N_13017,N_10888,N_10195);
nand U13018 (N_13018,N_10831,N_10768);
or U13019 (N_13019,N_10928,N_11485);
nand U13020 (N_13020,N_11154,N_10209);
nor U13021 (N_13021,N_11813,N_10733);
nand U13022 (N_13022,N_11940,N_10493);
nand U13023 (N_13023,N_11694,N_11680);
nor U13024 (N_13024,N_10671,N_10334);
or U13025 (N_13025,N_11032,N_10413);
or U13026 (N_13026,N_11388,N_10140);
nor U13027 (N_13027,N_10187,N_10485);
and U13028 (N_13028,N_11717,N_11204);
and U13029 (N_13029,N_10602,N_11292);
nand U13030 (N_13030,N_10380,N_10660);
or U13031 (N_13031,N_10770,N_10902);
nand U13032 (N_13032,N_11979,N_10186);
or U13033 (N_13033,N_10069,N_10270);
nor U13034 (N_13034,N_10769,N_10065);
and U13035 (N_13035,N_10390,N_10437);
nand U13036 (N_13036,N_11874,N_11539);
nand U13037 (N_13037,N_11198,N_11648);
and U13038 (N_13038,N_10471,N_10231);
nor U13039 (N_13039,N_11653,N_10088);
xor U13040 (N_13040,N_11379,N_10248);
or U13041 (N_13041,N_11213,N_10663);
nor U13042 (N_13042,N_11928,N_11818);
or U13043 (N_13043,N_10824,N_11622);
and U13044 (N_13044,N_11406,N_10890);
nor U13045 (N_13045,N_10752,N_11124);
nor U13046 (N_13046,N_10126,N_11836);
nor U13047 (N_13047,N_11701,N_10234);
or U13048 (N_13048,N_10525,N_11350);
nor U13049 (N_13049,N_11324,N_11463);
and U13050 (N_13050,N_10572,N_11410);
nor U13051 (N_13051,N_11692,N_11520);
xor U13052 (N_13052,N_11983,N_10788);
and U13053 (N_13053,N_11566,N_10039);
and U13054 (N_13054,N_10556,N_11581);
nand U13055 (N_13055,N_10434,N_11654);
or U13056 (N_13056,N_10503,N_11445);
nand U13057 (N_13057,N_11614,N_11753);
xor U13058 (N_13058,N_10101,N_11215);
xnor U13059 (N_13059,N_11319,N_10347);
or U13060 (N_13060,N_11232,N_11893);
nand U13061 (N_13061,N_10265,N_11391);
or U13062 (N_13062,N_11105,N_11610);
nand U13063 (N_13063,N_10953,N_11429);
and U13064 (N_13064,N_11034,N_10375);
nor U13065 (N_13065,N_11374,N_11618);
nor U13066 (N_13066,N_11313,N_11755);
nor U13067 (N_13067,N_11929,N_11323);
or U13068 (N_13068,N_10743,N_10232);
and U13069 (N_13069,N_11837,N_10975);
nor U13070 (N_13070,N_11550,N_10390);
nor U13071 (N_13071,N_10833,N_10507);
and U13072 (N_13072,N_10104,N_10800);
nand U13073 (N_13073,N_11853,N_11755);
xor U13074 (N_13074,N_10494,N_10082);
or U13075 (N_13075,N_10525,N_11390);
or U13076 (N_13076,N_10191,N_11061);
nor U13077 (N_13077,N_11844,N_11442);
nor U13078 (N_13078,N_10091,N_10691);
or U13079 (N_13079,N_11590,N_10545);
and U13080 (N_13080,N_10310,N_10795);
or U13081 (N_13081,N_10250,N_11828);
xor U13082 (N_13082,N_11232,N_10954);
nand U13083 (N_13083,N_10079,N_11280);
xor U13084 (N_13084,N_10682,N_11405);
or U13085 (N_13085,N_10203,N_11850);
or U13086 (N_13086,N_11950,N_11562);
nand U13087 (N_13087,N_11968,N_10441);
and U13088 (N_13088,N_10720,N_11869);
nor U13089 (N_13089,N_10382,N_11328);
nand U13090 (N_13090,N_10815,N_11714);
nor U13091 (N_13091,N_11369,N_11252);
nand U13092 (N_13092,N_10766,N_11395);
nand U13093 (N_13093,N_11758,N_10656);
nand U13094 (N_13094,N_10555,N_11786);
nor U13095 (N_13095,N_10479,N_10610);
or U13096 (N_13096,N_10912,N_11331);
nand U13097 (N_13097,N_11141,N_11642);
or U13098 (N_13098,N_10285,N_11190);
nor U13099 (N_13099,N_10519,N_11388);
and U13100 (N_13100,N_11750,N_11586);
nor U13101 (N_13101,N_10044,N_11398);
xnor U13102 (N_13102,N_10427,N_10438);
xor U13103 (N_13103,N_10313,N_10559);
xor U13104 (N_13104,N_10737,N_10309);
nand U13105 (N_13105,N_10240,N_10811);
or U13106 (N_13106,N_10331,N_10422);
nand U13107 (N_13107,N_10777,N_10370);
and U13108 (N_13108,N_10451,N_11723);
xor U13109 (N_13109,N_10363,N_11836);
or U13110 (N_13110,N_10198,N_11407);
nor U13111 (N_13111,N_11517,N_11594);
nand U13112 (N_13112,N_10631,N_10504);
xor U13113 (N_13113,N_11012,N_10725);
and U13114 (N_13114,N_10639,N_11940);
or U13115 (N_13115,N_11899,N_11618);
nand U13116 (N_13116,N_11667,N_11487);
and U13117 (N_13117,N_10239,N_10773);
nor U13118 (N_13118,N_11412,N_11077);
and U13119 (N_13119,N_10204,N_11586);
or U13120 (N_13120,N_10780,N_11734);
xor U13121 (N_13121,N_11167,N_11090);
or U13122 (N_13122,N_10387,N_11919);
and U13123 (N_13123,N_11921,N_11226);
nor U13124 (N_13124,N_10068,N_10802);
xor U13125 (N_13125,N_10595,N_11796);
and U13126 (N_13126,N_11986,N_10569);
and U13127 (N_13127,N_10800,N_11302);
and U13128 (N_13128,N_10134,N_11519);
nand U13129 (N_13129,N_10233,N_11256);
or U13130 (N_13130,N_11515,N_10344);
nor U13131 (N_13131,N_11611,N_11417);
and U13132 (N_13132,N_10713,N_10642);
or U13133 (N_13133,N_10645,N_11943);
nor U13134 (N_13134,N_11874,N_11300);
nor U13135 (N_13135,N_10001,N_11884);
or U13136 (N_13136,N_10830,N_11884);
nand U13137 (N_13137,N_10024,N_11260);
nand U13138 (N_13138,N_11987,N_11079);
nor U13139 (N_13139,N_11444,N_11247);
nor U13140 (N_13140,N_11073,N_11203);
nor U13141 (N_13141,N_11983,N_11367);
or U13142 (N_13142,N_11069,N_10677);
and U13143 (N_13143,N_10670,N_10477);
and U13144 (N_13144,N_11023,N_11297);
nand U13145 (N_13145,N_11861,N_10239);
and U13146 (N_13146,N_10798,N_11381);
or U13147 (N_13147,N_11311,N_10737);
nand U13148 (N_13148,N_11385,N_11737);
or U13149 (N_13149,N_11898,N_10599);
and U13150 (N_13150,N_11980,N_11364);
and U13151 (N_13151,N_10250,N_10203);
nand U13152 (N_13152,N_11852,N_11733);
nor U13153 (N_13153,N_10139,N_10726);
xor U13154 (N_13154,N_11239,N_10536);
and U13155 (N_13155,N_10050,N_11572);
and U13156 (N_13156,N_11169,N_11007);
or U13157 (N_13157,N_11687,N_11495);
nand U13158 (N_13158,N_11623,N_10416);
xor U13159 (N_13159,N_11302,N_11934);
nor U13160 (N_13160,N_10790,N_10414);
and U13161 (N_13161,N_11941,N_11449);
and U13162 (N_13162,N_10383,N_10695);
and U13163 (N_13163,N_10968,N_11178);
nor U13164 (N_13164,N_11039,N_10747);
nand U13165 (N_13165,N_10675,N_10409);
or U13166 (N_13166,N_10974,N_10930);
nand U13167 (N_13167,N_10491,N_10548);
nor U13168 (N_13168,N_10068,N_10933);
or U13169 (N_13169,N_11180,N_10387);
and U13170 (N_13170,N_10331,N_11564);
or U13171 (N_13171,N_11995,N_11411);
and U13172 (N_13172,N_10624,N_11046);
and U13173 (N_13173,N_11189,N_10796);
or U13174 (N_13174,N_11921,N_10673);
and U13175 (N_13175,N_11089,N_11295);
and U13176 (N_13176,N_10761,N_10747);
nor U13177 (N_13177,N_11997,N_10135);
nor U13178 (N_13178,N_11267,N_10700);
and U13179 (N_13179,N_11438,N_11874);
and U13180 (N_13180,N_11746,N_10963);
nand U13181 (N_13181,N_11095,N_11212);
nor U13182 (N_13182,N_11813,N_11171);
or U13183 (N_13183,N_11255,N_11523);
xor U13184 (N_13184,N_10669,N_11769);
and U13185 (N_13185,N_10808,N_11560);
or U13186 (N_13186,N_11558,N_10676);
nand U13187 (N_13187,N_11932,N_10203);
nand U13188 (N_13188,N_11140,N_10958);
nand U13189 (N_13189,N_11054,N_11992);
and U13190 (N_13190,N_11223,N_10242);
and U13191 (N_13191,N_11067,N_10137);
and U13192 (N_13192,N_11237,N_10887);
or U13193 (N_13193,N_10673,N_11059);
nand U13194 (N_13194,N_11593,N_10093);
xnor U13195 (N_13195,N_10013,N_10116);
nand U13196 (N_13196,N_10816,N_10514);
nand U13197 (N_13197,N_10501,N_10372);
nand U13198 (N_13198,N_11145,N_10796);
nand U13199 (N_13199,N_10751,N_10813);
or U13200 (N_13200,N_11173,N_11260);
and U13201 (N_13201,N_10861,N_10404);
nand U13202 (N_13202,N_11853,N_11800);
nor U13203 (N_13203,N_11040,N_10690);
and U13204 (N_13204,N_11396,N_11225);
and U13205 (N_13205,N_10615,N_10203);
nor U13206 (N_13206,N_11122,N_11918);
nand U13207 (N_13207,N_10840,N_10453);
and U13208 (N_13208,N_10210,N_11980);
nor U13209 (N_13209,N_11283,N_11713);
nand U13210 (N_13210,N_10107,N_10463);
nor U13211 (N_13211,N_11690,N_11972);
and U13212 (N_13212,N_11434,N_11954);
or U13213 (N_13213,N_11783,N_11100);
xor U13214 (N_13214,N_11913,N_11508);
nor U13215 (N_13215,N_10475,N_11585);
nand U13216 (N_13216,N_10167,N_10245);
nand U13217 (N_13217,N_11111,N_10565);
and U13218 (N_13218,N_10261,N_10071);
nand U13219 (N_13219,N_11566,N_11465);
nand U13220 (N_13220,N_11422,N_11156);
nor U13221 (N_13221,N_11101,N_10417);
and U13222 (N_13222,N_10819,N_11438);
nand U13223 (N_13223,N_10391,N_11832);
and U13224 (N_13224,N_11972,N_10160);
and U13225 (N_13225,N_10705,N_11831);
and U13226 (N_13226,N_10081,N_10029);
xnor U13227 (N_13227,N_10930,N_10564);
nor U13228 (N_13228,N_11150,N_11664);
nand U13229 (N_13229,N_11122,N_10890);
nor U13230 (N_13230,N_11730,N_11112);
nor U13231 (N_13231,N_11700,N_11925);
and U13232 (N_13232,N_11695,N_11773);
nor U13233 (N_13233,N_10581,N_11225);
and U13234 (N_13234,N_11620,N_10580);
nor U13235 (N_13235,N_11543,N_11289);
nand U13236 (N_13236,N_10340,N_10901);
or U13237 (N_13237,N_10461,N_11390);
nand U13238 (N_13238,N_10679,N_10412);
nor U13239 (N_13239,N_11593,N_10071);
and U13240 (N_13240,N_11969,N_11551);
nor U13241 (N_13241,N_11862,N_10024);
nand U13242 (N_13242,N_10601,N_10974);
nor U13243 (N_13243,N_10092,N_10455);
or U13244 (N_13244,N_10172,N_11090);
and U13245 (N_13245,N_10988,N_11925);
nand U13246 (N_13246,N_10117,N_10981);
xnor U13247 (N_13247,N_10755,N_10409);
and U13248 (N_13248,N_10855,N_10769);
or U13249 (N_13249,N_11019,N_10461);
and U13250 (N_13250,N_11058,N_10294);
or U13251 (N_13251,N_10877,N_10381);
and U13252 (N_13252,N_10334,N_10500);
nor U13253 (N_13253,N_11087,N_11377);
or U13254 (N_13254,N_11185,N_10631);
nor U13255 (N_13255,N_10203,N_11579);
and U13256 (N_13256,N_11742,N_11248);
nand U13257 (N_13257,N_11116,N_11139);
nor U13258 (N_13258,N_10389,N_11363);
nor U13259 (N_13259,N_11499,N_10163);
or U13260 (N_13260,N_11802,N_10977);
or U13261 (N_13261,N_11358,N_11043);
or U13262 (N_13262,N_11430,N_10870);
or U13263 (N_13263,N_10285,N_10115);
nand U13264 (N_13264,N_10126,N_11420);
or U13265 (N_13265,N_10243,N_11118);
xor U13266 (N_13266,N_11926,N_10944);
nand U13267 (N_13267,N_11485,N_10297);
nand U13268 (N_13268,N_11873,N_11071);
nand U13269 (N_13269,N_10084,N_11328);
or U13270 (N_13270,N_11358,N_11036);
and U13271 (N_13271,N_11072,N_10932);
or U13272 (N_13272,N_10240,N_11220);
and U13273 (N_13273,N_11471,N_10320);
nand U13274 (N_13274,N_11135,N_10116);
nor U13275 (N_13275,N_10562,N_10931);
nor U13276 (N_13276,N_10904,N_10726);
or U13277 (N_13277,N_10064,N_11597);
nor U13278 (N_13278,N_11468,N_10843);
nor U13279 (N_13279,N_11065,N_11975);
nand U13280 (N_13280,N_11008,N_10549);
xor U13281 (N_13281,N_11655,N_11448);
and U13282 (N_13282,N_10364,N_10031);
nor U13283 (N_13283,N_10708,N_10000);
and U13284 (N_13284,N_11119,N_11797);
nand U13285 (N_13285,N_10845,N_11965);
nor U13286 (N_13286,N_10242,N_10693);
nand U13287 (N_13287,N_10107,N_10148);
and U13288 (N_13288,N_11765,N_11147);
and U13289 (N_13289,N_10752,N_11566);
nor U13290 (N_13290,N_11310,N_11498);
or U13291 (N_13291,N_10311,N_10260);
or U13292 (N_13292,N_11388,N_10525);
and U13293 (N_13293,N_10170,N_10195);
or U13294 (N_13294,N_11557,N_11858);
and U13295 (N_13295,N_10558,N_10959);
nor U13296 (N_13296,N_10744,N_11723);
nor U13297 (N_13297,N_10683,N_10360);
nor U13298 (N_13298,N_10908,N_11031);
nand U13299 (N_13299,N_11929,N_11296);
nor U13300 (N_13300,N_10633,N_10282);
nand U13301 (N_13301,N_11096,N_10346);
nand U13302 (N_13302,N_11148,N_10996);
and U13303 (N_13303,N_11970,N_10029);
and U13304 (N_13304,N_11029,N_10016);
nand U13305 (N_13305,N_10598,N_10642);
nand U13306 (N_13306,N_10914,N_10003);
or U13307 (N_13307,N_10109,N_11434);
nor U13308 (N_13308,N_10326,N_10960);
nor U13309 (N_13309,N_10558,N_10620);
or U13310 (N_13310,N_11493,N_10641);
nor U13311 (N_13311,N_10157,N_10221);
and U13312 (N_13312,N_10190,N_11331);
nand U13313 (N_13313,N_10947,N_11772);
xnor U13314 (N_13314,N_11854,N_10208);
xor U13315 (N_13315,N_11633,N_10661);
or U13316 (N_13316,N_10434,N_10127);
and U13317 (N_13317,N_10056,N_10277);
xor U13318 (N_13318,N_10233,N_10406);
or U13319 (N_13319,N_11609,N_10841);
and U13320 (N_13320,N_10834,N_10520);
or U13321 (N_13321,N_10066,N_10382);
or U13322 (N_13322,N_10287,N_10309);
and U13323 (N_13323,N_11527,N_10676);
nand U13324 (N_13324,N_11784,N_11555);
xnor U13325 (N_13325,N_11661,N_10531);
or U13326 (N_13326,N_11609,N_11784);
and U13327 (N_13327,N_10613,N_10473);
and U13328 (N_13328,N_11255,N_10671);
and U13329 (N_13329,N_10015,N_10267);
nor U13330 (N_13330,N_11944,N_11862);
xor U13331 (N_13331,N_11868,N_11593);
nand U13332 (N_13332,N_10360,N_10052);
nor U13333 (N_13333,N_10417,N_10425);
and U13334 (N_13334,N_11075,N_11224);
and U13335 (N_13335,N_10493,N_10579);
nor U13336 (N_13336,N_10362,N_11489);
or U13337 (N_13337,N_11035,N_10014);
or U13338 (N_13338,N_11017,N_10416);
nand U13339 (N_13339,N_11591,N_10928);
and U13340 (N_13340,N_11477,N_10239);
nor U13341 (N_13341,N_10719,N_10844);
nand U13342 (N_13342,N_10280,N_11178);
xnor U13343 (N_13343,N_11023,N_10480);
or U13344 (N_13344,N_10032,N_10509);
nor U13345 (N_13345,N_11663,N_11124);
xor U13346 (N_13346,N_10366,N_11789);
and U13347 (N_13347,N_10059,N_11579);
nand U13348 (N_13348,N_10580,N_10467);
or U13349 (N_13349,N_10358,N_10524);
and U13350 (N_13350,N_11945,N_10405);
and U13351 (N_13351,N_10187,N_10293);
nor U13352 (N_13352,N_11904,N_11226);
nand U13353 (N_13353,N_11327,N_11913);
xor U13354 (N_13354,N_10414,N_10658);
or U13355 (N_13355,N_10255,N_11204);
xor U13356 (N_13356,N_10051,N_10908);
and U13357 (N_13357,N_11418,N_11979);
nand U13358 (N_13358,N_10593,N_11152);
and U13359 (N_13359,N_11753,N_11351);
and U13360 (N_13360,N_10291,N_10093);
nor U13361 (N_13361,N_11742,N_11284);
nor U13362 (N_13362,N_11842,N_10228);
and U13363 (N_13363,N_10991,N_11473);
nand U13364 (N_13364,N_11347,N_10603);
and U13365 (N_13365,N_10684,N_11381);
and U13366 (N_13366,N_11691,N_10088);
or U13367 (N_13367,N_10272,N_10681);
nand U13368 (N_13368,N_11612,N_11881);
or U13369 (N_13369,N_10257,N_10323);
or U13370 (N_13370,N_10966,N_11955);
xor U13371 (N_13371,N_10422,N_10047);
or U13372 (N_13372,N_11018,N_10796);
and U13373 (N_13373,N_10513,N_10611);
or U13374 (N_13374,N_10408,N_10430);
nand U13375 (N_13375,N_10488,N_11642);
nor U13376 (N_13376,N_11863,N_11352);
nand U13377 (N_13377,N_11487,N_11126);
and U13378 (N_13378,N_10376,N_10214);
nand U13379 (N_13379,N_10475,N_10516);
nand U13380 (N_13380,N_10375,N_10708);
nor U13381 (N_13381,N_10572,N_11594);
nor U13382 (N_13382,N_10437,N_10116);
and U13383 (N_13383,N_11744,N_10937);
nand U13384 (N_13384,N_10145,N_10120);
and U13385 (N_13385,N_10832,N_11428);
nor U13386 (N_13386,N_11611,N_11682);
nand U13387 (N_13387,N_11043,N_10628);
nor U13388 (N_13388,N_11359,N_11445);
nor U13389 (N_13389,N_11760,N_11681);
nor U13390 (N_13390,N_10077,N_10906);
nor U13391 (N_13391,N_10031,N_11586);
nand U13392 (N_13392,N_10896,N_10939);
or U13393 (N_13393,N_11012,N_11555);
or U13394 (N_13394,N_10597,N_11437);
xnor U13395 (N_13395,N_11293,N_11688);
nor U13396 (N_13396,N_11485,N_10899);
nor U13397 (N_13397,N_11043,N_11151);
nor U13398 (N_13398,N_11554,N_11094);
or U13399 (N_13399,N_10223,N_11724);
and U13400 (N_13400,N_10822,N_11789);
and U13401 (N_13401,N_11936,N_11930);
nand U13402 (N_13402,N_11679,N_11695);
nor U13403 (N_13403,N_11836,N_11372);
and U13404 (N_13404,N_11700,N_11051);
and U13405 (N_13405,N_10004,N_10979);
or U13406 (N_13406,N_11887,N_11815);
nand U13407 (N_13407,N_11825,N_10202);
and U13408 (N_13408,N_10704,N_10542);
nor U13409 (N_13409,N_11845,N_10747);
nor U13410 (N_13410,N_10847,N_10390);
xor U13411 (N_13411,N_11258,N_10543);
nor U13412 (N_13412,N_10883,N_10180);
and U13413 (N_13413,N_11726,N_11572);
nor U13414 (N_13414,N_10762,N_10232);
or U13415 (N_13415,N_11972,N_11473);
or U13416 (N_13416,N_10681,N_11439);
or U13417 (N_13417,N_10783,N_10635);
nand U13418 (N_13418,N_10499,N_11957);
nand U13419 (N_13419,N_10660,N_10407);
nand U13420 (N_13420,N_11408,N_11683);
nor U13421 (N_13421,N_10394,N_10095);
nor U13422 (N_13422,N_11404,N_11427);
nand U13423 (N_13423,N_11305,N_10277);
nand U13424 (N_13424,N_11729,N_11305);
or U13425 (N_13425,N_11876,N_11054);
nor U13426 (N_13426,N_10926,N_10049);
and U13427 (N_13427,N_10222,N_11462);
nand U13428 (N_13428,N_11927,N_10983);
nor U13429 (N_13429,N_10746,N_10343);
nand U13430 (N_13430,N_10066,N_10509);
or U13431 (N_13431,N_11575,N_10487);
xnor U13432 (N_13432,N_10024,N_11151);
or U13433 (N_13433,N_11523,N_11525);
nand U13434 (N_13434,N_11994,N_10991);
nor U13435 (N_13435,N_10202,N_11597);
and U13436 (N_13436,N_10236,N_10582);
nor U13437 (N_13437,N_10537,N_10807);
nand U13438 (N_13438,N_11652,N_10791);
nor U13439 (N_13439,N_11042,N_11423);
or U13440 (N_13440,N_11695,N_11815);
or U13441 (N_13441,N_10391,N_10617);
nand U13442 (N_13442,N_11536,N_10330);
nand U13443 (N_13443,N_11241,N_10758);
nor U13444 (N_13444,N_10656,N_10017);
and U13445 (N_13445,N_11708,N_11543);
nor U13446 (N_13446,N_11059,N_11139);
xor U13447 (N_13447,N_11400,N_10717);
nand U13448 (N_13448,N_10081,N_11192);
nor U13449 (N_13449,N_11278,N_11481);
nand U13450 (N_13450,N_11912,N_11823);
nor U13451 (N_13451,N_11397,N_11541);
nor U13452 (N_13452,N_10868,N_11650);
and U13453 (N_13453,N_11330,N_11155);
xor U13454 (N_13454,N_11270,N_11624);
and U13455 (N_13455,N_10419,N_11482);
and U13456 (N_13456,N_11422,N_11103);
or U13457 (N_13457,N_11787,N_10560);
or U13458 (N_13458,N_10705,N_10442);
or U13459 (N_13459,N_11922,N_10538);
and U13460 (N_13460,N_10870,N_11603);
nor U13461 (N_13461,N_10376,N_11755);
nor U13462 (N_13462,N_10206,N_11430);
nor U13463 (N_13463,N_11352,N_10054);
and U13464 (N_13464,N_10887,N_10340);
xnor U13465 (N_13465,N_11300,N_11352);
nor U13466 (N_13466,N_11397,N_10555);
nor U13467 (N_13467,N_10928,N_11049);
nand U13468 (N_13468,N_10175,N_10452);
and U13469 (N_13469,N_10829,N_11931);
and U13470 (N_13470,N_11588,N_10892);
or U13471 (N_13471,N_10091,N_10686);
or U13472 (N_13472,N_10766,N_10638);
or U13473 (N_13473,N_10101,N_10650);
nand U13474 (N_13474,N_10101,N_11025);
and U13475 (N_13475,N_10297,N_10498);
nor U13476 (N_13476,N_10036,N_11743);
or U13477 (N_13477,N_11248,N_10448);
nor U13478 (N_13478,N_11991,N_10976);
and U13479 (N_13479,N_10237,N_10801);
xnor U13480 (N_13480,N_10823,N_11610);
xnor U13481 (N_13481,N_10734,N_11282);
and U13482 (N_13482,N_11405,N_10387);
and U13483 (N_13483,N_11253,N_11709);
and U13484 (N_13484,N_11633,N_10591);
nand U13485 (N_13485,N_11640,N_11008);
nand U13486 (N_13486,N_11484,N_10459);
xnor U13487 (N_13487,N_10597,N_10761);
nor U13488 (N_13488,N_10297,N_11963);
or U13489 (N_13489,N_11812,N_10020);
or U13490 (N_13490,N_11422,N_11235);
nor U13491 (N_13491,N_11376,N_10393);
nor U13492 (N_13492,N_11995,N_10371);
nand U13493 (N_13493,N_10664,N_11202);
or U13494 (N_13494,N_10609,N_11786);
xor U13495 (N_13495,N_11453,N_10663);
or U13496 (N_13496,N_10120,N_10588);
and U13497 (N_13497,N_10276,N_11611);
or U13498 (N_13498,N_11325,N_10559);
nor U13499 (N_13499,N_11653,N_10994);
nor U13500 (N_13500,N_10316,N_11187);
or U13501 (N_13501,N_10358,N_11074);
nor U13502 (N_13502,N_11836,N_11072);
and U13503 (N_13503,N_10481,N_10171);
nor U13504 (N_13504,N_10489,N_10699);
nand U13505 (N_13505,N_10159,N_10146);
nand U13506 (N_13506,N_11390,N_10711);
nor U13507 (N_13507,N_11812,N_11705);
and U13508 (N_13508,N_11757,N_11831);
nand U13509 (N_13509,N_10388,N_10299);
nand U13510 (N_13510,N_10656,N_11609);
nand U13511 (N_13511,N_10416,N_10960);
and U13512 (N_13512,N_10901,N_10950);
and U13513 (N_13513,N_10615,N_10415);
nor U13514 (N_13514,N_10103,N_10650);
nor U13515 (N_13515,N_11689,N_10376);
nor U13516 (N_13516,N_10258,N_11231);
or U13517 (N_13517,N_10698,N_11743);
and U13518 (N_13518,N_11515,N_10258);
and U13519 (N_13519,N_11971,N_11937);
nand U13520 (N_13520,N_10862,N_10083);
nand U13521 (N_13521,N_10051,N_11879);
nor U13522 (N_13522,N_11466,N_10178);
nand U13523 (N_13523,N_11764,N_10327);
nor U13524 (N_13524,N_11227,N_11177);
nand U13525 (N_13525,N_11889,N_10517);
or U13526 (N_13526,N_11582,N_10307);
nand U13527 (N_13527,N_11592,N_10189);
and U13528 (N_13528,N_10730,N_10960);
or U13529 (N_13529,N_10617,N_10955);
nand U13530 (N_13530,N_10892,N_11848);
nor U13531 (N_13531,N_11628,N_11099);
and U13532 (N_13532,N_11398,N_10336);
nor U13533 (N_13533,N_10996,N_10339);
or U13534 (N_13534,N_10805,N_11827);
nand U13535 (N_13535,N_10677,N_11857);
nand U13536 (N_13536,N_10235,N_10396);
nor U13537 (N_13537,N_10233,N_11807);
nor U13538 (N_13538,N_10266,N_11419);
or U13539 (N_13539,N_11711,N_11552);
or U13540 (N_13540,N_10841,N_10440);
or U13541 (N_13541,N_11391,N_11420);
nor U13542 (N_13542,N_10113,N_11045);
nand U13543 (N_13543,N_11360,N_10020);
nor U13544 (N_13544,N_10272,N_11275);
and U13545 (N_13545,N_11555,N_10167);
or U13546 (N_13546,N_10826,N_11441);
or U13547 (N_13547,N_11162,N_10111);
nor U13548 (N_13548,N_10792,N_10615);
or U13549 (N_13549,N_10167,N_11287);
nor U13550 (N_13550,N_11648,N_11166);
nand U13551 (N_13551,N_11188,N_10534);
and U13552 (N_13552,N_10114,N_10058);
nor U13553 (N_13553,N_10943,N_10669);
or U13554 (N_13554,N_10402,N_11471);
and U13555 (N_13555,N_10316,N_10313);
and U13556 (N_13556,N_10533,N_11122);
xnor U13557 (N_13557,N_10321,N_10724);
xor U13558 (N_13558,N_10203,N_10597);
or U13559 (N_13559,N_10018,N_10019);
nand U13560 (N_13560,N_10024,N_11985);
nor U13561 (N_13561,N_11022,N_10317);
nand U13562 (N_13562,N_10522,N_10055);
xor U13563 (N_13563,N_11969,N_10893);
nand U13564 (N_13564,N_10650,N_11509);
or U13565 (N_13565,N_10678,N_10165);
nand U13566 (N_13566,N_11887,N_10051);
nor U13567 (N_13567,N_11161,N_11618);
xor U13568 (N_13568,N_10076,N_11277);
and U13569 (N_13569,N_11638,N_10007);
nor U13570 (N_13570,N_11152,N_11299);
or U13571 (N_13571,N_11094,N_11749);
nand U13572 (N_13572,N_11672,N_10361);
nor U13573 (N_13573,N_10312,N_11799);
nor U13574 (N_13574,N_10302,N_11630);
nor U13575 (N_13575,N_11648,N_10849);
or U13576 (N_13576,N_10205,N_10689);
nand U13577 (N_13577,N_10077,N_10342);
or U13578 (N_13578,N_10694,N_11491);
or U13579 (N_13579,N_10422,N_10146);
xor U13580 (N_13580,N_11313,N_10031);
and U13581 (N_13581,N_10904,N_10635);
nand U13582 (N_13582,N_11814,N_11516);
nor U13583 (N_13583,N_11288,N_10269);
and U13584 (N_13584,N_10343,N_10604);
nand U13585 (N_13585,N_10766,N_10224);
xnor U13586 (N_13586,N_10246,N_11413);
and U13587 (N_13587,N_11338,N_11546);
xor U13588 (N_13588,N_10967,N_11970);
or U13589 (N_13589,N_11659,N_11594);
and U13590 (N_13590,N_11107,N_10841);
nor U13591 (N_13591,N_11678,N_10256);
and U13592 (N_13592,N_11034,N_11283);
nor U13593 (N_13593,N_11976,N_11702);
nor U13594 (N_13594,N_11146,N_10172);
or U13595 (N_13595,N_11704,N_10496);
or U13596 (N_13596,N_11396,N_10965);
nand U13597 (N_13597,N_11613,N_11734);
nor U13598 (N_13598,N_10770,N_11109);
xnor U13599 (N_13599,N_11347,N_10857);
nor U13600 (N_13600,N_11810,N_11202);
or U13601 (N_13601,N_10552,N_10132);
nand U13602 (N_13602,N_11163,N_10265);
nand U13603 (N_13603,N_10150,N_10072);
nand U13604 (N_13604,N_10315,N_10070);
nor U13605 (N_13605,N_10777,N_11858);
or U13606 (N_13606,N_11750,N_10995);
and U13607 (N_13607,N_11799,N_10497);
or U13608 (N_13608,N_10757,N_11879);
nand U13609 (N_13609,N_10625,N_10265);
nand U13610 (N_13610,N_10063,N_11366);
and U13611 (N_13611,N_10846,N_10006);
or U13612 (N_13612,N_10422,N_11202);
xor U13613 (N_13613,N_11955,N_11714);
and U13614 (N_13614,N_11368,N_10312);
or U13615 (N_13615,N_10147,N_10442);
nand U13616 (N_13616,N_10421,N_11869);
or U13617 (N_13617,N_10269,N_11747);
nand U13618 (N_13618,N_11781,N_11252);
nor U13619 (N_13619,N_11338,N_11234);
nor U13620 (N_13620,N_10914,N_10658);
nand U13621 (N_13621,N_10274,N_11808);
and U13622 (N_13622,N_11868,N_11247);
or U13623 (N_13623,N_11420,N_10564);
or U13624 (N_13624,N_10225,N_11930);
nor U13625 (N_13625,N_11840,N_11665);
and U13626 (N_13626,N_10055,N_11236);
or U13627 (N_13627,N_11905,N_10265);
nand U13628 (N_13628,N_11459,N_11095);
or U13629 (N_13629,N_11770,N_11092);
or U13630 (N_13630,N_11809,N_10584);
and U13631 (N_13631,N_10649,N_11304);
nor U13632 (N_13632,N_11433,N_11839);
or U13633 (N_13633,N_11782,N_11489);
and U13634 (N_13634,N_10639,N_11414);
and U13635 (N_13635,N_10290,N_10055);
nor U13636 (N_13636,N_11207,N_11851);
nor U13637 (N_13637,N_11569,N_11435);
or U13638 (N_13638,N_11962,N_10344);
nand U13639 (N_13639,N_11455,N_11641);
and U13640 (N_13640,N_10971,N_10426);
nand U13641 (N_13641,N_11263,N_11803);
nor U13642 (N_13642,N_11727,N_10204);
nor U13643 (N_13643,N_11885,N_11236);
nor U13644 (N_13644,N_11119,N_11101);
nor U13645 (N_13645,N_11951,N_11476);
or U13646 (N_13646,N_10078,N_11986);
nor U13647 (N_13647,N_10592,N_11604);
xor U13648 (N_13648,N_11061,N_10372);
and U13649 (N_13649,N_10480,N_10554);
or U13650 (N_13650,N_10220,N_11400);
or U13651 (N_13651,N_10591,N_10313);
and U13652 (N_13652,N_11205,N_10386);
nand U13653 (N_13653,N_10489,N_11094);
and U13654 (N_13654,N_11435,N_11200);
xor U13655 (N_13655,N_11014,N_11359);
xnor U13656 (N_13656,N_11162,N_11249);
nand U13657 (N_13657,N_10702,N_10527);
and U13658 (N_13658,N_11777,N_10689);
nor U13659 (N_13659,N_10664,N_10227);
xor U13660 (N_13660,N_10505,N_11069);
nor U13661 (N_13661,N_11282,N_10470);
or U13662 (N_13662,N_10880,N_11781);
nand U13663 (N_13663,N_10349,N_10647);
or U13664 (N_13664,N_11732,N_10906);
nand U13665 (N_13665,N_10630,N_11859);
or U13666 (N_13666,N_11597,N_10993);
nand U13667 (N_13667,N_10166,N_11891);
and U13668 (N_13668,N_10289,N_10411);
nand U13669 (N_13669,N_10170,N_11418);
nand U13670 (N_13670,N_11544,N_11564);
nand U13671 (N_13671,N_11374,N_11156);
or U13672 (N_13672,N_10299,N_10025);
or U13673 (N_13673,N_10288,N_11701);
nand U13674 (N_13674,N_11346,N_10179);
or U13675 (N_13675,N_10524,N_11606);
nand U13676 (N_13676,N_11057,N_11127);
nor U13677 (N_13677,N_10716,N_11709);
nand U13678 (N_13678,N_11320,N_10975);
nand U13679 (N_13679,N_11561,N_10232);
nand U13680 (N_13680,N_11604,N_11957);
nand U13681 (N_13681,N_11909,N_11308);
xnor U13682 (N_13682,N_11748,N_11083);
or U13683 (N_13683,N_10497,N_11279);
nor U13684 (N_13684,N_10672,N_10423);
nand U13685 (N_13685,N_10440,N_11233);
nor U13686 (N_13686,N_11781,N_11299);
nand U13687 (N_13687,N_10249,N_11691);
and U13688 (N_13688,N_11960,N_11000);
nand U13689 (N_13689,N_11430,N_10502);
and U13690 (N_13690,N_10588,N_10024);
and U13691 (N_13691,N_10385,N_11635);
nand U13692 (N_13692,N_11839,N_10279);
or U13693 (N_13693,N_11535,N_11880);
or U13694 (N_13694,N_11007,N_10324);
nor U13695 (N_13695,N_11586,N_10026);
and U13696 (N_13696,N_11760,N_10181);
nor U13697 (N_13697,N_11754,N_10789);
nor U13698 (N_13698,N_11553,N_10315);
and U13699 (N_13699,N_11409,N_11689);
nand U13700 (N_13700,N_10718,N_11901);
nor U13701 (N_13701,N_11615,N_10132);
nand U13702 (N_13702,N_10027,N_11086);
nor U13703 (N_13703,N_11227,N_11092);
or U13704 (N_13704,N_11833,N_11740);
and U13705 (N_13705,N_10644,N_11656);
nor U13706 (N_13706,N_10072,N_11221);
or U13707 (N_13707,N_11930,N_11323);
nand U13708 (N_13708,N_11452,N_11560);
nand U13709 (N_13709,N_11280,N_11845);
nor U13710 (N_13710,N_11007,N_11593);
xnor U13711 (N_13711,N_11547,N_11369);
and U13712 (N_13712,N_10175,N_10870);
and U13713 (N_13713,N_10510,N_11665);
or U13714 (N_13714,N_10615,N_10248);
and U13715 (N_13715,N_10218,N_11336);
and U13716 (N_13716,N_11805,N_10984);
nor U13717 (N_13717,N_11660,N_10023);
nor U13718 (N_13718,N_10716,N_10803);
and U13719 (N_13719,N_10443,N_10807);
and U13720 (N_13720,N_10811,N_11929);
xnor U13721 (N_13721,N_10091,N_10742);
and U13722 (N_13722,N_11678,N_11551);
or U13723 (N_13723,N_10948,N_10701);
nor U13724 (N_13724,N_11682,N_11003);
or U13725 (N_13725,N_11161,N_10085);
nor U13726 (N_13726,N_11191,N_11613);
nor U13727 (N_13727,N_10419,N_10778);
or U13728 (N_13728,N_11439,N_11903);
or U13729 (N_13729,N_10977,N_10263);
and U13730 (N_13730,N_10683,N_10812);
nand U13731 (N_13731,N_10495,N_10106);
and U13732 (N_13732,N_11381,N_10514);
and U13733 (N_13733,N_10188,N_10990);
xnor U13734 (N_13734,N_10442,N_11245);
nor U13735 (N_13735,N_11013,N_11806);
and U13736 (N_13736,N_10214,N_11683);
nor U13737 (N_13737,N_11012,N_11909);
or U13738 (N_13738,N_10179,N_10482);
xor U13739 (N_13739,N_11453,N_11577);
nor U13740 (N_13740,N_11788,N_10689);
and U13741 (N_13741,N_10775,N_10090);
nor U13742 (N_13742,N_10153,N_11359);
nand U13743 (N_13743,N_11960,N_10264);
nor U13744 (N_13744,N_11082,N_11010);
or U13745 (N_13745,N_11406,N_10086);
nand U13746 (N_13746,N_10204,N_10112);
and U13747 (N_13747,N_11604,N_11246);
and U13748 (N_13748,N_11063,N_11229);
or U13749 (N_13749,N_11224,N_10638);
nor U13750 (N_13750,N_10496,N_10338);
and U13751 (N_13751,N_11204,N_11099);
nand U13752 (N_13752,N_11333,N_11917);
xnor U13753 (N_13753,N_11222,N_11022);
or U13754 (N_13754,N_11302,N_11200);
nand U13755 (N_13755,N_11032,N_10599);
and U13756 (N_13756,N_11952,N_10071);
or U13757 (N_13757,N_11932,N_11260);
nor U13758 (N_13758,N_11994,N_10510);
nand U13759 (N_13759,N_11213,N_11621);
and U13760 (N_13760,N_11073,N_11534);
or U13761 (N_13761,N_11514,N_10082);
nor U13762 (N_13762,N_11967,N_11592);
nor U13763 (N_13763,N_11199,N_11884);
nor U13764 (N_13764,N_10067,N_11671);
nand U13765 (N_13765,N_11234,N_11713);
or U13766 (N_13766,N_10856,N_10672);
nor U13767 (N_13767,N_10391,N_10071);
nor U13768 (N_13768,N_11368,N_10620);
and U13769 (N_13769,N_11256,N_11962);
or U13770 (N_13770,N_11935,N_11551);
nand U13771 (N_13771,N_10703,N_11543);
or U13772 (N_13772,N_11635,N_11802);
or U13773 (N_13773,N_11713,N_11940);
nand U13774 (N_13774,N_10157,N_11320);
nand U13775 (N_13775,N_10523,N_11749);
nor U13776 (N_13776,N_10453,N_11062);
nand U13777 (N_13777,N_10761,N_11606);
and U13778 (N_13778,N_11382,N_10429);
and U13779 (N_13779,N_10559,N_10286);
nor U13780 (N_13780,N_11145,N_11701);
or U13781 (N_13781,N_11117,N_11004);
xnor U13782 (N_13782,N_11040,N_11470);
and U13783 (N_13783,N_11641,N_11625);
nor U13784 (N_13784,N_11963,N_10689);
nand U13785 (N_13785,N_11689,N_10801);
nand U13786 (N_13786,N_11899,N_11843);
nand U13787 (N_13787,N_10609,N_11132);
xor U13788 (N_13788,N_10966,N_11198);
or U13789 (N_13789,N_11148,N_11927);
nand U13790 (N_13790,N_11569,N_11750);
nand U13791 (N_13791,N_10628,N_10919);
nor U13792 (N_13792,N_11364,N_11632);
nor U13793 (N_13793,N_10763,N_11991);
nand U13794 (N_13794,N_10895,N_10409);
nor U13795 (N_13795,N_11082,N_11085);
nand U13796 (N_13796,N_10574,N_10551);
nor U13797 (N_13797,N_11448,N_10932);
nor U13798 (N_13798,N_10087,N_11005);
and U13799 (N_13799,N_11202,N_10078);
xnor U13800 (N_13800,N_10327,N_11241);
or U13801 (N_13801,N_10581,N_10297);
nor U13802 (N_13802,N_10848,N_10031);
or U13803 (N_13803,N_10195,N_10086);
and U13804 (N_13804,N_11235,N_11987);
nand U13805 (N_13805,N_10528,N_10395);
nor U13806 (N_13806,N_11204,N_10658);
and U13807 (N_13807,N_11646,N_10271);
nand U13808 (N_13808,N_10311,N_11200);
nand U13809 (N_13809,N_10362,N_11140);
and U13810 (N_13810,N_10306,N_10536);
or U13811 (N_13811,N_10793,N_11188);
or U13812 (N_13812,N_11723,N_11916);
nand U13813 (N_13813,N_10760,N_11115);
nand U13814 (N_13814,N_10877,N_11600);
and U13815 (N_13815,N_11543,N_10014);
or U13816 (N_13816,N_10352,N_11379);
and U13817 (N_13817,N_10936,N_10747);
nor U13818 (N_13818,N_11736,N_10872);
nor U13819 (N_13819,N_10617,N_11076);
xnor U13820 (N_13820,N_11293,N_11184);
and U13821 (N_13821,N_11145,N_11248);
nor U13822 (N_13822,N_11941,N_10400);
nand U13823 (N_13823,N_11850,N_10432);
and U13824 (N_13824,N_11346,N_11334);
and U13825 (N_13825,N_11845,N_10435);
xnor U13826 (N_13826,N_11529,N_11739);
nand U13827 (N_13827,N_11612,N_11108);
or U13828 (N_13828,N_10647,N_10398);
and U13829 (N_13829,N_11136,N_10154);
or U13830 (N_13830,N_11130,N_11345);
nor U13831 (N_13831,N_10591,N_11030);
and U13832 (N_13832,N_10190,N_11054);
nor U13833 (N_13833,N_10879,N_11577);
nor U13834 (N_13834,N_10545,N_10118);
nor U13835 (N_13835,N_10764,N_11787);
nand U13836 (N_13836,N_11992,N_10476);
xor U13837 (N_13837,N_11296,N_10160);
and U13838 (N_13838,N_10637,N_11533);
or U13839 (N_13839,N_11262,N_10697);
nor U13840 (N_13840,N_10662,N_11212);
or U13841 (N_13841,N_11398,N_10361);
and U13842 (N_13842,N_11160,N_10743);
xor U13843 (N_13843,N_10862,N_10484);
nand U13844 (N_13844,N_11804,N_10512);
nand U13845 (N_13845,N_10968,N_11300);
and U13846 (N_13846,N_11868,N_10803);
xor U13847 (N_13847,N_10197,N_10531);
nand U13848 (N_13848,N_10020,N_10900);
or U13849 (N_13849,N_10058,N_10899);
and U13850 (N_13850,N_11206,N_10988);
nor U13851 (N_13851,N_11374,N_10716);
and U13852 (N_13852,N_11411,N_10684);
and U13853 (N_13853,N_10021,N_10737);
nand U13854 (N_13854,N_10009,N_11709);
nor U13855 (N_13855,N_10448,N_10596);
nor U13856 (N_13856,N_11753,N_11052);
or U13857 (N_13857,N_11603,N_10164);
nor U13858 (N_13858,N_11673,N_10262);
nand U13859 (N_13859,N_11999,N_11298);
or U13860 (N_13860,N_10915,N_10242);
nand U13861 (N_13861,N_11267,N_10608);
and U13862 (N_13862,N_11069,N_10480);
and U13863 (N_13863,N_10579,N_10154);
and U13864 (N_13864,N_11923,N_10264);
nand U13865 (N_13865,N_10206,N_11337);
nor U13866 (N_13866,N_10552,N_10071);
nand U13867 (N_13867,N_11528,N_11341);
or U13868 (N_13868,N_10253,N_10713);
or U13869 (N_13869,N_11076,N_11568);
nor U13870 (N_13870,N_11043,N_11345);
xor U13871 (N_13871,N_11979,N_10130);
and U13872 (N_13872,N_10256,N_11429);
and U13873 (N_13873,N_11795,N_10587);
or U13874 (N_13874,N_11700,N_10029);
nand U13875 (N_13875,N_11540,N_11575);
or U13876 (N_13876,N_11332,N_10991);
nor U13877 (N_13877,N_10062,N_11264);
nor U13878 (N_13878,N_11826,N_10196);
nor U13879 (N_13879,N_10202,N_10884);
nand U13880 (N_13880,N_10865,N_10213);
or U13881 (N_13881,N_10246,N_11280);
nand U13882 (N_13882,N_10318,N_11528);
and U13883 (N_13883,N_11447,N_10543);
or U13884 (N_13884,N_10826,N_10173);
and U13885 (N_13885,N_10204,N_11810);
nand U13886 (N_13886,N_10485,N_10106);
or U13887 (N_13887,N_11211,N_10192);
and U13888 (N_13888,N_10331,N_11038);
and U13889 (N_13889,N_10970,N_10050);
nand U13890 (N_13890,N_10831,N_10982);
nand U13891 (N_13891,N_11145,N_11676);
and U13892 (N_13892,N_11107,N_10788);
and U13893 (N_13893,N_11021,N_11755);
nor U13894 (N_13894,N_10503,N_11725);
nand U13895 (N_13895,N_11387,N_10625);
or U13896 (N_13896,N_10678,N_10273);
xor U13897 (N_13897,N_10087,N_11335);
or U13898 (N_13898,N_11605,N_10075);
or U13899 (N_13899,N_11053,N_11576);
and U13900 (N_13900,N_11405,N_10191);
nor U13901 (N_13901,N_10585,N_11626);
and U13902 (N_13902,N_10165,N_11558);
and U13903 (N_13903,N_10039,N_11479);
and U13904 (N_13904,N_11098,N_10094);
xnor U13905 (N_13905,N_10858,N_10499);
nor U13906 (N_13906,N_10561,N_11684);
xnor U13907 (N_13907,N_10459,N_10758);
and U13908 (N_13908,N_10793,N_11881);
nand U13909 (N_13909,N_11887,N_11892);
nand U13910 (N_13910,N_11997,N_10913);
xor U13911 (N_13911,N_11049,N_11291);
or U13912 (N_13912,N_10951,N_11747);
xnor U13913 (N_13913,N_11513,N_10301);
and U13914 (N_13914,N_11273,N_10330);
nor U13915 (N_13915,N_10444,N_10497);
xor U13916 (N_13916,N_11375,N_10504);
or U13917 (N_13917,N_10292,N_11481);
and U13918 (N_13918,N_10405,N_10194);
xnor U13919 (N_13919,N_10216,N_11180);
or U13920 (N_13920,N_11956,N_11991);
and U13921 (N_13921,N_11401,N_10875);
or U13922 (N_13922,N_10799,N_10476);
and U13923 (N_13923,N_11228,N_10163);
nor U13924 (N_13924,N_10660,N_10003);
or U13925 (N_13925,N_10519,N_10051);
nand U13926 (N_13926,N_11364,N_11280);
nor U13927 (N_13927,N_10336,N_10383);
xor U13928 (N_13928,N_11203,N_11811);
nor U13929 (N_13929,N_11497,N_11733);
nor U13930 (N_13930,N_11923,N_11550);
nand U13931 (N_13931,N_10538,N_11425);
nand U13932 (N_13932,N_11332,N_11953);
nand U13933 (N_13933,N_10295,N_11796);
and U13934 (N_13934,N_11850,N_10323);
nor U13935 (N_13935,N_10014,N_11762);
nand U13936 (N_13936,N_11247,N_10379);
and U13937 (N_13937,N_11362,N_10026);
nor U13938 (N_13938,N_11016,N_10060);
nand U13939 (N_13939,N_11787,N_10564);
or U13940 (N_13940,N_11599,N_10052);
nand U13941 (N_13941,N_10354,N_11052);
nor U13942 (N_13942,N_11932,N_10645);
nor U13943 (N_13943,N_10794,N_11855);
or U13944 (N_13944,N_11819,N_10538);
and U13945 (N_13945,N_11665,N_11311);
or U13946 (N_13946,N_10644,N_11689);
or U13947 (N_13947,N_10850,N_10128);
and U13948 (N_13948,N_10374,N_10471);
or U13949 (N_13949,N_11335,N_11380);
nor U13950 (N_13950,N_10967,N_11674);
and U13951 (N_13951,N_11953,N_11374);
and U13952 (N_13952,N_10427,N_10628);
or U13953 (N_13953,N_10581,N_10247);
nand U13954 (N_13954,N_10640,N_10207);
nand U13955 (N_13955,N_10246,N_10573);
xor U13956 (N_13956,N_11068,N_10106);
xnor U13957 (N_13957,N_11730,N_11119);
xnor U13958 (N_13958,N_11759,N_10365);
nand U13959 (N_13959,N_10048,N_11924);
nand U13960 (N_13960,N_10747,N_10014);
and U13961 (N_13961,N_11606,N_11054);
nor U13962 (N_13962,N_10157,N_11754);
and U13963 (N_13963,N_10070,N_10768);
or U13964 (N_13964,N_11488,N_10188);
nor U13965 (N_13965,N_10508,N_11890);
and U13966 (N_13966,N_10891,N_11211);
nand U13967 (N_13967,N_10366,N_10630);
nand U13968 (N_13968,N_11733,N_10782);
and U13969 (N_13969,N_11642,N_11542);
xor U13970 (N_13970,N_10453,N_11785);
or U13971 (N_13971,N_10227,N_11454);
xor U13972 (N_13972,N_10464,N_10203);
nand U13973 (N_13973,N_10346,N_11238);
nand U13974 (N_13974,N_11797,N_11326);
nand U13975 (N_13975,N_10799,N_10335);
and U13976 (N_13976,N_10622,N_10398);
or U13977 (N_13977,N_10638,N_11948);
nand U13978 (N_13978,N_10332,N_11900);
nor U13979 (N_13979,N_11561,N_11557);
nor U13980 (N_13980,N_10970,N_11719);
xnor U13981 (N_13981,N_10410,N_11321);
or U13982 (N_13982,N_10327,N_11027);
nor U13983 (N_13983,N_10094,N_10860);
and U13984 (N_13984,N_11698,N_11496);
or U13985 (N_13985,N_11509,N_11902);
nand U13986 (N_13986,N_10859,N_10819);
and U13987 (N_13987,N_10839,N_11619);
or U13988 (N_13988,N_11374,N_11249);
and U13989 (N_13989,N_11446,N_10522);
and U13990 (N_13990,N_10625,N_11575);
nand U13991 (N_13991,N_11490,N_11556);
and U13992 (N_13992,N_11074,N_10711);
and U13993 (N_13993,N_11935,N_11216);
and U13994 (N_13994,N_10940,N_10559);
nand U13995 (N_13995,N_11040,N_10493);
and U13996 (N_13996,N_10979,N_11339);
and U13997 (N_13997,N_10966,N_10230);
nor U13998 (N_13998,N_11235,N_11658);
or U13999 (N_13999,N_11296,N_10963);
xor U14000 (N_14000,N_12329,N_12196);
nand U14001 (N_14001,N_12253,N_12827);
nand U14002 (N_14002,N_13569,N_12554);
xor U14003 (N_14003,N_12027,N_12607);
xnor U14004 (N_14004,N_13063,N_12986);
nor U14005 (N_14005,N_12785,N_13923);
or U14006 (N_14006,N_13904,N_12793);
or U14007 (N_14007,N_13401,N_12468);
or U14008 (N_14008,N_12127,N_12474);
and U14009 (N_14009,N_13051,N_13842);
nand U14010 (N_14010,N_13599,N_13228);
nand U14011 (N_14011,N_13490,N_12997);
and U14012 (N_14012,N_12804,N_12859);
nor U14013 (N_14013,N_12886,N_13359);
xnor U14014 (N_14014,N_13552,N_12349);
nand U14015 (N_14015,N_12783,N_12299);
or U14016 (N_14016,N_13043,N_13493);
nor U14017 (N_14017,N_12972,N_12897);
nand U14018 (N_14018,N_13033,N_13297);
or U14019 (N_14019,N_13915,N_13361);
xor U14020 (N_14020,N_12824,N_13762);
xor U14021 (N_14021,N_13191,N_13554);
nor U14022 (N_14022,N_13933,N_13778);
and U14023 (N_14023,N_13965,N_13622);
or U14024 (N_14024,N_12216,N_12991);
nor U14025 (N_14025,N_13529,N_13294);
and U14026 (N_14026,N_12403,N_13031);
or U14027 (N_14027,N_12666,N_12985);
or U14028 (N_14028,N_13543,N_12105);
nand U14029 (N_14029,N_12614,N_13258);
or U14030 (N_14030,N_13626,N_13068);
and U14031 (N_14031,N_13208,N_13335);
or U14032 (N_14032,N_13917,N_13269);
nor U14033 (N_14033,N_12344,N_13365);
nor U14034 (N_14034,N_12906,N_12051);
nand U14035 (N_14035,N_13032,N_13832);
xnor U14036 (N_14036,N_12592,N_13675);
nand U14037 (N_14037,N_12097,N_13038);
xor U14038 (N_14038,N_12084,N_13467);
or U14039 (N_14039,N_13021,N_13541);
xnor U14040 (N_14040,N_13664,N_12915);
nand U14041 (N_14041,N_12655,N_13607);
or U14042 (N_14042,N_13851,N_13124);
nor U14043 (N_14043,N_12045,N_13942);
or U14044 (N_14044,N_13636,N_13586);
nand U14045 (N_14045,N_12810,N_13653);
or U14046 (N_14046,N_13057,N_13756);
and U14047 (N_14047,N_13134,N_12817);
xor U14048 (N_14048,N_12266,N_13557);
or U14049 (N_14049,N_12022,N_12619);
and U14050 (N_14050,N_13632,N_12589);
xnor U14051 (N_14051,N_13432,N_13555);
nor U14052 (N_14052,N_13873,N_13691);
or U14053 (N_14053,N_13864,N_13506);
nor U14054 (N_14054,N_13821,N_13396);
nor U14055 (N_14055,N_13265,N_13002);
nor U14056 (N_14056,N_12716,N_12364);
nand U14057 (N_14057,N_13517,N_12070);
or U14058 (N_14058,N_12860,N_12363);
and U14059 (N_14059,N_13480,N_13431);
xor U14060 (N_14060,N_12434,N_12085);
or U14061 (N_14061,N_13282,N_12375);
and U14062 (N_14062,N_13181,N_12815);
and U14063 (N_14063,N_13098,N_12422);
nand U14064 (N_14064,N_13822,N_13651);
nand U14065 (N_14065,N_12752,N_12709);
and U14066 (N_14066,N_12324,N_13340);
or U14067 (N_14067,N_12981,N_12534);
nand U14068 (N_14068,N_12365,N_13001);
nor U14069 (N_14069,N_12521,N_13080);
or U14070 (N_14070,N_13234,N_12994);
xnor U14071 (N_14071,N_12863,N_13852);
and U14072 (N_14072,N_13511,N_12154);
xor U14073 (N_14073,N_12703,N_12917);
or U14074 (N_14074,N_13833,N_12779);
nand U14075 (N_14075,N_12290,N_13922);
or U14076 (N_14076,N_13072,N_13302);
nor U14077 (N_14077,N_13966,N_13752);
xnor U14078 (N_14078,N_13266,N_13379);
or U14079 (N_14079,N_13790,N_12420);
or U14080 (N_14080,N_12932,N_12770);
or U14081 (N_14081,N_12499,N_12160);
nand U14082 (N_14082,N_13666,N_13686);
xnor U14083 (N_14083,N_13152,N_13947);
nor U14084 (N_14084,N_12660,N_13188);
xor U14085 (N_14085,N_13869,N_12242);
xor U14086 (N_14086,N_12472,N_12285);
nor U14087 (N_14087,N_12690,N_12314);
and U14088 (N_14088,N_13360,N_13699);
and U14089 (N_14089,N_13180,N_12901);
or U14090 (N_14090,N_13993,N_12280);
nor U14091 (N_14091,N_12912,N_12822);
nand U14092 (N_14092,N_12524,N_13624);
nand U14093 (N_14093,N_13680,N_12147);
nand U14094 (N_14094,N_13352,N_12203);
or U14095 (N_14095,N_13663,N_12724);
nor U14096 (N_14096,N_12899,N_13391);
or U14097 (N_14097,N_12020,N_12234);
nor U14098 (N_14098,N_13547,N_13542);
xnor U14099 (N_14099,N_13026,N_13217);
nand U14100 (N_14100,N_12872,N_13184);
nand U14101 (N_14101,N_12294,N_12565);
and U14102 (N_14102,N_12193,N_13908);
nor U14103 (N_14103,N_13816,N_12271);
and U14104 (N_14104,N_12381,N_12278);
nor U14105 (N_14105,N_13408,N_12327);
and U14106 (N_14106,N_13447,N_13924);
nand U14107 (N_14107,N_13956,N_13545);
nand U14108 (N_14108,N_13466,N_12388);
nand U14109 (N_14109,N_12223,N_12746);
xnor U14110 (N_14110,N_12797,N_12830);
and U14111 (N_14111,N_13201,N_12941);
xnor U14112 (N_14112,N_12118,N_13196);
and U14113 (N_14113,N_13795,N_13395);
or U14114 (N_14114,N_13958,N_13149);
nor U14115 (N_14115,N_12428,N_12873);
or U14116 (N_14116,N_13382,N_12228);
xor U14117 (N_14117,N_12615,N_12214);
or U14118 (N_14118,N_12251,N_13829);
xor U14119 (N_14119,N_12457,N_13327);
or U14120 (N_14120,N_13682,N_12158);
nor U14121 (N_14121,N_13276,N_12907);
and U14122 (N_14122,N_12588,N_13536);
or U14123 (N_14123,N_13847,N_12751);
nand U14124 (N_14124,N_12951,N_12865);
and U14125 (N_14125,N_13755,N_12777);
or U14126 (N_14126,N_13777,N_13830);
nor U14127 (N_14127,N_13916,N_12547);
or U14128 (N_14128,N_13433,N_12340);
nand U14129 (N_14129,N_12961,N_12958);
nor U14130 (N_14130,N_13377,N_13901);
and U14131 (N_14131,N_13561,N_13267);
nand U14132 (N_14132,N_12023,N_12689);
and U14133 (N_14133,N_12397,N_13350);
and U14134 (N_14134,N_12651,N_13837);
or U14135 (N_14135,N_12453,N_13040);
or U14136 (N_14136,N_12864,N_12210);
nor U14137 (N_14137,N_12080,N_12707);
or U14138 (N_14138,N_13619,N_12150);
nand U14139 (N_14139,N_12634,N_13973);
and U14140 (N_14140,N_13522,N_13528);
nor U14141 (N_14141,N_12957,N_12336);
or U14142 (N_14142,N_12106,N_13088);
or U14143 (N_14143,N_12055,N_13270);
and U14144 (N_14144,N_13415,N_13248);
nand U14145 (N_14145,N_12583,N_13027);
nand U14146 (N_14146,N_13419,N_13696);
and U14147 (N_14147,N_13717,N_12398);
nor U14148 (N_14148,N_12888,N_13252);
nor U14149 (N_14149,N_12005,N_12167);
nor U14150 (N_14150,N_12509,N_13605);
xnor U14151 (N_14151,N_13398,N_12878);
nor U14152 (N_14152,N_13338,N_12870);
or U14153 (N_14153,N_13113,N_12303);
xnor U14154 (N_14154,N_13598,N_13912);
xor U14155 (N_14155,N_13742,N_12676);
or U14156 (N_14156,N_12369,N_12247);
xor U14157 (N_14157,N_12169,N_12077);
xnor U14158 (N_14158,N_12302,N_12675);
or U14159 (N_14159,N_13858,N_13060);
nor U14160 (N_14160,N_13895,N_13714);
xnor U14161 (N_14161,N_12012,N_12177);
xnor U14162 (N_14162,N_12538,N_13123);
xor U14163 (N_14163,N_12248,N_13175);
or U14164 (N_14164,N_13865,N_13584);
or U14165 (N_14165,N_12699,N_13678);
and U14166 (N_14166,N_13962,N_13206);
nor U14167 (N_14167,N_12514,N_13483);
and U14168 (N_14168,N_13285,N_12416);
and U14169 (N_14169,N_13150,N_13177);
nand U14170 (N_14170,N_12125,N_12198);
or U14171 (N_14171,N_12652,N_13176);
and U14172 (N_14172,N_12025,N_12479);
or U14173 (N_14173,N_13496,N_13156);
nand U14174 (N_14174,N_12813,N_12663);
or U14175 (N_14175,N_13320,N_12325);
and U14176 (N_14176,N_13504,N_13676);
nand U14177 (N_14177,N_12575,N_13044);
and U14178 (N_14178,N_12673,N_13179);
nand U14179 (N_14179,N_13799,N_13512);
nor U14180 (N_14180,N_13802,N_13216);
nand U14181 (N_14181,N_13787,N_13418);
and U14182 (N_14182,N_13289,N_12979);
and U14183 (N_14183,N_13214,N_12421);
and U14184 (N_14184,N_13295,N_12180);
nor U14185 (N_14185,N_12747,N_12066);
xnor U14186 (N_14186,N_13107,N_12227);
xor U14187 (N_14187,N_13783,N_13929);
and U14188 (N_14188,N_12465,N_13960);
or U14189 (N_14189,N_12875,N_12186);
nand U14190 (N_14190,N_13478,N_13934);
and U14191 (N_14191,N_12535,N_13463);
and U14192 (N_14192,N_12636,N_13299);
and U14193 (N_14193,N_13951,N_13307);
nor U14194 (N_14194,N_13640,N_13715);
and U14195 (N_14195,N_13948,N_12653);
and U14196 (N_14196,N_13223,N_13709);
or U14197 (N_14197,N_12714,N_12750);
or U14198 (N_14198,N_12555,N_12502);
nand U14199 (N_14199,N_12123,N_12425);
or U14200 (N_14200,N_12343,N_13954);
or U14201 (N_14201,N_12373,N_12723);
and U14202 (N_14202,N_12182,N_13215);
and U14203 (N_14203,N_13079,N_12739);
xor U14204 (N_14204,N_12570,N_13355);
and U14205 (N_14205,N_13684,N_13913);
and U14206 (N_14206,N_13236,N_13314);
nor U14207 (N_14207,N_13066,N_12506);
xnor U14208 (N_14208,N_12181,N_12984);
and U14209 (N_14209,N_13878,N_13055);
nand U14210 (N_14210,N_12036,N_12389);
and U14211 (N_14211,N_12600,N_13747);
or U14212 (N_14212,N_13977,N_12530);
xor U14213 (N_14213,N_12488,N_12518);
nand U14214 (N_14214,N_12602,N_12871);
nor U14215 (N_14215,N_12862,N_13000);
or U14216 (N_14216,N_13671,N_13981);
nor U14217 (N_14217,N_13472,N_12031);
nand U14218 (N_14218,N_13311,N_13337);
xnor U14219 (N_14219,N_13053,N_13674);
or U14220 (N_14220,N_12613,N_13259);
and U14221 (N_14221,N_13054,N_13871);
nand U14222 (N_14222,N_13067,N_13559);
nor U14223 (N_14223,N_12441,N_13119);
nand U14224 (N_14224,N_13999,N_12047);
or U14225 (N_14225,N_13899,N_12372);
nor U14226 (N_14226,N_13754,N_13101);
or U14227 (N_14227,N_13109,N_12894);
nor U14228 (N_14228,N_13698,N_12069);
and U14229 (N_14229,N_13817,N_12470);
nand U14230 (N_14230,N_12559,N_13120);
xnor U14231 (N_14231,N_13527,N_12350);
and U14232 (N_14232,N_13994,N_12654);
and U14233 (N_14233,N_13660,N_12283);
nand U14234 (N_14234,N_12443,N_12816);
or U14235 (N_14235,N_13405,N_13105);
or U14236 (N_14236,N_13907,N_13597);
and U14237 (N_14237,N_12741,N_13481);
nor U14238 (N_14238,N_13708,N_12683);
nor U14239 (N_14239,N_13448,N_13313);
or U14240 (N_14240,N_13859,N_13260);
and U14241 (N_14241,N_13263,N_13157);
nor U14242 (N_14242,N_13500,N_13045);
and U14243 (N_14243,N_12409,N_12053);
xnor U14244 (N_14244,N_12522,N_12924);
nor U14245 (N_14245,N_12681,N_13465);
nand U14246 (N_14246,N_12543,N_13075);
nor U14247 (N_14247,N_13028,N_13036);
and U14248 (N_14248,N_12909,N_13016);
xor U14249 (N_14249,N_12200,N_12233);
nor U14250 (N_14250,N_13292,N_13892);
and U14251 (N_14251,N_13417,N_12260);
xor U14252 (N_14252,N_12209,N_12002);
xor U14253 (N_14253,N_13428,N_12202);
nor U14254 (N_14254,N_13946,N_13384);
xor U14255 (N_14255,N_12628,N_12406);
xor U14256 (N_14256,N_13071,N_13592);
nand U14257 (N_14257,N_12065,N_13608);
nor U14258 (N_14258,N_13798,N_12622);
or U14259 (N_14259,N_13891,N_12237);
nand U14260 (N_14260,N_13662,N_12659);
nand U14261 (N_14261,N_13690,N_13300);
or U14262 (N_14262,N_13239,N_12846);
nor U14263 (N_14263,N_12142,N_12262);
xor U14264 (N_14264,N_12826,N_12557);
nor U14265 (N_14265,N_12348,N_13262);
nand U14266 (N_14266,N_12183,N_12756);
xnor U14267 (N_14267,N_13761,N_12930);
nor U14268 (N_14268,N_12166,N_12934);
nor U14269 (N_14269,N_12853,N_13397);
and U14270 (N_14270,N_13571,N_13392);
nor U14271 (N_14271,N_12696,N_13643);
and U14272 (N_14272,N_12624,N_13585);
and U14273 (N_14273,N_12017,N_13731);
nand U14274 (N_14274,N_13210,N_13546);
nand U14275 (N_14275,N_12542,N_12353);
and U14276 (N_14276,N_13387,N_13301);
or U14277 (N_14277,N_13363,N_13792);
and U14278 (N_14278,N_13612,N_12844);
or U14279 (N_14279,N_12238,N_13928);
nand U14280 (N_14280,N_13730,N_12377);
nor U14281 (N_14281,N_13540,N_12438);
nand U14282 (N_14282,N_12787,N_13459);
nand U14283 (N_14283,N_13205,N_13484);
nor U14284 (N_14284,N_12046,N_12318);
nor U14285 (N_14285,N_12380,N_12946);
and U14286 (N_14286,N_13519,N_12639);
or U14287 (N_14287,N_13306,N_12737);
nor U14288 (N_14288,N_13861,N_13406);
or U14289 (N_14289,N_12366,N_12974);
nand U14290 (N_14290,N_13099,N_12698);
xor U14291 (N_14291,N_13930,N_13811);
nand U14292 (N_14292,N_13091,N_12308);
nand U14293 (N_14293,N_13220,N_13784);
or U14294 (N_14294,N_13544,N_13093);
nor U14295 (N_14295,N_12664,N_13775);
or U14296 (N_14296,N_13143,N_12286);
nor U14297 (N_14297,N_13159,N_12691);
and U14298 (N_14298,N_13280,N_12718);
and U14299 (N_14299,N_13009,N_13131);
nor U14300 (N_14300,N_12048,N_13436);
xnor U14301 (N_14301,N_12800,N_12379);
or U14302 (N_14302,N_12026,N_13921);
nand U14303 (N_14303,N_13160,N_13162);
xnor U14304 (N_14304,N_13812,N_12188);
and U14305 (N_14305,N_12500,N_13734);
and U14306 (N_14306,N_12914,N_12580);
and U14307 (N_14307,N_12791,N_12501);
and U14308 (N_14308,N_13641,N_12059);
and U14309 (N_14309,N_12030,N_13083);
nor U14310 (N_14310,N_13748,N_13750);
nand U14311 (N_14311,N_13429,N_13094);
nand U14312 (N_14312,N_13772,N_13827);
nand U14313 (N_14313,N_13342,N_13654);
nand U14314 (N_14314,N_12938,N_12254);
nor U14315 (N_14315,N_13414,N_12705);
and U14316 (N_14316,N_12774,N_13856);
and U14317 (N_14317,N_12149,N_13227);
or U14318 (N_14318,N_13343,N_12942);
nand U14319 (N_14319,N_13805,N_13114);
or U14320 (N_14320,N_13126,N_12679);
and U14321 (N_14321,N_12967,N_12568);
and U14322 (N_14322,N_13097,N_13982);
or U14323 (N_14323,N_12040,N_12728);
nand U14324 (N_14324,N_12650,N_12923);
and U14325 (N_14325,N_12205,N_13587);
or U14326 (N_14326,N_12481,N_12236);
nor U14327 (N_14327,N_12426,N_13834);
nor U14328 (N_14328,N_13739,N_12213);
nand U14329 (N_14329,N_12732,N_13305);
nor U14330 (N_14330,N_12847,N_13178);
and U14331 (N_14331,N_13796,N_13130);
and U14332 (N_14332,N_12141,N_12773);
nor U14333 (N_14333,N_13413,N_12802);
and U14334 (N_14334,N_13275,N_13041);
nor U14335 (N_14335,N_13839,N_13846);
nand U14336 (N_14336,N_13505,N_13074);
nor U14337 (N_14337,N_12476,N_12668);
nor U14338 (N_14338,N_12133,N_13737);
nand U14339 (N_14339,N_12098,N_13539);
nand U14340 (N_14340,N_13926,N_13024);
nand U14341 (N_14341,N_13766,N_12170);
nand U14342 (N_14342,N_13115,N_12587);
nor U14343 (N_14343,N_13025,N_12520);
and U14344 (N_14344,N_13997,N_12225);
nor U14345 (N_14345,N_13628,N_13017);
or U14346 (N_14346,N_13646,N_13169);
nor U14347 (N_14347,N_13254,N_12895);
nor U14348 (N_14348,N_12648,N_13583);
nor U14349 (N_14349,N_13147,N_12825);
and U14350 (N_14350,N_13964,N_12611);
nor U14351 (N_14351,N_13532,N_12110);
or U14352 (N_14352,N_12361,N_13870);
and U14353 (N_14353,N_13556,N_12099);
and U14354 (N_14354,N_12185,N_13970);
or U14355 (N_14355,N_13370,N_12337);
nor U14356 (N_14356,N_13745,N_13499);
and U14357 (N_14357,N_13095,N_13218);
and U14358 (N_14358,N_13046,N_13381);
or U14359 (N_14359,N_13441,N_12798);
xor U14360 (N_14360,N_13426,N_13146);
and U14361 (N_14361,N_13657,N_12843);
or U14362 (N_14362,N_13988,N_13578);
nor U14363 (N_14363,N_13848,N_13439);
xnor U14364 (N_14364,N_12569,N_13862);
nor U14365 (N_14365,N_12333,N_13797);
and U14366 (N_14366,N_13890,N_12669);
xor U14367 (N_14367,N_12165,N_13825);
or U14368 (N_14368,N_13005,N_13242);
nor U14369 (N_14369,N_12603,N_12606);
or U14370 (N_14370,N_12090,N_12952);
and U14371 (N_14371,N_13362,N_13336);
and U14372 (N_14372,N_13246,N_13341);
nor U14373 (N_14373,N_13650,N_13230);
nand U14374 (N_14374,N_13823,N_13371);
and U14375 (N_14375,N_13631,N_12109);
and U14376 (N_14376,N_13153,N_13108);
or U14377 (N_14377,N_13380,N_13132);
nor U14378 (N_14378,N_13331,N_12857);
or U14379 (N_14379,N_12539,N_13888);
nand U14380 (N_14380,N_12086,N_13503);
nand U14381 (N_14381,N_13118,N_13357);
nand U14382 (N_14382,N_12063,N_13356);
nand U14383 (N_14383,N_13525,N_13435);
or U14384 (N_14384,N_13444,N_13089);
and U14385 (N_14385,N_12304,N_12273);
nor U14386 (N_14386,N_12124,N_12781);
and U14387 (N_14387,N_12355,N_13015);
nor U14388 (N_14388,N_12755,N_12884);
nand U14389 (N_14389,N_12632,N_13740);
xor U14390 (N_14390,N_12473,N_12287);
nor U14391 (N_14391,N_13785,N_13279);
nand U14392 (N_14392,N_12903,N_13010);
or U14393 (N_14393,N_12761,N_13316);
nand U14394 (N_14394,N_13070,N_13329);
and U14395 (N_14395,N_12745,N_13667);
nand U14396 (N_14396,N_12338,N_13768);
nand U14397 (N_14397,N_12060,N_13138);
or U14398 (N_14398,N_13137,N_12401);
and U14399 (N_14399,N_13776,N_12370);
or U14400 (N_14400,N_13591,N_13471);
or U14401 (N_14401,N_12809,N_12328);
or U14402 (N_14402,N_13127,N_13758);
and U14403 (N_14403,N_13425,N_12711);
and U14404 (N_14404,N_13610,N_12342);
and U14405 (N_14405,N_12101,N_12631);
and U14406 (N_14406,N_13950,N_13037);
nor U14407 (N_14407,N_13272,N_13291);
and U14408 (N_14408,N_12784,N_12321);
nand U14409 (N_14409,N_13158,N_13403);
and U14410 (N_14410,N_12039,N_13151);
nand U14411 (N_14411,N_12740,N_13932);
and U14412 (N_14412,N_13207,N_13454);
or U14413 (N_14413,N_13468,N_12009);
nand U14414 (N_14414,N_12119,N_12001);
and U14415 (N_14415,N_13473,N_12117);
nor U14416 (N_14416,N_12194,N_12955);
and U14417 (N_14417,N_13635,N_12140);
nor U14418 (N_14418,N_13903,N_12392);
nor U14419 (N_14419,N_12497,N_13142);
nand U14420 (N_14420,N_13322,N_12232);
and U14421 (N_14421,N_13284,N_13389);
or U14422 (N_14422,N_13112,N_12913);
nand U14423 (N_14423,N_13082,N_12758);
nand U14424 (N_14424,N_13461,N_13298);
nor U14425 (N_14425,N_13976,N_12978);
and U14426 (N_14426,N_12764,N_12332);
nor U14427 (N_14427,N_13312,N_12627);
or U14428 (N_14428,N_13023,N_13039);
or U14429 (N_14429,N_13106,N_12116);
nor U14430 (N_14430,N_13479,N_12212);
xor U14431 (N_14431,N_13843,N_12179);
and U14432 (N_14432,N_13437,N_13164);
nor U14433 (N_14433,N_13535,N_13018);
or U14434 (N_14434,N_12464,N_13744);
xnor U14435 (N_14435,N_12074,N_13445);
and U14436 (N_14436,N_13121,N_13195);
or U14437 (N_14437,N_13765,N_12712);
nor U14438 (N_14438,N_13658,N_12818);
or U14439 (N_14439,N_12605,N_13974);
xnor U14440 (N_14440,N_13508,N_13875);
nor U14441 (N_14441,N_12028,N_12103);
and U14442 (N_14442,N_13779,N_12778);
nand U14443 (N_14443,N_12067,N_13354);
and U14444 (N_14444,N_12310,N_12451);
xnor U14445 (N_14445,N_13967,N_12162);
nand U14446 (N_14446,N_12962,N_12176);
xnor U14447 (N_14447,N_13824,N_12257);
and U14448 (N_14448,N_13482,N_13237);
nand U14449 (N_14449,N_12858,N_12840);
and U14450 (N_14450,N_12638,N_12667);
nor U14451 (N_14451,N_12931,N_13486);
or U14452 (N_14452,N_12970,N_12437);
or U14453 (N_14453,N_13412,N_13211);
nor U14454 (N_14454,N_12837,N_13661);
nor U14455 (N_14455,N_13111,N_13219);
nand U14456 (N_14456,N_13317,N_12192);
xnor U14457 (N_14457,N_12495,N_13491);
nand U14458 (N_14458,N_13268,N_13782);
xor U14459 (N_14459,N_12207,N_12869);
or U14460 (N_14460,N_13520,N_12111);
xnor U14461 (N_14461,N_13116,N_12436);
nand U14462 (N_14462,N_12269,N_12665);
nand U14463 (N_14463,N_12504,N_13198);
nor U14464 (N_14464,N_12657,N_13199);
nor U14465 (N_14465,N_12359,N_12567);
and U14466 (N_14466,N_12594,N_13558);
and U14467 (N_14467,N_13914,N_13702);
nand U14468 (N_14468,N_13086,N_12384);
nand U14469 (N_14469,N_12523,N_13987);
nand U14470 (N_14470,N_12073,N_13339);
and U14471 (N_14471,N_12289,N_13192);
and U14472 (N_14472,N_13732,N_13202);
or U14473 (N_14473,N_12315,N_13989);
xnor U14474 (N_14474,N_12450,N_13458);
nor U14475 (N_14475,N_12794,N_12694);
nor U14476 (N_14476,N_12172,N_13844);
nor U14477 (N_14477,N_13882,N_13972);
and U14478 (N_14478,N_13423,N_12033);
nor U14479 (N_14479,N_12529,N_12919);
nor U14480 (N_14480,N_13424,N_13623);
nand U14481 (N_14481,N_12126,N_13073);
or U14482 (N_14482,N_12995,N_13637);
nor U14483 (N_14483,N_13200,N_13058);
nand U14484 (N_14484,N_13617,N_12720);
xnor U14485 (N_14485,N_13936,N_12078);
nand U14486 (N_14486,N_13125,N_12277);
or U14487 (N_14487,N_12908,N_13369);
nor U14488 (N_14488,N_12973,N_12449);
nand U14489 (N_14489,N_12121,N_12713);
nand U14490 (N_14490,N_13850,N_12612);
nand U14491 (N_14491,N_13531,N_13986);
or U14492 (N_14492,N_13203,N_13047);
or U14493 (N_14493,N_12584,N_13820);
nor U14494 (N_14494,N_12035,N_13551);
or U14495 (N_14495,N_13286,N_13854);
or U14496 (N_14496,N_12219,N_12107);
nor U14497 (N_14497,N_13572,N_12259);
xnor U14498 (N_14498,N_13450,N_12331);
or U14499 (N_14499,N_13420,N_13385);
or U14500 (N_14500,N_13443,N_12134);
or U14501 (N_14501,N_12356,N_13806);
or U14502 (N_14502,N_13840,N_13814);
nor U14503 (N_14503,N_13809,N_13944);
xor U14504 (N_14504,N_12526,N_12593);
or U14505 (N_14505,N_12790,N_13524);
nor U14506 (N_14506,N_12485,N_13368);
nand U14507 (N_14507,N_12572,N_12037);
and U14508 (N_14508,N_12399,N_13594);
nor U14509 (N_14509,N_12968,N_12836);
nor U14510 (N_14510,N_12987,N_13774);
or U14511 (N_14511,N_12983,N_13438);
nor U14512 (N_14512,N_12255,N_12197);
or U14513 (N_14513,N_13885,N_12599);
nand U14514 (N_14514,N_12695,N_12990);
xor U14515 (N_14515,N_13853,N_13794);
nor U14516 (N_14516,N_12850,N_12102);
or U14517 (N_14517,N_12564,N_12034);
and U14518 (N_14518,N_12834,N_12295);
nor U14519 (N_14519,N_12267,N_12015);
xor U14520 (N_14520,N_12145,N_13510);
or U14521 (N_14521,N_12731,N_12680);
and U14522 (N_14522,N_12582,N_13133);
or U14523 (N_14523,N_12199,N_12643);
xnor U14524 (N_14524,N_13061,N_13102);
nor U14525 (N_14525,N_12391,N_12407);
xnor U14526 (N_14526,N_13400,N_12877);
nand U14527 (N_14527,N_12841,N_12831);
and U14528 (N_14528,N_12953,N_12852);
nor U14529 (N_14529,N_12108,N_12799);
or U14530 (N_14530,N_12459,N_13985);
xnor U14531 (N_14531,N_12748,N_12151);
or U14532 (N_14532,N_12419,N_13879);
and U14533 (N_14533,N_12014,N_12309);
xnor U14534 (N_14534,N_12229,N_13935);
nor U14535 (N_14535,N_12226,N_13096);
or U14536 (N_14536,N_12949,N_12068);
or U14537 (N_14537,N_13900,N_13815);
xnor U14538 (N_14538,N_12352,N_12729);
nor U14539 (N_14539,N_12656,N_13656);
and U14540 (N_14540,N_12905,N_12566);
and U14541 (N_14541,N_13876,N_13826);
and U14542 (N_14542,N_13485,N_13931);
nor U14543 (N_14543,N_12480,N_13918);
or U14544 (N_14544,N_13577,N_13893);
xor U14545 (N_14545,N_12856,N_13538);
nor U14546 (N_14546,N_12448,N_13326);
and U14547 (N_14547,N_12330,N_12410);
nor U14548 (N_14548,N_13866,N_13649);
xor U14549 (N_14549,N_12386,N_13706);
and U14550 (N_14550,N_13590,N_13804);
nor U14551 (N_14551,N_12491,N_13303);
or U14552 (N_14552,N_13501,N_12692);
and U14553 (N_14553,N_13287,N_13733);
xnor U14554 (N_14554,N_12936,N_13992);
and U14555 (N_14555,N_12418,N_12235);
nor U14556 (N_14556,N_12805,N_12563);
and U14557 (N_14557,N_12928,N_12064);
and U14558 (N_14558,N_12243,N_12757);
and U14559 (N_14559,N_12498,N_13257);
nor U14560 (N_14560,N_12156,N_13050);
nor U14561 (N_14561,N_13955,N_12463);
and U14562 (N_14562,N_12975,N_13048);
nor U14563 (N_14563,N_12918,N_13372);
or U14564 (N_14564,N_12835,N_12447);
nand U14565 (N_14565,N_12854,N_13721);
xor U14566 (N_14566,N_13390,N_13692);
nand U14567 (N_14567,N_13489,N_12394);
nor U14568 (N_14568,N_13564,N_12685);
and U14569 (N_14569,N_13148,N_12771);
or U14570 (N_14570,N_13736,N_12057);
or U14571 (N_14571,N_13897,N_12038);
nor U14572 (N_14572,N_13358,N_12088);
or U14573 (N_14573,N_12754,N_12306);
nor U14574 (N_14574,N_12661,N_13249);
nor U14575 (N_14575,N_13281,N_12417);
nor U14576 (N_14576,N_13659,N_12623);
xnor U14577 (N_14577,N_12054,N_13920);
and U14578 (N_14578,N_13753,N_12341);
and U14579 (N_14579,N_12335,N_12900);
and U14580 (N_14580,N_13881,N_13880);
and U14581 (N_14581,N_12440,N_12245);
nand U14582 (N_14582,N_12360,N_12788);
and U14583 (N_14583,N_13090,N_12921);
or U14584 (N_14584,N_12693,N_12112);
and U14585 (N_14585,N_13035,N_13672);
nand U14586 (N_14586,N_13399,N_13173);
or U14587 (N_14587,N_12275,N_12313);
or U14588 (N_14588,N_13255,N_12496);
nor U14589 (N_14589,N_13375,N_12532);
nor U14590 (N_14590,N_12829,N_13681);
or U14591 (N_14591,N_13470,N_12618);
and U14592 (N_14592,N_13278,N_13507);
nor U14593 (N_14593,N_13927,N_12722);
nand U14594 (N_14594,N_13344,N_13081);
and U14595 (N_14595,N_13128,N_12100);
and U14596 (N_14596,N_12159,N_12954);
nand U14597 (N_14597,N_13614,N_12029);
and U14598 (N_14598,N_12902,N_13144);
nor U14599 (N_14599,N_13062,N_12678);
and U14600 (N_14600,N_12795,N_12960);
and U14601 (N_14601,N_12780,N_12456);
and U14602 (N_14602,N_13738,N_12891);
nor U14603 (N_14603,N_13634,N_12519);
or U14604 (N_14604,N_13110,N_13321);
and U14605 (N_14605,N_13059,N_12833);
or U14606 (N_14606,N_13502,N_13533);
xor U14607 (N_14607,N_13100,N_12963);
nand U14608 (N_14608,N_13609,N_13451);
nand U14609 (N_14609,N_13022,N_13174);
nor U14610 (N_14610,N_13064,N_12702);
xor U14611 (N_14611,N_12024,N_12256);
or U14612 (N_14612,N_13225,N_12346);
nand U14613 (N_14613,N_13925,N_12494);
and U14614 (N_14614,N_13729,N_13245);
nor U14615 (N_14615,N_12562,N_13163);
and U14616 (N_14616,N_12855,N_13945);
and U14617 (N_14617,N_12489,N_12874);
and U14618 (N_14618,N_12230,N_12511);
nor U14619 (N_14619,N_13325,N_13957);
and U14620 (N_14620,N_13008,N_12556);
nand U14621 (N_14621,N_12487,N_12893);
or U14622 (N_14622,N_13409,N_12052);
nor U14623 (N_14623,N_13251,N_12431);
and U14624 (N_14624,N_12296,N_13884);
and U14625 (N_14625,N_12999,N_12429);
or U14626 (N_14626,N_12292,N_12146);
nand U14627 (N_14627,N_12976,N_13003);
nor U14628 (N_14628,N_12637,N_12832);
nand U14629 (N_14629,N_12537,N_12969);
nand U14630 (N_14630,N_13688,N_13004);
or U14631 (N_14631,N_13596,N_12966);
and U14632 (N_14632,N_13780,N_12076);
or U14633 (N_14633,N_13049,N_12044);
and U14634 (N_14634,N_13781,N_12455);
xnor U14635 (N_14635,N_13741,N_12404);
nor U14636 (N_14636,N_13446,N_12139);
or U14637 (N_14637,N_12191,N_12576);
nand U14638 (N_14638,N_12433,N_12435);
nor U14639 (N_14639,N_13477,N_13786);
or U14640 (N_14640,N_12719,N_12904);
nor U14641 (N_14641,N_12574,N_12776);
and U14642 (N_14642,N_13366,N_13652);
nor U14643 (N_14643,N_12423,N_13570);
and U14644 (N_14644,N_13209,N_13767);
and U14645 (N_14645,N_13185,N_13705);
nor U14646 (N_14646,N_12839,N_13788);
or U14647 (N_14647,N_12578,N_13562);
nor U14648 (N_14648,N_13052,N_12239);
nor U14649 (N_14649,N_13723,N_12189);
and U14650 (N_14650,N_13069,N_13092);
xnor U14651 (N_14651,N_12083,N_13763);
or U14652 (N_14652,N_13087,N_12959);
nand U14653 (N_14653,N_13581,N_13290);
xnor U14654 (N_14654,N_12400,N_13318);
or U14655 (N_14655,N_13595,N_13333);
nand U14656 (N_14656,N_13855,N_12927);
or U14657 (N_14657,N_13407,N_12467);
or U14658 (N_14658,N_13416,N_12319);
or U14659 (N_14659,N_13323,N_12626);
or U14660 (N_14660,N_12354,N_13980);
nor U14661 (N_14661,N_12708,N_12175);
and U14662 (N_14662,N_12446,N_13940);
or U14663 (N_14663,N_13867,N_13751);
nand U14664 (N_14664,N_13961,N_13042);
and U14665 (N_14665,N_12471,N_12677);
xnor U14666 (N_14666,N_13347,N_12195);
and U14667 (N_14667,N_12767,N_13434);
or U14668 (N_14668,N_13167,N_12130);
and U14669 (N_14669,N_12475,N_12276);
nand U14670 (N_14670,N_12686,N_13943);
nand U14671 (N_14671,N_13462,N_13601);
xor U14672 (N_14672,N_13703,N_12390);
nand U14673 (N_14673,N_13995,N_12760);
xor U14674 (N_14674,N_13274,N_12982);
xor U14675 (N_14675,N_13011,N_12744);
nand U14676 (N_14676,N_12581,N_13516);
or U14677 (N_14677,N_13902,N_13722);
nor U14678 (N_14678,N_12244,N_13085);
or U14679 (N_14679,N_13611,N_13449);
or U14680 (N_14680,N_12775,N_13373);
xnor U14681 (N_14681,N_13332,N_13668);
or U14682 (N_14682,N_13576,N_12772);
or U14683 (N_14683,N_13457,N_12881);
nand U14684 (N_14684,N_12838,N_12300);
or U14685 (N_14685,N_13579,N_12128);
or U14686 (N_14686,N_12546,N_12806);
and U14687 (N_14687,N_13978,N_13020);
nor U14688 (N_14688,N_12889,N_13233);
nor U14689 (N_14689,N_12345,N_12062);
or U14690 (N_14690,N_12153,N_12510);
nand U14691 (N_14691,N_12092,N_12413);
nor U14692 (N_14692,N_13243,N_13983);
or U14693 (N_14693,N_13716,N_13172);
or U14694 (N_14694,N_12885,N_12684);
nand U14695 (N_14695,N_13743,N_13749);
nor U14696 (N_14696,N_12882,N_12617);
nor U14697 (N_14697,N_13283,N_12374);
or U14698 (N_14698,N_12131,N_13488);
nor U14699 (N_14699,N_12081,N_12482);
nand U14700 (N_14700,N_13056,N_12241);
or U14701 (N_14701,N_12849,N_13919);
nor U14702 (N_14702,N_12114,N_13953);
and U14703 (N_14703,N_12743,N_12508);
nand U14704 (N_14704,N_12704,N_13474);
nor U14705 (N_14705,N_13939,N_13836);
nor U14706 (N_14706,N_13136,N_13523);
or U14707 (N_14707,N_12279,N_12948);
nand U14708 (N_14708,N_12503,N_12892);
or U14709 (N_14709,N_13029,N_13012);
nand U14710 (N_14710,N_13647,N_12071);
or U14711 (N_14711,N_12320,N_12807);
nor U14712 (N_14712,N_13841,N_13244);
nand U14713 (N_14713,N_12204,N_12042);
xnor U14714 (N_14714,N_13807,N_13883);
nor U14715 (N_14715,N_13013,N_12368);
and U14716 (N_14716,N_13757,N_12803);
nand U14717 (N_14717,N_12305,N_13166);
or U14718 (N_14718,N_12163,N_12896);
nor U14719 (N_14719,N_12270,N_13273);
nand U14720 (N_14720,N_13065,N_12935);
nor U14721 (N_14721,N_12992,N_13638);
or U14722 (N_14722,N_13746,N_12217);
or U14723 (N_14723,N_13694,N_12768);
nor U14724 (N_14724,N_13712,N_12004);
nand U14725 (N_14725,N_13606,N_12597);
nand U14726 (N_14726,N_13984,N_12079);
and U14727 (N_14727,N_12883,N_12640);
xor U14728 (N_14728,N_13271,N_13648);
or U14729 (N_14729,N_13568,N_12717);
nand U14730 (N_14730,N_13633,N_13831);
nand U14731 (N_14731,N_13304,N_13288);
nor U14732 (N_14732,N_13711,N_13849);
nand U14733 (N_14733,N_13835,N_12701);
nor U14734 (N_14734,N_12178,N_12734);
xor U14735 (N_14735,N_12898,N_12376);
or U14736 (N_14736,N_12322,N_12545);
or U14737 (N_14737,N_13665,N_13602);
and U14738 (N_14738,N_13253,N_12268);
and U14739 (N_14739,N_13963,N_12560);
nor U14740 (N_14740,N_12682,N_12157);
and U14741 (N_14741,N_12876,N_13145);
and U14742 (N_14742,N_12445,N_13549);
nand U14743 (N_14743,N_12544,N_13221);
nand U14744 (N_14744,N_12789,N_12828);
xnor U14745 (N_14745,N_13700,N_12408);
or U14746 (N_14746,N_12263,N_12879);
and U14747 (N_14747,N_12218,N_13348);
or U14748 (N_14748,N_13857,N_12887);
or U14749 (N_14749,N_13969,N_12706);
and U14750 (N_14750,N_13771,N_13238);
nor U14751 (N_14751,N_12821,N_13644);
and U14752 (N_14752,N_13695,N_13911);
xor U14753 (N_14753,N_13728,N_13625);
xnor U14754 (N_14754,N_12642,N_12742);
or U14755 (N_14755,N_13548,N_13386);
nand U14756 (N_14756,N_12484,N_13171);
nand U14757 (N_14757,N_13863,N_13725);
nor U14758 (N_14758,N_13212,N_12608);
nor U14759 (N_14759,N_12733,N_13492);
or U14760 (N_14760,N_12763,N_13034);
and U14761 (N_14761,N_13630,N_12649);
or U14762 (N_14762,N_13593,N_12383);
nand U14763 (N_14763,N_12980,N_12339);
nor U14764 (N_14764,N_13497,N_12541);
or U14765 (N_14765,N_12736,N_13673);
or U14766 (N_14766,N_12298,N_13639);
or U14767 (N_14767,N_13618,N_13324);
nor U14768 (N_14768,N_12796,N_13469);
xor U14769 (N_14769,N_12367,N_13213);
nor U14770 (N_14770,N_13642,N_13315);
nor U14771 (N_14771,N_12782,N_12006);
nand U14772 (N_14772,N_12610,N_13427);
nand U14773 (N_14773,N_12851,N_12861);
nor U14774 (N_14774,N_13084,N_13453);
nor U14775 (N_14775,N_12478,N_13949);
and U14776 (N_14776,N_12573,N_12670);
nor U14777 (N_14777,N_12122,N_13476);
or U14778 (N_14778,N_13007,N_12412);
or U14779 (N_14779,N_12129,N_13006);
nand U14780 (N_14780,N_13204,N_13627);
or U14781 (N_14781,N_13718,N_12075);
or U14782 (N_14782,N_13103,N_13388);
and U14783 (N_14783,N_13589,N_12016);
or U14784 (N_14784,N_12867,N_13604);
and U14785 (N_14785,N_12274,N_12240);
or U14786 (N_14786,N_12674,N_12442);
and U14787 (N_14787,N_13229,N_12819);
and U14788 (N_14788,N_13129,N_13707);
nor U14789 (N_14789,N_13910,N_12687);
or U14790 (N_14790,N_13193,N_12890);
xor U14791 (N_14791,N_13183,N_12517);
and U14792 (N_14792,N_13250,N_13521);
or U14793 (N_14793,N_13440,N_13308);
nand U14794 (N_14794,N_12385,N_12730);
nand U14795 (N_14795,N_12937,N_13990);
or U14796 (N_14796,N_13689,N_12011);
and U14797 (N_14797,N_12222,N_12926);
nand U14798 (N_14798,N_12281,N_12929);
nand U14799 (N_14799,N_13801,N_12598);
nand U14800 (N_14800,N_12144,N_13394);
xor U14801 (N_14801,N_13629,N_12452);
nor U14802 (N_14802,N_12738,N_13669);
and U14803 (N_14803,N_12823,N_12549);
nor U14804 (N_14804,N_12272,N_13526);
nor U14805 (N_14805,N_12021,N_13452);
and U14806 (N_14806,N_12621,N_12093);
nor U14807 (N_14807,N_12486,N_12000);
xor U14808 (N_14808,N_12944,N_13600);
nor U14809 (N_14809,N_13498,N_12910);
nand U14810 (N_14810,N_12842,N_13364);
or U14811 (N_14811,N_12591,N_13687);
nand U14812 (N_14812,N_13566,N_12671);
nor U14813 (N_14813,N_12427,N_13351);
nor U14814 (N_14814,N_13383,N_12462);
or U14815 (N_14815,N_13256,N_13979);
nor U14816 (N_14816,N_13621,N_12561);
nor U14817 (N_14817,N_12220,N_12988);
or U14818 (N_14818,N_12688,N_12492);
and U14819 (N_14819,N_12043,N_12137);
nor U14820 (N_14820,N_12507,N_12018);
nand U14821 (N_14821,N_12072,N_13971);
and U14822 (N_14822,N_12173,N_12184);
or U14823 (N_14823,N_12211,N_13190);
xnor U14824 (N_14824,N_12965,N_13226);
nor U14825 (N_14825,N_13860,N_12362);
nand U14826 (N_14826,N_12700,N_13810);
and U14827 (N_14827,N_13803,N_13693);
nor U14828 (N_14828,N_12493,N_12940);
and U14829 (N_14829,N_13330,N_12317);
nand U14830 (N_14830,N_13773,N_12553);
and U14831 (N_14831,N_13509,N_13819);
xnor U14832 (N_14832,N_13616,N_12174);
nand U14833 (N_14833,N_12993,N_12003);
xnor U14834 (N_14834,N_13573,N_12249);
xor U14835 (N_14835,N_13800,N_13460);
nor U14836 (N_14836,N_13906,N_13769);
nor U14837 (N_14837,N_13615,N_12007);
and U14838 (N_14838,N_12414,N_13104);
and U14839 (N_14839,N_13140,N_13422);
nand U14840 (N_14840,N_12288,N_13567);
or U14841 (N_14841,N_13349,N_12998);
and U14842 (N_14842,N_12432,N_13537);
or U14843 (N_14843,N_12152,N_12525);
nand U14844 (N_14844,N_13374,N_12801);
or U14845 (N_14845,N_12132,N_13704);
nor U14846 (N_14846,N_13534,N_13170);
nor U14847 (N_14847,N_12231,N_12224);
nand U14848 (N_14848,N_12947,N_13808);
or U14849 (N_14849,N_12552,N_12297);
nand U14850 (N_14850,N_12759,N_12120);
and U14851 (N_14851,N_12334,N_12515);
nor U14852 (N_14852,N_12089,N_13442);
or U14853 (N_14853,N_13560,N_13014);
nor U14854 (N_14854,N_13161,N_13563);
nor U14855 (N_14855,N_13231,N_12161);
nor U14856 (N_14856,N_12454,N_12477);
or U14857 (N_14857,N_12115,N_13530);
nand U14858 (N_14858,N_13353,N_12148);
nand U14859 (N_14859,N_12171,N_13764);
or U14860 (N_14860,N_12866,N_13937);
xor U14861 (N_14861,N_12550,N_12405);
xor U14862 (N_14862,N_12032,N_13393);
or U14863 (N_14863,N_13165,N_13247);
and U14864 (N_14864,N_12658,N_13224);
nand U14865 (N_14865,N_12540,N_12715);
nand U14866 (N_14866,N_12393,N_12187);
nor U14867 (N_14867,N_12820,N_12945);
nor U14868 (N_14868,N_13187,N_12964);
nand U14869 (N_14869,N_12460,N_12996);
xor U14870 (N_14870,N_12814,N_13655);
nand U14871 (N_14871,N_13701,N_12548);
nor U14872 (N_14872,N_12301,N_12956);
nor U14873 (N_14873,N_12326,N_12347);
and U14874 (N_14874,N_12933,N_12920);
and U14875 (N_14875,N_12351,N_13889);
nand U14876 (N_14876,N_12323,N_13495);
or U14877 (N_14877,N_12635,N_13588);
nor U14878 (N_14878,N_12136,N_12646);
and U14879 (N_14879,N_12812,N_13991);
nand U14880 (N_14880,N_12609,N_13828);
or U14881 (N_14881,N_12735,N_12911);
nand U14882 (N_14882,N_12792,N_12291);
and U14883 (N_14883,N_12943,N_12469);
nand U14884 (N_14884,N_12396,N_12135);
nand U14885 (N_14885,N_12293,N_13515);
nand U14886 (N_14886,N_12697,N_12307);
or U14887 (N_14887,N_13896,N_12721);
or U14888 (N_14888,N_13135,N_13550);
nand U14889 (N_14889,N_12087,N_13487);
and U14890 (N_14890,N_12094,N_12104);
and U14891 (N_14891,N_13998,N_12138);
nand U14892 (N_14892,N_13475,N_13938);
nand U14893 (N_14893,N_13404,N_12505);
or U14894 (N_14894,N_12662,N_12258);
and U14895 (N_14895,N_13182,N_12762);
and U14896 (N_14896,N_13410,N_13194);
or U14897 (N_14897,N_12644,N_12378);
nand U14898 (N_14898,N_12595,N_12411);
nor U14899 (N_14899,N_12811,N_12868);
nor U14900 (N_14900,N_12633,N_12625);
nand U14901 (N_14901,N_13886,N_13345);
nor U14902 (N_14902,N_13724,N_13277);
nand U14903 (N_14903,N_13367,N_12461);
nor U14904 (N_14904,N_13264,N_13679);
or U14905 (N_14905,N_12190,N_12710);
or U14906 (N_14906,N_12490,N_13235);
and U14907 (N_14907,N_13996,N_12358);
and U14908 (N_14908,N_12387,N_13494);
or U14909 (N_14909,N_12577,N_13813);
or U14910 (N_14910,N_13759,N_13232);
nor U14911 (N_14911,N_12726,N_12516);
and U14912 (N_14912,N_13334,N_12645);
nor U14913 (N_14913,N_12261,N_13456);
nand U14914 (N_14914,N_13189,N_13575);
nand U14915 (N_14915,N_12155,N_12483);
nor U14916 (N_14916,N_12725,N_12630);
nand U14917 (N_14917,N_13793,N_13580);
xnor U14918 (N_14918,N_12430,N_12439);
or U14919 (N_14919,N_13818,N_12265);
or U14920 (N_14920,N_13789,N_12513);
nand U14921 (N_14921,N_12512,N_12113);
and U14922 (N_14922,N_12458,N_12168);
xnor U14923 (N_14923,N_12536,N_12357);
and U14924 (N_14924,N_13122,N_13574);
nor U14925 (N_14925,N_12971,N_12629);
nand U14926 (N_14926,N_13293,N_13030);
nand U14927 (N_14927,N_12727,N_13872);
nor U14928 (N_14928,N_12056,N_12604);
nand U14929 (N_14929,N_13670,N_12312);
nor U14930 (N_14930,N_12201,N_13909);
or U14931 (N_14931,N_12585,N_13952);
or U14932 (N_14932,N_12206,N_12586);
or U14933 (N_14933,N_12672,N_12765);
nor U14934 (N_14934,N_13319,N_12916);
nor U14935 (N_14935,N_13514,N_12311);
or U14936 (N_14936,N_13685,N_12571);
or U14937 (N_14937,N_12246,N_12395);
nor U14938 (N_14938,N_13683,N_12590);
nor U14939 (N_14939,N_12528,N_13713);
nor U14940 (N_14940,N_13513,N_12845);
or U14941 (N_14941,N_12282,N_12466);
and U14942 (N_14942,N_12531,N_12749);
and U14943 (N_14943,N_12939,N_12620);
and U14944 (N_14944,N_13877,N_13553);
nand U14945 (N_14945,N_13735,N_13845);
and U14946 (N_14946,N_13309,N_13141);
and U14947 (N_14947,N_12082,N_12050);
or U14948 (N_14948,N_13455,N_13430);
nand U14949 (N_14949,N_12579,N_13296);
or U14950 (N_14950,N_13677,N_13726);
xnor U14951 (N_14951,N_12371,N_13959);
or U14952 (N_14952,N_13197,N_13968);
nand U14953 (N_14953,N_12922,N_12424);
xor U14954 (N_14954,N_13411,N_13760);
nor U14955 (N_14955,N_12284,N_13139);
nor U14956 (N_14956,N_13727,N_12977);
nand U14957 (N_14957,N_12786,N_12316);
nand U14958 (N_14958,N_12641,N_12143);
nand U14959 (N_14959,N_12808,N_12402);
nand U14960 (N_14960,N_12558,N_12221);
xnor U14961 (N_14961,N_12989,N_13770);
or U14962 (N_14962,N_12647,N_13898);
nor U14963 (N_14963,N_12950,N_12382);
and U14964 (N_14964,N_13346,N_13582);
nand U14965 (N_14965,N_13261,N_13240);
and U14966 (N_14966,N_13518,N_13975);
nand U14967 (N_14967,N_12527,N_12252);
or U14968 (N_14968,N_13376,N_13241);
or U14969 (N_14969,N_13464,N_13078);
and U14970 (N_14970,N_12848,N_12769);
nand U14971 (N_14971,N_13155,N_12058);
nand U14972 (N_14972,N_12096,N_12250);
nor U14973 (N_14973,N_13710,N_12061);
nor U14974 (N_14974,N_12596,N_12264);
nand U14975 (N_14975,N_13894,N_12095);
xnor U14976 (N_14976,N_12415,N_12444);
or U14977 (N_14977,N_12616,N_13645);
and U14978 (N_14978,N_13838,N_12010);
nor U14979 (N_14979,N_12533,N_13402);
nand U14980 (N_14980,N_13620,N_13077);
or U14981 (N_14981,N_13222,N_12925);
and U14982 (N_14982,N_13905,N_13186);
xor U14983 (N_14983,N_12215,N_12013);
xor U14984 (N_14984,N_13378,N_13791);
or U14985 (N_14985,N_13719,N_12164);
nor U14986 (N_14986,N_12601,N_13603);
or U14987 (N_14987,N_13565,N_12041);
nor U14988 (N_14988,N_12753,N_13874);
nand U14989 (N_14989,N_13168,N_13019);
nor U14990 (N_14990,N_13328,N_13868);
xor U14991 (N_14991,N_12049,N_13154);
nand U14992 (N_14992,N_13941,N_12019);
xor U14993 (N_14993,N_12008,N_13697);
and U14994 (N_14994,N_12208,N_12551);
xnor U14995 (N_14995,N_13720,N_13421);
xnor U14996 (N_14996,N_13887,N_12880);
nor U14997 (N_14997,N_13310,N_13117);
and U14998 (N_14998,N_13076,N_12091);
nand U14999 (N_14999,N_12766,N_13613);
nor U15000 (N_15000,N_13888,N_12100);
nor U15001 (N_15001,N_13242,N_13616);
and U15002 (N_15002,N_13828,N_13711);
and U15003 (N_15003,N_13493,N_13758);
or U15004 (N_15004,N_13435,N_12806);
nand U15005 (N_15005,N_12014,N_13722);
and U15006 (N_15006,N_13175,N_13972);
and U15007 (N_15007,N_12887,N_12252);
xor U15008 (N_15008,N_12082,N_12619);
nor U15009 (N_15009,N_13813,N_13551);
or U15010 (N_15010,N_13629,N_13195);
nor U15011 (N_15011,N_12973,N_13492);
nand U15012 (N_15012,N_13094,N_12690);
and U15013 (N_15013,N_12722,N_13898);
nor U15014 (N_15014,N_13305,N_13760);
or U15015 (N_15015,N_12185,N_12726);
nor U15016 (N_15016,N_12778,N_12144);
or U15017 (N_15017,N_13646,N_13861);
or U15018 (N_15018,N_13117,N_13609);
and U15019 (N_15019,N_13751,N_12802);
and U15020 (N_15020,N_13050,N_13801);
nand U15021 (N_15021,N_12639,N_12939);
nor U15022 (N_15022,N_12214,N_13706);
and U15023 (N_15023,N_12649,N_13159);
nand U15024 (N_15024,N_13601,N_12726);
xor U15025 (N_15025,N_13631,N_13223);
or U15026 (N_15026,N_12815,N_12509);
and U15027 (N_15027,N_12506,N_12227);
nand U15028 (N_15028,N_12845,N_13018);
nor U15029 (N_15029,N_13168,N_12760);
or U15030 (N_15030,N_13597,N_13078);
nor U15031 (N_15031,N_13507,N_13760);
nor U15032 (N_15032,N_13350,N_12478);
nor U15033 (N_15033,N_13941,N_12006);
nand U15034 (N_15034,N_12606,N_13270);
nand U15035 (N_15035,N_13230,N_12835);
nor U15036 (N_15036,N_12733,N_13652);
or U15037 (N_15037,N_12835,N_12805);
nand U15038 (N_15038,N_13840,N_13609);
and U15039 (N_15039,N_13727,N_13138);
nor U15040 (N_15040,N_12063,N_12555);
xor U15041 (N_15041,N_12988,N_12862);
xnor U15042 (N_15042,N_13686,N_13505);
and U15043 (N_15043,N_13716,N_12761);
nand U15044 (N_15044,N_13772,N_13893);
nor U15045 (N_15045,N_12043,N_13976);
nor U15046 (N_15046,N_13108,N_12510);
xnor U15047 (N_15047,N_13805,N_13917);
nand U15048 (N_15048,N_12131,N_13737);
nor U15049 (N_15049,N_13197,N_12066);
nand U15050 (N_15050,N_12605,N_13977);
xor U15051 (N_15051,N_13099,N_12296);
xnor U15052 (N_15052,N_13383,N_12800);
nand U15053 (N_15053,N_12832,N_13106);
nand U15054 (N_15054,N_13044,N_12832);
and U15055 (N_15055,N_12189,N_12585);
or U15056 (N_15056,N_12969,N_13539);
and U15057 (N_15057,N_12948,N_12956);
nor U15058 (N_15058,N_12298,N_12136);
nor U15059 (N_15059,N_12795,N_13106);
nor U15060 (N_15060,N_13655,N_12013);
or U15061 (N_15061,N_12682,N_12410);
or U15062 (N_15062,N_13305,N_12387);
xor U15063 (N_15063,N_13966,N_12209);
xor U15064 (N_15064,N_13118,N_12943);
nand U15065 (N_15065,N_13073,N_12335);
xor U15066 (N_15066,N_12804,N_12981);
and U15067 (N_15067,N_13722,N_12580);
or U15068 (N_15068,N_13925,N_12631);
nand U15069 (N_15069,N_12045,N_13596);
or U15070 (N_15070,N_12087,N_13472);
nor U15071 (N_15071,N_12135,N_13398);
nor U15072 (N_15072,N_12273,N_13767);
nand U15073 (N_15073,N_13844,N_12781);
nor U15074 (N_15074,N_13149,N_13867);
nor U15075 (N_15075,N_13444,N_13637);
or U15076 (N_15076,N_12676,N_12295);
or U15077 (N_15077,N_12488,N_13063);
nand U15078 (N_15078,N_12802,N_12304);
nor U15079 (N_15079,N_13485,N_12262);
nand U15080 (N_15080,N_12429,N_12435);
or U15081 (N_15081,N_13048,N_13453);
nor U15082 (N_15082,N_12557,N_12591);
nand U15083 (N_15083,N_13363,N_13354);
or U15084 (N_15084,N_13320,N_12767);
or U15085 (N_15085,N_12302,N_13613);
or U15086 (N_15086,N_13449,N_13702);
or U15087 (N_15087,N_13629,N_12949);
nor U15088 (N_15088,N_13859,N_12482);
nand U15089 (N_15089,N_13120,N_13384);
nand U15090 (N_15090,N_13724,N_13730);
nor U15091 (N_15091,N_13295,N_12680);
nand U15092 (N_15092,N_13313,N_12457);
nand U15093 (N_15093,N_12197,N_12875);
or U15094 (N_15094,N_13034,N_13386);
nand U15095 (N_15095,N_12860,N_12930);
or U15096 (N_15096,N_12971,N_13373);
or U15097 (N_15097,N_12496,N_12830);
nand U15098 (N_15098,N_12474,N_13002);
nor U15099 (N_15099,N_13074,N_12983);
nand U15100 (N_15100,N_12787,N_12673);
nor U15101 (N_15101,N_12975,N_13535);
nand U15102 (N_15102,N_13091,N_12922);
and U15103 (N_15103,N_12409,N_13284);
nor U15104 (N_15104,N_13825,N_12047);
nor U15105 (N_15105,N_12629,N_13321);
xor U15106 (N_15106,N_13943,N_13757);
nand U15107 (N_15107,N_13254,N_13515);
nand U15108 (N_15108,N_13132,N_12785);
nor U15109 (N_15109,N_12919,N_12080);
and U15110 (N_15110,N_12693,N_12271);
and U15111 (N_15111,N_13139,N_13645);
nor U15112 (N_15112,N_12677,N_13875);
nor U15113 (N_15113,N_13510,N_12331);
and U15114 (N_15114,N_12791,N_13045);
and U15115 (N_15115,N_13163,N_13425);
and U15116 (N_15116,N_12784,N_12728);
and U15117 (N_15117,N_13609,N_12752);
or U15118 (N_15118,N_13563,N_12583);
and U15119 (N_15119,N_13148,N_12503);
or U15120 (N_15120,N_12242,N_13354);
nand U15121 (N_15121,N_13757,N_13005);
nor U15122 (N_15122,N_12202,N_12692);
or U15123 (N_15123,N_12122,N_13926);
and U15124 (N_15124,N_12903,N_13545);
nor U15125 (N_15125,N_12068,N_12539);
or U15126 (N_15126,N_12512,N_13684);
nand U15127 (N_15127,N_12771,N_12512);
xnor U15128 (N_15128,N_12304,N_13420);
nand U15129 (N_15129,N_12936,N_13504);
nand U15130 (N_15130,N_13200,N_13990);
nor U15131 (N_15131,N_13574,N_12598);
nand U15132 (N_15132,N_13507,N_12411);
and U15133 (N_15133,N_13316,N_13072);
nand U15134 (N_15134,N_13415,N_13786);
nand U15135 (N_15135,N_13633,N_12223);
nor U15136 (N_15136,N_12402,N_13761);
and U15137 (N_15137,N_13016,N_12328);
or U15138 (N_15138,N_12562,N_13117);
nand U15139 (N_15139,N_13462,N_13531);
or U15140 (N_15140,N_13073,N_13478);
or U15141 (N_15141,N_13245,N_12572);
or U15142 (N_15142,N_12109,N_13847);
nor U15143 (N_15143,N_13758,N_13705);
nand U15144 (N_15144,N_13883,N_12491);
xor U15145 (N_15145,N_13800,N_13647);
and U15146 (N_15146,N_13886,N_12677);
nor U15147 (N_15147,N_12105,N_12182);
nor U15148 (N_15148,N_12942,N_12930);
or U15149 (N_15149,N_12336,N_12734);
or U15150 (N_15150,N_13387,N_12275);
and U15151 (N_15151,N_12443,N_12543);
nor U15152 (N_15152,N_12907,N_12794);
and U15153 (N_15153,N_13289,N_13590);
xor U15154 (N_15154,N_13878,N_12341);
nor U15155 (N_15155,N_12166,N_12311);
nand U15156 (N_15156,N_12238,N_12333);
and U15157 (N_15157,N_12798,N_12694);
or U15158 (N_15158,N_12482,N_13722);
or U15159 (N_15159,N_13360,N_12409);
nor U15160 (N_15160,N_13443,N_13939);
nand U15161 (N_15161,N_13986,N_13802);
and U15162 (N_15162,N_13773,N_13001);
and U15163 (N_15163,N_13806,N_12511);
nor U15164 (N_15164,N_13530,N_13068);
nand U15165 (N_15165,N_12110,N_12644);
nand U15166 (N_15166,N_12826,N_12309);
or U15167 (N_15167,N_13370,N_12245);
and U15168 (N_15168,N_12533,N_13348);
and U15169 (N_15169,N_12027,N_12738);
or U15170 (N_15170,N_13922,N_13215);
and U15171 (N_15171,N_12630,N_13653);
nand U15172 (N_15172,N_13844,N_12679);
xnor U15173 (N_15173,N_12284,N_12260);
nor U15174 (N_15174,N_13406,N_12943);
and U15175 (N_15175,N_13226,N_13049);
nor U15176 (N_15176,N_12680,N_12774);
xor U15177 (N_15177,N_12921,N_12601);
or U15178 (N_15178,N_12544,N_13015);
nor U15179 (N_15179,N_13206,N_13362);
and U15180 (N_15180,N_13471,N_12608);
or U15181 (N_15181,N_13126,N_13046);
and U15182 (N_15182,N_12942,N_13892);
or U15183 (N_15183,N_13191,N_13403);
nor U15184 (N_15184,N_12005,N_13012);
and U15185 (N_15185,N_12120,N_13039);
nand U15186 (N_15186,N_12199,N_12791);
nand U15187 (N_15187,N_12785,N_12951);
or U15188 (N_15188,N_13955,N_12904);
xnor U15189 (N_15189,N_13333,N_12554);
and U15190 (N_15190,N_13555,N_13038);
nor U15191 (N_15191,N_12992,N_12480);
nand U15192 (N_15192,N_12331,N_13276);
and U15193 (N_15193,N_12623,N_12074);
nor U15194 (N_15194,N_12569,N_12902);
and U15195 (N_15195,N_12290,N_12671);
nor U15196 (N_15196,N_13730,N_13807);
nor U15197 (N_15197,N_12848,N_12669);
xor U15198 (N_15198,N_13678,N_12451);
or U15199 (N_15199,N_12691,N_12211);
and U15200 (N_15200,N_12021,N_12202);
nor U15201 (N_15201,N_12927,N_12654);
and U15202 (N_15202,N_13821,N_12113);
or U15203 (N_15203,N_12406,N_12926);
or U15204 (N_15204,N_13113,N_12655);
xnor U15205 (N_15205,N_12904,N_12479);
nor U15206 (N_15206,N_13788,N_13005);
xnor U15207 (N_15207,N_13680,N_12702);
xor U15208 (N_15208,N_12422,N_12098);
nor U15209 (N_15209,N_13184,N_12521);
nand U15210 (N_15210,N_13517,N_12916);
and U15211 (N_15211,N_12533,N_12717);
or U15212 (N_15212,N_12447,N_13350);
or U15213 (N_15213,N_12113,N_13286);
nor U15214 (N_15214,N_13145,N_12761);
nor U15215 (N_15215,N_12515,N_12594);
nor U15216 (N_15216,N_13813,N_12867);
and U15217 (N_15217,N_12781,N_12836);
and U15218 (N_15218,N_13137,N_12990);
nor U15219 (N_15219,N_13628,N_13830);
or U15220 (N_15220,N_13621,N_12430);
and U15221 (N_15221,N_13596,N_12544);
or U15222 (N_15222,N_12533,N_13915);
or U15223 (N_15223,N_13603,N_12839);
or U15224 (N_15224,N_12272,N_12223);
nand U15225 (N_15225,N_12427,N_12176);
nand U15226 (N_15226,N_13829,N_12051);
nand U15227 (N_15227,N_12659,N_13835);
nand U15228 (N_15228,N_12413,N_13218);
nand U15229 (N_15229,N_13385,N_13723);
nand U15230 (N_15230,N_13560,N_13820);
and U15231 (N_15231,N_13971,N_13457);
or U15232 (N_15232,N_13636,N_12488);
nor U15233 (N_15233,N_13273,N_13380);
nor U15234 (N_15234,N_12816,N_12182);
nand U15235 (N_15235,N_13009,N_12158);
nor U15236 (N_15236,N_12023,N_12827);
and U15237 (N_15237,N_13130,N_13858);
xnor U15238 (N_15238,N_12135,N_12149);
xor U15239 (N_15239,N_13367,N_13962);
or U15240 (N_15240,N_12217,N_13090);
and U15241 (N_15241,N_12300,N_13616);
or U15242 (N_15242,N_13716,N_12074);
or U15243 (N_15243,N_12633,N_12374);
and U15244 (N_15244,N_13474,N_13847);
nor U15245 (N_15245,N_12109,N_12840);
or U15246 (N_15246,N_13685,N_13471);
nand U15247 (N_15247,N_12740,N_13031);
nand U15248 (N_15248,N_13659,N_12251);
or U15249 (N_15249,N_12362,N_12748);
and U15250 (N_15250,N_12196,N_12657);
or U15251 (N_15251,N_12705,N_13279);
nor U15252 (N_15252,N_12389,N_12336);
and U15253 (N_15253,N_12642,N_12281);
or U15254 (N_15254,N_12185,N_12813);
and U15255 (N_15255,N_13748,N_13164);
or U15256 (N_15256,N_12317,N_12435);
nor U15257 (N_15257,N_12801,N_13784);
nor U15258 (N_15258,N_12807,N_13717);
and U15259 (N_15259,N_13193,N_13571);
xnor U15260 (N_15260,N_12835,N_13986);
and U15261 (N_15261,N_13456,N_13157);
nand U15262 (N_15262,N_12596,N_12778);
and U15263 (N_15263,N_12978,N_13872);
xnor U15264 (N_15264,N_13326,N_12921);
nor U15265 (N_15265,N_13089,N_13909);
and U15266 (N_15266,N_12359,N_13901);
nor U15267 (N_15267,N_13739,N_12517);
xor U15268 (N_15268,N_12221,N_12829);
xor U15269 (N_15269,N_12089,N_13074);
or U15270 (N_15270,N_12450,N_13770);
xnor U15271 (N_15271,N_12865,N_12209);
nor U15272 (N_15272,N_13420,N_13390);
nor U15273 (N_15273,N_13976,N_12155);
and U15274 (N_15274,N_12641,N_12886);
or U15275 (N_15275,N_13568,N_12743);
nor U15276 (N_15276,N_13527,N_13149);
and U15277 (N_15277,N_12508,N_13556);
or U15278 (N_15278,N_13956,N_13929);
nand U15279 (N_15279,N_12962,N_13398);
nand U15280 (N_15280,N_12294,N_12428);
or U15281 (N_15281,N_13362,N_13233);
nor U15282 (N_15282,N_12615,N_12423);
and U15283 (N_15283,N_12699,N_12393);
nor U15284 (N_15284,N_13908,N_12983);
nor U15285 (N_15285,N_13926,N_12866);
nor U15286 (N_15286,N_12262,N_13819);
or U15287 (N_15287,N_12957,N_13955);
and U15288 (N_15288,N_13783,N_12659);
and U15289 (N_15289,N_13365,N_13245);
or U15290 (N_15290,N_13178,N_13297);
xor U15291 (N_15291,N_13003,N_12718);
nand U15292 (N_15292,N_13986,N_13124);
or U15293 (N_15293,N_12312,N_13851);
xor U15294 (N_15294,N_12650,N_12593);
or U15295 (N_15295,N_13626,N_12491);
nand U15296 (N_15296,N_12661,N_13096);
and U15297 (N_15297,N_13039,N_13672);
nor U15298 (N_15298,N_12834,N_13032);
nand U15299 (N_15299,N_13217,N_13262);
nor U15300 (N_15300,N_12403,N_12123);
nand U15301 (N_15301,N_12702,N_12359);
or U15302 (N_15302,N_12899,N_12706);
nor U15303 (N_15303,N_12696,N_12733);
and U15304 (N_15304,N_13975,N_13466);
and U15305 (N_15305,N_12664,N_13751);
xnor U15306 (N_15306,N_12769,N_13438);
and U15307 (N_15307,N_12717,N_13071);
and U15308 (N_15308,N_12134,N_12688);
and U15309 (N_15309,N_13027,N_13554);
nand U15310 (N_15310,N_12971,N_13411);
xor U15311 (N_15311,N_13654,N_12599);
or U15312 (N_15312,N_12824,N_12745);
or U15313 (N_15313,N_12224,N_13345);
or U15314 (N_15314,N_12258,N_12282);
or U15315 (N_15315,N_13868,N_13276);
or U15316 (N_15316,N_13511,N_13418);
nor U15317 (N_15317,N_12684,N_13465);
or U15318 (N_15318,N_13019,N_13002);
nand U15319 (N_15319,N_12679,N_12512);
nand U15320 (N_15320,N_13355,N_12387);
nor U15321 (N_15321,N_13701,N_12914);
nor U15322 (N_15322,N_12035,N_13330);
xnor U15323 (N_15323,N_13395,N_12758);
nand U15324 (N_15324,N_13691,N_12672);
nor U15325 (N_15325,N_13893,N_13489);
and U15326 (N_15326,N_13509,N_13702);
nand U15327 (N_15327,N_13843,N_13481);
or U15328 (N_15328,N_12952,N_13266);
or U15329 (N_15329,N_12294,N_12626);
or U15330 (N_15330,N_12987,N_12271);
nor U15331 (N_15331,N_12515,N_13086);
and U15332 (N_15332,N_13368,N_12308);
and U15333 (N_15333,N_12279,N_13475);
or U15334 (N_15334,N_12137,N_12294);
and U15335 (N_15335,N_13955,N_13279);
or U15336 (N_15336,N_13205,N_13815);
and U15337 (N_15337,N_13928,N_12241);
nand U15338 (N_15338,N_12619,N_12352);
and U15339 (N_15339,N_12953,N_13590);
nor U15340 (N_15340,N_13614,N_13251);
nand U15341 (N_15341,N_13853,N_12580);
nand U15342 (N_15342,N_12017,N_12226);
or U15343 (N_15343,N_13144,N_12299);
xor U15344 (N_15344,N_13984,N_13815);
nand U15345 (N_15345,N_12572,N_12958);
nor U15346 (N_15346,N_12809,N_12033);
and U15347 (N_15347,N_12436,N_13988);
nor U15348 (N_15348,N_13848,N_13179);
or U15349 (N_15349,N_13317,N_12638);
nor U15350 (N_15350,N_13985,N_12513);
and U15351 (N_15351,N_12264,N_12893);
and U15352 (N_15352,N_12716,N_12700);
or U15353 (N_15353,N_12553,N_13067);
and U15354 (N_15354,N_12391,N_13656);
xor U15355 (N_15355,N_12361,N_12195);
nor U15356 (N_15356,N_13906,N_13234);
and U15357 (N_15357,N_12069,N_12699);
and U15358 (N_15358,N_12989,N_12379);
nand U15359 (N_15359,N_13084,N_12694);
nor U15360 (N_15360,N_12239,N_13207);
or U15361 (N_15361,N_12805,N_12646);
xor U15362 (N_15362,N_13935,N_13694);
or U15363 (N_15363,N_13303,N_13107);
nand U15364 (N_15364,N_13613,N_12683);
nor U15365 (N_15365,N_12431,N_12909);
xor U15366 (N_15366,N_13951,N_12572);
nor U15367 (N_15367,N_13604,N_13962);
and U15368 (N_15368,N_13568,N_13497);
and U15369 (N_15369,N_13165,N_12710);
nand U15370 (N_15370,N_13669,N_13603);
or U15371 (N_15371,N_12818,N_13497);
nor U15372 (N_15372,N_12086,N_12573);
and U15373 (N_15373,N_13218,N_13786);
and U15374 (N_15374,N_12744,N_13752);
nand U15375 (N_15375,N_13450,N_13127);
nand U15376 (N_15376,N_13553,N_12865);
or U15377 (N_15377,N_13027,N_12921);
and U15378 (N_15378,N_13675,N_13431);
or U15379 (N_15379,N_13445,N_12805);
or U15380 (N_15380,N_13739,N_12117);
or U15381 (N_15381,N_12433,N_13830);
nand U15382 (N_15382,N_13902,N_12748);
and U15383 (N_15383,N_13927,N_13195);
and U15384 (N_15384,N_13653,N_13149);
and U15385 (N_15385,N_12028,N_12168);
or U15386 (N_15386,N_13868,N_12613);
and U15387 (N_15387,N_13127,N_13745);
or U15388 (N_15388,N_13320,N_13070);
or U15389 (N_15389,N_12741,N_12490);
and U15390 (N_15390,N_12077,N_12559);
or U15391 (N_15391,N_12865,N_12787);
nand U15392 (N_15392,N_12899,N_12499);
nand U15393 (N_15393,N_13438,N_13734);
nor U15394 (N_15394,N_12047,N_12604);
nand U15395 (N_15395,N_13636,N_13150);
nand U15396 (N_15396,N_12781,N_12561);
nand U15397 (N_15397,N_13567,N_12792);
nand U15398 (N_15398,N_12865,N_13815);
xnor U15399 (N_15399,N_13858,N_12274);
nor U15400 (N_15400,N_13119,N_12311);
nand U15401 (N_15401,N_13678,N_12706);
nand U15402 (N_15402,N_13540,N_12074);
nand U15403 (N_15403,N_12146,N_13065);
or U15404 (N_15404,N_13424,N_12416);
nor U15405 (N_15405,N_12592,N_13065);
nand U15406 (N_15406,N_13040,N_13111);
nor U15407 (N_15407,N_13402,N_12622);
and U15408 (N_15408,N_13161,N_12204);
and U15409 (N_15409,N_13526,N_13229);
and U15410 (N_15410,N_12735,N_12231);
xnor U15411 (N_15411,N_13852,N_12987);
nand U15412 (N_15412,N_12466,N_13442);
xnor U15413 (N_15413,N_12051,N_13157);
or U15414 (N_15414,N_12082,N_12743);
nand U15415 (N_15415,N_12755,N_12637);
nor U15416 (N_15416,N_13763,N_13570);
and U15417 (N_15417,N_13926,N_12840);
nand U15418 (N_15418,N_12055,N_13117);
nand U15419 (N_15419,N_12513,N_12138);
and U15420 (N_15420,N_13015,N_12508);
nor U15421 (N_15421,N_13156,N_13847);
and U15422 (N_15422,N_12455,N_12223);
nor U15423 (N_15423,N_12622,N_12924);
and U15424 (N_15424,N_12504,N_12173);
or U15425 (N_15425,N_12730,N_13755);
or U15426 (N_15426,N_13471,N_12451);
or U15427 (N_15427,N_12618,N_13956);
xor U15428 (N_15428,N_12689,N_12232);
or U15429 (N_15429,N_13394,N_13451);
or U15430 (N_15430,N_12100,N_12122);
nand U15431 (N_15431,N_12482,N_12423);
xor U15432 (N_15432,N_12828,N_12394);
nor U15433 (N_15433,N_13395,N_12125);
nand U15434 (N_15434,N_12677,N_13492);
xor U15435 (N_15435,N_13730,N_12227);
or U15436 (N_15436,N_12344,N_12477);
or U15437 (N_15437,N_13794,N_12841);
nor U15438 (N_15438,N_13635,N_12440);
nor U15439 (N_15439,N_12610,N_13590);
or U15440 (N_15440,N_13640,N_13119);
or U15441 (N_15441,N_12317,N_12206);
nor U15442 (N_15442,N_13442,N_13972);
and U15443 (N_15443,N_13761,N_13773);
and U15444 (N_15444,N_12593,N_12008);
nand U15445 (N_15445,N_13769,N_13344);
xor U15446 (N_15446,N_13636,N_13413);
and U15447 (N_15447,N_12804,N_12034);
and U15448 (N_15448,N_12903,N_12635);
nor U15449 (N_15449,N_12643,N_13701);
and U15450 (N_15450,N_13761,N_12293);
and U15451 (N_15451,N_13366,N_12384);
and U15452 (N_15452,N_13075,N_13100);
nand U15453 (N_15453,N_12832,N_12231);
and U15454 (N_15454,N_12324,N_13720);
nand U15455 (N_15455,N_12595,N_12781);
nor U15456 (N_15456,N_12239,N_13750);
nor U15457 (N_15457,N_12259,N_12339);
or U15458 (N_15458,N_12709,N_12549);
nor U15459 (N_15459,N_13324,N_13128);
or U15460 (N_15460,N_12485,N_12334);
or U15461 (N_15461,N_12256,N_13286);
xor U15462 (N_15462,N_13460,N_12432);
nor U15463 (N_15463,N_13301,N_13690);
and U15464 (N_15464,N_12705,N_13370);
and U15465 (N_15465,N_13588,N_12427);
and U15466 (N_15466,N_12412,N_12271);
or U15467 (N_15467,N_13879,N_12057);
and U15468 (N_15468,N_13237,N_13790);
nand U15469 (N_15469,N_12457,N_12477);
nand U15470 (N_15470,N_13170,N_12992);
nor U15471 (N_15471,N_13620,N_13403);
nor U15472 (N_15472,N_12771,N_12647);
nor U15473 (N_15473,N_12790,N_13238);
nand U15474 (N_15474,N_12780,N_13275);
nand U15475 (N_15475,N_13914,N_13077);
and U15476 (N_15476,N_13590,N_12004);
nand U15477 (N_15477,N_13896,N_12100);
and U15478 (N_15478,N_12615,N_12681);
nor U15479 (N_15479,N_13968,N_12900);
or U15480 (N_15480,N_13715,N_13371);
and U15481 (N_15481,N_12395,N_12805);
nor U15482 (N_15482,N_13818,N_12390);
nand U15483 (N_15483,N_12360,N_13484);
nand U15484 (N_15484,N_12232,N_13593);
and U15485 (N_15485,N_13340,N_13828);
nand U15486 (N_15486,N_12144,N_13264);
nand U15487 (N_15487,N_12549,N_12120);
xor U15488 (N_15488,N_13242,N_12933);
nor U15489 (N_15489,N_13394,N_12794);
nand U15490 (N_15490,N_12692,N_13183);
nand U15491 (N_15491,N_12807,N_13747);
and U15492 (N_15492,N_13291,N_13926);
or U15493 (N_15493,N_13549,N_13777);
nor U15494 (N_15494,N_13366,N_13376);
nor U15495 (N_15495,N_12110,N_12726);
nor U15496 (N_15496,N_12536,N_13239);
xor U15497 (N_15497,N_12989,N_12231);
or U15498 (N_15498,N_13687,N_12628);
and U15499 (N_15499,N_12165,N_13321);
or U15500 (N_15500,N_13388,N_13353);
nand U15501 (N_15501,N_13586,N_12545);
xnor U15502 (N_15502,N_12522,N_13983);
nand U15503 (N_15503,N_12225,N_13102);
nand U15504 (N_15504,N_12544,N_12507);
and U15505 (N_15505,N_12550,N_12725);
nor U15506 (N_15506,N_13925,N_13857);
xor U15507 (N_15507,N_13379,N_13293);
nand U15508 (N_15508,N_13815,N_12668);
and U15509 (N_15509,N_13233,N_12078);
or U15510 (N_15510,N_12360,N_13749);
nand U15511 (N_15511,N_13881,N_13451);
or U15512 (N_15512,N_13898,N_13104);
and U15513 (N_15513,N_12809,N_12443);
and U15514 (N_15514,N_12078,N_12312);
and U15515 (N_15515,N_13741,N_12933);
nand U15516 (N_15516,N_12043,N_12380);
or U15517 (N_15517,N_12632,N_13860);
nand U15518 (N_15518,N_13315,N_12323);
nor U15519 (N_15519,N_12000,N_13116);
or U15520 (N_15520,N_13897,N_12962);
or U15521 (N_15521,N_13612,N_12328);
or U15522 (N_15522,N_12046,N_12924);
or U15523 (N_15523,N_12737,N_13008);
nor U15524 (N_15524,N_13781,N_12794);
nand U15525 (N_15525,N_12917,N_13279);
nand U15526 (N_15526,N_12059,N_13521);
and U15527 (N_15527,N_12556,N_12381);
and U15528 (N_15528,N_13425,N_13740);
or U15529 (N_15529,N_13794,N_13184);
nor U15530 (N_15530,N_12314,N_13407);
xor U15531 (N_15531,N_12309,N_12213);
or U15532 (N_15532,N_13782,N_12921);
nor U15533 (N_15533,N_12775,N_12773);
nand U15534 (N_15534,N_13469,N_12230);
nand U15535 (N_15535,N_12879,N_13550);
nand U15536 (N_15536,N_12648,N_12149);
nand U15537 (N_15537,N_13043,N_13646);
and U15538 (N_15538,N_12367,N_12806);
nand U15539 (N_15539,N_13545,N_13702);
nor U15540 (N_15540,N_12685,N_12462);
xnor U15541 (N_15541,N_12641,N_12607);
or U15542 (N_15542,N_13541,N_13251);
nor U15543 (N_15543,N_13793,N_12502);
nand U15544 (N_15544,N_13115,N_13770);
and U15545 (N_15545,N_13722,N_12877);
nor U15546 (N_15546,N_12380,N_13381);
nor U15547 (N_15547,N_13625,N_12233);
nor U15548 (N_15548,N_12773,N_13828);
nand U15549 (N_15549,N_12333,N_13054);
and U15550 (N_15550,N_12451,N_13090);
or U15551 (N_15551,N_13868,N_13626);
or U15552 (N_15552,N_13195,N_12609);
nand U15553 (N_15553,N_12040,N_12008);
or U15554 (N_15554,N_13748,N_12897);
or U15555 (N_15555,N_13321,N_13537);
nand U15556 (N_15556,N_13943,N_12332);
nor U15557 (N_15557,N_13037,N_12637);
and U15558 (N_15558,N_13132,N_13148);
nor U15559 (N_15559,N_13731,N_13535);
xnor U15560 (N_15560,N_13216,N_12832);
nand U15561 (N_15561,N_12744,N_13430);
and U15562 (N_15562,N_13400,N_13237);
and U15563 (N_15563,N_13928,N_13391);
nor U15564 (N_15564,N_13648,N_13835);
or U15565 (N_15565,N_12495,N_13658);
nor U15566 (N_15566,N_13353,N_12573);
nor U15567 (N_15567,N_12309,N_13252);
or U15568 (N_15568,N_12390,N_13089);
or U15569 (N_15569,N_13652,N_12472);
nand U15570 (N_15570,N_12638,N_12945);
and U15571 (N_15571,N_13222,N_12009);
nor U15572 (N_15572,N_12881,N_12551);
nor U15573 (N_15573,N_12769,N_12187);
and U15574 (N_15574,N_12477,N_12214);
nand U15575 (N_15575,N_13909,N_12269);
or U15576 (N_15576,N_12514,N_13230);
nor U15577 (N_15577,N_12353,N_12362);
nor U15578 (N_15578,N_12929,N_13301);
or U15579 (N_15579,N_12922,N_12569);
nand U15580 (N_15580,N_12504,N_12309);
or U15581 (N_15581,N_13165,N_13420);
and U15582 (N_15582,N_13972,N_12779);
nor U15583 (N_15583,N_13170,N_12383);
nand U15584 (N_15584,N_12395,N_12396);
nand U15585 (N_15585,N_12605,N_12310);
or U15586 (N_15586,N_12995,N_12525);
xnor U15587 (N_15587,N_13515,N_12478);
nor U15588 (N_15588,N_13344,N_13065);
and U15589 (N_15589,N_12531,N_13665);
nor U15590 (N_15590,N_12429,N_13020);
and U15591 (N_15591,N_12254,N_12627);
nor U15592 (N_15592,N_12664,N_12441);
and U15593 (N_15593,N_12008,N_12180);
or U15594 (N_15594,N_13329,N_13386);
xor U15595 (N_15595,N_12332,N_12614);
and U15596 (N_15596,N_13520,N_13942);
nor U15597 (N_15597,N_13149,N_13302);
nor U15598 (N_15598,N_13693,N_13492);
nor U15599 (N_15599,N_13258,N_12246);
nand U15600 (N_15600,N_12985,N_12120);
or U15601 (N_15601,N_13295,N_13916);
or U15602 (N_15602,N_13427,N_12714);
and U15603 (N_15603,N_13430,N_13724);
and U15604 (N_15604,N_12114,N_13492);
nand U15605 (N_15605,N_13835,N_12121);
and U15606 (N_15606,N_13045,N_13942);
and U15607 (N_15607,N_12592,N_13376);
or U15608 (N_15608,N_12910,N_12413);
or U15609 (N_15609,N_12001,N_13888);
or U15610 (N_15610,N_12414,N_13582);
or U15611 (N_15611,N_13658,N_13386);
nor U15612 (N_15612,N_12328,N_13921);
nand U15613 (N_15613,N_12017,N_13536);
nor U15614 (N_15614,N_12949,N_12244);
nand U15615 (N_15615,N_12395,N_13947);
and U15616 (N_15616,N_12130,N_13076);
and U15617 (N_15617,N_13145,N_13479);
and U15618 (N_15618,N_13363,N_13310);
and U15619 (N_15619,N_13151,N_13092);
nand U15620 (N_15620,N_12312,N_12143);
and U15621 (N_15621,N_13478,N_13763);
and U15622 (N_15622,N_13593,N_12924);
or U15623 (N_15623,N_12996,N_12345);
nor U15624 (N_15624,N_13541,N_12843);
or U15625 (N_15625,N_12051,N_12114);
nor U15626 (N_15626,N_13606,N_12626);
and U15627 (N_15627,N_12357,N_12725);
and U15628 (N_15628,N_12838,N_12031);
xor U15629 (N_15629,N_12594,N_12453);
and U15630 (N_15630,N_13373,N_13431);
nor U15631 (N_15631,N_12707,N_12052);
or U15632 (N_15632,N_13224,N_13724);
nand U15633 (N_15633,N_13230,N_13568);
nand U15634 (N_15634,N_13767,N_13475);
and U15635 (N_15635,N_12435,N_12296);
or U15636 (N_15636,N_12602,N_12546);
nor U15637 (N_15637,N_12414,N_12180);
nor U15638 (N_15638,N_13052,N_13956);
nor U15639 (N_15639,N_12519,N_12589);
and U15640 (N_15640,N_13933,N_13196);
nand U15641 (N_15641,N_12576,N_12117);
nor U15642 (N_15642,N_12565,N_12533);
nor U15643 (N_15643,N_12753,N_13248);
nand U15644 (N_15644,N_12980,N_13888);
and U15645 (N_15645,N_13187,N_12498);
nand U15646 (N_15646,N_12167,N_13494);
nand U15647 (N_15647,N_13643,N_12369);
nor U15648 (N_15648,N_13722,N_13742);
nand U15649 (N_15649,N_12523,N_13318);
or U15650 (N_15650,N_12723,N_12388);
nand U15651 (N_15651,N_12714,N_12761);
and U15652 (N_15652,N_13758,N_12522);
nand U15653 (N_15653,N_12952,N_12627);
nand U15654 (N_15654,N_13402,N_12932);
and U15655 (N_15655,N_12350,N_13791);
and U15656 (N_15656,N_12940,N_12276);
and U15657 (N_15657,N_13991,N_13494);
xor U15658 (N_15658,N_12867,N_12488);
or U15659 (N_15659,N_13982,N_12385);
xnor U15660 (N_15660,N_12475,N_12069);
and U15661 (N_15661,N_13558,N_13192);
and U15662 (N_15662,N_13730,N_12278);
nor U15663 (N_15663,N_12092,N_12221);
nand U15664 (N_15664,N_12240,N_12043);
nand U15665 (N_15665,N_12005,N_13643);
nor U15666 (N_15666,N_13292,N_12878);
or U15667 (N_15667,N_12414,N_12217);
xnor U15668 (N_15668,N_13074,N_12647);
nand U15669 (N_15669,N_13566,N_12505);
nand U15670 (N_15670,N_12799,N_12747);
nand U15671 (N_15671,N_12475,N_12922);
nor U15672 (N_15672,N_13070,N_12775);
or U15673 (N_15673,N_13535,N_13158);
or U15674 (N_15674,N_13970,N_13525);
or U15675 (N_15675,N_13155,N_12376);
xor U15676 (N_15676,N_13210,N_12578);
nor U15677 (N_15677,N_13209,N_13450);
and U15678 (N_15678,N_12895,N_13322);
nand U15679 (N_15679,N_12000,N_12761);
nand U15680 (N_15680,N_12990,N_13081);
and U15681 (N_15681,N_13564,N_13277);
nor U15682 (N_15682,N_13922,N_13837);
nand U15683 (N_15683,N_13479,N_12425);
and U15684 (N_15684,N_13828,N_12305);
and U15685 (N_15685,N_12551,N_13658);
or U15686 (N_15686,N_13898,N_12909);
or U15687 (N_15687,N_13884,N_13815);
and U15688 (N_15688,N_13608,N_13836);
xor U15689 (N_15689,N_12842,N_13808);
and U15690 (N_15690,N_12345,N_13543);
or U15691 (N_15691,N_12684,N_13194);
nand U15692 (N_15692,N_13556,N_13750);
and U15693 (N_15693,N_12815,N_13349);
nor U15694 (N_15694,N_12820,N_13890);
xnor U15695 (N_15695,N_12834,N_13756);
nand U15696 (N_15696,N_13607,N_13825);
nor U15697 (N_15697,N_13473,N_13871);
nor U15698 (N_15698,N_12722,N_13099);
nor U15699 (N_15699,N_12239,N_12168);
or U15700 (N_15700,N_13394,N_13902);
xor U15701 (N_15701,N_13525,N_12775);
nand U15702 (N_15702,N_13973,N_13722);
nor U15703 (N_15703,N_13995,N_13517);
nor U15704 (N_15704,N_12608,N_13873);
nor U15705 (N_15705,N_12727,N_12626);
nand U15706 (N_15706,N_13953,N_13382);
xor U15707 (N_15707,N_12233,N_13425);
nor U15708 (N_15708,N_12514,N_12144);
or U15709 (N_15709,N_12292,N_13647);
xnor U15710 (N_15710,N_13764,N_13948);
and U15711 (N_15711,N_12882,N_12100);
and U15712 (N_15712,N_12992,N_13824);
or U15713 (N_15713,N_12056,N_12150);
xor U15714 (N_15714,N_12388,N_13606);
xnor U15715 (N_15715,N_12521,N_13320);
nand U15716 (N_15716,N_12089,N_12689);
nor U15717 (N_15717,N_12560,N_12478);
nand U15718 (N_15718,N_12180,N_13937);
or U15719 (N_15719,N_12861,N_13772);
nand U15720 (N_15720,N_13575,N_12042);
or U15721 (N_15721,N_12520,N_13609);
nand U15722 (N_15722,N_13208,N_13982);
or U15723 (N_15723,N_13661,N_13126);
nor U15724 (N_15724,N_13926,N_13955);
xor U15725 (N_15725,N_12023,N_13731);
or U15726 (N_15726,N_12602,N_13857);
or U15727 (N_15727,N_12713,N_13401);
xor U15728 (N_15728,N_13849,N_13932);
nand U15729 (N_15729,N_12113,N_12365);
nand U15730 (N_15730,N_13134,N_13231);
nand U15731 (N_15731,N_13729,N_12184);
nand U15732 (N_15732,N_13809,N_13106);
and U15733 (N_15733,N_12038,N_12219);
and U15734 (N_15734,N_13096,N_12943);
or U15735 (N_15735,N_12447,N_13687);
or U15736 (N_15736,N_13322,N_13515);
nand U15737 (N_15737,N_13884,N_12656);
and U15738 (N_15738,N_13161,N_12978);
nor U15739 (N_15739,N_12389,N_12010);
nor U15740 (N_15740,N_12144,N_13255);
and U15741 (N_15741,N_12086,N_12612);
and U15742 (N_15742,N_12332,N_12361);
or U15743 (N_15743,N_13390,N_12602);
nor U15744 (N_15744,N_12286,N_12475);
nand U15745 (N_15745,N_12077,N_12186);
xnor U15746 (N_15746,N_12588,N_12051);
nand U15747 (N_15747,N_13679,N_12570);
and U15748 (N_15748,N_13938,N_12249);
nand U15749 (N_15749,N_12909,N_12633);
and U15750 (N_15750,N_13243,N_12980);
or U15751 (N_15751,N_12336,N_12195);
or U15752 (N_15752,N_13890,N_13130);
nand U15753 (N_15753,N_13044,N_13523);
and U15754 (N_15754,N_12253,N_13330);
nand U15755 (N_15755,N_12480,N_12860);
nand U15756 (N_15756,N_13423,N_13676);
and U15757 (N_15757,N_13640,N_13801);
nor U15758 (N_15758,N_12197,N_13404);
nand U15759 (N_15759,N_12197,N_13683);
or U15760 (N_15760,N_12036,N_12480);
and U15761 (N_15761,N_13840,N_12485);
and U15762 (N_15762,N_12174,N_12806);
and U15763 (N_15763,N_12252,N_13606);
nor U15764 (N_15764,N_12356,N_13698);
and U15765 (N_15765,N_12988,N_12263);
xor U15766 (N_15766,N_13610,N_13408);
or U15767 (N_15767,N_12843,N_13330);
or U15768 (N_15768,N_12019,N_12934);
and U15769 (N_15769,N_13539,N_12421);
nor U15770 (N_15770,N_12706,N_13401);
nand U15771 (N_15771,N_12734,N_13188);
nor U15772 (N_15772,N_13063,N_12538);
xor U15773 (N_15773,N_13804,N_13390);
nor U15774 (N_15774,N_13859,N_13241);
and U15775 (N_15775,N_12856,N_12174);
nor U15776 (N_15776,N_12484,N_13599);
nor U15777 (N_15777,N_13468,N_13129);
and U15778 (N_15778,N_13220,N_12487);
xnor U15779 (N_15779,N_12615,N_12389);
nand U15780 (N_15780,N_13432,N_13810);
xor U15781 (N_15781,N_12982,N_12292);
nand U15782 (N_15782,N_12175,N_12051);
or U15783 (N_15783,N_13377,N_12537);
or U15784 (N_15784,N_13526,N_13146);
and U15785 (N_15785,N_13963,N_12420);
or U15786 (N_15786,N_12406,N_13315);
nor U15787 (N_15787,N_12220,N_12152);
xor U15788 (N_15788,N_12071,N_13381);
nand U15789 (N_15789,N_13851,N_12569);
or U15790 (N_15790,N_12122,N_13515);
or U15791 (N_15791,N_13456,N_12835);
nand U15792 (N_15792,N_12836,N_12488);
or U15793 (N_15793,N_12874,N_13029);
or U15794 (N_15794,N_13302,N_12999);
nand U15795 (N_15795,N_13967,N_12006);
nand U15796 (N_15796,N_13002,N_12932);
and U15797 (N_15797,N_12047,N_12206);
xor U15798 (N_15798,N_13039,N_13047);
and U15799 (N_15799,N_12780,N_13454);
or U15800 (N_15800,N_13976,N_13828);
and U15801 (N_15801,N_12887,N_13010);
nand U15802 (N_15802,N_12187,N_13902);
nor U15803 (N_15803,N_12783,N_12597);
and U15804 (N_15804,N_12083,N_13717);
nand U15805 (N_15805,N_12706,N_13831);
and U15806 (N_15806,N_12082,N_12471);
nand U15807 (N_15807,N_12735,N_12667);
and U15808 (N_15808,N_12765,N_13018);
nor U15809 (N_15809,N_13122,N_12570);
nand U15810 (N_15810,N_13752,N_13165);
nor U15811 (N_15811,N_13886,N_13052);
or U15812 (N_15812,N_12542,N_12144);
or U15813 (N_15813,N_13465,N_13995);
xor U15814 (N_15814,N_12978,N_13004);
nor U15815 (N_15815,N_12608,N_12518);
nor U15816 (N_15816,N_12670,N_13916);
or U15817 (N_15817,N_12240,N_13335);
nor U15818 (N_15818,N_12866,N_12575);
nor U15819 (N_15819,N_12113,N_13460);
and U15820 (N_15820,N_12504,N_12546);
nand U15821 (N_15821,N_13439,N_12529);
or U15822 (N_15822,N_13326,N_13706);
xor U15823 (N_15823,N_13519,N_12099);
nor U15824 (N_15824,N_12083,N_12095);
and U15825 (N_15825,N_12984,N_12952);
and U15826 (N_15826,N_12786,N_12264);
or U15827 (N_15827,N_12569,N_12672);
nor U15828 (N_15828,N_13857,N_13137);
nand U15829 (N_15829,N_13155,N_13924);
nand U15830 (N_15830,N_12973,N_12418);
nand U15831 (N_15831,N_12535,N_13988);
nand U15832 (N_15832,N_12403,N_12634);
and U15833 (N_15833,N_12505,N_13557);
nor U15834 (N_15834,N_13765,N_12366);
or U15835 (N_15835,N_13059,N_12089);
nor U15836 (N_15836,N_12237,N_13388);
nand U15837 (N_15837,N_13590,N_12088);
or U15838 (N_15838,N_13842,N_13710);
or U15839 (N_15839,N_13424,N_12473);
and U15840 (N_15840,N_12558,N_12528);
and U15841 (N_15841,N_13394,N_13568);
nor U15842 (N_15842,N_12965,N_12539);
and U15843 (N_15843,N_13438,N_12412);
nor U15844 (N_15844,N_13766,N_12499);
xnor U15845 (N_15845,N_13486,N_12806);
xor U15846 (N_15846,N_13728,N_13762);
or U15847 (N_15847,N_12626,N_13665);
nand U15848 (N_15848,N_13513,N_12258);
nor U15849 (N_15849,N_13594,N_13331);
and U15850 (N_15850,N_12406,N_13932);
nor U15851 (N_15851,N_13221,N_13700);
nand U15852 (N_15852,N_13457,N_12385);
nand U15853 (N_15853,N_13204,N_12139);
nor U15854 (N_15854,N_12752,N_12313);
nand U15855 (N_15855,N_12739,N_12077);
nand U15856 (N_15856,N_12498,N_12612);
nand U15857 (N_15857,N_12638,N_13134);
nor U15858 (N_15858,N_13384,N_12163);
or U15859 (N_15859,N_12402,N_12974);
or U15860 (N_15860,N_13808,N_12739);
and U15861 (N_15861,N_12474,N_13112);
or U15862 (N_15862,N_13144,N_13853);
or U15863 (N_15863,N_12199,N_12531);
nand U15864 (N_15864,N_12741,N_13597);
nand U15865 (N_15865,N_12569,N_12051);
nor U15866 (N_15866,N_13852,N_13052);
nand U15867 (N_15867,N_12622,N_13008);
or U15868 (N_15868,N_13537,N_13089);
or U15869 (N_15869,N_13149,N_13620);
nand U15870 (N_15870,N_12131,N_13623);
nor U15871 (N_15871,N_12814,N_13957);
nor U15872 (N_15872,N_13972,N_13551);
nand U15873 (N_15873,N_12376,N_13131);
nor U15874 (N_15874,N_13043,N_12739);
and U15875 (N_15875,N_13470,N_12216);
or U15876 (N_15876,N_12778,N_12497);
or U15877 (N_15877,N_13233,N_13103);
and U15878 (N_15878,N_13448,N_12930);
nor U15879 (N_15879,N_13775,N_12206);
xnor U15880 (N_15880,N_13078,N_13315);
xor U15881 (N_15881,N_12385,N_12211);
or U15882 (N_15882,N_12521,N_13188);
nand U15883 (N_15883,N_12339,N_13907);
or U15884 (N_15884,N_13392,N_12827);
or U15885 (N_15885,N_12222,N_13417);
or U15886 (N_15886,N_13584,N_13188);
xnor U15887 (N_15887,N_12124,N_12696);
and U15888 (N_15888,N_13283,N_12921);
and U15889 (N_15889,N_12511,N_12374);
nand U15890 (N_15890,N_13345,N_12435);
and U15891 (N_15891,N_12018,N_13867);
nor U15892 (N_15892,N_12916,N_13680);
or U15893 (N_15893,N_13961,N_13730);
nand U15894 (N_15894,N_12946,N_12149);
nand U15895 (N_15895,N_13969,N_12360);
or U15896 (N_15896,N_12456,N_12727);
and U15897 (N_15897,N_13801,N_12124);
xor U15898 (N_15898,N_12381,N_12217);
xnor U15899 (N_15899,N_12622,N_13908);
nand U15900 (N_15900,N_12014,N_13896);
nor U15901 (N_15901,N_12224,N_13310);
or U15902 (N_15902,N_12927,N_13657);
nand U15903 (N_15903,N_13715,N_13281);
xnor U15904 (N_15904,N_13692,N_13160);
or U15905 (N_15905,N_13072,N_13351);
xnor U15906 (N_15906,N_12012,N_12795);
or U15907 (N_15907,N_12510,N_13993);
and U15908 (N_15908,N_13796,N_13969);
nand U15909 (N_15909,N_13633,N_12805);
nand U15910 (N_15910,N_12833,N_13816);
and U15911 (N_15911,N_12334,N_13374);
and U15912 (N_15912,N_13360,N_13990);
nor U15913 (N_15913,N_12116,N_12568);
nand U15914 (N_15914,N_12632,N_12569);
nand U15915 (N_15915,N_12310,N_13931);
and U15916 (N_15916,N_13692,N_12975);
nor U15917 (N_15917,N_12393,N_12912);
or U15918 (N_15918,N_13475,N_13472);
xnor U15919 (N_15919,N_13336,N_12657);
or U15920 (N_15920,N_13247,N_13201);
or U15921 (N_15921,N_13399,N_12062);
nor U15922 (N_15922,N_13439,N_13720);
nand U15923 (N_15923,N_13231,N_12977);
and U15924 (N_15924,N_13373,N_13583);
and U15925 (N_15925,N_13263,N_12049);
nand U15926 (N_15926,N_13073,N_13042);
and U15927 (N_15927,N_13823,N_13982);
nand U15928 (N_15928,N_13843,N_12342);
nand U15929 (N_15929,N_12692,N_12424);
nand U15930 (N_15930,N_12095,N_12267);
or U15931 (N_15931,N_13457,N_12633);
xor U15932 (N_15932,N_13322,N_12824);
nor U15933 (N_15933,N_12687,N_13707);
or U15934 (N_15934,N_13191,N_12755);
nor U15935 (N_15935,N_13082,N_12228);
nor U15936 (N_15936,N_12673,N_13275);
xnor U15937 (N_15937,N_12815,N_13634);
nor U15938 (N_15938,N_13304,N_13024);
xnor U15939 (N_15939,N_13265,N_13014);
or U15940 (N_15940,N_12564,N_13688);
nor U15941 (N_15941,N_13589,N_12581);
nand U15942 (N_15942,N_13426,N_13253);
nor U15943 (N_15943,N_12652,N_13096);
or U15944 (N_15944,N_13708,N_12941);
nand U15945 (N_15945,N_13178,N_13521);
nand U15946 (N_15946,N_13233,N_13262);
nand U15947 (N_15947,N_12595,N_12930);
and U15948 (N_15948,N_13473,N_12535);
or U15949 (N_15949,N_12534,N_12600);
nor U15950 (N_15950,N_13497,N_13467);
nand U15951 (N_15951,N_12364,N_13104);
nand U15952 (N_15952,N_12480,N_12286);
or U15953 (N_15953,N_13393,N_12485);
or U15954 (N_15954,N_13996,N_13760);
or U15955 (N_15955,N_13187,N_12815);
and U15956 (N_15956,N_13481,N_12506);
nand U15957 (N_15957,N_13965,N_12445);
or U15958 (N_15958,N_12945,N_13377);
and U15959 (N_15959,N_12687,N_13883);
or U15960 (N_15960,N_12109,N_13729);
nand U15961 (N_15961,N_13619,N_13683);
nor U15962 (N_15962,N_13851,N_13532);
or U15963 (N_15963,N_13158,N_12334);
or U15964 (N_15964,N_12652,N_12805);
or U15965 (N_15965,N_13065,N_13261);
or U15966 (N_15966,N_13110,N_12767);
nor U15967 (N_15967,N_13466,N_12112);
nand U15968 (N_15968,N_13504,N_12696);
nand U15969 (N_15969,N_13737,N_12267);
and U15970 (N_15970,N_13733,N_12455);
nand U15971 (N_15971,N_12739,N_12180);
nand U15972 (N_15972,N_13479,N_13394);
and U15973 (N_15973,N_12739,N_12318);
and U15974 (N_15974,N_12947,N_13679);
and U15975 (N_15975,N_13967,N_12534);
xor U15976 (N_15976,N_13833,N_13159);
nand U15977 (N_15977,N_13608,N_13647);
nor U15978 (N_15978,N_12974,N_12794);
nand U15979 (N_15979,N_12910,N_13273);
or U15980 (N_15980,N_12546,N_12384);
nor U15981 (N_15981,N_13793,N_13515);
nand U15982 (N_15982,N_12721,N_12037);
and U15983 (N_15983,N_12379,N_12141);
nor U15984 (N_15984,N_12503,N_12687);
or U15985 (N_15985,N_13663,N_13449);
nand U15986 (N_15986,N_12579,N_12344);
or U15987 (N_15987,N_12861,N_13868);
nand U15988 (N_15988,N_13029,N_13618);
nand U15989 (N_15989,N_12250,N_12500);
and U15990 (N_15990,N_12247,N_13221);
nor U15991 (N_15991,N_13086,N_13990);
nand U15992 (N_15992,N_12227,N_12842);
nand U15993 (N_15993,N_13910,N_13117);
nand U15994 (N_15994,N_13906,N_12448);
nand U15995 (N_15995,N_12725,N_12372);
and U15996 (N_15996,N_12195,N_13664);
or U15997 (N_15997,N_12893,N_12118);
nor U15998 (N_15998,N_12757,N_13701);
and U15999 (N_15999,N_13432,N_13975);
nor U16000 (N_16000,N_14508,N_15246);
or U16001 (N_16001,N_15033,N_14201);
nor U16002 (N_16002,N_14826,N_14869);
and U16003 (N_16003,N_15771,N_15092);
and U16004 (N_16004,N_14657,N_14858);
xor U16005 (N_16005,N_15593,N_15020);
nor U16006 (N_16006,N_15902,N_14891);
nand U16007 (N_16007,N_15733,N_14428);
nand U16008 (N_16008,N_15428,N_15642);
nor U16009 (N_16009,N_14445,N_15349);
or U16010 (N_16010,N_15309,N_14388);
nand U16011 (N_16011,N_14713,N_15251);
nor U16012 (N_16012,N_15291,N_15795);
xnor U16013 (N_16013,N_14318,N_14410);
nor U16014 (N_16014,N_15609,N_15437);
nor U16015 (N_16015,N_15730,N_15748);
nor U16016 (N_16016,N_15207,N_14553);
nor U16017 (N_16017,N_14880,N_14310);
or U16018 (N_16018,N_14669,N_15624);
xnor U16019 (N_16019,N_14560,N_15169);
nor U16020 (N_16020,N_15659,N_14069);
and U16021 (N_16021,N_15355,N_14502);
nor U16022 (N_16022,N_14223,N_14649);
or U16023 (N_16023,N_14962,N_14889);
or U16024 (N_16024,N_15633,N_14945);
or U16025 (N_16025,N_15611,N_14395);
nor U16026 (N_16026,N_15921,N_15274);
and U16027 (N_16027,N_15107,N_14082);
and U16028 (N_16028,N_14363,N_14016);
or U16029 (N_16029,N_14013,N_15857);
or U16030 (N_16030,N_15629,N_14831);
nand U16031 (N_16031,N_14120,N_15940);
nor U16032 (N_16032,N_14865,N_15438);
or U16033 (N_16033,N_14421,N_15264);
nand U16034 (N_16034,N_14448,N_15380);
nor U16035 (N_16035,N_14026,N_15822);
or U16036 (N_16036,N_14609,N_15884);
xor U16037 (N_16037,N_14579,N_14511);
or U16038 (N_16038,N_15515,N_14357);
and U16039 (N_16039,N_15417,N_15526);
xor U16040 (N_16040,N_14796,N_14813);
nand U16041 (N_16041,N_14054,N_15031);
xnor U16042 (N_16042,N_14036,N_14050);
nor U16043 (N_16043,N_15385,N_14803);
nand U16044 (N_16044,N_15063,N_14847);
xnor U16045 (N_16045,N_15364,N_15821);
and U16046 (N_16046,N_14541,N_15057);
xnor U16047 (N_16047,N_14143,N_14663);
nand U16048 (N_16048,N_15279,N_14968);
nand U16049 (N_16049,N_14984,N_15358);
xnor U16050 (N_16050,N_15075,N_14885);
and U16051 (N_16051,N_15053,N_15718);
and U16052 (N_16052,N_14671,N_14212);
and U16053 (N_16053,N_14301,N_14070);
nand U16054 (N_16054,N_15000,N_14497);
nand U16055 (N_16055,N_15828,N_15338);
and U16056 (N_16056,N_15260,N_14309);
or U16057 (N_16057,N_15021,N_14987);
or U16058 (N_16058,N_15290,N_14126);
and U16059 (N_16059,N_15860,N_15851);
and U16060 (N_16060,N_15017,N_15086);
and U16061 (N_16061,N_15954,N_15323);
and U16062 (N_16062,N_14489,N_15465);
nand U16063 (N_16063,N_14008,N_15707);
nor U16064 (N_16064,N_15994,N_15466);
nand U16065 (N_16065,N_15464,N_14902);
or U16066 (N_16066,N_14398,N_14608);
and U16067 (N_16067,N_14299,N_14720);
xnor U16068 (N_16068,N_14462,N_15145);
or U16069 (N_16069,N_15142,N_15366);
nand U16070 (N_16070,N_15403,N_14386);
or U16071 (N_16071,N_15608,N_14990);
and U16072 (N_16072,N_14561,N_14271);
nand U16073 (N_16073,N_14660,N_14086);
nand U16074 (N_16074,N_14320,N_14898);
and U16075 (N_16075,N_15660,N_15651);
or U16076 (N_16076,N_15909,N_14371);
nor U16077 (N_16077,N_14444,N_14563);
and U16078 (N_16078,N_14806,N_15826);
or U16079 (N_16079,N_14650,N_14235);
and U16080 (N_16080,N_15143,N_14995);
and U16081 (N_16081,N_15335,N_14336);
xnor U16082 (N_16082,N_14273,N_15704);
nand U16083 (N_16083,N_14328,N_15722);
nand U16084 (N_16084,N_14569,N_15590);
nor U16085 (N_16085,N_15227,N_15334);
and U16086 (N_16086,N_15726,N_15667);
nand U16087 (N_16087,N_15875,N_14183);
or U16088 (N_16088,N_14258,N_14172);
xor U16089 (N_16089,N_15002,N_15024);
and U16090 (N_16090,N_15330,N_14789);
xor U16091 (N_16091,N_15044,N_14647);
or U16092 (N_16092,N_15357,N_14246);
nor U16093 (N_16093,N_14966,N_14245);
or U16094 (N_16094,N_15616,N_14930);
and U16095 (N_16095,N_15950,N_14918);
nor U16096 (N_16096,N_14046,N_15777);
nand U16097 (N_16097,N_15454,N_14837);
and U16098 (N_16098,N_15801,N_14754);
and U16099 (N_16099,N_15303,N_14287);
nor U16100 (N_16100,N_14332,N_14999);
and U16101 (N_16101,N_14150,N_14947);
nand U16102 (N_16102,N_14269,N_14236);
nand U16103 (N_16103,N_15635,N_14220);
nor U16104 (N_16104,N_15218,N_15026);
or U16105 (N_16105,N_14573,N_15287);
xnor U16106 (N_16106,N_14056,N_15672);
nor U16107 (N_16107,N_14524,N_14135);
and U16108 (N_16108,N_14280,N_15551);
nand U16109 (N_16109,N_15913,N_14384);
nor U16110 (N_16110,N_14267,N_14334);
or U16111 (N_16111,N_15090,N_15133);
and U16112 (N_16112,N_14331,N_15989);
and U16113 (N_16113,N_14073,N_14676);
nor U16114 (N_16114,N_15679,N_15962);
nor U16115 (N_16115,N_15758,N_15302);
and U16116 (N_16116,N_14510,N_15326);
nand U16117 (N_16117,N_14811,N_15534);
and U16118 (N_16118,N_14696,N_15193);
and U16119 (N_16119,N_14442,N_15240);
nor U16120 (N_16120,N_15621,N_15398);
or U16121 (N_16121,N_15705,N_14751);
or U16122 (N_16122,N_14862,N_15097);
and U16123 (N_16123,N_14459,N_14252);
nor U16124 (N_16124,N_14080,N_14124);
nand U16125 (N_16125,N_15029,N_15890);
nand U16126 (N_16126,N_14666,N_15541);
or U16127 (N_16127,N_14743,N_15981);
or U16128 (N_16128,N_15698,N_14856);
or U16129 (N_16129,N_14980,N_15779);
or U16130 (N_16130,N_15951,N_14830);
nand U16131 (N_16131,N_14540,N_15846);
and U16132 (N_16132,N_14719,N_14043);
nand U16133 (N_16133,N_14735,N_14499);
nor U16134 (N_16134,N_15304,N_15066);
and U16135 (N_16135,N_14290,N_14637);
and U16136 (N_16136,N_14387,N_15829);
or U16137 (N_16137,N_14810,N_14731);
or U16138 (N_16138,N_15373,N_15003);
nor U16139 (N_16139,N_15137,N_15662);
nor U16140 (N_16140,N_15396,N_14965);
and U16141 (N_16141,N_14170,N_14978);
nand U16142 (N_16142,N_14186,N_15037);
nand U16143 (N_16143,N_15160,N_14568);
nand U16144 (N_16144,N_15007,N_14780);
or U16145 (N_16145,N_14169,N_14602);
nor U16146 (N_16146,N_14943,N_15213);
xnor U16147 (N_16147,N_15342,N_15045);
nor U16148 (N_16148,N_14519,N_14030);
nand U16149 (N_16149,N_15391,N_15414);
and U16150 (N_16150,N_14618,N_14748);
or U16151 (N_16151,N_15778,N_14584);
xor U16152 (N_16152,N_15093,N_15471);
nor U16153 (N_16153,N_14634,N_14832);
nand U16154 (N_16154,N_14601,N_14338);
nand U16155 (N_16155,N_15286,N_15201);
and U16156 (N_16156,N_14373,N_15052);
or U16157 (N_16157,N_15501,N_14416);
nor U16158 (N_16158,N_15433,N_15721);
and U16159 (N_16159,N_14023,N_14296);
xnor U16160 (N_16160,N_15088,N_15410);
and U16161 (N_16161,N_15646,N_14304);
xor U16162 (N_16162,N_14821,N_14040);
nor U16163 (N_16163,N_15203,N_15583);
nand U16164 (N_16164,N_14171,N_15475);
nor U16165 (N_16165,N_14079,N_15917);
nand U16166 (N_16166,N_15839,N_15688);
nand U16167 (N_16167,N_14712,N_14533);
nand U16168 (N_16168,N_15379,N_14313);
nand U16169 (N_16169,N_14771,N_15710);
nor U16170 (N_16170,N_15571,N_15650);
nor U16171 (N_16171,N_14033,N_15640);
nor U16172 (N_16172,N_14717,N_14959);
xor U16173 (N_16173,N_15772,N_14059);
or U16174 (N_16174,N_14639,N_14153);
or U16175 (N_16175,N_15156,N_14615);
xor U16176 (N_16176,N_15210,N_15862);
nand U16177 (N_16177,N_14757,N_15485);
nor U16178 (N_16178,N_15337,N_14646);
or U16179 (N_16179,N_15577,N_15062);
nand U16180 (N_16180,N_15736,N_15987);
xor U16181 (N_16181,N_15830,N_15511);
and U16182 (N_16182,N_15663,N_15381);
and U16183 (N_16183,N_14512,N_14842);
or U16184 (N_16184,N_15861,N_14389);
xnor U16185 (N_16185,N_14006,N_14643);
or U16186 (N_16186,N_14193,N_14109);
and U16187 (N_16187,N_15176,N_14229);
or U16188 (N_16188,N_14651,N_14098);
and U16189 (N_16189,N_15209,N_15346);
or U16190 (N_16190,N_14668,N_14161);
nand U16191 (N_16191,N_14545,N_15897);
nand U16192 (N_16192,N_14544,N_15114);
or U16193 (N_16193,N_14931,N_15171);
and U16194 (N_16194,N_14430,N_14924);
nand U16195 (N_16195,N_15077,N_15301);
nand U16196 (N_16196,N_15390,N_14450);
and U16197 (N_16197,N_15903,N_15266);
nor U16198 (N_16198,N_14934,N_15386);
nor U16199 (N_16199,N_15675,N_14066);
or U16200 (N_16200,N_14706,N_15200);
nand U16201 (N_16201,N_14525,N_15299);
nor U16202 (N_16202,N_14325,N_15537);
and U16203 (N_16203,N_14225,N_14482);
and U16204 (N_16204,N_15181,N_15411);
and U16205 (N_16205,N_15673,N_15879);
xnor U16206 (N_16206,N_14045,N_15079);
nor U16207 (N_16207,N_15910,N_15329);
or U16208 (N_16208,N_15558,N_14372);
nand U16209 (N_16209,N_14722,N_14913);
nor U16210 (N_16210,N_14928,N_14173);
or U16211 (N_16211,N_14298,N_15850);
nor U16212 (N_16212,N_15306,N_15360);
and U16213 (N_16213,N_14094,N_14944);
or U16214 (N_16214,N_14460,N_15841);
and U16215 (N_16215,N_15854,N_15775);
and U16216 (N_16216,N_15770,N_15750);
and U16217 (N_16217,N_14973,N_14578);
nor U16218 (N_16218,N_14431,N_14951);
nand U16219 (N_16219,N_14204,N_14749);
or U16220 (N_16220,N_14805,N_14213);
nor U16221 (N_16221,N_14209,N_15574);
nor U16222 (N_16222,N_15192,N_14085);
or U16223 (N_16223,N_15654,N_14675);
nor U16224 (N_16224,N_14972,N_15333);
nor U16225 (N_16225,N_15056,N_15121);
nand U16226 (N_16226,N_14656,N_14382);
and U16227 (N_16227,N_15564,N_14134);
and U16228 (N_16228,N_15076,N_14443);
or U16229 (N_16229,N_14716,N_14364);
xnor U16230 (N_16230,N_14516,N_15588);
and U16231 (N_16231,N_14490,N_15996);
nand U16232 (N_16232,N_14255,N_14142);
and U16233 (N_16233,N_15273,N_14432);
nor U16234 (N_16234,N_14768,N_15392);
nor U16235 (N_16235,N_14518,N_15671);
nor U16236 (N_16236,N_14704,N_15528);
nand U16237 (N_16237,N_15489,N_15883);
nand U16238 (N_16238,N_14095,N_15252);
nor U16239 (N_16239,N_15376,N_15116);
and U16240 (N_16240,N_14390,N_15027);
and U16241 (N_16241,N_15999,N_15011);
xor U16242 (N_16242,N_14268,N_14264);
nor U16243 (N_16243,N_14061,N_14836);
xnor U16244 (N_16244,N_14282,N_14721);
and U16245 (N_16245,N_15870,N_15547);
or U16246 (N_16246,N_15891,N_15195);
nand U16247 (N_16247,N_14641,N_15325);
or U16248 (N_16248,N_14306,N_14697);
nand U16249 (N_16249,N_14483,N_15445);
xor U16250 (N_16250,N_14678,N_15948);
nand U16251 (N_16251,N_15047,N_14911);
nor U16252 (N_16252,N_15269,N_14595);
or U16253 (N_16253,N_15022,N_14202);
and U16254 (N_16254,N_14674,N_15233);
nand U16255 (N_16255,N_14597,N_15803);
nand U16256 (N_16256,N_15361,N_15794);
and U16257 (N_16257,N_15229,N_15185);
nor U16258 (N_16258,N_15078,N_15639);
and U16259 (N_16259,N_14509,N_14745);
nand U16260 (N_16260,N_14020,N_14393);
nor U16261 (N_16261,N_15243,N_15556);
or U16262 (N_16262,N_14447,N_14794);
nor U16263 (N_16263,N_15110,N_14871);
nor U16264 (N_16264,N_14791,N_14808);
and U16265 (N_16265,N_14103,N_15250);
nand U16266 (N_16266,N_14396,N_15668);
nand U16267 (N_16267,N_15964,N_15101);
or U16268 (N_16268,N_14542,N_14096);
nand U16269 (N_16269,N_14127,N_15050);
or U16270 (N_16270,N_15565,N_15103);
and U16271 (N_16271,N_14361,N_14698);
nor U16272 (N_16272,N_14740,N_15509);
nor U16273 (N_16273,N_14081,N_14164);
or U16274 (N_16274,N_15271,N_15068);
or U16275 (N_16275,N_14904,N_15741);
nand U16276 (N_16276,N_15261,N_14177);
or U16277 (N_16277,N_15425,N_14224);
nand U16278 (N_16278,N_15833,N_15180);
and U16279 (N_16279,N_14240,N_15628);
nor U16280 (N_16280,N_15277,N_15720);
nor U16281 (N_16281,N_14822,N_15960);
xnor U16282 (N_16282,N_15109,N_15742);
or U16283 (N_16283,N_15530,N_15695);
and U16284 (N_16284,N_14106,N_14146);
xor U16285 (N_16285,N_15106,N_15601);
or U16286 (N_16286,N_14184,N_14218);
nand U16287 (N_16287,N_14041,N_15518);
xor U16288 (N_16288,N_14732,N_14226);
nand U16289 (N_16289,N_14104,N_14607);
nand U16290 (N_16290,N_14162,N_15914);
and U16291 (N_16291,N_14585,N_14496);
or U16292 (N_16292,N_15263,N_14594);
or U16293 (N_16293,N_14158,N_15665);
and U16294 (N_16294,N_14778,N_14707);
or U16295 (N_16295,N_14348,N_15929);
or U16296 (N_16296,N_15389,N_15626);
nand U16297 (N_16297,N_15040,N_14293);
nor U16298 (N_16298,N_15328,N_15265);
nand U16299 (N_16299,N_15774,N_14292);
xor U16300 (N_16300,N_14548,N_14598);
and U16301 (N_16301,N_14974,N_15009);
and U16302 (N_16302,N_14097,N_15899);
nor U16303 (N_16303,N_14724,N_14192);
nor U16304 (N_16304,N_15276,N_15008);
or U16305 (N_16305,N_15932,N_14196);
nor U16306 (N_16306,N_14123,N_15925);
nand U16307 (N_16307,N_14378,N_15887);
nand U16308 (N_16308,N_15164,N_14690);
and U16309 (N_16309,N_14297,N_14039);
nand U16310 (N_16310,N_14956,N_14977);
or U16311 (N_16311,N_15533,N_14997);
nand U16312 (N_16312,N_15767,N_14031);
and U16313 (N_16313,N_14868,N_14329);
and U16314 (N_16314,N_15934,N_15591);
nor U16315 (N_16315,N_15782,N_14374);
nand U16316 (N_16316,N_14804,N_14469);
or U16317 (N_16317,N_15412,N_14322);
and U16318 (N_16318,N_14857,N_15219);
or U16319 (N_16319,N_15457,N_14905);
nor U16320 (N_16320,N_15042,N_14566);
nand U16321 (N_16321,N_14899,N_15566);
nand U16322 (N_16322,N_15488,N_15852);
or U16323 (N_16323,N_15716,N_14466);
nor U16324 (N_16324,N_14687,N_15248);
and U16325 (N_16325,N_15915,N_14018);
and U16326 (N_16326,N_15892,N_15872);
and U16327 (N_16327,N_14714,N_14558);
xnor U16328 (N_16328,N_15791,N_15529);
or U16329 (N_16329,N_15759,N_14938);
or U16330 (N_16330,N_15048,N_14537);
xor U16331 (N_16331,N_15163,N_15237);
nand U16332 (N_16332,N_15641,N_14588);
nor U16333 (N_16333,N_14688,N_15010);
nor U16334 (N_16334,N_14982,N_14993);
xor U16335 (N_16335,N_14185,N_15874);
or U16336 (N_16336,N_15280,N_15568);
or U16337 (N_16337,N_14790,N_15035);
and U16338 (N_16338,N_15815,N_14239);
nand U16339 (N_16339,N_15451,N_15254);
or U16340 (N_16340,N_14750,N_14189);
nand U16341 (N_16341,N_15963,N_15607);
and U16342 (N_16342,N_14691,N_15676);
nor U16343 (N_16343,N_15028,N_15431);
nor U16344 (N_16344,N_14700,N_15844);
and U16345 (N_16345,N_14181,N_15129);
nor U16346 (N_16346,N_15015,N_15498);
and U16347 (N_16347,N_15615,N_14785);
nor U16348 (N_16348,N_14961,N_15943);
or U16349 (N_16349,N_15552,N_14339);
nor U16350 (N_16350,N_15944,N_14488);
and U16351 (N_16351,N_15189,N_14795);
nor U16352 (N_16352,N_15531,N_14200);
nand U16353 (N_16353,N_15563,N_15298);
and U16354 (N_16354,N_14897,N_14640);
nand U16355 (N_16355,N_14479,N_14683);
or U16356 (N_16356,N_14950,N_14565);
and U16357 (N_16357,N_14067,N_14557);
nor U16358 (N_16358,N_14684,N_14385);
and U16359 (N_16359,N_15173,N_14077);
nand U16360 (N_16360,N_15377,N_14405);
or U16361 (N_16361,N_14487,N_15473);
or U16362 (N_16362,N_14344,N_15447);
and U16363 (N_16363,N_15647,N_14180);
nor U16364 (N_16364,N_15599,N_14093);
xor U16365 (N_16365,N_15728,N_15316);
and U16366 (N_16366,N_14621,N_14156);
nand U16367 (N_16367,N_15216,N_15442);
and U16368 (N_16368,N_15649,N_15188);
or U16369 (N_16369,N_15702,N_15873);
nand U16370 (N_16370,N_14729,N_14215);
xor U16371 (N_16371,N_14241,N_15555);
nand U16372 (N_16372,N_15148,N_15634);
nand U16373 (N_16373,N_14927,N_14957);
nor U16374 (N_16374,N_14333,N_15082);
and U16375 (N_16375,N_15920,N_15370);
nand U16376 (N_16376,N_14817,N_15980);
or U16377 (N_16377,N_15345,N_15843);
nand U16378 (N_16378,N_15468,N_14461);
nor U16379 (N_16379,N_14232,N_14251);
or U16380 (N_16380,N_15986,N_15919);
and U16381 (N_16381,N_14219,N_15916);
and U16382 (N_16382,N_15506,N_14397);
xnor U16383 (N_16383,N_15268,N_14010);
nor U16384 (N_16384,N_15524,N_15912);
nor U16385 (N_16385,N_14829,N_14802);
or U16386 (N_16386,N_14315,N_15395);
and U16387 (N_16387,N_15895,N_14379);
and U16388 (N_16388,N_15587,N_15941);
and U16389 (N_16389,N_15401,N_14556);
nand U16390 (N_16390,N_14368,N_14896);
or U16391 (N_16391,N_15939,N_14529);
or U16392 (N_16392,N_15618,N_14876);
nor U16393 (N_16393,N_14636,N_15288);
and U16394 (N_16394,N_15620,N_15926);
nand U16395 (N_16395,N_15091,N_14937);
or U16396 (N_16396,N_14032,N_15018);
and U16397 (N_16397,N_15115,N_15311);
xnor U16398 (N_16398,N_14929,N_15708);
nand U16399 (N_16399,N_15435,N_15074);
xor U16400 (N_16400,N_15384,N_14653);
and U16401 (N_16401,N_15908,N_14128);
and U16402 (N_16402,N_15049,N_14936);
nand U16403 (N_16403,N_15310,N_14424);
or U16404 (N_16404,N_15723,N_14132);
and U16405 (N_16405,N_15423,N_14591);
and U16406 (N_16406,N_15507,N_15762);
nand U16407 (N_16407,N_14839,N_14259);
and U16408 (N_16408,N_15039,N_15727);
nand U16409 (N_16409,N_15322,N_14933);
nor U16410 (N_16410,N_15985,N_14247);
or U16411 (N_16411,N_15835,N_14659);
nand U16412 (N_16412,N_14883,N_15224);
and U16413 (N_16413,N_14702,N_14622);
or U16414 (N_16414,N_14635,N_15735);
nand U16415 (N_16415,N_14816,N_14798);
and U16416 (N_16416,N_14480,N_15906);
or U16417 (N_16417,N_15592,N_15072);
xnor U16418 (N_16418,N_14216,N_14485);
and U16419 (N_16419,N_15836,N_15898);
nand U16420 (N_16420,N_15432,N_15289);
nand U16421 (N_16421,N_15644,N_14559);
or U16422 (N_16422,N_14029,N_14165);
nand U16423 (N_16423,N_15259,N_14491);
nand U16424 (N_16424,N_14715,N_14605);
xor U16425 (N_16425,N_15175,N_14507);
and U16426 (N_16426,N_15073,N_15174);
or U16427 (N_16427,N_14756,N_14890);
and U16428 (N_16428,N_15060,N_14231);
nand U16429 (N_16429,N_15096,N_14726);
xnor U16430 (N_16430,N_14417,N_15973);
or U16431 (N_16431,N_15598,N_14848);
nor U16432 (N_16432,N_15761,N_15832);
nor U16433 (N_16433,N_14900,N_15893);
nand U16434 (N_16434,N_15141,N_15694);
nor U16435 (N_16435,N_15636,N_15749);
and U16436 (N_16436,N_14157,N_14673);
xor U16437 (N_16437,N_15089,N_15363);
or U16438 (N_16438,N_15965,N_14823);
nor U16439 (N_16439,N_15658,N_15560);
and U16440 (N_16440,N_15455,N_14174);
or U16441 (N_16441,N_15128,N_14148);
nand U16442 (N_16442,N_14834,N_15135);
and U16443 (N_16443,N_15788,N_15512);
nand U16444 (N_16444,N_15383,N_15493);
and U16445 (N_16445,N_14088,N_15619);
nand U16446 (N_16446,N_14625,N_14807);
nor U16447 (N_16447,N_14910,N_14577);
or U16448 (N_16448,N_15371,N_14599);
nand U16449 (N_16449,N_15754,N_14818);
nand U16450 (N_16450,N_14501,N_14330);
nand U16451 (N_16451,N_15165,N_15119);
nand U16452 (N_16452,N_14383,N_15610);
nor U16453 (N_16453,N_14147,N_14582);
and U16454 (N_16454,N_14767,N_15623);
nand U16455 (N_16455,N_15789,N_14012);
nand U16456 (N_16456,N_14118,N_14217);
or U16457 (N_16457,N_15307,N_15812);
nand U16458 (N_16458,N_15613,N_15865);
nand U16459 (N_16459,N_15805,N_14612);
nand U16460 (N_16460,N_14176,N_14710);
and U16461 (N_16461,N_15312,N_15664);
nand U16462 (N_16462,N_15808,N_14763);
and U16463 (N_16463,N_15956,N_14270);
and U16464 (N_16464,N_14248,N_15474);
and U16465 (N_16465,N_15111,N_15458);
or U16466 (N_16466,N_14116,N_14841);
and U16467 (N_16467,N_14394,N_14846);
nand U16468 (N_16468,N_15845,N_14038);
and U16469 (N_16469,N_14187,N_14011);
nand U16470 (N_16470,N_14307,N_14346);
and U16471 (N_16471,N_15067,N_14828);
and U16472 (N_16472,N_14952,N_14278);
nor U16473 (N_16473,N_14948,N_15341);
xnor U16474 (N_16474,N_14590,N_15711);
and U16475 (N_16475,N_15627,N_14068);
nor U16476 (N_16476,N_14117,N_14679);
and U16477 (N_16477,N_14295,N_15426);
nand U16478 (N_16478,N_14981,N_15810);
nand U16479 (N_16479,N_15936,N_15559);
xor U16480 (N_16480,N_14755,N_15321);
nand U16481 (N_16481,N_14903,N_14439);
nor U16482 (N_16482,N_14034,N_15990);
nor U16483 (N_16483,N_14414,N_15146);
nor U16484 (N_16484,N_15510,N_14964);
xor U16485 (N_16485,N_15083,N_14210);
or U16486 (N_16486,N_14788,N_15282);
nand U16487 (N_16487,N_15689,N_15234);
nor U16488 (N_16488,N_14576,N_14976);
nand U16489 (N_16489,N_14616,N_15612);
and U16490 (N_16490,N_14454,N_15350);
and U16491 (N_16491,N_15098,N_15004);
nor U16492 (N_16492,N_15519,N_15586);
or U16493 (N_16493,N_15061,N_14058);
or U16494 (N_16494,N_15579,N_14228);
xor U16495 (N_16495,N_14303,N_15959);
or U16496 (N_16496,N_14354,N_15486);
nand U16497 (N_16497,N_15773,N_14703);
and U16498 (N_16498,N_14718,N_15983);
and U16499 (N_16499,N_14272,N_15998);
or U16500 (N_16500,N_14603,N_14492);
nor U16501 (N_16501,N_15525,N_14211);
and U16502 (N_16502,N_14992,N_15427);
and U16503 (N_16503,N_14672,N_14021);
or U16504 (N_16504,N_15924,N_14655);
nor U16505 (N_16505,N_14824,N_14327);
nand U16506 (N_16506,N_14915,N_14835);
and U16507 (N_16507,N_14286,N_15946);
xnor U16508 (N_16508,N_15840,N_14838);
or U16509 (N_16509,N_15172,N_15296);
or U16510 (N_16510,N_15054,N_15766);
nor U16511 (N_16511,N_15479,N_14326);
nand U16512 (N_16512,N_14484,N_15415);
nand U16513 (N_16513,N_14873,N_14110);
nand U16514 (N_16514,N_15480,N_15578);
or U16515 (N_16515,N_14520,N_15005);
or U16516 (N_16516,N_14131,N_14477);
and U16517 (N_16517,N_15215,N_14538);
xnor U16518 (N_16518,N_14581,N_15150);
and U16519 (N_16519,N_15630,N_15600);
or U16520 (N_16520,N_14665,N_14513);
or U16521 (N_16521,N_14670,N_15368);
or U16522 (N_16522,N_15422,N_15545);
nand U16523 (N_16523,N_15542,N_15896);
and U16524 (N_16524,N_14744,N_14705);
nand U16525 (N_16525,N_14630,N_15140);
nand U16526 (N_16526,N_14119,N_15800);
and U16527 (N_16527,N_14906,N_15747);
nor U16528 (N_16528,N_15546,N_14572);
or U16529 (N_16529,N_14478,N_15817);
and U16530 (N_16530,N_15155,N_15751);
and U16531 (N_16531,N_14404,N_14091);
nor U16532 (N_16532,N_15436,N_15809);
and U16533 (N_16533,N_14986,N_15570);
nor U16534 (N_16534,N_15484,N_15904);
or U16535 (N_16535,N_14644,N_15734);
nand U16536 (N_16536,N_15223,N_15538);
nor U16537 (N_16537,N_14628,N_15162);
or U16538 (N_16538,N_15043,N_14453);
nand U16539 (N_16539,N_15041,N_14206);
xnor U16540 (N_16540,N_14574,N_14547);
xor U16541 (N_16541,N_14878,N_15942);
and U16542 (N_16542,N_15970,N_15553);
nand U16543 (N_16543,N_14799,N_15888);
nand U16544 (N_16544,N_15257,N_14122);
nand U16545 (N_16545,N_14604,N_14052);
nor U16546 (N_16546,N_15604,N_15239);
xnor U16547 (N_16547,N_14527,N_14099);
and U16548 (N_16548,N_15961,N_15785);
and U16549 (N_16549,N_15118,N_14872);
or U16550 (N_16550,N_15806,N_15848);
nand U16551 (N_16551,N_15652,N_15167);
nor U16552 (N_16552,N_14552,N_14063);
nor U16553 (N_16553,N_15247,N_14851);
xor U16554 (N_16554,N_14254,N_14515);
nor U16555 (N_16555,N_15849,N_14275);
nor U16556 (N_16556,N_15949,N_15139);
nand U16557 (N_16557,N_14168,N_15369);
or U16558 (N_16558,N_14409,N_14882);
nor U16559 (N_16559,N_15988,N_15729);
nor U16560 (N_16560,N_14113,N_15179);
nor U16561 (N_16561,N_14337,N_14341);
or U16562 (N_16562,N_15557,N_15784);
nor U16563 (N_16563,N_14377,N_15847);
or U16564 (N_16564,N_15440,N_15992);
and U16565 (N_16565,N_14062,N_15933);
and U16566 (N_16566,N_15576,N_14941);
or U16567 (N_16567,N_15450,N_14107);
nand U16568 (N_16568,N_14892,N_15434);
and U16569 (N_16569,N_15543,N_15690);
nor U16570 (N_16570,N_15418,N_14770);
and U16571 (N_16571,N_14190,N_15460);
and U16572 (N_16572,N_14864,N_15409);
or U16573 (N_16573,N_14642,N_15931);
xor U16574 (N_16574,N_15977,N_15449);
and U16575 (N_16575,N_15187,N_14797);
xor U16576 (N_16576,N_14294,N_15997);
or U16577 (N_16577,N_14092,N_15134);
nor U16578 (N_16578,N_14742,N_14786);
nor U16579 (N_16579,N_14761,N_14543);
or U16580 (N_16580,N_14971,N_15947);
or U16581 (N_16581,N_14244,N_15006);
xor U16582 (N_16582,N_14486,N_14689);
or U16583 (N_16583,N_15419,N_15244);
or U16584 (N_16584,N_14053,N_14044);
and U16585 (N_16585,N_14376,N_15144);
nor U16586 (N_16586,N_14108,N_14160);
nand U16587 (N_16587,N_15256,N_15838);
nand U16588 (N_16588,N_15504,N_14495);
nand U16589 (N_16589,N_14288,N_14534);
nand U16590 (N_16590,N_15825,N_14551);
nand U16591 (N_16591,N_15781,N_15340);
nand U16592 (N_16592,N_14693,N_14888);
or U16593 (N_16593,N_14281,N_14633);
or U16594 (N_16594,N_14476,N_15157);
nor U16595 (N_16595,N_15685,N_14266);
nor U16596 (N_16596,N_15452,N_15225);
nor U16597 (N_16597,N_14437,N_14198);
and U16598 (N_16598,N_14523,N_14919);
nand U16599 (N_16599,N_14188,N_14592);
nand U16600 (N_16600,N_14449,N_14370);
or U16601 (N_16601,N_14855,N_15208);
nand U16602 (N_16602,N_15477,N_15231);
or U16603 (N_16603,N_14772,N_15780);
or U16604 (N_16604,N_15697,N_15463);
nand U16605 (N_16605,N_15562,N_14546);
nand U16606 (N_16606,N_15894,N_15126);
and U16607 (N_16607,N_15462,N_15802);
or U16608 (N_16608,N_14392,N_15740);
xor U16609 (N_16609,N_15211,N_14365);
nor U16610 (N_16610,N_15064,N_15297);
or U16611 (N_16611,N_15138,N_14154);
or U16612 (N_16612,N_14926,N_15945);
or U16613 (N_16613,N_15738,N_14844);
and U16614 (N_16614,N_15669,N_15918);
and U16615 (N_16615,N_15953,N_14163);
nand U16616 (N_16616,N_15393,N_14587);
nand U16617 (N_16617,N_14314,N_14658);
and U16618 (N_16618,N_15790,N_15617);
nor U16619 (N_16619,N_14238,N_14289);
and U16620 (N_16620,N_15399,N_14610);
nor U16621 (N_16621,N_15081,N_15153);
nand U16622 (N_16622,N_14129,N_15955);
nor U16623 (N_16623,N_15481,N_15842);
or U16624 (N_16624,N_15603,N_15262);
or U16625 (N_16625,N_15016,N_15127);
nor U16626 (N_16626,N_15717,N_14433);
nand U16627 (N_16627,N_15154,N_15957);
or U16628 (N_16628,N_15214,N_14814);
or U16629 (N_16629,N_14550,N_14182);
nor U16630 (N_16630,N_15285,N_15051);
or U16631 (N_16631,N_14783,N_15293);
nand U16632 (N_16632,N_14276,N_15561);
nand U16633 (N_16633,N_14440,N_15793);
nor U16634 (N_16634,N_15456,N_14921);
nand U16635 (N_16635,N_14422,N_14677);
or U16636 (N_16636,N_15575,N_14852);
and U16637 (N_16637,N_14854,N_14111);
and U16638 (N_16638,N_14342,N_15441);
nor U16639 (N_16639,N_14145,N_15927);
xor U16640 (N_16640,N_14415,N_14692);
and U16641 (N_16641,N_14531,N_14611);
nand U16642 (N_16642,N_14025,N_14014);
or U16643 (N_16643,N_15928,N_14407);
and U16644 (N_16644,N_15597,N_14886);
and U16645 (N_16645,N_14725,N_15152);
or U16646 (N_16646,N_15461,N_15232);
nand U16647 (N_16647,N_15292,N_15585);
xnor U16648 (N_16648,N_15969,N_14746);
or U16649 (N_16649,N_14623,N_14242);
and U16650 (N_16650,N_14850,N_14323);
xnor U16651 (N_16651,N_14411,N_14257);
or U16652 (N_16652,N_15241,N_15532);
nor U16653 (N_16653,N_14535,N_14105);
nand U16654 (N_16654,N_14090,N_15522);
nand U16655 (N_16655,N_15958,N_15573);
nand U16656 (N_16656,N_14249,N_14701);
or U16657 (N_16657,N_14521,N_14237);
nand U16658 (N_16658,N_14753,N_14391);
or U16659 (N_16659,N_15625,N_15681);
nand U16660 (N_16660,N_14435,N_15731);
and U16661 (N_16661,N_15356,N_14367);
and U16662 (N_16662,N_15683,N_15539);
or U16663 (N_16663,N_15347,N_15272);
and U16664 (N_16664,N_15459,N_15055);
nor U16665 (N_16665,N_14819,N_15242);
nand U16666 (N_16666,N_15295,N_15878);
or U16667 (N_16667,N_14347,N_15365);
xnor U16668 (N_16668,N_14925,N_15100);
nor U16669 (N_16669,N_14227,N_15589);
and U16670 (N_16670,N_14709,N_15058);
and U16671 (N_16671,N_14412,N_14057);
nor U16672 (N_16672,N_15827,N_14946);
xor U16673 (N_16673,N_15320,N_15424);
or U16674 (N_16674,N_14632,N_15132);
nor U16675 (N_16675,N_14825,N_14051);
xor U16676 (N_16676,N_14203,N_15972);
or U16677 (N_16677,N_15632,N_15343);
nand U16678 (N_16678,N_15375,N_14463);
nand U16679 (N_16679,N_15757,N_15420);
or U16680 (N_16680,N_15554,N_15478);
nand U16681 (N_16681,N_14600,N_15540);
or U16682 (N_16682,N_14940,N_14812);
nand U16683 (N_16683,N_14465,N_14564);
xor U16684 (N_16684,N_14685,N_15978);
and U16685 (N_16685,N_15182,N_14627);
and U16686 (N_16686,N_14074,N_14526);
nor U16687 (N_16687,N_14481,N_14881);
and U16688 (N_16688,N_14759,N_14782);
nand U16689 (N_16689,N_15655,N_15868);
nand U16690 (N_16690,N_14064,N_15275);
nand U16691 (N_16691,N_15786,N_14567);
and U16692 (N_16692,N_15503,N_14369);
nand U16693 (N_16693,N_15550,N_14849);
and U16694 (N_16694,N_14362,N_15443);
nand U16695 (N_16695,N_14539,N_15099);
xor U16696 (N_16696,N_15059,N_15703);
nor U16697 (N_16697,N_14352,N_14436);
or U16698 (N_16698,N_15643,N_14967);
or U16699 (N_16699,N_15645,N_14549);
or U16700 (N_16700,N_15388,N_15885);
nand U16701 (N_16701,N_15765,N_14274);
nor U16702 (N_16702,N_14208,N_15374);
nand U16703 (N_16703,N_14221,N_15661);
nor U16704 (N_16704,N_14195,N_15674);
or U16705 (N_16705,N_15732,N_14522);
nand U16706 (N_16706,N_15678,N_14472);
xnor U16707 (N_16707,N_14909,N_15858);
nand U16708 (N_16708,N_14350,N_14028);
and U16709 (N_16709,N_14413,N_14654);
nor U16710 (N_16710,N_15637,N_15768);
or U16711 (N_16711,N_14681,N_14914);
or U16712 (N_16712,N_14580,N_14024);
or U16713 (N_16713,N_15158,N_15813);
and U16714 (N_16714,N_14800,N_14988);
or U16715 (N_16715,N_14571,N_15976);
nor U16716 (N_16716,N_15448,N_15714);
xnor U16717 (N_16717,N_15161,N_14989);
and U16718 (N_16718,N_15406,N_14738);
nor U16719 (N_16719,N_14455,N_14159);
and U16720 (N_16720,N_14877,N_14233);
and U16721 (N_16721,N_14399,N_15811);
and U16722 (N_16722,N_14279,N_15353);
and U16723 (N_16723,N_15147,N_14733);
nor U16724 (N_16724,N_15413,N_15787);
and U16725 (N_16725,N_15535,N_14335);
and U16726 (N_16726,N_14002,N_15993);
nand U16727 (N_16727,N_14908,N_15038);
and U16728 (N_16728,N_15979,N_14935);
nor U16729 (N_16729,N_14809,N_14983);
or U16730 (N_16730,N_15467,N_14619);
and U16731 (N_16731,N_14758,N_15966);
and U16732 (N_16732,N_14214,N_14589);
xor U16733 (N_16733,N_14458,N_14317);
nand U16734 (N_16734,N_15974,N_14121);
or U16735 (N_16735,N_15876,N_15084);
nand U16736 (N_16736,N_14764,N_15930);
nand U16737 (N_16737,N_14167,N_14860);
nor U16738 (N_16738,N_14820,N_15184);
nor U16739 (N_16739,N_15869,N_14166);
and U16740 (N_16740,N_15190,N_14958);
nand U16741 (N_16741,N_15102,N_14312);
nand U16742 (N_16742,N_14979,N_15982);
and U16743 (N_16743,N_14500,N_14723);
nand U16744 (N_16744,N_14815,N_15255);
or U16745 (N_16745,N_14923,N_14949);
nand U16746 (N_16746,N_14631,N_15496);
nand U16747 (N_16747,N_14102,N_15238);
and U16748 (N_16748,N_14149,N_15816);
nand U16749 (N_16749,N_15378,N_14760);
xor U16750 (N_16750,N_14101,N_14076);
nor U16751 (N_16751,N_14356,N_15814);
nor U16752 (N_16752,N_15952,N_15344);
nand U16753 (N_16753,N_14353,N_14284);
or U16754 (N_16754,N_15866,N_15606);
and U16755 (N_16755,N_14060,N_14321);
nor U16756 (N_16756,N_14762,N_15351);
or U16757 (N_16757,N_15544,N_14253);
and U16758 (N_16758,N_15567,N_15820);
nand U16759 (N_16759,N_14452,N_15764);
or U16760 (N_16760,N_14833,N_15253);
or U16761 (N_16761,N_14570,N_15907);
or U16762 (N_16762,N_14699,N_14922);
nor U16763 (N_16763,N_14207,N_15105);
or U16764 (N_16764,N_14359,N_15104);
and U16765 (N_16765,N_14769,N_14985);
nand U16766 (N_16766,N_15682,N_15756);
or U16767 (N_16767,N_14451,N_14504);
nor U16768 (N_16768,N_15191,N_15905);
or U16769 (N_16769,N_15594,N_15476);
or U16770 (N_16770,N_14994,N_15117);
nor U16771 (N_16771,N_15514,N_14112);
and U16772 (N_16772,N_15753,N_15222);
or U16773 (N_16773,N_14355,N_15025);
nor U16774 (N_16774,N_15236,N_15911);
nand U16775 (N_16775,N_14528,N_14308);
nand U16776 (N_16776,N_15938,N_14100);
nand U16777 (N_16777,N_15725,N_14137);
and U16778 (N_16778,N_14536,N_15886);
nor U16779 (N_16779,N_15687,N_15968);
nand U16780 (N_16780,N_15249,N_15666);
nor U16781 (N_16781,N_14205,N_15019);
or U16782 (N_16782,N_14747,N_15743);
and U16783 (N_16783,N_15653,N_14801);
nand U16784 (N_16784,N_15439,N_15183);
and U16785 (N_16785,N_14517,N_14613);
nor U16786 (N_16786,N_14261,N_14340);
or U16787 (N_16787,N_14583,N_15070);
nand U16788 (N_16788,N_15023,N_14140);
nor U16789 (N_16789,N_14065,N_14381);
nand U16790 (N_16790,N_14360,N_14423);
nand U16791 (N_16791,N_14863,N_14875);
nor U16792 (N_16792,N_15497,N_14727);
and U16793 (N_16793,N_15001,N_15245);
xnor U16794 (N_16794,N_15715,N_14175);
nand U16795 (N_16795,N_14575,N_14624);
xnor U16796 (N_16796,N_14115,N_14954);
nand U16797 (N_16797,N_15030,N_15487);
nor U16798 (N_16798,N_15746,N_14004);
nor U16799 (N_16799,N_14055,N_15034);
nand U16800 (N_16800,N_15394,N_14506);
or U16801 (N_16801,N_15071,N_14774);
and U16802 (N_16802,N_14464,N_14305);
or U16803 (N_16803,N_14629,N_15159);
nor U16804 (N_16804,N_14017,N_15799);
or U16805 (N_16805,N_14645,N_14285);
nor U16806 (N_16806,N_14427,N_15517);
or U16807 (N_16807,N_14859,N_14861);
nand U16808 (N_16808,N_14457,N_15186);
and U16809 (N_16809,N_14136,N_15402);
nor U16810 (N_16810,N_14920,N_15446);
and U16811 (N_16811,N_14456,N_14402);
and U16812 (N_16812,N_15470,N_15124);
xor U16813 (N_16813,N_15429,N_14007);
nand U16814 (N_16814,N_14708,N_15324);
or U16815 (N_16815,N_14845,N_15331);
or U16816 (N_16816,N_15709,N_15724);
and U16817 (N_16817,N_15513,N_15125);
xnor U16818 (N_16818,N_15336,N_15228);
or U16819 (N_16819,N_14001,N_15700);
nor U16820 (N_16820,N_15278,N_14776);
nand U16821 (N_16821,N_15036,N_15548);
nand U16822 (N_16822,N_15212,N_15648);
and U16823 (N_16823,N_14728,N_14853);
nor U16824 (N_16824,N_15492,N_15739);
nand U16825 (N_16825,N_15226,N_15776);
nand U16826 (N_16826,N_14083,N_15168);
nand U16827 (N_16827,N_15798,N_15701);
nand U16828 (N_16828,N_14916,N_15080);
and U16829 (N_16829,N_14765,N_14250);
or U16830 (N_16830,N_14784,N_14638);
nor U16831 (N_16831,N_14695,N_15315);
nand U16832 (N_16832,N_14620,N_14019);
and U16833 (N_16833,N_15284,N_15991);
and U16834 (N_16834,N_14895,N_14498);
nand U16835 (N_16835,N_14400,N_14474);
xor U16836 (N_16836,N_14262,N_14737);
nor U16837 (N_16837,N_14152,N_15122);
nor U16838 (N_16838,N_14667,N_15871);
and U16839 (N_16839,N_14554,N_14626);
and U16840 (N_16840,N_15217,N_15831);
nor U16841 (N_16841,N_15752,N_15706);
and U16842 (N_16842,N_15677,N_15719);
and U16843 (N_16843,N_15900,N_15281);
nand U16844 (N_16844,N_14555,N_14441);
and U16845 (N_16845,N_15614,N_14827);
or U16846 (N_16846,N_14773,N_14901);
and U16847 (N_16847,N_14009,N_14197);
nand U16848 (N_16848,N_15205,N_14867);
nand U16849 (N_16849,N_14078,N_14766);
nand U16850 (N_16850,N_14711,N_15490);
nand U16851 (N_16851,N_15638,N_14503);
nand U16852 (N_16852,N_14141,N_15065);
and U16853 (N_16853,N_15580,N_15108);
nor U16854 (N_16854,N_14446,N_15359);
and U16855 (N_16855,N_14505,N_15755);
or U16856 (N_16856,N_14408,N_15408);
or U16857 (N_16857,N_14263,N_14256);
and U16858 (N_16858,N_15744,N_15483);
and U16859 (N_16859,N_15760,N_14302);
and U16860 (N_16860,N_15508,N_15837);
or U16861 (N_16861,N_15763,N_15975);
xor U16862 (N_16862,N_14752,N_15712);
nand U16863 (N_16863,N_15584,N_14230);
xor U16864 (N_16864,N_14035,N_15405);
or U16865 (N_16865,N_14779,N_14596);
nor U16866 (N_16866,N_14680,N_15859);
or U16867 (N_16867,N_14932,N_15258);
or U16868 (N_16868,N_14349,N_15984);
and U16869 (N_16869,N_14005,N_14027);
and U16870 (N_16870,N_15527,N_14114);
nor U16871 (N_16871,N_14260,N_15516);
nand U16872 (N_16872,N_15094,N_14151);
nand U16873 (N_16873,N_14048,N_15069);
xnor U16874 (N_16874,N_14781,N_14996);
nand U16875 (N_16875,N_15283,N_14562);
or U16876 (N_16876,N_15194,N_14955);
nor U16877 (N_16877,N_14291,N_14234);
nand U16878 (N_16878,N_14662,N_15348);
nand U16879 (N_16879,N_15792,N_14942);
nand U16880 (N_16880,N_15656,N_14139);
or U16881 (N_16881,N_14917,N_15313);
and U16882 (N_16882,N_15220,N_14138);
nor U16883 (N_16883,N_15367,N_15696);
xnor U16884 (N_16884,N_15482,N_15505);
or U16885 (N_16885,N_14071,N_14969);
nand U16886 (N_16886,N_14998,N_15317);
nor U16887 (N_16887,N_15523,N_14316);
nand U16888 (N_16888,N_14277,N_15469);
or U16889 (N_16889,N_15300,N_15318);
or U16890 (N_16890,N_15294,N_15494);
nor U16891 (N_16891,N_15495,N_15536);
nor U16892 (N_16892,N_14366,N_15499);
xnor U16893 (N_16893,N_14037,N_14343);
nand U16894 (N_16894,N_14493,N_15881);
or U16895 (N_16895,N_14467,N_14606);
nand U16896 (N_16896,N_14530,N_14191);
or U16897 (N_16897,N_14429,N_15270);
and U16898 (N_16898,N_14015,N_15877);
or U16899 (N_16899,N_14351,N_15834);
nand U16900 (N_16900,N_15131,N_15197);
or U16901 (N_16901,N_15500,N_15332);
nand U16902 (N_16902,N_15769,N_14840);
and U16903 (N_16903,N_14425,N_14907);
and U16904 (N_16904,N_15797,N_14022);
nand U16905 (N_16905,N_15319,N_15602);
nor U16906 (N_16906,N_14617,N_14866);
nand U16907 (N_16907,N_15995,N_14155);
nand U16908 (N_16908,N_15889,N_15521);
or U16909 (N_16909,N_15631,N_15937);
nor U16910 (N_16910,N_14243,N_15404);
nor U16911 (N_16911,N_14047,N_15686);
xor U16912 (N_16912,N_14793,N_14426);
and U16913 (N_16913,N_14893,N_15314);
and U16914 (N_16914,N_14075,N_14300);
and U16915 (N_16915,N_14741,N_14265);
nand U16916 (N_16916,N_15605,N_15397);
nand U16917 (N_16917,N_14593,N_14960);
nand U16918 (N_16918,N_15967,N_15196);
nand U16919 (N_16919,N_15823,N_14912);
or U16920 (N_16920,N_14661,N_15202);
nand U16921 (N_16921,N_15549,N_15581);
and U16922 (N_16922,N_15387,N_15818);
and U16923 (N_16923,N_14358,N_14125);
or U16924 (N_16924,N_15362,N_14475);
or U16925 (N_16925,N_14199,N_15199);
nand U16926 (N_16926,N_15198,N_14514);
nor U16927 (N_16927,N_14380,N_15804);
or U16928 (N_16928,N_15693,N_15382);
or U16929 (N_16929,N_15796,N_14087);
and U16930 (N_16930,N_15864,N_15657);
nor U16931 (N_16931,N_15853,N_14222);
xor U16932 (N_16932,N_14471,N_14953);
and U16933 (N_16933,N_14420,N_15680);
or U16934 (N_16934,N_15012,N_15308);
nand U16935 (N_16935,N_15204,N_14664);
and U16936 (N_16936,N_15327,N_15130);
nand U16937 (N_16937,N_14532,N_15691);
nand U16938 (N_16938,N_15882,N_15923);
xnor U16939 (N_16939,N_14401,N_15819);
and U16940 (N_16940,N_15014,N_15595);
nor U16941 (N_16941,N_15235,N_14000);
xor U16942 (N_16942,N_15622,N_14730);
xor U16943 (N_16943,N_15136,N_14319);
nand U16944 (N_16944,N_14963,N_14434);
nor U16945 (N_16945,N_15354,N_15444);
nor U16946 (N_16946,N_14879,N_15971);
nand U16947 (N_16947,N_15230,N_14894);
and U16948 (N_16948,N_14884,N_15901);
or U16949 (N_16949,N_14991,N_14792);
and U16950 (N_16950,N_14694,N_15922);
xnor U16951 (N_16951,N_14494,N_14682);
nand U16952 (N_16952,N_14283,N_15935);
xor U16953 (N_16953,N_15339,N_15692);
and U16954 (N_16954,N_14179,N_15596);
nand U16955 (N_16955,N_15178,N_15745);
nor U16956 (N_16956,N_14975,N_15582);
nor U16957 (N_16957,N_15046,N_15472);
nor U16958 (N_16958,N_14375,N_14049);
nand U16959 (N_16959,N_14734,N_14003);
or U16960 (N_16960,N_14419,N_15407);
xnor U16961 (N_16961,N_14777,N_15352);
or U16962 (N_16962,N_15085,N_15305);
nor U16963 (N_16963,N_14887,N_15112);
nor U16964 (N_16964,N_14470,N_14406);
or U16965 (N_16965,N_15856,N_15177);
and U16966 (N_16966,N_14084,N_15416);
nor U16967 (N_16967,N_14345,N_15166);
nor U16968 (N_16968,N_15572,N_14130);
nor U16969 (N_16969,N_15095,N_15087);
xnor U16970 (N_16970,N_15400,N_15421);
nand U16971 (N_16971,N_15867,N_15520);
or U16972 (N_16972,N_14178,N_15123);
or U16973 (N_16973,N_15032,N_15149);
nand U16974 (N_16974,N_15267,N_15863);
and U16975 (N_16975,N_14473,N_15880);
or U16976 (N_16976,N_15120,N_14736);
or U16977 (N_16977,N_14144,N_15855);
and U16978 (N_16978,N_15684,N_15170);
or U16979 (N_16979,N_14133,N_15569);
xnor U16980 (N_16980,N_14311,N_15670);
nor U16981 (N_16981,N_14648,N_14324);
or U16982 (N_16982,N_14970,N_14403);
xnor U16983 (N_16983,N_14939,N_15783);
or U16984 (N_16984,N_14438,N_15699);
or U16985 (N_16985,N_15372,N_14775);
or U16986 (N_16986,N_15491,N_15206);
nor U16987 (N_16987,N_15737,N_15713);
or U16988 (N_16988,N_15824,N_15113);
or U16989 (N_16989,N_14586,N_15807);
xor U16990 (N_16990,N_14194,N_14652);
xor U16991 (N_16991,N_14870,N_14843);
nor U16992 (N_16992,N_14686,N_14042);
nand U16993 (N_16993,N_14739,N_15221);
xor U16994 (N_16994,N_15013,N_14614);
xnor U16995 (N_16995,N_14418,N_14072);
and U16996 (N_16996,N_14089,N_15453);
xnor U16997 (N_16997,N_14468,N_14787);
xnor U16998 (N_16998,N_15151,N_15430);
nand U16999 (N_16999,N_14874,N_15502);
nand U17000 (N_17000,N_14957,N_14931);
nor U17001 (N_17001,N_15051,N_14492);
or U17002 (N_17002,N_14871,N_14925);
nand U17003 (N_17003,N_14671,N_14371);
nand U17004 (N_17004,N_15904,N_15576);
xor U17005 (N_17005,N_14429,N_15481);
and U17006 (N_17006,N_15027,N_14359);
nor U17007 (N_17007,N_15767,N_14869);
nand U17008 (N_17008,N_14873,N_14468);
or U17009 (N_17009,N_15794,N_14251);
nor U17010 (N_17010,N_15385,N_14556);
or U17011 (N_17011,N_14771,N_15925);
nor U17012 (N_17012,N_14748,N_14329);
or U17013 (N_17013,N_14060,N_14605);
and U17014 (N_17014,N_14988,N_15381);
and U17015 (N_17015,N_14843,N_15299);
or U17016 (N_17016,N_14076,N_15843);
xor U17017 (N_17017,N_14365,N_15760);
nor U17018 (N_17018,N_15922,N_15493);
nor U17019 (N_17019,N_14773,N_15908);
nor U17020 (N_17020,N_14012,N_15510);
nand U17021 (N_17021,N_14537,N_15746);
and U17022 (N_17022,N_14036,N_14986);
and U17023 (N_17023,N_15468,N_14180);
xnor U17024 (N_17024,N_15760,N_15120);
nor U17025 (N_17025,N_15579,N_14140);
nand U17026 (N_17026,N_14423,N_14913);
nand U17027 (N_17027,N_15582,N_14366);
xor U17028 (N_17028,N_14134,N_14816);
and U17029 (N_17029,N_15569,N_15116);
and U17030 (N_17030,N_14107,N_14021);
nor U17031 (N_17031,N_14122,N_15740);
nand U17032 (N_17032,N_15697,N_14547);
nor U17033 (N_17033,N_14761,N_14544);
nand U17034 (N_17034,N_14323,N_14479);
and U17035 (N_17035,N_14181,N_15715);
xnor U17036 (N_17036,N_14881,N_15569);
nor U17037 (N_17037,N_15176,N_15556);
nand U17038 (N_17038,N_15341,N_14694);
and U17039 (N_17039,N_14205,N_14196);
nor U17040 (N_17040,N_14247,N_14687);
or U17041 (N_17041,N_14505,N_15922);
xor U17042 (N_17042,N_15455,N_14863);
nand U17043 (N_17043,N_15797,N_15684);
nor U17044 (N_17044,N_14585,N_15229);
or U17045 (N_17045,N_15851,N_14064);
xor U17046 (N_17046,N_15234,N_15974);
nor U17047 (N_17047,N_14884,N_15912);
or U17048 (N_17048,N_14481,N_14987);
nor U17049 (N_17049,N_14142,N_14136);
or U17050 (N_17050,N_15370,N_14245);
nand U17051 (N_17051,N_15322,N_15903);
or U17052 (N_17052,N_14750,N_15019);
or U17053 (N_17053,N_14995,N_15684);
nor U17054 (N_17054,N_15110,N_14750);
nand U17055 (N_17055,N_15839,N_15601);
nand U17056 (N_17056,N_14323,N_15519);
nor U17057 (N_17057,N_15816,N_15589);
nor U17058 (N_17058,N_14383,N_14009);
xnor U17059 (N_17059,N_15974,N_14160);
or U17060 (N_17060,N_15945,N_14871);
or U17061 (N_17061,N_14883,N_14871);
and U17062 (N_17062,N_14912,N_14451);
nand U17063 (N_17063,N_15704,N_14323);
nand U17064 (N_17064,N_15090,N_15907);
nand U17065 (N_17065,N_14046,N_14778);
nand U17066 (N_17066,N_15499,N_15606);
nor U17067 (N_17067,N_15589,N_15655);
nand U17068 (N_17068,N_15911,N_14332);
nand U17069 (N_17069,N_15164,N_15157);
and U17070 (N_17070,N_15954,N_15956);
and U17071 (N_17071,N_15413,N_14667);
or U17072 (N_17072,N_15146,N_14840);
nor U17073 (N_17073,N_15793,N_14731);
and U17074 (N_17074,N_15060,N_14651);
nor U17075 (N_17075,N_14082,N_15132);
and U17076 (N_17076,N_14536,N_14106);
nand U17077 (N_17077,N_15969,N_15756);
nand U17078 (N_17078,N_14346,N_14874);
or U17079 (N_17079,N_15376,N_14619);
or U17080 (N_17080,N_14514,N_15731);
or U17081 (N_17081,N_15433,N_14695);
nor U17082 (N_17082,N_14839,N_14342);
and U17083 (N_17083,N_15926,N_15063);
nand U17084 (N_17084,N_15557,N_15516);
or U17085 (N_17085,N_15183,N_15431);
and U17086 (N_17086,N_15985,N_14211);
nor U17087 (N_17087,N_14146,N_14258);
nor U17088 (N_17088,N_15804,N_15439);
and U17089 (N_17089,N_15302,N_14390);
nand U17090 (N_17090,N_15406,N_14097);
nor U17091 (N_17091,N_14528,N_15221);
nor U17092 (N_17092,N_14718,N_14004);
nor U17093 (N_17093,N_14735,N_15645);
and U17094 (N_17094,N_14048,N_14213);
or U17095 (N_17095,N_14343,N_15897);
nand U17096 (N_17096,N_14361,N_14878);
or U17097 (N_17097,N_14954,N_15767);
nor U17098 (N_17098,N_14560,N_15775);
or U17099 (N_17099,N_15970,N_15007);
nor U17100 (N_17100,N_14837,N_14964);
or U17101 (N_17101,N_15547,N_14728);
and U17102 (N_17102,N_14384,N_15471);
nor U17103 (N_17103,N_15129,N_14262);
and U17104 (N_17104,N_15629,N_15742);
xor U17105 (N_17105,N_14347,N_15884);
nor U17106 (N_17106,N_14624,N_15452);
nand U17107 (N_17107,N_15718,N_15368);
nor U17108 (N_17108,N_14327,N_15905);
nand U17109 (N_17109,N_14938,N_15528);
nand U17110 (N_17110,N_14739,N_15017);
and U17111 (N_17111,N_14192,N_14364);
xor U17112 (N_17112,N_14759,N_14626);
and U17113 (N_17113,N_14871,N_14918);
nor U17114 (N_17114,N_14070,N_14462);
nand U17115 (N_17115,N_15927,N_15198);
or U17116 (N_17116,N_15312,N_15232);
nand U17117 (N_17117,N_14474,N_15124);
nor U17118 (N_17118,N_14915,N_15196);
nand U17119 (N_17119,N_14843,N_15845);
or U17120 (N_17120,N_15082,N_15900);
nor U17121 (N_17121,N_15196,N_15978);
nor U17122 (N_17122,N_15690,N_14573);
and U17123 (N_17123,N_15367,N_14660);
nand U17124 (N_17124,N_14663,N_14845);
nor U17125 (N_17125,N_15347,N_14476);
or U17126 (N_17126,N_14496,N_14142);
xor U17127 (N_17127,N_14636,N_14893);
or U17128 (N_17128,N_15482,N_14905);
or U17129 (N_17129,N_14937,N_15183);
nor U17130 (N_17130,N_15368,N_14092);
nor U17131 (N_17131,N_14719,N_15672);
and U17132 (N_17132,N_15630,N_15088);
or U17133 (N_17133,N_15487,N_15326);
and U17134 (N_17134,N_15809,N_15457);
or U17135 (N_17135,N_14099,N_15528);
nor U17136 (N_17136,N_14073,N_14016);
xor U17137 (N_17137,N_14987,N_14509);
or U17138 (N_17138,N_15312,N_14148);
xor U17139 (N_17139,N_14128,N_14198);
nor U17140 (N_17140,N_15078,N_14441);
or U17141 (N_17141,N_15121,N_15184);
and U17142 (N_17142,N_15152,N_15031);
nand U17143 (N_17143,N_14194,N_15006);
or U17144 (N_17144,N_15786,N_15638);
nor U17145 (N_17145,N_15235,N_15051);
nand U17146 (N_17146,N_14702,N_15639);
nor U17147 (N_17147,N_15388,N_15882);
and U17148 (N_17148,N_15940,N_14815);
nor U17149 (N_17149,N_14326,N_15060);
or U17150 (N_17150,N_15321,N_14448);
xor U17151 (N_17151,N_14456,N_15717);
or U17152 (N_17152,N_15517,N_14300);
and U17153 (N_17153,N_15964,N_15035);
and U17154 (N_17154,N_15974,N_15732);
nor U17155 (N_17155,N_15350,N_15670);
or U17156 (N_17156,N_14738,N_15086);
and U17157 (N_17157,N_14395,N_15070);
nand U17158 (N_17158,N_14767,N_15057);
nor U17159 (N_17159,N_14479,N_15424);
nand U17160 (N_17160,N_15562,N_15020);
nand U17161 (N_17161,N_14276,N_14150);
nor U17162 (N_17162,N_14809,N_15679);
and U17163 (N_17163,N_15628,N_15016);
nand U17164 (N_17164,N_14340,N_14539);
or U17165 (N_17165,N_14421,N_15851);
and U17166 (N_17166,N_15655,N_15552);
nand U17167 (N_17167,N_15148,N_15061);
nor U17168 (N_17168,N_15485,N_15512);
or U17169 (N_17169,N_14714,N_14052);
nand U17170 (N_17170,N_15651,N_15166);
or U17171 (N_17171,N_15505,N_15350);
nand U17172 (N_17172,N_14507,N_15129);
xor U17173 (N_17173,N_15145,N_15116);
nor U17174 (N_17174,N_15429,N_15029);
nand U17175 (N_17175,N_14787,N_14606);
or U17176 (N_17176,N_15035,N_14645);
xor U17177 (N_17177,N_15698,N_15550);
nor U17178 (N_17178,N_15090,N_14734);
and U17179 (N_17179,N_15913,N_15516);
nand U17180 (N_17180,N_15120,N_14356);
and U17181 (N_17181,N_15551,N_14079);
nand U17182 (N_17182,N_15414,N_14904);
or U17183 (N_17183,N_14144,N_14250);
nor U17184 (N_17184,N_14129,N_15587);
or U17185 (N_17185,N_15554,N_15222);
nand U17186 (N_17186,N_15235,N_15695);
nor U17187 (N_17187,N_14453,N_15255);
and U17188 (N_17188,N_15254,N_15857);
or U17189 (N_17189,N_15408,N_14236);
or U17190 (N_17190,N_15391,N_14220);
nor U17191 (N_17191,N_15182,N_14726);
nor U17192 (N_17192,N_14079,N_15200);
nand U17193 (N_17193,N_15273,N_15537);
or U17194 (N_17194,N_15328,N_15107);
nor U17195 (N_17195,N_14472,N_15936);
or U17196 (N_17196,N_14873,N_15450);
xnor U17197 (N_17197,N_15244,N_15755);
and U17198 (N_17198,N_15567,N_15824);
or U17199 (N_17199,N_14184,N_14151);
xnor U17200 (N_17200,N_14681,N_15355);
or U17201 (N_17201,N_15211,N_14127);
and U17202 (N_17202,N_15356,N_15331);
nor U17203 (N_17203,N_15712,N_15691);
and U17204 (N_17204,N_15398,N_15439);
nand U17205 (N_17205,N_15866,N_14031);
nand U17206 (N_17206,N_14210,N_14190);
or U17207 (N_17207,N_15184,N_14298);
and U17208 (N_17208,N_14832,N_14592);
or U17209 (N_17209,N_15617,N_14034);
or U17210 (N_17210,N_15597,N_14699);
nand U17211 (N_17211,N_14188,N_15241);
nor U17212 (N_17212,N_14150,N_14650);
and U17213 (N_17213,N_14937,N_15061);
nand U17214 (N_17214,N_14460,N_15683);
xnor U17215 (N_17215,N_14112,N_15139);
or U17216 (N_17216,N_14548,N_15469);
or U17217 (N_17217,N_15091,N_14549);
and U17218 (N_17218,N_14105,N_14348);
or U17219 (N_17219,N_14930,N_14553);
or U17220 (N_17220,N_14993,N_14396);
nand U17221 (N_17221,N_14334,N_14675);
xnor U17222 (N_17222,N_14249,N_14644);
and U17223 (N_17223,N_15529,N_14570);
xor U17224 (N_17224,N_14708,N_14165);
and U17225 (N_17225,N_14161,N_14717);
nor U17226 (N_17226,N_14349,N_14433);
or U17227 (N_17227,N_15913,N_15081);
and U17228 (N_17228,N_14512,N_14701);
and U17229 (N_17229,N_14407,N_15158);
nand U17230 (N_17230,N_15253,N_15223);
and U17231 (N_17231,N_14849,N_15451);
nand U17232 (N_17232,N_14261,N_14581);
nor U17233 (N_17233,N_14824,N_14443);
and U17234 (N_17234,N_15867,N_14775);
nor U17235 (N_17235,N_15297,N_15812);
or U17236 (N_17236,N_14597,N_15282);
and U17237 (N_17237,N_14578,N_14622);
nand U17238 (N_17238,N_15221,N_14774);
xnor U17239 (N_17239,N_14761,N_15685);
nor U17240 (N_17240,N_14493,N_14671);
or U17241 (N_17241,N_14441,N_15188);
or U17242 (N_17242,N_15350,N_14580);
and U17243 (N_17243,N_15445,N_14750);
nand U17244 (N_17244,N_14671,N_14920);
and U17245 (N_17245,N_15322,N_15479);
xnor U17246 (N_17246,N_15508,N_15709);
nor U17247 (N_17247,N_14063,N_14081);
nand U17248 (N_17248,N_15139,N_14595);
or U17249 (N_17249,N_14003,N_14897);
xor U17250 (N_17250,N_15833,N_15596);
nand U17251 (N_17251,N_15526,N_15171);
and U17252 (N_17252,N_14835,N_15005);
or U17253 (N_17253,N_15425,N_14394);
nand U17254 (N_17254,N_14278,N_14175);
or U17255 (N_17255,N_15539,N_15122);
and U17256 (N_17256,N_15146,N_14820);
xnor U17257 (N_17257,N_14086,N_14999);
or U17258 (N_17258,N_14837,N_14066);
nand U17259 (N_17259,N_14920,N_15150);
nand U17260 (N_17260,N_14845,N_15783);
or U17261 (N_17261,N_14997,N_15733);
nand U17262 (N_17262,N_14763,N_15335);
nor U17263 (N_17263,N_15247,N_14867);
nor U17264 (N_17264,N_15039,N_15342);
nand U17265 (N_17265,N_15636,N_14774);
nand U17266 (N_17266,N_14658,N_15083);
nand U17267 (N_17267,N_14530,N_14995);
nor U17268 (N_17268,N_14821,N_15556);
or U17269 (N_17269,N_14894,N_15355);
and U17270 (N_17270,N_14906,N_14246);
or U17271 (N_17271,N_14275,N_14347);
nand U17272 (N_17272,N_14684,N_15278);
and U17273 (N_17273,N_15237,N_14157);
xor U17274 (N_17274,N_14151,N_14281);
or U17275 (N_17275,N_15763,N_14754);
and U17276 (N_17276,N_14312,N_15166);
or U17277 (N_17277,N_14524,N_14920);
or U17278 (N_17278,N_14329,N_15753);
nor U17279 (N_17279,N_15994,N_14956);
nor U17280 (N_17280,N_15037,N_15736);
nor U17281 (N_17281,N_15359,N_15119);
nor U17282 (N_17282,N_15770,N_15644);
nand U17283 (N_17283,N_14748,N_14133);
or U17284 (N_17284,N_15705,N_14997);
or U17285 (N_17285,N_15193,N_15415);
xnor U17286 (N_17286,N_14879,N_15185);
or U17287 (N_17287,N_14296,N_15380);
and U17288 (N_17288,N_15235,N_15654);
and U17289 (N_17289,N_15052,N_14534);
nor U17290 (N_17290,N_14784,N_15183);
or U17291 (N_17291,N_15835,N_15996);
nor U17292 (N_17292,N_14183,N_15924);
nor U17293 (N_17293,N_15564,N_14738);
or U17294 (N_17294,N_15223,N_14303);
nand U17295 (N_17295,N_14646,N_15875);
xnor U17296 (N_17296,N_15680,N_15752);
and U17297 (N_17297,N_15468,N_15111);
nor U17298 (N_17298,N_14599,N_15957);
xor U17299 (N_17299,N_14431,N_15313);
nor U17300 (N_17300,N_14172,N_14293);
nor U17301 (N_17301,N_14913,N_14535);
and U17302 (N_17302,N_15100,N_14283);
or U17303 (N_17303,N_14550,N_14933);
nand U17304 (N_17304,N_15953,N_14827);
and U17305 (N_17305,N_14059,N_14001);
nor U17306 (N_17306,N_15659,N_14336);
nor U17307 (N_17307,N_14803,N_15617);
xnor U17308 (N_17308,N_15201,N_15697);
nand U17309 (N_17309,N_15076,N_14657);
nor U17310 (N_17310,N_14815,N_15880);
nand U17311 (N_17311,N_15199,N_14131);
or U17312 (N_17312,N_14363,N_15015);
and U17313 (N_17313,N_14947,N_14344);
or U17314 (N_17314,N_14404,N_14028);
nor U17315 (N_17315,N_14841,N_15669);
xor U17316 (N_17316,N_15026,N_15958);
nand U17317 (N_17317,N_15962,N_15379);
nor U17318 (N_17318,N_15379,N_14362);
nor U17319 (N_17319,N_15153,N_15120);
nand U17320 (N_17320,N_15677,N_15112);
and U17321 (N_17321,N_14330,N_14594);
and U17322 (N_17322,N_15586,N_15492);
and U17323 (N_17323,N_14464,N_15843);
or U17324 (N_17324,N_15368,N_14410);
and U17325 (N_17325,N_15299,N_15176);
nor U17326 (N_17326,N_14135,N_15065);
or U17327 (N_17327,N_15594,N_14105);
nand U17328 (N_17328,N_14843,N_15858);
and U17329 (N_17329,N_15874,N_14784);
nand U17330 (N_17330,N_15184,N_14150);
and U17331 (N_17331,N_15331,N_14635);
or U17332 (N_17332,N_15600,N_14926);
nand U17333 (N_17333,N_14439,N_15684);
or U17334 (N_17334,N_15251,N_15389);
nor U17335 (N_17335,N_15755,N_15652);
or U17336 (N_17336,N_14099,N_14777);
and U17337 (N_17337,N_15525,N_14115);
nand U17338 (N_17338,N_15965,N_15826);
nand U17339 (N_17339,N_15689,N_14271);
nand U17340 (N_17340,N_14701,N_15548);
or U17341 (N_17341,N_15139,N_14263);
or U17342 (N_17342,N_14180,N_14924);
nor U17343 (N_17343,N_15925,N_14800);
nand U17344 (N_17344,N_15412,N_14532);
nand U17345 (N_17345,N_14942,N_14276);
and U17346 (N_17346,N_15536,N_14162);
and U17347 (N_17347,N_14558,N_14079);
nand U17348 (N_17348,N_15052,N_15747);
and U17349 (N_17349,N_15620,N_15677);
nor U17350 (N_17350,N_14567,N_14047);
nor U17351 (N_17351,N_14000,N_14874);
or U17352 (N_17352,N_14375,N_14307);
nor U17353 (N_17353,N_15801,N_15586);
nand U17354 (N_17354,N_14130,N_14352);
nor U17355 (N_17355,N_14538,N_15252);
nor U17356 (N_17356,N_15861,N_14673);
nor U17357 (N_17357,N_15690,N_15590);
and U17358 (N_17358,N_15324,N_14186);
xnor U17359 (N_17359,N_14954,N_14742);
and U17360 (N_17360,N_14268,N_14405);
or U17361 (N_17361,N_15189,N_15261);
nand U17362 (N_17362,N_15562,N_14894);
nand U17363 (N_17363,N_15497,N_14664);
nand U17364 (N_17364,N_14436,N_14403);
and U17365 (N_17365,N_14551,N_14623);
and U17366 (N_17366,N_14103,N_14656);
nor U17367 (N_17367,N_15828,N_15466);
nor U17368 (N_17368,N_15216,N_15300);
and U17369 (N_17369,N_14707,N_14606);
and U17370 (N_17370,N_14915,N_15005);
nand U17371 (N_17371,N_14388,N_14918);
and U17372 (N_17372,N_14966,N_14892);
xor U17373 (N_17373,N_14824,N_14294);
nor U17374 (N_17374,N_15977,N_14404);
nor U17375 (N_17375,N_14969,N_15731);
nor U17376 (N_17376,N_14119,N_15416);
and U17377 (N_17377,N_15677,N_15332);
nor U17378 (N_17378,N_15063,N_15347);
and U17379 (N_17379,N_14850,N_15717);
xnor U17380 (N_17380,N_15087,N_14281);
or U17381 (N_17381,N_15084,N_14435);
or U17382 (N_17382,N_15440,N_15506);
nand U17383 (N_17383,N_15269,N_15217);
or U17384 (N_17384,N_14885,N_15570);
and U17385 (N_17385,N_14204,N_14708);
nand U17386 (N_17386,N_15655,N_15456);
and U17387 (N_17387,N_14620,N_14112);
xnor U17388 (N_17388,N_14477,N_15272);
and U17389 (N_17389,N_15607,N_15905);
and U17390 (N_17390,N_14819,N_14128);
or U17391 (N_17391,N_15694,N_14874);
or U17392 (N_17392,N_15807,N_14061);
and U17393 (N_17393,N_15403,N_14567);
nor U17394 (N_17394,N_14318,N_15646);
or U17395 (N_17395,N_15664,N_15275);
nor U17396 (N_17396,N_15777,N_14675);
xnor U17397 (N_17397,N_15543,N_15725);
or U17398 (N_17398,N_15768,N_15474);
nor U17399 (N_17399,N_14935,N_15468);
nor U17400 (N_17400,N_14501,N_14168);
or U17401 (N_17401,N_14572,N_14357);
and U17402 (N_17402,N_15820,N_14786);
nor U17403 (N_17403,N_14992,N_15970);
nor U17404 (N_17404,N_14344,N_14041);
or U17405 (N_17405,N_15695,N_15974);
and U17406 (N_17406,N_14193,N_14060);
nor U17407 (N_17407,N_14237,N_15011);
xnor U17408 (N_17408,N_14565,N_15766);
nor U17409 (N_17409,N_15917,N_15719);
xnor U17410 (N_17410,N_15084,N_14812);
nor U17411 (N_17411,N_15485,N_15619);
and U17412 (N_17412,N_14911,N_15795);
nor U17413 (N_17413,N_15511,N_14194);
and U17414 (N_17414,N_15465,N_15218);
nand U17415 (N_17415,N_14865,N_15428);
nor U17416 (N_17416,N_15968,N_15631);
and U17417 (N_17417,N_14466,N_14150);
nor U17418 (N_17418,N_15453,N_14759);
nor U17419 (N_17419,N_14073,N_15573);
or U17420 (N_17420,N_15840,N_14464);
and U17421 (N_17421,N_14938,N_14726);
nor U17422 (N_17422,N_14529,N_15742);
nor U17423 (N_17423,N_15778,N_14178);
nor U17424 (N_17424,N_15705,N_15837);
nand U17425 (N_17425,N_14560,N_15965);
or U17426 (N_17426,N_15251,N_14519);
nand U17427 (N_17427,N_15418,N_14260);
nor U17428 (N_17428,N_14616,N_14380);
or U17429 (N_17429,N_15515,N_14315);
or U17430 (N_17430,N_15981,N_14761);
and U17431 (N_17431,N_15834,N_14685);
or U17432 (N_17432,N_14525,N_15317);
nor U17433 (N_17433,N_15570,N_14061);
xnor U17434 (N_17434,N_14908,N_15953);
or U17435 (N_17435,N_14261,N_14652);
nor U17436 (N_17436,N_15457,N_14840);
or U17437 (N_17437,N_14508,N_15467);
nand U17438 (N_17438,N_14876,N_14678);
and U17439 (N_17439,N_14907,N_14128);
xor U17440 (N_17440,N_15636,N_15312);
xor U17441 (N_17441,N_14209,N_14122);
nor U17442 (N_17442,N_15813,N_15700);
and U17443 (N_17443,N_14986,N_15297);
nor U17444 (N_17444,N_14885,N_14775);
xor U17445 (N_17445,N_15190,N_15313);
or U17446 (N_17446,N_15431,N_14252);
and U17447 (N_17447,N_15621,N_14947);
nor U17448 (N_17448,N_15207,N_15426);
xor U17449 (N_17449,N_14435,N_15958);
and U17450 (N_17450,N_14982,N_14812);
nor U17451 (N_17451,N_15551,N_14488);
nor U17452 (N_17452,N_14252,N_14047);
or U17453 (N_17453,N_14875,N_15596);
nor U17454 (N_17454,N_14624,N_14791);
nand U17455 (N_17455,N_15722,N_15480);
nand U17456 (N_17456,N_15278,N_14394);
nor U17457 (N_17457,N_15011,N_15695);
and U17458 (N_17458,N_14334,N_15154);
nand U17459 (N_17459,N_15489,N_15651);
and U17460 (N_17460,N_14073,N_14186);
or U17461 (N_17461,N_15393,N_15504);
or U17462 (N_17462,N_14157,N_15729);
xnor U17463 (N_17463,N_15483,N_14430);
nor U17464 (N_17464,N_15391,N_14934);
nor U17465 (N_17465,N_14809,N_15233);
and U17466 (N_17466,N_14527,N_15508);
or U17467 (N_17467,N_15369,N_14197);
and U17468 (N_17468,N_15266,N_14687);
nor U17469 (N_17469,N_15364,N_14229);
or U17470 (N_17470,N_14224,N_14024);
nor U17471 (N_17471,N_15304,N_15497);
nor U17472 (N_17472,N_14878,N_15488);
and U17473 (N_17473,N_15924,N_15691);
xor U17474 (N_17474,N_15051,N_14074);
xnor U17475 (N_17475,N_14141,N_15821);
nor U17476 (N_17476,N_14898,N_14761);
and U17477 (N_17477,N_15373,N_14301);
and U17478 (N_17478,N_15605,N_14537);
or U17479 (N_17479,N_15990,N_14992);
nand U17480 (N_17480,N_14617,N_15975);
or U17481 (N_17481,N_15830,N_15756);
nand U17482 (N_17482,N_14797,N_14381);
nor U17483 (N_17483,N_14074,N_15973);
xor U17484 (N_17484,N_14333,N_15924);
and U17485 (N_17485,N_15041,N_14981);
and U17486 (N_17486,N_14556,N_14171);
or U17487 (N_17487,N_15348,N_14686);
nand U17488 (N_17488,N_15899,N_15259);
or U17489 (N_17489,N_14942,N_15123);
nor U17490 (N_17490,N_14126,N_15700);
nor U17491 (N_17491,N_14611,N_14563);
or U17492 (N_17492,N_15238,N_14353);
and U17493 (N_17493,N_15520,N_15119);
and U17494 (N_17494,N_14416,N_15627);
nor U17495 (N_17495,N_15242,N_14914);
or U17496 (N_17496,N_15289,N_15901);
nand U17497 (N_17497,N_14760,N_14822);
xor U17498 (N_17498,N_14975,N_15599);
xnor U17499 (N_17499,N_14866,N_14646);
nor U17500 (N_17500,N_14037,N_14598);
or U17501 (N_17501,N_15935,N_15852);
or U17502 (N_17502,N_14133,N_15957);
nor U17503 (N_17503,N_15768,N_14961);
or U17504 (N_17504,N_15808,N_14398);
nand U17505 (N_17505,N_14145,N_15144);
or U17506 (N_17506,N_15233,N_15120);
nand U17507 (N_17507,N_14872,N_14568);
nand U17508 (N_17508,N_15351,N_15033);
or U17509 (N_17509,N_15761,N_14677);
xor U17510 (N_17510,N_14283,N_14606);
and U17511 (N_17511,N_15034,N_15025);
nor U17512 (N_17512,N_15390,N_15300);
nand U17513 (N_17513,N_14188,N_15126);
nand U17514 (N_17514,N_14052,N_15507);
nor U17515 (N_17515,N_15199,N_14052);
and U17516 (N_17516,N_15123,N_15605);
xnor U17517 (N_17517,N_14025,N_15148);
or U17518 (N_17518,N_14280,N_14298);
nand U17519 (N_17519,N_14141,N_14261);
or U17520 (N_17520,N_15191,N_15766);
nor U17521 (N_17521,N_15943,N_14120);
and U17522 (N_17522,N_15901,N_15619);
nand U17523 (N_17523,N_15086,N_15267);
nand U17524 (N_17524,N_15223,N_15430);
or U17525 (N_17525,N_14702,N_15199);
nand U17526 (N_17526,N_15505,N_14896);
xnor U17527 (N_17527,N_14976,N_14133);
or U17528 (N_17528,N_14983,N_15942);
nand U17529 (N_17529,N_15484,N_14624);
or U17530 (N_17530,N_14437,N_14176);
or U17531 (N_17531,N_15465,N_14889);
and U17532 (N_17532,N_15770,N_14370);
and U17533 (N_17533,N_14442,N_15372);
or U17534 (N_17534,N_15090,N_15478);
and U17535 (N_17535,N_15043,N_14966);
xnor U17536 (N_17536,N_15466,N_14129);
xor U17537 (N_17537,N_15346,N_15294);
xor U17538 (N_17538,N_15629,N_15073);
nor U17539 (N_17539,N_14599,N_15273);
nand U17540 (N_17540,N_15968,N_14951);
xnor U17541 (N_17541,N_14056,N_15028);
and U17542 (N_17542,N_15919,N_14229);
or U17543 (N_17543,N_15918,N_14222);
nor U17544 (N_17544,N_14447,N_15463);
and U17545 (N_17545,N_15185,N_14722);
nand U17546 (N_17546,N_14623,N_14112);
or U17547 (N_17547,N_14184,N_15419);
or U17548 (N_17548,N_15221,N_15629);
and U17549 (N_17549,N_14723,N_15095);
xnor U17550 (N_17550,N_14925,N_15221);
nand U17551 (N_17551,N_14052,N_14452);
xnor U17552 (N_17552,N_15911,N_14992);
and U17553 (N_17553,N_14322,N_14000);
nor U17554 (N_17554,N_14624,N_15791);
or U17555 (N_17555,N_15266,N_14990);
nor U17556 (N_17556,N_15271,N_14403);
nor U17557 (N_17557,N_14622,N_15511);
or U17558 (N_17558,N_15399,N_14172);
or U17559 (N_17559,N_14483,N_15304);
or U17560 (N_17560,N_14629,N_14689);
nor U17561 (N_17561,N_14174,N_14440);
or U17562 (N_17562,N_14543,N_15859);
or U17563 (N_17563,N_14669,N_15767);
nor U17564 (N_17564,N_14904,N_14370);
or U17565 (N_17565,N_15677,N_15401);
nand U17566 (N_17566,N_14518,N_14907);
and U17567 (N_17567,N_15167,N_15392);
or U17568 (N_17568,N_14102,N_14674);
nor U17569 (N_17569,N_15163,N_14843);
nor U17570 (N_17570,N_14694,N_15287);
nand U17571 (N_17571,N_14387,N_15000);
nand U17572 (N_17572,N_15546,N_15358);
xor U17573 (N_17573,N_15494,N_15239);
nand U17574 (N_17574,N_15307,N_15490);
or U17575 (N_17575,N_15793,N_14225);
nor U17576 (N_17576,N_14096,N_14851);
nand U17577 (N_17577,N_15523,N_14252);
and U17578 (N_17578,N_14616,N_14697);
xor U17579 (N_17579,N_14680,N_15959);
xor U17580 (N_17580,N_15091,N_14650);
or U17581 (N_17581,N_14517,N_14143);
or U17582 (N_17582,N_14872,N_14537);
nor U17583 (N_17583,N_15452,N_15713);
and U17584 (N_17584,N_15040,N_14985);
or U17585 (N_17585,N_14372,N_14747);
and U17586 (N_17586,N_15474,N_14837);
nor U17587 (N_17587,N_14321,N_15373);
nand U17588 (N_17588,N_15130,N_14372);
or U17589 (N_17589,N_14207,N_14188);
nor U17590 (N_17590,N_15584,N_14985);
and U17591 (N_17591,N_15019,N_15713);
xor U17592 (N_17592,N_15788,N_14731);
or U17593 (N_17593,N_15026,N_14400);
nand U17594 (N_17594,N_15290,N_14536);
nor U17595 (N_17595,N_15246,N_15082);
xor U17596 (N_17596,N_15313,N_14735);
or U17597 (N_17597,N_15847,N_15967);
or U17598 (N_17598,N_14907,N_15716);
or U17599 (N_17599,N_14457,N_15916);
xor U17600 (N_17600,N_14310,N_15656);
nor U17601 (N_17601,N_15532,N_15681);
nand U17602 (N_17602,N_14848,N_15500);
and U17603 (N_17603,N_14887,N_15475);
nand U17604 (N_17604,N_15615,N_15718);
nand U17605 (N_17605,N_15597,N_15706);
or U17606 (N_17606,N_14838,N_14717);
nand U17607 (N_17607,N_14398,N_15591);
and U17608 (N_17608,N_15009,N_15040);
or U17609 (N_17609,N_14213,N_15577);
nand U17610 (N_17610,N_15173,N_15238);
and U17611 (N_17611,N_14550,N_14596);
or U17612 (N_17612,N_15805,N_15799);
nor U17613 (N_17613,N_15433,N_15664);
nor U17614 (N_17614,N_14002,N_14007);
and U17615 (N_17615,N_15773,N_15498);
nand U17616 (N_17616,N_15873,N_14533);
nand U17617 (N_17617,N_15742,N_14251);
xor U17618 (N_17618,N_15496,N_14401);
nor U17619 (N_17619,N_14538,N_15304);
nor U17620 (N_17620,N_15226,N_14374);
and U17621 (N_17621,N_15166,N_15396);
xor U17622 (N_17622,N_14759,N_14727);
or U17623 (N_17623,N_15712,N_14659);
and U17624 (N_17624,N_14324,N_14996);
and U17625 (N_17625,N_15854,N_15943);
nand U17626 (N_17626,N_15960,N_15783);
nand U17627 (N_17627,N_14910,N_14001);
nand U17628 (N_17628,N_14213,N_14097);
nor U17629 (N_17629,N_14275,N_15546);
or U17630 (N_17630,N_14922,N_15278);
nand U17631 (N_17631,N_14350,N_15611);
nor U17632 (N_17632,N_14231,N_15662);
and U17633 (N_17633,N_15022,N_15820);
nor U17634 (N_17634,N_14360,N_14789);
xnor U17635 (N_17635,N_14643,N_15313);
nor U17636 (N_17636,N_15928,N_15887);
nand U17637 (N_17637,N_15526,N_14742);
nor U17638 (N_17638,N_14681,N_14562);
nor U17639 (N_17639,N_15983,N_15021);
xnor U17640 (N_17640,N_15392,N_15477);
or U17641 (N_17641,N_14915,N_15679);
and U17642 (N_17642,N_14604,N_14458);
nand U17643 (N_17643,N_14078,N_15799);
nor U17644 (N_17644,N_15841,N_15395);
nand U17645 (N_17645,N_14069,N_14700);
nor U17646 (N_17646,N_14374,N_15917);
and U17647 (N_17647,N_15047,N_14476);
nor U17648 (N_17648,N_15726,N_14010);
nor U17649 (N_17649,N_15578,N_15902);
nand U17650 (N_17650,N_15496,N_14664);
nand U17651 (N_17651,N_15754,N_15006);
xnor U17652 (N_17652,N_15322,N_15159);
and U17653 (N_17653,N_15408,N_15048);
nor U17654 (N_17654,N_14373,N_15717);
and U17655 (N_17655,N_15159,N_14422);
nor U17656 (N_17656,N_14124,N_15559);
or U17657 (N_17657,N_14992,N_15396);
nand U17658 (N_17658,N_15810,N_15120);
or U17659 (N_17659,N_14631,N_14090);
or U17660 (N_17660,N_15758,N_15316);
and U17661 (N_17661,N_15505,N_14697);
and U17662 (N_17662,N_15949,N_15550);
nor U17663 (N_17663,N_14842,N_14197);
nor U17664 (N_17664,N_14160,N_14486);
or U17665 (N_17665,N_15762,N_14506);
or U17666 (N_17666,N_14362,N_15080);
or U17667 (N_17667,N_15129,N_14277);
xor U17668 (N_17668,N_15888,N_14707);
nor U17669 (N_17669,N_14298,N_15851);
and U17670 (N_17670,N_15145,N_15462);
and U17671 (N_17671,N_15137,N_14649);
or U17672 (N_17672,N_15967,N_15506);
nand U17673 (N_17673,N_15002,N_15487);
xnor U17674 (N_17674,N_14707,N_15975);
or U17675 (N_17675,N_14914,N_14687);
nor U17676 (N_17676,N_15189,N_14650);
nand U17677 (N_17677,N_14515,N_15254);
and U17678 (N_17678,N_14223,N_14493);
nor U17679 (N_17679,N_14761,N_14217);
and U17680 (N_17680,N_15070,N_15388);
nand U17681 (N_17681,N_14347,N_15408);
nand U17682 (N_17682,N_14181,N_14906);
nor U17683 (N_17683,N_14851,N_15963);
nor U17684 (N_17684,N_15886,N_15543);
nor U17685 (N_17685,N_15147,N_14213);
or U17686 (N_17686,N_15159,N_14078);
nand U17687 (N_17687,N_14541,N_15031);
nand U17688 (N_17688,N_15315,N_15019);
or U17689 (N_17689,N_15263,N_14266);
nor U17690 (N_17690,N_15568,N_14398);
and U17691 (N_17691,N_15559,N_15080);
and U17692 (N_17692,N_14780,N_14331);
or U17693 (N_17693,N_14732,N_14969);
nand U17694 (N_17694,N_14125,N_14433);
nand U17695 (N_17695,N_15909,N_15901);
or U17696 (N_17696,N_14809,N_14079);
nor U17697 (N_17697,N_14949,N_15018);
and U17698 (N_17698,N_15064,N_15939);
or U17699 (N_17699,N_15348,N_15090);
nand U17700 (N_17700,N_15005,N_15913);
nor U17701 (N_17701,N_14162,N_14083);
nand U17702 (N_17702,N_15200,N_15418);
nand U17703 (N_17703,N_14820,N_15626);
and U17704 (N_17704,N_15413,N_14704);
nand U17705 (N_17705,N_15714,N_14146);
nor U17706 (N_17706,N_14426,N_15224);
xnor U17707 (N_17707,N_14537,N_14470);
nor U17708 (N_17708,N_14051,N_14383);
or U17709 (N_17709,N_14970,N_14386);
nor U17710 (N_17710,N_15668,N_15275);
nand U17711 (N_17711,N_15346,N_14293);
or U17712 (N_17712,N_15760,N_15683);
nand U17713 (N_17713,N_15255,N_14349);
xnor U17714 (N_17714,N_14536,N_14045);
or U17715 (N_17715,N_14144,N_15705);
nor U17716 (N_17716,N_15034,N_15559);
nand U17717 (N_17717,N_15324,N_15406);
nand U17718 (N_17718,N_14102,N_14291);
and U17719 (N_17719,N_14763,N_15987);
nor U17720 (N_17720,N_14028,N_15220);
xnor U17721 (N_17721,N_15549,N_14219);
nand U17722 (N_17722,N_14548,N_15865);
xnor U17723 (N_17723,N_15294,N_14590);
nor U17724 (N_17724,N_14875,N_14883);
nand U17725 (N_17725,N_15640,N_14410);
nand U17726 (N_17726,N_15373,N_14514);
or U17727 (N_17727,N_14938,N_14936);
nor U17728 (N_17728,N_14460,N_14328);
nor U17729 (N_17729,N_14476,N_14620);
nand U17730 (N_17730,N_14490,N_14377);
and U17731 (N_17731,N_15610,N_15500);
and U17732 (N_17732,N_15604,N_15121);
nor U17733 (N_17733,N_14641,N_15984);
or U17734 (N_17734,N_14426,N_14088);
and U17735 (N_17735,N_14532,N_14703);
nor U17736 (N_17736,N_15311,N_15081);
and U17737 (N_17737,N_14004,N_14704);
and U17738 (N_17738,N_14089,N_14752);
and U17739 (N_17739,N_14941,N_15432);
and U17740 (N_17740,N_14059,N_15949);
nor U17741 (N_17741,N_15813,N_15625);
and U17742 (N_17742,N_15866,N_14774);
nand U17743 (N_17743,N_14481,N_15357);
and U17744 (N_17744,N_14551,N_15384);
nand U17745 (N_17745,N_14570,N_15697);
nor U17746 (N_17746,N_14373,N_15788);
nand U17747 (N_17747,N_15961,N_14790);
xor U17748 (N_17748,N_14004,N_15240);
and U17749 (N_17749,N_15575,N_14886);
or U17750 (N_17750,N_14723,N_14317);
or U17751 (N_17751,N_14698,N_14967);
or U17752 (N_17752,N_15228,N_14760);
nor U17753 (N_17753,N_15822,N_14292);
nand U17754 (N_17754,N_15282,N_15259);
nand U17755 (N_17755,N_15417,N_15915);
nand U17756 (N_17756,N_15265,N_14660);
nor U17757 (N_17757,N_14859,N_15003);
and U17758 (N_17758,N_15733,N_14234);
or U17759 (N_17759,N_14814,N_15437);
nand U17760 (N_17760,N_15842,N_15525);
xor U17761 (N_17761,N_14175,N_15019);
or U17762 (N_17762,N_15398,N_14654);
and U17763 (N_17763,N_15463,N_14160);
nand U17764 (N_17764,N_15807,N_15987);
nand U17765 (N_17765,N_15627,N_15510);
nor U17766 (N_17766,N_14187,N_14391);
nor U17767 (N_17767,N_15046,N_14654);
nor U17768 (N_17768,N_14559,N_15910);
or U17769 (N_17769,N_14769,N_15389);
and U17770 (N_17770,N_14989,N_15897);
or U17771 (N_17771,N_14843,N_14443);
or U17772 (N_17772,N_15748,N_15408);
and U17773 (N_17773,N_14361,N_14235);
or U17774 (N_17774,N_15651,N_14286);
nand U17775 (N_17775,N_14088,N_15103);
and U17776 (N_17776,N_14330,N_15963);
or U17777 (N_17777,N_15748,N_15826);
nor U17778 (N_17778,N_14300,N_15130);
and U17779 (N_17779,N_15131,N_15111);
and U17780 (N_17780,N_15050,N_14085);
xnor U17781 (N_17781,N_15674,N_14526);
or U17782 (N_17782,N_14682,N_14173);
nor U17783 (N_17783,N_15130,N_15488);
and U17784 (N_17784,N_15126,N_14204);
nor U17785 (N_17785,N_14415,N_14257);
xnor U17786 (N_17786,N_15344,N_14321);
nand U17787 (N_17787,N_14006,N_14144);
xor U17788 (N_17788,N_14706,N_14723);
nor U17789 (N_17789,N_15854,N_14424);
nand U17790 (N_17790,N_15304,N_15976);
xnor U17791 (N_17791,N_15325,N_15322);
or U17792 (N_17792,N_15148,N_14977);
nand U17793 (N_17793,N_15075,N_15054);
nor U17794 (N_17794,N_14675,N_15905);
nand U17795 (N_17795,N_15360,N_14986);
xor U17796 (N_17796,N_15105,N_15352);
nor U17797 (N_17797,N_14158,N_15437);
or U17798 (N_17798,N_15475,N_14051);
and U17799 (N_17799,N_15222,N_15011);
nand U17800 (N_17800,N_15801,N_14531);
nor U17801 (N_17801,N_15005,N_14429);
and U17802 (N_17802,N_14070,N_14491);
nand U17803 (N_17803,N_14158,N_14337);
nor U17804 (N_17804,N_15249,N_14671);
nor U17805 (N_17805,N_14008,N_15266);
and U17806 (N_17806,N_14066,N_15822);
nor U17807 (N_17807,N_15451,N_14834);
xnor U17808 (N_17808,N_15218,N_14751);
and U17809 (N_17809,N_14483,N_15441);
xnor U17810 (N_17810,N_15360,N_14300);
or U17811 (N_17811,N_14213,N_15319);
nand U17812 (N_17812,N_15638,N_15845);
nor U17813 (N_17813,N_15212,N_15898);
or U17814 (N_17814,N_15947,N_15951);
nand U17815 (N_17815,N_14933,N_15702);
and U17816 (N_17816,N_14673,N_15894);
or U17817 (N_17817,N_14139,N_15196);
xnor U17818 (N_17818,N_15896,N_15999);
nor U17819 (N_17819,N_15231,N_14606);
and U17820 (N_17820,N_14424,N_15159);
xnor U17821 (N_17821,N_15781,N_14722);
and U17822 (N_17822,N_14397,N_14706);
or U17823 (N_17823,N_14018,N_14367);
nand U17824 (N_17824,N_14824,N_14871);
and U17825 (N_17825,N_14366,N_15851);
and U17826 (N_17826,N_15707,N_15005);
or U17827 (N_17827,N_14027,N_15861);
or U17828 (N_17828,N_15101,N_15921);
and U17829 (N_17829,N_14945,N_15038);
nand U17830 (N_17830,N_15619,N_14826);
nor U17831 (N_17831,N_15082,N_15572);
or U17832 (N_17832,N_14414,N_15644);
nor U17833 (N_17833,N_14583,N_14142);
nand U17834 (N_17834,N_14905,N_15808);
and U17835 (N_17835,N_15981,N_14732);
and U17836 (N_17836,N_15401,N_15047);
xor U17837 (N_17837,N_14772,N_15033);
or U17838 (N_17838,N_15283,N_14428);
xor U17839 (N_17839,N_14737,N_15973);
nand U17840 (N_17840,N_15327,N_14002);
nand U17841 (N_17841,N_15284,N_14863);
and U17842 (N_17842,N_14272,N_15845);
or U17843 (N_17843,N_14903,N_15871);
nor U17844 (N_17844,N_15667,N_14740);
nand U17845 (N_17845,N_15191,N_15913);
nand U17846 (N_17846,N_15623,N_15725);
nand U17847 (N_17847,N_15622,N_15864);
nor U17848 (N_17848,N_15027,N_14733);
or U17849 (N_17849,N_14709,N_14918);
and U17850 (N_17850,N_15114,N_14846);
nand U17851 (N_17851,N_14817,N_15869);
nor U17852 (N_17852,N_14693,N_15288);
nor U17853 (N_17853,N_14718,N_15884);
nor U17854 (N_17854,N_14508,N_14321);
xnor U17855 (N_17855,N_15202,N_14158);
and U17856 (N_17856,N_15404,N_15446);
xnor U17857 (N_17857,N_14884,N_15726);
nand U17858 (N_17858,N_14677,N_14269);
nand U17859 (N_17859,N_14591,N_14863);
nor U17860 (N_17860,N_14880,N_15239);
nor U17861 (N_17861,N_14029,N_14494);
nand U17862 (N_17862,N_15218,N_15109);
or U17863 (N_17863,N_14239,N_15463);
and U17864 (N_17864,N_15690,N_14214);
nand U17865 (N_17865,N_14859,N_15652);
or U17866 (N_17866,N_14398,N_14354);
xnor U17867 (N_17867,N_14722,N_15255);
nand U17868 (N_17868,N_14260,N_14183);
nor U17869 (N_17869,N_14328,N_14620);
or U17870 (N_17870,N_14587,N_15984);
xnor U17871 (N_17871,N_14353,N_15625);
nand U17872 (N_17872,N_14431,N_15002);
or U17873 (N_17873,N_14166,N_15659);
and U17874 (N_17874,N_15974,N_14909);
or U17875 (N_17875,N_15148,N_15625);
nand U17876 (N_17876,N_14298,N_15552);
xor U17877 (N_17877,N_14254,N_14835);
and U17878 (N_17878,N_14848,N_14143);
and U17879 (N_17879,N_14625,N_15577);
nand U17880 (N_17880,N_14746,N_15606);
nor U17881 (N_17881,N_15255,N_15774);
and U17882 (N_17882,N_15218,N_15604);
nor U17883 (N_17883,N_15528,N_15916);
xnor U17884 (N_17884,N_15091,N_15237);
nor U17885 (N_17885,N_14774,N_14290);
xnor U17886 (N_17886,N_14700,N_15283);
nand U17887 (N_17887,N_15665,N_14471);
xor U17888 (N_17888,N_15427,N_15850);
and U17889 (N_17889,N_14074,N_14931);
nand U17890 (N_17890,N_14648,N_15577);
and U17891 (N_17891,N_15657,N_15425);
or U17892 (N_17892,N_15352,N_15171);
or U17893 (N_17893,N_15632,N_15309);
and U17894 (N_17894,N_15345,N_15674);
nor U17895 (N_17895,N_15502,N_14163);
or U17896 (N_17896,N_15814,N_15654);
or U17897 (N_17897,N_14041,N_15813);
or U17898 (N_17898,N_14199,N_15868);
nor U17899 (N_17899,N_15968,N_14992);
or U17900 (N_17900,N_15533,N_15311);
and U17901 (N_17901,N_15516,N_15428);
or U17902 (N_17902,N_14126,N_14692);
or U17903 (N_17903,N_14983,N_15212);
and U17904 (N_17904,N_14109,N_15220);
or U17905 (N_17905,N_15617,N_15370);
nor U17906 (N_17906,N_14468,N_14392);
nor U17907 (N_17907,N_14641,N_14644);
nand U17908 (N_17908,N_14271,N_15233);
and U17909 (N_17909,N_15631,N_15799);
or U17910 (N_17910,N_15863,N_15521);
nor U17911 (N_17911,N_15388,N_15252);
xor U17912 (N_17912,N_15003,N_15177);
and U17913 (N_17913,N_15856,N_14923);
nor U17914 (N_17914,N_15979,N_15377);
nor U17915 (N_17915,N_15816,N_15424);
nor U17916 (N_17916,N_15825,N_14830);
nor U17917 (N_17917,N_15048,N_14676);
and U17918 (N_17918,N_14553,N_14684);
and U17919 (N_17919,N_14469,N_15828);
or U17920 (N_17920,N_14689,N_14426);
xor U17921 (N_17921,N_15619,N_14223);
nand U17922 (N_17922,N_14461,N_14838);
and U17923 (N_17923,N_14149,N_15913);
nor U17924 (N_17924,N_14591,N_14097);
and U17925 (N_17925,N_15543,N_15813);
and U17926 (N_17926,N_14273,N_14629);
nor U17927 (N_17927,N_15064,N_15182);
nor U17928 (N_17928,N_14339,N_14491);
nand U17929 (N_17929,N_15096,N_15207);
and U17930 (N_17930,N_14341,N_15726);
nor U17931 (N_17931,N_15325,N_15471);
and U17932 (N_17932,N_14420,N_14511);
and U17933 (N_17933,N_15867,N_14201);
nor U17934 (N_17934,N_15719,N_15318);
and U17935 (N_17935,N_15433,N_15188);
and U17936 (N_17936,N_14405,N_14987);
and U17937 (N_17937,N_15447,N_15263);
nand U17938 (N_17938,N_15560,N_15461);
nand U17939 (N_17939,N_15991,N_14436);
or U17940 (N_17940,N_15179,N_14522);
or U17941 (N_17941,N_14728,N_15246);
and U17942 (N_17942,N_14470,N_14559);
and U17943 (N_17943,N_14547,N_14129);
nand U17944 (N_17944,N_15325,N_14822);
or U17945 (N_17945,N_15130,N_14738);
nand U17946 (N_17946,N_15919,N_15066);
nand U17947 (N_17947,N_15306,N_15597);
or U17948 (N_17948,N_14086,N_15079);
nor U17949 (N_17949,N_15587,N_14638);
nor U17950 (N_17950,N_14917,N_14473);
and U17951 (N_17951,N_14734,N_15330);
nand U17952 (N_17952,N_14563,N_15179);
nor U17953 (N_17953,N_15794,N_14491);
nor U17954 (N_17954,N_14886,N_15596);
or U17955 (N_17955,N_15807,N_14870);
and U17956 (N_17956,N_15739,N_14562);
or U17957 (N_17957,N_15447,N_15806);
and U17958 (N_17958,N_15897,N_15328);
nand U17959 (N_17959,N_14773,N_14685);
xnor U17960 (N_17960,N_14680,N_14996);
nor U17961 (N_17961,N_15199,N_14907);
xnor U17962 (N_17962,N_14750,N_14094);
and U17963 (N_17963,N_15640,N_15673);
and U17964 (N_17964,N_15266,N_15627);
or U17965 (N_17965,N_14088,N_15937);
nor U17966 (N_17966,N_15411,N_14043);
or U17967 (N_17967,N_14251,N_14719);
and U17968 (N_17968,N_14485,N_15534);
nor U17969 (N_17969,N_15008,N_15571);
or U17970 (N_17970,N_15044,N_15613);
xor U17971 (N_17971,N_14886,N_14019);
nand U17972 (N_17972,N_14912,N_15759);
and U17973 (N_17973,N_15956,N_14549);
nand U17974 (N_17974,N_14589,N_14975);
xnor U17975 (N_17975,N_15384,N_15302);
and U17976 (N_17976,N_14596,N_14502);
or U17977 (N_17977,N_14623,N_14659);
or U17978 (N_17978,N_14004,N_14950);
or U17979 (N_17979,N_14101,N_15484);
nand U17980 (N_17980,N_14069,N_14416);
or U17981 (N_17981,N_14174,N_14810);
or U17982 (N_17982,N_15712,N_15147);
and U17983 (N_17983,N_15159,N_15108);
nor U17984 (N_17984,N_15722,N_14704);
nand U17985 (N_17985,N_15557,N_15041);
and U17986 (N_17986,N_15442,N_14895);
and U17987 (N_17987,N_15115,N_14539);
or U17988 (N_17988,N_15161,N_15990);
nand U17989 (N_17989,N_14487,N_14546);
or U17990 (N_17990,N_15652,N_15482);
nand U17991 (N_17991,N_14618,N_14574);
nor U17992 (N_17992,N_15971,N_14747);
and U17993 (N_17993,N_14185,N_14553);
and U17994 (N_17994,N_14924,N_14232);
and U17995 (N_17995,N_14781,N_15987);
nor U17996 (N_17996,N_14495,N_14831);
or U17997 (N_17997,N_14400,N_14729);
nor U17998 (N_17998,N_15197,N_15680);
nand U17999 (N_17999,N_14813,N_14432);
and U18000 (N_18000,N_17807,N_16560);
nand U18001 (N_18001,N_17319,N_17800);
or U18002 (N_18002,N_16508,N_17304);
nand U18003 (N_18003,N_17863,N_17677);
nor U18004 (N_18004,N_17379,N_16610);
and U18005 (N_18005,N_16180,N_17516);
xor U18006 (N_18006,N_17995,N_16279);
and U18007 (N_18007,N_17078,N_16980);
and U18008 (N_18008,N_16233,N_16452);
nor U18009 (N_18009,N_16743,N_16339);
or U18010 (N_18010,N_16210,N_16244);
nor U18011 (N_18011,N_16993,N_17568);
nor U18012 (N_18012,N_16659,N_17281);
nand U18013 (N_18013,N_17954,N_16650);
xnor U18014 (N_18014,N_17385,N_16063);
and U18015 (N_18015,N_17802,N_17812);
or U18016 (N_18016,N_17463,N_17817);
nor U18017 (N_18017,N_16135,N_16264);
and U18018 (N_18018,N_16374,N_17896);
and U18019 (N_18019,N_16973,N_16534);
xnor U18020 (N_18020,N_17054,N_16300);
and U18021 (N_18021,N_17654,N_16075);
nor U18022 (N_18022,N_16608,N_16968);
or U18023 (N_18023,N_17309,N_17404);
nand U18024 (N_18024,N_17224,N_16584);
nand U18025 (N_18025,N_17183,N_16989);
nand U18026 (N_18026,N_17491,N_17259);
and U18027 (N_18027,N_17048,N_17950);
and U18028 (N_18028,N_16275,N_17306);
or U18029 (N_18029,N_17775,N_17887);
and U18030 (N_18030,N_16814,N_16910);
and U18031 (N_18031,N_16187,N_16904);
and U18032 (N_18032,N_16656,N_16462);
and U18033 (N_18033,N_17285,N_17408);
and U18034 (N_18034,N_16697,N_16791);
or U18035 (N_18035,N_17008,N_16850);
nor U18036 (N_18036,N_16157,N_17270);
and U18037 (N_18037,N_16047,N_16595);
xor U18038 (N_18038,N_17423,N_16485);
or U18039 (N_18039,N_17475,N_16478);
and U18040 (N_18040,N_16502,N_16683);
nand U18041 (N_18041,N_17032,N_16143);
nand U18042 (N_18042,N_17612,N_16809);
and U18043 (N_18043,N_17502,N_16556);
nor U18044 (N_18044,N_17198,N_17671);
nor U18045 (N_18045,N_16214,N_17001);
and U18046 (N_18046,N_17769,N_17640);
or U18047 (N_18047,N_17765,N_17993);
nand U18048 (N_18048,N_16375,N_16194);
nor U18049 (N_18049,N_16890,N_16321);
nor U18050 (N_18050,N_16440,N_16566);
nand U18051 (N_18051,N_16694,N_16444);
nor U18052 (N_18052,N_16184,N_17121);
or U18053 (N_18053,N_17715,N_16834);
nand U18054 (N_18054,N_16953,N_16223);
nor U18055 (N_18055,N_16874,N_16817);
xnor U18056 (N_18056,N_16905,N_16966);
and U18057 (N_18057,N_17342,N_16343);
and U18058 (N_18058,N_16597,N_16836);
nand U18059 (N_18059,N_16691,N_17790);
nand U18060 (N_18060,N_17696,N_16565);
nor U18061 (N_18061,N_17442,N_16951);
nor U18062 (N_18062,N_17543,N_16236);
or U18063 (N_18063,N_16745,N_16009);
nor U18064 (N_18064,N_17399,N_17865);
nor U18065 (N_18065,N_16921,N_16220);
nand U18066 (N_18066,N_16998,N_17165);
nand U18067 (N_18067,N_17426,N_16363);
or U18068 (N_18068,N_16093,N_17562);
nand U18069 (N_18069,N_17509,N_17301);
or U18070 (N_18070,N_16907,N_17551);
or U18071 (N_18071,N_17662,N_16901);
and U18072 (N_18072,N_17908,N_17197);
xnor U18073 (N_18073,N_17248,N_17360);
nor U18074 (N_18074,N_17272,N_17413);
and U18075 (N_18075,N_17446,N_17938);
nor U18076 (N_18076,N_16823,N_17965);
nand U18077 (N_18077,N_16253,N_16578);
and U18078 (N_18078,N_17033,N_17949);
or U18079 (N_18079,N_16420,N_17047);
and U18080 (N_18080,N_16765,N_16158);
nand U18081 (N_18081,N_16182,N_16119);
nor U18082 (N_18082,N_17981,N_17059);
nor U18083 (N_18083,N_16311,N_17030);
nor U18084 (N_18084,N_17407,N_17631);
xor U18085 (N_18085,N_17782,N_16794);
or U18086 (N_18086,N_16666,N_17526);
or U18087 (N_18087,N_17890,N_16131);
or U18088 (N_18088,N_17088,N_16642);
or U18089 (N_18089,N_17618,N_16107);
nand U18090 (N_18090,N_16759,N_16927);
nor U18091 (N_18091,N_17353,N_17928);
nor U18092 (N_18092,N_16407,N_17803);
nand U18093 (N_18093,N_16387,N_16755);
nor U18094 (N_18094,N_17756,N_16700);
nand U18095 (N_18095,N_17520,N_17736);
nand U18096 (N_18096,N_16050,N_16845);
nor U18097 (N_18097,N_17473,N_16055);
and U18098 (N_18098,N_16060,N_16322);
and U18099 (N_18099,N_17861,N_17398);
nand U18100 (N_18100,N_17395,N_17315);
xnor U18101 (N_18101,N_17713,N_16432);
or U18102 (N_18102,N_17739,N_17528);
or U18103 (N_18103,N_16630,N_16479);
or U18104 (N_18104,N_17341,N_17573);
or U18105 (N_18105,N_17441,N_16682);
nand U18106 (N_18106,N_16738,N_17916);
nor U18107 (N_18107,N_16766,N_17374);
and U18108 (N_18108,N_17042,N_16785);
and U18109 (N_18109,N_16494,N_17822);
or U18110 (N_18110,N_16764,N_17687);
and U18111 (N_18111,N_16709,N_17638);
and U18112 (N_18112,N_16971,N_17858);
or U18113 (N_18113,N_17091,N_17021);
and U18114 (N_18114,N_17286,N_16417);
or U18115 (N_18115,N_16978,N_16007);
nand U18116 (N_18116,N_16625,N_16357);
and U18117 (N_18117,N_17137,N_17770);
nor U18118 (N_18118,N_17621,N_16541);
and U18119 (N_18119,N_17280,N_17364);
and U18120 (N_18120,N_17912,N_16449);
or U18121 (N_18121,N_17962,N_17261);
or U18122 (N_18122,N_17120,N_17449);
xor U18123 (N_18123,N_17484,N_17829);
or U18124 (N_18124,N_16687,N_16672);
and U18125 (N_18125,N_16011,N_17875);
nor U18126 (N_18126,N_17716,N_16235);
and U18127 (N_18127,N_16928,N_17851);
or U18128 (N_18128,N_16170,N_17223);
nand U18129 (N_18129,N_17898,N_16199);
nor U18130 (N_18130,N_16392,N_17731);
xor U18131 (N_18131,N_17634,N_17682);
nor U18132 (N_18132,N_16990,N_16183);
nand U18133 (N_18133,N_16393,N_17106);
or U18134 (N_18134,N_17461,N_17658);
nand U18135 (N_18135,N_17542,N_16125);
xnor U18136 (N_18136,N_17324,N_16581);
nand U18137 (N_18137,N_17014,N_16090);
and U18138 (N_18138,N_17545,N_16287);
xor U18139 (N_18139,N_16999,N_17835);
and U18140 (N_18140,N_17531,N_16259);
nand U18141 (N_18141,N_17833,N_17102);
nand U18142 (N_18142,N_16269,N_17153);
xor U18143 (N_18143,N_16179,N_17480);
nor U18144 (N_18144,N_16692,N_16553);
nor U18145 (N_18145,N_16254,N_17348);
nor U18146 (N_18146,N_17410,N_17431);
nand U18147 (N_18147,N_17925,N_16832);
or U18148 (N_18148,N_17507,N_16081);
nand U18149 (N_18149,N_17086,N_17856);
or U18150 (N_18150,N_16028,N_16197);
or U18151 (N_18151,N_16885,N_16274);
nor U18152 (N_18152,N_17838,N_16395);
nor U18153 (N_18153,N_17874,N_17504);
nand U18154 (N_18154,N_16781,N_17171);
nor U18155 (N_18155,N_16493,N_17970);
or U18156 (N_18156,N_17750,N_17476);
nor U18157 (N_18157,N_17891,N_17845);
xor U18158 (N_18158,N_16883,N_17900);
nor U18159 (N_18159,N_17148,N_16870);
nand U18160 (N_18160,N_17037,N_17904);
nand U18161 (N_18161,N_17505,N_16974);
and U18162 (N_18162,N_17246,N_17295);
or U18163 (N_18163,N_16138,N_16078);
xnor U18164 (N_18164,N_16503,N_16835);
xor U18165 (N_18165,N_16021,N_16636);
nor U18166 (N_18166,N_17724,N_17237);
nor U18167 (N_18167,N_17494,N_16431);
xnor U18168 (N_18168,N_17847,N_17230);
nor U18169 (N_18169,N_16529,N_17038);
nand U18170 (N_18170,N_17514,N_17145);
and U18171 (N_18171,N_17337,N_17406);
or U18172 (N_18172,N_17955,N_17273);
or U18173 (N_18173,N_16278,N_16960);
nand U18174 (N_18174,N_17179,N_17496);
or U18175 (N_18175,N_17963,N_16389);
nor U18176 (N_18176,N_16411,N_17565);
nor U18177 (N_18177,N_17541,N_16286);
and U18178 (N_18178,N_16386,N_16139);
or U18179 (N_18179,N_17079,N_16470);
and U18180 (N_18180,N_16624,N_17396);
nand U18181 (N_18181,N_17058,N_17952);
nand U18182 (N_18182,N_16378,N_16342);
nand U18183 (N_18183,N_17241,N_17924);
nor U18184 (N_18184,N_17836,N_17308);
nor U18185 (N_18185,N_17255,N_17578);
xor U18186 (N_18186,N_17990,N_16576);
or U18187 (N_18187,N_16532,N_16903);
or U18188 (N_18188,N_16555,N_16171);
and U18189 (N_18189,N_17922,N_17068);
and U18190 (N_18190,N_17527,N_16314);
or U18191 (N_18191,N_16285,N_16002);
xor U18192 (N_18192,N_17331,N_16520);
nor U18193 (N_18193,N_17974,N_17643);
nor U18194 (N_18194,N_17109,N_17746);
nand U18195 (N_18195,N_17231,N_17683);
nand U18196 (N_18196,N_16875,N_16029);
nor U18197 (N_18197,N_17104,N_16318);
xnor U18198 (N_18198,N_17443,N_17848);
nor U18199 (N_18199,N_17667,N_17023);
nand U18200 (N_18200,N_16525,N_16705);
nand U18201 (N_18201,N_17244,N_17795);
or U18202 (N_18202,N_17436,N_16852);
and U18203 (N_18203,N_16162,N_17501);
nand U18204 (N_18204,N_17233,N_16773);
nor U18205 (N_18205,N_16716,N_17819);
nand U18206 (N_18206,N_16804,N_17809);
or U18207 (N_18207,N_16826,N_17783);
nor U18208 (N_18208,N_17370,N_17647);
nor U18209 (N_18209,N_17929,N_17992);
or U18210 (N_18210,N_17119,N_17701);
or U18211 (N_18211,N_17832,N_17036);
nand U18212 (N_18212,N_17753,N_16538);
and U18213 (N_18213,N_17823,N_17779);
or U18214 (N_18214,N_16023,N_16575);
or U18215 (N_18215,N_17227,N_16041);
nor U18216 (N_18216,N_17552,N_16327);
nor U18217 (N_18217,N_16186,N_17250);
nor U18218 (N_18218,N_17919,N_17905);
and U18219 (N_18219,N_16051,N_16326);
or U18220 (N_18220,N_17691,N_16001);
nand U18221 (N_18221,N_16092,N_16902);
nor U18222 (N_18222,N_17016,N_17204);
xor U18223 (N_18223,N_17983,N_16872);
or U18224 (N_18224,N_16984,N_16977);
and U18225 (N_18225,N_17382,N_16037);
nand U18226 (N_18226,N_17056,N_17646);
nand U18227 (N_18227,N_17401,N_17616);
and U18228 (N_18228,N_17367,N_16442);
nor U18229 (N_18229,N_16490,N_17140);
and U18230 (N_18230,N_16946,N_16152);
nand U18231 (N_18231,N_17866,N_16676);
xnor U18232 (N_18232,N_16718,N_17258);
xnor U18233 (N_18233,N_16748,N_17706);
nand U18234 (N_18234,N_17430,N_16406);
or U18235 (N_18235,N_16173,N_17697);
nor U18236 (N_18236,N_16784,N_17609);
nor U18237 (N_18237,N_16443,N_16871);
nand U18238 (N_18238,N_16886,N_16640);
or U18239 (N_18239,N_17810,N_17837);
nor U18240 (N_18240,N_17872,N_16600);
or U18241 (N_18241,N_16118,N_17125);
or U18242 (N_18242,N_17355,N_17296);
or U18243 (N_18243,N_16276,N_17266);
nor U18244 (N_18244,N_17584,N_17344);
xor U18245 (N_18245,N_16227,N_17070);
and U18246 (N_18246,N_16772,N_16088);
and U18247 (N_18247,N_17523,N_17346);
or U18248 (N_18248,N_17680,N_16097);
and U18249 (N_18249,N_16644,N_17740);
nor U18250 (N_18250,N_17567,N_17333);
nor U18251 (N_18251,N_16224,N_16238);
and U18252 (N_18252,N_16241,N_17641);
or U18253 (N_18253,N_16798,N_17672);
nand U18254 (N_18254,N_17347,N_16569);
nor U18255 (N_18255,N_16631,N_17143);
nand U18256 (N_18256,N_17967,N_16312);
nor U18257 (N_18257,N_17749,N_16113);
or U18258 (N_18258,N_17098,N_16937);
and U18259 (N_18259,N_17002,N_17608);
or U18260 (N_18260,N_16489,N_16195);
nand U18261 (N_18261,N_16364,N_16302);
nor U18262 (N_18262,N_17877,N_16100);
nor U18263 (N_18263,N_16935,N_16507);
xnor U18264 (N_18264,N_16572,N_16268);
or U18265 (N_18265,N_16251,N_17393);
or U18266 (N_18266,N_17936,N_16054);
or U18267 (N_18267,N_16258,N_17063);
and U18268 (N_18268,N_16371,N_16071);
nand U18269 (N_18269,N_17651,N_16667);
or U18270 (N_18270,N_16458,N_17524);
or U18271 (N_18271,N_17699,N_16067);
nor U18272 (N_18272,N_16196,N_17917);
nor U18273 (N_18273,N_17218,N_16942);
nor U18274 (N_18274,N_16154,N_16548);
nand U18275 (N_18275,N_16335,N_16669);
and U18276 (N_18276,N_16728,N_17852);
xnor U18277 (N_18277,N_17262,N_17359);
or U18278 (N_18278,N_17591,N_17689);
nor U18279 (N_18279,N_16609,N_16111);
nor U18280 (N_18280,N_17471,N_17320);
nand U18281 (N_18281,N_16463,N_16950);
or U18282 (N_18282,N_16505,N_17116);
nor U18283 (N_18283,N_17084,N_17458);
nor U18284 (N_18284,N_17225,N_17978);
xnor U18285 (N_18285,N_16737,N_16567);
xor U18286 (N_18286,N_16215,N_16715);
and U18287 (N_18287,N_16141,N_16559);
and U18288 (N_18288,N_17791,N_16109);
and U18289 (N_18289,N_16102,N_17416);
nand U18290 (N_18290,N_16517,N_16203);
or U18291 (N_18291,N_16844,N_17483);
and U18292 (N_18292,N_16104,N_17942);
and U18293 (N_18293,N_17208,N_17678);
nand U18294 (N_18294,N_16204,N_16024);
xnor U18295 (N_18295,N_17999,N_17422);
or U18296 (N_18296,N_16216,N_17944);
nand U18297 (N_18297,N_17610,N_16605);
and U18298 (N_18298,N_16592,N_17173);
and U18299 (N_18299,N_17708,N_17579);
nor U18300 (N_18300,N_17645,N_16218);
and U18301 (N_18301,N_16144,N_16382);
nor U18302 (N_18302,N_17652,N_16359);
nand U18303 (N_18303,N_16477,N_17433);
xnor U18304 (N_18304,N_16284,N_17044);
or U18305 (N_18305,N_17209,N_17011);
nand U18306 (N_18306,N_17323,N_16089);
or U18307 (N_18307,N_16723,N_16645);
xnor U18308 (N_18308,N_16762,N_16577);
xor U18309 (N_18309,N_16750,N_16132);
nand U18310 (N_18310,N_17558,N_17788);
xnor U18311 (N_18311,N_17139,N_16191);
or U18312 (N_18312,N_17655,N_17549);
nor U18313 (N_18313,N_16511,N_16263);
nor U18314 (N_18314,N_17611,N_16174);
or U18315 (N_18315,N_16026,N_16731);
xor U18316 (N_18316,N_16898,N_16945);
or U18317 (N_18317,N_16341,N_17768);
and U18318 (N_18318,N_17729,N_16776);
nand U18319 (N_18319,N_16954,N_17998);
or U18320 (N_18320,N_16615,N_17737);
or U18321 (N_18321,N_17217,N_17357);
or U18322 (N_18322,N_17006,N_17020);
xnor U18323 (N_18323,N_16512,N_17300);
nand U18324 (N_18324,N_16629,N_17214);
or U18325 (N_18325,N_16441,N_17221);
nor U18326 (N_18326,N_16424,N_16788);
nor U18327 (N_18327,N_17117,N_17155);
and U18328 (N_18328,N_16281,N_17821);
nor U18329 (N_18329,N_17450,N_17297);
nand U18330 (N_18330,N_17136,N_17580);
or U18331 (N_18331,N_17702,N_17299);
nand U18332 (N_18332,N_17384,N_16818);
and U18333 (N_18333,N_17964,N_17650);
nor U18334 (N_18334,N_17215,N_17329);
nand U18335 (N_18335,N_17151,N_16353);
and U18336 (N_18336,N_16879,N_16185);
nand U18337 (N_18337,N_17202,N_17097);
and U18338 (N_18338,N_16248,N_17168);
nand U18339 (N_18339,N_16652,N_17162);
and U18340 (N_18340,N_17681,N_17013);
nand U18341 (N_18341,N_17743,N_17878);
xnor U18342 (N_18342,N_17718,N_17825);
xor U18343 (N_18343,N_16077,N_16105);
nor U18344 (N_18344,N_16473,N_16841);
xor U18345 (N_18345,N_16775,N_17624);
nor U18346 (N_18346,N_16782,N_16146);
or U18347 (N_18347,N_16438,N_17532);
and U18348 (N_18348,N_17376,N_16367);
nand U18349 (N_18349,N_16733,N_16685);
xor U18350 (N_18350,N_17191,N_17553);
or U18351 (N_18351,N_17577,N_17445);
or U18352 (N_18352,N_16320,N_16213);
and U18353 (N_18353,N_16421,N_17727);
and U18354 (N_18354,N_16178,N_17670);
and U18355 (N_18355,N_17403,N_16291);
and U18356 (N_18356,N_16616,N_17115);
nor U18357 (N_18357,N_17004,N_16535);
nand U18358 (N_18358,N_17830,N_16803);
nand U18359 (N_18359,N_16433,N_17976);
and U18360 (N_18360,N_17247,N_16305);
nand U18361 (N_18361,N_17294,N_17675);
nor U18362 (N_18362,N_16134,N_16232);
nor U18363 (N_18363,N_16648,N_16668);
and U18364 (N_18364,N_17017,N_16448);
xnor U18365 (N_18365,N_16912,N_17457);
nand U18366 (N_18366,N_16777,N_16568);
xor U18367 (N_18367,N_16702,N_17419);
xor U18368 (N_18368,N_16713,N_16925);
xor U18369 (N_18369,N_16617,N_16126);
or U18370 (N_18370,N_17600,N_16040);
and U18371 (N_18371,N_17892,N_17585);
or U18372 (N_18372,N_16842,N_17535);
and U18373 (N_18373,N_16638,N_16074);
nand U18374 (N_18374,N_16365,N_17188);
or U18375 (N_18375,N_16727,N_17853);
nand U18376 (N_18376,N_16997,N_16416);
and U18377 (N_18377,N_16602,N_17635);
nand U18378 (N_18378,N_16524,N_17606);
and U18379 (N_18379,N_16779,N_16958);
and U18380 (N_18380,N_16317,N_17064);
and U18381 (N_18381,N_16770,N_16080);
or U18382 (N_18382,N_17291,N_16042);
nand U18383 (N_18383,N_17639,N_17172);
and U18384 (N_18384,N_16247,N_16255);
or U18385 (N_18385,N_17362,N_17328);
or U18386 (N_18386,N_17883,N_17050);
nand U18387 (N_18387,N_16988,N_17941);
or U18388 (N_18388,N_17862,N_17728);
nand U18389 (N_18389,N_17243,N_17688);
nor U18390 (N_18390,N_17096,N_16038);
and U18391 (N_18391,N_17642,N_16626);
nor U18392 (N_18392,N_16848,N_17538);
xnor U18393 (N_18393,N_16293,N_16588);
and U18394 (N_18394,N_17141,N_16720);
and U18395 (N_18395,N_16298,N_16456);
nor U18396 (N_18396,N_17519,N_16528);
nand U18397 (N_18397,N_16010,N_17622);
nor U18398 (N_18398,N_16551,N_17435);
nand U18399 (N_18399,N_17605,N_17045);
nand U18400 (N_18400,N_16379,N_17024);
nand U18401 (N_18401,N_17444,N_16159);
or U18402 (N_18402,N_16860,N_16108);
or U18403 (N_18403,N_16847,N_17991);
nor U18404 (N_18404,N_17888,N_16099);
nand U18405 (N_18405,N_16851,N_16915);
nor U18406 (N_18406,N_17763,N_16514);
and U18407 (N_18407,N_16543,N_16189);
nand U18408 (N_18408,N_16482,N_17659);
nand U18409 (N_18409,N_16033,N_17799);
nand U18410 (N_18410,N_16952,N_16854);
and U18411 (N_18411,N_16800,N_17040);
or U18412 (N_18412,N_16430,N_16604);
nor U18413 (N_18413,N_17870,N_16797);
or U18414 (N_18414,N_16563,N_16994);
nor U18415 (N_18415,N_16641,N_16896);
or U18416 (N_18416,N_17220,N_16061);
nand U18417 (N_18417,N_16603,N_16598);
xnor U18418 (N_18418,N_17897,N_16899);
xnor U18419 (N_18419,N_17871,N_16620);
or U18420 (N_18420,N_17352,N_16632);
nor U18421 (N_18421,N_16793,N_16426);
xnor U18422 (N_18422,N_16789,N_16969);
nor U18423 (N_18423,N_17010,N_17377);
or U18424 (N_18424,N_16714,N_17260);
and U18425 (N_18425,N_16995,N_17235);
xor U18426 (N_18426,N_16234,N_16192);
or U18427 (N_18427,N_17100,N_17118);
nand U18428 (N_18428,N_17705,N_17893);
xor U18429 (N_18429,N_17133,N_17177);
nand U18430 (N_18430,N_17147,N_16175);
or U18431 (N_18431,N_16283,N_16753);
nand U18432 (N_18432,N_17594,N_17182);
nor U18433 (N_18433,N_16758,N_17321);
nand U18434 (N_18434,N_16228,N_16405);
xnor U18435 (N_18435,N_17195,N_16265);
nand U18436 (N_18436,N_17498,N_17212);
and U18437 (N_18437,N_16140,N_17511);
or U18438 (N_18438,N_16701,N_17839);
and U18439 (N_18439,N_16231,N_17282);
or U18440 (N_18440,N_17387,N_17774);
and U18441 (N_18441,N_17012,N_17234);
nor U18442 (N_18442,N_17789,N_16892);
or U18443 (N_18443,N_17879,N_16025);
nand U18444 (N_18444,N_16926,N_16959);
or U18445 (N_18445,N_16309,N_16780);
nand U18446 (N_18446,N_17389,N_16006);
and U18447 (N_18447,N_17486,N_17583);
xnor U18448 (N_18448,N_16634,N_17603);
xor U18449 (N_18449,N_16976,N_17307);
xnor U18450 (N_18450,N_17864,N_16114);
and U18451 (N_18451,N_17161,N_16200);
and U18452 (N_18452,N_17284,N_17915);
nor U18453 (N_18453,N_17943,N_16744);
or U18454 (N_18454,N_16523,N_17424);
and U18455 (N_18455,N_16460,N_17095);
nor U18456 (N_18456,N_16461,N_17053);
and U18457 (N_18457,N_16334,N_16622);
nand U18458 (N_18458,N_16397,N_17434);
nor U18459 (N_18459,N_17757,N_17130);
nor U18460 (N_18460,N_16557,N_17249);
and U18461 (N_18461,N_17926,N_17719);
nor U18462 (N_18462,N_16437,N_17274);
nand U18463 (N_18463,N_16324,N_17025);
or U18464 (N_18464,N_16741,N_16229);
and U18465 (N_18465,N_17326,N_16065);
and U18466 (N_18466,N_16280,N_17813);
nor U18467 (N_18467,N_17717,N_17283);
nand U18468 (N_18468,N_17269,N_17150);
nor U18469 (N_18469,N_17894,N_16531);
xor U18470 (N_18470,N_16465,N_17834);
and U18471 (N_18471,N_16106,N_17418);
or U18472 (N_18472,N_17103,N_17420);
nand U18473 (N_18473,N_17889,N_17122);
and U18474 (N_18474,N_17907,N_16031);
nor U18475 (N_18475,N_16053,N_16661);
and U18476 (N_18476,N_17303,N_17164);
nor U18477 (N_18477,N_16816,N_17160);
nand U18478 (N_18478,N_16004,N_17707);
xnor U18479 (N_18479,N_16635,N_16708);
or U18480 (N_18480,N_16400,N_17167);
or U18481 (N_18481,N_16017,N_17134);
nand U18482 (N_18482,N_17128,N_17633);
xor U18483 (N_18483,N_16369,N_17325);
and U18484 (N_18484,N_16655,N_16085);
and U18485 (N_18485,N_16861,N_16344);
nor U18486 (N_18486,N_16756,N_17051);
nor U18487 (N_18487,N_17375,N_16190);
and U18488 (N_18488,N_17602,N_17007);
nor U18489 (N_18489,N_17415,N_16495);
and U18490 (N_18490,N_17203,N_17820);
xnor U18491 (N_18491,N_17158,N_16169);
nor U18492 (N_18492,N_17356,N_16066);
or U18493 (N_18493,N_17312,N_16121);
nor U18494 (N_18494,N_17236,N_16130);
xnor U18495 (N_18495,N_16868,N_17927);
and U18496 (N_18496,N_17945,N_17046);
or U18497 (N_18497,N_17674,N_17844);
or U18498 (N_18498,N_17588,N_16509);
nand U18499 (N_18499,N_16719,N_16880);
or U18500 (N_18500,N_16222,N_17625);
or U18501 (N_18501,N_17409,N_16404);
and U18502 (N_18502,N_17637,N_17777);
or U18503 (N_18503,N_16760,N_16574);
and U18504 (N_18504,N_16536,N_17684);
or U18505 (N_18505,N_16117,N_16355);
nor U18506 (N_18506,N_17206,N_17490);
nor U18507 (N_18507,N_17911,N_16689);
nor U18508 (N_18508,N_17318,N_16453);
or U18509 (N_18509,N_17525,N_16414);
nand U18510 (N_18510,N_16544,N_17190);
nand U18511 (N_18511,N_16752,N_17314);
nor U18512 (N_18512,N_16329,N_16252);
nor U18513 (N_18513,N_16332,N_17152);
nor U18514 (N_18514,N_16388,N_16153);
nor U18515 (N_18515,N_17482,N_17564);
and U18516 (N_18516,N_17730,N_16530);
nor U18517 (N_18517,N_16120,N_16558);
and U18518 (N_18518,N_16349,N_17453);
nand U18519 (N_18519,N_16472,N_16271);
and U18520 (N_18520,N_16221,N_17668);
nand U18521 (N_18521,N_17123,N_16142);
nand U18522 (N_18522,N_17003,N_17169);
and U18523 (N_18523,N_16331,N_17368);
nor U18524 (N_18524,N_17073,N_17163);
nand U18525 (N_18525,N_16891,N_16633);
nand U18526 (N_18526,N_16938,N_17953);
and U18527 (N_18527,N_16260,N_16706);
or U18528 (N_18528,N_17613,N_17439);
or U18529 (N_18529,N_17855,N_17586);
nand U18530 (N_18530,N_16916,N_16982);
nor U18531 (N_18531,N_16827,N_17752);
and U18532 (N_18532,N_17690,N_16579);
and U18533 (N_18533,N_17092,N_17636);
nor U18534 (N_18534,N_16427,N_16735);
and U18535 (N_18535,N_17210,N_16924);
and U18536 (N_18536,N_17029,N_17550);
or U18537 (N_18537,N_17723,N_16681);
and U18538 (N_18538,N_17714,N_16429);
and U18539 (N_18539,N_17288,N_16732);
and U18540 (N_18540,N_17869,N_17111);
and U18541 (N_18541,N_16979,N_17238);
xnor U18542 (N_18542,N_16129,N_16526);
nand U18543 (N_18543,N_16035,N_17110);
or U18544 (N_18544,N_16297,N_17448);
nor U18545 (N_18545,N_16445,N_16083);
and U18546 (N_18546,N_16864,N_16201);
or U18547 (N_18547,N_16815,N_17009);
and U18548 (N_18548,N_17517,N_17354);
or U18549 (N_18549,N_17087,N_16315);
xnor U18550 (N_18550,N_17910,N_16446);
nor U18551 (N_18551,N_17127,N_16580);
nand U18552 (N_18552,N_16292,N_16308);
and U18553 (N_18553,N_16778,N_17142);
nand U18554 (N_18554,N_17644,N_16516);
nand U18555 (N_18555,N_16267,N_16149);
and U18556 (N_18556,N_16671,N_16500);
and U18557 (N_18557,N_16394,N_16783);
nand U18558 (N_18558,N_16087,N_16436);
nor U18559 (N_18559,N_17090,N_17948);
xor U18560 (N_18560,N_16098,N_17544);
nand U18561 (N_18561,N_17057,N_17582);
xnor U18562 (N_18562,N_17432,N_17571);
nand U18563 (N_18563,N_16643,N_17868);
and U18564 (N_18564,N_17850,N_17921);
or U18565 (N_18565,N_17112,N_16361);
and U18566 (N_18566,N_17592,N_16821);
nor U18567 (N_18567,N_16045,N_16262);
and U18568 (N_18568,N_17530,N_17766);
nor U18569 (N_18569,N_16711,N_16920);
xor U18570 (N_18570,N_16722,N_17271);
and U18571 (N_18571,N_17597,N_16304);
nor U18572 (N_18572,N_16612,N_16887);
nand U18573 (N_18573,N_16351,N_17327);
or U18574 (N_18574,N_16936,N_16721);
or U18575 (N_18575,N_16628,N_17956);
and U18576 (N_18576,N_17598,N_16593);
nor U18577 (N_18577,N_17339,N_16552);
and U18578 (N_18578,N_16124,N_17960);
or U18579 (N_18579,N_16893,N_17539);
or U18580 (N_18580,N_17693,N_17885);
nand U18581 (N_18581,N_17289,N_16086);
nor U18582 (N_18582,N_16205,N_17559);
nand U18583 (N_18583,N_17028,N_17732);
nand U18584 (N_18584,N_17287,N_17604);
nor U18585 (N_18585,N_16545,N_16693);
or U18586 (N_18586,N_17762,N_16127);
nor U18587 (N_18587,N_17988,N_17614);
nor U18588 (N_18588,N_17465,N_17518);
or U18589 (N_18589,N_17977,N_17744);
nand U18590 (N_18590,N_16347,N_17797);
nand U18591 (N_18591,N_16751,N_17332);
or U18592 (N_18592,N_17213,N_17107);
and U18593 (N_18593,N_16813,N_17363);
nand U18594 (N_18594,N_17801,N_16792);
xnor U18595 (N_18595,N_16069,N_17947);
nand U18596 (N_18596,N_17411,N_16877);
nor U18597 (N_18597,N_16590,N_17184);
nand U18598 (N_18598,N_16742,N_16468);
nor U18599 (N_18599,N_17192,N_16328);
xor U18600 (N_18600,N_16016,N_16237);
and U18601 (N_18601,N_17089,N_17710);
xor U18602 (N_18602,N_16878,N_17229);
nor U18603 (N_18603,N_17378,N_17761);
and U18604 (N_18604,N_17648,N_16177);
and U18605 (N_18605,N_16145,N_16103);
and U18606 (N_18606,N_16282,N_16825);
or U18607 (N_18607,N_17781,N_17041);
and U18608 (N_18608,N_17468,N_17623);
nor U18609 (N_18609,N_16352,N_16418);
nor U18610 (N_18610,N_16164,N_16840);
nor U18611 (N_18611,N_16160,N_17176);
nand U18612 (N_18612,N_17469,N_16481);
nand U18613 (N_18613,N_16918,N_16601);
or U18614 (N_18614,N_17776,N_17239);
nor U18615 (N_18615,N_16225,N_16402);
or U18616 (N_18616,N_16934,N_17242);
and U18617 (N_18617,N_16261,N_16519);
or U18618 (N_18618,N_17540,N_17982);
or U18619 (N_18619,N_17316,N_17189);
nand U18620 (N_18620,N_16219,N_16325);
and U18621 (N_18621,N_16862,N_17913);
and U18622 (N_18622,N_16391,N_16790);
nand U18623 (N_18623,N_16450,N_16049);
nand U18624 (N_18624,N_16243,N_16385);
and U18625 (N_18625,N_17506,N_17267);
nor U18626 (N_18626,N_17589,N_17350);
nor U18627 (N_18627,N_17330,N_16521);
or U18628 (N_18628,N_16975,N_17816);
nand U18629 (N_18629,N_17735,N_17798);
or U18630 (N_18630,N_16455,N_16726);
and U18631 (N_18631,N_16469,N_16483);
and U18632 (N_18632,N_17201,N_17425);
nor U18633 (N_18633,N_17276,N_16467);
nor U18634 (N_18634,N_17254,N_16591);
nand U18635 (N_18635,N_17755,N_16699);
xnor U18636 (N_18636,N_17661,N_16039);
and U18637 (N_18637,N_17200,N_16206);
nor U18638 (N_18638,N_16340,N_16207);
and U18639 (N_18639,N_17778,N_16346);
and U18640 (N_18640,N_17811,N_17438);
and U18641 (N_18641,N_16857,N_16073);
or U18642 (N_18642,N_17388,N_16614);
or U18643 (N_18643,N_16774,N_16408);
nand U18644 (N_18644,N_16808,N_17828);
and U18645 (N_18645,N_16398,N_16176);
or U18646 (N_18646,N_16451,N_16005);
nor U18647 (N_18647,N_17488,N_17903);
xnor U18648 (N_18648,N_17909,N_16822);
or U18649 (N_18649,N_16647,N_17292);
and U18650 (N_18650,N_17178,N_17628);
or U18651 (N_18651,N_17806,N_16000);
and U18652 (N_18652,N_17669,N_17062);
xor U18653 (N_18653,N_17607,N_17031);
nor U18654 (N_18654,N_17181,N_16019);
nand U18655 (N_18655,N_17278,N_17521);
nand U18656 (N_18656,N_16704,N_17467);
nor U18657 (N_18657,N_16046,N_17961);
and U18658 (N_18658,N_16734,N_16381);
nor U18659 (N_18659,N_16044,N_16030);
nor U18660 (N_18660,N_17997,N_17000);
nor U18661 (N_18661,N_16707,N_16422);
xnor U18662 (N_18662,N_17773,N_17599);
and U18663 (N_18663,N_16674,N_16245);
nand U18664 (N_18664,N_16496,N_16337);
nor U18665 (N_18665,N_17489,N_17548);
and U18666 (N_18666,N_17593,N_16198);
xor U18667 (N_18667,N_16256,N_17219);
nor U18668 (N_18668,N_16048,N_16627);
nand U18669 (N_18669,N_16740,N_17940);
nand U18670 (N_18670,N_16819,N_17842);
xor U18671 (N_18671,N_17400,N_17815);
or U18672 (N_18672,N_16383,N_17787);
or U18673 (N_18673,N_16802,N_16853);
nand U18674 (N_18674,N_16837,N_17686);
nand U18675 (N_18675,N_16095,N_17066);
or U18676 (N_18676,N_17581,N_16831);
and U18677 (N_18677,N_16027,N_17345);
nand U18678 (N_18678,N_17185,N_16986);
and U18679 (N_18679,N_16486,N_16573);
and U18680 (N_18680,N_16812,N_16838);
xor U18681 (N_18681,N_16983,N_16717);
and U18682 (N_18682,N_17576,N_16323);
and U18683 (N_18683,N_17510,N_17015);
or U18684 (N_18684,N_16510,N_16101);
and U18685 (N_18685,N_17108,N_16466);
nor U18686 (N_18686,N_17786,N_17751);
nand U18687 (N_18687,N_16504,N_16410);
and U18688 (N_18688,N_17747,N_17764);
nand U18689 (N_18689,N_17754,N_17334);
nand U18690 (N_18690,N_17497,N_17222);
nor U18691 (N_18691,N_17487,N_17733);
and U18692 (N_18692,N_16447,N_16806);
xor U18693 (N_18693,N_16897,N_16922);
nand U18694 (N_18694,N_16646,N_16148);
nand U18695 (N_18695,N_16658,N_16582);
nor U18696 (N_18696,N_17698,N_16749);
nor U18697 (N_18697,N_17113,N_17666);
or U18698 (N_18698,N_16249,N_16739);
or U18699 (N_18699,N_16294,N_16796);
nor U18700 (N_18700,N_16246,N_16963);
xnor U18701 (N_18701,N_16833,N_16947);
nor U18702 (N_18702,N_16415,N_16606);
and U18703 (N_18703,N_17369,N_17481);
nand U18704 (N_18704,N_16677,N_16396);
nand U18705 (N_18705,N_16549,N_17338);
nand U18706 (N_18706,N_16497,N_16881);
nand U18707 (N_18707,N_17462,N_17402);
and U18708 (N_18708,N_17515,N_17043);
xor U18709 (N_18709,N_17060,N_16967);
nor U18710 (N_18710,N_17601,N_16539);
and U18711 (N_18711,N_17959,N_17027);
nand U18712 (N_18712,N_16226,N_17380);
xnor U18713 (N_18713,N_16824,N_17226);
or U18714 (N_18714,N_17796,N_17771);
nor U18715 (N_18715,N_17500,N_16068);
or U18716 (N_18716,N_17760,N_16079);
or U18717 (N_18717,N_17673,N_16457);
nor U18718 (N_18718,N_16515,N_17937);
or U18719 (N_18719,N_16895,N_16115);
nand U18720 (N_18720,N_17923,N_17154);
nand U18721 (N_18721,N_16356,N_17824);
and U18722 (N_18722,N_17554,N_16859);
nor U18723 (N_18723,N_16380,N_17094);
xnor U18724 (N_18724,N_17251,N_17493);
and U18725 (N_18725,N_17138,N_17302);
nor U18726 (N_18726,N_17022,N_16301);
nand U18727 (N_18727,N_17313,N_17067);
nor U18728 (N_18728,N_16761,N_16729);
or U18729 (N_18729,N_17159,N_16923);
xor U18730 (N_18730,N_16082,N_16242);
or U18731 (N_18731,N_16018,N_17703);
and U18732 (N_18732,N_16858,N_16763);
nor U18733 (N_18733,N_16172,N_17841);
nor U18734 (N_18734,N_17373,N_16319);
or U18735 (N_18735,N_17656,N_16948);
or U18736 (N_18736,N_16136,N_17694);
or U18737 (N_18737,N_17157,N_16801);
nor U18738 (N_18738,N_17649,N_16188);
or U18739 (N_18739,N_16116,N_16985);
or U18740 (N_18740,N_16849,N_16310);
and U18741 (N_18741,N_16811,N_16820);
or U18742 (N_18742,N_17186,N_16166);
nor U18743 (N_18743,N_16435,N_17005);
or U18744 (N_18744,N_17075,N_16856);
or U18745 (N_18745,N_16961,N_16059);
nand U18746 (N_18746,N_16202,N_16767);
or U18747 (N_18747,N_16649,N_16884);
and U18748 (N_18748,N_16955,N_16561);
nand U18749 (N_18749,N_17055,N_16064);
nor U18750 (N_18750,N_17322,N_16660);
nand U18751 (N_18751,N_17931,N_16015);
or U18752 (N_18752,N_16654,N_17720);
and U18753 (N_18753,N_17129,N_16939);
and U18754 (N_18754,N_17083,N_16621);
or U18755 (N_18755,N_17279,N_17405);
and U18756 (N_18756,N_16933,N_17767);
and U18757 (N_18757,N_16403,N_16688);
and U18758 (N_18758,N_17826,N_16419);
and U18759 (N_18759,N_16487,N_17629);
nor U18760 (N_18760,N_16680,N_17263);
and U18761 (N_18761,N_16499,N_17989);
xor U18762 (N_18762,N_16270,N_17149);
nand U18763 (N_18763,N_16014,N_17785);
nand U18764 (N_18764,N_17814,N_17440);
xor U18765 (N_18765,N_16795,N_17792);
xnor U18766 (N_18766,N_17725,N_17077);
and U18767 (N_18767,N_17704,N_17264);
xor U18768 (N_18768,N_17397,N_16637);
nand U18769 (N_18769,N_16163,N_16501);
nor U18770 (N_18770,N_17456,N_17293);
and U18771 (N_18771,N_16589,N_16554);
xnor U18772 (N_18772,N_17485,N_17882);
nand U18773 (N_18773,N_16583,N_16611);
or U18774 (N_18774,N_17709,N_16866);
nand U18775 (N_18775,N_16570,N_17726);
or U18776 (N_18776,N_17557,N_16888);
and U18777 (N_18777,N_17455,N_17886);
or U18778 (N_18778,N_17617,N_17076);
nand U18779 (N_18779,N_16345,N_16360);
nand U18780 (N_18780,N_17351,N_17657);
nand U18781 (N_18781,N_16736,N_17745);
nor U18782 (N_18782,N_16299,N_16156);
nor U18783 (N_18783,N_17340,N_16932);
nand U18784 (N_18784,N_17575,N_17758);
or U18785 (N_18785,N_17228,N_16412);
xnor U18786 (N_18786,N_16911,N_17881);
nand U18787 (N_18787,N_16863,N_16208);
nand U18788 (N_18788,N_16757,N_16333);
or U18789 (N_18789,N_16805,N_17187);
or U18790 (N_18790,N_17460,N_17536);
xor U18791 (N_18791,N_16972,N_17734);
or U18792 (N_18792,N_17563,N_16876);
nor U18793 (N_18793,N_17080,N_16846);
or U18794 (N_18794,N_17880,N_17857);
nand U18795 (N_18795,N_16913,N_17421);
and U18796 (N_18796,N_16623,N_16167);
and U18797 (N_18797,N_16390,N_16217);
nand U18798 (N_18798,N_16957,N_16571);
or U18799 (N_18799,N_17620,N_16919);
or U18800 (N_18800,N_16240,N_17166);
and U18801 (N_18801,N_17477,N_17619);
or U18802 (N_18802,N_16498,N_17759);
nand U18803 (N_18803,N_17459,N_16665);
xnor U18804 (N_18804,N_16348,N_16596);
or U18805 (N_18805,N_16072,N_16373);
and U18806 (N_18806,N_16193,N_16043);
nor U18807 (N_18807,N_17437,N_16786);
nand U18808 (N_18808,N_16506,N_17196);
and U18809 (N_18809,N_17700,N_17474);
nor U18810 (N_18810,N_16370,N_17211);
xnor U18811 (N_18811,N_17503,N_16056);
nand U18812 (N_18812,N_17906,N_16290);
nand U18813 (N_18813,N_16639,N_17537);
or U18814 (N_18814,N_17587,N_17335);
nand U18815 (N_18815,N_16076,N_16439);
or U18816 (N_18816,N_16869,N_16909);
or U18817 (N_18817,N_17843,N_16474);
or U18818 (N_18818,N_16613,N_16562);
nor U18819 (N_18819,N_16338,N_17895);
nand U18820 (N_18820,N_17804,N_17846);
or U18821 (N_18821,N_16965,N_17712);
and U18822 (N_18822,N_17365,N_16476);
and U18823 (N_18823,N_17546,N_17256);
nand U18824 (N_18824,N_16288,N_16542);
and U18825 (N_18825,N_17626,N_17918);
nor U18826 (N_18826,N_17170,N_16653);
nand U18827 (N_18827,N_17245,N_16155);
or U18828 (N_18828,N_16678,N_16316);
nor U18829 (N_18829,N_16358,N_16471);
and U18830 (N_18830,N_17268,N_17358);
or U18831 (N_18831,N_16585,N_17074);
and U18832 (N_18832,N_17772,N_16894);
or U18833 (N_18833,N_16366,N_17193);
and U18834 (N_18834,N_16829,N_16564);
nor U18835 (N_18835,N_16730,N_16272);
nand U18836 (N_18836,N_16949,N_16599);
or U18837 (N_18837,N_16303,N_16354);
nor U18838 (N_18838,N_16787,N_17513);
and U18839 (N_18839,N_17920,N_16799);
and U18840 (N_18840,N_17175,N_16810);
nor U18841 (N_18841,N_16434,N_16675);
nand U18842 (N_18842,N_17973,N_16698);
and U18843 (N_18843,N_16091,N_17180);
and U18844 (N_18844,N_17794,N_16929);
or U18845 (N_18845,N_17257,N_17232);
or U18846 (N_18846,N_16384,N_16133);
nand U18847 (N_18847,N_17381,N_16211);
nand U18848 (N_18848,N_16527,N_17464);
nand U18849 (N_18849,N_16996,N_16867);
nor U18850 (N_18850,N_16150,N_16768);
nand U18851 (N_18851,N_16096,N_16484);
or U18852 (N_18852,N_17572,N_17979);
nor U18853 (N_18853,N_17876,N_16032);
nor U18854 (N_18854,N_17305,N_16273);
nand U18855 (N_18855,N_17986,N_16034);
or U18856 (N_18856,N_17417,N_17093);
xnor U18857 (N_18857,N_17290,N_16754);
and U18858 (N_18858,N_16944,N_16664);
or U18859 (N_18859,N_17957,N_16662);
nor U18860 (N_18860,N_17566,N_17653);
and U18861 (N_18861,N_16917,N_17156);
xnor U18862 (N_18862,N_17065,N_17561);
nor U18863 (N_18863,N_17049,N_17722);
or U18864 (N_18864,N_16459,N_17996);
nor U18865 (N_18865,N_17026,N_16684);
or U18866 (N_18866,N_16425,N_16362);
nand U18867 (N_18867,N_17742,N_16058);
or U18868 (N_18868,N_16454,N_17522);
and U18869 (N_18869,N_17994,N_17311);
and U18870 (N_18870,N_17632,N_17854);
nor U18871 (N_18871,N_17132,N_16480);
nor U18872 (N_18872,N_16830,N_17529);
and U18873 (N_18873,N_16330,N_17741);
xnor U18874 (N_18874,N_17146,N_17061);
and U18875 (N_18875,N_16008,N_17034);
and U18876 (N_18876,N_16250,N_17664);
xor U18877 (N_18877,N_16930,N_17361);
and U18878 (N_18878,N_17867,N_16209);
nor U18879 (N_18879,N_16679,N_16546);
or U18880 (N_18880,N_17427,N_16873);
nand U18881 (N_18881,N_17277,N_16673);
nor U18882 (N_18882,N_16518,N_16307);
nand U18883 (N_18883,N_17679,N_16619);
nand U18884 (N_18884,N_16128,N_16540);
nor U18885 (N_18885,N_17534,N_16168);
and U18886 (N_18886,N_17721,N_17596);
nand U18887 (N_18887,N_17124,N_17072);
xor U18888 (N_18888,N_17972,N_16889);
or U18889 (N_18889,N_17207,N_16908);
and U18890 (N_18890,N_16306,N_16607);
nor U18891 (N_18891,N_16277,N_16401);
or U18892 (N_18892,N_17859,N_16257);
xnor U18893 (N_18893,N_17174,N_16491);
nor U18894 (N_18894,N_17884,N_17447);
or U18895 (N_18895,N_17738,N_17899);
nor U18896 (N_18896,N_17019,N_17429);
nor U18897 (N_18897,N_16052,N_17533);
and U18898 (N_18898,N_17383,N_17452);
nor U18899 (N_18899,N_16423,N_17349);
and U18900 (N_18900,N_17615,N_17939);
and U18901 (N_18901,N_17914,N_17071);
or U18902 (N_18902,N_17508,N_16239);
or U18903 (N_18903,N_16670,N_16724);
nand U18904 (N_18904,N_17194,N_17630);
nand U18905 (N_18905,N_16013,N_16062);
nor U18906 (N_18906,N_17574,N_16036);
nand U18907 (N_18907,N_17969,N_16533);
and U18908 (N_18908,N_16399,N_17479);
or U18909 (N_18909,N_16161,N_17695);
and U18910 (N_18910,N_17512,N_16022);
xnor U18911 (N_18911,N_17971,N_17470);
nand U18912 (N_18912,N_16376,N_16769);
nor U18913 (N_18913,N_17663,N_17499);
nor U18914 (N_18914,N_16212,N_17205);
nor U18915 (N_18915,N_17685,N_16122);
nand U18916 (N_18916,N_17343,N_16084);
nand U18917 (N_18917,N_16295,N_17391);
and U18918 (N_18918,N_17556,N_17873);
nand U18919 (N_18919,N_17085,N_17827);
and U18920 (N_18920,N_16943,N_16336);
nand U18921 (N_18921,N_16914,N_17114);
nor U18922 (N_18922,N_16587,N_17492);
nand U18923 (N_18923,N_16181,N_17126);
nor U18924 (N_18924,N_16981,N_17901);
nand U18925 (N_18925,N_17951,N_17252);
or U18926 (N_18926,N_16686,N_16475);
nor U18927 (N_18927,N_16464,N_16987);
xnor U18928 (N_18928,N_16537,N_17660);
or U18929 (N_18929,N_17560,N_16230);
nor U18930 (N_18930,N_17676,N_16725);
or U18931 (N_18931,N_16368,N_16651);
or U18932 (N_18932,N_16855,N_17860);
or U18933 (N_18933,N_16513,N_16941);
or U18934 (N_18934,N_17372,N_17987);
nor U18935 (N_18935,N_16618,N_17478);
nand U18936 (N_18936,N_16940,N_16070);
nand U18937 (N_18937,N_17933,N_17805);
nor U18938 (N_18938,N_17958,N_17935);
nand U18939 (N_18939,N_16828,N_17135);
or U18940 (N_18940,N_16428,N_16882);
nand U18941 (N_18941,N_16696,N_16488);
nor U18942 (N_18942,N_17985,N_16165);
nor U18943 (N_18943,N_17780,N_16992);
or U18944 (N_18944,N_17984,N_16313);
or U18945 (N_18945,N_17808,N_17265);
nor U18946 (N_18946,N_17966,N_16550);
nand U18947 (N_18947,N_16970,N_16094);
or U18948 (N_18948,N_17298,N_16900);
nor U18949 (N_18949,N_17932,N_16712);
and U18950 (N_18950,N_17082,N_17018);
nor U18951 (N_18951,N_17414,N_17495);
nor U18952 (N_18952,N_17101,N_17547);
or U18953 (N_18953,N_17472,N_16372);
or U18954 (N_18954,N_17692,N_17570);
nand U18955 (N_18955,N_17199,N_16151);
nand U18956 (N_18956,N_17081,N_16110);
xnor U18957 (N_18957,N_17934,N_16710);
nand U18958 (N_18958,N_17793,N_17390);
nand U18959 (N_18959,N_17451,N_16112);
and U18960 (N_18960,N_16522,N_16746);
or U18961 (N_18961,N_17216,N_17253);
xnor U18962 (N_18962,N_17946,N_17849);
nor U18963 (N_18963,N_16289,N_17555);
or U18964 (N_18964,N_17840,N_16843);
and U18965 (N_18965,N_16991,N_17569);
nand U18966 (N_18966,N_17454,N_16839);
and U18967 (N_18967,N_17310,N_16012);
nor U18968 (N_18968,N_16586,N_16147);
nor U18969 (N_18969,N_16865,N_17386);
or U18970 (N_18970,N_16690,N_16594);
or U18971 (N_18971,N_17930,N_16409);
and U18972 (N_18972,N_16807,N_17336);
nand U18973 (N_18973,N_17466,N_17590);
nand U18974 (N_18974,N_16695,N_17052);
or U18975 (N_18975,N_16350,N_17035);
and U18976 (N_18976,N_16747,N_17665);
nor U18977 (N_18977,N_16266,N_17627);
xor U18978 (N_18978,N_17131,N_16771);
nand U18979 (N_18979,N_16003,N_16296);
and U18980 (N_18980,N_17366,N_16547);
or U18981 (N_18981,N_16962,N_16964);
nor U18982 (N_18982,N_17240,N_17039);
or U18983 (N_18983,N_16413,N_17144);
and U18984 (N_18984,N_16492,N_17275);
nor U18985 (N_18985,N_17392,N_16931);
nand U18986 (N_18986,N_16020,N_16057);
and U18987 (N_18987,N_17394,N_17099);
and U18988 (N_18988,N_17428,N_17412);
nor U18989 (N_18989,N_16123,N_17784);
nor U18990 (N_18990,N_17748,N_17975);
nor U18991 (N_18991,N_17980,N_16703);
or U18992 (N_18992,N_17818,N_17371);
nor U18993 (N_18993,N_17069,N_17595);
and U18994 (N_18994,N_17831,N_17317);
nand U18995 (N_18995,N_17902,N_16377);
and U18996 (N_18996,N_16663,N_16956);
and U18997 (N_18997,N_16906,N_17968);
nor U18998 (N_18998,N_16137,N_17711);
nand U18999 (N_18999,N_16657,N_17105);
or U19000 (N_19000,N_17077,N_16536);
and U19001 (N_19001,N_17377,N_17292);
or U19002 (N_19002,N_17418,N_16473);
or U19003 (N_19003,N_17154,N_17149);
nand U19004 (N_19004,N_16616,N_16064);
nand U19005 (N_19005,N_16069,N_17760);
nand U19006 (N_19006,N_16956,N_17433);
and U19007 (N_19007,N_16870,N_17281);
and U19008 (N_19008,N_16091,N_17083);
or U19009 (N_19009,N_17236,N_16310);
xor U19010 (N_19010,N_16245,N_16668);
or U19011 (N_19011,N_16875,N_16765);
nand U19012 (N_19012,N_17525,N_17003);
and U19013 (N_19013,N_17440,N_17552);
nand U19014 (N_19014,N_16071,N_17533);
nor U19015 (N_19015,N_17500,N_17870);
nor U19016 (N_19016,N_17648,N_17966);
and U19017 (N_19017,N_16028,N_16524);
or U19018 (N_19018,N_17149,N_17636);
nor U19019 (N_19019,N_16460,N_17444);
or U19020 (N_19020,N_16097,N_17408);
and U19021 (N_19021,N_17876,N_17207);
xnor U19022 (N_19022,N_16434,N_17569);
and U19023 (N_19023,N_17934,N_17576);
xor U19024 (N_19024,N_16174,N_16258);
xnor U19025 (N_19025,N_17762,N_17482);
nor U19026 (N_19026,N_16817,N_17446);
and U19027 (N_19027,N_17846,N_16954);
nand U19028 (N_19028,N_17209,N_17838);
or U19029 (N_19029,N_16735,N_17616);
nand U19030 (N_19030,N_17478,N_17862);
and U19031 (N_19031,N_16426,N_16174);
nand U19032 (N_19032,N_17766,N_17250);
and U19033 (N_19033,N_16527,N_16852);
or U19034 (N_19034,N_17740,N_17894);
and U19035 (N_19035,N_17324,N_16254);
nor U19036 (N_19036,N_16632,N_16696);
nand U19037 (N_19037,N_17369,N_17935);
or U19038 (N_19038,N_17436,N_17028);
or U19039 (N_19039,N_16799,N_16175);
or U19040 (N_19040,N_16630,N_17138);
or U19041 (N_19041,N_16147,N_17177);
xor U19042 (N_19042,N_16794,N_17363);
and U19043 (N_19043,N_16040,N_16024);
nor U19044 (N_19044,N_17492,N_17013);
or U19045 (N_19045,N_17919,N_16315);
and U19046 (N_19046,N_16592,N_17786);
xnor U19047 (N_19047,N_16092,N_17171);
xnor U19048 (N_19048,N_16717,N_16675);
nor U19049 (N_19049,N_16035,N_17393);
nand U19050 (N_19050,N_16467,N_17661);
nand U19051 (N_19051,N_16008,N_16046);
or U19052 (N_19052,N_16674,N_17149);
and U19053 (N_19053,N_16478,N_17656);
or U19054 (N_19054,N_16617,N_17971);
or U19055 (N_19055,N_17306,N_17556);
nand U19056 (N_19056,N_16384,N_16540);
nand U19057 (N_19057,N_16879,N_16557);
nand U19058 (N_19058,N_17194,N_16223);
nand U19059 (N_19059,N_17855,N_16699);
nand U19060 (N_19060,N_16409,N_17187);
or U19061 (N_19061,N_16866,N_17225);
nor U19062 (N_19062,N_17966,N_16152);
and U19063 (N_19063,N_16996,N_16732);
and U19064 (N_19064,N_16473,N_17730);
xnor U19065 (N_19065,N_17046,N_17563);
xnor U19066 (N_19066,N_17748,N_17167);
and U19067 (N_19067,N_16310,N_16771);
and U19068 (N_19068,N_16264,N_16912);
nor U19069 (N_19069,N_16966,N_17873);
or U19070 (N_19070,N_16714,N_17470);
or U19071 (N_19071,N_17758,N_17060);
and U19072 (N_19072,N_17746,N_17868);
or U19073 (N_19073,N_17450,N_17215);
and U19074 (N_19074,N_17126,N_16342);
and U19075 (N_19075,N_17338,N_16548);
nand U19076 (N_19076,N_17365,N_16628);
nand U19077 (N_19077,N_16616,N_16572);
nor U19078 (N_19078,N_17342,N_17656);
nand U19079 (N_19079,N_17239,N_17091);
nand U19080 (N_19080,N_16108,N_16303);
nor U19081 (N_19081,N_17809,N_17511);
nor U19082 (N_19082,N_16151,N_17075);
or U19083 (N_19083,N_17165,N_16091);
nand U19084 (N_19084,N_16737,N_17130);
or U19085 (N_19085,N_16761,N_16470);
and U19086 (N_19086,N_17603,N_17870);
nor U19087 (N_19087,N_16515,N_16263);
xor U19088 (N_19088,N_16032,N_17047);
or U19089 (N_19089,N_17297,N_17724);
and U19090 (N_19090,N_17725,N_17591);
nand U19091 (N_19091,N_16724,N_16486);
xnor U19092 (N_19092,N_17297,N_16826);
and U19093 (N_19093,N_16535,N_17030);
nor U19094 (N_19094,N_16369,N_16641);
and U19095 (N_19095,N_17629,N_16679);
and U19096 (N_19096,N_17323,N_17973);
or U19097 (N_19097,N_16217,N_16699);
nor U19098 (N_19098,N_17274,N_16240);
nor U19099 (N_19099,N_16611,N_17480);
and U19100 (N_19100,N_16968,N_17605);
and U19101 (N_19101,N_16992,N_16284);
or U19102 (N_19102,N_16767,N_16727);
and U19103 (N_19103,N_16197,N_16213);
and U19104 (N_19104,N_17195,N_16996);
nand U19105 (N_19105,N_16180,N_17994);
xor U19106 (N_19106,N_17712,N_16384);
nor U19107 (N_19107,N_17334,N_17378);
nand U19108 (N_19108,N_17280,N_16288);
nor U19109 (N_19109,N_17784,N_16939);
and U19110 (N_19110,N_17968,N_17088);
and U19111 (N_19111,N_17235,N_16303);
nor U19112 (N_19112,N_17404,N_16556);
or U19113 (N_19113,N_17549,N_16019);
nand U19114 (N_19114,N_16755,N_16326);
nor U19115 (N_19115,N_17167,N_17021);
and U19116 (N_19116,N_16022,N_17668);
nand U19117 (N_19117,N_16899,N_16890);
nand U19118 (N_19118,N_17796,N_17177);
and U19119 (N_19119,N_16759,N_17741);
and U19120 (N_19120,N_16012,N_16122);
and U19121 (N_19121,N_16603,N_16860);
or U19122 (N_19122,N_16949,N_16978);
nor U19123 (N_19123,N_16015,N_17082);
nor U19124 (N_19124,N_17375,N_17613);
and U19125 (N_19125,N_16972,N_17706);
or U19126 (N_19126,N_16521,N_17220);
xnor U19127 (N_19127,N_16499,N_16591);
nand U19128 (N_19128,N_16562,N_17015);
nor U19129 (N_19129,N_16974,N_16639);
nor U19130 (N_19130,N_16748,N_17151);
and U19131 (N_19131,N_16854,N_16399);
and U19132 (N_19132,N_16942,N_16615);
or U19133 (N_19133,N_17500,N_16091);
nor U19134 (N_19134,N_17872,N_17699);
nor U19135 (N_19135,N_17540,N_16698);
and U19136 (N_19136,N_17196,N_17646);
or U19137 (N_19137,N_16685,N_17961);
or U19138 (N_19138,N_16663,N_17801);
nand U19139 (N_19139,N_17597,N_17385);
nand U19140 (N_19140,N_16342,N_16709);
xnor U19141 (N_19141,N_17128,N_16338);
and U19142 (N_19142,N_17929,N_17032);
nor U19143 (N_19143,N_17365,N_17260);
nand U19144 (N_19144,N_17633,N_17029);
xor U19145 (N_19145,N_16558,N_16539);
and U19146 (N_19146,N_16669,N_16874);
and U19147 (N_19147,N_17189,N_16996);
or U19148 (N_19148,N_16563,N_16906);
and U19149 (N_19149,N_17595,N_16104);
nand U19150 (N_19150,N_16398,N_16695);
or U19151 (N_19151,N_17699,N_16742);
and U19152 (N_19152,N_17537,N_16298);
nor U19153 (N_19153,N_17590,N_16109);
xnor U19154 (N_19154,N_17215,N_16583);
xnor U19155 (N_19155,N_17901,N_16398);
nor U19156 (N_19156,N_16512,N_16575);
or U19157 (N_19157,N_17932,N_17906);
and U19158 (N_19158,N_16839,N_17088);
nor U19159 (N_19159,N_17681,N_17804);
or U19160 (N_19160,N_16054,N_17523);
or U19161 (N_19161,N_17537,N_16514);
or U19162 (N_19162,N_17584,N_16612);
nand U19163 (N_19163,N_17924,N_16374);
nand U19164 (N_19164,N_16212,N_16597);
and U19165 (N_19165,N_16555,N_17526);
nand U19166 (N_19166,N_16664,N_16757);
nand U19167 (N_19167,N_16565,N_17213);
xor U19168 (N_19168,N_16352,N_17453);
or U19169 (N_19169,N_16639,N_16535);
or U19170 (N_19170,N_16252,N_17496);
nor U19171 (N_19171,N_17983,N_17156);
nor U19172 (N_19172,N_16300,N_16707);
xnor U19173 (N_19173,N_16733,N_17583);
xnor U19174 (N_19174,N_16908,N_17933);
or U19175 (N_19175,N_16030,N_17661);
or U19176 (N_19176,N_16267,N_17816);
nand U19177 (N_19177,N_16573,N_17529);
or U19178 (N_19178,N_16790,N_16184);
xnor U19179 (N_19179,N_16865,N_17835);
or U19180 (N_19180,N_16652,N_17813);
or U19181 (N_19181,N_16622,N_17271);
nand U19182 (N_19182,N_16525,N_17850);
nor U19183 (N_19183,N_17536,N_16784);
or U19184 (N_19184,N_17378,N_16895);
nand U19185 (N_19185,N_16091,N_17439);
or U19186 (N_19186,N_17495,N_16835);
nor U19187 (N_19187,N_16461,N_16698);
and U19188 (N_19188,N_16779,N_16411);
or U19189 (N_19189,N_17131,N_17107);
and U19190 (N_19190,N_16706,N_16496);
or U19191 (N_19191,N_17016,N_17796);
or U19192 (N_19192,N_16441,N_17113);
nor U19193 (N_19193,N_16174,N_16574);
and U19194 (N_19194,N_17686,N_17309);
nand U19195 (N_19195,N_16008,N_17307);
nand U19196 (N_19196,N_17104,N_16334);
xnor U19197 (N_19197,N_16911,N_17321);
xnor U19198 (N_19198,N_16116,N_17068);
nand U19199 (N_19199,N_17690,N_16981);
and U19200 (N_19200,N_16039,N_16289);
xnor U19201 (N_19201,N_17117,N_16736);
or U19202 (N_19202,N_16175,N_16323);
or U19203 (N_19203,N_16811,N_16216);
and U19204 (N_19204,N_17327,N_17040);
or U19205 (N_19205,N_17860,N_16553);
xor U19206 (N_19206,N_17097,N_17237);
or U19207 (N_19207,N_17377,N_16965);
nor U19208 (N_19208,N_17177,N_16862);
or U19209 (N_19209,N_17131,N_16813);
nand U19210 (N_19210,N_17966,N_17609);
or U19211 (N_19211,N_17043,N_16830);
and U19212 (N_19212,N_16522,N_17523);
nor U19213 (N_19213,N_17812,N_16906);
nand U19214 (N_19214,N_16825,N_16979);
and U19215 (N_19215,N_17148,N_16618);
or U19216 (N_19216,N_16410,N_17752);
and U19217 (N_19217,N_16173,N_16143);
and U19218 (N_19218,N_16928,N_17817);
nand U19219 (N_19219,N_16840,N_16945);
and U19220 (N_19220,N_16496,N_17384);
nor U19221 (N_19221,N_17287,N_17641);
or U19222 (N_19222,N_16834,N_17405);
nand U19223 (N_19223,N_16926,N_16943);
and U19224 (N_19224,N_16655,N_17785);
xnor U19225 (N_19225,N_17306,N_16819);
nor U19226 (N_19226,N_17916,N_16018);
nand U19227 (N_19227,N_16495,N_17455);
xor U19228 (N_19228,N_16648,N_16654);
and U19229 (N_19229,N_16364,N_16279);
and U19230 (N_19230,N_16344,N_17151);
nand U19231 (N_19231,N_17131,N_17346);
and U19232 (N_19232,N_17104,N_17368);
or U19233 (N_19233,N_17589,N_17925);
or U19234 (N_19234,N_16885,N_16523);
and U19235 (N_19235,N_16890,N_17025);
nor U19236 (N_19236,N_17142,N_17776);
nor U19237 (N_19237,N_17550,N_17126);
and U19238 (N_19238,N_16315,N_17564);
or U19239 (N_19239,N_16131,N_16469);
or U19240 (N_19240,N_17515,N_17248);
and U19241 (N_19241,N_17753,N_17288);
nor U19242 (N_19242,N_17534,N_17949);
and U19243 (N_19243,N_16180,N_16620);
xnor U19244 (N_19244,N_17413,N_17833);
nor U19245 (N_19245,N_17785,N_17526);
or U19246 (N_19246,N_16806,N_17954);
xnor U19247 (N_19247,N_17269,N_17909);
nand U19248 (N_19248,N_17509,N_16758);
and U19249 (N_19249,N_17007,N_17907);
and U19250 (N_19250,N_16147,N_16667);
or U19251 (N_19251,N_16803,N_16069);
and U19252 (N_19252,N_16887,N_16337);
and U19253 (N_19253,N_16380,N_17588);
xor U19254 (N_19254,N_16275,N_16798);
nor U19255 (N_19255,N_17739,N_17350);
or U19256 (N_19256,N_16293,N_16694);
and U19257 (N_19257,N_16257,N_17079);
nor U19258 (N_19258,N_16724,N_16286);
nand U19259 (N_19259,N_17240,N_17704);
nand U19260 (N_19260,N_17808,N_17833);
and U19261 (N_19261,N_16757,N_17929);
nand U19262 (N_19262,N_16926,N_17380);
and U19263 (N_19263,N_16150,N_16697);
nand U19264 (N_19264,N_16702,N_17398);
and U19265 (N_19265,N_16990,N_17760);
nand U19266 (N_19266,N_16339,N_17741);
nor U19267 (N_19267,N_16477,N_16442);
or U19268 (N_19268,N_16139,N_16967);
or U19269 (N_19269,N_16050,N_16798);
nor U19270 (N_19270,N_17414,N_17454);
nor U19271 (N_19271,N_16395,N_16027);
xor U19272 (N_19272,N_16316,N_17164);
nor U19273 (N_19273,N_16492,N_16708);
nor U19274 (N_19274,N_16805,N_16367);
nand U19275 (N_19275,N_17673,N_17807);
and U19276 (N_19276,N_17670,N_16586);
or U19277 (N_19277,N_17388,N_17650);
and U19278 (N_19278,N_17712,N_17388);
nor U19279 (N_19279,N_17871,N_16056);
xor U19280 (N_19280,N_16096,N_17777);
or U19281 (N_19281,N_16077,N_16061);
and U19282 (N_19282,N_17892,N_16602);
and U19283 (N_19283,N_17657,N_17600);
nand U19284 (N_19284,N_17772,N_17295);
nand U19285 (N_19285,N_17151,N_16176);
or U19286 (N_19286,N_16286,N_16870);
and U19287 (N_19287,N_16434,N_16046);
nor U19288 (N_19288,N_16773,N_16087);
xor U19289 (N_19289,N_17606,N_16049);
and U19290 (N_19290,N_17295,N_17962);
or U19291 (N_19291,N_16898,N_16863);
or U19292 (N_19292,N_17290,N_17318);
and U19293 (N_19293,N_17914,N_17967);
and U19294 (N_19294,N_16160,N_17313);
or U19295 (N_19295,N_16282,N_16766);
nand U19296 (N_19296,N_16292,N_16057);
nand U19297 (N_19297,N_16636,N_17926);
nand U19298 (N_19298,N_17804,N_16509);
and U19299 (N_19299,N_16070,N_17942);
or U19300 (N_19300,N_16770,N_17610);
nor U19301 (N_19301,N_17283,N_17934);
and U19302 (N_19302,N_17662,N_16428);
and U19303 (N_19303,N_17305,N_17204);
xor U19304 (N_19304,N_16403,N_16335);
and U19305 (N_19305,N_17992,N_17388);
and U19306 (N_19306,N_17417,N_17906);
nor U19307 (N_19307,N_17727,N_16560);
nand U19308 (N_19308,N_17251,N_17037);
nor U19309 (N_19309,N_17035,N_17983);
nand U19310 (N_19310,N_17112,N_16786);
or U19311 (N_19311,N_16741,N_16901);
nand U19312 (N_19312,N_17976,N_17730);
nor U19313 (N_19313,N_16759,N_16317);
nor U19314 (N_19314,N_17179,N_16759);
and U19315 (N_19315,N_17669,N_16360);
nor U19316 (N_19316,N_16086,N_16342);
and U19317 (N_19317,N_17989,N_17504);
nor U19318 (N_19318,N_16956,N_17731);
nand U19319 (N_19319,N_16457,N_16756);
or U19320 (N_19320,N_17314,N_17575);
and U19321 (N_19321,N_16314,N_17230);
or U19322 (N_19322,N_17059,N_17519);
and U19323 (N_19323,N_17730,N_17881);
or U19324 (N_19324,N_16458,N_16232);
or U19325 (N_19325,N_16753,N_16280);
xnor U19326 (N_19326,N_16085,N_17011);
xor U19327 (N_19327,N_17975,N_17784);
nor U19328 (N_19328,N_16780,N_17509);
xnor U19329 (N_19329,N_16707,N_16442);
xnor U19330 (N_19330,N_16167,N_16169);
xnor U19331 (N_19331,N_16970,N_17624);
xnor U19332 (N_19332,N_16920,N_16557);
nand U19333 (N_19333,N_17821,N_16066);
nor U19334 (N_19334,N_17307,N_17033);
nand U19335 (N_19335,N_17100,N_17857);
nand U19336 (N_19336,N_16575,N_17218);
nand U19337 (N_19337,N_16450,N_16460);
nor U19338 (N_19338,N_17831,N_16930);
and U19339 (N_19339,N_16560,N_17104);
or U19340 (N_19340,N_17966,N_16170);
and U19341 (N_19341,N_16629,N_16908);
or U19342 (N_19342,N_16642,N_16556);
or U19343 (N_19343,N_16167,N_16739);
or U19344 (N_19344,N_16755,N_17932);
xor U19345 (N_19345,N_17271,N_16751);
nor U19346 (N_19346,N_17356,N_16417);
or U19347 (N_19347,N_16872,N_16933);
and U19348 (N_19348,N_16906,N_17339);
or U19349 (N_19349,N_17978,N_16455);
nor U19350 (N_19350,N_16209,N_17084);
nor U19351 (N_19351,N_17862,N_17481);
nand U19352 (N_19352,N_16974,N_17334);
xnor U19353 (N_19353,N_17128,N_16088);
nor U19354 (N_19354,N_16716,N_17175);
nor U19355 (N_19355,N_16330,N_16474);
nand U19356 (N_19356,N_16708,N_16583);
and U19357 (N_19357,N_17285,N_17850);
nor U19358 (N_19358,N_16471,N_17168);
nor U19359 (N_19359,N_16443,N_17129);
nand U19360 (N_19360,N_17516,N_16884);
and U19361 (N_19361,N_17018,N_17716);
nor U19362 (N_19362,N_16683,N_17226);
nor U19363 (N_19363,N_17576,N_16166);
nor U19364 (N_19364,N_17862,N_16419);
nand U19365 (N_19365,N_16001,N_16597);
nand U19366 (N_19366,N_16093,N_16885);
nand U19367 (N_19367,N_16117,N_17258);
or U19368 (N_19368,N_17278,N_16185);
nand U19369 (N_19369,N_16210,N_16703);
nand U19370 (N_19370,N_16651,N_16362);
and U19371 (N_19371,N_16284,N_17669);
nand U19372 (N_19372,N_17793,N_16526);
nor U19373 (N_19373,N_16222,N_16257);
or U19374 (N_19374,N_16480,N_16649);
and U19375 (N_19375,N_16350,N_17279);
and U19376 (N_19376,N_16374,N_16227);
and U19377 (N_19377,N_17201,N_16992);
or U19378 (N_19378,N_17674,N_16342);
nor U19379 (N_19379,N_16179,N_17160);
nand U19380 (N_19380,N_16920,N_17703);
and U19381 (N_19381,N_17862,N_17686);
nand U19382 (N_19382,N_16446,N_17003);
xnor U19383 (N_19383,N_16593,N_17016);
nand U19384 (N_19384,N_16893,N_16115);
nor U19385 (N_19385,N_16551,N_17813);
nand U19386 (N_19386,N_16573,N_17219);
or U19387 (N_19387,N_17698,N_17165);
xnor U19388 (N_19388,N_16485,N_16544);
xor U19389 (N_19389,N_16060,N_17516);
nor U19390 (N_19390,N_16188,N_16846);
and U19391 (N_19391,N_17656,N_17116);
nand U19392 (N_19392,N_17411,N_17889);
nand U19393 (N_19393,N_16650,N_16310);
nand U19394 (N_19394,N_17491,N_16414);
xor U19395 (N_19395,N_16400,N_16310);
or U19396 (N_19396,N_16559,N_16402);
or U19397 (N_19397,N_16905,N_16909);
and U19398 (N_19398,N_16439,N_16063);
and U19399 (N_19399,N_17151,N_17036);
or U19400 (N_19400,N_17660,N_17860);
nor U19401 (N_19401,N_17023,N_16246);
nand U19402 (N_19402,N_17938,N_17934);
or U19403 (N_19403,N_16402,N_17728);
nor U19404 (N_19404,N_16123,N_17012);
and U19405 (N_19405,N_17150,N_16977);
nor U19406 (N_19406,N_16056,N_16293);
nor U19407 (N_19407,N_17649,N_17029);
nor U19408 (N_19408,N_16260,N_16619);
nor U19409 (N_19409,N_16754,N_17366);
nor U19410 (N_19410,N_16814,N_16965);
nand U19411 (N_19411,N_16439,N_16820);
nand U19412 (N_19412,N_16133,N_16829);
nand U19413 (N_19413,N_17452,N_17228);
nor U19414 (N_19414,N_16049,N_16652);
or U19415 (N_19415,N_16894,N_17574);
xnor U19416 (N_19416,N_17688,N_16025);
or U19417 (N_19417,N_16862,N_16322);
nand U19418 (N_19418,N_17311,N_16567);
and U19419 (N_19419,N_17108,N_17805);
nand U19420 (N_19420,N_17216,N_17451);
and U19421 (N_19421,N_17709,N_17012);
nand U19422 (N_19422,N_16531,N_17818);
nor U19423 (N_19423,N_16851,N_17802);
nor U19424 (N_19424,N_17870,N_16900);
or U19425 (N_19425,N_16571,N_17096);
or U19426 (N_19426,N_17897,N_17525);
and U19427 (N_19427,N_17147,N_16624);
xnor U19428 (N_19428,N_16779,N_16891);
nor U19429 (N_19429,N_17360,N_16309);
nor U19430 (N_19430,N_16907,N_16247);
and U19431 (N_19431,N_17976,N_17022);
nor U19432 (N_19432,N_17183,N_16588);
nand U19433 (N_19433,N_17458,N_16001);
xor U19434 (N_19434,N_16141,N_17880);
or U19435 (N_19435,N_17781,N_17558);
nand U19436 (N_19436,N_16111,N_16008);
or U19437 (N_19437,N_17131,N_16403);
nor U19438 (N_19438,N_17670,N_17695);
or U19439 (N_19439,N_16111,N_16993);
xor U19440 (N_19440,N_17876,N_17859);
xor U19441 (N_19441,N_16015,N_17274);
nand U19442 (N_19442,N_16142,N_17221);
nand U19443 (N_19443,N_17317,N_16715);
and U19444 (N_19444,N_16651,N_17879);
nand U19445 (N_19445,N_16469,N_17728);
nor U19446 (N_19446,N_16943,N_16483);
and U19447 (N_19447,N_16393,N_16352);
nand U19448 (N_19448,N_17744,N_17278);
nand U19449 (N_19449,N_16729,N_16891);
nand U19450 (N_19450,N_17106,N_16538);
xnor U19451 (N_19451,N_16139,N_17671);
or U19452 (N_19452,N_16646,N_16521);
or U19453 (N_19453,N_16014,N_17414);
or U19454 (N_19454,N_17432,N_17039);
or U19455 (N_19455,N_17728,N_17973);
and U19456 (N_19456,N_17019,N_16015);
nor U19457 (N_19457,N_17620,N_16473);
and U19458 (N_19458,N_17829,N_16575);
nand U19459 (N_19459,N_16809,N_17489);
and U19460 (N_19460,N_16851,N_16156);
nor U19461 (N_19461,N_16611,N_17053);
xnor U19462 (N_19462,N_16685,N_16939);
nor U19463 (N_19463,N_16649,N_17201);
nor U19464 (N_19464,N_17737,N_17307);
nand U19465 (N_19465,N_16840,N_17416);
and U19466 (N_19466,N_17616,N_16083);
or U19467 (N_19467,N_16689,N_17264);
nand U19468 (N_19468,N_16503,N_17415);
nand U19469 (N_19469,N_16764,N_17519);
or U19470 (N_19470,N_16822,N_16825);
or U19471 (N_19471,N_16225,N_16211);
xnor U19472 (N_19472,N_16921,N_17458);
xor U19473 (N_19473,N_17502,N_17309);
nand U19474 (N_19474,N_16853,N_17167);
nor U19475 (N_19475,N_16033,N_16073);
nor U19476 (N_19476,N_17428,N_16681);
nand U19477 (N_19477,N_16526,N_16012);
or U19478 (N_19478,N_17648,N_17382);
xor U19479 (N_19479,N_16249,N_17717);
and U19480 (N_19480,N_16595,N_17924);
or U19481 (N_19481,N_16347,N_17502);
nand U19482 (N_19482,N_16395,N_17634);
nand U19483 (N_19483,N_17466,N_16687);
and U19484 (N_19484,N_17714,N_16313);
nor U19485 (N_19485,N_17599,N_16453);
or U19486 (N_19486,N_16034,N_16529);
nor U19487 (N_19487,N_16212,N_17665);
and U19488 (N_19488,N_17764,N_16918);
xor U19489 (N_19489,N_17083,N_16545);
and U19490 (N_19490,N_16490,N_16739);
nand U19491 (N_19491,N_17408,N_16945);
or U19492 (N_19492,N_16815,N_16655);
nor U19493 (N_19493,N_17887,N_17503);
nand U19494 (N_19494,N_16846,N_17853);
nand U19495 (N_19495,N_16652,N_17751);
nor U19496 (N_19496,N_16354,N_17189);
xor U19497 (N_19497,N_16336,N_16286);
or U19498 (N_19498,N_16223,N_17292);
nand U19499 (N_19499,N_17610,N_16912);
or U19500 (N_19500,N_16244,N_16147);
nor U19501 (N_19501,N_16002,N_16226);
or U19502 (N_19502,N_16562,N_17356);
or U19503 (N_19503,N_16225,N_17283);
xnor U19504 (N_19504,N_16494,N_17469);
or U19505 (N_19505,N_17293,N_16762);
nor U19506 (N_19506,N_16831,N_17612);
and U19507 (N_19507,N_17176,N_16835);
xnor U19508 (N_19508,N_17946,N_17131);
and U19509 (N_19509,N_16814,N_16818);
xnor U19510 (N_19510,N_16981,N_17188);
nand U19511 (N_19511,N_17273,N_16245);
and U19512 (N_19512,N_17799,N_16139);
nand U19513 (N_19513,N_16041,N_16662);
nand U19514 (N_19514,N_16763,N_16639);
and U19515 (N_19515,N_17494,N_17953);
nor U19516 (N_19516,N_17066,N_17980);
or U19517 (N_19517,N_17900,N_16766);
and U19518 (N_19518,N_17586,N_16088);
or U19519 (N_19519,N_16646,N_16283);
nand U19520 (N_19520,N_16653,N_17518);
nor U19521 (N_19521,N_17727,N_16230);
and U19522 (N_19522,N_16498,N_17794);
nor U19523 (N_19523,N_16689,N_16921);
and U19524 (N_19524,N_16414,N_17076);
or U19525 (N_19525,N_17381,N_17426);
xnor U19526 (N_19526,N_17783,N_16609);
or U19527 (N_19527,N_16054,N_17452);
or U19528 (N_19528,N_16050,N_17043);
or U19529 (N_19529,N_16340,N_16458);
nor U19530 (N_19530,N_17400,N_17902);
or U19531 (N_19531,N_16367,N_16765);
nor U19532 (N_19532,N_17623,N_17032);
nor U19533 (N_19533,N_17579,N_16084);
nand U19534 (N_19534,N_16675,N_17975);
and U19535 (N_19535,N_16274,N_16719);
nand U19536 (N_19536,N_16624,N_17225);
xor U19537 (N_19537,N_16228,N_17050);
xor U19538 (N_19538,N_16890,N_17963);
nand U19539 (N_19539,N_17003,N_16566);
or U19540 (N_19540,N_17270,N_16492);
nand U19541 (N_19541,N_17474,N_17338);
or U19542 (N_19542,N_17683,N_17328);
xor U19543 (N_19543,N_16960,N_17918);
nand U19544 (N_19544,N_17659,N_16174);
and U19545 (N_19545,N_17306,N_17805);
and U19546 (N_19546,N_16005,N_17155);
and U19547 (N_19547,N_17071,N_16842);
or U19548 (N_19548,N_16375,N_16435);
or U19549 (N_19549,N_17718,N_17138);
nor U19550 (N_19550,N_16686,N_16076);
nor U19551 (N_19551,N_16534,N_17296);
nand U19552 (N_19552,N_17367,N_16344);
nor U19553 (N_19553,N_17940,N_17455);
or U19554 (N_19554,N_16502,N_17630);
or U19555 (N_19555,N_17855,N_17195);
or U19556 (N_19556,N_16651,N_16790);
nor U19557 (N_19557,N_17297,N_16049);
and U19558 (N_19558,N_17077,N_17121);
nand U19559 (N_19559,N_16470,N_16270);
nor U19560 (N_19560,N_17739,N_17573);
nor U19561 (N_19561,N_17568,N_16575);
and U19562 (N_19562,N_16180,N_16675);
nand U19563 (N_19563,N_16394,N_17056);
and U19564 (N_19564,N_17766,N_16412);
and U19565 (N_19565,N_17780,N_17751);
and U19566 (N_19566,N_17193,N_17840);
xnor U19567 (N_19567,N_16410,N_16228);
or U19568 (N_19568,N_17014,N_17000);
and U19569 (N_19569,N_17255,N_16819);
nand U19570 (N_19570,N_17681,N_16911);
nand U19571 (N_19571,N_16209,N_16164);
nand U19572 (N_19572,N_17051,N_16269);
nand U19573 (N_19573,N_16704,N_17524);
nor U19574 (N_19574,N_16897,N_16060);
or U19575 (N_19575,N_16862,N_16216);
and U19576 (N_19576,N_17738,N_17592);
or U19577 (N_19577,N_16524,N_16179);
and U19578 (N_19578,N_16802,N_16786);
nand U19579 (N_19579,N_16940,N_17884);
nor U19580 (N_19580,N_16676,N_17444);
nor U19581 (N_19581,N_16522,N_17927);
or U19582 (N_19582,N_16005,N_17531);
and U19583 (N_19583,N_16034,N_16668);
and U19584 (N_19584,N_16414,N_17043);
nor U19585 (N_19585,N_17243,N_16486);
or U19586 (N_19586,N_17570,N_17877);
or U19587 (N_19587,N_16589,N_17109);
or U19588 (N_19588,N_16831,N_16163);
nand U19589 (N_19589,N_17345,N_16702);
nand U19590 (N_19590,N_17530,N_16170);
nor U19591 (N_19591,N_16655,N_17246);
nand U19592 (N_19592,N_17469,N_16733);
or U19593 (N_19593,N_17041,N_17096);
and U19594 (N_19594,N_17093,N_16913);
xor U19595 (N_19595,N_16713,N_17557);
xnor U19596 (N_19596,N_17976,N_16811);
nor U19597 (N_19597,N_16649,N_16736);
xnor U19598 (N_19598,N_16434,N_17490);
xnor U19599 (N_19599,N_16815,N_16764);
and U19600 (N_19600,N_17552,N_16572);
nor U19601 (N_19601,N_16797,N_16349);
nor U19602 (N_19602,N_16822,N_16761);
or U19603 (N_19603,N_17841,N_16154);
nand U19604 (N_19604,N_16751,N_17829);
nor U19605 (N_19605,N_16062,N_17649);
nor U19606 (N_19606,N_17061,N_17005);
nand U19607 (N_19607,N_16942,N_17208);
and U19608 (N_19608,N_16603,N_17414);
nor U19609 (N_19609,N_16848,N_17470);
nor U19610 (N_19610,N_16645,N_16303);
nor U19611 (N_19611,N_16519,N_16180);
or U19612 (N_19612,N_16417,N_17313);
nor U19613 (N_19613,N_16810,N_17240);
and U19614 (N_19614,N_16171,N_16126);
nand U19615 (N_19615,N_16604,N_17677);
and U19616 (N_19616,N_16060,N_16963);
nor U19617 (N_19617,N_16559,N_17730);
or U19618 (N_19618,N_16965,N_17785);
nor U19619 (N_19619,N_17445,N_17027);
and U19620 (N_19620,N_16059,N_17969);
nand U19621 (N_19621,N_17757,N_16878);
or U19622 (N_19622,N_17816,N_17125);
and U19623 (N_19623,N_17451,N_16986);
nor U19624 (N_19624,N_16950,N_17270);
or U19625 (N_19625,N_17782,N_16855);
nand U19626 (N_19626,N_17924,N_17046);
and U19627 (N_19627,N_17581,N_17900);
and U19628 (N_19628,N_16168,N_17572);
nand U19629 (N_19629,N_16089,N_17952);
and U19630 (N_19630,N_16098,N_17585);
or U19631 (N_19631,N_17623,N_16518);
nor U19632 (N_19632,N_17383,N_16001);
and U19633 (N_19633,N_16922,N_17773);
or U19634 (N_19634,N_17319,N_16206);
and U19635 (N_19635,N_16077,N_16297);
or U19636 (N_19636,N_16124,N_17211);
or U19637 (N_19637,N_17871,N_16939);
nand U19638 (N_19638,N_17866,N_16737);
xor U19639 (N_19639,N_16821,N_16387);
nor U19640 (N_19640,N_16000,N_17934);
and U19641 (N_19641,N_17403,N_17215);
or U19642 (N_19642,N_17725,N_17360);
nor U19643 (N_19643,N_16254,N_16092);
nor U19644 (N_19644,N_16313,N_16907);
nor U19645 (N_19645,N_17571,N_16434);
or U19646 (N_19646,N_17420,N_17676);
xor U19647 (N_19647,N_16403,N_17239);
nand U19648 (N_19648,N_17659,N_17653);
and U19649 (N_19649,N_16047,N_16415);
and U19650 (N_19650,N_16930,N_17033);
nand U19651 (N_19651,N_16083,N_16962);
nand U19652 (N_19652,N_17482,N_16595);
nand U19653 (N_19653,N_17402,N_16863);
or U19654 (N_19654,N_16919,N_16503);
nor U19655 (N_19655,N_17489,N_16307);
nand U19656 (N_19656,N_17645,N_16428);
xor U19657 (N_19657,N_16119,N_17082);
or U19658 (N_19658,N_17029,N_16188);
and U19659 (N_19659,N_17557,N_16827);
nand U19660 (N_19660,N_16124,N_17521);
xnor U19661 (N_19661,N_17406,N_17437);
or U19662 (N_19662,N_16568,N_16962);
nand U19663 (N_19663,N_17475,N_16213);
nand U19664 (N_19664,N_17369,N_17842);
nor U19665 (N_19665,N_16288,N_16528);
nand U19666 (N_19666,N_16470,N_16969);
nand U19667 (N_19667,N_16855,N_16448);
nor U19668 (N_19668,N_17322,N_16787);
and U19669 (N_19669,N_16248,N_17803);
or U19670 (N_19670,N_16153,N_16301);
and U19671 (N_19671,N_17506,N_16057);
nand U19672 (N_19672,N_17064,N_17462);
and U19673 (N_19673,N_16972,N_17367);
nor U19674 (N_19674,N_17067,N_17093);
and U19675 (N_19675,N_17123,N_16328);
nand U19676 (N_19676,N_16976,N_17001);
nor U19677 (N_19677,N_16407,N_17771);
nor U19678 (N_19678,N_16968,N_16857);
nand U19679 (N_19679,N_16883,N_16499);
nand U19680 (N_19680,N_16414,N_16720);
or U19681 (N_19681,N_16908,N_17878);
nand U19682 (N_19682,N_16063,N_16295);
xnor U19683 (N_19683,N_17425,N_16631);
and U19684 (N_19684,N_17719,N_17862);
nand U19685 (N_19685,N_16334,N_17468);
or U19686 (N_19686,N_16840,N_16862);
nor U19687 (N_19687,N_17790,N_17398);
nand U19688 (N_19688,N_16190,N_16048);
nor U19689 (N_19689,N_16902,N_17062);
xnor U19690 (N_19690,N_17075,N_16237);
xor U19691 (N_19691,N_16732,N_16295);
and U19692 (N_19692,N_16340,N_16179);
and U19693 (N_19693,N_16887,N_16651);
nand U19694 (N_19694,N_17214,N_17425);
nor U19695 (N_19695,N_17357,N_17220);
nand U19696 (N_19696,N_16688,N_16742);
nor U19697 (N_19697,N_16452,N_16883);
nand U19698 (N_19698,N_16804,N_16234);
nand U19699 (N_19699,N_17098,N_16957);
or U19700 (N_19700,N_17142,N_17977);
or U19701 (N_19701,N_17086,N_16239);
or U19702 (N_19702,N_16829,N_16951);
xor U19703 (N_19703,N_17942,N_16002);
and U19704 (N_19704,N_17215,N_16314);
or U19705 (N_19705,N_17910,N_17232);
and U19706 (N_19706,N_16971,N_16663);
nor U19707 (N_19707,N_17146,N_16228);
xor U19708 (N_19708,N_16845,N_16862);
nand U19709 (N_19709,N_16975,N_17275);
nor U19710 (N_19710,N_16911,N_17699);
nor U19711 (N_19711,N_16900,N_16839);
and U19712 (N_19712,N_16177,N_17708);
nor U19713 (N_19713,N_16290,N_17241);
nor U19714 (N_19714,N_17572,N_16710);
and U19715 (N_19715,N_16242,N_17121);
xnor U19716 (N_19716,N_17421,N_17924);
xnor U19717 (N_19717,N_17894,N_17212);
nor U19718 (N_19718,N_16769,N_17282);
nor U19719 (N_19719,N_17927,N_17340);
and U19720 (N_19720,N_16905,N_16108);
nor U19721 (N_19721,N_16737,N_16040);
nor U19722 (N_19722,N_17654,N_17097);
nand U19723 (N_19723,N_16747,N_17216);
nand U19724 (N_19724,N_16851,N_17378);
or U19725 (N_19725,N_16373,N_17192);
and U19726 (N_19726,N_16514,N_17877);
or U19727 (N_19727,N_17236,N_16739);
xnor U19728 (N_19728,N_17130,N_16755);
xor U19729 (N_19729,N_17682,N_17154);
nor U19730 (N_19730,N_16266,N_16004);
and U19731 (N_19731,N_16824,N_17910);
or U19732 (N_19732,N_16550,N_17164);
nand U19733 (N_19733,N_16680,N_16765);
nor U19734 (N_19734,N_16502,N_17204);
and U19735 (N_19735,N_17575,N_16274);
nor U19736 (N_19736,N_16231,N_16506);
or U19737 (N_19737,N_17515,N_17012);
nand U19738 (N_19738,N_16113,N_17891);
xor U19739 (N_19739,N_16159,N_16441);
or U19740 (N_19740,N_16731,N_16240);
and U19741 (N_19741,N_17045,N_16871);
nand U19742 (N_19742,N_16724,N_16244);
xor U19743 (N_19743,N_16436,N_16560);
nand U19744 (N_19744,N_16840,N_16078);
and U19745 (N_19745,N_17673,N_16665);
and U19746 (N_19746,N_16159,N_16520);
nor U19747 (N_19747,N_17291,N_17175);
or U19748 (N_19748,N_17242,N_16211);
nor U19749 (N_19749,N_16707,N_16480);
nor U19750 (N_19750,N_17432,N_16526);
or U19751 (N_19751,N_16809,N_16375);
nor U19752 (N_19752,N_16078,N_17635);
xor U19753 (N_19753,N_17188,N_16298);
or U19754 (N_19754,N_17917,N_17115);
nor U19755 (N_19755,N_17810,N_17158);
nor U19756 (N_19756,N_16912,N_17491);
nand U19757 (N_19757,N_16758,N_17604);
and U19758 (N_19758,N_16172,N_17311);
nand U19759 (N_19759,N_17748,N_17350);
and U19760 (N_19760,N_16584,N_16752);
and U19761 (N_19761,N_16395,N_16030);
or U19762 (N_19762,N_16892,N_16454);
xnor U19763 (N_19763,N_16450,N_16128);
nor U19764 (N_19764,N_16118,N_17204);
and U19765 (N_19765,N_16085,N_16433);
nand U19766 (N_19766,N_17122,N_17323);
xnor U19767 (N_19767,N_17282,N_17443);
nor U19768 (N_19768,N_16526,N_16899);
nor U19769 (N_19769,N_16502,N_17394);
or U19770 (N_19770,N_16515,N_17020);
or U19771 (N_19771,N_16610,N_16085);
nand U19772 (N_19772,N_17669,N_16890);
nand U19773 (N_19773,N_16269,N_16875);
nand U19774 (N_19774,N_16078,N_16302);
and U19775 (N_19775,N_16569,N_16386);
and U19776 (N_19776,N_16919,N_17129);
or U19777 (N_19777,N_17580,N_17834);
nand U19778 (N_19778,N_17928,N_16810);
and U19779 (N_19779,N_16479,N_17203);
nor U19780 (N_19780,N_16417,N_17628);
nand U19781 (N_19781,N_17553,N_16959);
or U19782 (N_19782,N_16782,N_16712);
and U19783 (N_19783,N_17227,N_17176);
and U19784 (N_19784,N_16192,N_17214);
nor U19785 (N_19785,N_16897,N_17570);
nand U19786 (N_19786,N_17305,N_17296);
xnor U19787 (N_19787,N_16494,N_17949);
or U19788 (N_19788,N_17836,N_16079);
xnor U19789 (N_19789,N_17124,N_16948);
nand U19790 (N_19790,N_16787,N_16828);
nand U19791 (N_19791,N_17380,N_17711);
or U19792 (N_19792,N_17294,N_16785);
nor U19793 (N_19793,N_17457,N_17005);
and U19794 (N_19794,N_17186,N_17076);
nand U19795 (N_19795,N_17456,N_17884);
xor U19796 (N_19796,N_17746,N_17870);
xnor U19797 (N_19797,N_16724,N_16118);
or U19798 (N_19798,N_16500,N_16005);
and U19799 (N_19799,N_16229,N_16295);
or U19800 (N_19800,N_16878,N_17088);
nand U19801 (N_19801,N_16515,N_16759);
and U19802 (N_19802,N_17822,N_17631);
nor U19803 (N_19803,N_17566,N_16684);
and U19804 (N_19804,N_16672,N_16216);
and U19805 (N_19805,N_16548,N_16936);
and U19806 (N_19806,N_17571,N_17322);
and U19807 (N_19807,N_16719,N_16843);
nand U19808 (N_19808,N_16404,N_16291);
nor U19809 (N_19809,N_17458,N_16494);
nor U19810 (N_19810,N_16181,N_16914);
or U19811 (N_19811,N_16274,N_16478);
nor U19812 (N_19812,N_17927,N_17702);
and U19813 (N_19813,N_16823,N_16684);
nand U19814 (N_19814,N_16605,N_17807);
nand U19815 (N_19815,N_16690,N_16096);
or U19816 (N_19816,N_17366,N_16787);
nand U19817 (N_19817,N_17565,N_16806);
xor U19818 (N_19818,N_17251,N_17409);
or U19819 (N_19819,N_17094,N_16864);
xnor U19820 (N_19820,N_16980,N_16148);
or U19821 (N_19821,N_16726,N_16493);
nor U19822 (N_19822,N_17080,N_16274);
or U19823 (N_19823,N_16155,N_16900);
nor U19824 (N_19824,N_17317,N_16632);
xnor U19825 (N_19825,N_16970,N_16404);
nand U19826 (N_19826,N_16150,N_17566);
nand U19827 (N_19827,N_16713,N_17507);
or U19828 (N_19828,N_17668,N_16401);
or U19829 (N_19829,N_17931,N_16043);
nor U19830 (N_19830,N_17468,N_17142);
nand U19831 (N_19831,N_16928,N_17216);
nand U19832 (N_19832,N_16189,N_17648);
and U19833 (N_19833,N_16979,N_16188);
or U19834 (N_19834,N_16676,N_16870);
or U19835 (N_19835,N_16588,N_17070);
nand U19836 (N_19836,N_17335,N_16757);
xor U19837 (N_19837,N_16295,N_16342);
or U19838 (N_19838,N_16042,N_16483);
or U19839 (N_19839,N_17304,N_17844);
nor U19840 (N_19840,N_17344,N_17777);
nor U19841 (N_19841,N_16032,N_17933);
and U19842 (N_19842,N_16676,N_17891);
or U19843 (N_19843,N_17764,N_16121);
and U19844 (N_19844,N_16511,N_16889);
nand U19845 (N_19845,N_17902,N_17794);
nor U19846 (N_19846,N_17764,N_16556);
nand U19847 (N_19847,N_16696,N_17600);
or U19848 (N_19848,N_17716,N_17465);
and U19849 (N_19849,N_17167,N_17697);
nor U19850 (N_19850,N_17166,N_16892);
and U19851 (N_19851,N_17755,N_17983);
nor U19852 (N_19852,N_16372,N_16161);
or U19853 (N_19853,N_16447,N_17846);
nor U19854 (N_19854,N_16502,N_16646);
nand U19855 (N_19855,N_17448,N_16769);
nand U19856 (N_19856,N_17124,N_17355);
nand U19857 (N_19857,N_16577,N_16826);
nor U19858 (N_19858,N_16583,N_16343);
and U19859 (N_19859,N_16261,N_17641);
and U19860 (N_19860,N_16164,N_17513);
or U19861 (N_19861,N_17485,N_17579);
and U19862 (N_19862,N_17501,N_16833);
nor U19863 (N_19863,N_17960,N_16421);
nand U19864 (N_19864,N_17636,N_17347);
or U19865 (N_19865,N_17735,N_17196);
nor U19866 (N_19866,N_17167,N_17276);
and U19867 (N_19867,N_17397,N_16845);
or U19868 (N_19868,N_16278,N_17107);
nand U19869 (N_19869,N_16144,N_17432);
and U19870 (N_19870,N_17140,N_17914);
and U19871 (N_19871,N_17721,N_16063);
nand U19872 (N_19872,N_16313,N_17559);
and U19873 (N_19873,N_17218,N_16578);
nor U19874 (N_19874,N_17028,N_17452);
and U19875 (N_19875,N_17690,N_16610);
nor U19876 (N_19876,N_17708,N_16897);
and U19877 (N_19877,N_16662,N_17648);
and U19878 (N_19878,N_17968,N_17610);
xor U19879 (N_19879,N_17157,N_16667);
nand U19880 (N_19880,N_16672,N_17833);
nor U19881 (N_19881,N_16801,N_17038);
xnor U19882 (N_19882,N_17982,N_16600);
or U19883 (N_19883,N_16985,N_17218);
nand U19884 (N_19884,N_17812,N_16004);
nand U19885 (N_19885,N_17011,N_16196);
xor U19886 (N_19886,N_16943,N_17175);
or U19887 (N_19887,N_16447,N_17236);
and U19888 (N_19888,N_16128,N_17001);
and U19889 (N_19889,N_16035,N_16505);
nor U19890 (N_19890,N_16652,N_16346);
nand U19891 (N_19891,N_16799,N_17634);
or U19892 (N_19892,N_17346,N_16890);
nor U19893 (N_19893,N_16206,N_16505);
nor U19894 (N_19894,N_16551,N_16501);
nand U19895 (N_19895,N_17113,N_16126);
and U19896 (N_19896,N_16066,N_16821);
and U19897 (N_19897,N_16993,N_17290);
nor U19898 (N_19898,N_16692,N_16170);
nand U19899 (N_19899,N_16560,N_16863);
nand U19900 (N_19900,N_17378,N_17148);
and U19901 (N_19901,N_17429,N_17416);
nor U19902 (N_19902,N_17209,N_17975);
and U19903 (N_19903,N_17809,N_17077);
and U19904 (N_19904,N_16122,N_16494);
nand U19905 (N_19905,N_16510,N_16190);
and U19906 (N_19906,N_17361,N_16361);
and U19907 (N_19907,N_17100,N_17790);
nor U19908 (N_19908,N_17027,N_17233);
nand U19909 (N_19909,N_17123,N_16941);
nand U19910 (N_19910,N_17335,N_17112);
nand U19911 (N_19911,N_17048,N_17497);
nand U19912 (N_19912,N_16650,N_17442);
and U19913 (N_19913,N_16229,N_16113);
nand U19914 (N_19914,N_16531,N_17794);
or U19915 (N_19915,N_16308,N_17967);
or U19916 (N_19916,N_16741,N_16798);
nor U19917 (N_19917,N_16341,N_17261);
or U19918 (N_19918,N_17522,N_17171);
nand U19919 (N_19919,N_17174,N_17780);
or U19920 (N_19920,N_16504,N_16343);
nor U19921 (N_19921,N_16232,N_17381);
nor U19922 (N_19922,N_16496,N_17366);
or U19923 (N_19923,N_17756,N_16524);
and U19924 (N_19924,N_17591,N_17595);
and U19925 (N_19925,N_17683,N_16916);
or U19926 (N_19926,N_17285,N_16466);
and U19927 (N_19927,N_16822,N_16657);
and U19928 (N_19928,N_17955,N_17744);
or U19929 (N_19929,N_17933,N_16904);
nor U19930 (N_19930,N_17764,N_17956);
nand U19931 (N_19931,N_17899,N_16597);
nand U19932 (N_19932,N_16044,N_16965);
nor U19933 (N_19933,N_16025,N_16148);
xor U19934 (N_19934,N_17756,N_16261);
or U19935 (N_19935,N_17659,N_17065);
or U19936 (N_19936,N_16196,N_17902);
nor U19937 (N_19937,N_16700,N_17965);
and U19938 (N_19938,N_16059,N_16229);
xor U19939 (N_19939,N_16999,N_16271);
nor U19940 (N_19940,N_16042,N_17364);
or U19941 (N_19941,N_17344,N_17185);
nor U19942 (N_19942,N_16732,N_17138);
or U19943 (N_19943,N_17416,N_17973);
nor U19944 (N_19944,N_17258,N_17948);
and U19945 (N_19945,N_17685,N_16641);
or U19946 (N_19946,N_17938,N_16814);
nor U19947 (N_19947,N_17883,N_17785);
nand U19948 (N_19948,N_16307,N_17795);
and U19949 (N_19949,N_16145,N_17154);
nand U19950 (N_19950,N_17121,N_17518);
and U19951 (N_19951,N_17471,N_17968);
or U19952 (N_19952,N_17395,N_16624);
or U19953 (N_19953,N_17904,N_17634);
and U19954 (N_19954,N_17296,N_17093);
or U19955 (N_19955,N_16331,N_17797);
nor U19956 (N_19956,N_17883,N_17105);
and U19957 (N_19957,N_17737,N_17346);
nor U19958 (N_19958,N_16697,N_17828);
xor U19959 (N_19959,N_17390,N_17936);
nand U19960 (N_19960,N_17836,N_16994);
or U19961 (N_19961,N_16880,N_17953);
and U19962 (N_19962,N_16420,N_17140);
or U19963 (N_19963,N_16077,N_16484);
or U19964 (N_19964,N_16689,N_16485);
xor U19965 (N_19965,N_17502,N_17395);
nor U19966 (N_19966,N_17876,N_17525);
nor U19967 (N_19967,N_17455,N_17581);
nor U19968 (N_19968,N_16808,N_16568);
nor U19969 (N_19969,N_17234,N_17038);
nor U19970 (N_19970,N_16050,N_16812);
nor U19971 (N_19971,N_17068,N_17462);
nand U19972 (N_19972,N_17043,N_17677);
nand U19973 (N_19973,N_16606,N_17380);
and U19974 (N_19974,N_16939,N_17253);
nor U19975 (N_19975,N_17771,N_16963);
and U19976 (N_19976,N_16400,N_16226);
and U19977 (N_19977,N_17809,N_17721);
or U19978 (N_19978,N_16652,N_16478);
nand U19979 (N_19979,N_16874,N_17929);
nand U19980 (N_19980,N_17566,N_17666);
or U19981 (N_19981,N_16642,N_17641);
nor U19982 (N_19982,N_16985,N_17551);
nand U19983 (N_19983,N_16069,N_16046);
nor U19984 (N_19984,N_16209,N_17214);
xor U19985 (N_19985,N_16989,N_16770);
nor U19986 (N_19986,N_16654,N_17711);
xnor U19987 (N_19987,N_17302,N_17914);
or U19988 (N_19988,N_17376,N_16014);
or U19989 (N_19989,N_16463,N_16269);
nand U19990 (N_19990,N_16637,N_16970);
nand U19991 (N_19991,N_17961,N_17515);
or U19992 (N_19992,N_17084,N_16062);
nand U19993 (N_19993,N_16807,N_17964);
and U19994 (N_19994,N_17308,N_17609);
nand U19995 (N_19995,N_16049,N_16871);
nor U19996 (N_19996,N_17305,N_17945);
and U19997 (N_19997,N_17120,N_16485);
and U19998 (N_19998,N_16705,N_16436);
nand U19999 (N_19999,N_17103,N_16294);
nand UO_0 (O_0,N_18409,N_19100);
and UO_1 (O_1,N_19920,N_18349);
nand UO_2 (O_2,N_18187,N_19241);
and UO_3 (O_3,N_19779,N_19116);
or UO_4 (O_4,N_18656,N_19832);
nand UO_5 (O_5,N_18356,N_18703);
or UO_6 (O_6,N_18478,N_19618);
nand UO_7 (O_7,N_18692,N_18856);
or UO_8 (O_8,N_18093,N_19112);
nor UO_9 (O_9,N_18902,N_19184);
or UO_10 (O_10,N_18393,N_18251);
and UO_11 (O_11,N_19483,N_19398);
nand UO_12 (O_12,N_18921,N_19118);
or UO_13 (O_13,N_19639,N_19982);
nor UO_14 (O_14,N_19895,N_19185);
or UO_15 (O_15,N_19713,N_18009);
nor UO_16 (O_16,N_18842,N_19870);
or UO_17 (O_17,N_19901,N_19438);
xnor UO_18 (O_18,N_18639,N_18386);
nor UO_19 (O_19,N_18653,N_18406);
and UO_20 (O_20,N_18905,N_18184);
and UO_21 (O_21,N_18941,N_18029);
nor UO_22 (O_22,N_18199,N_19226);
and UO_23 (O_23,N_19166,N_18257);
nand UO_24 (O_24,N_18831,N_19355);
and UO_25 (O_25,N_19427,N_18577);
or UO_26 (O_26,N_19509,N_18723);
or UO_27 (O_27,N_18796,N_19972);
nand UO_28 (O_28,N_19403,N_19143);
and UO_29 (O_29,N_18085,N_19371);
nor UO_30 (O_30,N_19480,N_19090);
or UO_31 (O_31,N_19531,N_18550);
and UO_32 (O_32,N_19145,N_18351);
nand UO_33 (O_33,N_18272,N_19188);
nand UO_34 (O_34,N_19511,N_18479);
and UO_35 (O_35,N_18321,N_18866);
nand UO_36 (O_36,N_19921,N_18519);
or UO_37 (O_37,N_19503,N_19573);
nand UO_38 (O_38,N_19123,N_18245);
nand UO_39 (O_39,N_18769,N_18338);
and UO_40 (O_40,N_18400,N_18361);
nand UO_41 (O_41,N_18541,N_19668);
or UO_42 (O_42,N_19054,N_19887);
and UO_43 (O_43,N_18574,N_19691);
or UO_44 (O_44,N_18496,N_19368);
nor UO_45 (O_45,N_18868,N_19286);
nor UO_46 (O_46,N_19714,N_19893);
nand UO_47 (O_47,N_18489,N_19673);
and UO_48 (O_48,N_18504,N_18256);
nor UO_49 (O_49,N_18837,N_18976);
nor UO_50 (O_50,N_18357,N_19918);
or UO_51 (O_51,N_18940,N_18620);
or UO_52 (O_52,N_18657,N_18105);
or UO_53 (O_53,N_19314,N_19194);
nand UO_54 (O_54,N_19572,N_18755);
and UO_55 (O_55,N_19758,N_19720);
and UO_56 (O_56,N_18147,N_18697);
or UO_57 (O_57,N_19363,N_18185);
and UO_58 (O_58,N_19099,N_18224);
and UO_59 (O_59,N_19277,N_19923);
nand UO_60 (O_60,N_19603,N_19381);
or UO_61 (O_61,N_19827,N_18596);
or UO_62 (O_62,N_19141,N_19338);
or UO_63 (O_63,N_19683,N_18861);
nor UO_64 (O_64,N_18964,N_18287);
and UO_65 (O_65,N_19191,N_19174);
nor UO_66 (O_66,N_18246,N_19187);
or UO_67 (O_67,N_18672,N_18008);
or UO_68 (O_68,N_18883,N_19745);
xor UO_69 (O_69,N_19393,N_19125);
nor UO_70 (O_70,N_18456,N_18983);
and UO_71 (O_71,N_18616,N_18141);
or UO_72 (O_72,N_19769,N_18906);
and UO_73 (O_73,N_19919,N_18150);
or UO_74 (O_74,N_19809,N_19965);
or UO_75 (O_75,N_18714,N_18016);
nand UO_76 (O_76,N_19852,N_19929);
nand UO_77 (O_77,N_19791,N_18525);
and UO_78 (O_78,N_19937,N_19073);
and UO_79 (O_79,N_19866,N_19439);
xnor UO_80 (O_80,N_19130,N_19315);
and UO_81 (O_81,N_19131,N_19305);
nor UO_82 (O_82,N_18407,N_18365);
nand UO_83 (O_83,N_18335,N_19971);
and UO_84 (O_84,N_19447,N_18359);
or UO_85 (O_85,N_19012,N_18779);
or UO_86 (O_86,N_18043,N_19914);
nand UO_87 (O_87,N_18273,N_18982);
nor UO_88 (O_88,N_19493,N_18067);
nand UO_89 (O_89,N_19991,N_18355);
nor UO_90 (O_90,N_19756,N_19881);
xor UO_91 (O_91,N_19179,N_18670);
and UO_92 (O_92,N_19999,N_19486);
nand UO_93 (O_93,N_18939,N_19794);
xor UO_94 (O_94,N_19815,N_18735);
or UO_95 (O_95,N_18413,N_19193);
and UO_96 (O_96,N_18924,N_19489);
or UO_97 (O_97,N_18563,N_18743);
or UO_98 (O_98,N_18621,N_18996);
nor UO_99 (O_99,N_19181,N_19140);
and UO_100 (O_100,N_19906,N_18152);
nor UO_101 (O_101,N_19024,N_19276);
nand UO_102 (O_102,N_18310,N_18468);
nor UO_103 (O_103,N_18353,N_19458);
nor UO_104 (O_104,N_19859,N_18640);
nor UO_105 (O_105,N_19380,N_18193);
nand UO_106 (O_106,N_19886,N_18311);
or UO_107 (O_107,N_19762,N_19421);
nand UO_108 (O_108,N_19496,N_19149);
nand UO_109 (O_109,N_19821,N_18198);
nand UO_110 (O_110,N_19299,N_18342);
xnor UO_111 (O_111,N_18581,N_19308);
and UO_112 (O_112,N_19195,N_19165);
xor UO_113 (O_113,N_19258,N_18678);
or UO_114 (O_114,N_18696,N_19292);
or UO_115 (O_115,N_19443,N_18995);
nor UO_116 (O_116,N_18783,N_19153);
nand UO_117 (O_117,N_18225,N_19065);
nor UO_118 (O_118,N_19126,N_18605);
nand UO_119 (O_119,N_18918,N_18677);
and UO_120 (O_120,N_18417,N_19243);
nand UO_121 (O_121,N_19250,N_18891);
or UO_122 (O_122,N_19412,N_19750);
or UO_123 (O_123,N_18260,N_19932);
or UO_124 (O_124,N_19863,N_18740);
and UO_125 (O_125,N_18113,N_19465);
and UO_126 (O_126,N_19442,N_18623);
nand UO_127 (O_127,N_18717,N_19260);
nor UO_128 (O_128,N_18004,N_19210);
nor UO_129 (O_129,N_18431,N_18899);
nor UO_130 (O_130,N_18334,N_19346);
or UO_131 (O_131,N_18092,N_18764);
nor UO_132 (O_132,N_18711,N_18233);
xnor UO_133 (O_133,N_18477,N_18022);
nor UO_134 (O_134,N_19528,N_18585);
xnor UO_135 (O_135,N_18052,N_19601);
and UO_136 (O_136,N_19504,N_19175);
nand UO_137 (O_137,N_18002,N_19296);
or UO_138 (O_138,N_18425,N_19900);
nor UO_139 (O_139,N_18214,N_18427);
and UO_140 (O_140,N_19695,N_18915);
and UO_141 (O_141,N_18784,N_18049);
nand UO_142 (O_142,N_18348,N_18627);
and UO_143 (O_143,N_18299,N_19341);
or UO_144 (O_144,N_19703,N_19494);
and UO_145 (O_145,N_19606,N_19553);
nand UO_146 (O_146,N_18102,N_19506);
nor UO_147 (O_147,N_19671,N_18054);
xnor UO_148 (O_148,N_18155,N_19744);
xor UO_149 (O_149,N_19018,N_19416);
xor UO_150 (O_150,N_19613,N_18283);
or UO_151 (O_151,N_19177,N_18363);
nand UO_152 (O_152,N_18001,N_19422);
nand UO_153 (O_153,N_18775,N_18968);
nand UO_154 (O_154,N_19843,N_18178);
nand UO_155 (O_155,N_19765,N_19037);
or UO_156 (O_156,N_19641,N_18591);
nand UO_157 (O_157,N_18989,N_19556);
xnor UO_158 (O_158,N_19324,N_19415);
or UO_159 (O_159,N_19088,N_19868);
nor UO_160 (O_160,N_19616,N_19811);
xor UO_161 (O_161,N_18572,N_19955);
nand UO_162 (O_162,N_19708,N_19963);
and UO_163 (O_163,N_18452,N_19202);
nand UO_164 (O_164,N_18443,N_18462);
or UO_165 (O_165,N_19958,N_19013);
and UO_166 (O_166,N_19792,N_19726);
and UO_167 (O_167,N_18028,N_19059);
nand UO_168 (O_168,N_19807,N_18803);
and UO_169 (O_169,N_19294,N_19537);
or UO_170 (O_170,N_19559,N_19709);
and UO_171 (O_171,N_19017,N_19462);
nor UO_172 (O_172,N_18930,N_19798);
nand UO_173 (O_173,N_18588,N_18383);
and UO_174 (O_174,N_19425,N_19535);
nor UO_175 (O_175,N_18457,N_19461);
and UO_176 (O_176,N_18104,N_19977);
nand UO_177 (O_177,N_18998,N_19530);
nor UO_178 (O_178,N_19956,N_18833);
nor UO_179 (O_179,N_18910,N_18380);
or UO_180 (O_180,N_19446,N_19234);
xor UO_181 (O_181,N_19280,N_18534);
nor UO_182 (O_182,N_19678,N_19730);
or UO_183 (O_183,N_19636,N_18699);
nand UO_184 (O_184,N_19681,N_18858);
and UO_185 (O_185,N_18328,N_18231);
nand UO_186 (O_186,N_19625,N_18725);
and UO_187 (O_187,N_19101,N_18416);
xor UO_188 (O_188,N_18652,N_19563);
nor UO_189 (O_189,N_18241,N_18644);
nand UO_190 (O_190,N_19888,N_18451);
nor UO_191 (O_191,N_18073,N_18538);
and UO_192 (O_192,N_19097,N_18206);
and UO_193 (O_193,N_19871,N_19034);
and UO_194 (O_194,N_19208,N_19395);
nor UO_195 (O_195,N_19105,N_18798);
and UO_196 (O_196,N_19436,N_18838);
nor UO_197 (O_197,N_18539,N_18279);
xnor UO_198 (O_198,N_18481,N_19926);
and UO_199 (O_199,N_18999,N_18994);
nor UO_200 (O_200,N_19328,N_18947);
nand UO_201 (O_201,N_19160,N_19575);
or UO_202 (O_202,N_18292,N_18872);
and UO_203 (O_203,N_18773,N_18163);
or UO_204 (O_204,N_18038,N_19817);
nor UO_205 (O_205,N_19941,N_19089);
xor UO_206 (O_206,N_18601,N_18209);
and UO_207 (O_207,N_18254,N_19658);
nand UO_208 (O_208,N_19505,N_18592);
nor UO_209 (O_209,N_18165,N_19759);
nor UO_210 (O_210,N_18249,N_19220);
and UO_211 (O_211,N_18841,N_18221);
or UO_212 (O_212,N_19297,N_18689);
xnor UO_213 (O_213,N_18923,N_19468);
nor UO_214 (O_214,N_19864,N_19833);
nor UO_215 (O_215,N_19084,N_18414);
nor UO_216 (O_216,N_18810,N_18455);
xnor UO_217 (O_217,N_19384,N_19330);
and UO_218 (O_218,N_19488,N_19157);
nand UO_219 (O_219,N_19596,N_19580);
and UO_220 (O_220,N_18378,N_19567);
nor UO_221 (O_221,N_18985,N_18244);
nor UO_222 (O_222,N_18569,N_19312);
nand UO_223 (O_223,N_18617,N_18793);
nand UO_224 (O_224,N_18785,N_19102);
nand UO_225 (O_225,N_18761,N_18865);
nand UO_226 (O_226,N_19770,N_19410);
and UO_227 (O_227,N_19904,N_18878);
nand UO_228 (O_228,N_19644,N_18552);
xnor UO_229 (O_229,N_19359,N_19289);
nor UO_230 (O_230,N_19444,N_19058);
or UO_231 (O_231,N_19552,N_18745);
xor UO_232 (O_232,N_19109,N_19336);
or UO_233 (O_233,N_18682,N_18951);
or UO_234 (O_234,N_18240,N_19554);
nor UO_235 (O_235,N_19266,N_19699);
nand UO_236 (O_236,N_18958,N_18847);
nor UO_237 (O_237,N_19343,N_19285);
nor UO_238 (O_238,N_19772,N_19066);
and UO_239 (O_239,N_19722,N_19541);
nor UO_240 (O_240,N_18136,N_18753);
nor UO_241 (O_241,N_19516,N_19566);
nand UO_242 (O_242,N_18450,N_18173);
nor UO_243 (O_243,N_18718,N_18511);
or UO_244 (O_244,N_19902,N_19803);
nor UO_245 (O_245,N_18562,N_19263);
nor UO_246 (O_246,N_19753,N_18396);
nor UO_247 (O_247,N_19818,N_19041);
nand UO_248 (O_248,N_19682,N_18291);
and UO_249 (O_249,N_19274,N_18367);
nor UO_250 (O_250,N_18587,N_18015);
nor UO_251 (O_251,N_19916,N_18687);
xnor UO_252 (O_252,N_19764,N_18854);
or UO_253 (O_253,N_19874,N_19860);
or UO_254 (O_254,N_18663,N_19647);
xnor UO_255 (O_255,N_18467,N_18827);
and UO_256 (O_256,N_19850,N_18791);
nor UO_257 (O_257,N_18084,N_19056);
nand UO_258 (O_258,N_19590,N_19426);
nand UO_259 (O_259,N_18343,N_18253);
and UO_260 (O_260,N_19255,N_18024);
nor UO_261 (O_261,N_19627,N_18154);
nand UO_262 (O_262,N_18044,N_18758);
and UO_263 (O_263,N_19046,N_19044);
and UO_264 (O_264,N_19954,N_18545);
nor UO_265 (O_265,N_19478,N_19751);
and UO_266 (O_266,N_19755,N_18633);
and UO_267 (O_267,N_19674,N_18727);
nand UO_268 (O_268,N_19135,N_18146);
or UO_269 (O_269,N_18134,N_18611);
and UO_270 (O_270,N_19348,N_19071);
nand UO_271 (O_271,N_19477,N_19749);
xor UO_272 (O_272,N_18603,N_18835);
nor UO_273 (O_273,N_19408,N_19754);
nand UO_274 (O_274,N_19216,N_18629);
nor UO_275 (O_275,N_18341,N_18072);
or UO_276 (O_276,N_19829,N_19848);
nor UO_277 (O_277,N_19677,N_18634);
or UO_278 (O_278,N_19669,N_19108);
and UO_279 (O_279,N_19917,N_18109);
or UO_280 (O_280,N_19282,N_18327);
nor UO_281 (O_281,N_19544,N_18509);
or UO_282 (O_282,N_18884,N_19998);
nor UO_283 (O_283,N_19911,N_18867);
nor UO_284 (O_284,N_19020,N_18943);
nand UO_285 (O_285,N_18886,N_18993);
and UO_286 (O_286,N_19182,N_18120);
or UO_287 (O_287,N_19391,N_19409);
and UO_288 (O_288,N_19599,N_19736);
nand UO_289 (O_289,N_18060,N_19492);
and UO_290 (O_290,N_19600,N_19577);
and UO_291 (O_291,N_18688,N_18161);
xor UO_292 (O_292,N_18003,N_19473);
or UO_293 (O_293,N_18041,N_19161);
nor UO_294 (O_294,N_19679,N_18205);
and UO_295 (O_295,N_18919,N_18110);
nand UO_296 (O_296,N_19718,N_19912);
nor UO_297 (O_297,N_18473,N_19984);
nor UO_298 (O_298,N_19604,N_19705);
nand UO_299 (O_299,N_18051,N_18805);
or UO_300 (O_300,N_19783,N_18143);
nor UO_301 (O_301,N_18516,N_19448);
nor UO_302 (O_302,N_18666,N_18690);
or UO_303 (O_303,N_19248,N_19872);
nor UO_304 (O_304,N_18180,N_19347);
nand UO_305 (O_305,N_18502,N_18490);
nand UO_306 (O_306,N_19659,N_19378);
or UO_307 (O_307,N_19694,N_19428);
xor UO_308 (O_308,N_19091,N_18329);
nand UO_309 (O_309,N_18613,N_19574);
or UO_310 (O_310,N_18219,N_18920);
nand UO_311 (O_311,N_18290,N_18771);
and UO_312 (O_312,N_19351,N_19434);
nand UO_313 (O_313,N_18200,N_19386);
xor UO_314 (O_314,N_19275,N_18780);
nand UO_315 (O_315,N_18293,N_18966);
xor UO_316 (O_316,N_18956,N_18862);
or UO_317 (O_317,N_19164,N_18654);
xnor UO_318 (O_318,N_18503,N_18333);
nand UO_319 (O_319,N_18124,N_18598);
and UO_320 (O_320,N_18397,N_19651);
xor UO_321 (O_321,N_18521,N_19790);
nand UO_322 (O_322,N_19392,N_18307);
xnor UO_323 (O_323,N_18377,N_19610);
nor UO_324 (O_324,N_18536,N_19159);
nand UO_325 (O_325,N_19529,N_18974);
or UO_326 (O_326,N_19256,N_19212);
nand UO_327 (O_327,N_19799,N_19055);
nor UO_328 (O_328,N_18911,N_18314);
xnor UO_329 (O_329,N_19631,N_19376);
nor UO_330 (O_330,N_18801,N_19952);
nor UO_331 (O_331,N_18484,N_18626);
nand UO_332 (O_332,N_18444,N_19455);
or UO_333 (O_333,N_18843,N_18277);
or UO_334 (O_334,N_19546,N_18454);
or UO_335 (O_335,N_19092,N_18298);
nand UO_336 (O_336,N_19332,N_19086);
xnor UO_337 (O_337,N_19686,N_18375);
nor UO_338 (O_338,N_19288,N_19215);
nand UO_339 (O_339,N_18800,N_18816);
nand UO_340 (O_340,N_19967,N_18535);
nor UO_341 (O_341,N_19011,N_19615);
nor UO_342 (O_342,N_18701,N_19609);
and UO_343 (O_343,N_18848,N_18881);
or UO_344 (O_344,N_19508,N_18284);
xnor UO_345 (O_345,N_19278,N_18326);
and UO_346 (O_346,N_19252,N_18845);
and UO_347 (O_347,N_18495,N_19890);
and UO_348 (O_348,N_19320,N_18529);
nand UO_349 (O_349,N_19879,N_18709);
nor UO_350 (O_350,N_19085,N_19045);
and UO_351 (O_351,N_19635,N_19737);
or UO_352 (O_352,N_19549,N_18869);
nand UO_353 (O_353,N_19449,N_19626);
or UO_354 (O_354,N_18089,N_19362);
nor UO_355 (O_355,N_18568,N_19767);
or UO_356 (O_356,N_19329,N_19497);
or UO_357 (O_357,N_19935,N_19318);
or UO_358 (O_358,N_19562,N_19259);
xnor UO_359 (O_359,N_18339,N_18695);
nand UO_360 (O_360,N_19908,N_19325);
or UO_361 (O_361,N_19245,N_18961);
or UO_362 (O_362,N_19656,N_19978);
or UO_363 (O_363,N_19349,N_19632);
nand UO_364 (O_364,N_19374,N_18056);
or UO_365 (O_365,N_18373,N_19525);
or UO_366 (O_366,N_18969,N_19070);
nand UO_367 (O_367,N_19761,N_19238);
nand UO_368 (O_368,N_19230,N_18247);
or UO_369 (O_369,N_19898,N_19962);
nor UO_370 (O_370,N_19120,N_19290);
xnor UO_371 (O_371,N_19560,N_18074);
and UO_372 (O_372,N_18218,N_19028);
nand UO_373 (O_373,N_19533,N_18151);
or UO_374 (O_374,N_19479,N_18057);
or UO_375 (O_375,N_19413,N_18760);
and UO_376 (O_376,N_19614,N_18168);
or UO_377 (O_377,N_18220,N_19854);
or UO_378 (O_378,N_18645,N_19158);
and UO_379 (O_379,N_19352,N_19608);
and UO_380 (O_380,N_19653,N_19253);
and UO_381 (O_381,N_19162,N_19624);
or UO_382 (O_382,N_19979,N_18012);
and UO_383 (O_383,N_18300,N_18265);
and UO_384 (O_384,N_18636,N_19242);
or UO_385 (O_385,N_19420,N_18719);
nand UO_386 (O_386,N_19106,N_18759);
nand UO_387 (O_387,N_18935,N_19842);
nand UO_388 (O_388,N_19789,N_18561);
or UO_389 (O_389,N_19137,N_19414);
and UO_390 (O_390,N_19729,N_19339);
and UO_391 (O_391,N_19321,N_19734);
and UO_392 (O_392,N_18033,N_18418);
nor UO_393 (O_393,N_19096,N_19377);
or UO_394 (O_394,N_19005,N_19081);
nand UO_395 (O_395,N_18059,N_19640);
nor UO_396 (O_396,N_18807,N_19180);
nand UO_397 (O_397,N_18385,N_19570);
or UO_398 (O_398,N_19500,N_18594);
nor UO_399 (O_399,N_18737,N_18700);
nand UO_400 (O_400,N_19460,N_19057);
or UO_401 (O_401,N_19262,N_19113);
and UO_402 (O_402,N_18021,N_19155);
and UO_403 (O_403,N_19747,N_19814);
or UO_404 (O_404,N_19370,N_19974);
nor UO_405 (O_405,N_18019,N_19822);
nor UO_406 (O_406,N_18544,N_18691);
nand UO_407 (O_407,N_19796,N_18806);
xor UO_408 (O_408,N_18441,N_19132);
nor UO_409 (O_409,N_19246,N_18622);
and UO_410 (O_410,N_19670,N_19899);
and UO_411 (O_411,N_19813,N_18174);
and UO_412 (O_412,N_18204,N_18990);
nand UO_413 (O_413,N_19203,N_18181);
and UO_414 (O_414,N_19265,N_18111);
and UO_415 (O_415,N_18664,N_19358);
xnor UO_416 (O_416,N_18904,N_18515);
and UO_417 (O_417,N_18023,N_18227);
nand UO_418 (O_418,N_19828,N_19042);
nor UO_419 (O_419,N_19643,N_18903);
xnor UO_420 (O_420,N_18319,N_18037);
nand UO_421 (O_421,N_18765,N_19176);
and UO_422 (O_422,N_19660,N_19353);
nor UO_423 (O_423,N_19302,N_19701);
nor UO_424 (O_424,N_19568,N_19107);
nand UO_425 (O_425,N_18389,N_19450);
nor UO_426 (O_426,N_18813,N_18142);
or UO_427 (O_427,N_19602,N_18288);
nand UO_428 (O_428,N_19786,N_19236);
nand UO_429 (O_429,N_19069,N_19649);
or UO_430 (O_430,N_18324,N_19521);
nand UO_431 (O_431,N_18928,N_18453);
nand UO_432 (O_432,N_18762,N_18354);
nor UO_433 (O_433,N_19068,N_19960);
nand UO_434 (O_434,N_18039,N_19440);
or UO_435 (O_435,N_19016,N_19867);
or UO_436 (O_436,N_18295,N_19030);
nand UO_437 (O_437,N_18510,N_19032);
nor UO_438 (O_438,N_18907,N_18967);
or UO_439 (O_439,N_19469,N_19524);
or UO_440 (O_440,N_18997,N_19249);
and UO_441 (O_441,N_18212,N_18498);
and UO_442 (O_442,N_18533,N_18712);
nor UO_443 (O_443,N_18826,N_18487);
and UO_444 (O_444,N_19372,N_18020);
and UO_445 (O_445,N_19988,N_19424);
nand UO_446 (O_446,N_19061,N_18589);
nand UO_447 (O_447,N_18683,N_18062);
and UO_448 (O_448,N_19051,N_18635);
and UO_449 (O_449,N_18608,N_18446);
and UO_450 (O_450,N_18422,N_18088);
and UO_451 (O_451,N_18061,N_18957);
nor UO_452 (O_452,N_19950,N_19648);
or UO_453 (O_453,N_18223,N_18946);
xnor UO_454 (O_454,N_19499,N_19795);
or UO_455 (O_455,N_18305,N_18557);
or UO_456 (O_456,N_18937,N_18264);
or UO_457 (O_457,N_18252,N_18971);
nor UO_458 (O_458,N_18156,N_18882);
and UO_459 (O_459,N_19279,N_19877);
or UO_460 (O_460,N_18170,N_19802);
nor UO_461 (O_461,N_18391,N_18981);
or UO_462 (O_462,N_18469,N_19036);
xnor UO_463 (O_463,N_18875,N_19291);
nor UO_464 (O_464,N_18197,N_18660);
or UO_465 (O_465,N_19716,N_19665);
nor UO_466 (O_466,N_18790,N_19797);
nand UO_467 (O_467,N_19053,N_18528);
or UO_468 (O_468,N_19589,N_19283);
nor UO_469 (O_469,N_19951,N_19490);
or UO_470 (O_470,N_18650,N_19110);
xnor UO_471 (O_471,N_18984,N_18302);
nand UO_472 (O_472,N_19543,N_19839);
and UO_473 (O_473,N_18119,N_18694);
nor UO_474 (O_474,N_18280,N_19227);
and UO_475 (O_475,N_19471,N_19264);
or UO_476 (O_476,N_18722,N_18583);
and UO_477 (O_477,N_18226,N_18638);
xnor UO_478 (O_478,N_19419,N_19049);
nand UO_479 (O_479,N_18186,N_18742);
and UO_480 (O_480,N_18235,N_18420);
or UO_481 (O_481,N_18724,N_18447);
or UO_482 (O_482,N_18301,N_18017);
nand UO_483 (O_483,N_18079,N_18007);
xnor UO_484 (O_484,N_18025,N_18507);
or UO_485 (O_485,N_19183,N_18107);
nor UO_486 (O_486,N_19928,N_19732);
and UO_487 (O_487,N_18669,N_18318);
xor UO_488 (O_488,N_19808,N_18175);
or UO_489 (O_489,N_19768,N_18169);
or UO_490 (O_490,N_18744,N_19031);
xor UO_491 (O_491,N_18782,N_19922);
and UO_492 (O_492,N_19882,N_19388);
nand UO_493 (O_493,N_18849,N_18262);
or UO_494 (O_494,N_19949,N_18123);
or UO_495 (O_495,N_18485,N_18309);
and UO_496 (O_496,N_18286,N_19401);
or UO_497 (O_497,N_19819,N_18065);
nand UO_498 (O_498,N_19062,N_19327);
or UO_499 (O_499,N_19621,N_19316);
or UO_500 (O_500,N_18524,N_18948);
nand UO_501 (O_501,N_19214,N_19548);
nand UO_502 (O_502,N_19878,N_18148);
and UO_503 (O_503,N_19129,N_18208);
nand UO_504 (O_504,N_19856,N_19526);
nand UO_505 (O_505,N_18387,N_18242);
nor UO_506 (O_506,N_19119,N_19078);
nor UO_507 (O_507,N_18844,N_18532);
nor UO_508 (O_508,N_18312,N_18392);
or UO_509 (O_509,N_19633,N_18177);
nand UO_510 (O_510,N_18739,N_19379);
nor UO_511 (O_511,N_19752,N_18618);
and UO_512 (O_512,N_18461,N_18986);
nand UO_513 (O_513,N_18604,N_18708);
nand UO_514 (O_514,N_18750,N_18809);
and UO_515 (O_515,N_18424,N_19945);
xor UO_516 (O_516,N_19522,N_19170);
xor UO_517 (O_517,N_18316,N_18846);
nand UO_518 (O_518,N_19136,N_18560);
nand UO_519 (O_519,N_18860,N_18916);
nand UO_520 (O_520,N_18522,N_19739);
nor UO_521 (O_521,N_18306,N_19953);
or UO_522 (O_522,N_19557,N_19717);
nand UO_523 (O_523,N_18929,N_18121);
nor UO_524 (O_524,N_18135,N_19778);
nor UO_525 (O_525,N_19947,N_18571);
nor UO_526 (O_526,N_18384,N_18978);
and UO_527 (O_527,N_19777,N_19261);
xor UO_528 (O_528,N_18442,N_18767);
and UO_529 (O_529,N_19457,N_19800);
xor UO_530 (O_530,N_19989,N_19835);
and UO_531 (O_531,N_19710,N_18836);
and UO_532 (O_532,N_19801,N_19139);
xnor UO_533 (O_533,N_18258,N_18050);
xnor UO_534 (O_534,N_18144,N_19072);
and UO_535 (O_535,N_19698,N_19047);
or UO_536 (O_536,N_19689,N_19780);
nand UO_537 (O_537,N_19178,N_19225);
and UO_538 (O_538,N_19536,N_18628);
or UO_539 (O_539,N_19389,N_18125);
or UO_540 (O_540,N_18819,N_19731);
xor UO_541 (O_541,N_19233,N_19650);
and UO_542 (O_542,N_18248,N_18543);
or UO_543 (O_543,N_19437,N_18269);
and UO_544 (O_544,N_19663,N_19957);
or UO_545 (O_545,N_19931,N_19402);
or UO_546 (O_546,N_18526,N_18987);
xnor UO_547 (O_547,N_19117,N_18063);
or UO_548 (O_548,N_18681,N_19510);
nor UO_549 (O_549,N_18030,N_18756);
nor UO_550 (O_550,N_18595,N_18201);
nor UO_551 (O_551,N_18331,N_19350);
nor UO_552 (O_552,N_19093,N_19696);
nand UO_553 (O_553,N_18068,N_19333);
or UO_554 (O_554,N_19103,N_19806);
and UO_555 (O_555,N_18388,N_18897);
nand UO_556 (O_556,N_18194,N_18282);
and UO_557 (O_557,N_18963,N_19517);
nand UO_558 (O_558,N_19094,N_18207);
nor UO_559 (O_559,N_18275,N_19128);
and UO_560 (O_560,N_19724,N_19823);
or UO_561 (O_561,N_19907,N_18901);
nor UO_562 (O_562,N_19983,N_18076);
nor UO_563 (O_563,N_19002,N_19812);
nand UO_564 (O_564,N_19834,N_18347);
or UO_565 (O_565,N_18702,N_19990);
nor UO_566 (O_566,N_19326,N_19685);
and UO_567 (O_567,N_18716,N_19513);
and UO_568 (O_568,N_19507,N_19198);
nand UO_569 (O_569,N_18099,N_19142);
xor UO_570 (O_570,N_19172,N_18979);
nor UO_571 (O_571,N_18763,N_19862);
or UO_572 (O_572,N_18166,N_19331);
xnor UO_573 (O_573,N_18894,N_19592);
and UO_574 (O_574,N_19079,N_18895);
nand UO_575 (O_575,N_18297,N_18081);
nor UO_576 (O_576,N_19688,N_18733);
nor UO_577 (O_577,N_18953,N_18419);
xor UO_578 (O_578,N_18736,N_19788);
or UO_579 (O_579,N_18632,N_18766);
or UO_580 (O_580,N_18237,N_18641);
xor UO_581 (O_581,N_18922,N_19518);
and UO_582 (O_582,N_19022,N_18671);
nor UO_583 (O_583,N_18364,N_18781);
nor UO_584 (O_584,N_18285,N_18705);
xor UO_585 (O_585,N_18483,N_19441);
nor UO_586 (O_586,N_19869,N_19087);
nor UO_587 (O_587,N_19387,N_18133);
or UO_588 (O_588,N_18176,N_19781);
nand UO_589 (O_589,N_18236,N_19453);
nor UO_590 (O_590,N_18778,N_18491);
and UO_591 (O_591,N_18980,N_19317);
and UO_592 (O_592,N_19154,N_19199);
xnor UO_593 (O_593,N_19223,N_18655);
and UO_594 (O_594,N_19186,N_19723);
nand UO_595 (O_595,N_19976,N_18615);
nor UO_596 (O_596,N_18474,N_18789);
and UO_597 (O_597,N_19050,N_18751);
nor UO_598 (O_598,N_18651,N_19147);
and UO_599 (O_599,N_19970,N_18137);
or UO_600 (O_600,N_19373,N_19735);
or UO_601 (O_601,N_18195,N_18680);
and UO_602 (O_602,N_19251,N_18488);
xor UO_603 (O_603,N_18741,N_19579);
and UO_604 (O_604,N_18614,N_19254);
or UO_605 (O_605,N_18646,N_18497);
nand UO_606 (O_606,N_19021,N_19995);
nand UO_607 (O_607,N_19396,N_18259);
nor UO_608 (O_608,N_19303,N_19542);
or UO_609 (O_609,N_19470,N_18770);
nor UO_610 (O_610,N_19728,N_19630);
nor UO_611 (O_611,N_19122,N_19397);
nor UO_612 (O_612,N_18811,N_18210);
and UO_613 (O_613,N_18013,N_19934);
nor UO_614 (O_614,N_18547,N_19591);
and UO_615 (O_615,N_19993,N_18500);
nor UO_616 (O_616,N_19652,N_18429);
or UO_617 (O_617,N_18590,N_19189);
nor UO_618 (O_618,N_19433,N_18091);
or UO_619 (O_619,N_18693,N_18238);
nand UO_620 (O_620,N_19539,N_18470);
or UO_621 (O_621,N_19611,N_18567);
nand UO_622 (O_622,N_18821,N_19512);
nor UO_623 (O_623,N_19168,N_18877);
or UO_624 (O_624,N_19697,N_18320);
nand UO_625 (O_625,N_19733,N_18047);
or UO_626 (O_626,N_19712,N_18066);
nand UO_627 (O_627,N_18445,N_18374);
nor UO_628 (O_628,N_19925,N_18898);
nand UO_629 (O_629,N_19550,N_19273);
or UO_630 (O_630,N_18202,N_19968);
nand UO_631 (O_631,N_18787,N_18710);
xor UO_632 (O_632,N_18077,N_18619);
and UO_633 (O_633,N_19690,N_18662);
nor UO_634 (O_634,N_18975,N_18126);
or UO_635 (O_635,N_18160,N_18255);
and UO_636 (O_636,N_18370,N_19366);
or UO_637 (O_637,N_18350,N_18513);
nor UO_638 (O_638,N_19946,N_19076);
nand UO_639 (O_639,N_18578,N_19048);
and UO_640 (O_640,N_18399,N_18463);
nor UO_641 (O_641,N_19587,N_19035);
and UO_642 (O_642,N_18768,N_18243);
or UO_643 (O_643,N_18738,N_19304);
nand UO_644 (O_644,N_18885,N_19361);
and UO_645 (O_645,N_19146,N_18992);
and UO_646 (O_646,N_19623,N_19725);
and UO_647 (O_647,N_19672,N_18955);
xor UO_648 (O_648,N_19853,N_19661);
or UO_649 (O_649,N_18234,N_19309);
and UO_650 (O_650,N_18556,N_19948);
nor UO_651 (O_651,N_18433,N_18566);
or UO_652 (O_652,N_19354,N_18874);
nand UO_653 (O_653,N_19200,N_19607);
and UO_654 (O_654,N_19873,N_19295);
xnor UO_655 (O_655,N_18438,N_19742);
nand UO_656 (O_656,N_18428,N_18748);
or UO_657 (O_657,N_19565,N_19404);
and UO_658 (O_658,N_18159,N_19865);
xor UO_659 (O_659,N_18851,N_19231);
or UO_660 (O_660,N_18130,N_19619);
or UO_661 (O_661,N_18600,N_19896);
xnor UO_662 (O_662,N_19484,N_18830);
nand UO_663 (O_663,N_18101,N_18954);
or UO_664 (O_664,N_19287,N_18960);
or UO_665 (O_665,N_18962,N_19365);
nand UO_666 (O_666,N_19040,N_18095);
or UO_667 (O_667,N_19903,N_19400);
nand UO_668 (O_668,N_19959,N_18426);
nor UO_669 (O_669,N_19001,N_19235);
nand UO_670 (O_670,N_18912,N_18965);
nor UO_671 (O_671,N_18482,N_19313);
nand UO_672 (O_672,N_19875,N_19201);
nand UO_673 (O_673,N_18970,N_19004);
and UO_674 (O_674,N_18337,N_18679);
xnor UO_675 (O_675,N_18070,N_19464);
and UO_676 (O_676,N_18676,N_19715);
or UO_677 (O_677,N_18493,N_18075);
nand UO_678 (O_678,N_19007,N_19519);
nor UO_679 (O_679,N_18372,N_19704);
nor UO_680 (O_680,N_18196,N_19693);
and UO_681 (O_681,N_19284,N_18586);
and UO_682 (O_682,N_19239,N_18267);
or UO_683 (O_683,N_18749,N_19540);
or UO_684 (O_684,N_19944,N_19345);
nand UO_685 (O_685,N_18565,N_18673);
or UO_686 (O_686,N_19301,N_18162);
nor UO_687 (O_687,N_18840,N_18322);
or UO_688 (O_688,N_18352,N_19667);
xor UO_689 (O_689,N_19111,N_19482);
nor UO_690 (O_690,N_19064,N_18512);
nand UO_691 (O_691,N_18505,N_18706);
or UO_692 (O_692,N_19646,N_18818);
nand UO_693 (O_693,N_18046,N_19319);
or UO_694 (O_694,N_18116,N_19622);
nor UO_695 (O_695,N_18011,N_18158);
nand UO_696 (O_696,N_18642,N_19655);
nor UO_697 (O_697,N_18410,N_18381);
nor UO_698 (O_698,N_19127,N_19975);
xor UO_699 (O_699,N_19837,N_18517);
nor UO_700 (O_700,N_18839,N_18686);
nor UO_701 (O_701,N_19831,N_18820);
or UO_702 (O_702,N_18643,N_19620);
or UO_703 (O_703,N_19583,N_19675);
nor UO_704 (O_704,N_19052,N_19584);
and UO_705 (O_705,N_19156,N_19171);
or UO_706 (O_706,N_19008,N_18139);
nand UO_707 (O_707,N_19063,N_19545);
and UO_708 (O_708,N_18812,N_18232);
nand UO_709 (O_709,N_18870,N_19067);
or UO_710 (O_710,N_19190,N_19114);
and UO_711 (O_711,N_18434,N_19743);
nor UO_712 (O_712,N_19617,N_18048);
and UO_713 (O_713,N_19344,N_18713);
nor UO_714 (O_714,N_18228,N_19027);
xor UO_715 (O_715,N_19375,N_18358);
nor UO_716 (O_716,N_18157,N_18896);
xor UO_717 (O_717,N_18317,N_19322);
nand UO_718 (O_718,N_18546,N_18344);
xnor UO_719 (O_719,N_19593,N_18908);
nand UO_720 (O_720,N_19082,N_19417);
nand UO_721 (O_721,N_18058,N_18325);
nand UO_722 (O_722,N_19687,N_19151);
nand UO_723 (O_723,N_18944,N_19459);
or UO_724 (O_724,N_19961,N_18988);
or UO_725 (O_725,N_19367,N_19029);
and UO_726 (O_726,N_19083,N_18086);
nor UO_727 (O_727,N_19293,N_19740);
nand UO_728 (O_728,N_19271,N_18728);
nor UO_729 (O_729,N_18625,N_18630);
and UO_730 (O_730,N_18558,N_18936);
or UO_731 (O_731,N_19804,N_19985);
nor UO_732 (O_732,N_18747,N_18876);
nand UO_733 (O_733,N_18599,N_18612);
nand UO_734 (O_734,N_18131,N_19269);
and UO_735 (O_735,N_18403,N_19571);
or UO_736 (O_736,N_18476,N_19173);
or UO_737 (O_737,N_19487,N_19838);
or UO_738 (O_738,N_18730,N_18415);
xor UO_739 (O_739,N_18668,N_18707);
or UO_740 (O_740,N_19664,N_18078);
nor UO_741 (O_741,N_18053,N_18330);
nor UO_742 (O_742,N_19721,N_18859);
nor UO_743 (O_743,N_19826,N_18523);
xor UO_744 (O_744,N_19637,N_18368);
xnor UO_745 (O_745,N_19981,N_18440);
or UO_746 (O_746,N_18430,N_18890);
nor UO_747 (O_747,N_18229,N_18952);
xor UO_748 (O_748,N_19272,N_18777);
or UO_749 (O_749,N_18271,N_19836);
or UO_750 (O_750,N_18950,N_19335);
nand UO_751 (O_751,N_18336,N_18934);
and UO_752 (O_752,N_19406,N_19996);
and UO_753 (O_753,N_19927,N_18786);
or UO_754 (O_754,N_18667,N_19793);
and UO_755 (O_755,N_19910,N_18880);
nor UO_756 (O_756,N_18018,N_19980);
nand UO_757 (O_757,N_18213,N_19485);
and UO_758 (O_758,N_18715,N_19472);
nand UO_759 (O_759,N_18795,N_19657);
xnor UO_760 (O_760,N_19232,N_18499);
nand UO_761 (O_761,N_19431,N_18315);
nand UO_762 (O_762,N_19532,N_18927);
nand UO_763 (O_763,N_19538,N_18360);
nor UO_764 (O_764,N_18405,N_18045);
or UO_765 (O_765,N_18276,N_18822);
nor UO_766 (O_766,N_19432,N_19481);
nor UO_767 (O_767,N_19555,N_19023);
or UO_768 (O_768,N_18190,N_19942);
nand UO_769 (O_769,N_19095,N_19629);
and UO_770 (O_770,N_18752,N_18369);
nor UO_771 (O_771,N_18398,N_19787);
or UO_772 (O_772,N_18069,N_18530);
or UO_773 (O_773,N_19356,N_19986);
nand UO_774 (O_774,N_19551,N_18832);
or UO_775 (O_775,N_18035,N_19323);
nor UO_776 (O_776,N_18597,N_19399);
and UO_777 (O_777,N_18100,N_18346);
nor UO_778 (O_778,N_18892,N_19502);
xor UO_779 (O_779,N_19707,N_19152);
nor UO_780 (O_780,N_18087,N_19987);
xor UO_781 (O_781,N_19605,N_18250);
or UO_782 (O_782,N_19244,N_19534);
and UO_783 (O_783,N_18824,N_19845);
or UO_784 (O_784,N_19892,N_19849);
nand UO_785 (O_785,N_19973,N_18579);
nand UO_786 (O_786,N_19880,N_18893);
and UO_787 (O_787,N_19495,N_18863);
nand UO_788 (O_788,N_18439,N_19340);
xor UO_789 (O_789,N_18720,N_19080);
nor UO_790 (O_790,N_18034,N_19098);
or UO_791 (O_791,N_19766,N_18900);
and UO_792 (O_792,N_18404,N_19855);
and UO_793 (O_793,N_18458,N_19773);
nand UO_794 (O_794,N_18932,N_19169);
nor UO_795 (O_795,N_18850,N_18082);
nor UO_796 (O_796,N_19467,N_19014);
or UO_797 (O_797,N_18432,N_19706);
or UO_798 (O_798,N_18083,N_18659);
or UO_799 (O_799,N_19547,N_19846);
and UO_800 (O_800,N_18266,N_19586);
or UO_801 (O_801,N_18649,N_18217);
nor UO_802 (O_802,N_19825,N_18540);
nor UO_803 (O_803,N_19257,N_18118);
nor UO_804 (O_804,N_19039,N_19454);
nor UO_805 (O_805,N_18575,N_19144);
and UO_806 (O_806,N_18648,N_19390);
nor UO_807 (O_807,N_18323,N_19969);
nand UO_808 (O_808,N_19334,N_18390);
nor UO_809 (O_809,N_18580,N_19905);
xor UO_810 (O_810,N_19847,N_19133);
or UO_811 (O_811,N_19411,N_18857);
nand UO_812 (O_812,N_18506,N_19997);
or UO_813 (O_813,N_18274,N_19430);
nand UO_814 (O_814,N_18829,N_18010);
nor UO_815 (O_815,N_19582,N_18408);
or UO_816 (O_816,N_19206,N_18520);
nand UO_817 (O_817,N_19966,N_19452);
or UO_818 (O_818,N_18115,N_18684);
nand UO_819 (O_819,N_19498,N_18014);
and UO_820 (O_820,N_18027,N_19138);
nor UO_821 (O_821,N_19311,N_19043);
xor UO_822 (O_822,N_18129,N_18402);
nand UO_823 (O_823,N_19771,N_18551);
xnor UO_824 (O_824,N_19684,N_19913);
nand UO_825 (O_825,N_18480,N_18167);
and UO_826 (O_826,N_18239,N_19594);
or UO_827 (O_827,N_19940,N_19891);
and UO_828 (O_828,N_18804,N_18972);
and UO_829 (O_829,N_19435,N_18853);
and UO_830 (O_830,N_18977,N_19025);
nor UO_831 (O_831,N_18071,N_18917);
xor UO_832 (O_832,N_18026,N_19757);
and UO_833 (O_833,N_19746,N_19197);
xnor UO_834 (O_834,N_19357,N_18909);
nor UO_835 (O_835,N_19861,N_18658);
nor UO_836 (O_836,N_19196,N_19385);
xor UO_837 (O_837,N_18914,N_19474);
nand UO_838 (O_838,N_18754,N_19307);
nor UO_839 (O_839,N_19776,N_19298);
or UO_840 (O_840,N_19310,N_18973);
nor UO_841 (O_841,N_19463,N_18814);
nand UO_842 (O_842,N_19213,N_18776);
or UO_843 (O_843,N_18000,N_19578);
or UO_844 (O_844,N_18215,N_19015);
or UO_845 (O_845,N_18726,N_19281);
nand UO_846 (O_846,N_18991,N_19964);
or UO_847 (O_847,N_18179,N_19741);
and UO_848 (O_848,N_18889,N_19711);
nor UO_849 (O_849,N_19115,N_18925);
nor UO_850 (O_850,N_18808,N_18675);
and UO_851 (O_851,N_18542,N_18559);
nor UO_852 (O_852,N_18303,N_19192);
and UO_853 (O_853,N_19700,N_18294);
or UO_854 (O_854,N_19883,N_19909);
nor UO_855 (O_855,N_19595,N_18518);
nor UO_856 (O_856,N_19515,N_18815);
and UO_857 (O_857,N_19719,N_19876);
and UO_858 (O_858,N_19841,N_19000);
nand UO_859 (O_859,N_18624,N_18281);
and UO_860 (O_860,N_19247,N_19840);
xnor UO_861 (O_861,N_19816,N_19211);
and UO_862 (O_862,N_18959,N_19077);
nor UO_863 (O_863,N_19383,N_19810);
and UO_864 (O_864,N_18584,N_18492);
and UO_865 (O_865,N_18537,N_18261);
nor UO_866 (O_866,N_18797,N_18171);
and UO_867 (O_867,N_19581,N_18553);
nand UO_868 (O_868,N_19456,N_18128);
nand UO_869 (O_869,N_19204,N_19588);
and UO_870 (O_870,N_18345,N_19267);
and UO_871 (O_871,N_18421,N_18382);
and UO_872 (O_872,N_18127,N_18465);
and UO_873 (O_873,N_18098,N_19306);
nor UO_874 (O_874,N_18191,N_18040);
or UO_875 (O_875,N_18464,N_18887);
xor UO_876 (O_876,N_19857,N_19824);
nand UO_877 (O_877,N_19523,N_18230);
and UO_878 (O_878,N_19936,N_18411);
xnor UO_879 (O_879,N_18106,N_19337);
nor UO_880 (O_880,N_19520,N_19369);
and UO_881 (O_881,N_19060,N_19405);
and UO_882 (O_882,N_18090,N_19634);
or UO_883 (O_883,N_18731,N_18609);
nand UO_884 (O_884,N_18746,N_19598);
or UO_885 (O_885,N_18734,N_18189);
and UO_886 (O_886,N_19009,N_18460);
and UO_887 (O_887,N_18828,N_18606);
or UO_888 (O_888,N_19775,N_18108);
nor UO_889 (O_889,N_18732,N_19564);
and UO_890 (O_890,N_19897,N_18554);
nand UO_891 (O_891,N_19237,N_18792);
and UO_892 (O_892,N_18103,N_18379);
and UO_893 (O_893,N_19221,N_18549);
nor UO_894 (O_894,N_19666,N_19150);
xnor UO_895 (O_895,N_18032,N_18852);
and UO_896 (O_896,N_19476,N_19830);
xor UO_897 (O_897,N_18931,N_18423);
nand UO_898 (O_898,N_18871,N_18122);
or UO_899 (O_899,N_18448,N_18112);
nand UO_900 (O_900,N_19475,N_18270);
or UO_901 (O_901,N_18698,N_18942);
nand UO_902 (O_902,N_18945,N_18564);
or UO_903 (O_903,N_18602,N_19075);
xor UO_904 (O_904,N_18475,N_19676);
nor UO_905 (O_905,N_19124,N_18055);
nand UO_906 (O_906,N_18278,N_19939);
nand UO_907 (O_907,N_18582,N_19364);
nor UO_908 (O_908,N_19342,N_19167);
and UO_909 (O_909,N_19784,N_18064);
nor UO_910 (O_910,N_19992,N_19763);
nand UO_911 (O_911,N_19418,N_19163);
and UO_912 (O_912,N_18879,N_18501);
xor UO_913 (O_913,N_18437,N_18395);
xor UO_914 (O_914,N_18610,N_18774);
nor UO_915 (O_915,N_19738,N_19654);
nor UO_916 (O_916,N_19003,N_18674);
nor UO_917 (O_917,N_19994,N_19270);
nor UO_918 (O_918,N_18149,N_18607);
nand UO_919 (O_919,N_18412,N_18514);
or UO_920 (O_920,N_18926,N_18799);
nor UO_921 (O_921,N_19205,N_18145);
or UO_922 (O_922,N_19514,N_18313);
or UO_923 (O_923,N_19429,N_19930);
xor UO_924 (O_924,N_18685,N_18555);
nand UO_925 (O_925,N_19774,N_18182);
nand UO_926 (O_926,N_18665,N_19006);
nor UO_927 (O_927,N_18371,N_18114);
nand UO_928 (O_928,N_18304,N_19207);
or UO_929 (O_929,N_18855,N_19889);
nor UO_930 (O_930,N_19360,N_18006);
and UO_931 (O_931,N_18873,N_18459);
and UO_932 (O_932,N_18817,N_19228);
and UO_933 (O_933,N_18183,N_19217);
nand UO_934 (O_934,N_18729,N_19805);
or UO_935 (O_935,N_19680,N_18376);
or UO_936 (O_936,N_18508,N_19885);
or UO_937 (O_937,N_18153,N_19612);
nor UO_938 (O_938,N_18366,N_19558);
nand UO_939 (O_939,N_18794,N_18164);
nand UO_940 (O_940,N_19445,N_19382);
nor UO_941 (O_941,N_19218,N_18527);
nand UO_942 (O_942,N_18531,N_18548);
or UO_943 (O_943,N_18834,N_18938);
and UO_944 (O_944,N_18340,N_18471);
or UO_945 (O_945,N_18825,N_19466);
or UO_946 (O_946,N_18593,N_19209);
nor UO_947 (O_947,N_19074,N_18216);
and UO_948 (O_948,N_19628,N_19423);
nor UO_949 (O_949,N_19943,N_18203);
nand UO_950 (O_950,N_19851,N_18362);
nor UO_951 (O_951,N_19527,N_19148);
nand UO_952 (O_952,N_19576,N_18661);
nand UO_953 (O_953,N_18757,N_18080);
and UO_954 (O_954,N_18211,N_18949);
nand UO_955 (O_955,N_18823,N_19760);
or UO_956 (O_956,N_19748,N_18296);
nand UO_957 (O_957,N_18772,N_18042);
and UO_958 (O_958,N_18576,N_18864);
and UO_959 (O_959,N_18449,N_19019);
nor UO_960 (O_960,N_19645,N_18117);
nand UO_961 (O_961,N_19268,N_19121);
nor UO_962 (O_962,N_19219,N_18435);
nor UO_963 (O_963,N_18472,N_18308);
xor UO_964 (O_964,N_18031,N_18637);
and UO_965 (O_965,N_19844,N_18138);
and UO_966 (O_966,N_18140,N_19642);
xnor UO_967 (O_967,N_18570,N_19229);
nor UO_968 (O_968,N_19134,N_19394);
and UO_969 (O_969,N_18263,N_19491);
nor UO_970 (O_970,N_19894,N_19038);
nor UO_971 (O_971,N_19010,N_18005);
or UO_972 (O_972,N_18094,N_19727);
xor UO_973 (O_973,N_19638,N_19785);
and UO_974 (O_974,N_18188,N_18494);
and UO_975 (O_975,N_18401,N_18332);
nand UO_976 (O_976,N_19597,N_18394);
and UO_977 (O_977,N_19561,N_19820);
nand UO_978 (O_978,N_18036,N_18802);
or UO_979 (O_979,N_18486,N_19662);
nand UO_980 (O_980,N_18289,N_18631);
or UO_981 (O_981,N_19858,N_18096);
nand UO_982 (O_982,N_19692,N_19933);
nand UO_983 (O_983,N_19702,N_18097);
nor UO_984 (O_984,N_18192,N_18268);
xor UO_985 (O_985,N_18573,N_19938);
nor UO_986 (O_986,N_18436,N_18913);
xnor UO_987 (O_987,N_18888,N_19033);
nor UO_988 (O_988,N_19585,N_18704);
or UO_989 (O_989,N_19782,N_19222);
and UO_990 (O_990,N_19224,N_18788);
nor UO_991 (O_991,N_18132,N_19104);
nor UO_992 (O_992,N_18933,N_19569);
nand UO_993 (O_993,N_19240,N_19407);
and UO_994 (O_994,N_18222,N_19924);
nor UO_995 (O_995,N_19884,N_19501);
or UO_996 (O_996,N_18466,N_19300);
and UO_997 (O_997,N_18172,N_19451);
nand UO_998 (O_998,N_18647,N_18721);
xor UO_999 (O_999,N_19915,N_19026);
nor UO_1000 (O_1000,N_18974,N_19554);
and UO_1001 (O_1001,N_18176,N_18497);
or UO_1002 (O_1002,N_18925,N_19087);
nand UO_1003 (O_1003,N_19344,N_19029);
nand UO_1004 (O_1004,N_19344,N_18001);
or UO_1005 (O_1005,N_18585,N_19947);
and UO_1006 (O_1006,N_18868,N_18577);
and UO_1007 (O_1007,N_18086,N_18567);
nor UO_1008 (O_1008,N_18374,N_19232);
nand UO_1009 (O_1009,N_19723,N_19024);
nand UO_1010 (O_1010,N_18677,N_19892);
or UO_1011 (O_1011,N_18429,N_18983);
nor UO_1012 (O_1012,N_19229,N_19155);
nor UO_1013 (O_1013,N_18851,N_19607);
nand UO_1014 (O_1014,N_19696,N_18429);
xnor UO_1015 (O_1015,N_19790,N_19833);
nor UO_1016 (O_1016,N_19550,N_19189);
nor UO_1017 (O_1017,N_19476,N_19930);
and UO_1018 (O_1018,N_18623,N_18259);
and UO_1019 (O_1019,N_19755,N_19065);
nor UO_1020 (O_1020,N_19077,N_19980);
and UO_1021 (O_1021,N_19473,N_19725);
nand UO_1022 (O_1022,N_18459,N_18658);
or UO_1023 (O_1023,N_19698,N_19098);
xor UO_1024 (O_1024,N_19302,N_19812);
xor UO_1025 (O_1025,N_18615,N_19954);
nand UO_1026 (O_1026,N_18373,N_18809);
or UO_1027 (O_1027,N_19332,N_19614);
nand UO_1028 (O_1028,N_18088,N_19063);
and UO_1029 (O_1029,N_18884,N_18839);
nand UO_1030 (O_1030,N_18377,N_18108);
or UO_1031 (O_1031,N_18066,N_19661);
or UO_1032 (O_1032,N_19956,N_19622);
nor UO_1033 (O_1033,N_19087,N_18376);
nand UO_1034 (O_1034,N_19392,N_19774);
nor UO_1035 (O_1035,N_19156,N_18711);
nand UO_1036 (O_1036,N_18933,N_18785);
nand UO_1037 (O_1037,N_18298,N_18492);
nor UO_1038 (O_1038,N_18936,N_18732);
nor UO_1039 (O_1039,N_19495,N_19937);
or UO_1040 (O_1040,N_18236,N_18287);
or UO_1041 (O_1041,N_19577,N_18714);
and UO_1042 (O_1042,N_18167,N_19365);
or UO_1043 (O_1043,N_18857,N_19005);
and UO_1044 (O_1044,N_18109,N_19792);
nand UO_1045 (O_1045,N_19914,N_18164);
xor UO_1046 (O_1046,N_18833,N_18685);
xnor UO_1047 (O_1047,N_19325,N_19090);
and UO_1048 (O_1048,N_19344,N_18700);
nand UO_1049 (O_1049,N_18215,N_19075);
and UO_1050 (O_1050,N_19363,N_19725);
and UO_1051 (O_1051,N_18727,N_19034);
nand UO_1052 (O_1052,N_19674,N_19678);
and UO_1053 (O_1053,N_19945,N_18025);
nand UO_1054 (O_1054,N_18310,N_19718);
nand UO_1055 (O_1055,N_19832,N_19812);
or UO_1056 (O_1056,N_19393,N_18568);
or UO_1057 (O_1057,N_18085,N_19099);
nor UO_1058 (O_1058,N_18556,N_19240);
nor UO_1059 (O_1059,N_18702,N_18917);
and UO_1060 (O_1060,N_19355,N_18337);
or UO_1061 (O_1061,N_18117,N_19246);
nor UO_1062 (O_1062,N_19277,N_18180);
or UO_1063 (O_1063,N_18712,N_19282);
xor UO_1064 (O_1064,N_18886,N_18782);
or UO_1065 (O_1065,N_18001,N_19632);
nor UO_1066 (O_1066,N_18349,N_18458);
xor UO_1067 (O_1067,N_18364,N_18064);
nand UO_1068 (O_1068,N_18739,N_18916);
nor UO_1069 (O_1069,N_19831,N_19046);
or UO_1070 (O_1070,N_19029,N_18118);
nand UO_1071 (O_1071,N_18377,N_18703);
and UO_1072 (O_1072,N_18821,N_19661);
nand UO_1073 (O_1073,N_18254,N_19317);
and UO_1074 (O_1074,N_18761,N_19142);
or UO_1075 (O_1075,N_19531,N_18689);
nor UO_1076 (O_1076,N_18080,N_19128);
or UO_1077 (O_1077,N_19212,N_18222);
nor UO_1078 (O_1078,N_18902,N_18173);
nor UO_1079 (O_1079,N_19587,N_19352);
and UO_1080 (O_1080,N_19586,N_19984);
nand UO_1081 (O_1081,N_18048,N_19557);
and UO_1082 (O_1082,N_18877,N_18125);
nand UO_1083 (O_1083,N_19339,N_18864);
or UO_1084 (O_1084,N_19821,N_18885);
nand UO_1085 (O_1085,N_19683,N_19104);
or UO_1086 (O_1086,N_18793,N_18189);
nand UO_1087 (O_1087,N_18763,N_18130);
and UO_1088 (O_1088,N_18395,N_19153);
or UO_1089 (O_1089,N_19471,N_19780);
nor UO_1090 (O_1090,N_19927,N_18857);
or UO_1091 (O_1091,N_19591,N_18148);
and UO_1092 (O_1092,N_19074,N_19102);
and UO_1093 (O_1093,N_19497,N_18753);
or UO_1094 (O_1094,N_18819,N_18702);
or UO_1095 (O_1095,N_18952,N_18122);
or UO_1096 (O_1096,N_18921,N_19825);
nor UO_1097 (O_1097,N_19011,N_19062);
nand UO_1098 (O_1098,N_18389,N_19690);
xor UO_1099 (O_1099,N_19846,N_19814);
and UO_1100 (O_1100,N_19233,N_18218);
and UO_1101 (O_1101,N_18154,N_18567);
nor UO_1102 (O_1102,N_19877,N_18817);
or UO_1103 (O_1103,N_19985,N_19373);
nor UO_1104 (O_1104,N_18642,N_18901);
or UO_1105 (O_1105,N_19506,N_18182);
or UO_1106 (O_1106,N_19658,N_18149);
nor UO_1107 (O_1107,N_18014,N_18558);
nor UO_1108 (O_1108,N_19870,N_19162);
nand UO_1109 (O_1109,N_18141,N_18563);
or UO_1110 (O_1110,N_19808,N_19778);
nand UO_1111 (O_1111,N_18572,N_18633);
nand UO_1112 (O_1112,N_18804,N_18454);
nor UO_1113 (O_1113,N_19952,N_18763);
nor UO_1114 (O_1114,N_19067,N_19415);
nor UO_1115 (O_1115,N_18601,N_19649);
nor UO_1116 (O_1116,N_18965,N_19204);
nor UO_1117 (O_1117,N_19587,N_19091);
and UO_1118 (O_1118,N_18976,N_18464);
or UO_1119 (O_1119,N_19584,N_19170);
or UO_1120 (O_1120,N_18158,N_18481);
and UO_1121 (O_1121,N_19753,N_18355);
nor UO_1122 (O_1122,N_18580,N_18063);
xor UO_1123 (O_1123,N_18550,N_19928);
nor UO_1124 (O_1124,N_18848,N_18230);
nor UO_1125 (O_1125,N_19239,N_19181);
or UO_1126 (O_1126,N_18951,N_19749);
or UO_1127 (O_1127,N_19012,N_18551);
nor UO_1128 (O_1128,N_18161,N_18881);
or UO_1129 (O_1129,N_18650,N_19218);
xor UO_1130 (O_1130,N_19624,N_18935);
or UO_1131 (O_1131,N_18679,N_18877);
nor UO_1132 (O_1132,N_19309,N_19135);
and UO_1133 (O_1133,N_18822,N_19231);
nand UO_1134 (O_1134,N_18491,N_18323);
nand UO_1135 (O_1135,N_19598,N_18445);
and UO_1136 (O_1136,N_19423,N_18095);
or UO_1137 (O_1137,N_18498,N_19670);
nor UO_1138 (O_1138,N_19638,N_19344);
xnor UO_1139 (O_1139,N_18530,N_19770);
xnor UO_1140 (O_1140,N_18499,N_19596);
nand UO_1141 (O_1141,N_19379,N_18898);
nor UO_1142 (O_1142,N_19705,N_18123);
nand UO_1143 (O_1143,N_18123,N_19455);
nor UO_1144 (O_1144,N_18522,N_18357);
or UO_1145 (O_1145,N_18492,N_18933);
or UO_1146 (O_1146,N_18498,N_18046);
or UO_1147 (O_1147,N_19644,N_19116);
or UO_1148 (O_1148,N_19943,N_18729);
nand UO_1149 (O_1149,N_18460,N_18779);
and UO_1150 (O_1150,N_19006,N_18065);
xor UO_1151 (O_1151,N_18811,N_18736);
and UO_1152 (O_1152,N_18079,N_18761);
or UO_1153 (O_1153,N_19723,N_19472);
nand UO_1154 (O_1154,N_18236,N_19865);
and UO_1155 (O_1155,N_18750,N_19192);
xor UO_1156 (O_1156,N_18645,N_18996);
and UO_1157 (O_1157,N_19907,N_19716);
and UO_1158 (O_1158,N_19730,N_18019);
nor UO_1159 (O_1159,N_18496,N_19169);
or UO_1160 (O_1160,N_18114,N_18961);
nor UO_1161 (O_1161,N_18439,N_19696);
nor UO_1162 (O_1162,N_18336,N_18307);
or UO_1163 (O_1163,N_18409,N_18343);
and UO_1164 (O_1164,N_19304,N_18998);
and UO_1165 (O_1165,N_19191,N_18020);
nor UO_1166 (O_1166,N_18779,N_18295);
and UO_1167 (O_1167,N_18399,N_19981);
xnor UO_1168 (O_1168,N_18504,N_18606);
or UO_1169 (O_1169,N_18546,N_19502);
and UO_1170 (O_1170,N_19206,N_19293);
and UO_1171 (O_1171,N_18253,N_18383);
and UO_1172 (O_1172,N_19733,N_19126);
and UO_1173 (O_1173,N_18831,N_18553);
nor UO_1174 (O_1174,N_18267,N_18504);
nor UO_1175 (O_1175,N_18063,N_19870);
nor UO_1176 (O_1176,N_18022,N_18445);
or UO_1177 (O_1177,N_19712,N_19959);
nor UO_1178 (O_1178,N_19739,N_19553);
xor UO_1179 (O_1179,N_19366,N_18717);
and UO_1180 (O_1180,N_18025,N_19179);
and UO_1181 (O_1181,N_19466,N_18438);
and UO_1182 (O_1182,N_19702,N_19356);
nand UO_1183 (O_1183,N_19460,N_18597);
or UO_1184 (O_1184,N_19489,N_19323);
and UO_1185 (O_1185,N_19973,N_18891);
nand UO_1186 (O_1186,N_19914,N_18891);
nor UO_1187 (O_1187,N_19918,N_18057);
and UO_1188 (O_1188,N_18524,N_18250);
xor UO_1189 (O_1189,N_18906,N_19301);
xnor UO_1190 (O_1190,N_19096,N_19711);
nand UO_1191 (O_1191,N_19696,N_19131);
nor UO_1192 (O_1192,N_18598,N_18454);
nand UO_1193 (O_1193,N_18582,N_18697);
and UO_1194 (O_1194,N_19821,N_18945);
nor UO_1195 (O_1195,N_18203,N_19834);
xor UO_1196 (O_1196,N_19801,N_19438);
and UO_1197 (O_1197,N_19754,N_18101);
nand UO_1198 (O_1198,N_18590,N_19486);
or UO_1199 (O_1199,N_19728,N_18996);
nor UO_1200 (O_1200,N_19750,N_18195);
xnor UO_1201 (O_1201,N_19371,N_19317);
xnor UO_1202 (O_1202,N_19987,N_19387);
or UO_1203 (O_1203,N_19629,N_18516);
and UO_1204 (O_1204,N_18112,N_18586);
nand UO_1205 (O_1205,N_19286,N_19610);
xnor UO_1206 (O_1206,N_18007,N_18484);
nor UO_1207 (O_1207,N_18500,N_18954);
nor UO_1208 (O_1208,N_19450,N_18595);
nor UO_1209 (O_1209,N_19650,N_18210);
nor UO_1210 (O_1210,N_18942,N_18806);
nand UO_1211 (O_1211,N_19402,N_18593);
or UO_1212 (O_1212,N_18577,N_18520);
and UO_1213 (O_1213,N_18792,N_18069);
nor UO_1214 (O_1214,N_19103,N_19424);
nand UO_1215 (O_1215,N_19686,N_18467);
nand UO_1216 (O_1216,N_18600,N_18566);
and UO_1217 (O_1217,N_19218,N_18333);
and UO_1218 (O_1218,N_18616,N_18523);
nor UO_1219 (O_1219,N_18179,N_19025);
or UO_1220 (O_1220,N_19881,N_18824);
or UO_1221 (O_1221,N_19452,N_19833);
nor UO_1222 (O_1222,N_18134,N_18296);
or UO_1223 (O_1223,N_18814,N_18562);
nand UO_1224 (O_1224,N_18596,N_19289);
nor UO_1225 (O_1225,N_19592,N_18673);
nand UO_1226 (O_1226,N_19009,N_19522);
and UO_1227 (O_1227,N_18789,N_18687);
nand UO_1228 (O_1228,N_19563,N_18816);
or UO_1229 (O_1229,N_19261,N_19015);
xor UO_1230 (O_1230,N_18869,N_18993);
xnor UO_1231 (O_1231,N_18671,N_18430);
and UO_1232 (O_1232,N_19197,N_19687);
nor UO_1233 (O_1233,N_19332,N_18243);
nor UO_1234 (O_1234,N_19753,N_19077);
nand UO_1235 (O_1235,N_18574,N_18587);
xnor UO_1236 (O_1236,N_19644,N_18243);
or UO_1237 (O_1237,N_19402,N_18392);
and UO_1238 (O_1238,N_18897,N_19169);
nor UO_1239 (O_1239,N_19676,N_18006);
and UO_1240 (O_1240,N_18042,N_18476);
nand UO_1241 (O_1241,N_19314,N_18969);
nor UO_1242 (O_1242,N_18336,N_19710);
or UO_1243 (O_1243,N_18162,N_18261);
nand UO_1244 (O_1244,N_18192,N_18444);
nor UO_1245 (O_1245,N_19870,N_18214);
nand UO_1246 (O_1246,N_18810,N_19242);
xor UO_1247 (O_1247,N_18736,N_18261);
xor UO_1248 (O_1248,N_18247,N_19080);
and UO_1249 (O_1249,N_18202,N_18453);
and UO_1250 (O_1250,N_19064,N_18315);
or UO_1251 (O_1251,N_19509,N_19619);
or UO_1252 (O_1252,N_18237,N_19393);
nand UO_1253 (O_1253,N_18008,N_18593);
nand UO_1254 (O_1254,N_19021,N_19652);
xnor UO_1255 (O_1255,N_19453,N_18135);
and UO_1256 (O_1256,N_18765,N_18214);
xnor UO_1257 (O_1257,N_19819,N_18959);
or UO_1258 (O_1258,N_18623,N_18882);
or UO_1259 (O_1259,N_19449,N_19212);
or UO_1260 (O_1260,N_19621,N_18094);
or UO_1261 (O_1261,N_19550,N_18597);
and UO_1262 (O_1262,N_18613,N_18619);
and UO_1263 (O_1263,N_18619,N_19848);
nor UO_1264 (O_1264,N_18870,N_19952);
nor UO_1265 (O_1265,N_18166,N_18065);
nor UO_1266 (O_1266,N_19785,N_18340);
nand UO_1267 (O_1267,N_18587,N_19869);
and UO_1268 (O_1268,N_18441,N_19561);
or UO_1269 (O_1269,N_19283,N_19954);
nand UO_1270 (O_1270,N_19109,N_18051);
and UO_1271 (O_1271,N_18393,N_19042);
or UO_1272 (O_1272,N_19969,N_19641);
and UO_1273 (O_1273,N_19744,N_19652);
xnor UO_1274 (O_1274,N_18800,N_18953);
nor UO_1275 (O_1275,N_18861,N_19622);
and UO_1276 (O_1276,N_19220,N_19084);
nand UO_1277 (O_1277,N_19231,N_19995);
or UO_1278 (O_1278,N_18464,N_18069);
and UO_1279 (O_1279,N_19133,N_19268);
nand UO_1280 (O_1280,N_19819,N_19152);
or UO_1281 (O_1281,N_18163,N_18651);
and UO_1282 (O_1282,N_18897,N_18386);
and UO_1283 (O_1283,N_18658,N_19873);
or UO_1284 (O_1284,N_19964,N_19016);
or UO_1285 (O_1285,N_18644,N_19114);
and UO_1286 (O_1286,N_18442,N_18961);
or UO_1287 (O_1287,N_18910,N_18863);
or UO_1288 (O_1288,N_18221,N_18523);
and UO_1289 (O_1289,N_19367,N_18841);
and UO_1290 (O_1290,N_18893,N_19311);
nor UO_1291 (O_1291,N_18924,N_18405);
nor UO_1292 (O_1292,N_19353,N_18679);
xnor UO_1293 (O_1293,N_19770,N_18351);
xor UO_1294 (O_1294,N_19636,N_19690);
nand UO_1295 (O_1295,N_19017,N_18668);
nor UO_1296 (O_1296,N_19924,N_19724);
or UO_1297 (O_1297,N_18582,N_18830);
and UO_1298 (O_1298,N_19981,N_18640);
nor UO_1299 (O_1299,N_18479,N_18024);
xor UO_1300 (O_1300,N_19533,N_18220);
or UO_1301 (O_1301,N_19751,N_18822);
or UO_1302 (O_1302,N_19703,N_19354);
nand UO_1303 (O_1303,N_19853,N_18249);
nor UO_1304 (O_1304,N_19809,N_19627);
nand UO_1305 (O_1305,N_18515,N_18276);
nand UO_1306 (O_1306,N_19172,N_18998);
or UO_1307 (O_1307,N_18947,N_19879);
or UO_1308 (O_1308,N_18533,N_19455);
and UO_1309 (O_1309,N_18205,N_18929);
and UO_1310 (O_1310,N_18824,N_19943);
nor UO_1311 (O_1311,N_18022,N_18867);
nand UO_1312 (O_1312,N_19584,N_19273);
and UO_1313 (O_1313,N_19263,N_19559);
and UO_1314 (O_1314,N_18588,N_18313);
and UO_1315 (O_1315,N_18161,N_18810);
and UO_1316 (O_1316,N_19307,N_18729);
and UO_1317 (O_1317,N_18363,N_18278);
nand UO_1318 (O_1318,N_18334,N_19393);
xnor UO_1319 (O_1319,N_19348,N_18790);
nor UO_1320 (O_1320,N_19461,N_19972);
and UO_1321 (O_1321,N_19599,N_19630);
nand UO_1322 (O_1322,N_19412,N_18993);
xnor UO_1323 (O_1323,N_19555,N_19155);
or UO_1324 (O_1324,N_18718,N_19285);
nand UO_1325 (O_1325,N_19908,N_18894);
or UO_1326 (O_1326,N_19061,N_18573);
or UO_1327 (O_1327,N_18638,N_19363);
or UO_1328 (O_1328,N_18696,N_18805);
nor UO_1329 (O_1329,N_18674,N_18724);
xnor UO_1330 (O_1330,N_19271,N_19720);
and UO_1331 (O_1331,N_19935,N_19215);
nand UO_1332 (O_1332,N_19164,N_18872);
and UO_1333 (O_1333,N_18706,N_18326);
nor UO_1334 (O_1334,N_19430,N_19081);
and UO_1335 (O_1335,N_18360,N_18308);
and UO_1336 (O_1336,N_18439,N_19721);
nand UO_1337 (O_1337,N_19058,N_18199);
and UO_1338 (O_1338,N_19941,N_19681);
nand UO_1339 (O_1339,N_18470,N_18373);
nor UO_1340 (O_1340,N_19740,N_18976);
or UO_1341 (O_1341,N_19632,N_19792);
nand UO_1342 (O_1342,N_19083,N_18868);
nor UO_1343 (O_1343,N_19894,N_19711);
nand UO_1344 (O_1344,N_18477,N_18120);
nor UO_1345 (O_1345,N_18904,N_18612);
and UO_1346 (O_1346,N_18032,N_18656);
or UO_1347 (O_1347,N_18566,N_18172);
nand UO_1348 (O_1348,N_18671,N_18497);
nand UO_1349 (O_1349,N_18205,N_19169);
xor UO_1350 (O_1350,N_19981,N_18798);
nand UO_1351 (O_1351,N_19719,N_18663);
and UO_1352 (O_1352,N_18512,N_18174);
nand UO_1353 (O_1353,N_18129,N_18571);
nor UO_1354 (O_1354,N_18295,N_19724);
and UO_1355 (O_1355,N_19724,N_18119);
nand UO_1356 (O_1356,N_19314,N_19000);
and UO_1357 (O_1357,N_19661,N_18779);
or UO_1358 (O_1358,N_19852,N_19208);
nand UO_1359 (O_1359,N_19718,N_19982);
nor UO_1360 (O_1360,N_18635,N_19506);
nand UO_1361 (O_1361,N_19896,N_18234);
and UO_1362 (O_1362,N_19973,N_18411);
nand UO_1363 (O_1363,N_18299,N_18040);
or UO_1364 (O_1364,N_18893,N_19973);
or UO_1365 (O_1365,N_18390,N_18146);
nor UO_1366 (O_1366,N_19636,N_19413);
nor UO_1367 (O_1367,N_19069,N_18605);
or UO_1368 (O_1368,N_18212,N_19891);
or UO_1369 (O_1369,N_18295,N_19925);
or UO_1370 (O_1370,N_19030,N_19805);
and UO_1371 (O_1371,N_19855,N_19250);
nor UO_1372 (O_1372,N_18309,N_18051);
or UO_1373 (O_1373,N_19245,N_18600);
nor UO_1374 (O_1374,N_18067,N_19422);
and UO_1375 (O_1375,N_19202,N_18188);
nand UO_1376 (O_1376,N_19592,N_19834);
and UO_1377 (O_1377,N_18621,N_19120);
xor UO_1378 (O_1378,N_19884,N_18112);
and UO_1379 (O_1379,N_19179,N_19668);
nor UO_1380 (O_1380,N_18264,N_18626);
nand UO_1381 (O_1381,N_18104,N_18981);
nor UO_1382 (O_1382,N_18825,N_19725);
nor UO_1383 (O_1383,N_19419,N_19820);
and UO_1384 (O_1384,N_19943,N_19913);
xor UO_1385 (O_1385,N_19406,N_19940);
nor UO_1386 (O_1386,N_18068,N_19782);
and UO_1387 (O_1387,N_18238,N_18510);
nor UO_1388 (O_1388,N_19689,N_18270);
and UO_1389 (O_1389,N_18437,N_19178);
nand UO_1390 (O_1390,N_18650,N_19072);
or UO_1391 (O_1391,N_19524,N_19534);
and UO_1392 (O_1392,N_19953,N_19661);
or UO_1393 (O_1393,N_18212,N_18909);
nand UO_1394 (O_1394,N_18481,N_19507);
nor UO_1395 (O_1395,N_19175,N_19382);
or UO_1396 (O_1396,N_18944,N_19120);
and UO_1397 (O_1397,N_18238,N_19501);
and UO_1398 (O_1398,N_18883,N_18861);
and UO_1399 (O_1399,N_19892,N_18921);
nand UO_1400 (O_1400,N_18103,N_18033);
xor UO_1401 (O_1401,N_19231,N_19682);
nand UO_1402 (O_1402,N_18621,N_18140);
and UO_1403 (O_1403,N_18833,N_18924);
nor UO_1404 (O_1404,N_18090,N_19358);
nor UO_1405 (O_1405,N_18546,N_19080);
and UO_1406 (O_1406,N_19861,N_19548);
or UO_1407 (O_1407,N_19280,N_18816);
nand UO_1408 (O_1408,N_18427,N_18268);
nor UO_1409 (O_1409,N_19343,N_18289);
and UO_1410 (O_1410,N_19960,N_19942);
or UO_1411 (O_1411,N_19295,N_19317);
nor UO_1412 (O_1412,N_18552,N_19789);
and UO_1413 (O_1413,N_19571,N_19200);
and UO_1414 (O_1414,N_18578,N_19382);
xnor UO_1415 (O_1415,N_18387,N_19185);
nor UO_1416 (O_1416,N_19167,N_19302);
xnor UO_1417 (O_1417,N_19190,N_18360);
nand UO_1418 (O_1418,N_19883,N_19148);
or UO_1419 (O_1419,N_19974,N_18340);
and UO_1420 (O_1420,N_19829,N_19823);
nor UO_1421 (O_1421,N_18248,N_19474);
or UO_1422 (O_1422,N_19390,N_18582);
nand UO_1423 (O_1423,N_18542,N_18782);
and UO_1424 (O_1424,N_19017,N_19443);
xnor UO_1425 (O_1425,N_19107,N_19552);
xor UO_1426 (O_1426,N_18780,N_18258);
nand UO_1427 (O_1427,N_19455,N_19391);
or UO_1428 (O_1428,N_18014,N_19636);
nor UO_1429 (O_1429,N_18197,N_19962);
xor UO_1430 (O_1430,N_19396,N_19727);
or UO_1431 (O_1431,N_18270,N_19856);
or UO_1432 (O_1432,N_18460,N_18960);
nor UO_1433 (O_1433,N_19102,N_19740);
or UO_1434 (O_1434,N_18994,N_19407);
nand UO_1435 (O_1435,N_19980,N_19039);
or UO_1436 (O_1436,N_18643,N_19600);
nor UO_1437 (O_1437,N_18826,N_19772);
or UO_1438 (O_1438,N_18625,N_18446);
nor UO_1439 (O_1439,N_18179,N_18130);
nor UO_1440 (O_1440,N_18587,N_19284);
nand UO_1441 (O_1441,N_19931,N_19977);
and UO_1442 (O_1442,N_18963,N_19171);
nand UO_1443 (O_1443,N_18134,N_19112);
and UO_1444 (O_1444,N_19777,N_18279);
nor UO_1445 (O_1445,N_18031,N_18694);
xor UO_1446 (O_1446,N_18326,N_19900);
and UO_1447 (O_1447,N_19577,N_18156);
nor UO_1448 (O_1448,N_18691,N_19702);
or UO_1449 (O_1449,N_19305,N_19506);
nor UO_1450 (O_1450,N_18339,N_19889);
nor UO_1451 (O_1451,N_18626,N_19442);
nand UO_1452 (O_1452,N_18232,N_19870);
xnor UO_1453 (O_1453,N_18579,N_18005);
or UO_1454 (O_1454,N_19485,N_19244);
nand UO_1455 (O_1455,N_19959,N_19392);
or UO_1456 (O_1456,N_19976,N_19032);
nand UO_1457 (O_1457,N_19743,N_19681);
nor UO_1458 (O_1458,N_18450,N_19405);
and UO_1459 (O_1459,N_18002,N_18614);
nand UO_1460 (O_1460,N_19535,N_19397);
and UO_1461 (O_1461,N_18676,N_19662);
or UO_1462 (O_1462,N_18380,N_18257);
nand UO_1463 (O_1463,N_18698,N_18170);
xor UO_1464 (O_1464,N_19028,N_19632);
and UO_1465 (O_1465,N_19916,N_19623);
nand UO_1466 (O_1466,N_18202,N_19191);
or UO_1467 (O_1467,N_19216,N_19678);
and UO_1468 (O_1468,N_19082,N_19902);
or UO_1469 (O_1469,N_18996,N_18388);
nor UO_1470 (O_1470,N_18141,N_18996);
xor UO_1471 (O_1471,N_18174,N_19963);
nand UO_1472 (O_1472,N_18006,N_19282);
or UO_1473 (O_1473,N_18621,N_19148);
nand UO_1474 (O_1474,N_18123,N_19598);
nand UO_1475 (O_1475,N_18161,N_19629);
nor UO_1476 (O_1476,N_18074,N_19168);
and UO_1477 (O_1477,N_19950,N_18479);
xnor UO_1478 (O_1478,N_18372,N_19840);
or UO_1479 (O_1479,N_19421,N_18250);
nor UO_1480 (O_1480,N_19452,N_18908);
or UO_1481 (O_1481,N_19504,N_18491);
or UO_1482 (O_1482,N_18400,N_19426);
and UO_1483 (O_1483,N_19893,N_18026);
or UO_1484 (O_1484,N_18779,N_18190);
or UO_1485 (O_1485,N_19308,N_19897);
or UO_1486 (O_1486,N_18129,N_18608);
or UO_1487 (O_1487,N_18985,N_18994);
nand UO_1488 (O_1488,N_19273,N_19220);
and UO_1489 (O_1489,N_18396,N_19554);
nor UO_1490 (O_1490,N_19896,N_18151);
nand UO_1491 (O_1491,N_18935,N_18195);
and UO_1492 (O_1492,N_19986,N_19592);
nor UO_1493 (O_1493,N_18978,N_19589);
nand UO_1494 (O_1494,N_19915,N_19358);
or UO_1495 (O_1495,N_19594,N_19859);
xnor UO_1496 (O_1496,N_18943,N_18820);
nor UO_1497 (O_1497,N_19422,N_18293);
nand UO_1498 (O_1498,N_18139,N_18379);
or UO_1499 (O_1499,N_18342,N_18922);
nand UO_1500 (O_1500,N_18579,N_19286);
and UO_1501 (O_1501,N_18130,N_19506);
or UO_1502 (O_1502,N_18789,N_19975);
or UO_1503 (O_1503,N_19298,N_19421);
or UO_1504 (O_1504,N_19224,N_19707);
or UO_1505 (O_1505,N_19827,N_18424);
nor UO_1506 (O_1506,N_19728,N_19850);
and UO_1507 (O_1507,N_18357,N_19430);
and UO_1508 (O_1508,N_18313,N_18277);
or UO_1509 (O_1509,N_19822,N_18894);
nor UO_1510 (O_1510,N_18231,N_18824);
and UO_1511 (O_1511,N_18194,N_19130);
xor UO_1512 (O_1512,N_19582,N_18038);
nor UO_1513 (O_1513,N_19565,N_18922);
xor UO_1514 (O_1514,N_18650,N_18035);
or UO_1515 (O_1515,N_18896,N_19818);
xnor UO_1516 (O_1516,N_19222,N_18548);
nor UO_1517 (O_1517,N_18564,N_19576);
nor UO_1518 (O_1518,N_18299,N_19218);
nand UO_1519 (O_1519,N_18895,N_18694);
and UO_1520 (O_1520,N_18681,N_18538);
or UO_1521 (O_1521,N_19577,N_18266);
xnor UO_1522 (O_1522,N_19735,N_19135);
xnor UO_1523 (O_1523,N_19225,N_19297);
and UO_1524 (O_1524,N_19120,N_18048);
xnor UO_1525 (O_1525,N_19530,N_18836);
nor UO_1526 (O_1526,N_18458,N_18397);
or UO_1527 (O_1527,N_19591,N_19048);
or UO_1528 (O_1528,N_18101,N_19468);
nor UO_1529 (O_1529,N_19576,N_18569);
nor UO_1530 (O_1530,N_19607,N_19548);
nor UO_1531 (O_1531,N_19412,N_19122);
or UO_1532 (O_1532,N_18394,N_18402);
or UO_1533 (O_1533,N_19853,N_18981);
nand UO_1534 (O_1534,N_19789,N_19640);
nand UO_1535 (O_1535,N_18165,N_19841);
nor UO_1536 (O_1536,N_19840,N_18247);
or UO_1537 (O_1537,N_18634,N_19566);
nand UO_1538 (O_1538,N_19248,N_18384);
or UO_1539 (O_1539,N_18463,N_18689);
nor UO_1540 (O_1540,N_18855,N_19692);
xnor UO_1541 (O_1541,N_19836,N_19452);
and UO_1542 (O_1542,N_19781,N_19404);
xnor UO_1543 (O_1543,N_18801,N_19371);
or UO_1544 (O_1544,N_18651,N_19745);
nand UO_1545 (O_1545,N_18401,N_18185);
xor UO_1546 (O_1546,N_18835,N_19987);
nor UO_1547 (O_1547,N_19506,N_19398);
or UO_1548 (O_1548,N_19637,N_18949);
nor UO_1549 (O_1549,N_19738,N_19953);
and UO_1550 (O_1550,N_18882,N_18701);
and UO_1551 (O_1551,N_19052,N_19877);
nand UO_1552 (O_1552,N_18225,N_18720);
nor UO_1553 (O_1553,N_19608,N_18156);
and UO_1554 (O_1554,N_19133,N_18339);
or UO_1555 (O_1555,N_18656,N_19781);
xnor UO_1556 (O_1556,N_18482,N_19829);
and UO_1557 (O_1557,N_19830,N_18389);
nor UO_1558 (O_1558,N_19581,N_19892);
or UO_1559 (O_1559,N_19150,N_19361);
or UO_1560 (O_1560,N_18435,N_18223);
and UO_1561 (O_1561,N_18881,N_18632);
nand UO_1562 (O_1562,N_19852,N_18260);
nand UO_1563 (O_1563,N_18904,N_19129);
nor UO_1564 (O_1564,N_18744,N_19130);
or UO_1565 (O_1565,N_18077,N_19232);
nand UO_1566 (O_1566,N_19893,N_19316);
or UO_1567 (O_1567,N_18174,N_18010);
or UO_1568 (O_1568,N_19890,N_19147);
or UO_1569 (O_1569,N_19257,N_18670);
nor UO_1570 (O_1570,N_19259,N_18941);
nor UO_1571 (O_1571,N_18550,N_19345);
and UO_1572 (O_1572,N_19097,N_19073);
xor UO_1573 (O_1573,N_19254,N_18281);
nand UO_1574 (O_1574,N_18532,N_19291);
nor UO_1575 (O_1575,N_19242,N_19794);
nand UO_1576 (O_1576,N_19492,N_18737);
and UO_1577 (O_1577,N_18034,N_19818);
nand UO_1578 (O_1578,N_19616,N_19999);
and UO_1579 (O_1579,N_18123,N_19006);
or UO_1580 (O_1580,N_18983,N_18516);
nand UO_1581 (O_1581,N_18812,N_18766);
and UO_1582 (O_1582,N_18241,N_18004);
or UO_1583 (O_1583,N_18847,N_19967);
and UO_1584 (O_1584,N_18999,N_19031);
nor UO_1585 (O_1585,N_19255,N_18037);
xor UO_1586 (O_1586,N_18100,N_18232);
nor UO_1587 (O_1587,N_19130,N_19683);
nor UO_1588 (O_1588,N_18589,N_19723);
and UO_1589 (O_1589,N_19884,N_18705);
and UO_1590 (O_1590,N_19349,N_19555);
nand UO_1591 (O_1591,N_19350,N_18863);
and UO_1592 (O_1592,N_18697,N_18379);
nand UO_1593 (O_1593,N_19723,N_18758);
nand UO_1594 (O_1594,N_18746,N_19154);
xnor UO_1595 (O_1595,N_18434,N_19089);
and UO_1596 (O_1596,N_18190,N_19318);
and UO_1597 (O_1597,N_19750,N_19369);
and UO_1598 (O_1598,N_18940,N_19751);
xnor UO_1599 (O_1599,N_18589,N_19648);
nand UO_1600 (O_1600,N_18583,N_18700);
and UO_1601 (O_1601,N_18395,N_19081);
nand UO_1602 (O_1602,N_19642,N_19020);
nand UO_1603 (O_1603,N_18164,N_18855);
xnor UO_1604 (O_1604,N_18164,N_19731);
nand UO_1605 (O_1605,N_19604,N_18395);
and UO_1606 (O_1606,N_19141,N_18899);
and UO_1607 (O_1607,N_18563,N_19575);
nor UO_1608 (O_1608,N_19434,N_19560);
nand UO_1609 (O_1609,N_18339,N_19345);
and UO_1610 (O_1610,N_18846,N_19368);
nand UO_1611 (O_1611,N_18050,N_19100);
and UO_1612 (O_1612,N_18222,N_19349);
xor UO_1613 (O_1613,N_19027,N_19563);
nand UO_1614 (O_1614,N_18887,N_18752);
nand UO_1615 (O_1615,N_18837,N_18934);
and UO_1616 (O_1616,N_19275,N_18044);
nand UO_1617 (O_1617,N_18706,N_18937);
nand UO_1618 (O_1618,N_18561,N_18322);
and UO_1619 (O_1619,N_18847,N_19289);
or UO_1620 (O_1620,N_19652,N_19901);
nand UO_1621 (O_1621,N_19410,N_18575);
or UO_1622 (O_1622,N_18504,N_19922);
nor UO_1623 (O_1623,N_18710,N_18326);
nand UO_1624 (O_1624,N_19725,N_18244);
xor UO_1625 (O_1625,N_18820,N_18790);
or UO_1626 (O_1626,N_18830,N_18011);
nor UO_1627 (O_1627,N_19639,N_18122);
or UO_1628 (O_1628,N_18221,N_19062);
nand UO_1629 (O_1629,N_19372,N_18759);
xnor UO_1630 (O_1630,N_19433,N_19949);
or UO_1631 (O_1631,N_19206,N_18451);
and UO_1632 (O_1632,N_18881,N_18501);
nor UO_1633 (O_1633,N_19906,N_19115);
and UO_1634 (O_1634,N_19678,N_18792);
nor UO_1635 (O_1635,N_18870,N_18092);
nand UO_1636 (O_1636,N_18381,N_18409);
nor UO_1637 (O_1637,N_19419,N_19725);
or UO_1638 (O_1638,N_18534,N_18447);
nor UO_1639 (O_1639,N_19466,N_18373);
and UO_1640 (O_1640,N_19673,N_18703);
nor UO_1641 (O_1641,N_18489,N_19671);
or UO_1642 (O_1642,N_19518,N_19770);
or UO_1643 (O_1643,N_19448,N_19085);
nor UO_1644 (O_1644,N_19338,N_18449);
nand UO_1645 (O_1645,N_19125,N_19722);
and UO_1646 (O_1646,N_19392,N_18618);
and UO_1647 (O_1647,N_18408,N_19127);
xor UO_1648 (O_1648,N_18839,N_18038);
nand UO_1649 (O_1649,N_18429,N_19941);
nor UO_1650 (O_1650,N_19209,N_19219);
or UO_1651 (O_1651,N_19418,N_19473);
or UO_1652 (O_1652,N_19744,N_19330);
nand UO_1653 (O_1653,N_18236,N_18688);
and UO_1654 (O_1654,N_19123,N_18295);
nor UO_1655 (O_1655,N_19572,N_18431);
xnor UO_1656 (O_1656,N_19920,N_19938);
nand UO_1657 (O_1657,N_18645,N_18962);
nand UO_1658 (O_1658,N_19200,N_19795);
or UO_1659 (O_1659,N_18769,N_18150);
or UO_1660 (O_1660,N_19788,N_18419);
or UO_1661 (O_1661,N_19550,N_18314);
nand UO_1662 (O_1662,N_19042,N_19017);
nand UO_1663 (O_1663,N_18035,N_19144);
nor UO_1664 (O_1664,N_18369,N_19845);
xnor UO_1665 (O_1665,N_18920,N_18042);
and UO_1666 (O_1666,N_18709,N_18067);
and UO_1667 (O_1667,N_19840,N_18314);
nand UO_1668 (O_1668,N_19352,N_18151);
and UO_1669 (O_1669,N_19459,N_18587);
or UO_1670 (O_1670,N_18870,N_18603);
nor UO_1671 (O_1671,N_19317,N_18697);
and UO_1672 (O_1672,N_18304,N_18204);
or UO_1673 (O_1673,N_19267,N_19851);
and UO_1674 (O_1674,N_18432,N_18371);
xnor UO_1675 (O_1675,N_18984,N_18561);
or UO_1676 (O_1676,N_18769,N_18060);
nand UO_1677 (O_1677,N_18861,N_18024);
nand UO_1678 (O_1678,N_19111,N_18621);
nor UO_1679 (O_1679,N_19363,N_18468);
and UO_1680 (O_1680,N_19003,N_19274);
and UO_1681 (O_1681,N_18164,N_19068);
xnor UO_1682 (O_1682,N_18449,N_18164);
or UO_1683 (O_1683,N_19472,N_19797);
nor UO_1684 (O_1684,N_19896,N_19145);
or UO_1685 (O_1685,N_18154,N_19795);
and UO_1686 (O_1686,N_18941,N_19796);
or UO_1687 (O_1687,N_19504,N_19641);
nor UO_1688 (O_1688,N_19009,N_18678);
nand UO_1689 (O_1689,N_19301,N_19922);
nor UO_1690 (O_1690,N_19775,N_19448);
and UO_1691 (O_1691,N_18948,N_19001);
nor UO_1692 (O_1692,N_19044,N_18625);
nand UO_1693 (O_1693,N_18733,N_19607);
or UO_1694 (O_1694,N_18086,N_19067);
nand UO_1695 (O_1695,N_19267,N_18717);
or UO_1696 (O_1696,N_18283,N_18448);
or UO_1697 (O_1697,N_19751,N_18578);
or UO_1698 (O_1698,N_19397,N_19860);
xnor UO_1699 (O_1699,N_19632,N_19253);
and UO_1700 (O_1700,N_18634,N_18976);
and UO_1701 (O_1701,N_19842,N_18304);
and UO_1702 (O_1702,N_19671,N_18099);
nor UO_1703 (O_1703,N_19743,N_19483);
and UO_1704 (O_1704,N_18878,N_18954);
nor UO_1705 (O_1705,N_19720,N_18437);
nor UO_1706 (O_1706,N_18246,N_19818);
nor UO_1707 (O_1707,N_19356,N_19184);
nor UO_1708 (O_1708,N_18372,N_19380);
or UO_1709 (O_1709,N_19766,N_18805);
nor UO_1710 (O_1710,N_19968,N_19326);
or UO_1711 (O_1711,N_18984,N_18514);
nand UO_1712 (O_1712,N_18735,N_18875);
nor UO_1713 (O_1713,N_19499,N_18294);
or UO_1714 (O_1714,N_19828,N_19976);
nor UO_1715 (O_1715,N_19520,N_19357);
or UO_1716 (O_1716,N_19776,N_19363);
or UO_1717 (O_1717,N_19658,N_18069);
nand UO_1718 (O_1718,N_19950,N_19468);
or UO_1719 (O_1719,N_18051,N_19222);
nor UO_1720 (O_1720,N_19912,N_18086);
nor UO_1721 (O_1721,N_18836,N_19249);
or UO_1722 (O_1722,N_19235,N_19702);
or UO_1723 (O_1723,N_19308,N_18774);
nand UO_1724 (O_1724,N_18885,N_19499);
nor UO_1725 (O_1725,N_18602,N_18499);
nor UO_1726 (O_1726,N_19189,N_18793);
or UO_1727 (O_1727,N_18750,N_18304);
xnor UO_1728 (O_1728,N_18543,N_19386);
or UO_1729 (O_1729,N_19130,N_18220);
nor UO_1730 (O_1730,N_18018,N_19128);
or UO_1731 (O_1731,N_19808,N_19932);
and UO_1732 (O_1732,N_19554,N_19658);
xnor UO_1733 (O_1733,N_18401,N_19413);
nand UO_1734 (O_1734,N_18273,N_19828);
nand UO_1735 (O_1735,N_19394,N_19976);
nand UO_1736 (O_1736,N_18466,N_18765);
and UO_1737 (O_1737,N_18543,N_19910);
and UO_1738 (O_1738,N_18797,N_19955);
nand UO_1739 (O_1739,N_18656,N_19939);
or UO_1740 (O_1740,N_19078,N_18499);
nor UO_1741 (O_1741,N_18360,N_19413);
and UO_1742 (O_1742,N_18405,N_18691);
nor UO_1743 (O_1743,N_18190,N_19865);
xor UO_1744 (O_1744,N_18485,N_18285);
nor UO_1745 (O_1745,N_19629,N_18372);
or UO_1746 (O_1746,N_19333,N_19685);
nand UO_1747 (O_1747,N_19938,N_18052);
nor UO_1748 (O_1748,N_18275,N_18092);
nor UO_1749 (O_1749,N_19512,N_18651);
or UO_1750 (O_1750,N_19390,N_18211);
or UO_1751 (O_1751,N_19037,N_19865);
nor UO_1752 (O_1752,N_18837,N_19639);
nor UO_1753 (O_1753,N_19173,N_18880);
and UO_1754 (O_1754,N_18299,N_19848);
and UO_1755 (O_1755,N_19402,N_19755);
and UO_1756 (O_1756,N_19990,N_19139);
and UO_1757 (O_1757,N_19512,N_18405);
or UO_1758 (O_1758,N_19781,N_18088);
nor UO_1759 (O_1759,N_18971,N_18387);
and UO_1760 (O_1760,N_18390,N_18630);
and UO_1761 (O_1761,N_19229,N_18905);
nand UO_1762 (O_1762,N_18648,N_19672);
and UO_1763 (O_1763,N_18432,N_19253);
nor UO_1764 (O_1764,N_18074,N_19518);
or UO_1765 (O_1765,N_18731,N_19762);
or UO_1766 (O_1766,N_19204,N_19709);
nand UO_1767 (O_1767,N_18708,N_18816);
xnor UO_1768 (O_1768,N_18219,N_19770);
and UO_1769 (O_1769,N_19953,N_18651);
nor UO_1770 (O_1770,N_18826,N_18534);
or UO_1771 (O_1771,N_18821,N_18603);
and UO_1772 (O_1772,N_18937,N_19818);
and UO_1773 (O_1773,N_19005,N_18740);
nor UO_1774 (O_1774,N_19590,N_18749);
or UO_1775 (O_1775,N_19808,N_18711);
or UO_1776 (O_1776,N_19990,N_19141);
nand UO_1777 (O_1777,N_18535,N_18601);
and UO_1778 (O_1778,N_18698,N_19334);
xor UO_1779 (O_1779,N_19291,N_19777);
and UO_1780 (O_1780,N_18170,N_18178);
xor UO_1781 (O_1781,N_18062,N_18616);
and UO_1782 (O_1782,N_18163,N_19971);
and UO_1783 (O_1783,N_19295,N_19002);
nand UO_1784 (O_1784,N_18757,N_19435);
and UO_1785 (O_1785,N_18667,N_18683);
nand UO_1786 (O_1786,N_18712,N_18446);
or UO_1787 (O_1787,N_18792,N_19980);
and UO_1788 (O_1788,N_19145,N_19097);
or UO_1789 (O_1789,N_19052,N_18408);
and UO_1790 (O_1790,N_18584,N_19230);
nor UO_1791 (O_1791,N_19595,N_18712);
and UO_1792 (O_1792,N_18011,N_18515);
nor UO_1793 (O_1793,N_19278,N_18224);
and UO_1794 (O_1794,N_19324,N_19653);
xnor UO_1795 (O_1795,N_19886,N_18353);
or UO_1796 (O_1796,N_19820,N_19317);
and UO_1797 (O_1797,N_19460,N_19477);
nor UO_1798 (O_1798,N_19512,N_18694);
nor UO_1799 (O_1799,N_18908,N_18088);
and UO_1800 (O_1800,N_18720,N_19573);
and UO_1801 (O_1801,N_18206,N_18571);
nor UO_1802 (O_1802,N_19958,N_19500);
nor UO_1803 (O_1803,N_18035,N_19228);
or UO_1804 (O_1804,N_18085,N_18672);
or UO_1805 (O_1805,N_18208,N_19210);
and UO_1806 (O_1806,N_19709,N_19876);
and UO_1807 (O_1807,N_18669,N_18032);
xnor UO_1808 (O_1808,N_19504,N_18362);
nand UO_1809 (O_1809,N_18056,N_19083);
nor UO_1810 (O_1810,N_18501,N_19067);
xnor UO_1811 (O_1811,N_18583,N_18159);
nor UO_1812 (O_1812,N_18477,N_18429);
nand UO_1813 (O_1813,N_18849,N_19861);
or UO_1814 (O_1814,N_18010,N_18595);
or UO_1815 (O_1815,N_19122,N_19223);
or UO_1816 (O_1816,N_18956,N_19801);
nor UO_1817 (O_1817,N_19929,N_18452);
or UO_1818 (O_1818,N_19008,N_18886);
nand UO_1819 (O_1819,N_18198,N_19214);
xor UO_1820 (O_1820,N_18396,N_19596);
nand UO_1821 (O_1821,N_19809,N_18424);
nand UO_1822 (O_1822,N_19813,N_18748);
or UO_1823 (O_1823,N_18696,N_18483);
nor UO_1824 (O_1824,N_18872,N_19192);
nand UO_1825 (O_1825,N_19058,N_19351);
or UO_1826 (O_1826,N_19825,N_19194);
nand UO_1827 (O_1827,N_19759,N_18850);
nor UO_1828 (O_1828,N_19758,N_18643);
nand UO_1829 (O_1829,N_18927,N_18207);
xnor UO_1830 (O_1830,N_18233,N_19797);
nor UO_1831 (O_1831,N_18266,N_19210);
or UO_1832 (O_1832,N_19210,N_18205);
nand UO_1833 (O_1833,N_18819,N_19843);
and UO_1834 (O_1834,N_19833,N_19327);
nand UO_1835 (O_1835,N_18839,N_19329);
nor UO_1836 (O_1836,N_19123,N_19016);
or UO_1837 (O_1837,N_19167,N_18955);
or UO_1838 (O_1838,N_19547,N_19292);
or UO_1839 (O_1839,N_19661,N_19821);
nand UO_1840 (O_1840,N_19851,N_18462);
and UO_1841 (O_1841,N_19912,N_19009);
and UO_1842 (O_1842,N_18882,N_18104);
nand UO_1843 (O_1843,N_19406,N_19203);
nand UO_1844 (O_1844,N_19430,N_19385);
or UO_1845 (O_1845,N_19869,N_18381);
nor UO_1846 (O_1846,N_19316,N_18193);
nor UO_1847 (O_1847,N_19452,N_19601);
and UO_1848 (O_1848,N_19603,N_18140);
or UO_1849 (O_1849,N_19930,N_19967);
or UO_1850 (O_1850,N_18113,N_19970);
nand UO_1851 (O_1851,N_19202,N_19605);
nand UO_1852 (O_1852,N_18184,N_18877);
and UO_1853 (O_1853,N_19630,N_19992);
nand UO_1854 (O_1854,N_19876,N_19616);
nor UO_1855 (O_1855,N_18403,N_19834);
nand UO_1856 (O_1856,N_19990,N_18209);
nor UO_1857 (O_1857,N_18377,N_19155);
nor UO_1858 (O_1858,N_19947,N_19491);
nand UO_1859 (O_1859,N_19091,N_19926);
or UO_1860 (O_1860,N_19161,N_18254);
nor UO_1861 (O_1861,N_18353,N_18469);
nand UO_1862 (O_1862,N_18199,N_19475);
nand UO_1863 (O_1863,N_18656,N_18227);
nor UO_1864 (O_1864,N_18125,N_18711);
and UO_1865 (O_1865,N_18423,N_18308);
nand UO_1866 (O_1866,N_18687,N_18222);
nand UO_1867 (O_1867,N_19715,N_18144);
nand UO_1868 (O_1868,N_18859,N_18324);
or UO_1869 (O_1869,N_18210,N_19461);
and UO_1870 (O_1870,N_18550,N_18834);
nand UO_1871 (O_1871,N_18324,N_18318);
nand UO_1872 (O_1872,N_18385,N_18045);
and UO_1873 (O_1873,N_18801,N_18631);
or UO_1874 (O_1874,N_19457,N_18400);
nand UO_1875 (O_1875,N_18547,N_19701);
nand UO_1876 (O_1876,N_19474,N_18724);
nor UO_1877 (O_1877,N_18727,N_18794);
nand UO_1878 (O_1878,N_19772,N_19277);
nand UO_1879 (O_1879,N_18289,N_18966);
xor UO_1880 (O_1880,N_19787,N_18291);
nand UO_1881 (O_1881,N_19372,N_19301);
or UO_1882 (O_1882,N_18529,N_19173);
or UO_1883 (O_1883,N_19344,N_19621);
and UO_1884 (O_1884,N_18563,N_18040);
or UO_1885 (O_1885,N_19357,N_19613);
nand UO_1886 (O_1886,N_18998,N_19128);
and UO_1887 (O_1887,N_18435,N_19852);
or UO_1888 (O_1888,N_19980,N_18560);
and UO_1889 (O_1889,N_18658,N_19658);
and UO_1890 (O_1890,N_19538,N_18785);
or UO_1891 (O_1891,N_18693,N_18219);
nand UO_1892 (O_1892,N_19119,N_18487);
or UO_1893 (O_1893,N_19757,N_19731);
or UO_1894 (O_1894,N_19506,N_19527);
and UO_1895 (O_1895,N_19642,N_18372);
or UO_1896 (O_1896,N_18833,N_19666);
and UO_1897 (O_1897,N_19761,N_19131);
or UO_1898 (O_1898,N_18529,N_18808);
or UO_1899 (O_1899,N_18263,N_18206);
nand UO_1900 (O_1900,N_19140,N_18983);
xor UO_1901 (O_1901,N_19045,N_19142);
and UO_1902 (O_1902,N_18832,N_18593);
nand UO_1903 (O_1903,N_19122,N_19480);
nand UO_1904 (O_1904,N_18432,N_19065);
nor UO_1905 (O_1905,N_18087,N_19500);
xnor UO_1906 (O_1906,N_19652,N_19188);
nor UO_1907 (O_1907,N_18742,N_18912);
nor UO_1908 (O_1908,N_18855,N_19117);
xnor UO_1909 (O_1909,N_19089,N_19334);
xnor UO_1910 (O_1910,N_19598,N_18349);
nor UO_1911 (O_1911,N_19582,N_19021);
or UO_1912 (O_1912,N_19615,N_18492);
nor UO_1913 (O_1913,N_19592,N_19386);
and UO_1914 (O_1914,N_18144,N_19310);
nor UO_1915 (O_1915,N_19604,N_19543);
nand UO_1916 (O_1916,N_18526,N_19552);
nor UO_1917 (O_1917,N_19417,N_19244);
or UO_1918 (O_1918,N_18156,N_18514);
nor UO_1919 (O_1919,N_19549,N_18242);
nor UO_1920 (O_1920,N_18045,N_18306);
nand UO_1921 (O_1921,N_18981,N_18700);
and UO_1922 (O_1922,N_19435,N_19861);
and UO_1923 (O_1923,N_19515,N_18320);
nor UO_1924 (O_1924,N_18471,N_19602);
nand UO_1925 (O_1925,N_19040,N_19288);
or UO_1926 (O_1926,N_18960,N_18773);
nand UO_1927 (O_1927,N_19010,N_19011);
nor UO_1928 (O_1928,N_18273,N_18963);
and UO_1929 (O_1929,N_19271,N_19923);
nand UO_1930 (O_1930,N_19844,N_18066);
nor UO_1931 (O_1931,N_18410,N_18356);
and UO_1932 (O_1932,N_19579,N_19729);
nand UO_1933 (O_1933,N_18635,N_18802);
nand UO_1934 (O_1934,N_18718,N_18363);
nand UO_1935 (O_1935,N_18004,N_18189);
or UO_1936 (O_1936,N_18426,N_18201);
or UO_1937 (O_1937,N_19954,N_19125);
or UO_1938 (O_1938,N_19068,N_19855);
nand UO_1939 (O_1939,N_19433,N_18581);
xnor UO_1940 (O_1940,N_19327,N_19716);
nand UO_1941 (O_1941,N_19821,N_19231);
and UO_1942 (O_1942,N_19806,N_18365);
nand UO_1943 (O_1943,N_18640,N_18547);
and UO_1944 (O_1944,N_18990,N_19774);
xor UO_1945 (O_1945,N_18315,N_18291);
or UO_1946 (O_1946,N_19118,N_19744);
nor UO_1947 (O_1947,N_18215,N_18791);
or UO_1948 (O_1948,N_18037,N_18637);
xor UO_1949 (O_1949,N_18907,N_19975);
nand UO_1950 (O_1950,N_18260,N_19829);
nand UO_1951 (O_1951,N_19278,N_18107);
and UO_1952 (O_1952,N_18885,N_18647);
nor UO_1953 (O_1953,N_19956,N_18239);
nor UO_1954 (O_1954,N_18224,N_19598);
nor UO_1955 (O_1955,N_19243,N_19978);
nor UO_1956 (O_1956,N_18746,N_18901);
and UO_1957 (O_1957,N_19827,N_19777);
or UO_1958 (O_1958,N_19831,N_18207);
and UO_1959 (O_1959,N_18815,N_19289);
nand UO_1960 (O_1960,N_19033,N_18488);
nand UO_1961 (O_1961,N_18924,N_18922);
xor UO_1962 (O_1962,N_18455,N_19346);
or UO_1963 (O_1963,N_18999,N_19514);
and UO_1964 (O_1964,N_19244,N_18714);
nand UO_1965 (O_1965,N_18278,N_18715);
and UO_1966 (O_1966,N_18798,N_18143);
xnor UO_1967 (O_1967,N_19439,N_19397);
or UO_1968 (O_1968,N_18272,N_19886);
nand UO_1969 (O_1969,N_19253,N_19225);
nor UO_1970 (O_1970,N_18696,N_18592);
nand UO_1971 (O_1971,N_19739,N_18746);
or UO_1972 (O_1972,N_18298,N_19795);
nand UO_1973 (O_1973,N_19711,N_19815);
or UO_1974 (O_1974,N_19762,N_18848);
or UO_1975 (O_1975,N_19055,N_19904);
nand UO_1976 (O_1976,N_18320,N_19553);
nand UO_1977 (O_1977,N_18935,N_18327);
or UO_1978 (O_1978,N_19505,N_18447);
nor UO_1979 (O_1979,N_19651,N_18104);
or UO_1980 (O_1980,N_19552,N_19742);
or UO_1981 (O_1981,N_18054,N_18844);
nand UO_1982 (O_1982,N_19040,N_19118);
nor UO_1983 (O_1983,N_19367,N_18825);
nand UO_1984 (O_1984,N_18343,N_18222);
nand UO_1985 (O_1985,N_19035,N_19683);
xnor UO_1986 (O_1986,N_19915,N_18777);
and UO_1987 (O_1987,N_18429,N_18970);
and UO_1988 (O_1988,N_19916,N_18990);
and UO_1989 (O_1989,N_18853,N_18517);
nor UO_1990 (O_1990,N_19686,N_19799);
nor UO_1991 (O_1991,N_19423,N_18685);
or UO_1992 (O_1992,N_19203,N_19280);
or UO_1993 (O_1993,N_19491,N_19037);
and UO_1994 (O_1994,N_18842,N_19527);
and UO_1995 (O_1995,N_18267,N_19895);
and UO_1996 (O_1996,N_19037,N_19458);
nor UO_1997 (O_1997,N_18511,N_18764);
nor UO_1998 (O_1998,N_18809,N_18252);
nand UO_1999 (O_1999,N_19089,N_18785);
nand UO_2000 (O_2000,N_19038,N_19760);
and UO_2001 (O_2001,N_18877,N_18439);
or UO_2002 (O_2002,N_19831,N_18007);
or UO_2003 (O_2003,N_19931,N_19120);
xnor UO_2004 (O_2004,N_19026,N_18174);
or UO_2005 (O_2005,N_18972,N_18948);
or UO_2006 (O_2006,N_18201,N_18046);
and UO_2007 (O_2007,N_19162,N_18187);
xnor UO_2008 (O_2008,N_18324,N_19629);
xnor UO_2009 (O_2009,N_19392,N_19225);
and UO_2010 (O_2010,N_19745,N_18984);
nand UO_2011 (O_2011,N_18992,N_19810);
xor UO_2012 (O_2012,N_18616,N_18459);
or UO_2013 (O_2013,N_19505,N_19902);
nand UO_2014 (O_2014,N_18251,N_19396);
nand UO_2015 (O_2015,N_19276,N_18154);
or UO_2016 (O_2016,N_19603,N_19784);
nor UO_2017 (O_2017,N_18887,N_19237);
or UO_2018 (O_2018,N_19558,N_19526);
or UO_2019 (O_2019,N_19484,N_19289);
nor UO_2020 (O_2020,N_19395,N_18157);
and UO_2021 (O_2021,N_18006,N_19437);
or UO_2022 (O_2022,N_18022,N_19052);
or UO_2023 (O_2023,N_19951,N_18405);
or UO_2024 (O_2024,N_18175,N_18786);
nand UO_2025 (O_2025,N_18699,N_18971);
nor UO_2026 (O_2026,N_19469,N_19379);
nand UO_2027 (O_2027,N_19600,N_19131);
nand UO_2028 (O_2028,N_19346,N_19200);
and UO_2029 (O_2029,N_18624,N_18523);
xnor UO_2030 (O_2030,N_19187,N_19229);
nand UO_2031 (O_2031,N_19976,N_19169);
or UO_2032 (O_2032,N_19694,N_19108);
nor UO_2033 (O_2033,N_19088,N_18512);
nor UO_2034 (O_2034,N_19032,N_19677);
xnor UO_2035 (O_2035,N_18665,N_18839);
nand UO_2036 (O_2036,N_18702,N_18649);
or UO_2037 (O_2037,N_18251,N_19631);
nand UO_2038 (O_2038,N_18314,N_19703);
and UO_2039 (O_2039,N_19097,N_19505);
nand UO_2040 (O_2040,N_19080,N_18487);
and UO_2041 (O_2041,N_19884,N_18979);
nand UO_2042 (O_2042,N_18297,N_18138);
or UO_2043 (O_2043,N_18814,N_19663);
and UO_2044 (O_2044,N_18756,N_18757);
nand UO_2045 (O_2045,N_18982,N_19230);
nand UO_2046 (O_2046,N_19908,N_18613);
nand UO_2047 (O_2047,N_19318,N_19419);
or UO_2048 (O_2048,N_19620,N_18888);
or UO_2049 (O_2049,N_18784,N_19904);
xnor UO_2050 (O_2050,N_18794,N_19495);
nand UO_2051 (O_2051,N_19875,N_19672);
and UO_2052 (O_2052,N_19549,N_18514);
or UO_2053 (O_2053,N_19643,N_19662);
nand UO_2054 (O_2054,N_19133,N_18476);
and UO_2055 (O_2055,N_19661,N_18213);
xnor UO_2056 (O_2056,N_18072,N_18479);
nand UO_2057 (O_2057,N_18144,N_18127);
nand UO_2058 (O_2058,N_19865,N_19065);
or UO_2059 (O_2059,N_19412,N_18195);
nand UO_2060 (O_2060,N_19522,N_19123);
nor UO_2061 (O_2061,N_18204,N_19604);
nor UO_2062 (O_2062,N_19468,N_18412);
xnor UO_2063 (O_2063,N_19282,N_18326);
xor UO_2064 (O_2064,N_19937,N_18447);
or UO_2065 (O_2065,N_18626,N_19474);
nor UO_2066 (O_2066,N_18442,N_19588);
and UO_2067 (O_2067,N_19409,N_18917);
or UO_2068 (O_2068,N_18946,N_18895);
nor UO_2069 (O_2069,N_19723,N_19781);
nand UO_2070 (O_2070,N_18243,N_18108);
nor UO_2071 (O_2071,N_19344,N_19143);
nand UO_2072 (O_2072,N_19507,N_19518);
or UO_2073 (O_2073,N_18441,N_18159);
or UO_2074 (O_2074,N_18163,N_18445);
nor UO_2075 (O_2075,N_18331,N_19224);
or UO_2076 (O_2076,N_19772,N_19441);
nand UO_2077 (O_2077,N_19885,N_19253);
and UO_2078 (O_2078,N_19966,N_19797);
or UO_2079 (O_2079,N_19182,N_19557);
or UO_2080 (O_2080,N_19014,N_19654);
and UO_2081 (O_2081,N_19978,N_19765);
or UO_2082 (O_2082,N_18817,N_19349);
or UO_2083 (O_2083,N_18091,N_18211);
nor UO_2084 (O_2084,N_19871,N_18816);
nor UO_2085 (O_2085,N_19537,N_18130);
nand UO_2086 (O_2086,N_19387,N_18835);
nor UO_2087 (O_2087,N_19934,N_19943);
and UO_2088 (O_2088,N_19700,N_18725);
nand UO_2089 (O_2089,N_18954,N_18887);
xnor UO_2090 (O_2090,N_18969,N_18660);
and UO_2091 (O_2091,N_18213,N_19982);
nor UO_2092 (O_2092,N_18305,N_18857);
and UO_2093 (O_2093,N_18153,N_19444);
nand UO_2094 (O_2094,N_19898,N_19073);
nand UO_2095 (O_2095,N_19576,N_18785);
xor UO_2096 (O_2096,N_19488,N_18649);
and UO_2097 (O_2097,N_18642,N_18423);
nor UO_2098 (O_2098,N_19972,N_18756);
xor UO_2099 (O_2099,N_19156,N_19246);
nand UO_2100 (O_2100,N_18249,N_19931);
nor UO_2101 (O_2101,N_18990,N_18423);
or UO_2102 (O_2102,N_19842,N_19266);
nor UO_2103 (O_2103,N_18861,N_18730);
and UO_2104 (O_2104,N_18181,N_18994);
nand UO_2105 (O_2105,N_18518,N_19202);
nor UO_2106 (O_2106,N_19149,N_19164);
and UO_2107 (O_2107,N_18234,N_19126);
nand UO_2108 (O_2108,N_19471,N_19814);
or UO_2109 (O_2109,N_18377,N_18390);
and UO_2110 (O_2110,N_19774,N_19088);
and UO_2111 (O_2111,N_18103,N_18682);
and UO_2112 (O_2112,N_19137,N_19303);
nand UO_2113 (O_2113,N_18167,N_19133);
or UO_2114 (O_2114,N_18167,N_18283);
nand UO_2115 (O_2115,N_18585,N_19202);
nand UO_2116 (O_2116,N_19484,N_19100);
or UO_2117 (O_2117,N_18036,N_19966);
xnor UO_2118 (O_2118,N_19723,N_19577);
and UO_2119 (O_2119,N_18509,N_18255);
nand UO_2120 (O_2120,N_19938,N_18267);
xor UO_2121 (O_2121,N_19000,N_18645);
or UO_2122 (O_2122,N_18515,N_19744);
nand UO_2123 (O_2123,N_18866,N_18349);
nand UO_2124 (O_2124,N_19401,N_18384);
nand UO_2125 (O_2125,N_18785,N_19363);
xnor UO_2126 (O_2126,N_19857,N_18980);
nor UO_2127 (O_2127,N_19902,N_19343);
and UO_2128 (O_2128,N_18800,N_19842);
nand UO_2129 (O_2129,N_18998,N_18559);
or UO_2130 (O_2130,N_18670,N_19383);
nand UO_2131 (O_2131,N_18642,N_19374);
nor UO_2132 (O_2132,N_18310,N_19562);
and UO_2133 (O_2133,N_19477,N_18107);
and UO_2134 (O_2134,N_19182,N_18468);
or UO_2135 (O_2135,N_18105,N_18926);
nor UO_2136 (O_2136,N_19976,N_19319);
nand UO_2137 (O_2137,N_18801,N_18607);
nand UO_2138 (O_2138,N_19923,N_18380);
xnor UO_2139 (O_2139,N_18098,N_18940);
nand UO_2140 (O_2140,N_19919,N_19202);
or UO_2141 (O_2141,N_18247,N_18435);
nand UO_2142 (O_2142,N_18253,N_18233);
or UO_2143 (O_2143,N_19954,N_19491);
or UO_2144 (O_2144,N_19076,N_19170);
nand UO_2145 (O_2145,N_18086,N_19022);
or UO_2146 (O_2146,N_19306,N_19122);
and UO_2147 (O_2147,N_19111,N_18353);
xor UO_2148 (O_2148,N_19864,N_18125);
nand UO_2149 (O_2149,N_18193,N_18240);
or UO_2150 (O_2150,N_18895,N_19021);
and UO_2151 (O_2151,N_19491,N_19405);
or UO_2152 (O_2152,N_19511,N_18514);
nor UO_2153 (O_2153,N_18444,N_19695);
or UO_2154 (O_2154,N_18166,N_19139);
nand UO_2155 (O_2155,N_19817,N_18582);
xor UO_2156 (O_2156,N_19016,N_19917);
and UO_2157 (O_2157,N_18942,N_18747);
or UO_2158 (O_2158,N_18461,N_18449);
or UO_2159 (O_2159,N_18645,N_19235);
nor UO_2160 (O_2160,N_18392,N_18848);
and UO_2161 (O_2161,N_19037,N_19291);
or UO_2162 (O_2162,N_18247,N_19205);
nor UO_2163 (O_2163,N_19844,N_19272);
or UO_2164 (O_2164,N_19578,N_18289);
nand UO_2165 (O_2165,N_19640,N_18164);
and UO_2166 (O_2166,N_18621,N_19980);
nand UO_2167 (O_2167,N_19439,N_19758);
nand UO_2168 (O_2168,N_19485,N_18453);
or UO_2169 (O_2169,N_19826,N_19817);
and UO_2170 (O_2170,N_18823,N_18998);
nor UO_2171 (O_2171,N_18331,N_19544);
or UO_2172 (O_2172,N_19976,N_19387);
xor UO_2173 (O_2173,N_18112,N_18612);
and UO_2174 (O_2174,N_18946,N_19099);
and UO_2175 (O_2175,N_18946,N_19057);
nand UO_2176 (O_2176,N_18313,N_19093);
and UO_2177 (O_2177,N_18302,N_18299);
nor UO_2178 (O_2178,N_18786,N_18238);
and UO_2179 (O_2179,N_18842,N_18327);
and UO_2180 (O_2180,N_18999,N_19032);
nand UO_2181 (O_2181,N_18462,N_19436);
or UO_2182 (O_2182,N_18111,N_18561);
and UO_2183 (O_2183,N_19170,N_19849);
nand UO_2184 (O_2184,N_18180,N_18342);
and UO_2185 (O_2185,N_18359,N_18901);
nor UO_2186 (O_2186,N_19090,N_18798);
nand UO_2187 (O_2187,N_18982,N_18076);
nor UO_2188 (O_2188,N_18197,N_18644);
and UO_2189 (O_2189,N_18550,N_19630);
nand UO_2190 (O_2190,N_19470,N_19019);
nor UO_2191 (O_2191,N_18566,N_19623);
xor UO_2192 (O_2192,N_18173,N_19789);
xnor UO_2193 (O_2193,N_19877,N_18728);
nor UO_2194 (O_2194,N_18942,N_19869);
nor UO_2195 (O_2195,N_18146,N_18016);
nand UO_2196 (O_2196,N_18095,N_19612);
nor UO_2197 (O_2197,N_19911,N_19767);
or UO_2198 (O_2198,N_19738,N_19439);
and UO_2199 (O_2199,N_19937,N_19419);
nor UO_2200 (O_2200,N_19555,N_19527);
nor UO_2201 (O_2201,N_18150,N_19660);
or UO_2202 (O_2202,N_19748,N_19348);
nor UO_2203 (O_2203,N_18528,N_19519);
or UO_2204 (O_2204,N_19201,N_19752);
nor UO_2205 (O_2205,N_19331,N_18600);
or UO_2206 (O_2206,N_19228,N_18944);
and UO_2207 (O_2207,N_18807,N_18429);
nand UO_2208 (O_2208,N_19981,N_18269);
nor UO_2209 (O_2209,N_19382,N_19247);
nor UO_2210 (O_2210,N_18103,N_18785);
nand UO_2211 (O_2211,N_18514,N_19525);
and UO_2212 (O_2212,N_19177,N_18585);
and UO_2213 (O_2213,N_18684,N_18437);
and UO_2214 (O_2214,N_18491,N_19777);
nand UO_2215 (O_2215,N_18229,N_19895);
nor UO_2216 (O_2216,N_18488,N_19653);
and UO_2217 (O_2217,N_18355,N_18495);
nor UO_2218 (O_2218,N_18094,N_18385);
nand UO_2219 (O_2219,N_19968,N_18293);
xnor UO_2220 (O_2220,N_19822,N_19346);
and UO_2221 (O_2221,N_19800,N_18083);
or UO_2222 (O_2222,N_19003,N_18591);
nand UO_2223 (O_2223,N_18008,N_19193);
or UO_2224 (O_2224,N_19958,N_18564);
and UO_2225 (O_2225,N_18121,N_18893);
nor UO_2226 (O_2226,N_18403,N_19363);
nor UO_2227 (O_2227,N_18847,N_18890);
or UO_2228 (O_2228,N_19082,N_19020);
nor UO_2229 (O_2229,N_18558,N_19105);
xor UO_2230 (O_2230,N_18334,N_18539);
and UO_2231 (O_2231,N_18632,N_19671);
nor UO_2232 (O_2232,N_19995,N_18891);
nor UO_2233 (O_2233,N_19279,N_19787);
nand UO_2234 (O_2234,N_19886,N_18561);
or UO_2235 (O_2235,N_19666,N_19676);
nor UO_2236 (O_2236,N_19976,N_19858);
nand UO_2237 (O_2237,N_18231,N_19620);
and UO_2238 (O_2238,N_18330,N_19600);
and UO_2239 (O_2239,N_19422,N_19938);
or UO_2240 (O_2240,N_19743,N_19501);
and UO_2241 (O_2241,N_19753,N_18028);
or UO_2242 (O_2242,N_18820,N_19514);
and UO_2243 (O_2243,N_18056,N_18847);
nand UO_2244 (O_2244,N_19560,N_19246);
or UO_2245 (O_2245,N_18776,N_18978);
nand UO_2246 (O_2246,N_19933,N_19913);
xnor UO_2247 (O_2247,N_19842,N_18110);
or UO_2248 (O_2248,N_19662,N_18777);
or UO_2249 (O_2249,N_19682,N_18681);
nor UO_2250 (O_2250,N_19404,N_19402);
and UO_2251 (O_2251,N_19092,N_18089);
xor UO_2252 (O_2252,N_18142,N_18310);
or UO_2253 (O_2253,N_18164,N_19770);
nand UO_2254 (O_2254,N_18180,N_19261);
nor UO_2255 (O_2255,N_18176,N_19605);
xnor UO_2256 (O_2256,N_18456,N_18850);
nand UO_2257 (O_2257,N_18411,N_19377);
nand UO_2258 (O_2258,N_18119,N_19260);
and UO_2259 (O_2259,N_19776,N_18953);
nor UO_2260 (O_2260,N_18667,N_18778);
nor UO_2261 (O_2261,N_19850,N_18037);
nand UO_2262 (O_2262,N_18579,N_19185);
nand UO_2263 (O_2263,N_19084,N_18404);
nor UO_2264 (O_2264,N_19224,N_19859);
or UO_2265 (O_2265,N_19384,N_19083);
nand UO_2266 (O_2266,N_18768,N_19535);
or UO_2267 (O_2267,N_19643,N_18343);
or UO_2268 (O_2268,N_19118,N_19565);
and UO_2269 (O_2269,N_18184,N_19022);
xor UO_2270 (O_2270,N_19364,N_18709);
nand UO_2271 (O_2271,N_19057,N_19381);
or UO_2272 (O_2272,N_19928,N_19418);
nand UO_2273 (O_2273,N_19201,N_18358);
nand UO_2274 (O_2274,N_18337,N_18138);
or UO_2275 (O_2275,N_18690,N_19298);
nor UO_2276 (O_2276,N_18104,N_19242);
nand UO_2277 (O_2277,N_19633,N_18086);
or UO_2278 (O_2278,N_19323,N_19468);
and UO_2279 (O_2279,N_19098,N_18496);
nor UO_2280 (O_2280,N_18403,N_18970);
xnor UO_2281 (O_2281,N_18176,N_19946);
and UO_2282 (O_2282,N_19918,N_18386);
or UO_2283 (O_2283,N_18128,N_19063);
nor UO_2284 (O_2284,N_18312,N_19952);
nor UO_2285 (O_2285,N_19625,N_18076);
nand UO_2286 (O_2286,N_18106,N_18939);
nand UO_2287 (O_2287,N_18965,N_18468);
nand UO_2288 (O_2288,N_18772,N_18585);
nor UO_2289 (O_2289,N_19916,N_19379);
nor UO_2290 (O_2290,N_18483,N_19000);
or UO_2291 (O_2291,N_19926,N_19539);
or UO_2292 (O_2292,N_19339,N_18774);
and UO_2293 (O_2293,N_18888,N_18399);
and UO_2294 (O_2294,N_19340,N_18457);
and UO_2295 (O_2295,N_18129,N_18472);
and UO_2296 (O_2296,N_19233,N_18292);
nor UO_2297 (O_2297,N_18891,N_19010);
nand UO_2298 (O_2298,N_18064,N_18940);
nor UO_2299 (O_2299,N_18352,N_19554);
or UO_2300 (O_2300,N_19080,N_18499);
nand UO_2301 (O_2301,N_19774,N_19856);
xor UO_2302 (O_2302,N_18263,N_18542);
or UO_2303 (O_2303,N_19954,N_19130);
nand UO_2304 (O_2304,N_19967,N_19719);
xnor UO_2305 (O_2305,N_18447,N_19626);
or UO_2306 (O_2306,N_19145,N_19767);
and UO_2307 (O_2307,N_19284,N_19905);
nor UO_2308 (O_2308,N_18372,N_19236);
or UO_2309 (O_2309,N_19211,N_19151);
nand UO_2310 (O_2310,N_18612,N_18343);
and UO_2311 (O_2311,N_18499,N_19177);
nand UO_2312 (O_2312,N_18369,N_19632);
or UO_2313 (O_2313,N_18064,N_18411);
nor UO_2314 (O_2314,N_18425,N_19635);
nor UO_2315 (O_2315,N_19158,N_19666);
and UO_2316 (O_2316,N_19238,N_18258);
and UO_2317 (O_2317,N_19494,N_18808);
nand UO_2318 (O_2318,N_18106,N_18880);
nor UO_2319 (O_2319,N_18185,N_18997);
nor UO_2320 (O_2320,N_19034,N_18393);
xor UO_2321 (O_2321,N_18571,N_18935);
or UO_2322 (O_2322,N_18685,N_19553);
nand UO_2323 (O_2323,N_19269,N_18942);
nand UO_2324 (O_2324,N_18956,N_18499);
nand UO_2325 (O_2325,N_18083,N_19980);
and UO_2326 (O_2326,N_18667,N_19407);
xnor UO_2327 (O_2327,N_18150,N_19134);
or UO_2328 (O_2328,N_19761,N_19695);
and UO_2329 (O_2329,N_19139,N_19586);
nor UO_2330 (O_2330,N_18661,N_19567);
or UO_2331 (O_2331,N_18643,N_19289);
and UO_2332 (O_2332,N_18171,N_18785);
and UO_2333 (O_2333,N_18861,N_19742);
xor UO_2334 (O_2334,N_19008,N_19298);
nand UO_2335 (O_2335,N_18250,N_19675);
or UO_2336 (O_2336,N_18557,N_19935);
and UO_2337 (O_2337,N_18538,N_18720);
nor UO_2338 (O_2338,N_19691,N_18247);
nor UO_2339 (O_2339,N_19878,N_19131);
xnor UO_2340 (O_2340,N_19761,N_18531);
nand UO_2341 (O_2341,N_19845,N_19887);
and UO_2342 (O_2342,N_18355,N_18249);
or UO_2343 (O_2343,N_18365,N_19040);
and UO_2344 (O_2344,N_19276,N_19280);
nor UO_2345 (O_2345,N_18574,N_18329);
nor UO_2346 (O_2346,N_19946,N_18709);
nor UO_2347 (O_2347,N_19891,N_18258);
and UO_2348 (O_2348,N_18041,N_19616);
nand UO_2349 (O_2349,N_18096,N_18380);
xnor UO_2350 (O_2350,N_19987,N_18397);
nor UO_2351 (O_2351,N_19926,N_19963);
xor UO_2352 (O_2352,N_19650,N_19623);
or UO_2353 (O_2353,N_19324,N_19223);
or UO_2354 (O_2354,N_18914,N_19081);
or UO_2355 (O_2355,N_19168,N_19970);
nand UO_2356 (O_2356,N_18735,N_18870);
nand UO_2357 (O_2357,N_18312,N_18637);
nor UO_2358 (O_2358,N_18890,N_19669);
or UO_2359 (O_2359,N_19690,N_18764);
or UO_2360 (O_2360,N_19275,N_19072);
nand UO_2361 (O_2361,N_18000,N_19402);
nor UO_2362 (O_2362,N_19262,N_19316);
and UO_2363 (O_2363,N_19961,N_19299);
or UO_2364 (O_2364,N_18459,N_18917);
nor UO_2365 (O_2365,N_18767,N_19217);
xnor UO_2366 (O_2366,N_18461,N_19409);
nand UO_2367 (O_2367,N_18724,N_19040);
xnor UO_2368 (O_2368,N_19891,N_19423);
or UO_2369 (O_2369,N_18419,N_18609);
and UO_2370 (O_2370,N_18248,N_18266);
or UO_2371 (O_2371,N_18808,N_19321);
and UO_2372 (O_2372,N_19264,N_19554);
or UO_2373 (O_2373,N_18537,N_19175);
nor UO_2374 (O_2374,N_18117,N_19025);
xor UO_2375 (O_2375,N_18917,N_19465);
or UO_2376 (O_2376,N_18943,N_19488);
nand UO_2377 (O_2377,N_18747,N_18301);
or UO_2378 (O_2378,N_19461,N_18919);
xnor UO_2379 (O_2379,N_19763,N_18165);
xnor UO_2380 (O_2380,N_19256,N_18496);
nor UO_2381 (O_2381,N_19976,N_19437);
and UO_2382 (O_2382,N_19028,N_19687);
nor UO_2383 (O_2383,N_18357,N_18538);
nor UO_2384 (O_2384,N_19771,N_19397);
xnor UO_2385 (O_2385,N_18602,N_18279);
nor UO_2386 (O_2386,N_19681,N_19325);
and UO_2387 (O_2387,N_18874,N_18358);
or UO_2388 (O_2388,N_18762,N_18002);
xor UO_2389 (O_2389,N_19701,N_18909);
nand UO_2390 (O_2390,N_19578,N_19878);
nor UO_2391 (O_2391,N_19872,N_19643);
or UO_2392 (O_2392,N_18039,N_19181);
nand UO_2393 (O_2393,N_18849,N_19600);
or UO_2394 (O_2394,N_18893,N_19211);
and UO_2395 (O_2395,N_18556,N_19502);
or UO_2396 (O_2396,N_18392,N_19496);
nand UO_2397 (O_2397,N_18517,N_19021);
or UO_2398 (O_2398,N_19430,N_19448);
nor UO_2399 (O_2399,N_18199,N_19269);
or UO_2400 (O_2400,N_18468,N_18872);
xnor UO_2401 (O_2401,N_18601,N_18248);
nand UO_2402 (O_2402,N_19160,N_19328);
and UO_2403 (O_2403,N_19130,N_18938);
nor UO_2404 (O_2404,N_19877,N_19119);
nor UO_2405 (O_2405,N_19488,N_18701);
or UO_2406 (O_2406,N_19058,N_19646);
nor UO_2407 (O_2407,N_19616,N_18836);
nand UO_2408 (O_2408,N_18364,N_19870);
xor UO_2409 (O_2409,N_18979,N_19965);
nor UO_2410 (O_2410,N_18606,N_18996);
xor UO_2411 (O_2411,N_19613,N_18948);
or UO_2412 (O_2412,N_19460,N_19474);
xnor UO_2413 (O_2413,N_18974,N_18803);
nor UO_2414 (O_2414,N_18988,N_18846);
and UO_2415 (O_2415,N_18553,N_18083);
and UO_2416 (O_2416,N_18624,N_18063);
nand UO_2417 (O_2417,N_18718,N_19855);
nor UO_2418 (O_2418,N_19305,N_19463);
or UO_2419 (O_2419,N_19079,N_19747);
xor UO_2420 (O_2420,N_18069,N_19135);
nand UO_2421 (O_2421,N_18466,N_18733);
or UO_2422 (O_2422,N_18688,N_18297);
or UO_2423 (O_2423,N_18433,N_19892);
and UO_2424 (O_2424,N_19999,N_19972);
and UO_2425 (O_2425,N_18413,N_18336);
xor UO_2426 (O_2426,N_19728,N_18805);
nand UO_2427 (O_2427,N_18819,N_19024);
or UO_2428 (O_2428,N_18192,N_19388);
nor UO_2429 (O_2429,N_18092,N_18149);
xor UO_2430 (O_2430,N_19172,N_19648);
nand UO_2431 (O_2431,N_18340,N_18684);
nor UO_2432 (O_2432,N_19851,N_19025);
nand UO_2433 (O_2433,N_18216,N_19967);
and UO_2434 (O_2434,N_18445,N_18150);
and UO_2435 (O_2435,N_19614,N_19292);
and UO_2436 (O_2436,N_18891,N_18080);
nand UO_2437 (O_2437,N_18907,N_18774);
nand UO_2438 (O_2438,N_19710,N_19820);
nor UO_2439 (O_2439,N_19796,N_19991);
xor UO_2440 (O_2440,N_19796,N_19102);
xor UO_2441 (O_2441,N_19273,N_19464);
nor UO_2442 (O_2442,N_18407,N_19586);
and UO_2443 (O_2443,N_18217,N_18256);
and UO_2444 (O_2444,N_19811,N_19500);
and UO_2445 (O_2445,N_19379,N_18776);
nor UO_2446 (O_2446,N_18029,N_19188);
nor UO_2447 (O_2447,N_19910,N_18052);
nand UO_2448 (O_2448,N_18356,N_19187);
or UO_2449 (O_2449,N_18033,N_19172);
and UO_2450 (O_2450,N_19853,N_19643);
nor UO_2451 (O_2451,N_19177,N_18623);
xnor UO_2452 (O_2452,N_18124,N_18244);
nor UO_2453 (O_2453,N_19424,N_19969);
or UO_2454 (O_2454,N_18673,N_19153);
or UO_2455 (O_2455,N_19519,N_19683);
nor UO_2456 (O_2456,N_19226,N_19097);
nand UO_2457 (O_2457,N_18157,N_18314);
xnor UO_2458 (O_2458,N_18902,N_18293);
and UO_2459 (O_2459,N_18445,N_19162);
and UO_2460 (O_2460,N_19210,N_18286);
nand UO_2461 (O_2461,N_19052,N_18688);
and UO_2462 (O_2462,N_19507,N_19651);
and UO_2463 (O_2463,N_19315,N_19609);
or UO_2464 (O_2464,N_19654,N_18985);
nand UO_2465 (O_2465,N_18388,N_19388);
nand UO_2466 (O_2466,N_18525,N_18392);
and UO_2467 (O_2467,N_18686,N_18028);
nor UO_2468 (O_2468,N_19223,N_18803);
or UO_2469 (O_2469,N_18230,N_18821);
nor UO_2470 (O_2470,N_18907,N_18629);
or UO_2471 (O_2471,N_18455,N_19825);
xor UO_2472 (O_2472,N_18125,N_19414);
and UO_2473 (O_2473,N_19034,N_18565);
nand UO_2474 (O_2474,N_18783,N_18802);
and UO_2475 (O_2475,N_19431,N_19214);
or UO_2476 (O_2476,N_19639,N_18150);
xor UO_2477 (O_2477,N_19229,N_19270);
nand UO_2478 (O_2478,N_19884,N_19374);
and UO_2479 (O_2479,N_18481,N_18906);
nor UO_2480 (O_2480,N_19106,N_19637);
nand UO_2481 (O_2481,N_18085,N_19837);
and UO_2482 (O_2482,N_18435,N_19532);
nor UO_2483 (O_2483,N_19166,N_19096);
nor UO_2484 (O_2484,N_19417,N_18661);
nor UO_2485 (O_2485,N_19979,N_19975);
or UO_2486 (O_2486,N_18209,N_18343);
or UO_2487 (O_2487,N_18128,N_18206);
or UO_2488 (O_2488,N_19807,N_19900);
or UO_2489 (O_2489,N_19814,N_18260);
and UO_2490 (O_2490,N_18052,N_18388);
nor UO_2491 (O_2491,N_18743,N_18527);
nor UO_2492 (O_2492,N_18163,N_18356);
nand UO_2493 (O_2493,N_18357,N_19290);
nand UO_2494 (O_2494,N_19858,N_18552);
and UO_2495 (O_2495,N_19878,N_19247);
or UO_2496 (O_2496,N_19355,N_18533);
nor UO_2497 (O_2497,N_19533,N_19262);
nand UO_2498 (O_2498,N_18904,N_19943);
and UO_2499 (O_2499,N_18677,N_19123);
endmodule