module basic_3000_30000_3500_6_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_143,In_1986);
or U1 (N_1,In_2993,In_1599);
or U2 (N_2,In_2893,In_2674);
nand U3 (N_3,In_2482,In_2684);
or U4 (N_4,In_2611,In_2169);
nand U5 (N_5,In_2422,In_2954);
xor U6 (N_6,In_1027,In_276);
or U7 (N_7,In_1265,In_263);
and U8 (N_8,In_596,In_2093);
nor U9 (N_9,In_1271,In_858);
nor U10 (N_10,In_2428,In_2170);
and U11 (N_11,In_2449,In_1054);
and U12 (N_12,In_1138,In_1245);
or U13 (N_13,In_364,In_701);
or U14 (N_14,In_1284,In_1009);
nor U15 (N_15,In_525,In_2889);
xor U16 (N_16,In_1725,In_422);
xor U17 (N_17,In_726,In_2410);
nand U18 (N_18,In_2007,In_308);
and U19 (N_19,In_2155,In_1662);
and U20 (N_20,In_1189,In_1329);
and U21 (N_21,In_2388,In_524);
and U22 (N_22,In_1642,In_1434);
nor U23 (N_23,In_1942,In_341);
nand U24 (N_24,In_1678,In_13);
or U25 (N_25,In_666,In_1626);
nand U26 (N_26,In_786,In_2631);
and U27 (N_27,In_2650,In_1338);
nor U28 (N_28,In_1336,In_1476);
or U29 (N_29,In_80,In_744);
nand U30 (N_30,In_380,In_476);
nand U31 (N_31,In_2283,In_1891);
or U32 (N_32,In_386,In_2799);
and U33 (N_33,In_1342,In_1471);
or U34 (N_34,In_1282,In_248);
nor U35 (N_35,In_2721,In_2232);
xnor U36 (N_36,In_1323,In_874);
xor U37 (N_37,In_384,In_401);
nand U38 (N_38,In_1967,In_256);
nand U39 (N_39,In_2301,In_2393);
xnor U40 (N_40,In_2182,In_1635);
and U41 (N_41,In_1077,In_618);
xor U42 (N_42,In_678,In_1168);
and U43 (N_43,In_2369,In_1739);
xnor U44 (N_44,In_1477,In_2264);
nor U45 (N_45,In_2885,In_2425);
xor U46 (N_46,In_1359,In_354);
xor U47 (N_47,In_120,In_1107);
and U48 (N_48,In_2612,In_1930);
nand U49 (N_49,In_2198,In_432);
xor U50 (N_50,In_351,In_1534);
xor U51 (N_51,In_1079,In_2278);
and U52 (N_52,In_2959,In_128);
nor U53 (N_53,In_792,In_1367);
and U54 (N_54,In_2836,In_1877);
nand U55 (N_55,In_2065,In_2277);
xor U56 (N_56,In_54,In_2978);
nor U57 (N_57,In_1208,In_2246);
xnor U58 (N_58,In_684,In_1497);
nand U59 (N_59,In_2771,In_1718);
or U60 (N_60,In_1893,In_544);
or U61 (N_61,In_514,In_134);
and U62 (N_62,In_379,In_2759);
and U63 (N_63,In_702,In_1822);
nand U64 (N_64,In_2082,In_250);
or U65 (N_65,In_1597,In_1907);
and U66 (N_66,In_1745,In_557);
nand U67 (N_67,In_1064,In_2298);
nand U68 (N_68,In_1920,In_1843);
nand U69 (N_69,In_2568,In_862);
nand U70 (N_70,In_615,In_1674);
nand U71 (N_71,In_1663,In_2347);
or U72 (N_72,In_267,In_2116);
nand U73 (N_73,In_2874,In_1790);
nand U74 (N_74,In_1896,In_721);
nand U75 (N_75,In_1428,In_901);
nand U76 (N_76,In_1972,In_2451);
xnor U77 (N_77,In_1254,In_581);
and U78 (N_78,In_444,In_1179);
xor U79 (N_79,In_753,In_1902);
xnor U80 (N_80,In_1393,In_2747);
or U81 (N_81,In_1129,In_1363);
nand U82 (N_82,In_783,In_1550);
nor U83 (N_83,In_2215,In_1037);
xnor U84 (N_84,In_1389,In_472);
nor U85 (N_85,In_2560,In_1078);
nor U86 (N_86,In_1517,In_2900);
and U87 (N_87,In_2976,In_1086);
nand U88 (N_88,In_1622,In_2312);
xnor U89 (N_89,In_961,In_2296);
or U90 (N_90,In_712,In_489);
nand U91 (N_91,In_1101,In_808);
nor U92 (N_92,In_1303,In_2702);
nor U93 (N_93,In_2273,In_1708);
nand U94 (N_94,In_907,In_685);
nor U95 (N_95,In_1144,In_183);
nor U96 (N_96,In_2104,In_1031);
or U97 (N_97,In_225,In_945);
or U98 (N_98,In_2980,In_1895);
xor U99 (N_99,In_2250,In_919);
or U100 (N_100,In_1785,In_2546);
nand U101 (N_101,In_1696,In_1257);
and U102 (N_102,In_2829,In_2647);
xor U103 (N_103,In_1536,In_621);
and U104 (N_104,In_1001,In_2081);
xor U105 (N_105,In_1084,In_583);
xor U106 (N_106,In_2257,In_1108);
xnor U107 (N_107,In_1447,In_2816);
and U108 (N_108,In_2964,In_1201);
or U109 (N_109,In_1118,In_601);
and U110 (N_110,In_2586,In_1504);
xor U111 (N_111,In_1924,In_879);
or U112 (N_112,In_2107,In_2968);
and U113 (N_113,In_1210,In_922);
xor U114 (N_114,In_1430,In_2772);
and U115 (N_115,In_193,In_2991);
or U116 (N_116,In_2371,In_2032);
and U117 (N_117,In_793,In_2497);
or U118 (N_118,In_1897,In_960);
nor U119 (N_119,In_2746,In_90);
nor U120 (N_120,In_2117,In_2585);
nor U121 (N_121,In_1308,In_146);
nor U122 (N_122,In_2867,In_587);
xor U123 (N_123,In_1005,In_2092);
nand U124 (N_124,In_1246,In_280);
nand U125 (N_125,In_287,In_719);
and U126 (N_126,In_2963,In_403);
xnor U127 (N_127,In_1831,In_2915);
and U128 (N_128,In_2554,In_2691);
nor U129 (N_129,In_638,In_2779);
and U130 (N_130,In_2988,In_1780);
or U131 (N_131,In_2583,In_2110);
nor U132 (N_132,In_25,In_1844);
and U133 (N_133,In_2005,In_2628);
or U134 (N_134,In_2433,In_1703);
and U135 (N_135,In_2548,In_156);
or U136 (N_136,In_979,In_2706);
and U137 (N_137,In_1668,In_478);
nand U138 (N_138,In_2933,In_2488);
xnor U139 (N_139,In_2059,In_967);
and U140 (N_140,In_71,In_2290);
or U141 (N_141,In_1651,In_2417);
xnor U142 (N_142,In_1029,In_1861);
xnor U143 (N_143,In_400,In_437);
or U144 (N_144,In_2525,In_2971);
nor U145 (N_145,In_1773,In_1518);
and U146 (N_146,In_1052,In_1111);
and U147 (N_147,In_1012,In_2552);
nand U148 (N_148,In_2,In_1180);
and U149 (N_149,In_1561,In_2673);
or U150 (N_150,In_2641,In_409);
nor U151 (N_151,In_2941,In_532);
or U152 (N_152,In_5,In_2756);
nand U153 (N_153,In_2187,In_1253);
xnor U154 (N_154,In_1485,In_2330);
xor U155 (N_155,In_307,In_606);
or U156 (N_156,In_485,In_16);
nand U157 (N_157,In_2837,In_2821);
or U158 (N_158,In_595,In_1914);
and U159 (N_159,In_2467,In_445);
or U160 (N_160,In_2513,In_1821);
xor U161 (N_161,In_1787,In_645);
and U162 (N_162,In_681,In_2138);
nor U163 (N_163,In_2131,In_515);
and U164 (N_164,In_2492,In_1598);
nor U165 (N_165,In_1579,In_980);
nor U166 (N_166,In_1681,In_229);
and U167 (N_167,In_1417,In_1243);
and U168 (N_168,In_1815,In_772);
xor U169 (N_169,In_2502,In_1713);
nor U170 (N_170,In_1612,In_2135);
xor U171 (N_171,In_95,In_2935);
or U172 (N_172,In_2851,In_1949);
nor U173 (N_173,In_1131,In_1295);
nor U174 (N_174,In_1824,In_1370);
and U175 (N_175,In_2532,In_2094);
nand U176 (N_176,In_1071,In_2887);
or U177 (N_177,In_112,In_1124);
nor U178 (N_178,In_1484,In_1595);
nand U179 (N_179,In_1742,In_2768);
or U180 (N_180,In_1605,In_2656);
nand U181 (N_181,In_2056,In_872);
xor U182 (N_182,In_2389,In_1938);
xor U183 (N_183,In_2106,In_2563);
nor U184 (N_184,In_881,In_2786);
and U185 (N_185,In_2953,In_2260);
or U186 (N_186,In_210,In_2668);
nand U187 (N_187,In_1957,In_1412);
or U188 (N_188,In_1672,In_531);
xnor U189 (N_189,In_1456,In_2326);
and U190 (N_190,In_1887,In_619);
nand U191 (N_191,In_41,In_851);
or U192 (N_192,In_1796,In_318);
xnor U193 (N_193,In_886,In_2681);
or U194 (N_194,In_1998,In_2778);
or U195 (N_195,In_1817,In_1617);
and U196 (N_196,In_2929,In_818);
nor U197 (N_197,In_39,In_836);
and U198 (N_198,In_878,In_2237);
nor U199 (N_199,In_1454,In_711);
or U200 (N_200,In_197,In_668);
xor U201 (N_201,In_1919,In_1867);
and U202 (N_202,In_260,In_2152);
or U203 (N_203,In_1377,In_2919);
or U204 (N_204,In_623,In_1686);
nor U205 (N_205,In_501,In_92);
or U206 (N_206,In_1994,In_1307);
nand U207 (N_207,In_1842,In_240);
and U208 (N_208,In_413,In_2648);
nor U209 (N_209,In_2434,In_2649);
xor U210 (N_210,In_1406,In_10);
and U211 (N_211,In_1305,In_325);
or U212 (N_212,In_2033,In_1234);
nor U213 (N_213,In_426,In_174);
nand U214 (N_214,In_129,In_56);
or U215 (N_215,In_513,In_117);
or U216 (N_216,In_329,In_125);
and U217 (N_217,In_2419,In_1446);
xnor U218 (N_218,In_870,In_2420);
nand U219 (N_219,In_368,In_1298);
nand U220 (N_220,In_2536,In_1343);
or U221 (N_221,In_2604,In_1231);
and U222 (N_222,In_1464,In_297);
nand U223 (N_223,In_843,In_1847);
or U224 (N_224,In_2391,In_288);
and U225 (N_225,In_1571,In_2950);
and U226 (N_226,In_2374,In_264);
and U227 (N_227,In_1075,In_2342);
nand U228 (N_228,In_2233,In_1218);
nor U229 (N_229,In_1576,In_194);
and U230 (N_230,In_434,In_2698);
or U231 (N_231,In_254,In_2561);
xnor U232 (N_232,In_419,In_1378);
xnor U233 (N_233,In_1051,In_1206);
xnor U234 (N_234,In_937,In_1699);
nor U235 (N_235,In_1838,In_2584);
and U236 (N_236,In_2564,In_1682);
nor U237 (N_237,In_1149,In_2745);
nand U238 (N_238,In_1969,In_2809);
and U239 (N_239,In_40,In_2876);
nor U240 (N_240,In_1399,In_24);
nor U241 (N_241,In_160,In_2992);
xor U242 (N_242,In_1007,In_326);
xnor U243 (N_243,In_1392,In_2784);
or U244 (N_244,In_184,In_633);
nand U245 (N_245,In_2735,In_1448);
nor U246 (N_246,In_69,In_1373);
nor U247 (N_247,In_588,In_2080);
nand U248 (N_248,In_337,In_1185);
and U249 (N_249,In_454,In_1368);
and U250 (N_250,In_2239,In_1755);
nand U251 (N_251,In_2173,In_138);
nand U252 (N_252,In_2426,In_2589);
or U253 (N_253,In_2531,In_372);
and U254 (N_254,In_1496,In_1936);
nor U255 (N_255,In_6,In_2710);
nor U256 (N_256,In_2366,In_825);
nor U257 (N_257,In_739,In_199);
xnor U258 (N_258,In_2234,In_1082);
and U259 (N_259,In_1886,In_776);
nand U260 (N_260,In_2742,In_2118);
xor U261 (N_261,In_1687,In_1870);
nand U262 (N_262,In_1570,In_2252);
or U263 (N_263,In_1322,In_2060);
or U264 (N_264,In_630,In_96);
nand U265 (N_265,In_1935,In_867);
nand U266 (N_266,In_1053,In_765);
xor U267 (N_267,In_1016,In_584);
nand U268 (N_268,In_2195,In_2466);
or U269 (N_269,In_833,In_1981);
or U270 (N_270,In_677,In_2798);
and U271 (N_271,In_2639,In_2986);
nand U272 (N_272,In_1350,In_698);
or U273 (N_273,In_1801,In_130);
or U274 (N_274,In_294,In_1292);
xnor U275 (N_275,In_2794,In_1833);
nand U276 (N_276,In_2248,In_2856);
and U277 (N_277,In_187,In_1724);
and U278 (N_278,In_154,In_1784);
xnor U279 (N_279,In_1814,In_1743);
and U280 (N_280,In_2275,In_2593);
and U281 (N_281,In_1973,In_756);
nand U282 (N_282,In_889,In_847);
or U283 (N_283,In_1038,In_1993);
nand U284 (N_284,In_1069,In_2063);
nor U285 (N_285,In_535,In_1911);
nor U286 (N_286,In_849,In_2154);
or U287 (N_287,In_652,In_468);
nor U288 (N_288,In_2960,In_2379);
nor U289 (N_289,In_2262,In_2207);
nand U290 (N_290,In_1553,In_757);
xnor U291 (N_291,In_1564,In_2453);
or U292 (N_292,In_2670,In_2375);
nand U293 (N_293,In_2902,In_2640);
nor U294 (N_294,In_854,In_2361);
xor U295 (N_295,In_1148,In_2223);
nor U296 (N_296,In_722,In_2643);
nor U297 (N_297,In_163,In_2946);
xor U298 (N_298,In_1530,In_281);
nand U299 (N_299,In_2834,In_2334);
and U300 (N_300,In_1424,In_2089);
nand U301 (N_301,In_2962,In_1065);
xor U302 (N_302,In_1033,In_597);
or U303 (N_303,In_2027,In_1106);
nor U304 (N_304,In_568,In_1278);
or U305 (N_305,In_1804,In_2003);
or U306 (N_306,In_141,In_2922);
nand U307 (N_307,In_2981,In_1638);
xnor U308 (N_308,In_21,In_2000);
nor U309 (N_309,In_2675,In_1503);
or U310 (N_310,In_1892,In_305);
xnor U311 (N_311,In_1590,In_1491);
xnor U312 (N_312,In_2061,In_1791);
xor U313 (N_313,In_1238,In_1629);
nor U314 (N_314,In_2789,In_2731);
nor U315 (N_315,In_605,In_607);
nor U316 (N_316,In_2622,In_1960);
or U317 (N_317,In_2454,In_2945);
nand U318 (N_318,In_2679,In_1963);
nand U319 (N_319,In_933,In_344);
nand U320 (N_320,In_111,In_797);
nand U321 (N_321,In_1156,In_1019);
nor U322 (N_322,In_1056,In_119);
xor U323 (N_323,In_1618,In_74);
nand U324 (N_324,In_799,In_2229);
nor U325 (N_325,In_529,In_1432);
nor U326 (N_326,In_2814,In_1976);
nor U327 (N_327,In_827,In_1970);
and U328 (N_328,In_2338,In_830);
or U329 (N_329,In_1829,In_2261);
nand U330 (N_330,In_763,In_1975);
and U331 (N_331,In_2225,In_1992);
nand U332 (N_332,In_392,In_1355);
or U333 (N_333,In_1685,In_2174);
or U334 (N_334,In_2443,In_1722);
xnor U335 (N_335,In_1566,In_1905);
nor U336 (N_336,In_2490,In_1912);
and U337 (N_337,In_1750,In_1020);
and U338 (N_338,In_2997,In_1068);
xor U339 (N_339,In_2214,In_834);
or U340 (N_340,In_731,In_2284);
nand U341 (N_341,In_2509,In_1311);
xor U342 (N_342,In_133,In_244);
nor U343 (N_343,In_2787,In_2409);
and U344 (N_344,In_1091,In_1883);
xnor U345 (N_345,In_752,In_78);
xor U346 (N_346,In_2692,In_1939);
xnor U347 (N_347,In_494,In_1145);
xor U348 (N_348,In_2925,In_2730);
nand U349 (N_349,In_2791,In_1630);
nand U350 (N_350,In_1803,In_784);
nand U351 (N_351,In_1737,In_207);
nor U352 (N_352,In_1182,In_1580);
or U353 (N_353,In_1772,In_2448);
xnor U354 (N_354,In_1439,In_1495);
or U355 (N_355,In_227,In_569);
or U356 (N_356,In_2455,In_2271);
nor U357 (N_357,In_2528,In_304);
or U358 (N_358,In_2069,In_905);
and U359 (N_359,In_1244,In_469);
nor U360 (N_360,In_1481,In_1139);
or U361 (N_361,In_1213,In_1903);
nor U362 (N_362,In_279,In_104);
nand U363 (N_363,In_2242,In_1586);
nand U364 (N_364,In_1711,In_309);
nor U365 (N_365,In_692,In_34);
and U366 (N_366,In_123,In_1562);
xor U367 (N_367,In_2411,In_2358);
xnor U368 (N_368,In_2311,In_1006);
or U369 (N_369,In_2635,In_2952);
or U370 (N_370,In_2857,In_2947);
xnor U371 (N_371,In_819,In_640);
nand U372 (N_372,In_795,In_1247);
nor U373 (N_373,In_769,In_550);
and U374 (N_374,In_1289,In_2892);
nor U375 (N_375,In_2217,In_2603);
nor U376 (N_376,In_1807,In_2325);
or U377 (N_377,In_2119,In_1362);
xor U378 (N_378,In_211,In_2587);
xor U379 (N_379,In_462,In_2295);
or U380 (N_380,In_759,In_271);
nand U381 (N_381,In_1693,In_2468);
xnor U382 (N_382,In_2018,In_598);
and U383 (N_383,In_2370,In_2045);
nor U384 (N_384,In_2767,In_1411);
nor U385 (N_385,In_1493,In_2352);
nor U386 (N_386,In_1050,In_2833);
and U387 (N_387,In_2123,In_1395);
nand U388 (N_388,In_2348,In_972);
or U389 (N_389,In_209,In_1061);
and U390 (N_390,In_777,In_779);
nor U391 (N_391,In_2253,In_1863);
xnor U392 (N_392,In_2321,In_2943);
and U393 (N_393,In_2303,In_2363);
nor U394 (N_394,In_1030,In_147);
nor U395 (N_395,In_26,In_1782);
xnor U396 (N_396,In_450,In_913);
xor U397 (N_397,In_2510,In_932);
xor U398 (N_398,In_620,In_1354);
xor U399 (N_399,In_941,In_1418);
and U400 (N_400,In_2073,In_1151);
xor U401 (N_401,In_2588,In_706);
or U402 (N_402,In_36,In_452);
or U403 (N_403,In_106,In_665);
nand U404 (N_404,In_393,In_1057);
and U405 (N_405,In_2686,In_1172);
or U406 (N_406,In_230,In_578);
or U407 (N_407,In_2499,In_1953);
nand U408 (N_408,In_2773,In_1537);
and U409 (N_409,In_1190,In_2581);
nand U410 (N_410,In_2208,In_821);
nand U411 (N_411,In_1134,In_1966);
or U412 (N_412,In_464,In_2359);
nand U413 (N_413,In_1300,In_1003);
or U414 (N_414,In_667,In_993);
or U415 (N_415,In_773,In_949);
and U416 (N_416,In_1394,In_1717);
nand U417 (N_417,In_1494,In_1955);
or U418 (N_418,In_1256,In_1684);
nor U419 (N_419,In_1081,In_2383);
nor U420 (N_420,In_1070,In_567);
and U421 (N_421,In_1800,In_971);
nand U422 (N_422,In_1375,In_1024);
and U423 (N_423,In_824,In_2481);
xor U424 (N_424,In_2346,In_1459);
or U425 (N_425,In_1632,In_2013);
nand U426 (N_426,In_1192,In_1540);
or U427 (N_427,In_2267,In_1239);
xor U428 (N_428,In_2895,In_1734);
nor U429 (N_429,In_2543,In_912);
xor U430 (N_430,In_1525,In_212);
xnor U431 (N_431,In_1689,In_284);
or U432 (N_432,In_2351,In_2539);
and U433 (N_433,In_2412,In_1132);
or U434 (N_434,In_2500,In_1716);
or U435 (N_435,In_2636,In_2637);
nor U436 (N_436,In_2595,In_2245);
xnor U437 (N_437,In_802,In_429);
nor U438 (N_438,In_2785,In_998);
nor U439 (N_439,In_1288,In_1653);
nand U440 (N_440,In_1022,In_277);
and U441 (N_441,In_2875,In_840);
xnor U442 (N_442,In_2004,In_1733);
nand U443 (N_443,In_1974,In_2827);
nand U444 (N_444,In_2313,In_2802);
xor U445 (N_445,In_2697,In_2218);
nand U446 (N_446,In_2219,In_1162);
and U447 (N_447,In_2011,In_1285);
nor U448 (N_448,In_2803,In_237);
nor U449 (N_449,In_365,In_2699);
nand U450 (N_450,In_1552,In_302);
and U451 (N_451,In_298,In_576);
xor U452 (N_452,In_2621,In_660);
nand U453 (N_453,In_1607,In_1871);
or U454 (N_454,In_2987,In_2396);
xor U455 (N_455,In_2306,In_746);
xor U456 (N_456,In_837,In_149);
xor U457 (N_457,In_2105,In_2285);
nand U458 (N_458,In_1062,In_2146);
or U459 (N_459,In_1879,In_2645);
nor U460 (N_460,In_1868,In_1263);
or U461 (N_461,In_2906,In_807);
and U462 (N_462,In_1788,In_87);
or U463 (N_463,In_1478,In_735);
and U464 (N_464,In_2353,In_1421);
xor U465 (N_465,In_860,In_1296);
and U466 (N_466,In_2038,In_2682);
nand U467 (N_467,In_1425,In_688);
nor U468 (N_468,In_2101,In_2416);
nor U469 (N_469,In_2537,In_2270);
nor U470 (N_470,In_1461,In_604);
or U471 (N_471,In_1140,In_547);
xor U472 (N_472,In_512,In_1698);
nand U473 (N_473,In_369,In_755);
xor U474 (N_474,In_334,In_2855);
or U475 (N_475,In_1209,In_2203);
or U476 (N_476,In_2797,In_911);
nor U477 (N_477,In_2506,In_1876);
xor U478 (N_478,In_2286,In_2776);
nor U479 (N_479,In_290,In_2415);
or U480 (N_480,In_2211,In_608);
and U481 (N_481,In_1215,In_2620);
nor U482 (N_482,In_2888,In_1273);
nand U483 (N_483,In_2614,In_1812);
nor U484 (N_484,In_1109,In_2990);
nand U485 (N_485,In_2164,In_1982);
nor U486 (N_486,In_1453,In_2852);
nand U487 (N_487,In_651,In_1827);
nor U488 (N_488,In_1175,In_2818);
nor U489 (N_489,In_1979,In_460);
xor U490 (N_490,In_1319,In_1252);
xor U491 (N_491,In_2144,In_2293);
and U492 (N_492,In_1123,In_1055);
nor U493 (N_493,In_2826,In_2464);
nand U494 (N_494,In_2258,In_1968);
nor U495 (N_495,In_1715,In_2255);
xnor U496 (N_496,In_497,In_1694);
and U497 (N_497,In_2542,In_1881);
xnor U498 (N_498,In_1152,In_2324);
xnor U499 (N_499,In_299,In_536);
and U500 (N_500,In_2349,In_1014);
xnor U501 (N_501,In_1444,In_1904);
nand U502 (N_502,In_1313,In_1501);
nand U503 (N_503,In_2220,In_2512);
xnor U504 (N_504,In_394,In_543);
or U505 (N_505,In_984,In_1726);
nor U506 (N_506,In_2367,In_2801);
nand U507 (N_507,In_2951,In_609);
nand U508 (N_508,In_1223,In_2427);
or U509 (N_509,In_1908,In_2127);
nand U510 (N_510,In_1203,In_1173);
nand U511 (N_511,In_1872,In_540);
xor U512 (N_512,In_1945,In_1783);
and U513 (N_513,In_1648,In_2457);
nand U514 (N_514,In_2569,In_314);
xor U515 (N_515,In_91,In_2143);
xnor U516 (N_516,In_274,In_545);
or U517 (N_517,In_891,In_383);
xor U518 (N_518,In_316,In_1269);
xor U519 (N_519,In_2088,In_813);
nand U520 (N_520,In_816,In_1660);
or U521 (N_521,In_969,In_602);
nand U522 (N_522,In_1588,In_2533);
xor U523 (N_523,In_1353,In_357);
or U524 (N_524,In_1858,In_213);
and U525 (N_525,In_1971,In_2165);
or U526 (N_526,In_2758,In_2613);
and U527 (N_527,In_148,In_1039);
and U528 (N_528,In_1828,In_1352);
or U529 (N_529,In_1126,In_2084);
and U530 (N_530,In_1087,In_953);
nor U531 (N_531,In_978,In_2103);
or U532 (N_532,In_1183,In_136);
and U533 (N_533,In_50,In_2734);
xor U534 (N_534,In_2133,In_1775);
and U535 (N_535,In_990,In_336);
xnor U536 (N_536,In_1122,In_2753);
xor U537 (N_537,In_2024,In_100);
xnor U538 (N_538,In_2824,In_2266);
nor U539 (N_539,In_2209,In_79);
xnor U540 (N_540,In_1422,In_656);
nor U541 (N_541,In_1864,In_1249);
and U542 (N_542,In_1513,In_2590);
and U543 (N_543,In_2337,In_1529);
xor U544 (N_544,In_7,In_2177);
nor U545 (N_545,In_1042,In_345);
xor U546 (N_546,In_644,In_1695);
xnor U547 (N_547,In_155,In_2197);
nor U548 (N_548,In_2654,In_323);
xnor U549 (N_549,In_1382,In_1554);
nor U550 (N_550,In_1002,In_1608);
nor U551 (N_551,In_1542,In_1511);
nor U552 (N_552,In_58,In_1736);
and U553 (N_553,In_1977,In_1627);
or U554 (N_554,In_1700,In_315);
xnor U555 (N_555,In_2810,In_324);
nor U556 (N_556,In_2297,In_2870);
or U557 (N_557,In_1339,In_2701);
nand U558 (N_558,In_1654,In_1926);
or U559 (N_559,In_1702,In_2397);
nor U560 (N_560,In_2871,In_1187);
nand U561 (N_561,In_1806,In_500);
nor U562 (N_562,In_2651,In_1846);
nor U563 (N_563,In_1752,In_2905);
and U564 (N_564,In_1468,In_2486);
nand U565 (N_565,In_884,In_689);
xnor U566 (N_566,In_2766,In_2861);
nor U567 (N_567,In_750,In_2469);
and U568 (N_568,In_533,In_1596);
nand U569 (N_569,In_2700,In_2134);
and U570 (N_570,In_2901,In_2849);
and U571 (N_571,In_1522,In_114);
or U572 (N_572,In_553,In_203);
nand U573 (N_573,In_246,In_1749);
and U574 (N_574,In_2578,In_272);
and U575 (N_575,In_865,In_1741);
xnor U576 (N_576,In_632,In_9);
nor U577 (N_577,In_2471,In_2148);
nand U578 (N_578,In_558,In_1415);
or U579 (N_579,In_1344,In_1345);
xor U580 (N_580,In_1809,In_671);
nor U581 (N_581,In_2037,In_1366);
and U582 (N_582,In_831,In_2339);
xor U583 (N_583,In_2357,In_1349);
nor U584 (N_584,In_2664,In_1125);
or U585 (N_585,In_389,In_2881);
nor U586 (N_586,In_2141,In_1202);
and U587 (N_587,In_2811,In_1952);
or U588 (N_588,In_538,In_164);
or U589 (N_589,In_2908,In_1856);
nor U590 (N_590,In_1874,In_2846);
and U591 (N_591,In_740,In_2377);
or U592 (N_592,In_275,In_1291);
nor U593 (N_593,In_2831,In_1933);
or U594 (N_594,In_1441,In_1194);
or U595 (N_595,In_699,In_2014);
nor U596 (N_596,In_407,In_1241);
or U597 (N_597,In_2708,In_950);
nor U598 (N_598,In_2764,In_42);
nand U599 (N_599,In_734,In_2869);
or U600 (N_600,In_1221,In_2555);
xnor U601 (N_601,In_2452,In_1516);
xnor U602 (N_602,In_2688,In_1925);
nand U603 (N_603,In_1890,In_1306);
and U604 (N_604,In_1317,In_648);
xnor U605 (N_605,In_2049,In_1777);
or U606 (N_606,In_812,In_231);
xor U607 (N_607,In_1121,In_98);
xnor U608 (N_608,In_1442,In_2596);
xor U609 (N_609,In_457,In_1793);
xor U610 (N_610,In_2392,In_340);
and U611 (N_611,In_1665,In_467);
or U612 (N_612,In_2320,In_2178);
or U613 (N_613,In_343,In_2395);
and U614 (N_614,In_218,In_977);
nand U615 (N_615,In_1677,In_2292);
or U616 (N_616,In_2210,In_2083);
nor U617 (N_617,In_2387,In_2384);
nor U618 (N_618,In_770,In_2001);
nor U619 (N_619,In_2345,In_2329);
or U620 (N_620,In_1443,In_803);
nor U621 (N_621,In_1414,In_853);
and U622 (N_622,In_1230,In_1514);
or U623 (N_623,In_1620,In_390);
nor U624 (N_624,In_1059,In_996);
and U625 (N_625,In_245,In_815);
nor U626 (N_626,In_2400,In_2189);
nand U627 (N_627,In_2168,In_1859);
and U628 (N_628,In_2473,In_347);
nand U629 (N_629,In_2461,In_2519);
xor U630 (N_630,In_319,In_131);
nor U631 (N_631,In_1889,In_1102);
or U632 (N_632,In_931,In_360);
or U633 (N_633,In_2115,In_1774);
and U634 (N_634,In_1191,In_2385);
nor U635 (N_635,In_2336,In_1384);
and U636 (N_636,In_1470,In_2690);
and U637 (N_637,In_1035,In_1171);
nor U638 (N_638,In_2254,In_2970);
nor U639 (N_639,In_1232,In_1880);
and U640 (N_640,In_2432,In_817);
nor U641 (N_641,In_1917,In_381);
and U642 (N_642,In_842,In_1652);
nor U643 (N_643,In_892,In_1819);
and U644 (N_644,In_1862,In_1707);
nor U645 (N_645,In_2331,In_1929);
xnor U646 (N_646,In_105,In_2414);
or U647 (N_647,In_1766,In_747);
nand U648 (N_648,In_762,In_2256);
xnor U649 (N_649,In_508,In_2047);
or U650 (N_650,In_2465,In_2494);
nor U651 (N_651,In_68,In_1021);
xnor U652 (N_652,In_2557,In_890);
xnor U653 (N_653,In_2230,In_859);
nor U654 (N_654,In_47,In_1017);
and U655 (N_655,In_966,In_2937);
xnor U656 (N_656,In_1810,In_989);
nand U657 (N_657,In_2288,In_2090);
nor U658 (N_658,In_1947,In_423);
or U659 (N_659,In_1985,In_2711);
nor U660 (N_660,In_1163,In_1427);
or U661 (N_661,In_659,In_2983);
nor U662 (N_662,In_253,In_12);
nand U663 (N_663,In_1199,In_1593);
and U664 (N_664,In_2156,In_2407);
nor U665 (N_665,In_661,In_2068);
nor U666 (N_666,In_1198,In_2194);
and U667 (N_667,In_868,In_374);
and U668 (N_668,In_258,In_1710);
nor U669 (N_669,In_2850,In_1110);
xor U670 (N_670,In_1839,In_1820);
nand U671 (N_671,In_952,In_848);
xor U672 (N_672,In_1402,In_1299);
xor U673 (N_673,In_2276,In_723);
and U674 (N_674,In_814,In_1747);
or U675 (N_675,In_2709,In_2860);
or U676 (N_676,In_1740,In_355);
or U677 (N_677,In_2501,In_2485);
nand U678 (N_678,In_2025,In_2793);
or U679 (N_679,In_574,In_774);
or U680 (N_680,In_441,In_805);
or U681 (N_681,In_2316,In_83);
and U682 (N_682,In_1980,In_1761);
nor U683 (N_683,In_1997,In_2973);
nand U684 (N_684,In_2795,In_2862);
or U685 (N_685,In_81,In_1837);
or U686 (N_686,In_625,In_2279);
or U687 (N_687,In_1096,In_674);
nor U688 (N_688,In_906,In_1645);
xnor U689 (N_689,In_2835,In_2130);
nor U690 (N_690,In_1888,In_456);
xnor U691 (N_691,In_2677,In_2848);
or U692 (N_692,In_2841,In_242);
and U693 (N_693,In_252,In_2010);
and U694 (N_694,In_733,In_1851);
and U695 (N_695,In_863,In_590);
nor U696 (N_696,In_1331,In_612);
nand U697 (N_697,In_1950,In_2522);
nor U698 (N_698,In_943,In_479);
nand U699 (N_699,In_591,In_301);
nand U700 (N_700,In_742,In_506);
or U701 (N_701,In_17,In_534);
or U702 (N_702,In_73,In_480);
nor U703 (N_703,In_1048,In_788);
nand U704 (N_704,In_103,In_1176);
or U705 (N_705,In_766,In_2097);
or U706 (N_706,In_2315,In_169);
or U707 (N_707,In_958,In_1878);
xnor U708 (N_708,In_646,In_2865);
nor U709 (N_709,In_519,In_2920);
nor U710 (N_710,In_2023,In_2854);
nor U711 (N_711,In_1834,In_431);
or U712 (N_712,In_1991,In_2044);
nand U713 (N_713,In_1532,In_2491);
or U714 (N_714,In_1600,In_1099);
or U715 (N_715,In_2939,In_1396);
nor U716 (N_716,In_503,In_1988);
and U717 (N_717,In_2565,In_2880);
nor U718 (N_718,In_2122,In_1808);
xor U719 (N_719,In_387,In_322);
and U720 (N_720,In_2226,In_2240);
nand U721 (N_721,In_975,In_176);
nor U722 (N_722,In_1527,In_771);
or U723 (N_723,In_142,In_708);
and U724 (N_724,In_1623,In_2399);
and U725 (N_725,In_2029,In_703);
or U726 (N_726,In_973,In_1885);
and U727 (N_727,In_2300,In_2549);
nor U728 (N_728,In_2401,In_397);
or U729 (N_729,In_1130,In_1429);
nand U730 (N_730,In_1509,In_1135);
nor U731 (N_731,In_1435,In_527);
nand U732 (N_732,In_161,In_2944);
and U733 (N_733,In_15,In_1076);
or U734 (N_734,In_66,In_1410);
nor U735 (N_735,In_1340,In_22);
nand U736 (N_736,In_158,In_1114);
nand U737 (N_737,In_2489,In_201);
or U738 (N_738,In_2936,In_938);
or U739 (N_739,In_934,In_636);
nand U740 (N_740,In_2932,In_2440);
xor U741 (N_741,In_2221,In_2805);
nor U742 (N_742,In_628,In_1267);
or U743 (N_743,In_624,In_2496);
nor U744 (N_744,In_1523,In_2601);
xor U745 (N_745,In_165,In_1697);
nor U746 (N_746,In_1921,In_2040);
nor U747 (N_747,In_2012,In_1763);
nand U748 (N_748,In_492,In_616);
nor U749 (N_749,In_2227,In_992);
xor U750 (N_750,In_1753,In_1222);
xor U751 (N_751,In_1692,In_124);
nand U752 (N_752,In_2333,In_985);
and U753 (N_753,In_86,In_1433);
and U754 (N_754,In_570,In_2354);
or U755 (N_755,In_241,In_2483);
or U756 (N_756,In_613,In_2934);
or U757 (N_757,In_221,In_416);
nand U758 (N_758,In_2404,In_614);
or U759 (N_759,In_964,In_1852);
nand U760 (N_760,In_2518,In_1128);
xnor U761 (N_761,In_1512,In_180);
nand U762 (N_762,In_2739,In_1419);
nor U763 (N_763,In_1840,In_1089);
nor U764 (N_764,In_2355,In_2535);
nor U765 (N_765,In_243,In_2918);
or U766 (N_766,In_2072,In_2599);
or U767 (N_767,In_2205,In_170);
nor U768 (N_768,In_518,In_2281);
xor U769 (N_769,In_1541,In_2703);
or U770 (N_770,In_709,In_2322);
and U771 (N_771,In_367,In_2626);
nor U772 (N_772,In_1732,In_2580);
xnor U773 (N_773,In_2160,In_2180);
and U774 (N_774,In_72,In_2036);
or U775 (N_775,In_361,In_2696);
nand U776 (N_776,In_436,In_2150);
or U777 (N_777,In_1909,In_1910);
or U778 (N_778,In_555,In_1758);
and U779 (N_779,In_1631,In_48);
and U780 (N_780,In_2884,In_226);
or U781 (N_781,In_806,In_101);
xor U782 (N_782,In_2538,In_713);
xor U783 (N_783,In_303,In_2890);
and U784 (N_784,In_2547,In_171);
nor U785 (N_785,In_1964,In_186);
nor U786 (N_786,In_801,In_887);
nand U787 (N_787,In_846,In_2924);
xor U788 (N_788,In_1592,In_1);
xnor U789 (N_789,In_940,In_1644);
nand U790 (N_790,In_561,In_477);
nor U791 (N_791,In_2942,In_1487);
and U792 (N_792,In_552,In_2238);
nor U793 (N_793,In_2598,In_2607);
nor U794 (N_794,In_1049,In_2605);
nor U795 (N_795,In_2408,In_593);
nor U796 (N_796,In_110,In_1407);
and U797 (N_797,In_2820,In_1073);
nor U798 (N_798,In_1990,In_55);
nand U799 (N_799,In_113,In_2031);
or U800 (N_800,In_2762,In_791);
or U801 (N_801,In_883,In_2204);
nand U802 (N_802,In_2897,In_1473);
or U803 (N_803,In_2931,In_1259);
or U804 (N_804,In_321,In_2940);
nand U805 (N_805,In_310,In_1236);
nor U806 (N_806,In_1304,In_175);
and U807 (N_807,In_2062,In_2441);
xnor U808 (N_808,In_546,In_1538);
nor U809 (N_809,In_2558,In_1364);
and U810 (N_810,In_2479,In_2685);
and U811 (N_811,In_1334,In_2576);
xor U812 (N_812,In_2938,In_238);
nand U813 (N_813,In_438,In_398);
and U814 (N_814,In_2825,In_2228);
nor U815 (N_815,In_2308,In_2423);
xnor U816 (N_816,In_395,In_424);
or U817 (N_817,In_2026,In_2577);
nor U818 (N_818,In_1701,In_1460);
nor U819 (N_819,In_1549,In_269);
nand U820 (N_820,In_2048,In_1941);
or U821 (N_821,In_1455,In_2843);
nor U822 (N_822,In_2602,In_433);
xnor U823 (N_823,In_2317,In_1764);
and U824 (N_824,In_179,In_826);
xnor U825 (N_825,In_1835,In_2592);
and U826 (N_826,In_459,In_880);
and U827 (N_827,In_331,In_1594);
xor U828 (N_828,In_944,In_592);
nor U829 (N_829,In_2200,In_330);
nand U830 (N_830,In_1142,In_2175);
and U831 (N_831,In_1146,In_2176);
nand U832 (N_832,In_2002,In_1611);
or U833 (N_833,In_700,In_947);
or U834 (N_834,In_2616,In_278);
and U835 (N_835,In_718,In_2186);
nand U836 (N_836,In_1526,In_2961);
nand U837 (N_837,In_1869,In_1400);
and U838 (N_838,In_2800,In_2913);
nand U839 (N_839,In_2495,In_673);
xnor U840 (N_840,In_178,In_694);
and U841 (N_841,In_2161,In_2078);
xor U842 (N_842,In_417,In_517);
nand U843 (N_843,In_2665,In_2043);
nand U844 (N_844,In_2761,In_1776);
and U845 (N_845,In_370,In_2365);
nand U846 (N_846,In_781,In_1195);
xor U847 (N_847,In_1274,In_1388);
nand U848 (N_848,In_2715,In_1312);
or U849 (N_849,In_844,In_2188);
and U850 (N_850,In_2571,In_1255);
xnor U851 (N_851,In_610,In_2879);
and U852 (N_852,In_2373,In_2424);
nor U853 (N_853,In_220,In_962);
nand U854 (N_854,In_728,In_440);
and U855 (N_855,In_1272,In_839);
nor U856 (N_856,In_1898,In_232);
nor U857 (N_857,In_575,In_1769);
xnor U858 (N_858,In_2694,In_838);
or U859 (N_859,In_122,In_994);
and U860 (N_860,In_2368,In_1679);
or U861 (N_861,In_49,In_629);
and U862 (N_862,In_2095,In_888);
or U863 (N_863,In_2524,In_2859);
nand U864 (N_864,In_1560,In_1664);
xor U865 (N_865,In_1301,In_2749);
or U866 (N_866,In_2566,In_2140);
xor U867 (N_867,In_1823,In_2085);
and U868 (N_868,In_2630,In_2927);
or U869 (N_869,In_296,In_228);
nand U870 (N_870,In_2019,In_976);
nor U871 (N_871,In_1018,In_939);
nand U872 (N_872,In_2840,In_151);
xnor U873 (N_873,In_1572,In_1141);
or U874 (N_874,In_1634,In_1639);
nand U875 (N_875,In_2975,In_2398);
or U876 (N_876,In_687,In_1376);
xnor U877 (N_877,In_273,In_19);
xnor U878 (N_878,In_2725,In_2574);
and U879 (N_879,In_317,In_2022);
nand U880 (N_880,In_1591,In_473);
and U881 (N_881,In_1452,In_2907);
nor U882 (N_882,In_1161,In_67);
nand U883 (N_883,In_1845,In_2435);
and U884 (N_884,In_391,In_2100);
nor U885 (N_885,In_716,In_2294);
xnor U886 (N_886,In_1333,In_2274);
nor U887 (N_887,In_177,In_1046);
nor U888 (N_888,In_481,In_2792);
nor U889 (N_889,In_1060,In_2926);
or U890 (N_890,In_453,In_1738);
nand U891 (N_891,In_2327,In_1490);
and U892 (N_892,In_1899,In_2808);
nand U893 (N_893,In_116,In_2193);
nand U894 (N_894,In_2224,In_929);
nor U895 (N_895,In_402,In_2600);
and U896 (N_896,In_52,In_77);
nor U897 (N_897,In_809,In_2845);
nand U898 (N_898,In_1219,In_224);
xor U899 (N_899,In_2573,In_2579);
or U900 (N_900,In_850,In_1436);
nand U901 (N_901,In_1094,In_1405);
xnor U902 (N_902,In_2693,In_1507);
and U903 (N_903,In_30,In_873);
and U904 (N_904,In_335,In_1258);
or U905 (N_905,In_1104,In_921);
or U906 (N_906,In_2163,In_63);
nor U907 (N_907,In_1403,In_2493);
nor U908 (N_908,In_2185,In_463);
and U909 (N_909,In_2015,In_562);
and U910 (N_910,In_2567,In_2087);
xor U911 (N_911,In_1381,In_474);
or U912 (N_912,In_31,In_2319);
and U913 (N_913,In_2074,In_2340);
xnor U914 (N_914,In_2832,In_782);
nand U915 (N_915,In_1445,In_62);
or U916 (N_916,In_2508,In_1583);
or U917 (N_917,In_2477,In_2462);
and U918 (N_918,In_1066,In_1900);
and U919 (N_919,In_20,In_1721);
nor U920 (N_920,In_109,In_2891);
xor U921 (N_921,In_51,In_2842);
nor U922 (N_922,In_895,In_107);
xor U923 (N_923,In_1356,In_504);
nand U924 (N_924,In_172,In_2111);
or U925 (N_925,In_778,In_1603);
or U926 (N_926,In_2247,In_1347);
xnor U927 (N_927,In_600,In_2191);
nand U928 (N_928,In_1587,In_2125);
or U929 (N_929,In_2179,In_2545);
nor U930 (N_930,In_1999,In_1423);
nand U931 (N_931,In_2719,In_2658);
or U932 (N_932,In_268,In_363);
and U933 (N_933,In_1647,In_585);
or U934 (N_934,In_1137,In_871);
nand U935 (N_935,In_2623,In_137);
nor U936 (N_936,In_1637,In_1276);
and U937 (N_937,In_856,In_2153);
or U938 (N_938,In_732,In_1853);
nor U939 (N_939,In_1937,In_2521);
or U940 (N_940,In_2886,In_2956);
and U941 (N_941,In_559,In_2763);
nor U942 (N_942,In_2807,In_657);
or U943 (N_943,In_1416,In_523);
or U944 (N_944,In_1948,In_93);
nand U945 (N_945,In_153,In_754);
nand U946 (N_946,In_1535,In_1266);
or U947 (N_947,In_2982,In_1420);
nand U948 (N_948,In_1646,In_1667);
or U949 (N_949,In_1413,In_1556);
and U950 (N_950,In_421,In_2460);
nor U951 (N_951,In_265,In_1321);
xnor U952 (N_952,In_2183,In_430);
and U953 (N_953,In_1619,In_126);
nor U954 (N_954,In_2644,In_1013);
nand U955 (N_955,In_1324,In_2741);
or U956 (N_956,In_2738,In_261);
nand U957 (N_957,In_1440,In_1242);
or U958 (N_958,In_751,In_2847);
nor U959 (N_959,In_1458,In_1602);
nor U960 (N_960,In_1943,In_490);
nand U961 (N_961,In_1480,In_2661);
nand U962 (N_962,In_1770,In_1882);
nand U963 (N_963,In_2475,In_311);
nand U964 (N_964,In_2657,In_1781);
and U965 (N_965,In_1719,In_1211);
or U966 (N_966,In_1335,In_925);
nor U967 (N_967,In_1989,In_663);
nor U968 (N_968,In_2609,In_2655);
and U969 (N_969,In_157,In_121);
and U970 (N_970,In_676,In_470);
nor U971 (N_971,In_76,In_1916);
nor U972 (N_972,In_537,In_1860);
or U973 (N_973,In_1727,In_1524);
or U974 (N_974,In_2222,In_2145);
and U975 (N_975,In_948,In_852);
xor U976 (N_976,In_1577,In_639);
xnor U977 (N_977,In_1797,In_1640);
xor U978 (N_978,In_686,In_511);
and U979 (N_979,In_145,In_1928);
nand U980 (N_980,In_1962,In_611);
nand U981 (N_981,In_2732,In_150);
or U982 (N_982,In_2765,In_2403);
xor U983 (N_983,In_449,In_2431);
nand U984 (N_984,In_1063,In_2894);
and U985 (N_985,In_2137,In_1283);
and U986 (N_986,In_1260,In_375);
xnor U987 (N_987,In_841,In_1792);
nand U988 (N_988,In_2394,In_1160);
xor U989 (N_989,In_2124,In_461);
or U990 (N_990,In_1227,In_1044);
or U991 (N_991,In_893,In_987);
nor U992 (N_992,In_2863,In_1510);
nor U993 (N_993,In_291,In_2541);
nor U994 (N_994,In_882,In_2877);
or U995 (N_995,In_915,In_2804);
or U996 (N_996,In_1216,In_2627);
and U997 (N_997,In_1351,In_1723);
nor U998 (N_998,In_1978,In_1836);
nor U999 (N_999,In_572,In_691);
nor U1000 (N_1000,In_1996,In_510);
xor U1001 (N_1001,In_1825,In_1636);
nor U1002 (N_1002,In_2202,In_579);
nor U1003 (N_1003,In_1705,In_1028);
nand U1004 (N_1004,In_2966,In_2064);
or U1005 (N_1005,In_499,In_1116);
xor U1006 (N_1006,In_970,In_448);
nand U1007 (N_1007,In_2206,In_196);
xor U1008 (N_1008,In_900,In_2171);
nand U1009 (N_1009,In_215,In_2139);
nor U1010 (N_1010,In_1369,In_1167);
nor U1011 (N_1011,In_554,In_2268);
and U1012 (N_1012,In_1371,In_439);
or U1013 (N_1013,In_1671,In_496);
or U1014 (N_1014,In_2343,In_1372);
or U1015 (N_1015,In_1922,In_2903);
or U1016 (N_1016,In_295,In_857);
and U1017 (N_1017,In_1113,In_2591);
xnor U1018 (N_1018,In_904,In_516);
nand U1019 (N_1019,In_1609,In_1760);
xor U1020 (N_1020,In_2476,In_2683);
and U1021 (N_1021,In_2653,In_2783);
and U1022 (N_1022,In_2498,In_577);
and U1023 (N_1023,In_2916,In_2444);
and U1024 (N_1024,In_675,In_2705);
or U1025 (N_1025,In_1262,In_563);
or U1026 (N_1026,In_1628,In_486);
and U1027 (N_1027,In_97,In_658);
nor U1028 (N_1028,In_484,In_724);
or U1029 (N_1029,In_2760,In_1728);
xor U1030 (N_1030,In_2305,In_564);
nor U1031 (N_1031,In_2967,In_1251);
or U1032 (N_1032,In_1505,In_1196);
xor U1033 (N_1033,In_1676,In_234);
nor U1034 (N_1034,In_1894,In_1043);
xnor U1035 (N_1035,In_2291,In_1169);
nand U1036 (N_1036,In_1565,In_715);
and U1037 (N_1037,In_2830,In_2899);
nand U1038 (N_1038,In_346,In_910);
or U1039 (N_1039,In_2487,In_2838);
or U1040 (N_1040,In_2718,In_2615);
xnor U1041 (N_1041,In_1515,In_2430);
xnor U1042 (N_1042,In_2091,In_1004);
xnor U1043 (N_1043,In_152,In_59);
or U1044 (N_1044,In_968,In_1212);
or U1045 (N_1045,In_1673,In_1984);
xnor U1046 (N_1046,In_1466,In_1100);
nand U1047 (N_1047,In_1469,In_560);
and U1048 (N_1048,In_2474,In_2516);
or U1049 (N_1049,In_353,In_2021);
nor U1050 (N_1050,In_412,In_1794);
xnor U1051 (N_1051,In_2328,In_1621);
and U1052 (N_1052,In_957,In_2780);
xor U1053 (N_1053,In_217,In_2041);
xor U1054 (N_1054,In_2520,In_1080);
nor U1055 (N_1055,In_682,In_565);
xnor U1056 (N_1056,In_594,In_166);
or U1057 (N_1057,In_2666,In_1154);
nand U1058 (N_1058,In_2617,In_866);
and U1059 (N_1059,In_2438,In_2096);
nor U1060 (N_1060,In_428,In_2823);
and U1061 (N_1061,In_2231,In_1959);
nor U1062 (N_1062,In_1483,In_2921);
nand U1063 (N_1063,In_1217,In_804);
and U1064 (N_1064,In_1398,In_2086);
xor U1065 (N_1065,In_760,In_1961);
xor U1066 (N_1066,In_285,In_1569);
xor U1067 (N_1067,In_28,In_2624);
and U1068 (N_1068,In_1090,In_1467);
or U1069 (N_1069,In_643,In_359);
and U1070 (N_1070,In_2594,In_2463);
and U1071 (N_1071,In_2672,In_2909);
or U1072 (N_1072,In_338,In_1088);
xor U1073 (N_1073,In_2035,In_2687);
xor U1074 (N_1074,In_1805,In_2196);
xnor U1075 (N_1075,In_810,In_1813);
nor U1076 (N_1076,In_1818,In_1946);
nor U1077 (N_1077,In_2911,In_2530);
and U1078 (N_1078,In_2129,In_1751);
xnor U1079 (N_1079,In_2309,In_235);
or U1080 (N_1080,In_603,In_2844);
nand U1081 (N_1081,In_1379,In_188);
and U1082 (N_1082,In_1528,In_981);
nor U1083 (N_1083,In_1475,In_2619);
or U1084 (N_1084,In_2484,In_2166);
nor U1085 (N_1085,In_1757,In_2009);
xnor U1086 (N_1086,In_995,In_1557);
nand U1087 (N_1087,In_266,In_270);
and U1088 (N_1088,In_927,In_690);
nor U1089 (N_1089,In_2067,In_983);
or U1090 (N_1090,In_1127,In_259);
or U1091 (N_1091,In_2099,In_2356);
xnor U1092 (N_1092,In_1729,In_566);
and U1093 (N_1093,In_352,In_1093);
or U1094 (N_1094,In_286,In_1248);
nand U1095 (N_1095,In_2076,In_2503);
nor U1096 (N_1096,In_2972,In_1492);
xor U1097 (N_1097,In_2695,In_1235);
nand U1098 (N_1098,In_1275,In_2259);
nand U1099 (N_1099,In_251,In_551);
or U1100 (N_1100,In_2055,In_43);
xor U1101 (N_1101,In_118,In_717);
nand U1102 (N_1102,In_2470,In_549);
and U1103 (N_1103,In_1143,In_956);
nand U1104 (N_1104,In_1041,In_1606);
nand U1105 (N_1105,In_822,In_167);
xor U1106 (N_1106,In_1956,In_1120);
and U1107 (N_1107,In_2517,In_1506);
or U1108 (N_1108,In_936,In_875);
or U1109 (N_1109,In_2659,In_2873);
nand U1110 (N_1110,In_1474,In_2149);
or U1111 (N_1111,In_1906,In_2241);
nor U1112 (N_1112,In_586,In_647);
and U1113 (N_1113,In_1932,In_1720);
or U1114 (N_1114,In_385,In_1573);
nand U1115 (N_1115,In_1112,In_521);
and U1116 (N_1116,In_1361,In_2606);
nand U1117 (N_1117,In_542,In_2979);
or U1118 (N_1118,In_2625,In_2638);
xnor U1119 (N_1119,In_526,In_1170);
and U1120 (N_1120,In_1830,In_35);
or U1121 (N_1121,In_1604,In_672);
nor U1122 (N_1122,In_425,In_1220);
nand U1123 (N_1123,In_1649,In_823);
nor U1124 (N_1124,In_920,In_1934);
xnor U1125 (N_1125,In_2201,In_1582);
xor U1126 (N_1126,In_2446,In_1669);
or U1127 (N_1127,In_1754,In_2556);
and U1128 (N_1128,In_2350,In_2190);
nor U1129 (N_1129,In_705,In_1326);
nor U1130 (N_1130,In_1559,In_1083);
and U1131 (N_1131,In_1186,In_2796);
nor U1132 (N_1132,In_2109,In_339);
xnor U1133 (N_1133,In_2332,In_1714);
xnor U1134 (N_1134,In_2714,In_2151);
or U1135 (N_1135,In_1795,In_356);
nand U1136 (N_1136,In_204,In_820);
or U1137 (N_1137,In_2642,In_2447);
xnor U1138 (N_1138,In_1601,In_53);
nor U1139 (N_1139,In_2437,In_342);
nand U1140 (N_1140,In_2472,In_2608);
nand U1141 (N_1141,In_2562,In_447);
nand U1142 (N_1142,In_1940,In_509);
xnor U1143 (N_1143,In_641,In_1133);
or U1144 (N_1144,In_1184,In_1584);
nor U1145 (N_1145,In_127,In_2928);
nand U1146 (N_1146,In_1207,In_82);
nand U1147 (N_1147,In_2965,In_2559);
and U1148 (N_1148,In_1408,In_902);
nand U1149 (N_1149,In_60,In_1731);
xor U1150 (N_1150,In_1045,In_223);
and U1151 (N_1151,In_1771,In_2866);
and U1152 (N_1152,In_761,In_2480);
nor U1153 (N_1153,In_917,In_46);
or U1154 (N_1154,In_2912,In_768);
or U1155 (N_1155,In_2727,In_293);
and U1156 (N_1156,In_1310,In_2016);
nand U1157 (N_1157,In_1040,In_2421);
nor U1158 (N_1158,In_800,In_2828);
nor U1159 (N_1159,In_1995,In_1438);
or U1160 (N_1160,In_1854,In_1585);
nand U1161 (N_1161,In_2671,In_1615);
xor U1162 (N_1162,In_855,In_1341);
nor U1163 (N_1163,In_1204,In_2676);
nor U1164 (N_1164,In_94,In_2335);
nand U1165 (N_1165,In_483,In_446);
nor U1166 (N_1166,In_102,In_650);
nor U1167 (N_1167,In_1250,In_348);
xor U1168 (N_1168,In_548,In_1655);
xnor U1169 (N_1169,In_1330,In_2071);
nand U1170 (N_1170,In_1387,In_1798);
nand U1171 (N_1171,In_1548,In_2289);
and U1172 (N_1172,In_2034,In_829);
nor U1173 (N_1173,In_1098,In_236);
nand U1174 (N_1174,In_1931,In_653);
nand U1175 (N_1175,In_2729,In_2550);
nand U1176 (N_1176,In_2898,In_205);
xnor U1177 (N_1177,In_192,In_1270);
or U1178 (N_1178,In_45,In_1802);
xnor U1179 (N_1179,In_1023,In_1983);
nor U1180 (N_1180,In_2723,In_190);
xnor U1181 (N_1181,In_1616,In_306);
nor U1182 (N_1182,In_916,In_159);
nand U1183 (N_1183,In_2478,In_64);
and U1184 (N_1184,In_1136,In_1614);
xnor U1185 (N_1185,In_2112,In_930);
xnor U1186 (N_1186,In_1181,In_2740);
nand U1187 (N_1187,In_2632,In_505);
or U1188 (N_1188,In_300,In_1380);
or U1189 (N_1189,In_332,In_1449);
and U1190 (N_1190,In_1085,In_378);
nor U1191 (N_1191,In_1025,In_2633);
nand U1192 (N_1192,In_1463,In_1811);
nand U1193 (N_1193,In_2304,In_2142);
nor U1194 (N_1194,In_2812,In_1730);
nor U1195 (N_1195,In_1287,In_1661);
nand U1196 (N_1196,In_794,In_1092);
nor U1197 (N_1197,In_785,In_1302);
nand U1198 (N_1198,In_2439,In_181);
and U1199 (N_1199,In_1294,In_2751);
or U1200 (N_1200,In_2629,In_189);
or U1201 (N_1201,In_1290,In_2597);
nand U1202 (N_1202,In_2957,In_2402);
or U1203 (N_1203,In_57,In_2770);
xor U1204 (N_1204,In_589,In_38);
nor U1205 (N_1205,In_1712,In_1704);
or U1206 (N_1206,In_2181,In_1404);
nor U1207 (N_1207,In_1913,In_1547);
or U1208 (N_1208,In_2235,In_404);
xor U1209 (N_1209,In_714,In_2977);
nand U1210 (N_1210,In_2052,In_2057);
nand U1211 (N_1211,In_2669,In_487);
nor U1212 (N_1212,In_2781,In_1884);
nor U1213 (N_1213,In_2724,In_914);
nor U1214 (N_1214,In_2923,In_1610);
nand U1215 (N_1215,In_488,In_2610);
and U1216 (N_1216,In_627,In_530);
nor U1217 (N_1217,In_491,In_2529);
or U1218 (N_1218,In_955,In_1832);
xnor U1219 (N_1219,In_1281,In_2917);
or U1220 (N_1220,In_541,In_1767);
or U1221 (N_1221,In_2755,In_282);
xor U1222 (N_1222,In_2712,In_2704);
nor U1223 (N_1223,In_2507,In_1759);
or U1224 (N_1224,In_710,In_1346);
or U1225 (N_1225,In_1200,In_2713);
nor U1226 (N_1226,In_2299,In_2042);
nand U1227 (N_1227,In_1386,In_2030);
xnor U1228 (N_1228,In_1927,In_1500);
and U1229 (N_1229,In_1670,In_1348);
and U1230 (N_1230,In_2442,In_1237);
xnor U1231 (N_1231,In_70,In_946);
and U1232 (N_1232,In_442,In_1578);
nand U1233 (N_1233,In_382,In_1225);
and U1234 (N_1234,In_89,In_1318);
and U1235 (N_1235,In_214,In_1567);
xnor U1236 (N_1236,In_1451,In_1965);
and U1237 (N_1237,In_1465,In_2006);
or U1238 (N_1238,In_896,In_200);
xor U1239 (N_1239,In_1865,In_2020);
nand U1240 (N_1240,In_2380,In_2505);
or U1241 (N_1241,In_1850,In_1309);
nand U1242 (N_1242,In_2192,In_2743);
and U1243 (N_1243,In_2102,In_1401);
xor U1244 (N_1244,In_2958,In_2075);
xnor U1245 (N_1245,In_23,In_2323);
or U1246 (N_1246,In_435,In_1643);
nand U1247 (N_1247,In_655,In_2660);
xor U1248 (N_1248,In_2390,In_2930);
nor U1249 (N_1249,In_1650,In_1233);
and U1250 (N_1250,In_2243,In_2344);
xor U1251 (N_1251,In_963,In_2378);
nand U1252 (N_1252,In_1519,In_2077);
xor U1253 (N_1253,In_1875,In_1365);
and U1254 (N_1254,In_2418,In_1316);
or U1255 (N_1255,In_664,In_923);
xor U1256 (N_1256,In_764,In_1240);
xnor U1257 (N_1257,In_1735,In_2456);
nand U1258 (N_1258,In_2722,In_1325);
and U1259 (N_1259,In_2167,In_2386);
nor U1260 (N_1260,In_2039,In_1849);
and U1261 (N_1261,In_528,In_75);
xor U1262 (N_1262,In_376,In_2868);
or U1263 (N_1263,In_634,In_2511);
nand U1264 (N_1264,In_2280,In_502);
or U1265 (N_1265,In_2307,In_1297);
xor U1266 (N_1266,In_418,In_2646);
nor U1267 (N_1267,In_247,In_1067);
or U1268 (N_1268,In_704,In_1659);
and U1269 (N_1269,In_2819,In_182);
xnor U1270 (N_1270,In_206,In_2806);
nor U1271 (N_1271,In_14,In_2680);
xnor U1272 (N_1272,In_1666,In_1115);
xor U1273 (N_1273,In_1848,In_1103);
or U1274 (N_1274,In_2995,In_2458);
or U1275 (N_1275,In_924,In_999);
xnor U1276 (N_1276,In_2079,In_1074);
xor U1277 (N_1277,In_909,In_405);
xnor U1278 (N_1278,In_1280,In_255);
xor U1279 (N_1279,In_37,In_495);
nand U1280 (N_1280,In_2526,In_2572);
xor U1281 (N_1281,In_135,In_1789);
or U1282 (N_1282,In_1164,In_2364);
xor U1283 (N_1283,In_366,In_697);
or U1284 (N_1284,In_2540,In_1165);
or U1285 (N_1285,In_4,In_649);
nor U1286 (N_1286,In_982,In_1177);
xnor U1287 (N_1287,In_1521,In_539);
and U1288 (N_1288,In_2381,In_399);
nor U1289 (N_1289,In_1866,In_2046);
xnor U1290 (N_1290,In_1479,In_864);
and U1291 (N_1291,In_482,In_465);
xnor U1292 (N_1292,In_2058,In_580);
xnor U1293 (N_1293,In_1097,In_1499);
xor U1294 (N_1294,In_997,In_115);
or U1295 (N_1295,In_599,In_1954);
and U1296 (N_1296,In_1688,In_2878);
or U1297 (N_1297,In_1779,In_1105);
xor U1298 (N_1298,In_2126,In_2162);
nor U1299 (N_1299,In_2028,In_1545);
nand U1300 (N_1300,In_451,In_2147);
and U1301 (N_1301,In_2199,In_198);
nor U1302 (N_1302,In_796,In_1159);
xor U1303 (N_1303,In_1709,In_1539);
or U1304 (N_1304,In_2570,In_1158);
and U1305 (N_1305,In_2544,In_377);
or U1306 (N_1306,In_1918,In_1374);
nor U1307 (N_1307,In_2459,In_239);
nor U1308 (N_1308,In_2302,In_2382);
nor U1309 (N_1309,In_2948,In_2413);
or U1310 (N_1310,In_626,In_1746);
xnor U1311 (N_1311,In_749,In_313);
or U1312 (N_1312,In_2858,In_410);
xnor U1313 (N_1313,In_1337,In_845);
and U1314 (N_1314,In_1958,In_1462);
and U1315 (N_1315,In_2782,In_1826);
nor U1316 (N_1316,In_388,In_1426);
xor U1317 (N_1317,In_219,In_1409);
nand U1318 (N_1318,In_876,In_1756);
or U1319 (N_1319,In_65,In_2108);
nand U1320 (N_1320,In_139,In_2914);
or U1321 (N_1321,In_2689,In_475);
or U1322 (N_1322,In_582,In_427);
and U1323 (N_1323,In_1987,In_669);
or U1324 (N_1324,In_2236,In_411);
nand U1325 (N_1325,In_173,In_371);
and U1326 (N_1326,In_2974,In_443);
or U1327 (N_1327,In_2515,In_2872);
or U1328 (N_1328,In_832,In_729);
nand U1329 (N_1329,In_2717,In_1520);
nand U1330 (N_1330,In_988,In_898);
nand U1331 (N_1331,In_2817,In_262);
nand U1332 (N_1332,In_1015,In_2667);
and U1333 (N_1333,In_2822,In_1036);
xor U1334 (N_1334,In_1008,In_918);
and U1335 (N_1335,In_1157,In_11);
or U1336 (N_1336,In_1613,In_741);
xnor U1337 (N_1337,In_1489,In_1119);
nor U1338 (N_1338,In_2752,In_1657);
xor U1339 (N_1339,In_61,In_670);
or U1340 (N_1340,In_185,In_458);
and U1341 (N_1341,In_2534,In_642);
nor U1342 (N_1342,In_622,In_2158);
nor U1343 (N_1343,In_408,In_2969);
or U1344 (N_1344,In_2882,In_233);
or U1345 (N_1345,In_2287,In_8);
xnor U1346 (N_1346,In_2984,In_965);
or U1347 (N_1347,In_2989,In_2053);
nand U1348 (N_1348,In_2750,In_2996);
nor U1349 (N_1349,In_2114,In_2136);
nand U1350 (N_1350,In_2341,In_935);
or U1351 (N_1351,In_2904,In_1816);
and U1352 (N_1352,In_1472,In_1034);
nand U1353 (N_1353,In_662,In_2318);
or U1354 (N_1354,In_29,In_1026);
or U1355 (N_1355,In_897,In_727);
nand U1356 (N_1356,In_2372,In_1923);
xor U1357 (N_1357,In_1658,In_1011);
or U1358 (N_1358,In_2128,In_2265);
or U1359 (N_1359,In_1589,In_1841);
or U1360 (N_1360,In_748,In_2272);
nor U1361 (N_1361,In_1327,In_2244);
xnor U1362 (N_1362,In_1625,In_737);
and U1363 (N_1363,In_249,In_208);
and U1364 (N_1364,In_811,In_1383);
nor U1365 (N_1365,In_2054,In_790);
xor U1366 (N_1366,In_1551,In_780);
nor U1367 (N_1367,In_1765,In_2017);
and U1368 (N_1368,In_2429,In_695);
or U1369 (N_1369,In_654,In_835);
nor U1370 (N_1370,In_1574,In_1197);
xnor U1371 (N_1371,In_1450,In_928);
nand U1372 (N_1372,In_1315,In_1457);
and U1373 (N_1373,In_775,In_27);
nor U1374 (N_1374,In_420,In_2790);
nand U1375 (N_1375,In_1680,In_635);
nor U1376 (N_1376,In_373,In_1032);
and U1377 (N_1377,In_680,In_2360);
xnor U1378 (N_1378,In_1214,In_2910);
nand U1379 (N_1379,In_1544,In_1328);
or U1380 (N_1380,In_2051,In_1166);
nand U1381 (N_1381,In_2184,In_903);
and U1382 (N_1382,In_1205,In_2896);
xor U1383 (N_1383,In_292,In_2994);
and U1384 (N_1384,In_736,In_2066);
xnor U1385 (N_1385,In_2582,In_899);
xor U1386 (N_1386,In_1360,In_1951);
nor U1387 (N_1387,In_2551,In_1174);
nand U1388 (N_1388,In_1691,In_498);
and U1389 (N_1389,In_720,In_869);
nor U1390 (N_1390,In_1581,In_926);
and U1391 (N_1391,In_2864,In_1286);
or U1392 (N_1392,In_2172,In_2883);
or U1393 (N_1393,In_693,In_885);
nand U1394 (N_1394,In_1944,In_1675);
and U1395 (N_1395,In_195,In_2788);
nand U1396 (N_1396,In_222,In_986);
nand U1397 (N_1397,In_327,In_1748);
nand U1398 (N_1398,In_2249,In_2757);
and U1399 (N_1399,In_828,In_2406);
nor U1400 (N_1400,In_1575,In_99);
or U1401 (N_1401,In_758,In_1690);
or U1402 (N_1402,In_362,In_406);
or U1403 (N_1403,In_2132,In_32);
nor U1404 (N_1404,In_2815,In_168);
or U1405 (N_1405,In_637,In_1357);
or U1406 (N_1406,In_1486,In_2955);
nor U1407 (N_1407,In_84,In_2008);
xnor U1408 (N_1408,In_2050,In_2553);
xor U1409 (N_1409,In_2728,In_1010);
nor U1410 (N_1410,In_877,In_350);
nand U1411 (N_1411,In_951,In_2405);
nand U1412 (N_1412,In_2504,In_415);
or U1413 (N_1413,In_1555,In_358);
xor U1414 (N_1414,In_2213,In_2263);
xor U1415 (N_1415,In_1320,In_2070);
or U1416 (N_1416,In_1095,In_2853);
nand U1417 (N_1417,In_1228,In_787);
xnor U1418 (N_1418,In_696,In_974);
or U1419 (N_1419,In_349,In_1224);
nor U1420 (N_1420,In_2949,In_140);
nand U1421 (N_1421,In_1498,In_1624);
nor U1422 (N_1422,In_2436,In_455);
or U1423 (N_1423,In_798,In_328);
nand U1424 (N_1424,In_2720,In_1706);
nand U1425 (N_1425,In_2652,In_2121);
xor U1426 (N_1426,In_954,In_44);
nand U1427 (N_1427,In_396,In_1155);
and U1428 (N_1428,In_631,In_2527);
or U1429 (N_1429,In_2998,In_466);
nand U1430 (N_1430,In_18,In_2777);
and U1431 (N_1431,In_1901,In_571);
and U1432 (N_1432,In_1431,In_2113);
xor U1433 (N_1433,In_1744,In_894);
nand U1434 (N_1434,In_312,In_1558);
and U1435 (N_1435,In_2736,In_1683);
xnor U1436 (N_1436,In_1261,In_2634);
or U1437 (N_1437,In_683,In_320);
nor U1438 (N_1438,In_861,In_1857);
or U1439 (N_1439,In_2251,In_2120);
xor U1440 (N_1440,In_1147,In_493);
and U1441 (N_1441,In_216,In_1226);
and U1442 (N_1442,In_1385,In_33);
nor U1443 (N_1443,In_1768,In_1279);
nor U1444 (N_1444,In_1568,In_2662);
or U1445 (N_1445,In_108,In_1358);
nand U1446 (N_1446,In_2376,In_1778);
nand U1447 (N_1447,In_1437,In_1188);
nand U1448 (N_1448,In_144,In_85);
xnor U1449 (N_1449,In_745,In_942);
or U1450 (N_1450,In_333,In_2754);
and U1451 (N_1451,In_1264,In_1397);
nor U1452 (N_1452,In_2618,In_283);
nand U1453 (N_1453,In_1193,In_767);
nand U1454 (N_1454,In_1502,In_191);
or U1455 (N_1455,In_1641,In_471);
nand U1456 (N_1456,In_88,In_2314);
nand U1457 (N_1457,In_2716,In_2707);
nor U1458 (N_1458,In_2678,In_617);
nand U1459 (N_1459,In_1799,In_2737);
xor U1460 (N_1460,In_522,In_707);
xnor U1461 (N_1461,In_789,In_520);
and U1462 (N_1462,In_2269,In_1058);
xor U1463 (N_1463,In_908,In_991);
nor U1464 (N_1464,In_3,In_1915);
nor U1465 (N_1465,In_730,In_2726);
nor U1466 (N_1466,In_573,In_1391);
xnor U1467 (N_1467,In_2159,In_1508);
or U1468 (N_1468,In_2362,In_1762);
nor U1469 (N_1469,In_1531,In_1873);
nor U1470 (N_1470,In_257,In_2663);
nor U1471 (N_1471,In_1563,In_679);
and U1472 (N_1472,In_1390,In_289);
nand U1473 (N_1473,In_1543,In_1047);
or U1474 (N_1474,In_1546,In_738);
and U1475 (N_1475,In_2523,In_1229);
xnor U1476 (N_1476,In_1178,In_2310);
and U1477 (N_1477,In_2748,In_2813);
nor U1478 (N_1478,In_1153,In_1150);
xnor U1479 (N_1479,In_1533,In_2157);
or U1480 (N_1480,In_2744,In_2098);
nor U1481 (N_1481,In_1488,In_2575);
and U1482 (N_1482,In_1293,In_556);
nor U1483 (N_1483,In_1277,In_1332);
nand U1484 (N_1484,In_2282,In_1633);
and U1485 (N_1485,In_414,In_1786);
or U1486 (N_1486,In_2999,In_2445);
nor U1487 (N_1487,In_202,In_743);
or U1488 (N_1488,In_725,In_2775);
and U1489 (N_1489,In_2514,In_2450);
nand U1490 (N_1490,In_2212,In_2774);
xnor U1491 (N_1491,In_2985,In_1268);
and U1492 (N_1492,In_2733,In_132);
and U1493 (N_1493,In_1117,In_959);
and U1494 (N_1494,In_2216,In_1855);
or U1495 (N_1495,In_2839,In_2769);
or U1496 (N_1496,In_1656,In_507);
or U1497 (N_1497,In_162,In_1072);
nor U1498 (N_1498,In_1482,In_0);
nor U1499 (N_1499,In_1314,In_1000);
or U1500 (N_1500,In_997,In_1296);
nor U1501 (N_1501,In_1895,In_1660);
nand U1502 (N_1502,In_1405,In_604);
or U1503 (N_1503,In_2830,In_625);
or U1504 (N_1504,In_2763,In_605);
or U1505 (N_1505,In_2642,In_2957);
or U1506 (N_1506,In_638,In_2527);
or U1507 (N_1507,In_2721,In_686);
or U1508 (N_1508,In_2853,In_1254);
or U1509 (N_1509,In_2275,In_484);
or U1510 (N_1510,In_1736,In_320);
nand U1511 (N_1511,In_501,In_2012);
nor U1512 (N_1512,In_1319,In_2751);
nand U1513 (N_1513,In_49,In_1786);
xnor U1514 (N_1514,In_523,In_2027);
xnor U1515 (N_1515,In_1170,In_2184);
nor U1516 (N_1516,In_40,In_2995);
nand U1517 (N_1517,In_1177,In_707);
and U1518 (N_1518,In_2805,In_1662);
nand U1519 (N_1519,In_2507,In_1590);
nor U1520 (N_1520,In_1530,In_450);
xnor U1521 (N_1521,In_1872,In_728);
or U1522 (N_1522,In_1528,In_1288);
or U1523 (N_1523,In_1185,In_1821);
nand U1524 (N_1524,In_286,In_2970);
and U1525 (N_1525,In_443,In_2734);
nand U1526 (N_1526,In_1188,In_524);
nand U1527 (N_1527,In_1438,In_2260);
nor U1528 (N_1528,In_2577,In_2300);
xnor U1529 (N_1529,In_1834,In_135);
and U1530 (N_1530,In_2394,In_29);
and U1531 (N_1531,In_1535,In_76);
nand U1532 (N_1532,In_2732,In_2080);
or U1533 (N_1533,In_2923,In_1351);
nor U1534 (N_1534,In_2605,In_2862);
nor U1535 (N_1535,In_473,In_259);
nand U1536 (N_1536,In_1413,In_931);
and U1537 (N_1537,In_2754,In_235);
xor U1538 (N_1538,In_1600,In_2490);
nor U1539 (N_1539,In_2813,In_359);
nor U1540 (N_1540,In_1458,In_2710);
nor U1541 (N_1541,In_1875,In_2452);
or U1542 (N_1542,In_2166,In_2379);
nand U1543 (N_1543,In_898,In_2507);
nor U1544 (N_1544,In_401,In_2146);
or U1545 (N_1545,In_1648,In_1431);
or U1546 (N_1546,In_2398,In_1590);
or U1547 (N_1547,In_885,In_372);
xnor U1548 (N_1548,In_1362,In_692);
or U1549 (N_1549,In_2383,In_2360);
xor U1550 (N_1550,In_1545,In_1932);
nor U1551 (N_1551,In_695,In_2963);
nor U1552 (N_1552,In_2411,In_1404);
xnor U1553 (N_1553,In_734,In_182);
xor U1554 (N_1554,In_2379,In_868);
nor U1555 (N_1555,In_440,In_1339);
and U1556 (N_1556,In_937,In_2723);
or U1557 (N_1557,In_2989,In_808);
nor U1558 (N_1558,In_2575,In_2651);
xnor U1559 (N_1559,In_466,In_1254);
nor U1560 (N_1560,In_249,In_325);
or U1561 (N_1561,In_2351,In_2532);
nor U1562 (N_1562,In_12,In_629);
or U1563 (N_1563,In_1387,In_474);
nand U1564 (N_1564,In_2495,In_2803);
xor U1565 (N_1565,In_2745,In_2593);
xor U1566 (N_1566,In_1861,In_1737);
and U1567 (N_1567,In_1359,In_1661);
or U1568 (N_1568,In_305,In_1365);
nand U1569 (N_1569,In_1852,In_1084);
nand U1570 (N_1570,In_2777,In_423);
nand U1571 (N_1571,In_1280,In_2377);
nand U1572 (N_1572,In_1815,In_1778);
nor U1573 (N_1573,In_1880,In_1784);
or U1574 (N_1574,In_2151,In_1093);
nand U1575 (N_1575,In_2233,In_2888);
and U1576 (N_1576,In_953,In_1231);
or U1577 (N_1577,In_1277,In_1025);
or U1578 (N_1578,In_1391,In_633);
xnor U1579 (N_1579,In_2213,In_148);
nor U1580 (N_1580,In_761,In_959);
nor U1581 (N_1581,In_959,In_2147);
or U1582 (N_1582,In_353,In_2865);
and U1583 (N_1583,In_1324,In_91);
xnor U1584 (N_1584,In_2903,In_62);
nand U1585 (N_1585,In_2093,In_2160);
xnor U1586 (N_1586,In_1427,In_2798);
xnor U1587 (N_1587,In_698,In_1867);
or U1588 (N_1588,In_2848,In_2614);
nand U1589 (N_1589,In_2533,In_753);
and U1590 (N_1590,In_2774,In_2806);
nand U1591 (N_1591,In_2264,In_308);
or U1592 (N_1592,In_2513,In_1146);
xnor U1593 (N_1593,In_1447,In_2222);
or U1594 (N_1594,In_2038,In_2769);
xnor U1595 (N_1595,In_396,In_2221);
nand U1596 (N_1596,In_2194,In_1075);
or U1597 (N_1597,In_102,In_1947);
xnor U1598 (N_1598,In_1133,In_1642);
or U1599 (N_1599,In_24,In_513);
nor U1600 (N_1600,In_1654,In_2831);
xnor U1601 (N_1601,In_1475,In_561);
or U1602 (N_1602,In_918,In_1987);
nor U1603 (N_1603,In_454,In_200);
nand U1604 (N_1604,In_22,In_2304);
or U1605 (N_1605,In_118,In_457);
nor U1606 (N_1606,In_2346,In_1866);
nor U1607 (N_1607,In_2766,In_2105);
and U1608 (N_1608,In_2587,In_1693);
and U1609 (N_1609,In_2954,In_1893);
or U1610 (N_1610,In_2346,In_60);
or U1611 (N_1611,In_1322,In_1469);
or U1612 (N_1612,In_926,In_1239);
nor U1613 (N_1613,In_1616,In_313);
nor U1614 (N_1614,In_788,In_2545);
nor U1615 (N_1615,In_2656,In_709);
xor U1616 (N_1616,In_1342,In_849);
and U1617 (N_1617,In_401,In_254);
and U1618 (N_1618,In_2598,In_2655);
and U1619 (N_1619,In_1792,In_2817);
or U1620 (N_1620,In_1949,In_1952);
and U1621 (N_1621,In_1568,In_335);
and U1622 (N_1622,In_806,In_626);
xnor U1623 (N_1623,In_1216,In_2797);
nor U1624 (N_1624,In_2338,In_1933);
or U1625 (N_1625,In_2170,In_2118);
nor U1626 (N_1626,In_1000,In_693);
xor U1627 (N_1627,In_1540,In_212);
or U1628 (N_1628,In_153,In_913);
or U1629 (N_1629,In_2586,In_1025);
nor U1630 (N_1630,In_1788,In_2510);
or U1631 (N_1631,In_1186,In_909);
nand U1632 (N_1632,In_987,In_2569);
nand U1633 (N_1633,In_1563,In_2657);
nor U1634 (N_1634,In_2811,In_1587);
nand U1635 (N_1635,In_2032,In_948);
and U1636 (N_1636,In_1856,In_985);
nand U1637 (N_1637,In_1309,In_519);
nor U1638 (N_1638,In_2914,In_2290);
nand U1639 (N_1639,In_1463,In_139);
and U1640 (N_1640,In_1233,In_2230);
and U1641 (N_1641,In_999,In_2831);
nand U1642 (N_1642,In_625,In_2394);
or U1643 (N_1643,In_2081,In_552);
nand U1644 (N_1644,In_2773,In_1057);
or U1645 (N_1645,In_2342,In_2104);
nor U1646 (N_1646,In_727,In_1898);
nor U1647 (N_1647,In_2931,In_767);
nand U1648 (N_1648,In_628,In_991);
and U1649 (N_1649,In_908,In_1384);
xor U1650 (N_1650,In_169,In_2120);
xor U1651 (N_1651,In_2588,In_2304);
or U1652 (N_1652,In_1359,In_942);
nor U1653 (N_1653,In_2294,In_1627);
xor U1654 (N_1654,In_1577,In_891);
nand U1655 (N_1655,In_518,In_467);
xnor U1656 (N_1656,In_997,In_1226);
nor U1657 (N_1657,In_614,In_1669);
xnor U1658 (N_1658,In_1186,In_1676);
or U1659 (N_1659,In_2710,In_1093);
nand U1660 (N_1660,In_2619,In_2065);
and U1661 (N_1661,In_548,In_1261);
and U1662 (N_1662,In_658,In_2697);
and U1663 (N_1663,In_1894,In_2696);
or U1664 (N_1664,In_1433,In_1829);
xnor U1665 (N_1665,In_2285,In_112);
or U1666 (N_1666,In_721,In_1371);
xnor U1667 (N_1667,In_1900,In_1596);
or U1668 (N_1668,In_614,In_1437);
xnor U1669 (N_1669,In_1572,In_2450);
nand U1670 (N_1670,In_2963,In_2884);
or U1671 (N_1671,In_1210,In_2933);
xor U1672 (N_1672,In_921,In_306);
nor U1673 (N_1673,In_647,In_2877);
xor U1674 (N_1674,In_2782,In_584);
xor U1675 (N_1675,In_803,In_2558);
xor U1676 (N_1676,In_1487,In_2969);
and U1677 (N_1677,In_436,In_925);
and U1678 (N_1678,In_2361,In_254);
and U1679 (N_1679,In_258,In_1945);
or U1680 (N_1680,In_1372,In_1625);
or U1681 (N_1681,In_750,In_1533);
xor U1682 (N_1682,In_2893,In_744);
xnor U1683 (N_1683,In_892,In_696);
nor U1684 (N_1684,In_1271,In_1505);
nor U1685 (N_1685,In_2384,In_1645);
xnor U1686 (N_1686,In_351,In_1188);
xnor U1687 (N_1687,In_2671,In_2129);
nor U1688 (N_1688,In_2309,In_2641);
nand U1689 (N_1689,In_1911,In_1561);
or U1690 (N_1690,In_1023,In_96);
or U1691 (N_1691,In_810,In_2965);
or U1692 (N_1692,In_1987,In_2419);
and U1693 (N_1693,In_868,In_1791);
and U1694 (N_1694,In_1239,In_2858);
or U1695 (N_1695,In_1586,In_2159);
nand U1696 (N_1696,In_2994,In_798);
nor U1697 (N_1697,In_1843,In_1633);
and U1698 (N_1698,In_1910,In_222);
or U1699 (N_1699,In_1287,In_2709);
nand U1700 (N_1700,In_2937,In_2280);
xor U1701 (N_1701,In_1773,In_328);
or U1702 (N_1702,In_1354,In_2966);
nand U1703 (N_1703,In_92,In_1695);
xor U1704 (N_1704,In_1456,In_2926);
nand U1705 (N_1705,In_646,In_1628);
and U1706 (N_1706,In_146,In_2977);
nor U1707 (N_1707,In_2291,In_283);
xnor U1708 (N_1708,In_2187,In_1983);
nand U1709 (N_1709,In_59,In_2932);
and U1710 (N_1710,In_157,In_2416);
and U1711 (N_1711,In_2376,In_1527);
nor U1712 (N_1712,In_2466,In_139);
nor U1713 (N_1713,In_1693,In_233);
nor U1714 (N_1714,In_116,In_306);
xor U1715 (N_1715,In_1207,In_2090);
and U1716 (N_1716,In_1808,In_2653);
nand U1717 (N_1717,In_2498,In_2108);
xor U1718 (N_1718,In_2078,In_2812);
and U1719 (N_1719,In_1842,In_1652);
nand U1720 (N_1720,In_2977,In_2325);
xor U1721 (N_1721,In_788,In_2702);
or U1722 (N_1722,In_1737,In_994);
xnor U1723 (N_1723,In_792,In_1536);
nor U1724 (N_1724,In_1119,In_2686);
nor U1725 (N_1725,In_2044,In_1852);
nand U1726 (N_1726,In_2497,In_1669);
or U1727 (N_1727,In_2346,In_1446);
nor U1728 (N_1728,In_1156,In_2);
or U1729 (N_1729,In_1862,In_984);
and U1730 (N_1730,In_1957,In_2751);
nor U1731 (N_1731,In_893,In_1419);
or U1732 (N_1732,In_1746,In_2049);
or U1733 (N_1733,In_2705,In_1798);
xor U1734 (N_1734,In_2184,In_1211);
and U1735 (N_1735,In_201,In_515);
or U1736 (N_1736,In_570,In_2287);
nand U1737 (N_1737,In_1993,In_2944);
nor U1738 (N_1738,In_940,In_2816);
nor U1739 (N_1739,In_2797,In_401);
nand U1740 (N_1740,In_214,In_1431);
nand U1741 (N_1741,In_2524,In_1896);
nor U1742 (N_1742,In_236,In_1335);
xor U1743 (N_1743,In_2470,In_2309);
or U1744 (N_1744,In_1576,In_2849);
or U1745 (N_1745,In_2519,In_2265);
or U1746 (N_1746,In_1821,In_726);
nor U1747 (N_1747,In_1083,In_2629);
and U1748 (N_1748,In_1913,In_1457);
nand U1749 (N_1749,In_1211,In_2823);
nor U1750 (N_1750,In_1489,In_2057);
nor U1751 (N_1751,In_1189,In_818);
xor U1752 (N_1752,In_366,In_2238);
xnor U1753 (N_1753,In_1687,In_796);
and U1754 (N_1754,In_607,In_1475);
xnor U1755 (N_1755,In_1325,In_1182);
or U1756 (N_1756,In_1,In_1224);
or U1757 (N_1757,In_495,In_73);
and U1758 (N_1758,In_2102,In_838);
and U1759 (N_1759,In_2807,In_2307);
and U1760 (N_1760,In_1621,In_467);
nor U1761 (N_1761,In_1632,In_1638);
xnor U1762 (N_1762,In_139,In_780);
and U1763 (N_1763,In_840,In_2447);
or U1764 (N_1764,In_1203,In_1129);
xor U1765 (N_1765,In_843,In_2144);
nand U1766 (N_1766,In_1822,In_1113);
xnor U1767 (N_1767,In_795,In_2978);
xnor U1768 (N_1768,In_2454,In_1346);
nand U1769 (N_1769,In_2769,In_2984);
xor U1770 (N_1770,In_2656,In_1500);
xor U1771 (N_1771,In_2236,In_1946);
xnor U1772 (N_1772,In_1812,In_944);
nor U1773 (N_1773,In_1235,In_2679);
nand U1774 (N_1774,In_1527,In_1098);
or U1775 (N_1775,In_2665,In_2995);
nand U1776 (N_1776,In_1112,In_753);
or U1777 (N_1777,In_2139,In_2298);
xor U1778 (N_1778,In_2395,In_732);
xnor U1779 (N_1779,In_2344,In_2385);
and U1780 (N_1780,In_2070,In_377);
nor U1781 (N_1781,In_177,In_1995);
or U1782 (N_1782,In_897,In_2849);
and U1783 (N_1783,In_2020,In_2219);
xnor U1784 (N_1784,In_1587,In_637);
or U1785 (N_1785,In_1585,In_1777);
nor U1786 (N_1786,In_2405,In_388);
nor U1787 (N_1787,In_1579,In_942);
nand U1788 (N_1788,In_425,In_2459);
nand U1789 (N_1789,In_801,In_2719);
or U1790 (N_1790,In_1051,In_1132);
or U1791 (N_1791,In_2338,In_2735);
nand U1792 (N_1792,In_838,In_55);
xor U1793 (N_1793,In_2011,In_243);
nand U1794 (N_1794,In_2178,In_1325);
or U1795 (N_1795,In_2272,In_2562);
nand U1796 (N_1796,In_995,In_2900);
nand U1797 (N_1797,In_1185,In_2260);
nand U1798 (N_1798,In_2997,In_825);
xnor U1799 (N_1799,In_635,In_2612);
and U1800 (N_1800,In_691,In_254);
and U1801 (N_1801,In_1911,In_474);
xor U1802 (N_1802,In_2578,In_2739);
or U1803 (N_1803,In_2239,In_2875);
and U1804 (N_1804,In_2019,In_2118);
nand U1805 (N_1805,In_399,In_2657);
nand U1806 (N_1806,In_2656,In_1617);
nand U1807 (N_1807,In_1426,In_713);
xnor U1808 (N_1808,In_2022,In_1999);
and U1809 (N_1809,In_1080,In_2894);
and U1810 (N_1810,In_1452,In_71);
nor U1811 (N_1811,In_54,In_105);
and U1812 (N_1812,In_759,In_2695);
or U1813 (N_1813,In_2295,In_976);
or U1814 (N_1814,In_1011,In_2971);
and U1815 (N_1815,In_2588,In_1384);
and U1816 (N_1816,In_2176,In_1302);
and U1817 (N_1817,In_168,In_349);
nor U1818 (N_1818,In_2989,In_2233);
nand U1819 (N_1819,In_2733,In_1571);
and U1820 (N_1820,In_844,In_2371);
nor U1821 (N_1821,In_1993,In_1040);
and U1822 (N_1822,In_2510,In_722);
xnor U1823 (N_1823,In_1972,In_2372);
and U1824 (N_1824,In_2177,In_140);
nand U1825 (N_1825,In_36,In_2929);
nand U1826 (N_1826,In_1156,In_52);
xnor U1827 (N_1827,In_2721,In_1167);
and U1828 (N_1828,In_550,In_1621);
xnor U1829 (N_1829,In_249,In_1289);
nand U1830 (N_1830,In_1688,In_2744);
or U1831 (N_1831,In_833,In_529);
xor U1832 (N_1832,In_537,In_2877);
and U1833 (N_1833,In_1260,In_2515);
nor U1834 (N_1834,In_465,In_2964);
nand U1835 (N_1835,In_598,In_261);
and U1836 (N_1836,In_835,In_1730);
nand U1837 (N_1837,In_2179,In_1146);
or U1838 (N_1838,In_1485,In_2794);
nand U1839 (N_1839,In_2256,In_133);
nor U1840 (N_1840,In_2602,In_1692);
nor U1841 (N_1841,In_2327,In_1489);
nor U1842 (N_1842,In_1985,In_774);
or U1843 (N_1843,In_2589,In_651);
nand U1844 (N_1844,In_1442,In_491);
or U1845 (N_1845,In_2169,In_632);
nand U1846 (N_1846,In_2351,In_1477);
nor U1847 (N_1847,In_1693,In_2849);
nand U1848 (N_1848,In_2640,In_1575);
nor U1849 (N_1849,In_941,In_1413);
xor U1850 (N_1850,In_1143,In_1541);
xnor U1851 (N_1851,In_2947,In_1203);
nand U1852 (N_1852,In_1502,In_2838);
nand U1853 (N_1853,In_1088,In_342);
nor U1854 (N_1854,In_1074,In_2790);
xor U1855 (N_1855,In_2569,In_2100);
or U1856 (N_1856,In_2952,In_780);
xor U1857 (N_1857,In_301,In_1774);
nand U1858 (N_1858,In_1415,In_2291);
nand U1859 (N_1859,In_298,In_987);
and U1860 (N_1860,In_27,In_391);
nor U1861 (N_1861,In_903,In_1569);
xor U1862 (N_1862,In_556,In_126);
nand U1863 (N_1863,In_752,In_1036);
and U1864 (N_1864,In_1482,In_1346);
nor U1865 (N_1865,In_2469,In_527);
nor U1866 (N_1866,In_277,In_647);
xor U1867 (N_1867,In_1107,In_406);
nor U1868 (N_1868,In_497,In_266);
nor U1869 (N_1869,In_1818,In_1465);
or U1870 (N_1870,In_478,In_115);
xnor U1871 (N_1871,In_2837,In_1853);
xnor U1872 (N_1872,In_1537,In_1877);
nor U1873 (N_1873,In_571,In_2798);
and U1874 (N_1874,In_1711,In_2275);
or U1875 (N_1875,In_1526,In_87);
and U1876 (N_1876,In_1808,In_978);
nand U1877 (N_1877,In_2404,In_1818);
xor U1878 (N_1878,In_922,In_1141);
xor U1879 (N_1879,In_1091,In_171);
or U1880 (N_1880,In_1100,In_435);
or U1881 (N_1881,In_1530,In_922);
nor U1882 (N_1882,In_2975,In_2799);
nand U1883 (N_1883,In_1913,In_2453);
nand U1884 (N_1884,In_2035,In_1782);
nand U1885 (N_1885,In_1139,In_1065);
xnor U1886 (N_1886,In_2008,In_2988);
nor U1887 (N_1887,In_2945,In_1952);
xnor U1888 (N_1888,In_1386,In_612);
and U1889 (N_1889,In_997,In_2075);
nor U1890 (N_1890,In_372,In_1209);
nor U1891 (N_1891,In_2379,In_2519);
and U1892 (N_1892,In_232,In_2218);
nand U1893 (N_1893,In_717,In_59);
or U1894 (N_1894,In_202,In_2049);
nor U1895 (N_1895,In_353,In_2520);
nor U1896 (N_1896,In_450,In_2199);
or U1897 (N_1897,In_1188,In_2734);
nor U1898 (N_1898,In_1320,In_628);
xor U1899 (N_1899,In_444,In_1215);
xor U1900 (N_1900,In_1989,In_2602);
nor U1901 (N_1901,In_1191,In_2740);
or U1902 (N_1902,In_2928,In_2749);
or U1903 (N_1903,In_2279,In_1209);
xnor U1904 (N_1904,In_521,In_366);
nand U1905 (N_1905,In_1899,In_456);
nor U1906 (N_1906,In_2794,In_2611);
nor U1907 (N_1907,In_2469,In_1380);
xnor U1908 (N_1908,In_268,In_2663);
and U1909 (N_1909,In_45,In_235);
or U1910 (N_1910,In_2464,In_2473);
or U1911 (N_1911,In_1178,In_2949);
nand U1912 (N_1912,In_542,In_739);
or U1913 (N_1913,In_1312,In_1181);
nand U1914 (N_1914,In_713,In_624);
or U1915 (N_1915,In_2763,In_2634);
and U1916 (N_1916,In_904,In_2343);
nor U1917 (N_1917,In_2668,In_1917);
xor U1918 (N_1918,In_2471,In_1458);
and U1919 (N_1919,In_2167,In_194);
or U1920 (N_1920,In_2606,In_554);
nand U1921 (N_1921,In_3,In_831);
nand U1922 (N_1922,In_547,In_1213);
and U1923 (N_1923,In_1200,In_2310);
nand U1924 (N_1924,In_1905,In_2411);
nand U1925 (N_1925,In_1155,In_1499);
and U1926 (N_1926,In_174,In_910);
and U1927 (N_1927,In_824,In_1790);
and U1928 (N_1928,In_2597,In_1851);
nand U1929 (N_1929,In_1267,In_1307);
xor U1930 (N_1930,In_968,In_548);
or U1931 (N_1931,In_2011,In_2210);
nand U1932 (N_1932,In_2750,In_1246);
and U1933 (N_1933,In_766,In_311);
or U1934 (N_1934,In_214,In_1115);
nand U1935 (N_1935,In_1315,In_1023);
nand U1936 (N_1936,In_108,In_1269);
nor U1937 (N_1937,In_2654,In_2726);
nor U1938 (N_1938,In_1396,In_1905);
or U1939 (N_1939,In_104,In_1454);
or U1940 (N_1940,In_2762,In_1485);
xnor U1941 (N_1941,In_102,In_501);
and U1942 (N_1942,In_1614,In_2259);
and U1943 (N_1943,In_59,In_2105);
xnor U1944 (N_1944,In_2729,In_2694);
xnor U1945 (N_1945,In_2191,In_2435);
nor U1946 (N_1946,In_2289,In_2488);
xnor U1947 (N_1947,In_925,In_34);
xnor U1948 (N_1948,In_2888,In_2449);
xnor U1949 (N_1949,In_342,In_2110);
nor U1950 (N_1950,In_2780,In_1996);
and U1951 (N_1951,In_1556,In_2250);
nand U1952 (N_1952,In_1865,In_855);
nor U1953 (N_1953,In_191,In_1991);
nor U1954 (N_1954,In_955,In_462);
nand U1955 (N_1955,In_884,In_1328);
xnor U1956 (N_1956,In_2915,In_1105);
nand U1957 (N_1957,In_1805,In_1479);
or U1958 (N_1958,In_1771,In_2988);
nor U1959 (N_1959,In_2847,In_194);
nor U1960 (N_1960,In_2412,In_2346);
or U1961 (N_1961,In_630,In_641);
and U1962 (N_1962,In_628,In_1283);
and U1963 (N_1963,In_717,In_698);
nor U1964 (N_1964,In_1486,In_234);
and U1965 (N_1965,In_1333,In_1542);
and U1966 (N_1966,In_328,In_274);
nor U1967 (N_1967,In_2688,In_620);
and U1968 (N_1968,In_633,In_2994);
nand U1969 (N_1969,In_1659,In_1242);
xor U1970 (N_1970,In_2352,In_1943);
or U1971 (N_1971,In_1926,In_2081);
xnor U1972 (N_1972,In_1006,In_261);
or U1973 (N_1973,In_824,In_491);
and U1974 (N_1974,In_1651,In_570);
xor U1975 (N_1975,In_572,In_50);
xnor U1976 (N_1976,In_2155,In_2011);
and U1977 (N_1977,In_2196,In_197);
nor U1978 (N_1978,In_2998,In_1058);
and U1979 (N_1979,In_275,In_2400);
or U1980 (N_1980,In_2062,In_595);
nor U1981 (N_1981,In_1280,In_1617);
or U1982 (N_1982,In_633,In_847);
or U1983 (N_1983,In_729,In_2560);
and U1984 (N_1984,In_1996,In_52);
nand U1985 (N_1985,In_2521,In_1929);
or U1986 (N_1986,In_1973,In_220);
xor U1987 (N_1987,In_1880,In_2356);
nand U1988 (N_1988,In_1719,In_2351);
nand U1989 (N_1989,In_2024,In_1989);
and U1990 (N_1990,In_855,In_2159);
nor U1991 (N_1991,In_1035,In_687);
xor U1992 (N_1992,In_331,In_1901);
xor U1993 (N_1993,In_2917,In_551);
or U1994 (N_1994,In_2430,In_1798);
and U1995 (N_1995,In_2783,In_2338);
xor U1996 (N_1996,In_2356,In_2239);
nor U1997 (N_1997,In_253,In_793);
nor U1998 (N_1998,In_1036,In_2612);
or U1999 (N_1999,In_762,In_831);
xor U2000 (N_2000,In_2839,In_2816);
nand U2001 (N_2001,In_97,In_392);
nor U2002 (N_2002,In_1049,In_1405);
or U2003 (N_2003,In_2531,In_540);
nand U2004 (N_2004,In_1636,In_2325);
and U2005 (N_2005,In_413,In_885);
xor U2006 (N_2006,In_2219,In_643);
nand U2007 (N_2007,In_2373,In_1224);
and U2008 (N_2008,In_1723,In_1076);
and U2009 (N_2009,In_1429,In_34);
and U2010 (N_2010,In_2376,In_2741);
nor U2011 (N_2011,In_521,In_2109);
nand U2012 (N_2012,In_694,In_457);
nand U2013 (N_2013,In_1413,In_1888);
xnor U2014 (N_2014,In_2006,In_2107);
nand U2015 (N_2015,In_1143,In_910);
or U2016 (N_2016,In_499,In_1186);
nor U2017 (N_2017,In_324,In_1183);
and U2018 (N_2018,In_146,In_1739);
or U2019 (N_2019,In_1748,In_1417);
nor U2020 (N_2020,In_60,In_817);
or U2021 (N_2021,In_1872,In_2517);
and U2022 (N_2022,In_2734,In_1916);
nand U2023 (N_2023,In_1463,In_355);
and U2024 (N_2024,In_337,In_2885);
xnor U2025 (N_2025,In_878,In_2934);
and U2026 (N_2026,In_2882,In_2381);
nand U2027 (N_2027,In_2076,In_231);
nand U2028 (N_2028,In_1513,In_1602);
and U2029 (N_2029,In_733,In_1508);
xor U2030 (N_2030,In_327,In_1723);
and U2031 (N_2031,In_543,In_1336);
or U2032 (N_2032,In_1555,In_1724);
and U2033 (N_2033,In_491,In_2832);
xnor U2034 (N_2034,In_1554,In_2589);
xnor U2035 (N_2035,In_1680,In_1045);
nor U2036 (N_2036,In_1831,In_2977);
nor U2037 (N_2037,In_1720,In_421);
xor U2038 (N_2038,In_908,In_1110);
and U2039 (N_2039,In_68,In_2555);
xor U2040 (N_2040,In_2686,In_2807);
xor U2041 (N_2041,In_1444,In_1753);
xnor U2042 (N_2042,In_2174,In_1763);
and U2043 (N_2043,In_104,In_1116);
and U2044 (N_2044,In_890,In_2978);
nor U2045 (N_2045,In_2929,In_1678);
and U2046 (N_2046,In_1757,In_475);
and U2047 (N_2047,In_2728,In_1923);
or U2048 (N_2048,In_533,In_7);
xnor U2049 (N_2049,In_2671,In_183);
xor U2050 (N_2050,In_2047,In_932);
or U2051 (N_2051,In_1078,In_2324);
nor U2052 (N_2052,In_2203,In_1559);
nor U2053 (N_2053,In_269,In_213);
or U2054 (N_2054,In_367,In_814);
xor U2055 (N_2055,In_683,In_6);
xor U2056 (N_2056,In_247,In_531);
or U2057 (N_2057,In_828,In_2190);
nor U2058 (N_2058,In_315,In_1260);
nand U2059 (N_2059,In_642,In_1573);
or U2060 (N_2060,In_1933,In_1697);
and U2061 (N_2061,In_281,In_864);
xnor U2062 (N_2062,In_833,In_740);
nand U2063 (N_2063,In_2159,In_1533);
xnor U2064 (N_2064,In_1805,In_2038);
nand U2065 (N_2065,In_2529,In_421);
and U2066 (N_2066,In_1563,In_2079);
nand U2067 (N_2067,In_2955,In_2184);
xnor U2068 (N_2068,In_2764,In_1384);
or U2069 (N_2069,In_2580,In_1320);
nand U2070 (N_2070,In_1701,In_1935);
nand U2071 (N_2071,In_1817,In_1535);
nand U2072 (N_2072,In_1523,In_329);
xor U2073 (N_2073,In_1948,In_2740);
nor U2074 (N_2074,In_1933,In_2624);
or U2075 (N_2075,In_484,In_2754);
nor U2076 (N_2076,In_1191,In_589);
xnor U2077 (N_2077,In_699,In_2397);
xor U2078 (N_2078,In_2610,In_2623);
or U2079 (N_2079,In_2682,In_746);
or U2080 (N_2080,In_909,In_631);
and U2081 (N_2081,In_1340,In_2732);
xor U2082 (N_2082,In_1965,In_1969);
and U2083 (N_2083,In_500,In_957);
xor U2084 (N_2084,In_2016,In_913);
nand U2085 (N_2085,In_506,In_451);
xor U2086 (N_2086,In_2713,In_1185);
nand U2087 (N_2087,In_1412,In_1348);
and U2088 (N_2088,In_2587,In_2183);
xor U2089 (N_2089,In_1194,In_2490);
nand U2090 (N_2090,In_2821,In_1059);
nor U2091 (N_2091,In_2681,In_1859);
xor U2092 (N_2092,In_2846,In_184);
or U2093 (N_2093,In_2673,In_1871);
nand U2094 (N_2094,In_1501,In_347);
and U2095 (N_2095,In_1408,In_1007);
nand U2096 (N_2096,In_1822,In_2395);
nor U2097 (N_2097,In_870,In_1646);
nand U2098 (N_2098,In_2046,In_1614);
and U2099 (N_2099,In_1856,In_1679);
nand U2100 (N_2100,In_723,In_176);
nand U2101 (N_2101,In_2174,In_2222);
nand U2102 (N_2102,In_2064,In_834);
nand U2103 (N_2103,In_2915,In_108);
and U2104 (N_2104,In_438,In_1512);
xor U2105 (N_2105,In_2832,In_376);
or U2106 (N_2106,In_2601,In_197);
or U2107 (N_2107,In_2118,In_537);
or U2108 (N_2108,In_987,In_2907);
or U2109 (N_2109,In_1979,In_445);
xnor U2110 (N_2110,In_102,In_191);
nor U2111 (N_2111,In_733,In_2118);
nand U2112 (N_2112,In_2017,In_2945);
xnor U2113 (N_2113,In_2656,In_1210);
or U2114 (N_2114,In_1062,In_109);
and U2115 (N_2115,In_1835,In_1789);
nand U2116 (N_2116,In_1688,In_2653);
nand U2117 (N_2117,In_1327,In_991);
and U2118 (N_2118,In_2171,In_2877);
nor U2119 (N_2119,In_438,In_1802);
or U2120 (N_2120,In_1863,In_2743);
nor U2121 (N_2121,In_2126,In_620);
nor U2122 (N_2122,In_1058,In_2131);
or U2123 (N_2123,In_2963,In_1646);
nor U2124 (N_2124,In_899,In_2788);
or U2125 (N_2125,In_2082,In_2536);
and U2126 (N_2126,In_1412,In_2801);
or U2127 (N_2127,In_238,In_2532);
nand U2128 (N_2128,In_744,In_235);
and U2129 (N_2129,In_1787,In_1338);
nor U2130 (N_2130,In_1651,In_1725);
xnor U2131 (N_2131,In_602,In_134);
or U2132 (N_2132,In_1966,In_2117);
and U2133 (N_2133,In_1278,In_1349);
nand U2134 (N_2134,In_593,In_1605);
nand U2135 (N_2135,In_2780,In_2834);
nor U2136 (N_2136,In_1748,In_2809);
or U2137 (N_2137,In_2863,In_754);
or U2138 (N_2138,In_1713,In_2548);
xor U2139 (N_2139,In_961,In_2290);
nand U2140 (N_2140,In_2654,In_733);
xnor U2141 (N_2141,In_2089,In_98);
and U2142 (N_2142,In_1791,In_1856);
nor U2143 (N_2143,In_21,In_188);
nand U2144 (N_2144,In_92,In_2797);
and U2145 (N_2145,In_768,In_2633);
nand U2146 (N_2146,In_2735,In_821);
and U2147 (N_2147,In_738,In_2495);
nor U2148 (N_2148,In_2336,In_371);
xnor U2149 (N_2149,In_1463,In_1028);
or U2150 (N_2150,In_164,In_2276);
nor U2151 (N_2151,In_2224,In_1331);
xor U2152 (N_2152,In_1807,In_2275);
nor U2153 (N_2153,In_549,In_217);
and U2154 (N_2154,In_205,In_487);
and U2155 (N_2155,In_341,In_1346);
and U2156 (N_2156,In_1490,In_390);
nand U2157 (N_2157,In_53,In_2835);
and U2158 (N_2158,In_1,In_219);
xor U2159 (N_2159,In_1230,In_2237);
xnor U2160 (N_2160,In_1029,In_1318);
and U2161 (N_2161,In_678,In_1686);
nor U2162 (N_2162,In_1140,In_932);
xnor U2163 (N_2163,In_1877,In_1442);
and U2164 (N_2164,In_2843,In_2203);
xnor U2165 (N_2165,In_2910,In_2481);
or U2166 (N_2166,In_2857,In_185);
and U2167 (N_2167,In_1850,In_825);
or U2168 (N_2168,In_2063,In_617);
or U2169 (N_2169,In_2592,In_1797);
or U2170 (N_2170,In_2368,In_1228);
nor U2171 (N_2171,In_2454,In_1040);
or U2172 (N_2172,In_840,In_443);
or U2173 (N_2173,In_1141,In_545);
nand U2174 (N_2174,In_754,In_877);
xor U2175 (N_2175,In_439,In_2914);
xor U2176 (N_2176,In_2883,In_317);
nand U2177 (N_2177,In_1463,In_619);
nand U2178 (N_2178,In_2551,In_828);
or U2179 (N_2179,In_914,In_1767);
or U2180 (N_2180,In_1614,In_2561);
nor U2181 (N_2181,In_108,In_88);
or U2182 (N_2182,In_2493,In_210);
or U2183 (N_2183,In_2382,In_1964);
or U2184 (N_2184,In_345,In_2004);
xor U2185 (N_2185,In_923,In_1916);
and U2186 (N_2186,In_588,In_291);
nand U2187 (N_2187,In_2829,In_2240);
nor U2188 (N_2188,In_2897,In_2472);
or U2189 (N_2189,In_206,In_1151);
nand U2190 (N_2190,In_1128,In_2654);
nor U2191 (N_2191,In_2439,In_1663);
xor U2192 (N_2192,In_2705,In_870);
nand U2193 (N_2193,In_2747,In_690);
xor U2194 (N_2194,In_637,In_177);
and U2195 (N_2195,In_2884,In_2612);
nor U2196 (N_2196,In_2920,In_2163);
nor U2197 (N_2197,In_289,In_274);
or U2198 (N_2198,In_2212,In_2444);
nor U2199 (N_2199,In_795,In_1019);
xnor U2200 (N_2200,In_397,In_1349);
nand U2201 (N_2201,In_2732,In_2873);
and U2202 (N_2202,In_1660,In_1010);
or U2203 (N_2203,In_546,In_2315);
nand U2204 (N_2204,In_2443,In_340);
xor U2205 (N_2205,In_623,In_2600);
xor U2206 (N_2206,In_1457,In_729);
and U2207 (N_2207,In_854,In_2818);
xor U2208 (N_2208,In_1366,In_2418);
nand U2209 (N_2209,In_795,In_403);
nor U2210 (N_2210,In_2560,In_1535);
and U2211 (N_2211,In_2646,In_2594);
nor U2212 (N_2212,In_1484,In_1817);
and U2213 (N_2213,In_2270,In_1383);
or U2214 (N_2214,In_326,In_980);
nand U2215 (N_2215,In_2409,In_2897);
and U2216 (N_2216,In_2422,In_341);
xor U2217 (N_2217,In_2105,In_69);
or U2218 (N_2218,In_1807,In_855);
nand U2219 (N_2219,In_1684,In_151);
and U2220 (N_2220,In_1359,In_1713);
nor U2221 (N_2221,In_1805,In_2953);
xnor U2222 (N_2222,In_2123,In_2536);
nor U2223 (N_2223,In_767,In_934);
nand U2224 (N_2224,In_1397,In_2626);
or U2225 (N_2225,In_1438,In_2709);
and U2226 (N_2226,In_2380,In_1283);
nand U2227 (N_2227,In_1503,In_1813);
or U2228 (N_2228,In_2703,In_627);
xnor U2229 (N_2229,In_266,In_666);
or U2230 (N_2230,In_2604,In_316);
nand U2231 (N_2231,In_2640,In_1376);
or U2232 (N_2232,In_440,In_86);
and U2233 (N_2233,In_957,In_47);
or U2234 (N_2234,In_1935,In_438);
nor U2235 (N_2235,In_729,In_634);
and U2236 (N_2236,In_605,In_409);
and U2237 (N_2237,In_934,In_294);
or U2238 (N_2238,In_2142,In_2943);
nor U2239 (N_2239,In_837,In_2927);
xor U2240 (N_2240,In_841,In_695);
nand U2241 (N_2241,In_2704,In_799);
nand U2242 (N_2242,In_1429,In_1443);
and U2243 (N_2243,In_1474,In_605);
and U2244 (N_2244,In_2458,In_1646);
or U2245 (N_2245,In_1087,In_1420);
nor U2246 (N_2246,In_1357,In_1015);
or U2247 (N_2247,In_708,In_2434);
or U2248 (N_2248,In_869,In_933);
and U2249 (N_2249,In_112,In_1975);
xnor U2250 (N_2250,In_1807,In_2641);
nor U2251 (N_2251,In_1978,In_889);
nand U2252 (N_2252,In_1547,In_1786);
nand U2253 (N_2253,In_596,In_2617);
nor U2254 (N_2254,In_2983,In_478);
nor U2255 (N_2255,In_1973,In_633);
nand U2256 (N_2256,In_505,In_112);
or U2257 (N_2257,In_2615,In_1823);
nand U2258 (N_2258,In_47,In_2486);
xnor U2259 (N_2259,In_2891,In_2828);
nor U2260 (N_2260,In_2406,In_2112);
xor U2261 (N_2261,In_2119,In_274);
or U2262 (N_2262,In_1731,In_492);
xnor U2263 (N_2263,In_1948,In_2327);
nand U2264 (N_2264,In_727,In_330);
and U2265 (N_2265,In_1296,In_2664);
or U2266 (N_2266,In_891,In_2528);
nand U2267 (N_2267,In_2023,In_1137);
nand U2268 (N_2268,In_1434,In_1317);
xor U2269 (N_2269,In_288,In_2812);
or U2270 (N_2270,In_2890,In_1315);
nor U2271 (N_2271,In_119,In_1749);
and U2272 (N_2272,In_820,In_2732);
nand U2273 (N_2273,In_1308,In_2741);
and U2274 (N_2274,In_498,In_1842);
and U2275 (N_2275,In_1484,In_1291);
nand U2276 (N_2276,In_484,In_645);
and U2277 (N_2277,In_123,In_486);
and U2278 (N_2278,In_2724,In_2437);
xnor U2279 (N_2279,In_830,In_2179);
nor U2280 (N_2280,In_1098,In_404);
nand U2281 (N_2281,In_560,In_2673);
nor U2282 (N_2282,In_2437,In_327);
and U2283 (N_2283,In_2303,In_690);
and U2284 (N_2284,In_2272,In_2612);
nand U2285 (N_2285,In_768,In_1460);
xor U2286 (N_2286,In_765,In_847);
xnor U2287 (N_2287,In_2744,In_1558);
xnor U2288 (N_2288,In_1365,In_763);
nor U2289 (N_2289,In_1067,In_2813);
xnor U2290 (N_2290,In_2635,In_1099);
or U2291 (N_2291,In_1355,In_1345);
nor U2292 (N_2292,In_581,In_807);
xor U2293 (N_2293,In_2452,In_1345);
nand U2294 (N_2294,In_101,In_88);
or U2295 (N_2295,In_449,In_347);
or U2296 (N_2296,In_2349,In_1644);
xor U2297 (N_2297,In_2307,In_2162);
xnor U2298 (N_2298,In_1699,In_1538);
nand U2299 (N_2299,In_2855,In_1505);
and U2300 (N_2300,In_1078,In_393);
nand U2301 (N_2301,In_2268,In_1528);
and U2302 (N_2302,In_769,In_1634);
nor U2303 (N_2303,In_123,In_2599);
nand U2304 (N_2304,In_1263,In_1931);
nor U2305 (N_2305,In_1786,In_2231);
and U2306 (N_2306,In_1241,In_890);
or U2307 (N_2307,In_450,In_995);
or U2308 (N_2308,In_1150,In_2610);
nand U2309 (N_2309,In_2326,In_565);
nor U2310 (N_2310,In_686,In_1737);
nand U2311 (N_2311,In_324,In_175);
xor U2312 (N_2312,In_1868,In_1625);
nand U2313 (N_2313,In_2515,In_2598);
nor U2314 (N_2314,In_1058,In_2751);
or U2315 (N_2315,In_2643,In_1005);
nand U2316 (N_2316,In_2169,In_86);
and U2317 (N_2317,In_2327,In_2376);
or U2318 (N_2318,In_1556,In_1563);
or U2319 (N_2319,In_2464,In_1464);
or U2320 (N_2320,In_144,In_2552);
xor U2321 (N_2321,In_1643,In_2818);
and U2322 (N_2322,In_307,In_1017);
xor U2323 (N_2323,In_1732,In_2369);
xor U2324 (N_2324,In_1886,In_470);
and U2325 (N_2325,In_596,In_1356);
nor U2326 (N_2326,In_908,In_1250);
xor U2327 (N_2327,In_2445,In_1006);
nor U2328 (N_2328,In_55,In_1291);
or U2329 (N_2329,In_1487,In_1216);
nand U2330 (N_2330,In_109,In_590);
and U2331 (N_2331,In_1595,In_1583);
xnor U2332 (N_2332,In_2414,In_1892);
nand U2333 (N_2333,In_2638,In_891);
xnor U2334 (N_2334,In_2248,In_1030);
nand U2335 (N_2335,In_1679,In_2040);
nor U2336 (N_2336,In_1135,In_1710);
and U2337 (N_2337,In_2918,In_2701);
nand U2338 (N_2338,In_1782,In_1243);
nand U2339 (N_2339,In_2324,In_884);
nor U2340 (N_2340,In_1105,In_1151);
nor U2341 (N_2341,In_1447,In_839);
nand U2342 (N_2342,In_2521,In_2345);
xnor U2343 (N_2343,In_366,In_2864);
nand U2344 (N_2344,In_2100,In_2734);
nor U2345 (N_2345,In_2559,In_2014);
nand U2346 (N_2346,In_574,In_1742);
xor U2347 (N_2347,In_246,In_591);
nor U2348 (N_2348,In_2289,In_2990);
and U2349 (N_2349,In_2686,In_2101);
or U2350 (N_2350,In_1474,In_586);
xnor U2351 (N_2351,In_814,In_728);
nor U2352 (N_2352,In_1188,In_1175);
xor U2353 (N_2353,In_749,In_2014);
xnor U2354 (N_2354,In_168,In_1082);
nor U2355 (N_2355,In_2793,In_2990);
and U2356 (N_2356,In_1320,In_1727);
xor U2357 (N_2357,In_123,In_560);
xnor U2358 (N_2358,In_1385,In_1105);
or U2359 (N_2359,In_2974,In_644);
xnor U2360 (N_2360,In_1019,In_2009);
nor U2361 (N_2361,In_2619,In_2314);
nand U2362 (N_2362,In_1109,In_2249);
and U2363 (N_2363,In_2746,In_2336);
xnor U2364 (N_2364,In_861,In_2090);
or U2365 (N_2365,In_1943,In_597);
and U2366 (N_2366,In_447,In_2081);
nand U2367 (N_2367,In_70,In_2483);
nand U2368 (N_2368,In_1746,In_2169);
nor U2369 (N_2369,In_277,In_2177);
or U2370 (N_2370,In_2056,In_2010);
and U2371 (N_2371,In_619,In_1386);
or U2372 (N_2372,In_1084,In_2810);
nand U2373 (N_2373,In_1156,In_1068);
nand U2374 (N_2374,In_463,In_1448);
nor U2375 (N_2375,In_2538,In_1058);
xnor U2376 (N_2376,In_928,In_1996);
nand U2377 (N_2377,In_983,In_2461);
or U2378 (N_2378,In_207,In_952);
nor U2379 (N_2379,In_2134,In_294);
nand U2380 (N_2380,In_1041,In_704);
and U2381 (N_2381,In_1755,In_261);
nor U2382 (N_2382,In_302,In_2614);
nand U2383 (N_2383,In_1782,In_550);
xnor U2384 (N_2384,In_112,In_1894);
or U2385 (N_2385,In_1234,In_2115);
nor U2386 (N_2386,In_759,In_2413);
xnor U2387 (N_2387,In_453,In_2038);
xnor U2388 (N_2388,In_1078,In_2532);
nor U2389 (N_2389,In_524,In_1753);
nand U2390 (N_2390,In_987,In_1780);
xnor U2391 (N_2391,In_2540,In_432);
nand U2392 (N_2392,In_600,In_1384);
nor U2393 (N_2393,In_500,In_1727);
or U2394 (N_2394,In_369,In_2924);
xnor U2395 (N_2395,In_1957,In_1934);
nand U2396 (N_2396,In_2742,In_1586);
xnor U2397 (N_2397,In_570,In_1912);
or U2398 (N_2398,In_2469,In_1456);
and U2399 (N_2399,In_20,In_2758);
nor U2400 (N_2400,In_1036,In_1722);
nand U2401 (N_2401,In_2379,In_351);
and U2402 (N_2402,In_1884,In_1620);
xnor U2403 (N_2403,In_1767,In_1964);
or U2404 (N_2404,In_2166,In_2197);
xnor U2405 (N_2405,In_1326,In_647);
xor U2406 (N_2406,In_2414,In_2174);
xor U2407 (N_2407,In_2366,In_2489);
or U2408 (N_2408,In_2417,In_441);
xor U2409 (N_2409,In_278,In_739);
xnor U2410 (N_2410,In_352,In_1939);
xor U2411 (N_2411,In_1683,In_2553);
xor U2412 (N_2412,In_125,In_2832);
and U2413 (N_2413,In_2585,In_105);
and U2414 (N_2414,In_1157,In_2246);
nand U2415 (N_2415,In_701,In_712);
or U2416 (N_2416,In_2195,In_1945);
xnor U2417 (N_2417,In_603,In_1395);
nor U2418 (N_2418,In_2535,In_1081);
or U2419 (N_2419,In_1197,In_1149);
or U2420 (N_2420,In_1022,In_1813);
nand U2421 (N_2421,In_2315,In_209);
nand U2422 (N_2422,In_1526,In_2987);
and U2423 (N_2423,In_2005,In_2622);
or U2424 (N_2424,In_2154,In_410);
nor U2425 (N_2425,In_2962,In_384);
nor U2426 (N_2426,In_2180,In_1518);
nor U2427 (N_2427,In_1084,In_2836);
or U2428 (N_2428,In_1163,In_1833);
or U2429 (N_2429,In_537,In_2040);
nor U2430 (N_2430,In_476,In_358);
or U2431 (N_2431,In_881,In_134);
nand U2432 (N_2432,In_1279,In_2495);
xor U2433 (N_2433,In_21,In_1565);
xor U2434 (N_2434,In_1052,In_2002);
nand U2435 (N_2435,In_1685,In_1938);
and U2436 (N_2436,In_2195,In_852);
nor U2437 (N_2437,In_2243,In_2902);
xor U2438 (N_2438,In_2245,In_2062);
xnor U2439 (N_2439,In_2965,In_1672);
and U2440 (N_2440,In_1394,In_1162);
nand U2441 (N_2441,In_1094,In_255);
and U2442 (N_2442,In_769,In_2407);
nand U2443 (N_2443,In_1118,In_2908);
or U2444 (N_2444,In_1354,In_924);
nor U2445 (N_2445,In_2734,In_1696);
xnor U2446 (N_2446,In_694,In_2030);
and U2447 (N_2447,In_2857,In_119);
xor U2448 (N_2448,In_2196,In_1791);
nor U2449 (N_2449,In_598,In_2381);
nand U2450 (N_2450,In_1473,In_1089);
nand U2451 (N_2451,In_2595,In_737);
or U2452 (N_2452,In_1193,In_1315);
or U2453 (N_2453,In_1585,In_2770);
or U2454 (N_2454,In_1356,In_625);
or U2455 (N_2455,In_1660,In_2609);
nor U2456 (N_2456,In_2508,In_2729);
xor U2457 (N_2457,In_1827,In_1272);
nor U2458 (N_2458,In_4,In_961);
nor U2459 (N_2459,In_82,In_728);
nor U2460 (N_2460,In_1434,In_1908);
and U2461 (N_2461,In_695,In_2806);
or U2462 (N_2462,In_2381,In_2919);
xnor U2463 (N_2463,In_2035,In_2305);
or U2464 (N_2464,In_738,In_441);
and U2465 (N_2465,In_19,In_769);
xnor U2466 (N_2466,In_2473,In_2618);
xnor U2467 (N_2467,In_710,In_1656);
and U2468 (N_2468,In_575,In_757);
nor U2469 (N_2469,In_1102,In_1624);
or U2470 (N_2470,In_817,In_305);
nand U2471 (N_2471,In_2389,In_76);
xor U2472 (N_2472,In_1267,In_2201);
xnor U2473 (N_2473,In_1945,In_2123);
or U2474 (N_2474,In_311,In_72);
nand U2475 (N_2475,In_810,In_1818);
xnor U2476 (N_2476,In_1168,In_2378);
and U2477 (N_2477,In_401,In_1717);
nor U2478 (N_2478,In_2500,In_1573);
nor U2479 (N_2479,In_717,In_548);
nand U2480 (N_2480,In_1690,In_836);
and U2481 (N_2481,In_2314,In_2893);
or U2482 (N_2482,In_602,In_725);
nand U2483 (N_2483,In_492,In_277);
nand U2484 (N_2484,In_277,In_2265);
xnor U2485 (N_2485,In_2929,In_276);
xnor U2486 (N_2486,In_2825,In_2522);
nor U2487 (N_2487,In_102,In_2275);
nor U2488 (N_2488,In_2262,In_168);
nor U2489 (N_2489,In_700,In_2310);
nand U2490 (N_2490,In_478,In_492);
nor U2491 (N_2491,In_1236,In_1430);
nand U2492 (N_2492,In_1312,In_263);
nor U2493 (N_2493,In_1713,In_2503);
xnor U2494 (N_2494,In_1933,In_180);
and U2495 (N_2495,In_1754,In_2358);
xor U2496 (N_2496,In_1273,In_305);
nand U2497 (N_2497,In_1755,In_1044);
xor U2498 (N_2498,In_1512,In_1655);
or U2499 (N_2499,In_2776,In_2918);
or U2500 (N_2500,In_2542,In_295);
nor U2501 (N_2501,In_2892,In_2326);
xor U2502 (N_2502,In_1007,In_249);
nand U2503 (N_2503,In_2259,In_1813);
nand U2504 (N_2504,In_2384,In_1446);
and U2505 (N_2505,In_1776,In_1737);
nor U2506 (N_2506,In_1817,In_693);
nor U2507 (N_2507,In_1795,In_2655);
and U2508 (N_2508,In_2140,In_1606);
xor U2509 (N_2509,In_75,In_2035);
nand U2510 (N_2510,In_632,In_2016);
and U2511 (N_2511,In_1016,In_2022);
or U2512 (N_2512,In_2236,In_1854);
xor U2513 (N_2513,In_1672,In_2624);
nand U2514 (N_2514,In_836,In_925);
nand U2515 (N_2515,In_1092,In_1942);
nor U2516 (N_2516,In_24,In_33);
nor U2517 (N_2517,In_1703,In_1319);
nand U2518 (N_2518,In_1548,In_1094);
xnor U2519 (N_2519,In_2398,In_1566);
xnor U2520 (N_2520,In_382,In_1063);
nand U2521 (N_2521,In_2966,In_2649);
nor U2522 (N_2522,In_50,In_2764);
and U2523 (N_2523,In_2362,In_1028);
nor U2524 (N_2524,In_1227,In_2456);
xnor U2525 (N_2525,In_1669,In_990);
or U2526 (N_2526,In_1242,In_520);
xor U2527 (N_2527,In_302,In_1854);
nand U2528 (N_2528,In_1789,In_1032);
xnor U2529 (N_2529,In_815,In_812);
nor U2530 (N_2530,In_1786,In_1085);
nor U2531 (N_2531,In_415,In_2014);
xnor U2532 (N_2532,In_2105,In_921);
or U2533 (N_2533,In_1484,In_1059);
nor U2534 (N_2534,In_1667,In_134);
xnor U2535 (N_2535,In_471,In_1127);
and U2536 (N_2536,In_2815,In_1687);
and U2537 (N_2537,In_1169,In_1858);
or U2538 (N_2538,In_1249,In_2553);
nand U2539 (N_2539,In_1147,In_1053);
nand U2540 (N_2540,In_1097,In_2882);
xnor U2541 (N_2541,In_1010,In_2266);
nor U2542 (N_2542,In_1559,In_2434);
xnor U2543 (N_2543,In_2976,In_2395);
or U2544 (N_2544,In_653,In_895);
and U2545 (N_2545,In_65,In_6);
or U2546 (N_2546,In_742,In_2532);
and U2547 (N_2547,In_2679,In_2518);
nand U2548 (N_2548,In_2266,In_787);
nand U2549 (N_2549,In_2530,In_2350);
nor U2550 (N_2550,In_154,In_2249);
nand U2551 (N_2551,In_1017,In_2256);
xnor U2552 (N_2552,In_1252,In_369);
or U2553 (N_2553,In_2541,In_2056);
nand U2554 (N_2554,In_153,In_2284);
nand U2555 (N_2555,In_2368,In_1569);
and U2556 (N_2556,In_2134,In_28);
and U2557 (N_2557,In_567,In_980);
nand U2558 (N_2558,In_2585,In_7);
nand U2559 (N_2559,In_490,In_1466);
or U2560 (N_2560,In_1887,In_282);
nor U2561 (N_2561,In_1859,In_2097);
xor U2562 (N_2562,In_1830,In_1374);
nand U2563 (N_2563,In_829,In_2299);
and U2564 (N_2564,In_2273,In_128);
and U2565 (N_2565,In_2859,In_582);
and U2566 (N_2566,In_1796,In_679);
or U2567 (N_2567,In_629,In_2059);
and U2568 (N_2568,In_455,In_316);
or U2569 (N_2569,In_1420,In_769);
nor U2570 (N_2570,In_368,In_576);
nor U2571 (N_2571,In_799,In_2848);
nor U2572 (N_2572,In_1691,In_31);
nand U2573 (N_2573,In_2820,In_365);
nand U2574 (N_2574,In_2574,In_1910);
nand U2575 (N_2575,In_350,In_846);
xnor U2576 (N_2576,In_336,In_503);
nor U2577 (N_2577,In_1339,In_2985);
nor U2578 (N_2578,In_1618,In_2628);
nand U2579 (N_2579,In_2919,In_1483);
and U2580 (N_2580,In_1284,In_1421);
and U2581 (N_2581,In_2723,In_264);
and U2582 (N_2582,In_1357,In_1796);
nand U2583 (N_2583,In_1310,In_1421);
and U2584 (N_2584,In_82,In_849);
and U2585 (N_2585,In_1035,In_2775);
and U2586 (N_2586,In_1541,In_1962);
or U2587 (N_2587,In_575,In_1644);
nor U2588 (N_2588,In_990,In_1656);
xnor U2589 (N_2589,In_1301,In_2937);
nor U2590 (N_2590,In_1745,In_1997);
and U2591 (N_2591,In_1883,In_2222);
and U2592 (N_2592,In_2425,In_1487);
nor U2593 (N_2593,In_2897,In_571);
nand U2594 (N_2594,In_1254,In_375);
nand U2595 (N_2595,In_1263,In_2124);
or U2596 (N_2596,In_160,In_1530);
or U2597 (N_2597,In_104,In_694);
xor U2598 (N_2598,In_561,In_1298);
xor U2599 (N_2599,In_1658,In_1810);
xor U2600 (N_2600,In_2865,In_2219);
and U2601 (N_2601,In_2418,In_69);
and U2602 (N_2602,In_618,In_2032);
nand U2603 (N_2603,In_1223,In_2552);
or U2604 (N_2604,In_1217,In_1401);
nand U2605 (N_2605,In_1349,In_2131);
nand U2606 (N_2606,In_1298,In_1070);
nor U2607 (N_2607,In_887,In_2082);
nor U2608 (N_2608,In_1946,In_1562);
nor U2609 (N_2609,In_1734,In_1639);
nor U2610 (N_2610,In_1362,In_511);
nor U2611 (N_2611,In_1915,In_1556);
nor U2612 (N_2612,In_2754,In_1208);
nor U2613 (N_2613,In_506,In_2881);
nor U2614 (N_2614,In_886,In_1568);
xor U2615 (N_2615,In_1736,In_24);
xor U2616 (N_2616,In_2046,In_676);
and U2617 (N_2617,In_534,In_1771);
nand U2618 (N_2618,In_1659,In_2328);
nand U2619 (N_2619,In_2914,In_2567);
nand U2620 (N_2620,In_1351,In_971);
or U2621 (N_2621,In_634,In_367);
and U2622 (N_2622,In_1014,In_310);
nor U2623 (N_2623,In_734,In_2854);
nor U2624 (N_2624,In_1105,In_2637);
and U2625 (N_2625,In_1970,In_545);
xor U2626 (N_2626,In_848,In_547);
or U2627 (N_2627,In_1419,In_1061);
xor U2628 (N_2628,In_1716,In_932);
nand U2629 (N_2629,In_1685,In_1389);
xor U2630 (N_2630,In_2470,In_1406);
or U2631 (N_2631,In_1276,In_2279);
and U2632 (N_2632,In_1995,In_1497);
and U2633 (N_2633,In_2017,In_2990);
xor U2634 (N_2634,In_2794,In_2616);
nand U2635 (N_2635,In_455,In_1770);
xnor U2636 (N_2636,In_2403,In_2500);
or U2637 (N_2637,In_604,In_510);
nor U2638 (N_2638,In_2327,In_348);
nand U2639 (N_2639,In_2926,In_1394);
or U2640 (N_2640,In_2594,In_514);
or U2641 (N_2641,In_1019,In_627);
xnor U2642 (N_2642,In_7,In_767);
or U2643 (N_2643,In_1225,In_44);
xor U2644 (N_2644,In_431,In_2013);
nor U2645 (N_2645,In_510,In_767);
xor U2646 (N_2646,In_2357,In_490);
nor U2647 (N_2647,In_1301,In_2585);
nand U2648 (N_2648,In_2603,In_2302);
or U2649 (N_2649,In_497,In_2569);
nor U2650 (N_2650,In_1992,In_2719);
nand U2651 (N_2651,In_1779,In_2040);
and U2652 (N_2652,In_1961,In_2443);
nand U2653 (N_2653,In_1826,In_1649);
nor U2654 (N_2654,In_1891,In_311);
nor U2655 (N_2655,In_982,In_2089);
nand U2656 (N_2656,In_367,In_2915);
and U2657 (N_2657,In_2144,In_592);
or U2658 (N_2658,In_110,In_2806);
nand U2659 (N_2659,In_1479,In_636);
xnor U2660 (N_2660,In_1686,In_2107);
or U2661 (N_2661,In_2593,In_1082);
or U2662 (N_2662,In_938,In_1730);
xnor U2663 (N_2663,In_996,In_1891);
nor U2664 (N_2664,In_935,In_2552);
nand U2665 (N_2665,In_2030,In_1758);
and U2666 (N_2666,In_2109,In_1266);
xor U2667 (N_2667,In_2442,In_1091);
xnor U2668 (N_2668,In_2056,In_440);
nor U2669 (N_2669,In_293,In_1401);
or U2670 (N_2670,In_308,In_568);
xnor U2671 (N_2671,In_2908,In_1663);
xor U2672 (N_2672,In_472,In_342);
or U2673 (N_2673,In_1023,In_2879);
nand U2674 (N_2674,In_1517,In_2065);
and U2675 (N_2675,In_1543,In_2792);
or U2676 (N_2676,In_1449,In_32);
nand U2677 (N_2677,In_2842,In_877);
and U2678 (N_2678,In_2134,In_1382);
and U2679 (N_2679,In_1640,In_2014);
or U2680 (N_2680,In_2599,In_2889);
nor U2681 (N_2681,In_1645,In_695);
nor U2682 (N_2682,In_2082,In_2404);
nand U2683 (N_2683,In_2598,In_1917);
and U2684 (N_2684,In_2423,In_121);
and U2685 (N_2685,In_1775,In_1997);
nor U2686 (N_2686,In_1931,In_1844);
and U2687 (N_2687,In_2116,In_1172);
xnor U2688 (N_2688,In_2675,In_1508);
nor U2689 (N_2689,In_461,In_1694);
and U2690 (N_2690,In_1046,In_1481);
xor U2691 (N_2691,In_321,In_289);
nand U2692 (N_2692,In_893,In_726);
nor U2693 (N_2693,In_2773,In_2150);
and U2694 (N_2694,In_1563,In_563);
or U2695 (N_2695,In_941,In_1175);
or U2696 (N_2696,In_2456,In_1366);
xor U2697 (N_2697,In_1385,In_1531);
nor U2698 (N_2698,In_2111,In_2546);
xor U2699 (N_2699,In_834,In_40);
nor U2700 (N_2700,In_2622,In_41);
xor U2701 (N_2701,In_2825,In_509);
nand U2702 (N_2702,In_509,In_1747);
xnor U2703 (N_2703,In_1298,In_915);
or U2704 (N_2704,In_1239,In_602);
nor U2705 (N_2705,In_1055,In_2967);
or U2706 (N_2706,In_2727,In_2554);
xnor U2707 (N_2707,In_2002,In_1727);
or U2708 (N_2708,In_1569,In_309);
or U2709 (N_2709,In_2078,In_131);
nor U2710 (N_2710,In_2461,In_604);
nor U2711 (N_2711,In_215,In_2999);
or U2712 (N_2712,In_2349,In_1165);
xor U2713 (N_2713,In_390,In_700);
nor U2714 (N_2714,In_2923,In_670);
nand U2715 (N_2715,In_1495,In_1022);
and U2716 (N_2716,In_176,In_2995);
xor U2717 (N_2717,In_262,In_2289);
nand U2718 (N_2718,In_1347,In_1461);
nand U2719 (N_2719,In_98,In_2371);
xor U2720 (N_2720,In_1404,In_2398);
and U2721 (N_2721,In_718,In_2714);
nor U2722 (N_2722,In_834,In_1872);
nand U2723 (N_2723,In_2392,In_309);
xnor U2724 (N_2724,In_1492,In_1009);
nor U2725 (N_2725,In_2761,In_191);
and U2726 (N_2726,In_1306,In_949);
nor U2727 (N_2727,In_141,In_404);
and U2728 (N_2728,In_1320,In_1285);
xnor U2729 (N_2729,In_2949,In_2190);
nand U2730 (N_2730,In_2336,In_664);
or U2731 (N_2731,In_1036,In_1768);
and U2732 (N_2732,In_2471,In_1849);
or U2733 (N_2733,In_130,In_881);
or U2734 (N_2734,In_34,In_1885);
xor U2735 (N_2735,In_1515,In_2140);
nor U2736 (N_2736,In_2853,In_1073);
and U2737 (N_2737,In_2098,In_2045);
nand U2738 (N_2738,In_2331,In_1358);
and U2739 (N_2739,In_708,In_193);
or U2740 (N_2740,In_2037,In_1074);
nand U2741 (N_2741,In_2085,In_1700);
nand U2742 (N_2742,In_2874,In_960);
nor U2743 (N_2743,In_2281,In_546);
or U2744 (N_2744,In_623,In_652);
nor U2745 (N_2745,In_2628,In_2099);
and U2746 (N_2746,In_692,In_1148);
nand U2747 (N_2747,In_2102,In_740);
and U2748 (N_2748,In_1031,In_1298);
nor U2749 (N_2749,In_249,In_2357);
or U2750 (N_2750,In_2263,In_2926);
or U2751 (N_2751,In_1305,In_2502);
and U2752 (N_2752,In_1926,In_1588);
and U2753 (N_2753,In_2402,In_1184);
nor U2754 (N_2754,In_2401,In_1982);
xnor U2755 (N_2755,In_908,In_2051);
nand U2756 (N_2756,In_1946,In_2334);
xor U2757 (N_2757,In_708,In_180);
and U2758 (N_2758,In_1126,In_1337);
and U2759 (N_2759,In_790,In_1629);
xnor U2760 (N_2760,In_1522,In_2262);
or U2761 (N_2761,In_963,In_2762);
nand U2762 (N_2762,In_1574,In_772);
nand U2763 (N_2763,In_2935,In_194);
nor U2764 (N_2764,In_626,In_1530);
nand U2765 (N_2765,In_2333,In_884);
xnor U2766 (N_2766,In_919,In_2082);
and U2767 (N_2767,In_2166,In_1523);
nand U2768 (N_2768,In_2164,In_1679);
or U2769 (N_2769,In_933,In_2889);
or U2770 (N_2770,In_750,In_2624);
xor U2771 (N_2771,In_1759,In_2776);
and U2772 (N_2772,In_1329,In_1289);
nor U2773 (N_2773,In_408,In_1503);
or U2774 (N_2774,In_2396,In_1971);
nor U2775 (N_2775,In_1852,In_1312);
and U2776 (N_2776,In_1133,In_1758);
nand U2777 (N_2777,In_1381,In_259);
nor U2778 (N_2778,In_885,In_1560);
xor U2779 (N_2779,In_2414,In_1352);
nor U2780 (N_2780,In_2670,In_1581);
xor U2781 (N_2781,In_20,In_974);
nor U2782 (N_2782,In_1346,In_2128);
and U2783 (N_2783,In_584,In_726);
and U2784 (N_2784,In_834,In_964);
or U2785 (N_2785,In_2576,In_2418);
xor U2786 (N_2786,In_1342,In_1270);
and U2787 (N_2787,In_2386,In_2932);
and U2788 (N_2788,In_1474,In_2724);
nor U2789 (N_2789,In_2331,In_955);
nor U2790 (N_2790,In_213,In_14);
nand U2791 (N_2791,In_2071,In_2305);
xnor U2792 (N_2792,In_1495,In_548);
and U2793 (N_2793,In_1718,In_1943);
nand U2794 (N_2794,In_1489,In_2363);
or U2795 (N_2795,In_723,In_2334);
xnor U2796 (N_2796,In_1929,In_2527);
or U2797 (N_2797,In_2313,In_2915);
nand U2798 (N_2798,In_910,In_1627);
nor U2799 (N_2799,In_2900,In_1635);
nand U2800 (N_2800,In_530,In_2646);
nor U2801 (N_2801,In_2166,In_279);
nand U2802 (N_2802,In_1420,In_1793);
or U2803 (N_2803,In_2906,In_2798);
and U2804 (N_2804,In_639,In_1594);
or U2805 (N_2805,In_194,In_509);
nand U2806 (N_2806,In_351,In_1340);
or U2807 (N_2807,In_1924,In_2516);
nor U2808 (N_2808,In_966,In_543);
and U2809 (N_2809,In_163,In_1477);
nand U2810 (N_2810,In_1122,In_1543);
nand U2811 (N_2811,In_2064,In_2933);
xor U2812 (N_2812,In_8,In_1403);
or U2813 (N_2813,In_520,In_2225);
or U2814 (N_2814,In_686,In_407);
or U2815 (N_2815,In_2431,In_2967);
nand U2816 (N_2816,In_1928,In_766);
and U2817 (N_2817,In_1459,In_949);
and U2818 (N_2818,In_1004,In_1844);
nor U2819 (N_2819,In_2402,In_2603);
or U2820 (N_2820,In_100,In_1033);
nand U2821 (N_2821,In_476,In_1454);
xnor U2822 (N_2822,In_197,In_303);
and U2823 (N_2823,In_2286,In_2392);
and U2824 (N_2824,In_1208,In_2731);
or U2825 (N_2825,In_2862,In_450);
nand U2826 (N_2826,In_2997,In_796);
xor U2827 (N_2827,In_587,In_228);
nand U2828 (N_2828,In_1201,In_1893);
or U2829 (N_2829,In_2729,In_2111);
nor U2830 (N_2830,In_1395,In_916);
nor U2831 (N_2831,In_1347,In_2577);
xnor U2832 (N_2832,In_1027,In_1676);
and U2833 (N_2833,In_2865,In_389);
or U2834 (N_2834,In_175,In_1427);
and U2835 (N_2835,In_1803,In_247);
nand U2836 (N_2836,In_236,In_233);
and U2837 (N_2837,In_2339,In_2913);
or U2838 (N_2838,In_988,In_2633);
and U2839 (N_2839,In_305,In_994);
or U2840 (N_2840,In_1454,In_2927);
nand U2841 (N_2841,In_1869,In_282);
xor U2842 (N_2842,In_446,In_576);
or U2843 (N_2843,In_2562,In_2363);
nand U2844 (N_2844,In_380,In_1329);
and U2845 (N_2845,In_320,In_1519);
nor U2846 (N_2846,In_2681,In_1668);
and U2847 (N_2847,In_234,In_2715);
xor U2848 (N_2848,In_1557,In_1676);
nand U2849 (N_2849,In_643,In_1726);
nor U2850 (N_2850,In_2813,In_2533);
nor U2851 (N_2851,In_2519,In_1184);
nor U2852 (N_2852,In_1471,In_2335);
xor U2853 (N_2853,In_808,In_2636);
or U2854 (N_2854,In_320,In_115);
nand U2855 (N_2855,In_129,In_2184);
and U2856 (N_2856,In_404,In_1757);
xor U2857 (N_2857,In_674,In_2362);
nand U2858 (N_2858,In_2847,In_551);
nand U2859 (N_2859,In_2581,In_2641);
or U2860 (N_2860,In_1602,In_2270);
nand U2861 (N_2861,In_784,In_1293);
nor U2862 (N_2862,In_399,In_304);
nor U2863 (N_2863,In_53,In_1409);
nor U2864 (N_2864,In_2269,In_92);
or U2865 (N_2865,In_393,In_966);
nor U2866 (N_2866,In_537,In_2529);
xnor U2867 (N_2867,In_659,In_449);
and U2868 (N_2868,In_2077,In_2405);
and U2869 (N_2869,In_1978,In_1412);
or U2870 (N_2870,In_2841,In_361);
or U2871 (N_2871,In_2676,In_422);
nor U2872 (N_2872,In_866,In_441);
or U2873 (N_2873,In_2139,In_1299);
nand U2874 (N_2874,In_1811,In_530);
and U2875 (N_2875,In_330,In_2314);
or U2876 (N_2876,In_1854,In_2633);
xnor U2877 (N_2877,In_1699,In_2352);
nand U2878 (N_2878,In_1246,In_2395);
xnor U2879 (N_2879,In_720,In_338);
nand U2880 (N_2880,In_2141,In_2179);
nor U2881 (N_2881,In_526,In_99);
or U2882 (N_2882,In_1081,In_2484);
xnor U2883 (N_2883,In_187,In_568);
nand U2884 (N_2884,In_232,In_2132);
and U2885 (N_2885,In_1566,In_2220);
or U2886 (N_2886,In_805,In_210);
nor U2887 (N_2887,In_169,In_286);
xor U2888 (N_2888,In_2726,In_582);
nand U2889 (N_2889,In_1956,In_1181);
nor U2890 (N_2890,In_2436,In_514);
xor U2891 (N_2891,In_763,In_2560);
or U2892 (N_2892,In_44,In_1506);
xnor U2893 (N_2893,In_2586,In_1370);
nand U2894 (N_2894,In_889,In_2090);
nor U2895 (N_2895,In_2600,In_788);
nor U2896 (N_2896,In_2866,In_2633);
or U2897 (N_2897,In_1801,In_160);
or U2898 (N_2898,In_185,In_1595);
or U2899 (N_2899,In_669,In_1489);
nor U2900 (N_2900,In_2749,In_2276);
or U2901 (N_2901,In_2329,In_384);
xor U2902 (N_2902,In_2233,In_1759);
and U2903 (N_2903,In_2653,In_2174);
or U2904 (N_2904,In_1956,In_223);
or U2905 (N_2905,In_885,In_349);
or U2906 (N_2906,In_1597,In_1410);
xnor U2907 (N_2907,In_2295,In_665);
and U2908 (N_2908,In_1961,In_2403);
nand U2909 (N_2909,In_1352,In_415);
nor U2910 (N_2910,In_1338,In_1476);
or U2911 (N_2911,In_1968,In_2113);
nor U2912 (N_2912,In_1976,In_679);
and U2913 (N_2913,In_1421,In_421);
or U2914 (N_2914,In_2495,In_2258);
nor U2915 (N_2915,In_2682,In_1880);
nor U2916 (N_2916,In_2824,In_2899);
xnor U2917 (N_2917,In_1700,In_2907);
or U2918 (N_2918,In_95,In_619);
nor U2919 (N_2919,In_31,In_1266);
nand U2920 (N_2920,In_113,In_2894);
xnor U2921 (N_2921,In_133,In_2307);
nand U2922 (N_2922,In_1663,In_1483);
and U2923 (N_2923,In_2406,In_2984);
xor U2924 (N_2924,In_34,In_1336);
xnor U2925 (N_2925,In_969,In_821);
nand U2926 (N_2926,In_1491,In_293);
nand U2927 (N_2927,In_1460,In_732);
and U2928 (N_2928,In_1013,In_901);
nor U2929 (N_2929,In_2111,In_1246);
nor U2930 (N_2930,In_1809,In_528);
nor U2931 (N_2931,In_1446,In_168);
xor U2932 (N_2932,In_80,In_745);
or U2933 (N_2933,In_2705,In_1502);
or U2934 (N_2934,In_390,In_686);
nand U2935 (N_2935,In_2511,In_723);
or U2936 (N_2936,In_1743,In_274);
nand U2937 (N_2937,In_547,In_330);
nand U2938 (N_2938,In_1003,In_880);
xor U2939 (N_2939,In_2946,In_2156);
nand U2940 (N_2940,In_1336,In_97);
and U2941 (N_2941,In_106,In_269);
xnor U2942 (N_2942,In_2527,In_2919);
xor U2943 (N_2943,In_496,In_2041);
nand U2944 (N_2944,In_1050,In_1702);
nand U2945 (N_2945,In_1011,In_2771);
and U2946 (N_2946,In_800,In_1660);
or U2947 (N_2947,In_2298,In_1814);
nor U2948 (N_2948,In_1872,In_2611);
and U2949 (N_2949,In_678,In_2726);
or U2950 (N_2950,In_2135,In_587);
nand U2951 (N_2951,In_2254,In_145);
nor U2952 (N_2952,In_240,In_943);
nand U2953 (N_2953,In_427,In_1574);
and U2954 (N_2954,In_2384,In_1747);
nand U2955 (N_2955,In_772,In_138);
and U2956 (N_2956,In_409,In_1410);
or U2957 (N_2957,In_1282,In_1468);
nor U2958 (N_2958,In_243,In_1713);
or U2959 (N_2959,In_2358,In_1083);
and U2960 (N_2960,In_1327,In_2521);
xnor U2961 (N_2961,In_1552,In_62);
or U2962 (N_2962,In_1095,In_60);
xnor U2963 (N_2963,In_1820,In_1399);
xnor U2964 (N_2964,In_235,In_2355);
nand U2965 (N_2965,In_563,In_2801);
and U2966 (N_2966,In_1953,In_2423);
or U2967 (N_2967,In_1666,In_881);
nand U2968 (N_2968,In_2649,In_2384);
and U2969 (N_2969,In_15,In_252);
nor U2970 (N_2970,In_2561,In_2839);
and U2971 (N_2971,In_1670,In_257);
xor U2972 (N_2972,In_2576,In_208);
or U2973 (N_2973,In_2272,In_2257);
nor U2974 (N_2974,In_785,In_2910);
and U2975 (N_2975,In_1278,In_1742);
and U2976 (N_2976,In_1077,In_2973);
or U2977 (N_2977,In_2001,In_1635);
xnor U2978 (N_2978,In_2094,In_1539);
xnor U2979 (N_2979,In_1557,In_2211);
and U2980 (N_2980,In_2276,In_293);
nand U2981 (N_2981,In_1041,In_431);
nor U2982 (N_2982,In_1587,In_1844);
and U2983 (N_2983,In_659,In_2461);
and U2984 (N_2984,In_1156,In_2022);
nor U2985 (N_2985,In_1348,In_661);
and U2986 (N_2986,In_1671,In_2149);
nand U2987 (N_2987,In_2919,In_2813);
and U2988 (N_2988,In_888,In_722);
and U2989 (N_2989,In_436,In_414);
xnor U2990 (N_2990,In_615,In_2859);
xnor U2991 (N_2991,In_2328,In_2335);
nor U2992 (N_2992,In_2517,In_204);
nor U2993 (N_2993,In_646,In_1276);
nor U2994 (N_2994,In_2333,In_172);
nor U2995 (N_2995,In_597,In_2455);
nand U2996 (N_2996,In_1865,In_2595);
or U2997 (N_2997,In_1779,In_895);
nor U2998 (N_2998,In_166,In_14);
nand U2999 (N_2999,In_1860,In_1133);
and U3000 (N_3000,In_1974,In_1180);
nand U3001 (N_3001,In_427,In_811);
and U3002 (N_3002,In_1483,In_2610);
xor U3003 (N_3003,In_697,In_1484);
xor U3004 (N_3004,In_1210,In_2921);
nand U3005 (N_3005,In_1954,In_2410);
and U3006 (N_3006,In_1768,In_69);
or U3007 (N_3007,In_929,In_1745);
nor U3008 (N_3008,In_699,In_388);
or U3009 (N_3009,In_2477,In_1349);
and U3010 (N_3010,In_744,In_977);
nor U3011 (N_3011,In_2238,In_2644);
and U3012 (N_3012,In_165,In_607);
nand U3013 (N_3013,In_863,In_2384);
nand U3014 (N_3014,In_2174,In_1989);
and U3015 (N_3015,In_1684,In_2881);
xnor U3016 (N_3016,In_2566,In_2058);
nand U3017 (N_3017,In_1715,In_1648);
xnor U3018 (N_3018,In_1027,In_45);
and U3019 (N_3019,In_1326,In_719);
nor U3020 (N_3020,In_1976,In_1155);
xnor U3021 (N_3021,In_2376,In_2453);
and U3022 (N_3022,In_2048,In_2092);
or U3023 (N_3023,In_2544,In_2467);
xor U3024 (N_3024,In_2892,In_1733);
and U3025 (N_3025,In_1318,In_542);
nand U3026 (N_3026,In_167,In_291);
or U3027 (N_3027,In_2663,In_1830);
nor U3028 (N_3028,In_268,In_2274);
nand U3029 (N_3029,In_1823,In_821);
xnor U3030 (N_3030,In_1515,In_234);
nand U3031 (N_3031,In_910,In_2240);
nor U3032 (N_3032,In_1633,In_1173);
nor U3033 (N_3033,In_58,In_1576);
and U3034 (N_3034,In_2592,In_165);
nor U3035 (N_3035,In_1950,In_436);
and U3036 (N_3036,In_2263,In_1571);
nor U3037 (N_3037,In_2062,In_884);
or U3038 (N_3038,In_1292,In_836);
nor U3039 (N_3039,In_113,In_1243);
nand U3040 (N_3040,In_300,In_1018);
xor U3041 (N_3041,In_52,In_904);
nand U3042 (N_3042,In_90,In_920);
nor U3043 (N_3043,In_184,In_1109);
nand U3044 (N_3044,In_2380,In_1524);
or U3045 (N_3045,In_199,In_469);
and U3046 (N_3046,In_2363,In_1075);
nand U3047 (N_3047,In_2885,In_330);
and U3048 (N_3048,In_2162,In_2276);
nor U3049 (N_3049,In_1527,In_46);
and U3050 (N_3050,In_2962,In_2692);
or U3051 (N_3051,In_535,In_2076);
nor U3052 (N_3052,In_2018,In_1530);
nand U3053 (N_3053,In_1109,In_1330);
nor U3054 (N_3054,In_2427,In_2691);
nand U3055 (N_3055,In_120,In_869);
and U3056 (N_3056,In_2938,In_1451);
and U3057 (N_3057,In_1628,In_2574);
nor U3058 (N_3058,In_2123,In_2506);
or U3059 (N_3059,In_2131,In_2018);
nor U3060 (N_3060,In_2714,In_746);
or U3061 (N_3061,In_1251,In_269);
nor U3062 (N_3062,In_1716,In_2133);
nor U3063 (N_3063,In_633,In_75);
nand U3064 (N_3064,In_201,In_121);
and U3065 (N_3065,In_194,In_2669);
nor U3066 (N_3066,In_878,In_1079);
xnor U3067 (N_3067,In_2476,In_1898);
xor U3068 (N_3068,In_344,In_1364);
nor U3069 (N_3069,In_2631,In_897);
and U3070 (N_3070,In_777,In_126);
and U3071 (N_3071,In_2938,In_1153);
xnor U3072 (N_3072,In_2535,In_913);
or U3073 (N_3073,In_1096,In_1672);
nor U3074 (N_3074,In_1504,In_138);
or U3075 (N_3075,In_1744,In_463);
xor U3076 (N_3076,In_387,In_1739);
and U3077 (N_3077,In_806,In_2544);
or U3078 (N_3078,In_2239,In_886);
nand U3079 (N_3079,In_2130,In_2290);
xor U3080 (N_3080,In_484,In_595);
or U3081 (N_3081,In_2141,In_2880);
xor U3082 (N_3082,In_2036,In_603);
and U3083 (N_3083,In_691,In_2414);
and U3084 (N_3084,In_2386,In_2211);
nand U3085 (N_3085,In_1359,In_1756);
nor U3086 (N_3086,In_605,In_1477);
nor U3087 (N_3087,In_2618,In_1013);
or U3088 (N_3088,In_2162,In_2963);
or U3089 (N_3089,In_1004,In_1424);
nand U3090 (N_3090,In_769,In_1409);
or U3091 (N_3091,In_870,In_2164);
nor U3092 (N_3092,In_217,In_2978);
and U3093 (N_3093,In_195,In_1401);
xnor U3094 (N_3094,In_2659,In_1184);
or U3095 (N_3095,In_785,In_2405);
and U3096 (N_3096,In_2146,In_973);
and U3097 (N_3097,In_1019,In_471);
or U3098 (N_3098,In_613,In_2392);
nor U3099 (N_3099,In_2069,In_2110);
or U3100 (N_3100,In_1661,In_1043);
and U3101 (N_3101,In_1031,In_1877);
or U3102 (N_3102,In_2255,In_1210);
nand U3103 (N_3103,In_1683,In_2351);
nand U3104 (N_3104,In_513,In_1539);
nor U3105 (N_3105,In_1850,In_489);
xnor U3106 (N_3106,In_2013,In_284);
xnor U3107 (N_3107,In_2818,In_2587);
nor U3108 (N_3108,In_1326,In_1002);
xor U3109 (N_3109,In_1464,In_189);
or U3110 (N_3110,In_1089,In_309);
and U3111 (N_3111,In_1062,In_1021);
nand U3112 (N_3112,In_1736,In_1037);
and U3113 (N_3113,In_1906,In_2525);
nand U3114 (N_3114,In_586,In_2838);
nand U3115 (N_3115,In_1900,In_1243);
nand U3116 (N_3116,In_1061,In_1611);
xor U3117 (N_3117,In_1201,In_2525);
or U3118 (N_3118,In_820,In_513);
xnor U3119 (N_3119,In_2141,In_1404);
or U3120 (N_3120,In_729,In_2576);
and U3121 (N_3121,In_791,In_1364);
xor U3122 (N_3122,In_912,In_774);
or U3123 (N_3123,In_1009,In_532);
or U3124 (N_3124,In_1427,In_2316);
and U3125 (N_3125,In_1826,In_2551);
nor U3126 (N_3126,In_1592,In_2969);
and U3127 (N_3127,In_859,In_552);
xor U3128 (N_3128,In_2418,In_661);
nor U3129 (N_3129,In_1773,In_2560);
nand U3130 (N_3130,In_122,In_1802);
and U3131 (N_3131,In_1731,In_1013);
nand U3132 (N_3132,In_2558,In_487);
xor U3133 (N_3133,In_200,In_497);
nand U3134 (N_3134,In_902,In_1739);
nand U3135 (N_3135,In_2332,In_277);
or U3136 (N_3136,In_715,In_2243);
nand U3137 (N_3137,In_1122,In_235);
xor U3138 (N_3138,In_591,In_1547);
nand U3139 (N_3139,In_2764,In_1849);
or U3140 (N_3140,In_1200,In_2113);
xnor U3141 (N_3141,In_2338,In_511);
and U3142 (N_3142,In_1458,In_2989);
nor U3143 (N_3143,In_2740,In_914);
xnor U3144 (N_3144,In_998,In_1540);
and U3145 (N_3145,In_852,In_2622);
xor U3146 (N_3146,In_1353,In_2078);
or U3147 (N_3147,In_1208,In_100);
or U3148 (N_3148,In_1924,In_1874);
and U3149 (N_3149,In_734,In_1072);
or U3150 (N_3150,In_2076,In_778);
or U3151 (N_3151,In_1296,In_807);
xnor U3152 (N_3152,In_1585,In_2038);
or U3153 (N_3153,In_674,In_1161);
or U3154 (N_3154,In_2148,In_1002);
or U3155 (N_3155,In_686,In_964);
nand U3156 (N_3156,In_2861,In_2128);
or U3157 (N_3157,In_2124,In_2699);
nor U3158 (N_3158,In_1391,In_789);
nand U3159 (N_3159,In_1745,In_2718);
or U3160 (N_3160,In_1818,In_414);
or U3161 (N_3161,In_167,In_2793);
nand U3162 (N_3162,In_1334,In_957);
or U3163 (N_3163,In_142,In_547);
or U3164 (N_3164,In_435,In_2633);
xnor U3165 (N_3165,In_1906,In_1619);
xor U3166 (N_3166,In_2221,In_1180);
and U3167 (N_3167,In_2506,In_2818);
xor U3168 (N_3168,In_2453,In_2467);
and U3169 (N_3169,In_148,In_3);
xnor U3170 (N_3170,In_2754,In_2685);
nor U3171 (N_3171,In_1399,In_2221);
and U3172 (N_3172,In_1786,In_368);
or U3173 (N_3173,In_2936,In_501);
nor U3174 (N_3174,In_2868,In_1115);
nand U3175 (N_3175,In_1653,In_2302);
xnor U3176 (N_3176,In_2762,In_1797);
xnor U3177 (N_3177,In_135,In_217);
nor U3178 (N_3178,In_1448,In_1718);
xor U3179 (N_3179,In_2587,In_1907);
and U3180 (N_3180,In_1539,In_2064);
or U3181 (N_3181,In_803,In_2778);
nor U3182 (N_3182,In_2627,In_2606);
nand U3183 (N_3183,In_1037,In_2695);
nor U3184 (N_3184,In_2874,In_115);
or U3185 (N_3185,In_2702,In_1132);
or U3186 (N_3186,In_146,In_883);
xor U3187 (N_3187,In_1114,In_447);
and U3188 (N_3188,In_673,In_889);
or U3189 (N_3189,In_1445,In_2058);
nor U3190 (N_3190,In_1876,In_1277);
xor U3191 (N_3191,In_827,In_654);
nand U3192 (N_3192,In_2801,In_703);
or U3193 (N_3193,In_2956,In_717);
nor U3194 (N_3194,In_2989,In_1224);
or U3195 (N_3195,In_311,In_2611);
or U3196 (N_3196,In_1877,In_436);
or U3197 (N_3197,In_1433,In_386);
xor U3198 (N_3198,In_76,In_1404);
nand U3199 (N_3199,In_2490,In_40);
or U3200 (N_3200,In_1611,In_1526);
xnor U3201 (N_3201,In_617,In_2702);
xor U3202 (N_3202,In_2166,In_669);
xor U3203 (N_3203,In_2375,In_3);
nor U3204 (N_3204,In_1369,In_2083);
nor U3205 (N_3205,In_290,In_2140);
or U3206 (N_3206,In_2305,In_366);
nor U3207 (N_3207,In_2983,In_2788);
and U3208 (N_3208,In_1919,In_291);
xnor U3209 (N_3209,In_2948,In_1265);
nor U3210 (N_3210,In_569,In_1353);
xnor U3211 (N_3211,In_2739,In_2112);
or U3212 (N_3212,In_1122,In_1793);
nor U3213 (N_3213,In_978,In_264);
or U3214 (N_3214,In_1165,In_730);
or U3215 (N_3215,In_2463,In_1164);
or U3216 (N_3216,In_2142,In_1391);
nand U3217 (N_3217,In_2958,In_1690);
or U3218 (N_3218,In_450,In_2340);
nand U3219 (N_3219,In_1051,In_1705);
and U3220 (N_3220,In_132,In_470);
nand U3221 (N_3221,In_876,In_1202);
nand U3222 (N_3222,In_2356,In_2629);
and U3223 (N_3223,In_346,In_2301);
nor U3224 (N_3224,In_426,In_1942);
and U3225 (N_3225,In_2012,In_1535);
and U3226 (N_3226,In_1626,In_1521);
xor U3227 (N_3227,In_1756,In_1175);
and U3228 (N_3228,In_1994,In_1279);
nor U3229 (N_3229,In_546,In_1863);
nand U3230 (N_3230,In_1036,In_2187);
xor U3231 (N_3231,In_2971,In_1880);
nor U3232 (N_3232,In_987,In_1946);
nor U3233 (N_3233,In_2127,In_1604);
or U3234 (N_3234,In_2197,In_1824);
and U3235 (N_3235,In_1020,In_364);
xnor U3236 (N_3236,In_2208,In_1512);
xnor U3237 (N_3237,In_1416,In_1420);
nand U3238 (N_3238,In_327,In_1225);
and U3239 (N_3239,In_551,In_80);
or U3240 (N_3240,In_645,In_2410);
or U3241 (N_3241,In_1080,In_2085);
nand U3242 (N_3242,In_1509,In_2991);
xnor U3243 (N_3243,In_2476,In_475);
nand U3244 (N_3244,In_1570,In_2209);
nand U3245 (N_3245,In_1038,In_2303);
xnor U3246 (N_3246,In_2287,In_676);
nand U3247 (N_3247,In_174,In_1406);
nor U3248 (N_3248,In_611,In_2642);
and U3249 (N_3249,In_1777,In_739);
or U3250 (N_3250,In_1521,In_185);
xor U3251 (N_3251,In_462,In_2473);
and U3252 (N_3252,In_1862,In_1314);
xor U3253 (N_3253,In_2260,In_2693);
nor U3254 (N_3254,In_1400,In_2820);
and U3255 (N_3255,In_1922,In_2127);
and U3256 (N_3256,In_2840,In_1992);
nor U3257 (N_3257,In_457,In_715);
and U3258 (N_3258,In_179,In_707);
xnor U3259 (N_3259,In_954,In_2749);
and U3260 (N_3260,In_2265,In_1470);
nor U3261 (N_3261,In_821,In_1921);
nor U3262 (N_3262,In_2163,In_2338);
xnor U3263 (N_3263,In_1930,In_35);
nor U3264 (N_3264,In_1229,In_2671);
nand U3265 (N_3265,In_1814,In_1399);
and U3266 (N_3266,In_25,In_302);
and U3267 (N_3267,In_1140,In_1723);
and U3268 (N_3268,In_2280,In_915);
nand U3269 (N_3269,In_1486,In_2269);
nor U3270 (N_3270,In_603,In_2750);
and U3271 (N_3271,In_1299,In_862);
and U3272 (N_3272,In_1762,In_2117);
and U3273 (N_3273,In_2906,In_628);
nand U3274 (N_3274,In_582,In_836);
and U3275 (N_3275,In_1079,In_465);
nand U3276 (N_3276,In_2659,In_690);
xnor U3277 (N_3277,In_839,In_605);
nor U3278 (N_3278,In_1931,In_1979);
xnor U3279 (N_3279,In_1357,In_1949);
nand U3280 (N_3280,In_2775,In_317);
xnor U3281 (N_3281,In_1684,In_1184);
nand U3282 (N_3282,In_495,In_1164);
xor U3283 (N_3283,In_1752,In_1618);
and U3284 (N_3284,In_2233,In_2334);
or U3285 (N_3285,In_1279,In_1194);
and U3286 (N_3286,In_1562,In_695);
and U3287 (N_3287,In_1406,In_1393);
xor U3288 (N_3288,In_292,In_2037);
xnor U3289 (N_3289,In_2495,In_2711);
nor U3290 (N_3290,In_2311,In_769);
nor U3291 (N_3291,In_1286,In_1847);
and U3292 (N_3292,In_364,In_933);
and U3293 (N_3293,In_1892,In_2794);
or U3294 (N_3294,In_441,In_2772);
and U3295 (N_3295,In_2701,In_1128);
nor U3296 (N_3296,In_527,In_2731);
or U3297 (N_3297,In_1979,In_375);
nor U3298 (N_3298,In_2532,In_1727);
nor U3299 (N_3299,In_2926,In_2465);
nor U3300 (N_3300,In_556,In_2519);
and U3301 (N_3301,In_2582,In_2279);
xor U3302 (N_3302,In_2338,In_1117);
xnor U3303 (N_3303,In_2438,In_1777);
nor U3304 (N_3304,In_495,In_734);
nand U3305 (N_3305,In_1697,In_2460);
nor U3306 (N_3306,In_2586,In_499);
and U3307 (N_3307,In_835,In_1507);
and U3308 (N_3308,In_931,In_2508);
xnor U3309 (N_3309,In_387,In_2733);
or U3310 (N_3310,In_570,In_2608);
nor U3311 (N_3311,In_437,In_635);
nand U3312 (N_3312,In_2183,In_1856);
nand U3313 (N_3313,In_2906,In_172);
nor U3314 (N_3314,In_992,In_601);
nand U3315 (N_3315,In_394,In_1482);
and U3316 (N_3316,In_245,In_180);
nor U3317 (N_3317,In_2495,In_1383);
nand U3318 (N_3318,In_1554,In_489);
xor U3319 (N_3319,In_480,In_1910);
or U3320 (N_3320,In_2499,In_2101);
xnor U3321 (N_3321,In_2101,In_2955);
nand U3322 (N_3322,In_2996,In_987);
and U3323 (N_3323,In_935,In_2017);
or U3324 (N_3324,In_2573,In_2572);
xnor U3325 (N_3325,In_2131,In_608);
and U3326 (N_3326,In_1179,In_1489);
or U3327 (N_3327,In_484,In_2142);
nor U3328 (N_3328,In_1601,In_949);
xor U3329 (N_3329,In_228,In_2443);
xor U3330 (N_3330,In_1661,In_882);
and U3331 (N_3331,In_1890,In_2496);
xnor U3332 (N_3332,In_538,In_2778);
nand U3333 (N_3333,In_1644,In_2408);
nor U3334 (N_3334,In_714,In_1830);
xnor U3335 (N_3335,In_2993,In_1723);
nand U3336 (N_3336,In_2807,In_2070);
xnor U3337 (N_3337,In_2707,In_2592);
nand U3338 (N_3338,In_2170,In_813);
nor U3339 (N_3339,In_1532,In_2912);
or U3340 (N_3340,In_2301,In_2919);
nand U3341 (N_3341,In_286,In_185);
or U3342 (N_3342,In_2678,In_1665);
xor U3343 (N_3343,In_123,In_2842);
or U3344 (N_3344,In_2124,In_2453);
nor U3345 (N_3345,In_1413,In_2348);
and U3346 (N_3346,In_2650,In_427);
and U3347 (N_3347,In_1015,In_784);
xor U3348 (N_3348,In_354,In_2947);
xor U3349 (N_3349,In_2145,In_2687);
nor U3350 (N_3350,In_1779,In_2270);
nand U3351 (N_3351,In_1256,In_538);
xnor U3352 (N_3352,In_2590,In_1986);
nor U3353 (N_3353,In_2854,In_1220);
nand U3354 (N_3354,In_2767,In_1975);
xnor U3355 (N_3355,In_721,In_2970);
nor U3356 (N_3356,In_774,In_638);
and U3357 (N_3357,In_552,In_1476);
nand U3358 (N_3358,In_1389,In_1807);
and U3359 (N_3359,In_875,In_645);
or U3360 (N_3360,In_1300,In_608);
xor U3361 (N_3361,In_2986,In_1171);
xnor U3362 (N_3362,In_1500,In_804);
and U3363 (N_3363,In_205,In_2589);
nor U3364 (N_3364,In_830,In_607);
nor U3365 (N_3365,In_1100,In_270);
nand U3366 (N_3366,In_2633,In_2086);
nand U3367 (N_3367,In_868,In_2945);
nand U3368 (N_3368,In_2778,In_1329);
nor U3369 (N_3369,In_2402,In_1273);
nand U3370 (N_3370,In_661,In_1705);
and U3371 (N_3371,In_128,In_1771);
nor U3372 (N_3372,In_2693,In_1444);
nor U3373 (N_3373,In_1485,In_324);
nor U3374 (N_3374,In_1867,In_2684);
nand U3375 (N_3375,In_2500,In_508);
xnor U3376 (N_3376,In_614,In_1807);
and U3377 (N_3377,In_883,In_2375);
or U3378 (N_3378,In_2328,In_240);
xnor U3379 (N_3379,In_2430,In_1767);
or U3380 (N_3380,In_1746,In_2379);
or U3381 (N_3381,In_1772,In_2579);
or U3382 (N_3382,In_745,In_2310);
nor U3383 (N_3383,In_2488,In_2459);
nand U3384 (N_3384,In_163,In_990);
nand U3385 (N_3385,In_159,In_502);
and U3386 (N_3386,In_2894,In_981);
nand U3387 (N_3387,In_821,In_1272);
xor U3388 (N_3388,In_2387,In_1956);
nor U3389 (N_3389,In_1560,In_2019);
nand U3390 (N_3390,In_471,In_773);
and U3391 (N_3391,In_577,In_85);
nand U3392 (N_3392,In_2655,In_460);
nand U3393 (N_3393,In_2621,In_1532);
nand U3394 (N_3394,In_212,In_1936);
and U3395 (N_3395,In_1731,In_1432);
nand U3396 (N_3396,In_217,In_1268);
nand U3397 (N_3397,In_2908,In_1760);
or U3398 (N_3398,In_2322,In_664);
xor U3399 (N_3399,In_823,In_319);
and U3400 (N_3400,In_154,In_899);
and U3401 (N_3401,In_289,In_37);
xnor U3402 (N_3402,In_442,In_400);
xor U3403 (N_3403,In_339,In_1086);
nand U3404 (N_3404,In_1363,In_827);
nand U3405 (N_3405,In_2323,In_302);
xor U3406 (N_3406,In_362,In_869);
nand U3407 (N_3407,In_164,In_2189);
nand U3408 (N_3408,In_2565,In_1475);
xnor U3409 (N_3409,In_1681,In_1049);
xor U3410 (N_3410,In_1671,In_1668);
xor U3411 (N_3411,In_72,In_2143);
xor U3412 (N_3412,In_1892,In_1737);
nor U3413 (N_3413,In_1230,In_1656);
xnor U3414 (N_3414,In_2638,In_1123);
or U3415 (N_3415,In_2545,In_2107);
or U3416 (N_3416,In_2957,In_775);
and U3417 (N_3417,In_2411,In_2820);
and U3418 (N_3418,In_647,In_1874);
and U3419 (N_3419,In_1062,In_2209);
nand U3420 (N_3420,In_94,In_762);
or U3421 (N_3421,In_1318,In_813);
or U3422 (N_3422,In_1058,In_1229);
xnor U3423 (N_3423,In_775,In_2718);
and U3424 (N_3424,In_2408,In_205);
and U3425 (N_3425,In_2077,In_2059);
nand U3426 (N_3426,In_242,In_1666);
or U3427 (N_3427,In_391,In_2159);
or U3428 (N_3428,In_2068,In_438);
xnor U3429 (N_3429,In_1358,In_2409);
nor U3430 (N_3430,In_298,In_951);
nor U3431 (N_3431,In_880,In_1494);
nand U3432 (N_3432,In_81,In_531);
nand U3433 (N_3433,In_1996,In_345);
nand U3434 (N_3434,In_1122,In_1917);
nand U3435 (N_3435,In_1477,In_12);
xor U3436 (N_3436,In_2794,In_400);
xnor U3437 (N_3437,In_1357,In_641);
and U3438 (N_3438,In_269,In_1216);
xor U3439 (N_3439,In_1512,In_1060);
xnor U3440 (N_3440,In_529,In_2887);
or U3441 (N_3441,In_692,In_484);
and U3442 (N_3442,In_1396,In_2607);
or U3443 (N_3443,In_1998,In_2000);
or U3444 (N_3444,In_315,In_2881);
nand U3445 (N_3445,In_1865,In_2571);
xnor U3446 (N_3446,In_2564,In_2302);
nor U3447 (N_3447,In_2562,In_2966);
xnor U3448 (N_3448,In_542,In_582);
and U3449 (N_3449,In_1717,In_1006);
nor U3450 (N_3450,In_289,In_821);
nor U3451 (N_3451,In_2309,In_346);
and U3452 (N_3452,In_743,In_1392);
nor U3453 (N_3453,In_2629,In_1753);
nor U3454 (N_3454,In_2420,In_580);
xor U3455 (N_3455,In_1172,In_1628);
nor U3456 (N_3456,In_1451,In_1778);
xor U3457 (N_3457,In_2973,In_1534);
nand U3458 (N_3458,In_2390,In_1446);
or U3459 (N_3459,In_843,In_1690);
and U3460 (N_3460,In_933,In_221);
and U3461 (N_3461,In_351,In_1992);
nand U3462 (N_3462,In_912,In_2435);
xor U3463 (N_3463,In_2460,In_1009);
and U3464 (N_3464,In_457,In_513);
or U3465 (N_3465,In_2268,In_2894);
nand U3466 (N_3466,In_409,In_240);
nand U3467 (N_3467,In_1088,In_1086);
xor U3468 (N_3468,In_2612,In_2148);
or U3469 (N_3469,In_2760,In_1229);
or U3470 (N_3470,In_2105,In_2185);
and U3471 (N_3471,In_1177,In_52);
and U3472 (N_3472,In_159,In_2004);
or U3473 (N_3473,In_1996,In_854);
and U3474 (N_3474,In_1351,In_758);
or U3475 (N_3475,In_605,In_2620);
nor U3476 (N_3476,In_339,In_292);
and U3477 (N_3477,In_1002,In_2441);
or U3478 (N_3478,In_1677,In_294);
nand U3479 (N_3479,In_1396,In_2519);
xnor U3480 (N_3480,In_1580,In_75);
and U3481 (N_3481,In_1916,In_1642);
or U3482 (N_3482,In_2159,In_907);
nand U3483 (N_3483,In_942,In_1298);
nand U3484 (N_3484,In_360,In_850);
or U3485 (N_3485,In_2067,In_1673);
xnor U3486 (N_3486,In_1300,In_2048);
xnor U3487 (N_3487,In_2665,In_719);
nor U3488 (N_3488,In_1227,In_957);
and U3489 (N_3489,In_2099,In_1779);
nor U3490 (N_3490,In_328,In_2361);
and U3491 (N_3491,In_2566,In_1565);
nand U3492 (N_3492,In_2459,In_793);
nand U3493 (N_3493,In_2304,In_2476);
nor U3494 (N_3494,In_2352,In_1853);
xnor U3495 (N_3495,In_2199,In_2331);
or U3496 (N_3496,In_819,In_1772);
or U3497 (N_3497,In_947,In_1911);
xor U3498 (N_3498,In_2930,In_1104);
or U3499 (N_3499,In_2533,In_1432);
nor U3500 (N_3500,In_164,In_1706);
nor U3501 (N_3501,In_2987,In_1048);
or U3502 (N_3502,In_1052,In_1446);
or U3503 (N_3503,In_129,In_1174);
or U3504 (N_3504,In_2341,In_483);
and U3505 (N_3505,In_1000,In_1260);
and U3506 (N_3506,In_780,In_350);
and U3507 (N_3507,In_2388,In_201);
xor U3508 (N_3508,In_2376,In_777);
and U3509 (N_3509,In_1625,In_545);
nor U3510 (N_3510,In_564,In_2693);
nor U3511 (N_3511,In_1289,In_2975);
and U3512 (N_3512,In_97,In_1395);
nand U3513 (N_3513,In_1639,In_1318);
xnor U3514 (N_3514,In_819,In_2779);
xor U3515 (N_3515,In_1074,In_193);
or U3516 (N_3516,In_2777,In_1567);
or U3517 (N_3517,In_2772,In_2961);
nand U3518 (N_3518,In_1760,In_2097);
nor U3519 (N_3519,In_31,In_2898);
xnor U3520 (N_3520,In_229,In_696);
nand U3521 (N_3521,In_1541,In_1018);
xnor U3522 (N_3522,In_2240,In_489);
nand U3523 (N_3523,In_781,In_1909);
nand U3524 (N_3524,In_1934,In_2951);
nand U3525 (N_3525,In_315,In_795);
and U3526 (N_3526,In_2886,In_1499);
and U3527 (N_3527,In_1790,In_1835);
xnor U3528 (N_3528,In_1517,In_620);
nor U3529 (N_3529,In_347,In_2355);
nand U3530 (N_3530,In_1666,In_1921);
and U3531 (N_3531,In_2430,In_1596);
xor U3532 (N_3532,In_2849,In_1174);
xor U3533 (N_3533,In_2320,In_2395);
or U3534 (N_3534,In_659,In_1196);
or U3535 (N_3535,In_445,In_2780);
nor U3536 (N_3536,In_1076,In_2829);
xor U3537 (N_3537,In_2241,In_393);
or U3538 (N_3538,In_354,In_2529);
or U3539 (N_3539,In_2461,In_673);
nor U3540 (N_3540,In_2504,In_1288);
and U3541 (N_3541,In_950,In_2192);
nor U3542 (N_3542,In_2242,In_2175);
nand U3543 (N_3543,In_758,In_1756);
xor U3544 (N_3544,In_2281,In_189);
xnor U3545 (N_3545,In_2592,In_1071);
nand U3546 (N_3546,In_1972,In_2560);
xor U3547 (N_3547,In_1537,In_1804);
and U3548 (N_3548,In_911,In_2608);
or U3549 (N_3549,In_506,In_321);
or U3550 (N_3550,In_333,In_1644);
or U3551 (N_3551,In_2992,In_729);
and U3552 (N_3552,In_1335,In_420);
nand U3553 (N_3553,In_94,In_574);
nor U3554 (N_3554,In_1878,In_1870);
and U3555 (N_3555,In_2513,In_2524);
nor U3556 (N_3556,In_1235,In_2526);
nand U3557 (N_3557,In_1873,In_529);
nand U3558 (N_3558,In_2075,In_2193);
nand U3559 (N_3559,In_723,In_1090);
nor U3560 (N_3560,In_1012,In_689);
and U3561 (N_3561,In_908,In_2808);
nor U3562 (N_3562,In_2021,In_2199);
and U3563 (N_3563,In_2858,In_128);
and U3564 (N_3564,In_1285,In_42);
nand U3565 (N_3565,In_1334,In_1131);
nand U3566 (N_3566,In_2218,In_309);
or U3567 (N_3567,In_1184,In_2681);
and U3568 (N_3568,In_606,In_1940);
or U3569 (N_3569,In_581,In_1267);
or U3570 (N_3570,In_1578,In_2697);
and U3571 (N_3571,In_1485,In_1507);
nor U3572 (N_3572,In_501,In_519);
or U3573 (N_3573,In_802,In_1105);
nand U3574 (N_3574,In_371,In_1574);
nand U3575 (N_3575,In_2276,In_2492);
and U3576 (N_3576,In_1849,In_2970);
xnor U3577 (N_3577,In_844,In_568);
xnor U3578 (N_3578,In_20,In_137);
or U3579 (N_3579,In_107,In_48);
xor U3580 (N_3580,In_2024,In_2155);
nand U3581 (N_3581,In_495,In_1746);
xnor U3582 (N_3582,In_463,In_2584);
or U3583 (N_3583,In_1425,In_1808);
xnor U3584 (N_3584,In_1687,In_2438);
nor U3585 (N_3585,In_2908,In_1235);
or U3586 (N_3586,In_1710,In_2956);
nand U3587 (N_3587,In_1938,In_2691);
nand U3588 (N_3588,In_2078,In_569);
nor U3589 (N_3589,In_2913,In_1163);
nand U3590 (N_3590,In_2899,In_1551);
nand U3591 (N_3591,In_601,In_507);
xnor U3592 (N_3592,In_1371,In_2892);
nor U3593 (N_3593,In_706,In_1108);
nor U3594 (N_3594,In_1988,In_2485);
nor U3595 (N_3595,In_1375,In_2531);
and U3596 (N_3596,In_1563,In_2490);
and U3597 (N_3597,In_2201,In_72);
xnor U3598 (N_3598,In_2450,In_723);
and U3599 (N_3599,In_1990,In_821);
and U3600 (N_3600,In_2913,In_2838);
nor U3601 (N_3601,In_1877,In_966);
nor U3602 (N_3602,In_2212,In_1408);
and U3603 (N_3603,In_2449,In_1418);
nor U3604 (N_3604,In_1530,In_2464);
nor U3605 (N_3605,In_848,In_1974);
nor U3606 (N_3606,In_1126,In_1664);
or U3607 (N_3607,In_83,In_1708);
xor U3608 (N_3608,In_1121,In_2822);
and U3609 (N_3609,In_2239,In_267);
nor U3610 (N_3610,In_2873,In_1083);
or U3611 (N_3611,In_320,In_1561);
nor U3612 (N_3612,In_1305,In_882);
or U3613 (N_3613,In_1382,In_1586);
xnor U3614 (N_3614,In_2418,In_2004);
xor U3615 (N_3615,In_1659,In_1952);
and U3616 (N_3616,In_606,In_884);
nor U3617 (N_3617,In_736,In_696);
xor U3618 (N_3618,In_119,In_123);
nor U3619 (N_3619,In_1070,In_25);
or U3620 (N_3620,In_1203,In_418);
nand U3621 (N_3621,In_2194,In_1303);
nand U3622 (N_3622,In_2278,In_534);
xnor U3623 (N_3623,In_2301,In_132);
xor U3624 (N_3624,In_73,In_1170);
or U3625 (N_3625,In_2243,In_2292);
nand U3626 (N_3626,In_1670,In_1174);
nand U3627 (N_3627,In_147,In_2651);
and U3628 (N_3628,In_1186,In_762);
xor U3629 (N_3629,In_999,In_2809);
nor U3630 (N_3630,In_242,In_2235);
and U3631 (N_3631,In_478,In_1613);
xor U3632 (N_3632,In_604,In_2144);
nand U3633 (N_3633,In_2768,In_1950);
nand U3634 (N_3634,In_86,In_2970);
nand U3635 (N_3635,In_991,In_1822);
or U3636 (N_3636,In_723,In_2967);
nand U3637 (N_3637,In_685,In_401);
nor U3638 (N_3638,In_1148,In_203);
xor U3639 (N_3639,In_2691,In_1059);
and U3640 (N_3640,In_2679,In_327);
xor U3641 (N_3641,In_582,In_583);
nand U3642 (N_3642,In_963,In_258);
nor U3643 (N_3643,In_375,In_87);
nand U3644 (N_3644,In_1973,In_1074);
nand U3645 (N_3645,In_2977,In_2809);
or U3646 (N_3646,In_1047,In_1645);
and U3647 (N_3647,In_465,In_1562);
nand U3648 (N_3648,In_2257,In_2174);
and U3649 (N_3649,In_1812,In_1646);
nor U3650 (N_3650,In_2187,In_2768);
xnor U3651 (N_3651,In_470,In_2647);
xor U3652 (N_3652,In_2272,In_2140);
or U3653 (N_3653,In_2436,In_767);
or U3654 (N_3654,In_2996,In_2349);
nand U3655 (N_3655,In_1226,In_365);
or U3656 (N_3656,In_2019,In_13);
or U3657 (N_3657,In_1340,In_611);
xor U3658 (N_3658,In_1467,In_176);
and U3659 (N_3659,In_1371,In_483);
and U3660 (N_3660,In_68,In_2766);
xor U3661 (N_3661,In_1477,In_1227);
nand U3662 (N_3662,In_420,In_1896);
xnor U3663 (N_3663,In_2062,In_1041);
nor U3664 (N_3664,In_1314,In_746);
nor U3665 (N_3665,In_1138,In_279);
xnor U3666 (N_3666,In_2221,In_1051);
nand U3667 (N_3667,In_424,In_2555);
xnor U3668 (N_3668,In_290,In_1270);
nand U3669 (N_3669,In_208,In_2285);
xnor U3670 (N_3670,In_185,In_609);
nor U3671 (N_3671,In_2817,In_1616);
or U3672 (N_3672,In_561,In_2772);
xor U3673 (N_3673,In_2032,In_39);
nor U3674 (N_3674,In_999,In_1487);
nor U3675 (N_3675,In_617,In_1520);
or U3676 (N_3676,In_1307,In_1789);
or U3677 (N_3677,In_572,In_1733);
and U3678 (N_3678,In_1597,In_119);
xnor U3679 (N_3679,In_2577,In_887);
nand U3680 (N_3680,In_2282,In_2038);
xor U3681 (N_3681,In_2558,In_2809);
xor U3682 (N_3682,In_2103,In_2336);
and U3683 (N_3683,In_811,In_1000);
nor U3684 (N_3684,In_964,In_1296);
xnor U3685 (N_3685,In_510,In_453);
or U3686 (N_3686,In_566,In_402);
xnor U3687 (N_3687,In_1961,In_1139);
nor U3688 (N_3688,In_89,In_463);
nor U3689 (N_3689,In_1785,In_1495);
nand U3690 (N_3690,In_2849,In_1874);
nand U3691 (N_3691,In_862,In_1058);
nor U3692 (N_3692,In_709,In_1665);
and U3693 (N_3693,In_163,In_474);
xnor U3694 (N_3694,In_787,In_961);
nor U3695 (N_3695,In_988,In_2598);
nand U3696 (N_3696,In_1512,In_2079);
nand U3697 (N_3697,In_847,In_1539);
nand U3698 (N_3698,In_2083,In_2913);
nor U3699 (N_3699,In_2167,In_584);
or U3700 (N_3700,In_740,In_2667);
and U3701 (N_3701,In_220,In_62);
xnor U3702 (N_3702,In_2385,In_872);
or U3703 (N_3703,In_2012,In_1331);
and U3704 (N_3704,In_2324,In_2800);
or U3705 (N_3705,In_2372,In_1692);
and U3706 (N_3706,In_980,In_2381);
and U3707 (N_3707,In_2844,In_1180);
nand U3708 (N_3708,In_2475,In_1205);
nand U3709 (N_3709,In_1930,In_1503);
nor U3710 (N_3710,In_2183,In_1730);
nor U3711 (N_3711,In_368,In_906);
xnor U3712 (N_3712,In_1293,In_448);
or U3713 (N_3713,In_2661,In_1778);
or U3714 (N_3714,In_736,In_660);
and U3715 (N_3715,In_2713,In_2649);
nor U3716 (N_3716,In_2446,In_187);
and U3717 (N_3717,In_1938,In_2047);
or U3718 (N_3718,In_2313,In_899);
nand U3719 (N_3719,In_668,In_1419);
nand U3720 (N_3720,In_1860,In_2824);
xnor U3721 (N_3721,In_1928,In_325);
or U3722 (N_3722,In_1902,In_831);
nor U3723 (N_3723,In_1930,In_2043);
or U3724 (N_3724,In_2032,In_1870);
nand U3725 (N_3725,In_2142,In_1991);
and U3726 (N_3726,In_463,In_1354);
nand U3727 (N_3727,In_1960,In_850);
and U3728 (N_3728,In_2352,In_2763);
nor U3729 (N_3729,In_2353,In_2076);
nor U3730 (N_3730,In_2885,In_2300);
nand U3731 (N_3731,In_2343,In_370);
and U3732 (N_3732,In_2820,In_63);
nor U3733 (N_3733,In_1502,In_2465);
and U3734 (N_3734,In_1935,In_1879);
xnor U3735 (N_3735,In_1110,In_1564);
or U3736 (N_3736,In_1424,In_2797);
nand U3737 (N_3737,In_2071,In_1206);
xnor U3738 (N_3738,In_2636,In_2092);
xnor U3739 (N_3739,In_469,In_1302);
nor U3740 (N_3740,In_2344,In_678);
and U3741 (N_3741,In_841,In_2428);
nand U3742 (N_3742,In_2874,In_1765);
nand U3743 (N_3743,In_2053,In_2951);
nor U3744 (N_3744,In_2943,In_234);
nor U3745 (N_3745,In_1543,In_139);
nand U3746 (N_3746,In_2926,In_1809);
nor U3747 (N_3747,In_429,In_2743);
nor U3748 (N_3748,In_1603,In_2281);
nand U3749 (N_3749,In_344,In_2571);
and U3750 (N_3750,In_438,In_1560);
and U3751 (N_3751,In_539,In_284);
or U3752 (N_3752,In_988,In_233);
nand U3753 (N_3753,In_2546,In_1115);
or U3754 (N_3754,In_853,In_2720);
nand U3755 (N_3755,In_1149,In_795);
nor U3756 (N_3756,In_2020,In_2515);
or U3757 (N_3757,In_293,In_2138);
nand U3758 (N_3758,In_277,In_2715);
and U3759 (N_3759,In_847,In_2982);
nand U3760 (N_3760,In_2871,In_108);
nand U3761 (N_3761,In_2030,In_2005);
xor U3762 (N_3762,In_2695,In_1237);
xor U3763 (N_3763,In_1141,In_732);
or U3764 (N_3764,In_1502,In_2359);
or U3765 (N_3765,In_1969,In_859);
xnor U3766 (N_3766,In_788,In_865);
and U3767 (N_3767,In_2390,In_453);
and U3768 (N_3768,In_2933,In_1188);
and U3769 (N_3769,In_1817,In_2698);
or U3770 (N_3770,In_2793,In_2116);
nand U3771 (N_3771,In_1857,In_1934);
nor U3772 (N_3772,In_2840,In_2049);
xnor U3773 (N_3773,In_2997,In_2201);
or U3774 (N_3774,In_2056,In_615);
nor U3775 (N_3775,In_2590,In_1416);
and U3776 (N_3776,In_696,In_163);
or U3777 (N_3777,In_1480,In_377);
or U3778 (N_3778,In_2876,In_2077);
or U3779 (N_3779,In_2489,In_2790);
xor U3780 (N_3780,In_845,In_191);
nand U3781 (N_3781,In_18,In_2115);
and U3782 (N_3782,In_2716,In_2805);
and U3783 (N_3783,In_726,In_1375);
nor U3784 (N_3784,In_575,In_2674);
nand U3785 (N_3785,In_2850,In_704);
and U3786 (N_3786,In_2724,In_2397);
xnor U3787 (N_3787,In_1431,In_1112);
and U3788 (N_3788,In_2421,In_2104);
nand U3789 (N_3789,In_348,In_1883);
nand U3790 (N_3790,In_1797,In_989);
or U3791 (N_3791,In_1886,In_2790);
nor U3792 (N_3792,In_2601,In_1703);
xnor U3793 (N_3793,In_2153,In_818);
nand U3794 (N_3794,In_898,In_182);
nor U3795 (N_3795,In_469,In_1575);
nor U3796 (N_3796,In_1607,In_855);
or U3797 (N_3797,In_1335,In_2713);
and U3798 (N_3798,In_43,In_154);
and U3799 (N_3799,In_961,In_1651);
nand U3800 (N_3800,In_833,In_2045);
xor U3801 (N_3801,In_2064,In_354);
nand U3802 (N_3802,In_928,In_605);
or U3803 (N_3803,In_2734,In_1791);
nor U3804 (N_3804,In_2834,In_1762);
nand U3805 (N_3805,In_801,In_634);
xor U3806 (N_3806,In_2847,In_2324);
and U3807 (N_3807,In_1998,In_2666);
nor U3808 (N_3808,In_2419,In_885);
xnor U3809 (N_3809,In_1788,In_1275);
xnor U3810 (N_3810,In_2876,In_364);
nor U3811 (N_3811,In_2951,In_624);
nand U3812 (N_3812,In_1166,In_2039);
nand U3813 (N_3813,In_2275,In_1544);
or U3814 (N_3814,In_2592,In_2116);
nor U3815 (N_3815,In_546,In_2319);
xor U3816 (N_3816,In_1149,In_1324);
or U3817 (N_3817,In_1388,In_2448);
nand U3818 (N_3818,In_532,In_2359);
xnor U3819 (N_3819,In_901,In_2747);
xor U3820 (N_3820,In_2876,In_2354);
nand U3821 (N_3821,In_1143,In_1213);
xnor U3822 (N_3822,In_2375,In_2132);
xor U3823 (N_3823,In_1739,In_2902);
nand U3824 (N_3824,In_2145,In_727);
xor U3825 (N_3825,In_414,In_2898);
xnor U3826 (N_3826,In_299,In_934);
xnor U3827 (N_3827,In_134,In_2204);
nand U3828 (N_3828,In_1418,In_493);
nand U3829 (N_3829,In_1470,In_2923);
nor U3830 (N_3830,In_2094,In_357);
xor U3831 (N_3831,In_1590,In_2051);
or U3832 (N_3832,In_1620,In_2848);
and U3833 (N_3833,In_908,In_2381);
nand U3834 (N_3834,In_1817,In_1278);
nor U3835 (N_3835,In_1987,In_2114);
nand U3836 (N_3836,In_1801,In_904);
or U3837 (N_3837,In_992,In_2006);
xor U3838 (N_3838,In_246,In_1036);
xnor U3839 (N_3839,In_2151,In_1447);
xnor U3840 (N_3840,In_2002,In_1951);
and U3841 (N_3841,In_875,In_1234);
or U3842 (N_3842,In_1395,In_2888);
and U3843 (N_3843,In_2186,In_972);
xnor U3844 (N_3844,In_386,In_1123);
or U3845 (N_3845,In_2071,In_724);
nand U3846 (N_3846,In_2358,In_667);
and U3847 (N_3847,In_2970,In_2955);
xor U3848 (N_3848,In_2712,In_2054);
or U3849 (N_3849,In_2415,In_688);
xor U3850 (N_3850,In_1301,In_819);
nand U3851 (N_3851,In_1400,In_2569);
xnor U3852 (N_3852,In_1470,In_2980);
and U3853 (N_3853,In_1624,In_153);
nand U3854 (N_3854,In_295,In_537);
nor U3855 (N_3855,In_1943,In_1233);
xnor U3856 (N_3856,In_39,In_1884);
or U3857 (N_3857,In_2322,In_441);
nand U3858 (N_3858,In_1025,In_14);
nor U3859 (N_3859,In_909,In_58);
xnor U3860 (N_3860,In_891,In_446);
xor U3861 (N_3861,In_1010,In_139);
xor U3862 (N_3862,In_1853,In_2718);
and U3863 (N_3863,In_1590,In_224);
xnor U3864 (N_3864,In_996,In_749);
or U3865 (N_3865,In_2881,In_2857);
nor U3866 (N_3866,In_1860,In_2730);
and U3867 (N_3867,In_2637,In_772);
xnor U3868 (N_3868,In_1250,In_350);
nand U3869 (N_3869,In_742,In_2219);
nor U3870 (N_3870,In_1635,In_547);
xnor U3871 (N_3871,In_2795,In_721);
nor U3872 (N_3872,In_859,In_2017);
nand U3873 (N_3873,In_2461,In_2215);
nor U3874 (N_3874,In_822,In_1522);
nor U3875 (N_3875,In_2181,In_1234);
and U3876 (N_3876,In_1393,In_2290);
or U3877 (N_3877,In_2961,In_1610);
or U3878 (N_3878,In_1485,In_1047);
or U3879 (N_3879,In_723,In_2702);
or U3880 (N_3880,In_320,In_572);
xor U3881 (N_3881,In_345,In_482);
or U3882 (N_3882,In_1608,In_1307);
or U3883 (N_3883,In_2332,In_2990);
and U3884 (N_3884,In_2087,In_2227);
and U3885 (N_3885,In_2140,In_1057);
xnor U3886 (N_3886,In_2128,In_2067);
or U3887 (N_3887,In_2300,In_2801);
and U3888 (N_3888,In_450,In_1727);
or U3889 (N_3889,In_1928,In_1437);
or U3890 (N_3890,In_2549,In_361);
nand U3891 (N_3891,In_2892,In_251);
nand U3892 (N_3892,In_219,In_442);
or U3893 (N_3893,In_351,In_1337);
or U3894 (N_3894,In_2174,In_1402);
or U3895 (N_3895,In_2478,In_425);
nor U3896 (N_3896,In_468,In_1260);
or U3897 (N_3897,In_1438,In_1927);
xor U3898 (N_3898,In_2821,In_2034);
nand U3899 (N_3899,In_418,In_950);
nor U3900 (N_3900,In_2285,In_2812);
nor U3901 (N_3901,In_2652,In_2890);
and U3902 (N_3902,In_1280,In_769);
xor U3903 (N_3903,In_1052,In_2060);
nor U3904 (N_3904,In_14,In_2827);
xnor U3905 (N_3905,In_22,In_2314);
nor U3906 (N_3906,In_825,In_1776);
nor U3907 (N_3907,In_2148,In_2797);
or U3908 (N_3908,In_2060,In_768);
nor U3909 (N_3909,In_1855,In_243);
nand U3910 (N_3910,In_1258,In_1497);
xor U3911 (N_3911,In_2967,In_2391);
nor U3912 (N_3912,In_157,In_1115);
nor U3913 (N_3913,In_1647,In_826);
or U3914 (N_3914,In_1699,In_2143);
nor U3915 (N_3915,In_2958,In_1656);
nand U3916 (N_3916,In_2821,In_2115);
or U3917 (N_3917,In_453,In_1313);
xor U3918 (N_3918,In_2685,In_295);
nand U3919 (N_3919,In_2558,In_1776);
nand U3920 (N_3920,In_2992,In_875);
nand U3921 (N_3921,In_1347,In_957);
nand U3922 (N_3922,In_2209,In_222);
nor U3923 (N_3923,In_2184,In_2514);
xnor U3924 (N_3924,In_857,In_1309);
and U3925 (N_3925,In_1977,In_1786);
and U3926 (N_3926,In_2391,In_290);
nor U3927 (N_3927,In_27,In_2460);
nor U3928 (N_3928,In_2255,In_2368);
nand U3929 (N_3929,In_744,In_2880);
nand U3930 (N_3930,In_1129,In_270);
and U3931 (N_3931,In_182,In_1831);
or U3932 (N_3932,In_1418,In_2350);
and U3933 (N_3933,In_28,In_2908);
nor U3934 (N_3934,In_2604,In_2522);
xnor U3935 (N_3935,In_1327,In_2171);
xnor U3936 (N_3936,In_2818,In_1738);
xor U3937 (N_3937,In_1732,In_795);
and U3938 (N_3938,In_2950,In_83);
and U3939 (N_3939,In_2565,In_359);
nand U3940 (N_3940,In_2194,In_432);
and U3941 (N_3941,In_268,In_1614);
xnor U3942 (N_3942,In_2704,In_2042);
nor U3943 (N_3943,In_621,In_1706);
or U3944 (N_3944,In_120,In_2038);
or U3945 (N_3945,In_1480,In_1778);
nor U3946 (N_3946,In_22,In_2151);
nand U3947 (N_3947,In_655,In_391);
nand U3948 (N_3948,In_1325,In_1862);
xnor U3949 (N_3949,In_1274,In_2244);
xnor U3950 (N_3950,In_1216,In_702);
and U3951 (N_3951,In_1559,In_2035);
and U3952 (N_3952,In_2656,In_0);
and U3953 (N_3953,In_1381,In_1751);
nor U3954 (N_3954,In_1442,In_1040);
nor U3955 (N_3955,In_1699,In_1256);
and U3956 (N_3956,In_1888,In_758);
or U3957 (N_3957,In_159,In_166);
nor U3958 (N_3958,In_685,In_449);
and U3959 (N_3959,In_2915,In_2066);
or U3960 (N_3960,In_408,In_69);
nand U3961 (N_3961,In_1948,In_1654);
and U3962 (N_3962,In_513,In_2873);
xnor U3963 (N_3963,In_2100,In_1749);
xor U3964 (N_3964,In_404,In_1343);
nor U3965 (N_3965,In_1427,In_821);
nor U3966 (N_3966,In_1367,In_814);
xnor U3967 (N_3967,In_496,In_2290);
xor U3968 (N_3968,In_1823,In_1469);
nor U3969 (N_3969,In_1255,In_1485);
nor U3970 (N_3970,In_2689,In_1196);
nand U3971 (N_3971,In_548,In_897);
nand U3972 (N_3972,In_350,In_2048);
nor U3973 (N_3973,In_731,In_1613);
nand U3974 (N_3974,In_138,In_2948);
or U3975 (N_3975,In_2400,In_573);
nor U3976 (N_3976,In_1667,In_858);
nand U3977 (N_3977,In_1434,In_1184);
and U3978 (N_3978,In_1804,In_1192);
xor U3979 (N_3979,In_2568,In_2176);
xnor U3980 (N_3980,In_3,In_16);
xor U3981 (N_3981,In_2452,In_1223);
nand U3982 (N_3982,In_2473,In_1837);
nor U3983 (N_3983,In_879,In_221);
nand U3984 (N_3984,In_154,In_1260);
nand U3985 (N_3985,In_427,In_1583);
xor U3986 (N_3986,In_114,In_554);
or U3987 (N_3987,In_1386,In_396);
nor U3988 (N_3988,In_1432,In_557);
nor U3989 (N_3989,In_383,In_498);
xnor U3990 (N_3990,In_1620,In_1604);
xnor U3991 (N_3991,In_2845,In_2051);
nand U3992 (N_3992,In_1953,In_667);
nand U3993 (N_3993,In_2241,In_686);
or U3994 (N_3994,In_1459,In_1758);
or U3995 (N_3995,In_1945,In_2631);
nor U3996 (N_3996,In_2173,In_2418);
and U3997 (N_3997,In_1265,In_2603);
or U3998 (N_3998,In_1597,In_392);
or U3999 (N_3999,In_1171,In_1757);
nor U4000 (N_4000,In_379,In_2118);
or U4001 (N_4001,In_988,In_1867);
xor U4002 (N_4002,In_1761,In_1208);
or U4003 (N_4003,In_940,In_2938);
nand U4004 (N_4004,In_296,In_353);
nand U4005 (N_4005,In_2859,In_2287);
nor U4006 (N_4006,In_678,In_2242);
and U4007 (N_4007,In_521,In_1553);
xnor U4008 (N_4008,In_2632,In_1806);
nand U4009 (N_4009,In_639,In_2175);
and U4010 (N_4010,In_631,In_2785);
xor U4011 (N_4011,In_610,In_673);
and U4012 (N_4012,In_197,In_2712);
nor U4013 (N_4013,In_2049,In_1791);
xor U4014 (N_4014,In_549,In_1706);
or U4015 (N_4015,In_1584,In_2978);
or U4016 (N_4016,In_1768,In_1429);
or U4017 (N_4017,In_1510,In_2007);
or U4018 (N_4018,In_1174,In_2396);
xnor U4019 (N_4019,In_2569,In_652);
nand U4020 (N_4020,In_688,In_1344);
xor U4021 (N_4021,In_519,In_2533);
nand U4022 (N_4022,In_1314,In_1367);
xor U4023 (N_4023,In_448,In_2474);
nor U4024 (N_4024,In_179,In_2062);
xnor U4025 (N_4025,In_302,In_2783);
nor U4026 (N_4026,In_449,In_2052);
or U4027 (N_4027,In_2554,In_53);
xnor U4028 (N_4028,In_2849,In_1199);
xnor U4029 (N_4029,In_851,In_1646);
nor U4030 (N_4030,In_2028,In_1185);
nand U4031 (N_4031,In_1709,In_162);
nand U4032 (N_4032,In_2726,In_610);
xnor U4033 (N_4033,In_572,In_855);
nand U4034 (N_4034,In_135,In_288);
nor U4035 (N_4035,In_660,In_2401);
and U4036 (N_4036,In_2021,In_1657);
xnor U4037 (N_4037,In_2906,In_1434);
nor U4038 (N_4038,In_1514,In_783);
nor U4039 (N_4039,In_187,In_2709);
or U4040 (N_4040,In_17,In_1881);
nor U4041 (N_4041,In_1895,In_728);
or U4042 (N_4042,In_257,In_425);
xnor U4043 (N_4043,In_1648,In_707);
and U4044 (N_4044,In_994,In_2380);
nand U4045 (N_4045,In_2079,In_657);
and U4046 (N_4046,In_1757,In_586);
or U4047 (N_4047,In_2142,In_2686);
and U4048 (N_4048,In_17,In_1703);
nor U4049 (N_4049,In_2800,In_224);
nor U4050 (N_4050,In_616,In_238);
nor U4051 (N_4051,In_1465,In_418);
and U4052 (N_4052,In_808,In_2689);
xnor U4053 (N_4053,In_1914,In_2820);
or U4054 (N_4054,In_1946,In_2053);
and U4055 (N_4055,In_1109,In_980);
or U4056 (N_4056,In_1702,In_1747);
or U4057 (N_4057,In_1643,In_909);
nand U4058 (N_4058,In_2161,In_1590);
or U4059 (N_4059,In_818,In_2465);
nand U4060 (N_4060,In_951,In_2019);
nor U4061 (N_4061,In_2800,In_434);
xnor U4062 (N_4062,In_1885,In_1732);
nand U4063 (N_4063,In_223,In_961);
xor U4064 (N_4064,In_1561,In_2732);
nor U4065 (N_4065,In_1238,In_1964);
xnor U4066 (N_4066,In_2791,In_2157);
and U4067 (N_4067,In_1717,In_1016);
and U4068 (N_4068,In_1447,In_1808);
nor U4069 (N_4069,In_1456,In_934);
xnor U4070 (N_4070,In_917,In_518);
nor U4071 (N_4071,In_1898,In_144);
xor U4072 (N_4072,In_890,In_673);
nor U4073 (N_4073,In_2176,In_2573);
nor U4074 (N_4074,In_1692,In_198);
nand U4075 (N_4075,In_2579,In_317);
nand U4076 (N_4076,In_1683,In_1496);
or U4077 (N_4077,In_382,In_2854);
xor U4078 (N_4078,In_412,In_1918);
nor U4079 (N_4079,In_1557,In_550);
xnor U4080 (N_4080,In_1980,In_2759);
nand U4081 (N_4081,In_1298,In_1640);
nand U4082 (N_4082,In_1204,In_400);
nand U4083 (N_4083,In_13,In_815);
nor U4084 (N_4084,In_2503,In_829);
nor U4085 (N_4085,In_88,In_1986);
nand U4086 (N_4086,In_1293,In_1046);
nand U4087 (N_4087,In_2471,In_2015);
or U4088 (N_4088,In_751,In_28);
and U4089 (N_4089,In_524,In_603);
and U4090 (N_4090,In_2265,In_2372);
xor U4091 (N_4091,In_2992,In_2371);
nor U4092 (N_4092,In_7,In_234);
and U4093 (N_4093,In_1431,In_2554);
or U4094 (N_4094,In_2982,In_1098);
or U4095 (N_4095,In_159,In_120);
and U4096 (N_4096,In_956,In_1446);
or U4097 (N_4097,In_769,In_1721);
or U4098 (N_4098,In_2385,In_2521);
or U4099 (N_4099,In_1486,In_2575);
and U4100 (N_4100,In_1375,In_498);
nand U4101 (N_4101,In_2378,In_2415);
xnor U4102 (N_4102,In_1698,In_960);
xor U4103 (N_4103,In_2472,In_1110);
nor U4104 (N_4104,In_530,In_2402);
nand U4105 (N_4105,In_1595,In_2785);
xnor U4106 (N_4106,In_501,In_1096);
nor U4107 (N_4107,In_1504,In_2077);
xnor U4108 (N_4108,In_1000,In_1801);
xnor U4109 (N_4109,In_26,In_1140);
or U4110 (N_4110,In_1934,In_2906);
nand U4111 (N_4111,In_1543,In_2677);
and U4112 (N_4112,In_719,In_232);
and U4113 (N_4113,In_120,In_189);
nor U4114 (N_4114,In_724,In_1879);
nor U4115 (N_4115,In_476,In_926);
and U4116 (N_4116,In_2487,In_2394);
nand U4117 (N_4117,In_2689,In_1536);
xor U4118 (N_4118,In_1334,In_2682);
nor U4119 (N_4119,In_84,In_2616);
nand U4120 (N_4120,In_1061,In_2116);
or U4121 (N_4121,In_143,In_1638);
xor U4122 (N_4122,In_390,In_388);
xor U4123 (N_4123,In_1350,In_1634);
xnor U4124 (N_4124,In_1262,In_451);
nor U4125 (N_4125,In_1700,In_2035);
and U4126 (N_4126,In_2211,In_1933);
nand U4127 (N_4127,In_2682,In_1242);
and U4128 (N_4128,In_1559,In_2819);
nand U4129 (N_4129,In_722,In_1001);
xnor U4130 (N_4130,In_2509,In_769);
nand U4131 (N_4131,In_802,In_681);
nor U4132 (N_4132,In_582,In_827);
xor U4133 (N_4133,In_128,In_560);
or U4134 (N_4134,In_351,In_1162);
or U4135 (N_4135,In_2728,In_1310);
xor U4136 (N_4136,In_1488,In_2625);
and U4137 (N_4137,In_2376,In_227);
xor U4138 (N_4138,In_54,In_2230);
nor U4139 (N_4139,In_2388,In_2839);
xor U4140 (N_4140,In_849,In_2788);
nor U4141 (N_4141,In_2274,In_2607);
or U4142 (N_4142,In_598,In_2197);
nor U4143 (N_4143,In_1044,In_1917);
and U4144 (N_4144,In_1065,In_247);
and U4145 (N_4145,In_1333,In_592);
xor U4146 (N_4146,In_2543,In_2210);
and U4147 (N_4147,In_646,In_1603);
and U4148 (N_4148,In_2383,In_1996);
nand U4149 (N_4149,In_485,In_1822);
xnor U4150 (N_4150,In_640,In_1850);
nand U4151 (N_4151,In_2889,In_2649);
and U4152 (N_4152,In_2577,In_112);
nand U4153 (N_4153,In_2345,In_1842);
nor U4154 (N_4154,In_2911,In_223);
and U4155 (N_4155,In_2938,In_2539);
nand U4156 (N_4156,In_244,In_165);
nand U4157 (N_4157,In_187,In_2456);
nor U4158 (N_4158,In_655,In_340);
and U4159 (N_4159,In_705,In_856);
xnor U4160 (N_4160,In_189,In_2826);
xnor U4161 (N_4161,In_1301,In_1586);
nand U4162 (N_4162,In_2876,In_1554);
nor U4163 (N_4163,In_2772,In_2102);
or U4164 (N_4164,In_2399,In_1301);
nor U4165 (N_4165,In_800,In_567);
and U4166 (N_4166,In_1058,In_1496);
nor U4167 (N_4167,In_1630,In_1651);
or U4168 (N_4168,In_158,In_1868);
or U4169 (N_4169,In_1289,In_2338);
and U4170 (N_4170,In_2144,In_974);
xnor U4171 (N_4171,In_1904,In_776);
xor U4172 (N_4172,In_1484,In_1532);
xor U4173 (N_4173,In_1211,In_2161);
or U4174 (N_4174,In_112,In_1260);
xor U4175 (N_4175,In_1787,In_2911);
nor U4176 (N_4176,In_1,In_944);
nand U4177 (N_4177,In_735,In_2218);
xnor U4178 (N_4178,In_750,In_2562);
nor U4179 (N_4179,In_581,In_2865);
and U4180 (N_4180,In_2961,In_406);
and U4181 (N_4181,In_192,In_935);
xnor U4182 (N_4182,In_1081,In_1881);
nand U4183 (N_4183,In_1585,In_2923);
and U4184 (N_4184,In_2914,In_131);
or U4185 (N_4185,In_1863,In_1418);
xnor U4186 (N_4186,In_1649,In_1672);
and U4187 (N_4187,In_1879,In_214);
and U4188 (N_4188,In_1623,In_413);
or U4189 (N_4189,In_2791,In_1855);
nor U4190 (N_4190,In_1220,In_675);
xor U4191 (N_4191,In_2272,In_1060);
nand U4192 (N_4192,In_277,In_1303);
or U4193 (N_4193,In_1412,In_1826);
xor U4194 (N_4194,In_2130,In_2599);
xor U4195 (N_4195,In_1098,In_1111);
and U4196 (N_4196,In_2659,In_470);
and U4197 (N_4197,In_257,In_1356);
xor U4198 (N_4198,In_761,In_936);
nor U4199 (N_4199,In_2867,In_629);
or U4200 (N_4200,In_1124,In_271);
or U4201 (N_4201,In_1452,In_867);
nand U4202 (N_4202,In_2732,In_980);
nand U4203 (N_4203,In_2315,In_635);
nand U4204 (N_4204,In_2610,In_665);
xnor U4205 (N_4205,In_2795,In_667);
or U4206 (N_4206,In_698,In_1065);
and U4207 (N_4207,In_1542,In_1653);
or U4208 (N_4208,In_2939,In_225);
xnor U4209 (N_4209,In_1991,In_426);
and U4210 (N_4210,In_804,In_690);
or U4211 (N_4211,In_1803,In_2098);
nor U4212 (N_4212,In_1639,In_1006);
nand U4213 (N_4213,In_817,In_340);
nand U4214 (N_4214,In_2983,In_612);
and U4215 (N_4215,In_814,In_2645);
and U4216 (N_4216,In_497,In_1698);
nor U4217 (N_4217,In_2379,In_1873);
xnor U4218 (N_4218,In_1493,In_1609);
and U4219 (N_4219,In_363,In_2879);
or U4220 (N_4220,In_1805,In_454);
xnor U4221 (N_4221,In_2793,In_882);
nor U4222 (N_4222,In_2705,In_2805);
or U4223 (N_4223,In_2253,In_2794);
xor U4224 (N_4224,In_1498,In_102);
and U4225 (N_4225,In_2824,In_2389);
nand U4226 (N_4226,In_69,In_2306);
xor U4227 (N_4227,In_378,In_380);
xnor U4228 (N_4228,In_1247,In_2082);
and U4229 (N_4229,In_2250,In_1393);
xnor U4230 (N_4230,In_994,In_913);
nand U4231 (N_4231,In_582,In_2426);
nor U4232 (N_4232,In_666,In_2643);
nand U4233 (N_4233,In_2188,In_357);
xor U4234 (N_4234,In_1679,In_1784);
and U4235 (N_4235,In_144,In_2006);
or U4236 (N_4236,In_2836,In_2425);
xnor U4237 (N_4237,In_2110,In_2482);
nand U4238 (N_4238,In_1346,In_2431);
or U4239 (N_4239,In_1091,In_1352);
or U4240 (N_4240,In_1682,In_1301);
nor U4241 (N_4241,In_1680,In_2654);
or U4242 (N_4242,In_609,In_2491);
xor U4243 (N_4243,In_1017,In_2468);
nand U4244 (N_4244,In_1733,In_1541);
or U4245 (N_4245,In_19,In_1878);
xnor U4246 (N_4246,In_1246,In_880);
nor U4247 (N_4247,In_1625,In_2635);
and U4248 (N_4248,In_847,In_1242);
xnor U4249 (N_4249,In_2817,In_2702);
or U4250 (N_4250,In_651,In_2363);
xor U4251 (N_4251,In_2043,In_2427);
xor U4252 (N_4252,In_2066,In_1124);
and U4253 (N_4253,In_2797,In_2011);
and U4254 (N_4254,In_79,In_2813);
nand U4255 (N_4255,In_1106,In_2766);
and U4256 (N_4256,In_276,In_1864);
nand U4257 (N_4257,In_916,In_2522);
or U4258 (N_4258,In_1773,In_27);
xnor U4259 (N_4259,In_2366,In_1191);
nand U4260 (N_4260,In_2307,In_1029);
or U4261 (N_4261,In_970,In_2391);
nand U4262 (N_4262,In_843,In_1250);
and U4263 (N_4263,In_2831,In_1300);
nor U4264 (N_4264,In_1132,In_2956);
xor U4265 (N_4265,In_1107,In_775);
nand U4266 (N_4266,In_2961,In_972);
or U4267 (N_4267,In_1360,In_1631);
and U4268 (N_4268,In_2432,In_2218);
xnor U4269 (N_4269,In_890,In_1474);
and U4270 (N_4270,In_1761,In_1928);
nand U4271 (N_4271,In_2543,In_2624);
or U4272 (N_4272,In_29,In_1832);
and U4273 (N_4273,In_2965,In_1800);
nor U4274 (N_4274,In_1761,In_242);
nand U4275 (N_4275,In_989,In_2920);
xor U4276 (N_4276,In_2798,In_1870);
xor U4277 (N_4277,In_2496,In_2235);
or U4278 (N_4278,In_692,In_2455);
nor U4279 (N_4279,In_2153,In_108);
nor U4280 (N_4280,In_1305,In_2130);
or U4281 (N_4281,In_1883,In_2856);
nor U4282 (N_4282,In_1453,In_1782);
or U4283 (N_4283,In_1854,In_1598);
nor U4284 (N_4284,In_1130,In_855);
nand U4285 (N_4285,In_196,In_1275);
nand U4286 (N_4286,In_319,In_850);
xnor U4287 (N_4287,In_2058,In_902);
nand U4288 (N_4288,In_1912,In_2713);
nand U4289 (N_4289,In_2880,In_2463);
or U4290 (N_4290,In_1049,In_834);
xor U4291 (N_4291,In_730,In_1351);
nor U4292 (N_4292,In_397,In_2994);
nand U4293 (N_4293,In_2305,In_2731);
or U4294 (N_4294,In_1551,In_2130);
xnor U4295 (N_4295,In_756,In_1456);
nor U4296 (N_4296,In_468,In_832);
nor U4297 (N_4297,In_1430,In_412);
nand U4298 (N_4298,In_1057,In_2325);
nand U4299 (N_4299,In_482,In_1042);
xor U4300 (N_4300,In_345,In_2673);
xor U4301 (N_4301,In_613,In_114);
and U4302 (N_4302,In_729,In_1451);
nor U4303 (N_4303,In_1760,In_2425);
nand U4304 (N_4304,In_2747,In_42);
nand U4305 (N_4305,In_2319,In_2405);
or U4306 (N_4306,In_726,In_311);
nor U4307 (N_4307,In_1169,In_2301);
and U4308 (N_4308,In_1187,In_2040);
and U4309 (N_4309,In_482,In_1607);
xnor U4310 (N_4310,In_557,In_1531);
nand U4311 (N_4311,In_2471,In_2016);
xnor U4312 (N_4312,In_2560,In_2832);
or U4313 (N_4313,In_342,In_584);
nand U4314 (N_4314,In_114,In_2650);
and U4315 (N_4315,In_2316,In_2702);
xor U4316 (N_4316,In_1901,In_498);
nand U4317 (N_4317,In_2438,In_1676);
and U4318 (N_4318,In_205,In_137);
or U4319 (N_4319,In_869,In_1447);
nor U4320 (N_4320,In_1517,In_798);
xor U4321 (N_4321,In_882,In_2731);
nand U4322 (N_4322,In_2465,In_1394);
or U4323 (N_4323,In_2330,In_1245);
and U4324 (N_4324,In_1963,In_2426);
nor U4325 (N_4325,In_241,In_848);
nor U4326 (N_4326,In_1139,In_1801);
and U4327 (N_4327,In_156,In_1625);
or U4328 (N_4328,In_2697,In_2830);
nand U4329 (N_4329,In_2757,In_1155);
nor U4330 (N_4330,In_2206,In_449);
and U4331 (N_4331,In_166,In_2883);
and U4332 (N_4332,In_802,In_1137);
nor U4333 (N_4333,In_2396,In_2448);
xnor U4334 (N_4334,In_1351,In_2127);
xnor U4335 (N_4335,In_494,In_1604);
nor U4336 (N_4336,In_2951,In_1085);
or U4337 (N_4337,In_2716,In_2437);
or U4338 (N_4338,In_766,In_945);
nor U4339 (N_4339,In_814,In_1910);
and U4340 (N_4340,In_2650,In_1254);
xor U4341 (N_4341,In_2268,In_313);
nand U4342 (N_4342,In_2843,In_2941);
nand U4343 (N_4343,In_71,In_1643);
nor U4344 (N_4344,In_347,In_2814);
nand U4345 (N_4345,In_2211,In_1676);
or U4346 (N_4346,In_2003,In_1938);
nor U4347 (N_4347,In_1806,In_1477);
nor U4348 (N_4348,In_1418,In_157);
or U4349 (N_4349,In_2543,In_1357);
xor U4350 (N_4350,In_1295,In_1108);
and U4351 (N_4351,In_2057,In_2369);
and U4352 (N_4352,In_1841,In_2676);
and U4353 (N_4353,In_1713,In_1708);
xor U4354 (N_4354,In_1101,In_2805);
xnor U4355 (N_4355,In_1206,In_1808);
nor U4356 (N_4356,In_2914,In_2502);
nand U4357 (N_4357,In_745,In_859);
nor U4358 (N_4358,In_282,In_329);
nor U4359 (N_4359,In_2342,In_1360);
and U4360 (N_4360,In_1319,In_75);
or U4361 (N_4361,In_528,In_1386);
nand U4362 (N_4362,In_1662,In_728);
nand U4363 (N_4363,In_2390,In_1684);
nand U4364 (N_4364,In_2744,In_2320);
nor U4365 (N_4365,In_2580,In_2524);
nor U4366 (N_4366,In_1225,In_2209);
or U4367 (N_4367,In_2687,In_18);
nand U4368 (N_4368,In_1080,In_1221);
and U4369 (N_4369,In_2139,In_2533);
nor U4370 (N_4370,In_2929,In_1007);
xnor U4371 (N_4371,In_1837,In_2336);
or U4372 (N_4372,In_2930,In_2209);
nand U4373 (N_4373,In_715,In_2628);
nand U4374 (N_4374,In_2655,In_1956);
nand U4375 (N_4375,In_1342,In_218);
nand U4376 (N_4376,In_1814,In_1114);
or U4377 (N_4377,In_328,In_434);
and U4378 (N_4378,In_2638,In_404);
and U4379 (N_4379,In_1301,In_346);
or U4380 (N_4380,In_1432,In_1063);
nor U4381 (N_4381,In_472,In_1305);
and U4382 (N_4382,In_2156,In_1155);
nand U4383 (N_4383,In_385,In_2077);
xor U4384 (N_4384,In_322,In_1162);
and U4385 (N_4385,In_2346,In_1045);
nor U4386 (N_4386,In_1568,In_2364);
nand U4387 (N_4387,In_2854,In_1504);
or U4388 (N_4388,In_493,In_161);
xor U4389 (N_4389,In_1652,In_1562);
nand U4390 (N_4390,In_2159,In_271);
xnor U4391 (N_4391,In_2035,In_1913);
xor U4392 (N_4392,In_1068,In_738);
nor U4393 (N_4393,In_1851,In_2569);
nor U4394 (N_4394,In_1636,In_2633);
nor U4395 (N_4395,In_2791,In_2593);
or U4396 (N_4396,In_2248,In_2786);
nand U4397 (N_4397,In_2559,In_129);
nor U4398 (N_4398,In_64,In_968);
nor U4399 (N_4399,In_2452,In_2726);
xnor U4400 (N_4400,In_1398,In_1929);
nand U4401 (N_4401,In_2133,In_986);
nand U4402 (N_4402,In_1704,In_2575);
nand U4403 (N_4403,In_52,In_2038);
or U4404 (N_4404,In_1739,In_48);
nor U4405 (N_4405,In_2344,In_2712);
xnor U4406 (N_4406,In_2837,In_464);
or U4407 (N_4407,In_1000,In_1241);
xor U4408 (N_4408,In_1285,In_1223);
or U4409 (N_4409,In_1453,In_485);
or U4410 (N_4410,In_1028,In_2245);
xor U4411 (N_4411,In_1776,In_127);
xnor U4412 (N_4412,In_1623,In_286);
or U4413 (N_4413,In_609,In_336);
nand U4414 (N_4414,In_2479,In_1776);
xnor U4415 (N_4415,In_639,In_75);
nor U4416 (N_4416,In_2451,In_2384);
and U4417 (N_4417,In_1822,In_1876);
nand U4418 (N_4418,In_2284,In_1617);
nand U4419 (N_4419,In_1685,In_1124);
nor U4420 (N_4420,In_867,In_2649);
nand U4421 (N_4421,In_2072,In_300);
nor U4422 (N_4422,In_2269,In_2465);
nor U4423 (N_4423,In_1774,In_2233);
nor U4424 (N_4424,In_454,In_1430);
nand U4425 (N_4425,In_2378,In_1810);
or U4426 (N_4426,In_2414,In_1535);
xnor U4427 (N_4427,In_226,In_1621);
nor U4428 (N_4428,In_2097,In_1586);
nor U4429 (N_4429,In_254,In_1052);
xnor U4430 (N_4430,In_1189,In_2798);
nand U4431 (N_4431,In_2104,In_2947);
and U4432 (N_4432,In_973,In_2021);
nor U4433 (N_4433,In_870,In_355);
and U4434 (N_4434,In_38,In_1900);
nor U4435 (N_4435,In_512,In_1191);
nand U4436 (N_4436,In_573,In_1649);
or U4437 (N_4437,In_2893,In_547);
and U4438 (N_4438,In_2389,In_916);
or U4439 (N_4439,In_379,In_998);
and U4440 (N_4440,In_787,In_2435);
or U4441 (N_4441,In_2834,In_1399);
and U4442 (N_4442,In_1089,In_1821);
nor U4443 (N_4443,In_1799,In_2963);
and U4444 (N_4444,In_2294,In_1818);
nor U4445 (N_4445,In_1147,In_625);
xor U4446 (N_4446,In_2388,In_1941);
or U4447 (N_4447,In_1822,In_1117);
and U4448 (N_4448,In_2935,In_2681);
or U4449 (N_4449,In_1864,In_2795);
nor U4450 (N_4450,In_2801,In_358);
nand U4451 (N_4451,In_2176,In_746);
nand U4452 (N_4452,In_1810,In_320);
and U4453 (N_4453,In_1148,In_534);
and U4454 (N_4454,In_2216,In_1338);
nor U4455 (N_4455,In_1140,In_1580);
nor U4456 (N_4456,In_2297,In_1736);
nor U4457 (N_4457,In_1626,In_273);
nand U4458 (N_4458,In_247,In_76);
and U4459 (N_4459,In_1984,In_1741);
xor U4460 (N_4460,In_2309,In_1088);
or U4461 (N_4461,In_2439,In_673);
nand U4462 (N_4462,In_442,In_382);
or U4463 (N_4463,In_1536,In_1833);
or U4464 (N_4464,In_713,In_2707);
xnor U4465 (N_4465,In_1222,In_19);
xnor U4466 (N_4466,In_1734,In_166);
nand U4467 (N_4467,In_2443,In_312);
and U4468 (N_4468,In_1458,In_1960);
or U4469 (N_4469,In_710,In_1916);
nor U4470 (N_4470,In_2789,In_202);
or U4471 (N_4471,In_1189,In_302);
or U4472 (N_4472,In_2557,In_2930);
or U4473 (N_4473,In_1655,In_1216);
or U4474 (N_4474,In_302,In_2556);
nor U4475 (N_4475,In_2,In_2935);
or U4476 (N_4476,In_1314,In_2743);
or U4477 (N_4477,In_1994,In_460);
and U4478 (N_4478,In_2702,In_2304);
nor U4479 (N_4479,In_557,In_121);
nor U4480 (N_4480,In_2386,In_670);
and U4481 (N_4481,In_308,In_331);
nand U4482 (N_4482,In_920,In_2014);
nor U4483 (N_4483,In_2842,In_810);
or U4484 (N_4484,In_2951,In_768);
or U4485 (N_4485,In_2295,In_1500);
nor U4486 (N_4486,In_2781,In_26);
and U4487 (N_4487,In_1428,In_1867);
xor U4488 (N_4488,In_639,In_347);
xor U4489 (N_4489,In_188,In_382);
or U4490 (N_4490,In_1626,In_1491);
xor U4491 (N_4491,In_2168,In_979);
nor U4492 (N_4492,In_643,In_1309);
nand U4493 (N_4493,In_462,In_2965);
nand U4494 (N_4494,In_207,In_1180);
and U4495 (N_4495,In_451,In_1471);
nand U4496 (N_4496,In_2381,In_1749);
or U4497 (N_4497,In_2528,In_2478);
and U4498 (N_4498,In_2408,In_864);
nand U4499 (N_4499,In_1224,In_764);
or U4500 (N_4500,In_1492,In_1856);
xnor U4501 (N_4501,In_868,In_1251);
and U4502 (N_4502,In_2063,In_2572);
or U4503 (N_4503,In_2873,In_1820);
nor U4504 (N_4504,In_2052,In_2975);
nor U4505 (N_4505,In_263,In_1838);
and U4506 (N_4506,In_1699,In_1169);
nor U4507 (N_4507,In_2012,In_941);
or U4508 (N_4508,In_2145,In_2680);
nor U4509 (N_4509,In_1334,In_32);
and U4510 (N_4510,In_1112,In_407);
and U4511 (N_4511,In_1488,In_304);
nand U4512 (N_4512,In_299,In_2816);
and U4513 (N_4513,In_478,In_2504);
and U4514 (N_4514,In_1636,In_1935);
nor U4515 (N_4515,In_741,In_1226);
or U4516 (N_4516,In_1922,In_1045);
xnor U4517 (N_4517,In_194,In_2627);
and U4518 (N_4518,In_1692,In_526);
nor U4519 (N_4519,In_2169,In_249);
or U4520 (N_4520,In_425,In_433);
xnor U4521 (N_4521,In_1105,In_2671);
or U4522 (N_4522,In_2831,In_1529);
and U4523 (N_4523,In_2724,In_823);
or U4524 (N_4524,In_2681,In_2912);
xnor U4525 (N_4525,In_159,In_1216);
or U4526 (N_4526,In_2681,In_1889);
nor U4527 (N_4527,In_101,In_1437);
nand U4528 (N_4528,In_2997,In_1430);
nor U4529 (N_4529,In_1895,In_268);
or U4530 (N_4530,In_1187,In_392);
nor U4531 (N_4531,In_1489,In_1535);
or U4532 (N_4532,In_193,In_2222);
nand U4533 (N_4533,In_1974,In_2250);
and U4534 (N_4534,In_1418,In_2203);
and U4535 (N_4535,In_1044,In_1182);
nor U4536 (N_4536,In_2803,In_2872);
nor U4537 (N_4537,In_55,In_2250);
and U4538 (N_4538,In_1816,In_2963);
nor U4539 (N_4539,In_2628,In_566);
nor U4540 (N_4540,In_2256,In_796);
and U4541 (N_4541,In_1982,In_1474);
nand U4542 (N_4542,In_2461,In_249);
and U4543 (N_4543,In_2082,In_2406);
xor U4544 (N_4544,In_1551,In_2173);
or U4545 (N_4545,In_7,In_572);
xnor U4546 (N_4546,In_376,In_34);
xor U4547 (N_4547,In_2241,In_723);
xnor U4548 (N_4548,In_2637,In_2246);
nor U4549 (N_4549,In_1938,In_689);
nand U4550 (N_4550,In_1398,In_1071);
nor U4551 (N_4551,In_2662,In_1842);
nor U4552 (N_4552,In_401,In_80);
xor U4553 (N_4553,In_732,In_853);
and U4554 (N_4554,In_1444,In_2699);
xnor U4555 (N_4555,In_827,In_797);
nor U4556 (N_4556,In_89,In_2862);
nor U4557 (N_4557,In_2412,In_162);
nor U4558 (N_4558,In_1019,In_2038);
or U4559 (N_4559,In_10,In_2929);
nand U4560 (N_4560,In_981,In_1358);
and U4561 (N_4561,In_1905,In_2747);
or U4562 (N_4562,In_2972,In_2633);
or U4563 (N_4563,In_1921,In_912);
and U4564 (N_4564,In_2515,In_297);
or U4565 (N_4565,In_1867,In_9);
and U4566 (N_4566,In_2498,In_671);
nand U4567 (N_4567,In_1052,In_679);
xnor U4568 (N_4568,In_1879,In_1732);
xor U4569 (N_4569,In_2940,In_907);
and U4570 (N_4570,In_384,In_1441);
or U4571 (N_4571,In_1088,In_721);
nor U4572 (N_4572,In_2904,In_2077);
and U4573 (N_4573,In_1876,In_2257);
or U4574 (N_4574,In_498,In_2815);
or U4575 (N_4575,In_951,In_283);
and U4576 (N_4576,In_2273,In_2225);
or U4577 (N_4577,In_1638,In_2624);
nor U4578 (N_4578,In_2959,In_896);
nand U4579 (N_4579,In_2620,In_1708);
xor U4580 (N_4580,In_1341,In_78);
and U4581 (N_4581,In_1636,In_1158);
nor U4582 (N_4582,In_1339,In_2952);
or U4583 (N_4583,In_746,In_541);
nand U4584 (N_4584,In_2432,In_136);
nor U4585 (N_4585,In_1822,In_1722);
nor U4586 (N_4586,In_2797,In_2799);
and U4587 (N_4587,In_570,In_2065);
nand U4588 (N_4588,In_1542,In_2323);
and U4589 (N_4589,In_2841,In_507);
nand U4590 (N_4590,In_1488,In_18);
nand U4591 (N_4591,In_2660,In_1486);
nor U4592 (N_4592,In_1031,In_249);
and U4593 (N_4593,In_637,In_2446);
and U4594 (N_4594,In_278,In_2847);
nor U4595 (N_4595,In_718,In_429);
or U4596 (N_4596,In_1551,In_2436);
and U4597 (N_4597,In_305,In_1635);
xnor U4598 (N_4598,In_200,In_1605);
nor U4599 (N_4599,In_1021,In_967);
nand U4600 (N_4600,In_2241,In_2062);
xnor U4601 (N_4601,In_523,In_974);
and U4602 (N_4602,In_1254,In_2610);
and U4603 (N_4603,In_2976,In_274);
or U4604 (N_4604,In_1108,In_2506);
nor U4605 (N_4605,In_1118,In_2345);
nor U4606 (N_4606,In_1634,In_1881);
or U4607 (N_4607,In_2057,In_307);
and U4608 (N_4608,In_2286,In_638);
or U4609 (N_4609,In_905,In_452);
xor U4610 (N_4610,In_1765,In_244);
and U4611 (N_4611,In_2469,In_265);
or U4612 (N_4612,In_2316,In_2447);
nand U4613 (N_4613,In_2248,In_1211);
xnor U4614 (N_4614,In_517,In_2165);
and U4615 (N_4615,In_310,In_2182);
xnor U4616 (N_4616,In_2436,In_1131);
nor U4617 (N_4617,In_676,In_1993);
and U4618 (N_4618,In_649,In_700);
nand U4619 (N_4619,In_1263,In_2139);
and U4620 (N_4620,In_361,In_1377);
nand U4621 (N_4621,In_1913,In_2956);
nand U4622 (N_4622,In_1427,In_895);
nand U4623 (N_4623,In_304,In_1211);
nor U4624 (N_4624,In_2464,In_71);
nand U4625 (N_4625,In_2621,In_959);
or U4626 (N_4626,In_2536,In_1184);
nand U4627 (N_4627,In_2017,In_714);
nor U4628 (N_4628,In_1882,In_341);
xor U4629 (N_4629,In_1360,In_467);
or U4630 (N_4630,In_2929,In_1140);
and U4631 (N_4631,In_2884,In_1228);
or U4632 (N_4632,In_2232,In_780);
and U4633 (N_4633,In_1351,In_1037);
and U4634 (N_4634,In_2794,In_2886);
or U4635 (N_4635,In_1854,In_2765);
nand U4636 (N_4636,In_1613,In_2301);
nor U4637 (N_4637,In_2712,In_2320);
nor U4638 (N_4638,In_973,In_983);
xor U4639 (N_4639,In_1730,In_57);
xor U4640 (N_4640,In_2015,In_2651);
xor U4641 (N_4641,In_1711,In_51);
nor U4642 (N_4642,In_1021,In_2566);
and U4643 (N_4643,In_155,In_452);
nor U4644 (N_4644,In_2249,In_112);
or U4645 (N_4645,In_680,In_2004);
nand U4646 (N_4646,In_816,In_1274);
nand U4647 (N_4647,In_287,In_458);
xor U4648 (N_4648,In_1349,In_496);
or U4649 (N_4649,In_2243,In_2291);
and U4650 (N_4650,In_2172,In_2398);
nor U4651 (N_4651,In_2483,In_335);
nand U4652 (N_4652,In_1972,In_1907);
or U4653 (N_4653,In_2975,In_1005);
and U4654 (N_4654,In_2505,In_2346);
xnor U4655 (N_4655,In_1245,In_114);
nor U4656 (N_4656,In_2985,In_2394);
and U4657 (N_4657,In_2479,In_176);
nor U4658 (N_4658,In_2907,In_71);
nor U4659 (N_4659,In_1511,In_2633);
nand U4660 (N_4660,In_2435,In_1764);
xor U4661 (N_4661,In_118,In_476);
xor U4662 (N_4662,In_1873,In_78);
nor U4663 (N_4663,In_1128,In_489);
nor U4664 (N_4664,In_1584,In_278);
and U4665 (N_4665,In_1808,In_1999);
and U4666 (N_4666,In_2487,In_421);
nor U4667 (N_4667,In_305,In_271);
and U4668 (N_4668,In_2960,In_3);
xor U4669 (N_4669,In_1403,In_2859);
or U4670 (N_4670,In_850,In_1636);
xor U4671 (N_4671,In_2360,In_1609);
nand U4672 (N_4672,In_2686,In_2278);
or U4673 (N_4673,In_1631,In_868);
nor U4674 (N_4674,In_1001,In_2017);
nor U4675 (N_4675,In_2436,In_583);
and U4676 (N_4676,In_381,In_1698);
nor U4677 (N_4677,In_1794,In_1295);
or U4678 (N_4678,In_244,In_1099);
nand U4679 (N_4679,In_475,In_2946);
nor U4680 (N_4680,In_225,In_2174);
xor U4681 (N_4681,In_1226,In_580);
or U4682 (N_4682,In_1962,In_603);
nand U4683 (N_4683,In_726,In_373);
and U4684 (N_4684,In_2083,In_1305);
or U4685 (N_4685,In_632,In_919);
nor U4686 (N_4686,In_1207,In_1336);
or U4687 (N_4687,In_876,In_2662);
nand U4688 (N_4688,In_2664,In_2957);
and U4689 (N_4689,In_2526,In_1381);
nor U4690 (N_4690,In_1429,In_1014);
and U4691 (N_4691,In_2405,In_1731);
or U4692 (N_4692,In_557,In_2511);
xor U4693 (N_4693,In_1284,In_2067);
and U4694 (N_4694,In_806,In_648);
xnor U4695 (N_4695,In_2504,In_2623);
nand U4696 (N_4696,In_2450,In_463);
nand U4697 (N_4697,In_2660,In_1650);
xor U4698 (N_4698,In_495,In_961);
or U4699 (N_4699,In_1407,In_695);
or U4700 (N_4700,In_339,In_369);
nand U4701 (N_4701,In_1790,In_1705);
nand U4702 (N_4702,In_441,In_2251);
nor U4703 (N_4703,In_2871,In_1290);
xnor U4704 (N_4704,In_1582,In_1940);
and U4705 (N_4705,In_2103,In_1170);
or U4706 (N_4706,In_1394,In_1834);
or U4707 (N_4707,In_2124,In_1678);
and U4708 (N_4708,In_715,In_442);
nor U4709 (N_4709,In_1873,In_154);
and U4710 (N_4710,In_1987,In_2744);
nor U4711 (N_4711,In_966,In_2308);
or U4712 (N_4712,In_632,In_1078);
nand U4713 (N_4713,In_1299,In_1412);
nand U4714 (N_4714,In_1432,In_2004);
nand U4715 (N_4715,In_2765,In_815);
and U4716 (N_4716,In_2978,In_222);
and U4717 (N_4717,In_2586,In_783);
nand U4718 (N_4718,In_2628,In_1306);
xnor U4719 (N_4719,In_2355,In_1001);
xor U4720 (N_4720,In_2786,In_1952);
or U4721 (N_4721,In_2138,In_2204);
nand U4722 (N_4722,In_1480,In_2410);
xnor U4723 (N_4723,In_520,In_873);
nor U4724 (N_4724,In_2829,In_2206);
or U4725 (N_4725,In_1200,In_1251);
nor U4726 (N_4726,In_988,In_520);
or U4727 (N_4727,In_1761,In_891);
or U4728 (N_4728,In_301,In_59);
nor U4729 (N_4729,In_1899,In_373);
and U4730 (N_4730,In_2989,In_1646);
nor U4731 (N_4731,In_1369,In_1693);
xor U4732 (N_4732,In_1392,In_1653);
nand U4733 (N_4733,In_1033,In_1553);
nor U4734 (N_4734,In_845,In_1922);
or U4735 (N_4735,In_2700,In_2153);
nor U4736 (N_4736,In_2281,In_220);
xor U4737 (N_4737,In_929,In_813);
nand U4738 (N_4738,In_1209,In_1550);
and U4739 (N_4739,In_1669,In_2362);
xnor U4740 (N_4740,In_556,In_462);
and U4741 (N_4741,In_1091,In_7);
and U4742 (N_4742,In_799,In_475);
nand U4743 (N_4743,In_2718,In_269);
xor U4744 (N_4744,In_1045,In_1105);
nand U4745 (N_4745,In_2151,In_831);
and U4746 (N_4746,In_896,In_965);
or U4747 (N_4747,In_1701,In_818);
xnor U4748 (N_4748,In_2506,In_2049);
or U4749 (N_4749,In_2291,In_2082);
xor U4750 (N_4750,In_457,In_1839);
nand U4751 (N_4751,In_1275,In_2373);
nor U4752 (N_4752,In_2602,In_1738);
xor U4753 (N_4753,In_324,In_2767);
nor U4754 (N_4754,In_1454,In_1278);
and U4755 (N_4755,In_513,In_1495);
xnor U4756 (N_4756,In_1100,In_612);
nand U4757 (N_4757,In_2124,In_560);
nand U4758 (N_4758,In_2888,In_286);
or U4759 (N_4759,In_1898,In_2125);
and U4760 (N_4760,In_1749,In_171);
and U4761 (N_4761,In_1992,In_19);
and U4762 (N_4762,In_1917,In_1552);
and U4763 (N_4763,In_2918,In_277);
and U4764 (N_4764,In_578,In_2210);
nand U4765 (N_4765,In_2696,In_1149);
nor U4766 (N_4766,In_793,In_358);
xor U4767 (N_4767,In_2796,In_71);
xor U4768 (N_4768,In_1539,In_1460);
nor U4769 (N_4769,In_1275,In_1688);
nand U4770 (N_4770,In_2047,In_1827);
or U4771 (N_4771,In_1341,In_1028);
or U4772 (N_4772,In_1060,In_2264);
nor U4773 (N_4773,In_1552,In_969);
and U4774 (N_4774,In_2025,In_667);
nor U4775 (N_4775,In_2607,In_2158);
and U4776 (N_4776,In_2426,In_832);
xnor U4777 (N_4777,In_1781,In_2556);
or U4778 (N_4778,In_376,In_2466);
and U4779 (N_4779,In_2882,In_195);
nor U4780 (N_4780,In_2946,In_1290);
xnor U4781 (N_4781,In_222,In_203);
or U4782 (N_4782,In_2335,In_38);
or U4783 (N_4783,In_1090,In_2307);
xor U4784 (N_4784,In_1368,In_2723);
and U4785 (N_4785,In_248,In_707);
nor U4786 (N_4786,In_1288,In_2653);
or U4787 (N_4787,In_2630,In_863);
or U4788 (N_4788,In_517,In_1260);
and U4789 (N_4789,In_2767,In_233);
nor U4790 (N_4790,In_1676,In_2922);
xnor U4791 (N_4791,In_1657,In_610);
nand U4792 (N_4792,In_1810,In_737);
and U4793 (N_4793,In_2289,In_2001);
xor U4794 (N_4794,In_767,In_2860);
and U4795 (N_4795,In_543,In_721);
and U4796 (N_4796,In_1595,In_7);
and U4797 (N_4797,In_1941,In_1215);
and U4798 (N_4798,In_1992,In_186);
nor U4799 (N_4799,In_1281,In_2678);
nand U4800 (N_4800,In_2945,In_2152);
nor U4801 (N_4801,In_1013,In_779);
xor U4802 (N_4802,In_1898,In_540);
xnor U4803 (N_4803,In_471,In_2836);
xor U4804 (N_4804,In_250,In_2851);
and U4805 (N_4805,In_2564,In_986);
or U4806 (N_4806,In_2319,In_1864);
or U4807 (N_4807,In_2254,In_1276);
or U4808 (N_4808,In_1796,In_1041);
or U4809 (N_4809,In_1927,In_2398);
xor U4810 (N_4810,In_2592,In_1966);
or U4811 (N_4811,In_1696,In_434);
xnor U4812 (N_4812,In_2997,In_2775);
or U4813 (N_4813,In_950,In_772);
and U4814 (N_4814,In_515,In_2682);
nor U4815 (N_4815,In_1346,In_87);
xor U4816 (N_4816,In_2381,In_497);
xnor U4817 (N_4817,In_2810,In_983);
or U4818 (N_4818,In_647,In_1028);
xnor U4819 (N_4819,In_2273,In_1467);
and U4820 (N_4820,In_203,In_1002);
nor U4821 (N_4821,In_992,In_77);
or U4822 (N_4822,In_2266,In_983);
xor U4823 (N_4823,In_2277,In_325);
xor U4824 (N_4824,In_2912,In_2326);
nor U4825 (N_4825,In_796,In_79);
or U4826 (N_4826,In_2448,In_1877);
nor U4827 (N_4827,In_2074,In_1431);
xnor U4828 (N_4828,In_2525,In_1403);
or U4829 (N_4829,In_1691,In_874);
nor U4830 (N_4830,In_2440,In_2240);
xnor U4831 (N_4831,In_2382,In_2189);
xor U4832 (N_4832,In_1083,In_1649);
nor U4833 (N_4833,In_2419,In_498);
or U4834 (N_4834,In_1450,In_215);
and U4835 (N_4835,In_706,In_1105);
xnor U4836 (N_4836,In_682,In_1739);
or U4837 (N_4837,In_2206,In_4);
xor U4838 (N_4838,In_2241,In_2999);
nor U4839 (N_4839,In_1590,In_324);
xor U4840 (N_4840,In_2090,In_1610);
or U4841 (N_4841,In_1487,In_2616);
nor U4842 (N_4842,In_218,In_97);
nand U4843 (N_4843,In_2446,In_2199);
nor U4844 (N_4844,In_814,In_2530);
xnor U4845 (N_4845,In_2900,In_1054);
nand U4846 (N_4846,In_2843,In_2029);
and U4847 (N_4847,In_1221,In_2351);
nand U4848 (N_4848,In_2168,In_1600);
and U4849 (N_4849,In_358,In_442);
and U4850 (N_4850,In_1006,In_2265);
or U4851 (N_4851,In_2622,In_1816);
and U4852 (N_4852,In_2435,In_2935);
and U4853 (N_4853,In_2982,In_1286);
nor U4854 (N_4854,In_2573,In_1846);
nand U4855 (N_4855,In_653,In_1045);
nor U4856 (N_4856,In_2265,In_2095);
and U4857 (N_4857,In_2318,In_74);
nor U4858 (N_4858,In_1083,In_2503);
xnor U4859 (N_4859,In_827,In_2687);
or U4860 (N_4860,In_992,In_2488);
nand U4861 (N_4861,In_1991,In_2369);
and U4862 (N_4862,In_1000,In_849);
xor U4863 (N_4863,In_43,In_1921);
or U4864 (N_4864,In_909,In_346);
or U4865 (N_4865,In_1941,In_1742);
and U4866 (N_4866,In_2449,In_1734);
nor U4867 (N_4867,In_1692,In_1738);
or U4868 (N_4868,In_510,In_1243);
nand U4869 (N_4869,In_1075,In_141);
nand U4870 (N_4870,In_2290,In_229);
nor U4871 (N_4871,In_1191,In_1152);
xor U4872 (N_4872,In_567,In_2693);
or U4873 (N_4873,In_1523,In_2856);
xor U4874 (N_4874,In_1698,In_2353);
and U4875 (N_4875,In_257,In_544);
xor U4876 (N_4876,In_649,In_1191);
and U4877 (N_4877,In_856,In_1681);
nor U4878 (N_4878,In_2423,In_2337);
nor U4879 (N_4879,In_2907,In_2659);
nor U4880 (N_4880,In_1712,In_377);
or U4881 (N_4881,In_1422,In_569);
nand U4882 (N_4882,In_1124,In_2487);
and U4883 (N_4883,In_477,In_534);
or U4884 (N_4884,In_760,In_667);
nand U4885 (N_4885,In_1992,In_245);
nor U4886 (N_4886,In_1502,In_2200);
and U4887 (N_4887,In_906,In_1695);
nor U4888 (N_4888,In_223,In_2082);
nor U4889 (N_4889,In_434,In_91);
nor U4890 (N_4890,In_870,In_523);
nor U4891 (N_4891,In_988,In_1049);
xnor U4892 (N_4892,In_2388,In_16);
or U4893 (N_4893,In_1704,In_1361);
xor U4894 (N_4894,In_260,In_1042);
nand U4895 (N_4895,In_1058,In_108);
nor U4896 (N_4896,In_1988,In_1237);
nand U4897 (N_4897,In_2909,In_2947);
or U4898 (N_4898,In_805,In_1719);
nor U4899 (N_4899,In_2516,In_806);
nor U4900 (N_4900,In_1216,In_2181);
and U4901 (N_4901,In_2256,In_1825);
and U4902 (N_4902,In_355,In_2687);
nor U4903 (N_4903,In_1354,In_1538);
nand U4904 (N_4904,In_665,In_802);
or U4905 (N_4905,In_1313,In_2070);
nand U4906 (N_4906,In_1682,In_2290);
and U4907 (N_4907,In_103,In_2844);
nand U4908 (N_4908,In_366,In_987);
xor U4909 (N_4909,In_371,In_2957);
xnor U4910 (N_4910,In_1547,In_2375);
and U4911 (N_4911,In_1443,In_3);
xnor U4912 (N_4912,In_2057,In_1503);
or U4913 (N_4913,In_2507,In_2050);
or U4914 (N_4914,In_1925,In_2556);
and U4915 (N_4915,In_2359,In_298);
and U4916 (N_4916,In_115,In_234);
nor U4917 (N_4917,In_977,In_2762);
xor U4918 (N_4918,In_1221,In_2296);
or U4919 (N_4919,In_1171,In_1770);
or U4920 (N_4920,In_820,In_185);
nand U4921 (N_4921,In_2886,In_2583);
nor U4922 (N_4922,In_1151,In_2333);
nand U4923 (N_4923,In_2820,In_2581);
nor U4924 (N_4924,In_959,In_2221);
or U4925 (N_4925,In_2687,In_619);
nand U4926 (N_4926,In_1043,In_2702);
and U4927 (N_4927,In_121,In_1796);
nand U4928 (N_4928,In_2309,In_1028);
nor U4929 (N_4929,In_1988,In_1295);
nand U4930 (N_4930,In_708,In_939);
or U4931 (N_4931,In_728,In_299);
xor U4932 (N_4932,In_2664,In_1953);
and U4933 (N_4933,In_2085,In_261);
or U4934 (N_4934,In_1007,In_2083);
xor U4935 (N_4935,In_2074,In_2354);
nor U4936 (N_4936,In_549,In_769);
and U4937 (N_4937,In_1292,In_2633);
nor U4938 (N_4938,In_1062,In_1989);
xor U4939 (N_4939,In_2156,In_480);
nand U4940 (N_4940,In_2394,In_711);
nand U4941 (N_4941,In_194,In_940);
nor U4942 (N_4942,In_1962,In_276);
and U4943 (N_4943,In_321,In_2690);
nor U4944 (N_4944,In_1025,In_467);
nor U4945 (N_4945,In_505,In_287);
nor U4946 (N_4946,In_2737,In_2672);
nor U4947 (N_4947,In_1859,In_473);
xnor U4948 (N_4948,In_2515,In_2945);
and U4949 (N_4949,In_1795,In_692);
nor U4950 (N_4950,In_1031,In_1404);
nor U4951 (N_4951,In_1865,In_467);
xor U4952 (N_4952,In_724,In_1133);
nand U4953 (N_4953,In_1134,In_2873);
and U4954 (N_4954,In_296,In_180);
or U4955 (N_4955,In_2555,In_1697);
xor U4956 (N_4956,In_2145,In_2940);
or U4957 (N_4957,In_2590,In_2846);
nor U4958 (N_4958,In_2366,In_2674);
and U4959 (N_4959,In_706,In_2753);
or U4960 (N_4960,In_2140,In_39);
nor U4961 (N_4961,In_1557,In_1217);
xor U4962 (N_4962,In_2161,In_2483);
xnor U4963 (N_4963,In_2583,In_1441);
or U4964 (N_4964,In_2213,In_1590);
nor U4965 (N_4965,In_382,In_1938);
xor U4966 (N_4966,In_1946,In_1753);
xnor U4967 (N_4967,In_2254,In_2693);
nor U4968 (N_4968,In_1717,In_211);
and U4969 (N_4969,In_2749,In_284);
xor U4970 (N_4970,In_803,In_452);
xor U4971 (N_4971,In_2140,In_427);
and U4972 (N_4972,In_1989,In_488);
and U4973 (N_4973,In_1901,In_744);
nor U4974 (N_4974,In_1803,In_879);
xor U4975 (N_4975,In_287,In_753);
xnor U4976 (N_4976,In_2539,In_2005);
nand U4977 (N_4977,In_1612,In_2719);
xor U4978 (N_4978,In_1432,In_2739);
nand U4979 (N_4979,In_812,In_263);
and U4980 (N_4980,In_2109,In_574);
or U4981 (N_4981,In_1733,In_1149);
nor U4982 (N_4982,In_330,In_205);
nand U4983 (N_4983,In_2605,In_1208);
nand U4984 (N_4984,In_1673,In_310);
xor U4985 (N_4985,In_1217,In_609);
or U4986 (N_4986,In_2627,In_69);
nand U4987 (N_4987,In_2291,In_2920);
xnor U4988 (N_4988,In_2988,In_952);
nor U4989 (N_4989,In_18,In_912);
xor U4990 (N_4990,In_1087,In_687);
nand U4991 (N_4991,In_1210,In_814);
or U4992 (N_4992,In_1210,In_1135);
nor U4993 (N_4993,In_955,In_2806);
xnor U4994 (N_4994,In_577,In_1581);
and U4995 (N_4995,In_134,In_2129);
or U4996 (N_4996,In_1251,In_1001);
or U4997 (N_4997,In_1859,In_514);
xor U4998 (N_4998,In_105,In_1905);
nor U4999 (N_4999,In_1307,In_419);
and U5000 (N_5000,N_1603,N_2263);
xor U5001 (N_5001,N_1754,N_243);
nand U5002 (N_5002,N_2938,N_1973);
or U5003 (N_5003,N_801,N_3298);
and U5004 (N_5004,N_386,N_560);
nand U5005 (N_5005,N_1861,N_4552);
and U5006 (N_5006,N_670,N_722);
or U5007 (N_5007,N_3900,N_4508);
and U5008 (N_5008,N_2043,N_1422);
and U5009 (N_5009,N_3536,N_4251);
xnor U5010 (N_5010,N_4503,N_3751);
or U5011 (N_5011,N_3540,N_2494);
and U5012 (N_5012,N_2234,N_3210);
or U5013 (N_5013,N_3743,N_4634);
nor U5014 (N_5014,N_3926,N_1550);
or U5015 (N_5015,N_1386,N_3613);
or U5016 (N_5016,N_417,N_3214);
and U5017 (N_5017,N_453,N_4456);
xnor U5018 (N_5018,N_4506,N_1736);
and U5019 (N_5019,N_2436,N_1114);
xor U5020 (N_5020,N_2703,N_1119);
nor U5021 (N_5021,N_2470,N_1172);
and U5022 (N_5022,N_1845,N_3941);
nand U5023 (N_5023,N_3645,N_2911);
or U5024 (N_5024,N_2142,N_2438);
or U5025 (N_5025,N_975,N_418);
or U5026 (N_5026,N_2073,N_1489);
or U5027 (N_5027,N_2336,N_2616);
and U5028 (N_5028,N_3428,N_816);
xor U5029 (N_5029,N_4910,N_4366);
or U5030 (N_5030,N_1131,N_2052);
and U5031 (N_5031,N_3239,N_2491);
xnor U5032 (N_5032,N_2759,N_319);
nor U5033 (N_5033,N_1077,N_110);
and U5034 (N_5034,N_885,N_3993);
and U5035 (N_5035,N_4039,N_498);
and U5036 (N_5036,N_1370,N_1536);
nor U5037 (N_5037,N_1539,N_1642);
xor U5038 (N_5038,N_2187,N_1856);
or U5039 (N_5039,N_836,N_3716);
and U5040 (N_5040,N_732,N_4472);
nor U5041 (N_5041,N_313,N_3960);
nor U5042 (N_5042,N_1883,N_4502);
and U5043 (N_5043,N_4872,N_4498);
nand U5044 (N_5044,N_2049,N_389);
xnor U5045 (N_5045,N_1915,N_1769);
and U5046 (N_5046,N_3190,N_2023);
nand U5047 (N_5047,N_4428,N_3184);
xor U5048 (N_5048,N_2634,N_989);
xnor U5049 (N_5049,N_4580,N_4709);
nand U5050 (N_5050,N_3476,N_1208);
nor U5051 (N_5051,N_4857,N_4220);
and U5052 (N_5052,N_4296,N_3970);
and U5053 (N_5053,N_1542,N_1535);
and U5054 (N_5054,N_3124,N_24);
nand U5055 (N_5055,N_3162,N_2762);
or U5056 (N_5056,N_3107,N_4632);
xnor U5057 (N_5057,N_2763,N_3882);
or U5058 (N_5058,N_4358,N_3050);
nand U5059 (N_5059,N_101,N_667);
or U5060 (N_5060,N_233,N_3617);
and U5061 (N_5061,N_3318,N_596);
or U5062 (N_5062,N_1663,N_1433);
nor U5063 (N_5063,N_574,N_3314);
and U5064 (N_5064,N_2445,N_912);
xnor U5065 (N_5065,N_261,N_617);
and U5066 (N_5066,N_1320,N_4254);
xor U5067 (N_5067,N_2061,N_370);
nand U5068 (N_5068,N_3752,N_4411);
and U5069 (N_5069,N_705,N_628);
nand U5070 (N_5070,N_1302,N_390);
nor U5071 (N_5071,N_723,N_4669);
and U5072 (N_5072,N_3279,N_1864);
nor U5073 (N_5073,N_3120,N_3505);
or U5074 (N_5074,N_2287,N_4998);
nor U5075 (N_5075,N_803,N_982);
nand U5076 (N_5076,N_3383,N_22);
xnor U5077 (N_5077,N_2104,N_4953);
nand U5078 (N_5078,N_4515,N_2385);
xor U5079 (N_5079,N_4949,N_3621);
or U5080 (N_5080,N_2246,N_127);
xnor U5081 (N_5081,N_3666,N_3434);
and U5082 (N_5082,N_1155,N_3932);
xor U5083 (N_5083,N_4501,N_1288);
xor U5084 (N_5084,N_4255,N_1718);
and U5085 (N_5085,N_4952,N_1504);
nor U5086 (N_5086,N_2890,N_3290);
and U5087 (N_5087,N_1395,N_1076);
xor U5088 (N_5088,N_4649,N_2272);
nor U5089 (N_5089,N_1073,N_2513);
or U5090 (N_5090,N_2308,N_3856);
nor U5091 (N_5091,N_4627,N_2907);
and U5092 (N_5092,N_4828,N_1026);
xor U5093 (N_5093,N_1782,N_4664);
and U5094 (N_5094,N_3216,N_4215);
xnor U5095 (N_5095,N_4125,N_4321);
nand U5096 (N_5096,N_4435,N_1831);
or U5097 (N_5097,N_655,N_4665);
nor U5098 (N_5098,N_2430,N_4855);
nor U5099 (N_5099,N_3069,N_2376);
or U5100 (N_5100,N_1707,N_4354);
xor U5101 (N_5101,N_232,N_762);
and U5102 (N_5102,N_4914,N_778);
or U5103 (N_5103,N_1356,N_3879);
nor U5104 (N_5104,N_4858,N_4476);
and U5105 (N_5105,N_303,N_4920);
or U5106 (N_5106,N_624,N_2047);
or U5107 (N_5107,N_606,N_2783);
xor U5108 (N_5108,N_179,N_4063);
xnor U5109 (N_5109,N_3673,N_2526);
or U5110 (N_5110,N_1733,N_2480);
nand U5111 (N_5111,N_3165,N_2887);
or U5112 (N_5112,N_831,N_3683);
nand U5113 (N_5113,N_4058,N_2979);
xor U5114 (N_5114,N_1054,N_1417);
and U5115 (N_5115,N_3401,N_4120);
nand U5116 (N_5116,N_2975,N_4462);
xnor U5117 (N_5117,N_2454,N_4530);
xnor U5118 (N_5118,N_766,N_1963);
nand U5119 (N_5119,N_2925,N_4014);
and U5120 (N_5120,N_3459,N_2476);
xor U5121 (N_5121,N_2229,N_2578);
xor U5122 (N_5122,N_1450,N_3034);
or U5123 (N_5123,N_3692,N_2443);
nand U5124 (N_5124,N_4198,N_586);
xor U5125 (N_5125,N_4277,N_3320);
nor U5126 (N_5126,N_33,N_549);
and U5127 (N_5127,N_1239,N_266);
or U5128 (N_5128,N_822,N_4110);
nand U5129 (N_5129,N_966,N_2138);
and U5130 (N_5130,N_1652,N_3354);
nor U5131 (N_5131,N_2331,N_4942);
nand U5132 (N_5132,N_3491,N_3470);
and U5133 (N_5133,N_1388,N_4867);
xnor U5134 (N_5134,N_4201,N_4104);
nand U5135 (N_5135,N_113,N_2825);
xnor U5136 (N_5136,N_951,N_4599);
nand U5137 (N_5137,N_4809,N_1237);
nor U5138 (N_5138,N_3352,N_3292);
and U5139 (N_5139,N_4701,N_3251);
nand U5140 (N_5140,N_2201,N_2420);
nand U5141 (N_5141,N_4688,N_891);
nor U5142 (N_5142,N_1464,N_1214);
nor U5143 (N_5143,N_1621,N_1123);
nor U5144 (N_5144,N_534,N_4094);
nor U5145 (N_5145,N_868,N_1735);
nor U5146 (N_5146,N_2679,N_1454);
xnor U5147 (N_5147,N_2714,N_581);
and U5148 (N_5148,N_2481,N_1381);
xnor U5149 (N_5149,N_2275,N_1322);
xor U5150 (N_5150,N_2717,N_1284);
and U5151 (N_5151,N_1108,N_3146);
and U5152 (N_5152,N_553,N_1605);
nand U5153 (N_5153,N_1778,N_2561);
and U5154 (N_5154,N_2942,N_3535);
and U5155 (N_5155,N_4533,N_4330);
nand U5156 (N_5156,N_308,N_4438);
xnor U5157 (N_5157,N_3492,N_1439);
or U5158 (N_5158,N_2035,N_2670);
or U5159 (N_5159,N_3293,N_1483);
nand U5160 (N_5160,N_3227,N_4240);
and U5161 (N_5161,N_3614,N_3112);
or U5162 (N_5162,N_2610,N_282);
xnor U5163 (N_5163,N_2784,N_1136);
nand U5164 (N_5164,N_324,N_4864);
nand U5165 (N_5165,N_4710,N_4234);
nand U5166 (N_5166,N_4360,N_945);
or U5167 (N_5167,N_2317,N_4990);
nor U5168 (N_5168,N_1360,N_2678);
nor U5169 (N_5169,N_1798,N_2901);
and U5170 (N_5170,N_58,N_2909);
xnor U5171 (N_5171,N_3678,N_784);
nor U5172 (N_5172,N_4304,N_4658);
or U5173 (N_5173,N_4854,N_3129);
xnor U5174 (N_5174,N_2007,N_582);
nand U5175 (N_5175,N_4291,N_4294);
nor U5176 (N_5176,N_3894,N_3807);
and U5177 (N_5177,N_1152,N_2194);
and U5178 (N_5178,N_395,N_347);
and U5179 (N_5179,N_4008,N_3203);
xor U5180 (N_5180,N_2843,N_2130);
xnor U5181 (N_5181,N_1977,N_3761);
xnor U5182 (N_5182,N_1293,N_3878);
nor U5183 (N_5183,N_4205,N_4779);
nor U5184 (N_5184,N_1746,N_3113);
nor U5185 (N_5185,N_4243,N_218);
and U5186 (N_5186,N_4547,N_3631);
or U5187 (N_5187,N_1955,N_988);
or U5188 (N_5188,N_2163,N_4421);
and U5189 (N_5189,N_4763,N_163);
or U5190 (N_5190,N_1757,N_4662);
xor U5191 (N_5191,N_1255,N_387);
xnor U5192 (N_5192,N_2583,N_2562);
or U5193 (N_5193,N_4646,N_2157);
nor U5194 (N_5194,N_341,N_1683);
or U5195 (N_5195,N_2434,N_1497);
nand U5196 (N_5196,N_3606,N_1412);
xor U5197 (N_5197,N_4225,N_3099);
xnor U5198 (N_5198,N_3179,N_713);
and U5199 (N_5199,N_4250,N_4651);
and U5200 (N_5200,N_383,N_4168);
and U5201 (N_5201,N_1227,N_877);
nor U5202 (N_5202,N_4538,N_787);
nand U5203 (N_5203,N_4762,N_964);
nor U5204 (N_5204,N_4932,N_149);
nor U5205 (N_5205,N_3779,N_2820);
and U5206 (N_5206,N_1,N_3685);
xor U5207 (N_5207,N_597,N_1133);
nor U5208 (N_5208,N_2193,N_2700);
nand U5209 (N_5209,N_3147,N_4066);
and U5210 (N_5210,N_2113,N_2642);
and U5211 (N_5211,N_62,N_1614);
or U5212 (N_5212,N_3035,N_753);
nand U5213 (N_5213,N_694,N_1870);
xor U5214 (N_5214,N_3705,N_1547);
nor U5215 (N_5215,N_4208,N_4761);
xor U5216 (N_5216,N_3925,N_941);
nand U5217 (N_5217,N_4299,N_2335);
nand U5218 (N_5218,N_806,N_1444);
xor U5219 (N_5219,N_804,N_16);
nand U5220 (N_5220,N_2511,N_4442);
or U5221 (N_5221,N_1598,N_2903);
or U5222 (N_5222,N_2731,N_2852);
xnor U5223 (N_5223,N_4846,N_2015);
nand U5224 (N_5224,N_2967,N_4840);
nand U5225 (N_5225,N_981,N_933);
xnor U5226 (N_5226,N_1256,N_2953);
or U5227 (N_5227,N_819,N_554);
nand U5228 (N_5228,N_176,N_2338);
and U5229 (N_5229,N_3132,N_2145);
nand U5230 (N_5230,N_3054,N_2000);
xnor U5231 (N_5231,N_2917,N_4001);
xor U5232 (N_5232,N_1341,N_3805);
or U5233 (N_5233,N_4405,N_1771);
nand U5234 (N_5234,N_4466,N_3951);
and U5235 (N_5235,N_2400,N_2257);
or U5236 (N_5236,N_4954,N_1587);
nor U5237 (N_5237,N_707,N_2418);
or U5238 (N_5238,N_2854,N_4043);
nand U5239 (N_5239,N_3379,N_3188);
xor U5240 (N_5240,N_283,N_870);
nand U5241 (N_5241,N_4751,N_2960);
nand U5242 (N_5242,N_4156,N_4876);
xnor U5243 (N_5243,N_4578,N_284);
xor U5244 (N_5244,N_4320,N_807);
nand U5245 (N_5245,N_4248,N_2318);
xor U5246 (N_5246,N_4326,N_3018);
and U5247 (N_5247,N_1182,N_1801);
nand U5248 (N_5248,N_4672,N_4592);
xor U5249 (N_5249,N_2259,N_3710);
and U5250 (N_5250,N_2726,N_3270);
nand U5251 (N_5251,N_2254,N_1717);
nand U5252 (N_5252,N_2880,N_2196);
or U5253 (N_5253,N_633,N_3398);
nor U5254 (N_5254,N_3387,N_2135);
and U5255 (N_5255,N_4244,N_639);
nor U5256 (N_5256,N_4222,N_1626);
xnor U5257 (N_5257,N_493,N_2785);
or U5258 (N_5258,N_1634,N_866);
or U5259 (N_5259,N_971,N_1151);
nand U5260 (N_5260,N_1996,N_768);
nor U5261 (N_5261,N_4095,N_858);
xor U5262 (N_5262,N_2098,N_3062);
nand U5263 (N_5263,N_4021,N_4415);
nor U5264 (N_5264,N_748,N_446);
or U5265 (N_5265,N_4084,N_2268);
and U5266 (N_5266,N_1203,N_4929);
xnor U5267 (N_5267,N_1134,N_2122);
and U5268 (N_5268,N_2732,N_643);
and U5269 (N_5269,N_4830,N_448);
nand U5270 (N_5270,N_1638,N_1958);
and U5271 (N_5271,N_3944,N_350);
xor U5272 (N_5272,N_2985,N_2691);
nor U5273 (N_5273,N_1460,N_3757);
nor U5274 (N_5274,N_3711,N_3565);
xor U5275 (N_5275,N_2984,N_1065);
xnor U5276 (N_5276,N_3080,N_2197);
or U5277 (N_5277,N_3820,N_4049);
xor U5278 (N_5278,N_3955,N_2564);
and U5279 (N_5279,N_1471,N_2111);
and U5280 (N_5280,N_367,N_2674);
xor U5281 (N_5281,N_1919,N_1327);
nor U5282 (N_5282,N_3369,N_3224);
and U5283 (N_5283,N_3356,N_3760);
or U5284 (N_5284,N_603,N_1546);
nand U5285 (N_5285,N_193,N_4605);
and U5286 (N_5286,N_1879,N_754);
nand U5287 (N_5287,N_364,N_1223);
or U5288 (N_5288,N_2151,N_1466);
xnor U5289 (N_5289,N_1616,N_1731);
and U5290 (N_5290,N_2154,N_1581);
nor U5291 (N_5291,N_4433,N_345);
and U5292 (N_5292,N_136,N_4102);
or U5293 (N_5293,N_4394,N_4841);
nor U5294 (N_5294,N_3867,N_4406);
nand U5295 (N_5295,N_1301,N_2776);
and U5296 (N_5296,N_528,N_1312);
nor U5297 (N_5297,N_4612,N_3774);
nand U5298 (N_5298,N_467,N_3664);
or U5299 (N_5299,N_4484,N_380);
nor U5300 (N_5300,N_644,N_561);
and U5301 (N_5301,N_1991,N_1138);
nor U5302 (N_5302,N_3472,N_3885);
or U5303 (N_5303,N_3667,N_2657);
or U5304 (N_5304,N_4911,N_541);
nor U5305 (N_5305,N_4455,N_1154);
or U5306 (N_5306,N_1604,N_4853);
and U5307 (N_5307,N_2805,N_857);
nand U5308 (N_5308,N_985,N_3351);
xor U5309 (N_5309,N_4280,N_2036);
or U5310 (N_5310,N_4713,N_2658);
and U5311 (N_5311,N_1825,N_2651);
nand U5312 (N_5312,N_247,N_1687);
or U5313 (N_5313,N_2830,N_627);
xnor U5314 (N_5314,N_4711,N_3136);
xnor U5315 (N_5315,N_1384,N_135);
nor U5316 (N_5316,N_2577,N_4670);
nor U5317 (N_5317,N_4888,N_2581);
nand U5318 (N_5318,N_4844,N_3432);
nor U5319 (N_5319,N_1946,N_1226);
nand U5320 (N_5320,N_3304,N_3204);
nand U5321 (N_5321,N_3178,N_1660);
and U5322 (N_5322,N_3501,N_2373);
and U5323 (N_5323,N_3082,N_1531);
xor U5324 (N_5324,N_3886,N_2757);
and U5325 (N_5325,N_4226,N_4544);
and U5326 (N_5326,N_4631,N_4884);
or U5327 (N_5327,N_2845,N_1708);
and U5328 (N_5328,N_1308,N_1376);
or U5329 (N_5329,N_1647,N_4359);
nor U5330 (N_5330,N_436,N_3923);
or U5331 (N_5331,N_536,N_2472);
nor U5332 (N_5332,N_407,N_433);
nand U5333 (N_5333,N_3015,N_1624);
xor U5334 (N_5334,N_4504,N_2375);
nand U5335 (N_5335,N_1636,N_3185);
nor U5336 (N_5336,N_3707,N_4989);
xnor U5337 (N_5337,N_1096,N_4388);
or U5338 (N_5338,N_4047,N_3229);
nor U5339 (N_5339,N_2001,N_3530);
or U5340 (N_5340,N_4774,N_2221);
xor U5341 (N_5341,N_2238,N_2332);
or U5342 (N_5342,N_4402,N_965);
and U5343 (N_5343,N_2598,N_2878);
or U5344 (N_5344,N_3608,N_539);
or U5345 (N_5345,N_3969,N_575);
nand U5346 (N_5346,N_4069,N_1995);
nor U5347 (N_5347,N_1519,N_3708);
or U5348 (N_5348,N_2815,N_1704);
xnor U5349 (N_5349,N_4370,N_2681);
nor U5350 (N_5350,N_4568,N_2499);
nor U5351 (N_5351,N_691,N_3934);
xnor U5352 (N_5352,N_1601,N_1276);
and U5353 (N_5353,N_4965,N_2223);
nor U5354 (N_5354,N_3950,N_4787);
or U5355 (N_5355,N_2993,N_4906);
or U5356 (N_5356,N_1305,N_4374);
and U5357 (N_5357,N_1538,N_2068);
nand U5358 (N_5358,N_4452,N_4556);
or U5359 (N_5359,N_3482,N_683);
nand U5360 (N_5360,N_2628,N_1416);
or U5361 (N_5361,N_3755,N_1415);
or U5362 (N_5362,N_1016,N_287);
nor U5363 (N_5363,N_2339,N_1495);
xnor U5364 (N_5364,N_1374,N_3556);
nor U5365 (N_5365,N_2702,N_702);
nand U5366 (N_5366,N_4186,N_2675);
and U5367 (N_5367,N_4868,N_4349);
nor U5368 (N_5368,N_4390,N_3338);
xnor U5369 (N_5369,N_906,N_2233);
nor U5370 (N_5370,N_1661,N_4939);
nand U5371 (N_5371,N_3390,N_379);
xnor U5372 (N_5372,N_4837,N_3948);
nand U5373 (N_5373,N_229,N_3739);
nor U5374 (N_5374,N_1455,N_4702);
or U5375 (N_5375,N_3713,N_2032);
nand U5376 (N_5376,N_3759,N_4542);
xnor U5377 (N_5377,N_1901,N_4909);
and U5378 (N_5378,N_2319,N_177);
nor U5379 (N_5379,N_3087,N_3674);
nand U5380 (N_5380,N_1938,N_2667);
and U5381 (N_5381,N_4931,N_4015);
and U5382 (N_5382,N_4142,N_2698);
nand U5383 (N_5383,N_1418,N_957);
nor U5384 (N_5384,N_1741,N_85);
nand U5385 (N_5385,N_2071,N_1499);
xnor U5386 (N_5386,N_2758,N_2977);
xor U5387 (N_5387,N_96,N_2416);
nand U5388 (N_5388,N_4306,N_4356);
nor U5389 (N_5389,N_1654,N_3931);
nand U5390 (N_5390,N_1025,N_2378);
nand U5391 (N_5391,N_3093,N_356);
nand U5392 (N_5392,N_4959,N_144);
xor U5393 (N_5393,N_3873,N_2177);
nand U5394 (N_5394,N_788,N_4573);
xor U5395 (N_5395,N_2837,N_2247);
or U5396 (N_5396,N_860,N_3478);
or U5397 (N_5397,N_1484,N_211);
nand U5398 (N_5398,N_1192,N_66);
nor U5399 (N_5399,N_4625,N_4179);
and U5400 (N_5400,N_2755,N_2540);
and U5401 (N_5401,N_990,N_3189);
and U5402 (N_5402,N_974,N_4159);
or U5403 (N_5403,N_2364,N_4068);
nand U5404 (N_5404,N_4564,N_993);
or U5405 (N_5405,N_550,N_2870);
xor U5406 (N_5406,N_4293,N_4638);
xor U5407 (N_5407,N_246,N_589);
xor U5408 (N_5408,N_2112,N_1997);
xnor U5409 (N_5409,N_3975,N_3067);
or U5410 (N_5410,N_3850,N_2970);
xnor U5411 (N_5411,N_2595,N_2884);
xnor U5412 (N_5412,N_422,N_3231);
nor U5413 (N_5413,N_786,N_2764);
and U5414 (N_5414,N_286,N_2627);
nor U5415 (N_5415,N_4913,N_2411);
xor U5416 (N_5416,N_1569,N_1074);
nor U5417 (N_5417,N_240,N_2871);
nand U5418 (N_5418,N_2467,N_1591);
nand U5419 (N_5419,N_1622,N_2095);
xnor U5420 (N_5420,N_2934,N_484);
or U5421 (N_5421,N_3972,N_4712);
and U5422 (N_5422,N_4726,N_1665);
nor U5423 (N_5423,N_4727,N_4975);
nand U5424 (N_5424,N_1606,N_2790);
nand U5425 (N_5425,N_1103,N_1004);
xnor U5426 (N_5426,N_882,N_4191);
nand U5427 (N_5427,N_4447,N_1045);
and U5428 (N_5428,N_2300,N_2180);
and U5429 (N_5429,N_4811,N_4941);
xor U5430 (N_5430,N_2816,N_3377);
nand U5431 (N_5431,N_1878,N_4901);
nor U5432 (N_5432,N_3966,N_2722);
nor U5433 (N_5433,N_1686,N_1165);
and U5434 (N_5434,N_3819,N_2127);
or U5435 (N_5435,N_1029,N_1545);
and U5436 (N_5436,N_3722,N_2106);
xnor U5437 (N_5437,N_717,N_4892);
nor U5438 (N_5438,N_1964,N_3717);
and U5439 (N_5439,N_120,N_2159);
and U5440 (N_5440,N_2281,N_3917);
xor U5441 (N_5441,N_1582,N_3471);
nand U5442 (N_5442,N_2236,N_2639);
nand U5443 (N_5443,N_3776,N_393);
or U5444 (N_5444,N_692,N_689);
nand U5445 (N_5445,N_419,N_506);
nand U5446 (N_5446,N_2524,N_3289);
xor U5447 (N_5447,N_4778,N_3801);
xor U5448 (N_5448,N_532,N_432);
or U5449 (N_5449,N_3983,N_3542);
nor U5450 (N_5450,N_155,N_139);
xor U5451 (N_5451,N_4917,N_874);
or U5452 (N_5452,N_2767,N_607);
xnor U5453 (N_5453,N_3104,N_796);
nor U5454 (N_5454,N_2539,N_832);
xnor U5455 (N_5455,N_3594,N_4806);
nand U5456 (N_5456,N_2584,N_799);
nand U5457 (N_5457,N_4823,N_917);
and U5458 (N_5458,N_2077,N_526);
xnor U5459 (N_5459,N_4164,N_3832);
and U5460 (N_5460,N_464,N_2220);
nor U5461 (N_5461,N_1570,N_71);
nand U5462 (N_5462,N_2192,N_2525);
nand U5463 (N_5463,N_2795,N_4005);
and U5464 (N_5464,N_1984,N_3840);
xnor U5465 (N_5465,N_594,N_3083);
and U5466 (N_5466,N_4100,N_3174);
xor U5467 (N_5467,N_1148,N_2791);
nor U5468 (N_5468,N_3008,N_3989);
or U5469 (N_5469,N_1910,N_4964);
or U5470 (N_5470,N_783,N_1724);
or U5471 (N_5471,N_846,N_4567);
or U5472 (N_5472,N_2661,N_4736);
nor U5473 (N_5473,N_317,N_2063);
xnor U5474 (N_5474,N_1815,N_97);
xnor U5475 (N_5475,N_4571,N_973);
nor U5476 (N_5476,N_2136,N_4849);
and U5477 (N_5477,N_4147,N_1770);
and U5478 (N_5478,N_4622,N_3340);
nor U5479 (N_5479,N_86,N_1270);
or U5480 (N_5480,N_2304,N_133);
nor U5481 (N_5481,N_2478,N_1153);
or U5482 (N_5482,N_280,N_7);
or U5483 (N_5483,N_4256,N_3953);
or U5484 (N_5484,N_248,N_89);
nor U5485 (N_5485,N_3603,N_4741);
or U5486 (N_5486,N_1058,N_3183);
nor U5487 (N_5487,N_3901,N_599);
nand U5488 (N_5488,N_3172,N_4417);
or U5489 (N_5489,N_165,N_2950);
and U5490 (N_5490,N_443,N_710);
nor U5491 (N_5491,N_3553,N_759);
or U5492 (N_5492,N_4816,N_626);
or U5493 (N_5493,N_1564,N_833);
nor U5494 (N_5494,N_2946,N_1989);
xnor U5495 (N_5495,N_909,N_4597);
nand U5496 (N_5496,N_1458,N_4686);
or U5497 (N_5497,N_26,N_2040);
and U5498 (N_5498,N_4130,N_3503);
and U5499 (N_5499,N_3072,N_4797);
and U5500 (N_5500,N_291,N_751);
xor U5501 (N_5501,N_4050,N_361);
nand U5502 (N_5502,N_2649,N_820);
and U5503 (N_5503,N_3477,N_494);
nor U5504 (N_5504,N_1530,N_4165);
or U5505 (N_5505,N_756,N_2349);
or U5506 (N_5506,N_2372,N_2270);
nand U5507 (N_5507,N_2060,N_2920);
or U5508 (N_5508,N_2274,N_910);
nand U5509 (N_5509,N_1674,N_3475);
and U5510 (N_5510,N_4733,N_2365);
and U5511 (N_5511,N_3566,N_1446);
nand U5512 (N_5512,N_3910,N_1027);
or U5513 (N_5513,N_2775,N_2786);
nand U5514 (N_5514,N_4292,N_4743);
or U5515 (N_5515,N_300,N_4451);
nor U5516 (N_5516,N_3731,N_2744);
or U5517 (N_5517,N_3528,N_1889);
xor U5518 (N_5518,N_2141,N_1445);
xnor U5519 (N_5519,N_1857,N_3437);
or U5520 (N_5520,N_3388,N_1574);
xor U5521 (N_5521,N_3527,N_81);
and U5522 (N_5522,N_3794,N_2167);
nor U5523 (N_5523,N_4079,N_1679);
nor U5524 (N_5524,N_68,N_2357);
and U5525 (N_5525,N_1084,N_416);
xor U5526 (N_5526,N_4124,N_1498);
nand U5527 (N_5527,N_2527,N_3287);
and U5528 (N_5528,N_1988,N_905);
or U5529 (N_5529,N_637,N_2718);
or U5530 (N_5530,N_3762,N_2463);
nand U5531 (N_5531,N_3904,N_3391);
nor U5532 (N_5532,N_1809,N_3332);
or U5533 (N_5533,N_1286,N_2738);
and U5534 (N_5534,N_236,N_2160);
nor U5535 (N_5535,N_46,N_3533);
xor U5536 (N_5536,N_2126,N_3205);
xor U5537 (N_5537,N_3091,N_4080);
or U5538 (N_5538,N_1143,N_3257);
or U5539 (N_5539,N_3607,N_2682);
or U5540 (N_5540,N_454,N_476);
nor U5541 (N_5541,N_2659,N_1635);
xor U5542 (N_5542,N_1744,N_2643);
nor U5543 (N_5543,N_2173,N_154);
nor U5544 (N_5544,N_578,N_1111);
or U5545 (N_5545,N_182,N_170);
and U5546 (N_5546,N_4540,N_969);
or U5547 (N_5547,N_2632,N_2389);
nor U5548 (N_5548,N_3235,N_2105);
nor U5549 (N_5549,N_1281,N_4000);
xnor U5550 (N_5550,N_4269,N_1462);
or U5551 (N_5551,N_2260,N_1933);
or U5552 (N_5552,N_1730,N_8);
or U5553 (N_5553,N_2079,N_3310);
nand U5554 (N_5554,N_188,N_3590);
xor U5555 (N_5555,N_2264,N_3191);
or U5556 (N_5556,N_326,N_1482);
and U5557 (N_5557,N_4896,N_4224);
and U5558 (N_5558,N_2161,N_662);
nor U5559 (N_5559,N_1125,N_4082);
nand U5560 (N_5560,N_636,N_4372);
nand U5561 (N_5561,N_3845,N_3373);
nor U5562 (N_5562,N_1619,N_3698);
xnor U5563 (N_5563,N_1408,N_3002);
xnor U5564 (N_5564,N_3396,N_256);
or U5565 (N_5565,N_2498,N_2883);
nor U5566 (N_5566,N_2591,N_972);
and U5567 (N_5567,N_3258,N_749);
and U5568 (N_5568,N_1869,N_3570);
nand U5569 (N_5569,N_3144,N_3079);
and U5570 (N_5570,N_4109,N_641);
or U5571 (N_5571,N_3126,N_1365);
and U5572 (N_5572,N_1922,N_825);
and U5573 (N_5573,N_3756,N_3835);
or U5574 (N_5574,N_577,N_1020);
nor U5575 (N_5575,N_653,N_2501);
nand U5576 (N_5576,N_590,N_2303);
or U5577 (N_5577,N_699,N_1487);
and U5578 (N_5578,N_830,N_4875);
nand U5579 (N_5579,N_1745,N_3336);
or U5580 (N_5580,N_2743,N_41);
nor U5581 (N_5581,N_2889,N_414);
xor U5582 (N_5582,N_1578,N_764);
nor U5583 (N_5583,N_2439,N_4740);
xnor U5584 (N_5584,N_369,N_4520);
or U5585 (N_5585,N_142,N_3851);
nand U5586 (N_5586,N_4138,N_1212);
nand U5587 (N_5587,N_4945,N_2109);
and U5588 (N_5588,N_4759,N_2461);
nand U5589 (N_5589,N_760,N_4771);
xnor U5590 (N_5590,N_1917,N_67);
nand U5591 (N_5591,N_4380,N_2696);
nor U5592 (N_5592,N_3922,N_3111);
nand U5593 (N_5593,N_2886,N_4985);
or U5594 (N_5594,N_4531,N_2861);
xor U5595 (N_5595,N_3274,N_3443);
nand U5596 (N_5596,N_4392,N_3935);
or U5597 (N_5597,N_3577,N_3959);
nand U5598 (N_5598,N_40,N_4583);
nor U5599 (N_5599,N_4881,N_2102);
or U5600 (N_5600,N_3094,N_327);
nand U5601 (N_5601,N_102,N_3157);
xor U5602 (N_5602,N_2803,N_3230);
nand U5603 (N_5603,N_4317,N_1858);
or U5604 (N_5604,N_4286,N_488);
and U5605 (N_5605,N_3395,N_2271);
and U5606 (N_5606,N_676,N_4947);
xnor U5607 (N_5607,N_721,N_3254);
nand U5608 (N_5608,N_1195,N_1292);
or U5609 (N_5609,N_1206,N_1748);
nor U5610 (N_5610,N_1219,N_2118);
xnor U5611 (N_5611,N_1298,N_3550);
nand U5612 (N_5612,N_2875,N_2708);
or U5613 (N_5613,N_1932,N_1871);
nand U5614 (N_5614,N_2965,N_2864);
nand U5615 (N_5615,N_1367,N_3221);
nor U5616 (N_5616,N_1118,N_2415);
nand U5617 (N_5617,N_3694,N_1034);
or U5618 (N_5618,N_162,N_1555);
nor U5619 (N_5619,N_3141,N_4522);
nor U5620 (N_5620,N_1608,N_2693);
nor U5621 (N_5621,N_3447,N_2110);
nand U5622 (N_5622,N_3220,N_4033);
nand U5623 (N_5623,N_4148,N_2156);
nor U5624 (N_5624,N_4873,N_1324);
nor U5625 (N_5625,N_435,N_4559);
and U5626 (N_5626,N_2802,N_4847);
nor U5627 (N_5627,N_4154,N_851);
xor U5628 (N_5628,N_4692,N_255);
or U5629 (N_5629,N_880,N_1723);
nor U5630 (N_5630,N_2766,N_1044);
nor U5631 (N_5631,N_4899,N_4818);
or U5632 (N_5632,N_3877,N_2479);
or U5633 (N_5633,N_4783,N_1773);
nand U5634 (N_5634,N_711,N_87);
nor U5635 (N_5635,N_373,N_1700);
nand U5636 (N_5636,N_1732,N_269);
nor U5637 (N_5637,N_84,N_2053);
and U5638 (N_5638,N_1411,N_4002);
or U5639 (N_5639,N_4334,N_3746);
or U5640 (N_5640,N_587,N_4675);
and U5641 (N_5641,N_3770,N_3211);
and U5642 (N_5642,N_3119,N_2429);
nand U5643 (N_5643,N_4971,N_2404);
xor U5644 (N_5644,N_718,N_4022);
xor U5645 (N_5645,N_1524,N_3309);
xnor U5646 (N_5646,N_634,N_3322);
and U5647 (N_5647,N_2655,N_4157);
nor U5648 (N_5648,N_4303,N_1918);
xor U5649 (N_5649,N_231,N_4199);
nor U5650 (N_5650,N_4838,N_197);
and U5651 (N_5651,N_3635,N_198);
and U5652 (N_5652,N_129,N_955);
nand U5653 (N_5653,N_1254,N_1548);
nand U5654 (N_5654,N_3266,N_304);
nand U5655 (N_5655,N_2533,N_3367);
or U5656 (N_5656,N_2637,N_1565);
nor U5657 (N_5657,N_2371,N_2314);
or U5658 (N_5658,N_337,N_2559);
and U5659 (N_5659,N_1434,N_4499);
nand U5660 (N_5660,N_939,N_4683);
xor U5661 (N_5661,N_2166,N_1897);
or U5662 (N_5662,N_3822,N_223);
nand U5663 (N_5663,N_2504,N_3646);
nand U5664 (N_5664,N_4851,N_4078);
nor U5665 (N_5665,N_452,N_4934);
nand U5666 (N_5666,N_1821,N_2407);
nand U5667 (N_5667,N_1189,N_3084);
xnor U5668 (N_5668,N_1962,N_385);
nor U5669 (N_5669,N_3888,N_4337);
xor U5670 (N_5670,N_4071,N_1262);
or U5671 (N_5671,N_3037,N_3860);
xnor U5672 (N_5672,N_679,N_1640);
and U5673 (N_5673,N_405,N_1257);
or U5674 (N_5674,N_3732,N_1211);
or U5675 (N_5675,N_3508,N_4764);
or U5676 (N_5676,N_4158,N_4297);
or U5677 (N_5677,N_4668,N_3625);
nor U5678 (N_5678,N_4273,N_3142);
nor U5679 (N_5679,N_53,N_4758);
nor U5680 (N_5680,N_3182,N_3244);
and U5681 (N_5681,N_3783,N_3232);
nor U5682 (N_5682,N_954,N_316);
nor U5683 (N_5683,N_4122,N_3815);
or U5684 (N_5684,N_2387,N_1721);
nand U5685 (N_5685,N_406,N_1107);
or U5686 (N_5686,N_2368,N_2893);
xor U5687 (N_5687,N_2989,N_4362);
or U5688 (N_5688,N_2804,N_4791);
xnor U5689 (N_5689,N_4852,N_4135);
nand U5690 (N_5690,N_1643,N_1345);
nor U5691 (N_5691,N_2968,N_2927);
nor U5692 (N_5692,N_3372,N_3942);
nand U5693 (N_5693,N_2360,N_3486);
nand U5694 (N_5694,N_1957,N_3308);
nand U5695 (N_5695,N_262,N_4993);
and U5696 (N_5696,N_323,N_4272);
or U5697 (N_5697,N_3370,N_507);
xor U5698 (N_5698,N_1970,N_2388);
and U5699 (N_5699,N_2851,N_2280);
nor U5700 (N_5700,N_137,N_64);
or U5701 (N_5701,N_920,N_761);
nand U5702 (N_5702,N_4903,N_4257);
or U5703 (N_5703,N_3357,N_1062);
xnor U5704 (N_5704,N_4591,N_1438);
xnor U5705 (N_5705,N_4173,N_377);
or U5706 (N_5706,N_1552,N_1480);
nand U5707 (N_5707,N_203,N_1502);
xor U5708 (N_5708,N_1142,N_674);
or U5709 (N_5709,N_616,N_4637);
or U5710 (N_5710,N_992,N_2057);
and U5711 (N_5711,N_353,N_357);
or U5712 (N_5712,N_4261,N_2296);
and U5713 (N_5713,N_4194,N_3642);
and U5714 (N_5714,N_1611,N_4871);
xnor U5715 (N_5715,N_3439,N_1491);
xnor U5716 (N_5716,N_3341,N_27);
nand U5717 (N_5717,N_3321,N_4861);
xnor U5718 (N_5718,N_2945,N_74);
nand U5719 (N_5719,N_272,N_2971);
xnor U5720 (N_5720,N_461,N_3777);
xor U5721 (N_5721,N_4643,N_2624);
nand U5722 (N_5722,N_4663,N_1453);
nand U5723 (N_5723,N_2568,N_2798);
nand U5724 (N_5724,N_2178,N_1843);
nand U5725 (N_5725,N_1672,N_2408);
xnor U5726 (N_5726,N_3516,N_4606);
nand U5727 (N_5727,N_4543,N_1776);
and U5728 (N_5728,N_937,N_3325);
and U5729 (N_5729,N_400,N_3792);
and U5730 (N_5730,N_4289,N_4629);
xor U5731 (N_5731,N_1980,N_4409);
xor U5732 (N_5732,N_2297,N_3282);
xor U5733 (N_5733,N_3562,N_1911);
or U5734 (N_5734,N_30,N_2261);
nor U5735 (N_5735,N_4982,N_1091);
or U5736 (N_5736,N_2916,N_1999);
or U5737 (N_5737,N_1650,N_2810);
nand U5738 (N_5738,N_810,N_3490);
nand U5739 (N_5739,N_372,N_3468);
nand U5740 (N_5740,N_4101,N_503);
nor U5741 (N_5741,N_758,N_1777);
xor U5742 (N_5742,N_4908,N_4107);
nor U5743 (N_5743,N_4919,N_4943);
or U5744 (N_5744,N_2064,N_1339);
xnor U5745 (N_5745,N_2941,N_925);
xor U5746 (N_5746,N_249,N_727);
nor U5747 (N_5747,N_1326,N_3300);
nand U5748 (N_5748,N_2520,N_1913);
xor U5749 (N_5749,N_2951,N_1948);
nand U5750 (N_5750,N_1244,N_2301);
xnor U5751 (N_5751,N_3628,N_1532);
nand U5752 (N_5752,N_3134,N_2705);
and U5753 (N_5753,N_1824,N_3800);
nor U5754 (N_5754,N_2565,N_3048);
nand U5755 (N_5755,N_3591,N_1924);
or U5756 (N_5756,N_1862,N_2034);
nand U5757 (N_5757,N_1005,N_948);
nor U5758 (N_5758,N_2716,N_3033);
and U5759 (N_5759,N_648,N_1023);
or U5760 (N_5760,N_998,N_3197);
nand U5761 (N_5761,N_257,N_4325);
nand U5762 (N_5762,N_4718,N_1201);
xnor U5763 (N_5763,N_2252,N_4836);
or U5764 (N_5764,N_3151,N_2273);
and U5765 (N_5765,N_3267,N_1609);
or U5766 (N_5766,N_1246,N_1140);
nand U5767 (N_5767,N_3748,N_2730);
and U5768 (N_5768,N_2913,N_4704);
nand U5769 (N_5769,N_252,N_2914);
nor U5770 (N_5770,N_4070,N_1204);
and U5771 (N_5771,N_3557,N_3825);
nand U5772 (N_5772,N_4785,N_2973);
and U5773 (N_5773,N_3358,N_1022);
xnor U5774 (N_5774,N_3896,N_2369);
nor U5775 (N_5775,N_3303,N_1000);
and U5776 (N_5776,N_525,N_2468);
or U5777 (N_5777,N_1873,N_3610);
and U5778 (N_5778,N_2666,N_1765);
nand U5779 (N_5779,N_1515,N_250);
and U5780 (N_5780,N_1505,N_2955);
xnor U5781 (N_5781,N_979,N_1275);
or U5782 (N_5782,N_3056,N_613);
and U5783 (N_5783,N_932,N_3241);
nand U5784 (N_5784,N_3811,N_352);
or U5785 (N_5785,N_2390,N_398);
nand U5786 (N_5786,N_2751,N_3727);
nor U5787 (N_5787,N_3633,N_1556);
and U5788 (N_5788,N_771,N_4333);
nand U5789 (N_5789,N_1559,N_2330);
and U5790 (N_5790,N_2181,N_890);
xnor U5791 (N_5791,N_1343,N_3638);
or U5792 (N_5792,N_2222,N_312);
or U5793 (N_5793,N_4593,N_1633);
and U5794 (N_5794,N_663,N_3510);
xnor U5795 (N_5795,N_4979,N_4346);
nor U5796 (N_5796,N_3507,N_3782);
xor U5797 (N_5797,N_4782,N_2437);
or U5798 (N_5798,N_4035,N_2011);
xnor U5799 (N_5799,N_2787,N_2862);
xnor U5800 (N_5800,N_3077,N_3719);
nand U5801 (N_5801,N_3865,N_4983);
or U5802 (N_5802,N_1692,N_2176);
nor U5803 (N_5803,N_4719,N_3675);
or U5804 (N_5804,N_3747,N_3101);
nor U5805 (N_5805,N_1666,N_3463);
and U5806 (N_5806,N_2028,N_580);
nand U5807 (N_5807,N_745,N_222);
or U5808 (N_5808,N_649,N_4161);
or U5809 (N_5809,N_3005,N_1268);
xor U5810 (N_5810,N_4569,N_4900);
and U5811 (N_5811,N_863,N_1925);
or U5812 (N_5812,N_456,N_1580);
xnor U5813 (N_5813,N_978,N_1347);
xor U5814 (N_5814,N_3166,N_995);
nor U5815 (N_5815,N_1247,N_1470);
xor U5816 (N_5816,N_4616,N_164);
nor U5817 (N_5817,N_3161,N_4518);
xnor U5818 (N_5818,N_3047,N_4389);
nor U5819 (N_5819,N_4601,N_4162);
or U5820 (N_5820,N_1725,N_1787);
or U5821 (N_5821,N_4430,N_4367);
or U5822 (N_5822,N_421,N_3780);
and U5823 (N_5823,N_187,N_4075);
nand U5824 (N_5824,N_1304,N_2752);
nand U5825 (N_5825,N_1959,N_1463);
nand U5826 (N_5826,N_4471,N_2185);
xnor U5827 (N_5827,N_1130,N_4536);
xor U5828 (N_5828,N_290,N_105);
nor U5829 (N_5829,N_2444,N_1414);
nor U5830 (N_5830,N_195,N_4314);
nor U5831 (N_5831,N_3691,N_2442);
xnor U5832 (N_5832,N_2779,N_2038);
xor U5833 (N_5833,N_2827,N_823);
nor U5834 (N_5834,N_2635,N_4807);
or U5835 (N_5835,N_180,N_3194);
nor U5836 (N_5836,N_194,N_1442);
nand U5837 (N_5837,N_1842,N_2781);
or U5838 (N_5838,N_2515,N_3561);
nand U5839 (N_5839,N_3689,N_873);
xor U5840 (N_5840,N_798,N_1209);
xor U5841 (N_5841,N_2922,N_408);
nand U5842 (N_5842,N_78,N_4987);
nand U5843 (N_5843,N_3135,N_2239);
xor U5844 (N_5844,N_463,N_128);
xor U5845 (N_5845,N_901,N_4229);
nand U5846 (N_5846,N_2423,N_2114);
xnor U5847 (N_5847,N_3127,N_3871);
or U5848 (N_5848,N_4046,N_277);
nand U5849 (N_5849,N_1081,N_1517);
or U5850 (N_5850,N_396,N_1812);
nand U5851 (N_5851,N_2522,N_3295);
xor U5852 (N_5852,N_234,N_2753);
or U5853 (N_5853,N_9,N_2143);
or U5854 (N_5854,N_1124,N_1676);
nor U5855 (N_5855,N_224,N_986);
nand U5856 (N_5856,N_3964,N_499);
or U5857 (N_5857,N_3788,N_3778);
nor U5858 (N_5858,N_2029,N_1278);
nor U5859 (N_5859,N_869,N_1908);
nor U5860 (N_5860,N_486,N_878);
nand U5861 (N_5861,N_1553,N_1920);
and U5862 (N_5862,N_3416,N_1173);
or U5863 (N_5863,N_3911,N_1287);
xnor U5864 (N_5864,N_2027,N_2972);
nor U5865 (N_5865,N_259,N_976);
nand U5866 (N_5866,N_29,N_4548);
nand U5867 (N_5867,N_4946,N_3096);
nor U5868 (N_5868,N_4152,N_1085);
nand U5869 (N_5869,N_3866,N_1567);
nor U5870 (N_5870,N_174,N_1644);
and U5871 (N_5871,N_934,N_3987);
or U5872 (N_5872,N_1818,N_4106);
or U5873 (N_5873,N_2356,N_4516);
nand U5874 (N_5874,N_2957,N_3848);
nor U5875 (N_5875,N_2995,N_923);
xnor U5876 (N_5876,N_2380,N_3488);
nor U5877 (N_5877,N_3253,N_3281);
xor U5878 (N_5878,N_3092,N_2799);
and U5879 (N_5879,N_4697,N_1050);
or U5880 (N_5880,N_482,N_245);
xor U5881 (N_5881,N_4413,N_1351);
or U5882 (N_5882,N_1348,N_1937);
or U5883 (N_5883,N_1793,N_3360);
xnor U5884 (N_5884,N_462,N_3497);
nand U5885 (N_5885,N_635,N_4815);
or U5886 (N_5886,N_849,N_1405);
xor U5887 (N_5887,N_88,N_2146);
or U5888 (N_5888,N_2012,N_3286);
or U5889 (N_5889,N_3741,N_3494);
and U5890 (N_5890,N_2062,N_3806);
nand U5891 (N_5891,N_2489,N_2981);
xnor U5892 (N_5892,N_2747,N_1052);
and U5893 (N_5893,N_3417,N_2606);
nand U5894 (N_5894,N_3479,N_1572);
nor U5895 (N_5895,N_3611,N_1313);
and U5896 (N_5896,N_3409,N_4212);
nand U5897 (N_5897,N_4933,N_693);
nand U5898 (N_5898,N_3496,N_2644);
and U5899 (N_5899,N_2424,N_1053);
nor U5900 (N_5900,N_4477,N_1366);
and U5901 (N_5901,N_4203,N_517);
xnor U5902 (N_5902,N_3017,N_2812);
or U5903 (N_5903,N_2367,N_1835);
and U5904 (N_5904,N_779,N_3271);
xnor U5905 (N_5905,N_1008,N_1509);
nor U5906 (N_5906,N_1872,N_3376);
or U5907 (N_5907,N_4748,N_3915);
or U5908 (N_5908,N_1690,N_3399);
nor U5909 (N_5909,N_2966,N_3869);
nand U5910 (N_5910,N_1215,N_3299);
nand U5911 (N_5911,N_514,N_1896);
xnor U5912 (N_5912,N_4209,N_3378);
xnor U5913 (N_5913,N_647,N_2538);
or U5914 (N_5914,N_4960,N_3842);
nand U5915 (N_5915,N_3721,N_706);
and U5916 (N_5916,N_4368,N_4822);
or U5917 (N_5917,N_2619,N_2727);
and U5918 (N_5918,N_1840,N_3167);
xor U5919 (N_5919,N_776,N_2823);
or U5920 (N_5920,N_777,N_1075);
and U5921 (N_5921,N_4562,N_4776);
and U5922 (N_5922,N_4940,N_143);
xnor U5923 (N_5923,N_2888,N_2980);
or U5924 (N_5924,N_3273,N_285);
nand U5925 (N_5925,N_3656,N_1252);
xor U5926 (N_5926,N_795,N_4721);
nor U5927 (N_5927,N_3240,N_3582);
xnor U5928 (N_5928,N_1363,N_190);
or U5929 (N_5929,N_1540,N_4603);
xnor U5930 (N_5930,N_1393,N_3545);
nand U5931 (N_5931,N_301,N_2725);
nand U5932 (N_5932,N_2379,N_2226);
nor U5933 (N_5933,N_1597,N_209);
and U5934 (N_5934,N_4796,N_2943);
or U5935 (N_5935,N_2282,N_4619);
xor U5936 (N_5936,N_4385,N_3715);
xor U5937 (N_5937,N_3246,N_3028);
or U5938 (N_5938,N_3580,N_530);
and U5939 (N_5939,N_4928,N_3296);
or U5940 (N_5940,N_585,N_4185);
nor U5941 (N_5941,N_363,N_652);
or U5942 (N_5942,N_1496,N_2749);
or U5943 (N_5943,N_473,N_3938);
or U5944 (N_5944,N_1120,N_4654);
or U5945 (N_5945,N_340,N_659);
or U5946 (N_5946,N_2289,N_1241);
xor U5947 (N_5947,N_4794,N_716);
nor U5948 (N_5948,N_2821,N_3604);
or U5949 (N_5949,N_3546,N_3957);
xnor U5950 (N_5950,N_1575,N_3154);
nand U5951 (N_5951,N_853,N_4155);
and U5952 (N_5952,N_1041,N_3828);
or U5953 (N_5953,N_936,N_3583);
and U5954 (N_5954,N_4980,N_3361);
and U5955 (N_5955,N_3916,N_4340);
or U5956 (N_5956,N_2542,N_3823);
and U5957 (N_5957,N_2701,N_1145);
xnor U5958 (N_5958,N_242,N_2928);
and U5959 (N_5959,N_2431,N_1168);
or U5960 (N_5960,N_1169,N_3597);
and U5961 (N_5961,N_1891,N_3764);
xnor U5962 (N_5962,N_4128,N_1866);
nand U5963 (N_5963,N_3651,N_2518);
nand U5964 (N_5964,N_1653,N_1967);
nand U5965 (N_5965,N_4792,N_881);
and U5966 (N_5966,N_4765,N_1251);
nor U5967 (N_5967,N_2100,N_1456);
or U5968 (N_5968,N_3445,N_2069);
and U5969 (N_5969,N_1909,N_1234);
xor U5970 (N_5970,N_2432,N_4798);
nand U5971 (N_5971,N_3198,N_4492);
or U5972 (N_5972,N_1001,N_339);
and U5973 (N_5973,N_2179,N_1432);
nand U5974 (N_5974,N_2599,N_2541);
and U5975 (N_5975,N_583,N_2760);
nor U5976 (N_5976,N_2310,N_4090);
and U5977 (N_5977,N_4353,N_2394);
nor U5978 (N_5978,N_935,N_214);
nand U5979 (N_5979,N_1299,N_2174);
or U5980 (N_5980,N_4527,N_709);
nor U5981 (N_5981,N_3520,N_1887);
nor U5982 (N_5982,N_3402,N_4077);
nand U5983 (N_5983,N_1954,N_3059);
or U5984 (N_5984,N_4927,N_2334);
and U5985 (N_5985,N_450,N_3121);
nor U5986 (N_5986,N_2736,N_4309);
or U5987 (N_5987,N_2313,N_3316);
nor U5988 (N_5988,N_2872,N_1881);
xnor U5989 (N_5989,N_2919,N_2088);
and U5990 (N_5990,N_1248,N_2370);
nand U5991 (N_5991,N_2084,N_115);
xnor U5992 (N_5992,N_382,N_805);
and U5993 (N_5993,N_3990,N_3585);
and U5994 (N_5994,N_2419,N_4870);
nor U5995 (N_5995,N_2051,N_3665);
nor U5996 (N_5996,N_3599,N_814);
xnor U5997 (N_5997,N_172,N_2516);
nor U5998 (N_5998,N_2039,N_2780);
nor U5999 (N_5999,N_403,N_4245);
and U6000 (N_6000,N_690,N_1722);
nand U6001 (N_6001,N_3979,N_227);
or U6002 (N_6002,N_2347,N_2083);
and U6003 (N_6003,N_3070,N_1492);
or U6004 (N_6004,N_984,N_258);
xor U6005 (N_6005,N_150,N_4777);
nor U6006 (N_6006,N_672,N_2969);
nor U6007 (N_6007,N_485,N_4267);
and U6008 (N_6008,N_3837,N_3998);
or U6009 (N_6009,N_2609,N_4617);
nand U6010 (N_6010,N_829,N_1267);
or U6011 (N_6011,N_4393,N_1651);
nor U6012 (N_6012,N_519,N_2555);
or U6013 (N_6013,N_1588,N_2414);
xor U6014 (N_6014,N_1344,N_1359);
or U6015 (N_6015,N_1655,N_3392);
and U6016 (N_6016,N_4862,N_2572);
nand U6017 (N_6017,N_1952,N_4448);
xor U6018 (N_6018,N_4604,N_1756);
or U6019 (N_6019,N_1419,N_466);
nand U6020 (N_6020,N_4151,N_4004);
or U6021 (N_6021,N_2677,N_2853);
nand U6022 (N_6022,N_3994,N_1447);
xnor U6023 (N_6023,N_2398,N_2552);
and U6024 (N_6024,N_4495,N_1271);
xor U6025 (N_6025,N_4324,N_348);
and U6026 (N_6026,N_265,N_2248);
and U6027 (N_6027,N_207,N_2800);
nor U6028 (N_6028,N_926,N_4988);
or U6029 (N_6029,N_4012,N_608);
nand U6030 (N_6030,N_4805,N_915);
and U6031 (N_6031,N_2202,N_2484);
and U6032 (N_6032,N_4264,N_336);
nor U6033 (N_6033,N_3618,N_2709);
and U6034 (N_6034,N_199,N_908);
and U6035 (N_6035,N_1936,N_3148);
nor U6036 (N_6036,N_4786,N_1051);
xnor U6037 (N_6037,N_2745,N_4705);
xnor U6038 (N_6038,N_1894,N_2952);
nand U6039 (N_6039,N_4652,N_3331);
nand U6040 (N_6040,N_410,N_2309);
or U6041 (N_6041,N_3255,N_3519);
xor U6042 (N_6042,N_1092,N_3889);
nor U6043 (N_6043,N_2508,N_1698);
xnor U6044 (N_6044,N_1028,N_512);
nand U6045 (N_6045,N_3066,N_552);
xor U6046 (N_6046,N_918,N_1449);
or U6047 (N_6047,N_358,N_3106);
or U6048 (N_6048,N_2004,N_3049);
nor U6049 (N_6049,N_1207,N_3637);
or U6050 (N_6050,N_3870,N_4700);
and U6051 (N_6051,N_1335,N_235);
nand U6052 (N_6052,N_1380,N_3682);
and U6053 (N_6053,N_2721,N_2237);
and U6054 (N_6054,N_3250,N_360);
nor U6055 (N_6055,N_28,N_3639);
and U6056 (N_6056,N_2921,N_736);
or U6057 (N_6057,N_3259,N_2393);
nand U6058 (N_6058,N_1766,N_4276);
nor U6059 (N_6059,N_4999,N_3415);
or U6060 (N_6060,N_4551,N_559);
or U6061 (N_6061,N_469,N_1855);
or U6062 (N_6062,N_2003,N_3829);
or U6063 (N_6063,N_297,N_2486);
nand U6064 (N_6064,N_1753,N_747);
nor U6065 (N_6065,N_1714,N_1078);
xor U6066 (N_6066,N_2648,N_1198);
nand U6067 (N_6067,N_3064,N_505);
nor U6068 (N_6068,N_2750,N_4766);
nand U6069 (N_6069,N_1541,N_944);
and U6070 (N_6070,N_2850,N_573);
or U6071 (N_6071,N_4131,N_1794);
nor U6072 (N_6072,N_3734,N_3543);
nor U6073 (N_6073,N_3128,N_3787);
or U6074 (N_6074,N_3485,N_455);
nand U6075 (N_6075,N_4027,N_3329);
and U6076 (N_6076,N_3237,N_1823);
nor U6077 (N_6077,N_1639,N_3818);
nand U6078 (N_6078,N_3380,N_1783);
nor U6079 (N_6079,N_4832,N_3305);
xor U6080 (N_6080,N_4054,N_4378);
xnor U6081 (N_6081,N_2704,N_1220);
nand U6082 (N_6082,N_4478,N_824);
nand U6083 (N_6083,N_3988,N_4420);
and U6084 (N_6084,N_2250,N_4488);
xnor U6085 (N_6085,N_430,N_1537);
xnor U6086 (N_6086,N_2550,N_2048);
xnor U6087 (N_6087,N_668,N_3041);
xnor U6088 (N_6088,N_3624,N_431);
or U6089 (N_6089,N_15,N_4307);
or U6090 (N_6090,N_1425,N_2094);
and U6091 (N_6091,N_4313,N_1017);
nor U6092 (N_6092,N_4319,N_1761);
or U6093 (N_6093,N_715,N_2140);
and U6094 (N_6094,N_3140,N_1972);
and U6095 (N_6095,N_3575,N_3937);
nand U6096 (N_6096,N_3348,N_2519);
nor U6097 (N_6097,N_1737,N_2251);
nand U6098 (N_6098,N_2587,N_2024);
and U6099 (N_6099,N_3199,N_3986);
or U6100 (N_6100,N_4403,N_1139);
nand U6101 (N_6101,N_76,N_4720);
xnor U6102 (N_6102,N_509,N_263);
xnor U6103 (N_6103,N_1242,N_4013);
nor U6104 (N_6104,N_1978,N_3192);
or U6105 (N_6105,N_4301,N_3462);
nor U6106 (N_6106,N_4770,N_3419);
xnor U6107 (N_6107,N_1094,N_513);
xor U6108 (N_6108,N_3384,N_2694);
nand U6109 (N_6109,N_3887,N_733);
xnor U6110 (N_6110,N_4994,N_4661);
xnor U6111 (N_6111,N_1784,N_2528);
xnor U6112 (N_6112,N_3302,N_3426);
xor U6113 (N_6113,N_4772,N_4316);
xnor U6114 (N_6114,N_1563,N_2832);
xnor U6115 (N_6115,N_3576,N_4802);
or U6116 (N_6116,N_3578,N_3600);
nor U6117 (N_6117,N_3324,N_4693);
nor U6118 (N_6118,N_2348,N_1620);
nor U6119 (N_6119,N_4938,N_2944);
xor U6120 (N_6120,N_2507,N_3785);
nand U6121 (N_6121,N_598,N_4098);
and U6122 (N_6122,N_3652,N_4882);
and U6123 (N_6123,N_2536,N_1088);
or U6124 (N_6124,N_4750,N_3265);
or U6125 (N_6125,N_1990,N_859);
or U6126 (N_6126,N_2413,N_2288);
and U6127 (N_6127,N_4833,N_2580);
nand U6128 (N_6128,N_2482,N_4136);
xor U6129 (N_6129,N_3143,N_3118);
or U6130 (N_6130,N_4026,N_4967);
xor U6131 (N_6131,N_4757,N_2216);
and U6132 (N_6132,N_4037,N_3701);
or U6133 (N_6133,N_3342,N_4284);
xnor U6134 (N_6134,N_4656,N_1739);
nand U6135 (N_6135,N_2152,N_2841);
nand U6136 (N_6136,N_4895,N_4081);
nor U6137 (N_6137,N_2182,N_842);
and U6138 (N_6138,N_719,N_4174);
xnor U6139 (N_6139,N_1033,N_1159);
nand U6140 (N_6140,N_1628,N_1488);
nor U6141 (N_6141,N_57,N_2175);
nor U6142 (N_6142,N_834,N_907);
nor U6143 (N_6143,N_4626,N_4554);
nor U6144 (N_6144,N_2720,N_2556);
xor U6145 (N_6145,N_3880,N_4561);
and U6146 (N_6146,N_4793,N_4444);
and U6147 (N_6147,N_3025,N_1658);
nand U6148 (N_6148,N_276,N_2462);
nand U6149 (N_6149,N_2517,N_1478);
nand U6150 (N_6150,N_4768,N_2050);
and U6151 (N_6151,N_3130,N_1311);
xor U6152 (N_6152,N_2796,N_2692);
or U6153 (N_6153,N_2343,N_4731);
nand U6154 (N_6154,N_3999,N_3030);
nor U6155 (N_6155,N_1087,N_3602);
nor U6156 (N_6156,N_3804,N_2108);
and U6157 (N_6157,N_1595,N_3524);
xor U6158 (N_6158,N_1832,N_1342);
or U6159 (N_6159,N_1637,N_2904);
nand U6160 (N_6160,N_1338,N_1992);
nand U6161 (N_6161,N_970,N_4408);
xnor U6162 (N_6162,N_3853,N_94);
and U6163 (N_6163,N_2361,N_2867);
and U6164 (N_6164,N_797,N_1331);
nor U6165 (N_6165,N_940,N_3264);
or U6166 (N_6166,N_4422,N_459);
xor U6167 (N_6167,N_2191,N_4615);
or U6168 (N_6168,N_2195,N_6);
xnor U6169 (N_6169,N_2933,N_3381);
nor U6170 (N_6170,N_2842,N_3152);
nand U6171 (N_6171,N_4202,N_4991);
nor U6172 (N_6172,N_4371,N_1554);
xor U6173 (N_6173,N_4948,N_1314);
and U6174 (N_6174,N_173,N_1056);
or U6175 (N_6175,N_4874,N_2131);
nand U6176 (N_6176,N_1013,N_595);
or U6177 (N_6177,N_3156,N_2607);
or U6178 (N_6178,N_4623,N_1877);
nor U6179 (N_6179,N_1610,N_556);
or U6180 (N_6180,N_741,N_2269);
nand U6181 (N_6181,N_809,N_2203);
nor U6182 (N_6182,N_4446,N_2982);
nor U6183 (N_6183,N_4715,N_1792);
nand U6184 (N_6184,N_3429,N_1378);
nand U6185 (N_6185,N_424,N_1307);
nand U6186 (N_6186,N_1632,N_835);
and U6187 (N_6187,N_579,N_2460);
or U6188 (N_6188,N_1975,N_1323);
or U6189 (N_6189,N_4992,N_4801);
xor U6190 (N_6190,N_1011,N_11);
and U6191 (N_6191,N_3996,N_1228);
nor U6192 (N_6192,N_2092,N_2198);
nand U6193 (N_6193,N_4464,N_4714);
xnor U6194 (N_6194,N_3408,N_4877);
or U6195 (N_6195,N_889,N_4572);
or U6196 (N_6196,N_1061,N_1325);
xor U6197 (N_6197,N_3125,N_4821);
or U6198 (N_6198,N_960,N_4474);
nand U6199 (N_6199,N_213,N_1368);
nor U6200 (N_6200,N_1394,N_2395);
nand U6201 (N_6201,N_1024,N_3180);
nand U6202 (N_6202,N_3927,N_2090);
nor U6203 (N_6203,N_3902,N_119);
and U6204 (N_6204,N_2474,N_1137);
and U6205 (N_6205,N_3857,N_4647);
xor U6206 (N_6206,N_1971,N_3374);
and U6207 (N_6207,N_2325,N_3262);
xor U6208 (N_6208,N_4804,N_4379);
nand U6209 (N_6209,N_1785,N_2588);
nor U6210 (N_6210,N_2604,N_3364);
xor U6211 (N_6211,N_1836,N_1510);
and U6212 (N_6212,N_2406,N_566);
and U6213 (N_6213,N_3404,N_2085);
or U6214 (N_6214,N_1799,N_790);
nor U6215 (N_6215,N_3744,N_4950);
and U6216 (N_6216,N_2576,N_537);
or U6217 (N_6217,N_95,N_2740);
nor U6218 (N_6218,N_171,N_4912);
or U6219 (N_6219,N_2808,N_3085);
or U6220 (N_6220,N_1002,N_497);
nand U6221 (N_6221,N_1385,N_2493);
and U6222 (N_6222,N_855,N_1003);
xnor U6223 (N_6223,N_1093,N_3584);
nor U6224 (N_6224,N_332,N_2352);
and U6225 (N_6225,N_847,N_4278);
nor U6226 (N_6226,N_2629,N_3109);
or U6227 (N_6227,N_253,N_765);
nor U6228 (N_6228,N_1518,N_4088);
xor U6229 (N_6229,N_930,N_938);
or U6230 (N_6230,N_1115,N_3834);
and U6231 (N_6231,N_23,N_3671);
nor U6232 (N_6232,N_4529,N_3252);
and U6233 (N_6233,N_2549,N_1618);
and U6234 (N_6234,N_757,N_687);
and U6235 (N_6235,N_4086,N_4553);
nor U6236 (N_6236,N_4338,N_1719);
nor U6237 (N_6237,N_1321,N_1850);
or U6238 (N_6238,N_132,N_3436);
xnor U6239 (N_6239,N_1500,N_837);
or U6240 (N_6240,N_3225,N_2267);
nand U6241 (N_6241,N_1329,N_2612);
nor U6242 (N_6242,N_3040,N_3238);
or U6243 (N_6243,N_445,N_1720);
xnor U6244 (N_6244,N_4576,N_3242);
nand U6245 (N_6245,N_1899,N_4924);
and U6246 (N_6246,N_2031,N_3596);
nor U6247 (N_6247,N_3903,N_1230);
nand U6248 (N_6248,N_3058,N_1494);
xor U6249 (N_6249,N_959,N_2892);
xor U6250 (N_6250,N_2774,N_4211);
nand U6251 (N_6251,N_3514,N_2044);
nor U6252 (N_6252,N_1080,N_3046);
xor U6253 (N_6253,N_3891,N_893);
nand U6254 (N_6254,N_4419,N_1749);
nor U6255 (N_6255,N_3452,N_3024);
nor U6256 (N_6256,N_3844,N_3961);
or U6257 (N_6257,N_3695,N_4144);
and U6258 (N_6258,N_540,N_4747);
and U6259 (N_6259,N_546,N_3859);
nor U6260 (N_6260,N_3319,N_4703);
xnor U6261 (N_6261,N_14,N_1615);
xnor U6262 (N_6262,N_2125,N_4756);
nand U6263 (N_6263,N_3958,N_3858);
xor U6264 (N_6264,N_1834,N_884);
nand U6265 (N_6265,N_1334,N_3767);
nor U6266 (N_6266,N_1352,N_4737);
and U6267 (N_6267,N_4898,N_2490);
or U6268 (N_6268,N_1805,N_763);
nor U6269 (N_6269,N_2448,N_2);
nand U6270 (N_6270,N_3444,N_3483);
nor U6271 (N_6271,N_449,N_3297);
xnor U6272 (N_6272,N_299,N_2353);
xor U6273 (N_6273,N_496,N_2469);
and U6274 (N_6274,N_4407,N_3574);
nand U6275 (N_6275,N_1659,N_1584);
and U6276 (N_6276,N_4424,N_2328);
nand U6277 (N_6277,N_1711,N_2446);
or U6278 (N_6278,N_4365,N_3493);
and U6279 (N_6279,N_1669,N_991);
nand U6280 (N_6280,N_4384,N_2600);
nor U6281 (N_6281,N_2543,N_840);
nor U6282 (N_6282,N_4698,N_3766);
nand U6283 (N_6283,N_1059,N_4398);
nor U6284 (N_6284,N_911,N_2396);
and U6285 (N_6285,N_4734,N_1122);
nand U6286 (N_6286,N_3029,N_334);
and U6287 (N_6287,N_3688,N_338);
and U6288 (N_6288,N_1551,N_2976);
nor U6289 (N_6289,N_3045,N_3729);
xnor U6290 (N_6290,N_3330,N_1833);
nand U6291 (N_6291,N_688,N_59);
nor U6292 (N_6292,N_660,N_4453);
nand U6293 (N_6293,N_3648,N_1183);
xor U6294 (N_6294,N_1859,N_4820);
xor U6295 (N_6295,N_3884,N_2586);
or U6296 (N_6296,N_2509,N_4139);
and U6297 (N_6297,N_3413,N_4582);
nand U6298 (N_6298,N_2155,N_1340);
or U6299 (N_6299,N_2523,N_2477);
or U6300 (N_6300,N_4323,N_852);
nand U6301 (N_6301,N_4645,N_3458);
and U6302 (N_6302,N_856,N_4206);
nor U6303 (N_6303,N_962,N_4829);
nor U6304 (N_6304,N_2954,N_4352);
nor U6305 (N_6305,N_3831,N_1612);
or U6306 (N_6306,N_4650,N_983);
xor U6307 (N_6307,N_1860,N_3217);
or U6308 (N_6308,N_4404,N_225);
or U6309 (N_6309,N_714,N_2046);
xnor U6310 (N_6310,N_1596,N_4509);
xnor U6311 (N_6311,N_558,N_2617);
xor U6312 (N_6312,N_4003,N_3662);
and U6313 (N_6313,N_1573,N_3572);
or U6314 (N_6314,N_4610,N_333);
nor U6315 (N_6315,N_4200,N_2530);
and U6316 (N_6316,N_2451,N_3769);
nand U6317 (N_6317,N_1803,N_4570);
nor U6318 (N_6318,N_4607,N_202);
nor U6319 (N_6319,N_2856,N_2190);
xor U6320 (N_6320,N_2932,N_2107);
xnor U6321 (N_6321,N_4843,N_2650);
or U6322 (N_6322,N_4996,N_572);
or U6323 (N_6323,N_1185,N_43);
nand U6324 (N_6324,N_4613,N_3386);
xor U6325 (N_6325,N_3939,N_2689);
and U6326 (N_6326,N_4496,N_4789);
nand U6327 (N_6327,N_4585,N_664);
nor U6328 (N_6328,N_576,N_2362);
and U6329 (N_6329,N_896,N_3312);
xor U6330 (N_6330,N_3228,N_4944);
nor U6331 (N_6331,N_4657,N_772);
xnor U6332 (N_6332,N_1021,N_2626);
xor U6333 (N_6333,N_3549,N_708);
nand U6334 (N_6334,N_3864,N_4784);
xor U6335 (N_6335,N_956,N_2735);
and U6336 (N_6336,N_2734,N_2514);
or U6337 (N_6337,N_681,N_642);
xor U6338 (N_6338,N_4119,N_1848);
nor U6339 (N_6339,N_2345,N_4099);
nand U6340 (N_6340,N_1009,N_72);
nand U6341 (N_6341,N_4219,N_2712);
xor U6342 (N_6342,N_117,N_4062);
or U6343 (N_6343,N_800,N_1600);
or U6344 (N_6344,N_3521,N_1116);
or U6345 (N_6345,N_1160,N_1121);
and U6346 (N_6346,N_1516,N_2715);
nor U6347 (N_6347,N_4382,N_4391);
nor U6348 (N_6348,N_4028,N_4118);
nand U6349 (N_6349,N_3019,N_4621);
xor U6350 (N_6350,N_1807,N_1012);
and U6351 (N_6351,N_697,N_3013);
nor U6352 (N_6352,N_3171,N_3326);
or U6353 (N_6353,N_2258,N_1513);
nor U6354 (N_6354,N_2227,N_1906);
or U6355 (N_6355,N_879,N_3740);
xnor U6356 (N_6356,N_2547,N_1533);
or U6357 (N_6357,N_4247,N_2421);
nor U6358 (N_6358,N_320,N_80);
nand U6359 (N_6359,N_2433,N_4620);
nor U6360 (N_6360,N_2761,N_2278);
nor U6361 (N_6361,N_4233,N_588);
nand U6362 (N_6362,N_605,N_3108);
or U6363 (N_6363,N_815,N_623);
and U6364 (N_6364,N_4505,N_2217);
xor U6365 (N_6365,N_3981,N_4848);
nor U6366 (N_6366,N_1740,N_3974);
nand U6367 (N_6367,N_271,N_4470);
xnor U6368 (N_6368,N_1048,N_4537);
xnor U6369 (N_6369,N_3841,N_2579);
and U6370 (N_6370,N_3353,N_2189);
and U6371 (N_6371,N_314,N_2002);
xor U6372 (N_6372,N_3919,N_1358);
and U6373 (N_6373,N_123,N_2510);
and U6374 (N_6374,N_4817,N_3963);
or U6375 (N_6375,N_4017,N_2502);
nor U6376 (N_6376,N_1981,N_3219);
nor U6377 (N_6377,N_4197,N_746);
or U6378 (N_6378,N_440,N_3791);
nand U6379 (N_6379,N_5,N_2881);
or U6380 (N_6380,N_4628,N_3623);
nor U6381 (N_6381,N_4925,N_3658);
nand U6382 (N_6382,N_4923,N_4825);
and U6383 (N_6383,N_2532,N_3307);
and U6384 (N_6384,N_1486,N_950);
and U6385 (N_6385,N_2158,N_1528);
or U6386 (N_6386,N_2153,N_1072);
and U6387 (N_6387,N_1571,N_426);
nor U6388 (N_6388,N_2243,N_206);
nand U6389 (N_6389,N_3511,N_4594);
or U6390 (N_6390,N_2874,N_121);
nor U6391 (N_6391,N_2497,N_4282);
xnor U6392 (N_6392,N_4074,N_4915);
and U6393 (N_6393,N_2215,N_3991);
nand U6394 (N_6394,N_1263,N_4055);
nor U6395 (N_6395,N_4300,N_1960);
nand U6396 (N_6396,N_161,N_2312);
or U6397 (N_6397,N_1813,N_899);
xor U6398 (N_6398,N_3817,N_3657);
nor U6399 (N_6399,N_2631,N_3010);
or U6400 (N_6400,N_2384,N_3907);
and U6401 (N_6401,N_2844,N_750);
nor U6402 (N_6402,N_2204,N_3222);
nand U6403 (N_6403,N_1747,N_2924);
and U6404 (N_6404,N_4287,N_3696);
nand U6405 (N_6405,N_3647,N_4897);
and U6406 (N_6406,N_2399,N_4454);
nand U6407 (N_6407,N_2457,N_4238);
nand U6408 (N_6408,N_3389,N_3784);
nand U6409 (N_6409,N_4016,N_1826);
nand U6410 (N_6410,N_2899,N_3412);
and U6411 (N_6411,N_274,N_1435);
nor U6412 (N_6412,N_2754,N_2128);
nor U6413 (N_6413,N_4609,N_2230);
or U6414 (N_6414,N_2863,N_2569);
and U6415 (N_6415,N_565,N_329);
xnor U6416 (N_6416,N_3272,N_914);
xnor U6417 (N_6417,N_4644,N_275);
nor U6418 (N_6418,N_2206,N_237);
or U6419 (N_6419,N_4600,N_2656);
nor U6420 (N_6420,N_1294,N_1942);
nand U6421 (N_6421,N_1890,N_1038);
nor U6422 (N_6422,N_4137,N_4132);
xnor U6423 (N_6423,N_212,N_4581);
or U6424 (N_6424,N_2422,N_1382);
nand U6425 (N_6425,N_2341,N_2082);
or U6426 (N_6426,N_4322,N_2582);
xnor U6427 (N_6427,N_4230,N_219);
xor U6428 (N_6428,N_2013,N_1357);
nand U6429 (N_6429,N_362,N_1982);
xor U6430 (N_6430,N_4788,N_3517);
and U6431 (N_6431,N_3513,N_2869);
or U6432 (N_6432,N_780,N_1863);
xor U6433 (N_6433,N_1743,N_4036);
xnor U6434 (N_6434,N_3809,N_2923);
xnor U6435 (N_6435,N_3813,N_3874);
or U6436 (N_6436,N_470,N_4866);
nor U6437 (N_6437,N_4029,N_2665);
or U6438 (N_6438,N_2822,N_1927);
xor U6439 (N_6439,N_2441,N_3195);
or U6440 (N_6440,N_871,N_1333);
nor U6441 (N_6441,N_153,N_1199);
xnor U6442 (N_6442,N_4308,N_4956);
and U6443 (N_6443,N_279,N_4145);
nor U6444 (N_6444,N_2299,N_3824);
and U6445 (N_6445,N_1452,N_489);
nor U6446 (N_6446,N_4641,N_1375);
nand U6447 (N_6447,N_2488,N_3003);
nand U6448 (N_6448,N_3863,N_1126);
or U6449 (N_6449,N_429,N_782);
nor U6450 (N_6450,N_922,N_4974);
xor U6451 (N_6451,N_2771,N_1649);
nor U6452 (N_6452,N_201,N_2014);
nor U6453 (N_6453,N_4754,N_802);
or U6454 (N_6454,N_3913,N_872);
nand U6455 (N_6455,N_658,N_3260);
xnor U6456 (N_6456,N_2613,N_4376);
xnor U6457 (N_6457,N_1775,N_4810);
or U6458 (N_6458,N_4717,N_2807);
xnor U6459 (N_6459,N_2835,N_1902);
nor U6460 (N_6460,N_2266,N_208);
and U6461 (N_6461,N_1867,N_3763);
or U6462 (N_6462,N_1162,N_1613);
and U6463 (N_6463,N_458,N_21);
or U6464 (N_6464,N_704,N_1882);
xnor U6465 (N_6465,N_439,N_1673);
nor U6466 (N_6466,N_4534,N_3337);
xnor U6467 (N_6467,N_567,N_3334);
and U6468 (N_6468,N_3968,N_3797);
or U6469 (N_6469,N_4995,N_402);
and U6470 (N_6470,N_1916,N_3589);
and U6471 (N_6471,N_654,N_4893);
nand U6472 (N_6472,N_1437,N_1057);
xor U6473 (N_6473,N_2847,N_1837);
or U6474 (N_6474,N_3943,N_4633);
nand U6475 (N_6475,N_100,N_4973);
nor U6476 (N_6476,N_4497,N_4275);
nand U6477 (N_6477,N_2458,N_3796);
or U6478 (N_6478,N_1297,N_325);
nor U6479 (N_6479,N_32,N_1068);
nand U6480 (N_6480,N_4729,N_3073);
and U6481 (N_6481,N_4369,N_533);
xnor U6482 (N_6482,N_116,N_2056);
and U6483 (N_6483,N_1945,N_4096);
or U6484 (N_6484,N_2428,N_1474);
or U6485 (N_6485,N_2276,N_2865);
nor U6486 (N_6486,N_3114,N_3284);
nand U6487 (N_6487,N_4545,N_785);
or U6488 (N_6488,N_2447,N_1904);
and U6489 (N_6489,N_4381,N_4023);
nor U6490 (N_6490,N_4596,N_4739);
xor U6491 (N_6491,N_427,N_2896);
xnor U6492 (N_6492,N_4249,N_4468);
or U6493 (N_6493,N_3414,N_447);
or U6494 (N_6494,N_4057,N_518);
nand U6495 (N_6495,N_2374,N_2566);
and U6496 (N_6496,N_1309,N_2846);
nand U6497 (N_6497,N_569,N_1694);
nand U6498 (N_6498,N_289,N_1193);
or U6499 (N_6499,N_4977,N_2563);
nand U6500 (N_6500,N_3954,N_1560);
or U6501 (N_6501,N_3169,N_1816);
or U6502 (N_6502,N_3420,N_4800);
and U6503 (N_6503,N_4691,N_307);
nor U6504 (N_6504,N_2030,N_391);
nor U6505 (N_6505,N_1508,N_4064);
and U6506 (N_6506,N_2435,N_2132);
xnor U6507 (N_6507,N_4416,N_1224);
or U6508 (N_6508,N_1179,N_1135);
and U6509 (N_6509,N_3679,N_2664);
nand U6510 (N_6510,N_2008,N_1039);
or U6511 (N_6511,N_2828,N_4557);
nand U6512 (N_6512,N_79,N_789);
xor U6513 (N_6513,N_1950,N_1186);
nand U6514 (N_6514,N_3032,N_384);
xor U6515 (N_6515,N_4682,N_166);
nand U6516 (N_6516,N_2575,N_1213);
or U6517 (N_6517,N_1205,N_146);
xor U6518 (N_6518,N_1987,N_2391);
xor U6519 (N_6519,N_2492,N_3512);
and U6520 (N_6520,N_2996,N_3564);
xor U6521 (N_6521,N_4549,N_791);
nand U6522 (N_6522,N_609,N_3031);
and U6523 (N_6523,N_2840,N_4863);
or U6524 (N_6524,N_3995,N_1231);
and U6525 (N_6525,N_3382,N_1752);
and U6526 (N_6526,N_2723,N_862);
nand U6527 (N_6527,N_1389,N_3315);
xor U6528 (N_6528,N_4490,N_929);
nor U6529 (N_6529,N_2344,N_3208);
or U6530 (N_6530,N_3480,N_4163);
and U6531 (N_6531,N_4204,N_3668);
and U6532 (N_6532,N_3616,N_4259);
nor U6533 (N_6533,N_1664,N_1903);
and U6534 (N_6534,N_3872,N_4449);
and U6535 (N_6535,N_2019,N_56);
nor U6536 (N_6536,N_4790,N_1951);
or U6537 (N_6537,N_3418,N_2589);
or U6538 (N_6538,N_2596,N_1210);
nand U6539 (N_6539,N_4044,N_571);
xor U6540 (N_6540,N_3256,N_3992);
xnor U6541 (N_6541,N_3153,N_1641);
nand U6542 (N_6542,N_3725,N_895);
and U6543 (N_6543,N_3810,N_584);
nor U6544 (N_6544,N_1892,N_2873);
and U6545 (N_6545,N_3973,N_2412);
and U6546 (N_6546,N_3531,N_2742);
nand U6547 (N_6547,N_4311,N_2839);
nor U6548 (N_6548,N_3078,N_34);
nor U6549 (N_6549,N_4655,N_3821);
xor U6550 (N_6550,N_4177,N_3655);
nand U6551 (N_6551,N_1279,N_1156);
or U6552 (N_6552,N_1036,N_3406);
xor U6553 (N_6553,N_4396,N_3687);
or U6554 (N_6554,N_1774,N_55);
xor U6555 (N_6555,N_2882,N_4962);
nor U6556 (N_6556,N_1400,N_2560);
xnor U6557 (N_6557,N_2326,N_2120);
xor U6558 (N_6558,N_3173,N_63);
xnor U6559 (N_6559,N_2962,N_4707);
nand U6560 (N_6560,N_1390,N_1285);
xor U6561 (N_6561,N_3102,N_3515);
xnor U6562 (N_6562,N_3421,N_4341);
or U6563 (N_6563,N_1874,N_3103);
or U6564 (N_6564,N_3629,N_4539);
and U6565 (N_6565,N_2183,N_4373);
nand U6566 (N_6566,N_701,N_4653);
xor U6567 (N_6567,N_4242,N_811);
xnor U6568 (N_6568,N_2831,N_1944);
nor U6569 (N_6569,N_2058,N_729);
and U6570 (N_6570,N_666,N_4441);
or U6571 (N_6571,N_4266,N_4363);
nand U6572 (N_6572,N_2324,N_310);
nand U6573 (N_6573,N_4041,N_4059);
xnor U6574 (N_6574,N_3997,N_1589);
xnor U6575 (N_6575,N_1657,N_2255);
nor U6576 (N_6576,N_3736,N_543);
nor U6577 (N_6577,N_4172,N_2307);
and U6578 (N_6578,N_2149,N_3598);
nor U6579 (N_6579,N_2593,N_1273);
and U6580 (N_6580,N_112,N_2858);
nand U6581 (N_6581,N_864,N_1353);
nand U6582 (N_6582,N_730,N_4357);
xor U6583 (N_6583,N_4827,N_2283);
or U6584 (N_6584,N_2103,N_1630);
nor U6585 (N_6585,N_3684,N_4085);
and U6586 (N_6586,N_3952,N_3726);
and U6587 (N_6587,N_953,N_1667);
or U6588 (N_6588,N_108,N_522);
or U6589 (N_6589,N_2065,N_4060);
and U6590 (N_6590,N_1648,N_2879);
and U6591 (N_6591,N_270,N_2164);
or U6592 (N_6592,N_3457,N_4869);
and U6593 (N_6593,N_2770,N_2535);
xor U6594 (N_6594,N_997,N_2685);
xor U6595 (N_6595,N_4386,N_949);
and U6596 (N_6596,N_861,N_2381);
or U6597 (N_6597,N_2729,N_4150);
nor U6598 (N_6598,N_4263,N_306);
and U6599 (N_6599,N_3723,N_35);
xor U6600 (N_6600,N_4831,N_4429);
or U6601 (N_6601,N_4887,N_4239);
or U6602 (N_6602,N_570,N_2150);
or U6603 (N_6603,N_615,N_1629);
nand U6604 (N_6604,N_3021,N_4921);
xnor U6605 (N_6605,N_4507,N_883);
nor U6606 (N_6606,N_3714,N_1399);
nand U6607 (N_6607,N_2172,N_4262);
xnor U6608 (N_6608,N_2548,N_3454);
xnor U6609 (N_6609,N_1976,N_4);
or U6610 (N_6610,N_18,N_646);
or U6611 (N_6611,N_3920,N_3946);
or U6612 (N_6612,N_99,N_4427);
or U6613 (N_6613,N_2930,N_4595);
nor U6614 (N_6614,N_2366,N_3733);
or U6615 (N_6615,N_2711,N_2690);
xor U6616 (N_6616,N_547,N_1282);
xor U6617 (N_6617,N_1627,N_1373);
or U6618 (N_6618,N_1949,N_4984);
or U6619 (N_6619,N_4926,N_2346);
nor U6620 (N_6620,N_4587,N_1791);
and U6621 (N_6621,N_1728,N_1592);
xnor U6622 (N_6622,N_958,N_700);
nand U6623 (N_6623,N_913,N_2940);
nand U6624 (N_6624,N_3742,N_4936);
xnor U6625 (N_6625,N_1712,N_1238);
and U6626 (N_6626,N_2772,N_817);
and U6627 (N_6627,N_4460,N_524);
and U6628 (N_6628,N_2134,N_3898);
nand U6629 (N_6629,N_159,N_1781);
xor U6630 (N_6630,N_2284,N_378);
nand U6631 (N_6631,N_1264,N_3481);
xor U6632 (N_6632,N_1112,N_4694);
and U6633 (N_6633,N_444,N_542);
nand U6634 (N_6634,N_3593,N_4706);
nand U6635 (N_6635,N_2939,N_826);
nor U6636 (N_6636,N_4986,N_1804);
nor U6637 (N_6637,N_2662,N_1930);
nand U6638 (N_6638,N_3177,N_2315);
or U6639 (N_6639,N_1846,N_4981);
nand U6640 (N_6640,N_1225,N_409);
xor U6641 (N_6641,N_720,N_3020);
and U6642 (N_6642,N_1527,N_318);
xnor U6643 (N_6643,N_343,N_611);
and U6644 (N_6644,N_4475,N_1082);
xor U6645 (N_6645,N_1066,N_354);
nand U6646 (N_6646,N_1682,N_4461);
nor U6647 (N_6647,N_4241,N_2686);
and U6648 (N_6648,N_2005,N_4976);
nand U6649 (N_6649,N_3588,N_4550);
and U6650 (N_6650,N_1602,N_2877);
and U6651 (N_6651,N_3213,N_3893);
or U6652 (N_6652,N_527,N_2212);
nand U6653 (N_6653,N_3350,N_3363);
and U6654 (N_6654,N_4799,N_4842);
xnor U6655 (N_6655,N_2782,N_4716);
or U6656 (N_6656,N_3160,N_1035);
nand U6657 (N_6657,N_3775,N_3672);
nand U6658 (N_6658,N_4951,N_1040);
or U6659 (N_6659,N_4590,N_2990);
or U6660 (N_6660,N_2209,N_294);
nor U6661 (N_6661,N_3223,N_4886);
nor U6662 (N_6662,N_3830,N_2570);
nor U6663 (N_6663,N_3654,N_1939);
nand U6664 (N_6664,N_2342,N_4108);
and U6665 (N_6665,N_2086,N_2403);
nand U6666 (N_6666,N_3247,N_3936);
xor U6667 (N_6667,N_4775,N_1830);
nor U6668 (N_6668,N_2354,N_4076);
nand U6669 (N_6669,N_1841,N_4972);
nor U6670 (N_6670,N_2235,N_4486);
and U6671 (N_6671,N_2676,N_3945);
and U6672 (N_6672,N_2848,N_1409);
nand U6673 (N_6673,N_2295,N_850);
nor U6674 (N_6674,N_4918,N_1191);
or U6675 (N_6675,N_1800,N_192);
nor U6676 (N_6676,N_2017,N_3001);
or U6677 (N_6677,N_4961,N_1645);
nor U6678 (N_6678,N_2773,N_1269);
nand U6679 (N_6679,N_2397,N_114);
nand U6680 (N_6680,N_160,N_2625);
or U6681 (N_6681,N_4814,N_1507);
nor U6682 (N_6682,N_3730,N_994);
and U6683 (N_6683,N_3558,N_4753);
nor U6684 (N_6684,N_2630,N_1401);
and U6685 (N_6685,N_4193,N_1102);
or U6686 (N_6686,N_3139,N_0);
and U6687 (N_6687,N_1819,N_1750);
nor U6688 (N_6688,N_281,N_1149);
and U6689 (N_6689,N_2453,N_3659);
xor U6690 (N_6690,N_629,N_4436);
nor U6691 (N_6691,N_4678,N_2958);
nand U6692 (N_6692,N_1678,N_1689);
nor U6693 (N_6693,N_10,N_1788);
xor U6694 (N_6694,N_4190,N_2789);
nor U6695 (N_6695,N_696,N_4061);
and U6696 (N_6696,N_359,N_1986);
or U6697 (N_6697,N_1106,N_1300);
or U6698 (N_6698,N_2680,N_1501);
nand U6699 (N_6699,N_4839,N_3209);
and U6700 (N_6700,N_3619,N_1089);
xor U6701 (N_6701,N_4812,N_3263);
xor U6702 (N_6702,N_298,N_1079);
nor U6703 (N_6703,N_4690,N_2641);
and U6704 (N_6704,N_1295,N_1176);
nor U6705 (N_6705,N_2495,N_2653);
nand U6706 (N_6706,N_2647,N_157);
or U6707 (N_6707,N_3906,N_4231);
or U6708 (N_6708,N_963,N_3451);
and U6709 (N_6709,N_4457,N_1662);
nand U6710 (N_6710,N_3368,N_3897);
and U6711 (N_6711,N_3023,N_2045);
or U6712 (N_6712,N_4565,N_3275);
or U6713 (N_6713,N_2093,N_3768);
or U6714 (N_6714,N_1235,N_625);
and U6715 (N_6715,N_4695,N_2991);
nand U6716 (N_6716,N_3495,N_4355);
and U6717 (N_6717,N_4667,N_3311);
nand U6718 (N_6718,N_3410,N_4526);
nand U6719 (N_6719,N_3567,N_38);
and U6720 (N_6720,N_3798,N_3644);
xnor U6721 (N_6721,N_1579,N_1767);
and U6722 (N_6722,N_1876,N_593);
nand U6723 (N_6723,N_892,N_4103);
and U6724 (N_6724,N_1907,N_592);
nand U6725 (N_6725,N_1623,N_848);
and U6726 (N_6726,N_744,N_4089);
nand U6727 (N_6727,N_3245,N_2987);
nor U6728 (N_6728,N_3393,N_3268);
xnor U6729 (N_6729,N_4056,N_3626);
nor U6730 (N_6730,N_3609,N_1202);
nor U6731 (N_6731,N_185,N_2801);
or U6732 (N_6732,N_3339,N_1705);
or U6733 (N_6733,N_2602,N_1319);
xor U6734 (N_6734,N_4439,N_2426);
and U6735 (N_6735,N_4685,N_3461);
and U6736 (N_6736,N_1607,N_2512);
and U6737 (N_6737,N_903,N_2997);
xnor U6738 (N_6738,N_1441,N_2241);
nor U6739 (N_6739,N_4860,N_4541);
nand U6740 (N_6740,N_2768,N_1355);
xnor U6741 (N_6741,N_1758,N_1178);
xor U6742 (N_6742,N_3044,N_521);
and U6743 (N_6743,N_1161,N_104);
or U6744 (N_6744,N_4134,N_1656);
or U6745 (N_6745,N_4426,N_3039);
nor U6746 (N_6746,N_158,N_2737);
xor U6747 (N_6747,N_4051,N_4397);
nand U6748 (N_6748,N_1983,N_1557);
xor U6749 (N_6749,N_2949,N_2868);
nor U6750 (N_6750,N_1424,N_106);
nor U6751 (N_6751,N_460,N_1046);
or U6752 (N_6752,N_3249,N_671);
and U6753 (N_6753,N_1568,N_698);
nand U6754 (N_6754,N_3875,N_1387);
nand U6755 (N_6755,N_1371,N_3548);
nand U6756 (N_6756,N_1475,N_1921);
or U6757 (N_6757,N_4123,N_1383);
xor U6758 (N_6758,N_3022,N_2806);
nor U6759 (N_6759,N_4865,N_3423);
nand U6760 (N_6760,N_1197,N_3758);
nor U6761 (N_6761,N_2792,N_2956);
nand U6762 (N_6762,N_4824,N_2739);
or U6763 (N_6763,N_3397,N_742);
or U6764 (N_6764,N_564,N_2225);
nand U6765 (N_6765,N_2741,N_437);
nor U6766 (N_6766,N_2099,N_1064);
and U6767 (N_6767,N_4491,N_927);
or U6768 (N_6768,N_2855,N_2506);
nand U6769 (N_6769,N_183,N_2894);
nand U6770 (N_6770,N_2809,N_2963);
or U6771 (N_6771,N_501,N_773);
nor U6772 (N_6772,N_1900,N_77);
nor U6773 (N_6773,N_1760,N_4143);
nor U6774 (N_6774,N_3074,N_1232);
xor U6775 (N_6775,N_349,N_371);
nor U6776 (N_6776,N_1364,N_4265);
nand U6777 (N_6777,N_4114,N_39);
or U6778 (N_6778,N_3518,N_4383);
and U6779 (N_6779,N_54,N_3441);
nand U6780 (N_6780,N_1095,N_4053);
xnor U6781 (N_6781,N_1726,N_4093);
nor U6782 (N_6782,N_124,N_4246);
nand U6783 (N_6783,N_529,N_1194);
nand U6784 (N_6784,N_1233,N_737);
nand U6785 (N_6785,N_3168,N_412);
and U6786 (N_6786,N_602,N_2320);
nand U6787 (N_6787,N_365,N_2285);
and U6788 (N_6788,N_620,N_1691);
xor U6789 (N_6789,N_394,N_865);
or U6790 (N_6790,N_1188,N_483);
and U6791 (N_6791,N_3940,N_1055);
or U6792 (N_6792,N_2900,N_4237);
nor U6793 (N_6793,N_4732,N_1420);
nand U6794 (N_6794,N_4038,N_296);
nor U6795 (N_6795,N_1190,N_739);
and U6796 (N_6796,N_267,N_2117);
and U6797 (N_6797,N_3949,N_4465);
nand U6798 (N_6798,N_3745,N_4642);
and U6799 (N_6799,N_3615,N_555);
or U6800 (N_6800,N_4011,N_3261);
and U6801 (N_6801,N_4006,N_1431);
nor U6802 (N_6802,N_500,N_1469);
xor U6803 (N_6803,N_987,N_2228);
nor U6804 (N_6804,N_1184,N_3187);
nor U6805 (N_6805,N_204,N_3690);
xnor U6806 (N_6806,N_1283,N_2983);
nor U6807 (N_6807,N_4290,N_3455);
nand U6808 (N_6808,N_1956,N_3343);
and U6809 (N_6809,N_3138,N_3057);
xor U6810 (N_6810,N_3883,N_1961);
xnor U6811 (N_6811,N_4019,N_1354);
nor U6812 (N_6812,N_2733,N_47);
and U6813 (N_6813,N_2072,N_3207);
xor U6814 (N_6814,N_1272,N_4253);
nand U6815 (N_6815,N_2119,N_3504);
xnor U6816 (N_6816,N_2756,N_4510);
and U6817 (N_6817,N_1250,N_4052);
nor U6818 (N_6818,N_3038,N_239);
or U6819 (N_6819,N_4563,N_4310);
xor U6820 (N_6820,N_3568,N_3502);
or U6821 (N_6821,N_3899,N_1772);
xor U6822 (N_6822,N_4760,N_728);
or U6823 (N_6823,N_1010,N_91);
nor U6824 (N_6824,N_640,N_2245);
and U6825 (N_6825,N_2214,N_4679);
or U6826 (N_6826,N_4689,N_2253);
xnor U6827 (N_6827,N_4566,N_1688);
nor U6828 (N_6828,N_1696,N_4318);
xnor U6829 (N_6829,N_3544,N_843);
xor U6830 (N_6830,N_3097,N_17);
and U6831 (N_6831,N_3226,N_1763);
nand U6832 (N_6832,N_1993,N_4315);
or U6833 (N_6833,N_2623,N_3881);
and U6834 (N_6834,N_3000,N_844);
xor U6835 (N_6835,N_888,N_1994);
and U6836 (N_6836,N_1175,N_1566);
nand U6837 (N_6837,N_3474,N_968);
nand U6838 (N_6838,N_1680,N_3571);
nor U6839 (N_6839,N_4187,N_4252);
and U6840 (N_6840,N_4525,N_4517);
nor U6841 (N_6841,N_392,N_2184);
xnor U6842 (N_6842,N_2405,N_3465);
nand U6843 (N_6843,N_4434,N_3411);
or U6844 (N_6844,N_3702,N_4024);
or U6845 (N_6845,N_2290,N_61);
or U6846 (N_6846,N_4116,N_898);
and U6847 (N_6847,N_1477,N_1520);
xnor U6848 (N_6848,N_1525,N_1476);
nand U6849 (N_6849,N_3781,N_3976);
nand U6850 (N_6850,N_818,N_3276);
or U6851 (N_6851,N_4513,N_1844);
nand U6852 (N_6852,N_2574,N_3110);
and U6853 (N_6853,N_3509,N_2713);
nand U6854 (N_6854,N_1943,N_1128);
or U6855 (N_6855,N_1880,N_3176);
or U6856 (N_6856,N_4227,N_4803);
xnor U6857 (N_6857,N_1030,N_3838);
nor U6858 (N_6858,N_4213,N_4511);
or U6859 (N_6859,N_1317,N_2456);
nor U6860 (N_6860,N_1479,N_2551);
nand U6861 (N_6861,N_254,N_2417);
or U6862 (N_6862,N_630,N_2076);
and U6863 (N_6863,N_4579,N_2978);
and U6864 (N_6864,N_792,N_3612);
nand U6865 (N_6865,N_4228,N_3573);
and U6866 (N_6866,N_3636,N_3632);
nand U6867 (N_6867,N_867,N_1105);
nor U6868 (N_6868,N_631,N_1144);
nand U6869 (N_6869,N_4048,N_3346);
xor U6870 (N_6870,N_3277,N_3155);
nor U6871 (N_6871,N_3718,N_2620);
nor U6872 (N_6872,N_3676,N_2697);
xnor U6873 (N_6873,N_3827,N_3537);
nand U6874 (N_6874,N_397,N_4584);
xnor U6875 (N_6875,N_3622,N_854);
nand U6876 (N_6876,N_2123,N_1086);
and U6877 (N_6877,N_1289,N_1221);
or U6878 (N_6878,N_1738,N_3786);
and U6879 (N_6879,N_4336,N_442);
or U6880 (N_6880,N_1336,N_4146);
or U6881 (N_6881,N_3301,N_661);
xnor U6882 (N_6882,N_1473,N_3422);
or U6883 (N_6883,N_1410,N_2554);
nand U6884 (N_6884,N_3909,N_4684);
xor U6885 (N_6885,N_3849,N_1260);
nor U6886 (N_6886,N_2673,N_1849);
and U6887 (N_6887,N_4905,N_381);
nand U6888 (N_6888,N_828,N_3773);
and U6889 (N_6889,N_2033,N_4916);
xnor U6890 (N_6890,N_2410,N_12);
and U6891 (N_6891,N_875,N_4045);
and U6892 (N_6892,N_2096,N_3641);
nand U6893 (N_6893,N_743,N_36);
or U6894 (N_6894,N_1709,N_1413);
and U6895 (N_6895,N_2054,N_2200);
nor U6896 (N_6896,N_680,N_3795);
nand U6897 (N_6897,N_1820,N_2386);
or U6898 (N_6898,N_2459,N_2475);
nor U6899 (N_6899,N_1291,N_4575);
nand U6900 (N_6900,N_4268,N_2906);
xnor U6901 (N_6901,N_4969,N_1243);
nor U6902 (N_6902,N_2496,N_2905);
nor U6903 (N_6903,N_1396,N_2986);
xor U6904 (N_6904,N_3703,N_4749);
and U6905 (N_6905,N_1468,N_2277);
and U6906 (N_6906,N_1941,N_4032);
xnor U6907 (N_6907,N_4073,N_3333);
and U6908 (N_6908,N_2256,N_1940);
or U6909 (N_6909,N_3233,N_1015);
or U6910 (N_6910,N_2427,N_3098);
and U6911 (N_6911,N_2359,N_3435);
and U6912 (N_6912,N_2672,N_3349);
xor U6913 (N_6913,N_3100,N_1007);
and U6914 (N_6914,N_169,N_2208);
nand U6915 (N_6915,N_1177,N_3697);
xnor U6916 (N_6916,N_3359,N_1583);
nor U6917 (N_6917,N_4214,N_2129);
or U6918 (N_6918,N_3500,N_669);
nor U6919 (N_6919,N_508,N_4523);
nand U6920 (N_6920,N_2262,N_2931);
xnor U6921 (N_6921,N_3116,N_3269);
and U6922 (N_6922,N_1795,N_2935);
or U6923 (N_6923,N_1702,N_4639);
xor U6924 (N_6924,N_1167,N_1923);
nor U6925 (N_6925,N_1147,N_3630);
nor U6926 (N_6926,N_961,N_1522);
nand U6927 (N_6927,N_4083,N_2059);
and U6928 (N_6928,N_3181,N_3555);
or U6929 (N_6929,N_4260,N_4674);
and U6930 (N_6930,N_3812,N_1755);
xnor U6931 (N_6931,N_3833,N_210);
or U6932 (N_6932,N_4350,N_1847);
nand U6933 (N_6933,N_156,N_19);
nand U6934 (N_6934,N_1303,N_4970);
xor U6935 (N_6935,N_278,N_4752);
nor U6936 (N_6936,N_2961,N_138);
xor U6937 (N_6937,N_2926,N_601);
nor U6938 (N_6938,N_4375,N_4630);
nand U6939 (N_6939,N_1914,N_1141);
nor U6940 (N_6940,N_2471,N_1259);
and U6941 (N_6941,N_3487,N_3620);
and U6942 (N_6942,N_2026,N_775);
nor U6943 (N_6943,N_70,N_465);
xnor U6944 (N_6944,N_2329,N_4400);
nor U6945 (N_6945,N_2293,N_4735);
and U6946 (N_6946,N_3405,N_4232);
xnor U6947 (N_6947,N_4602,N_3006);
nor U6948 (N_6948,N_4410,N_3446);
and U6949 (N_6949,N_2291,N_604);
xnor U6950 (N_6950,N_4728,N_3947);
nor U6951 (N_6951,N_3669,N_3442);
nand U6952 (N_6952,N_3288,N_3862);
or U6953 (N_6953,N_4614,N_4636);
nor U6954 (N_6954,N_2402,N_1695);
nor U6955 (N_6955,N_2813,N_3347);
nor U6956 (N_6956,N_4677,N_4399);
or U6957 (N_6957,N_924,N_3212);
or U6958 (N_6958,N_2553,N_2265);
and U6959 (N_6959,N_1814,N_480);
or U6960 (N_6960,N_645,N_591);
and U6961 (N_6961,N_712,N_3460);
xnor U6962 (N_6962,N_2688,N_3163);
nand U6963 (N_6963,N_2382,N_2218);
or U6964 (N_6964,N_4218,N_1407);
xnor U6965 (N_6965,N_1063,N_3918);
nor U6966 (N_6966,N_900,N_1561);
xor U6967 (N_6967,N_4819,N_3704);
xnor U6968 (N_6968,N_3014,N_4188);
xnor U6969 (N_6969,N_3053,N_3450);
xor U6970 (N_6970,N_2959,N_2401);
xnor U6971 (N_6971,N_490,N_1150);
nor U6972 (N_6972,N_2363,N_481);
and U6973 (N_6973,N_425,N_3175);
xor U6974 (N_6974,N_44,N_2936);
or U6975 (N_6975,N_1158,N_4521);
and U6976 (N_6976,N_774,N_1998);
and U6977 (N_6977,N_2016,N_1671);
xor U6978 (N_6978,N_3371,N_3643);
xor U6979 (N_6979,N_1886,N_943);
or U6980 (N_6980,N_3327,N_4878);
nand U6981 (N_6981,N_3720,N_2455);
nor U6982 (N_6982,N_1764,N_4018);
and U6983 (N_6983,N_4494,N_3855);
or U6984 (N_6984,N_4283,N_1779);
xor U6985 (N_6985,N_4067,N_477);
xnor U6986 (N_6986,N_769,N_342);
and U6987 (N_6987,N_1100,N_1083);
nor U6988 (N_6988,N_1222,N_1727);
or U6989 (N_6989,N_226,N_2594);
nor U6990 (N_6990,N_1526,N_3592);
xnor U6991 (N_6991,N_4724,N_3965);
and U6992 (N_6992,N_2833,N_894);
nand U6993 (N_6993,N_4660,N_2654);
or U6994 (N_6994,N_1362,N_472);
xnor U6995 (N_6995,N_523,N_181);
or U6996 (N_6996,N_4480,N_2333);
nand U6997 (N_6997,N_3750,N_2067);
nand U6998 (N_6998,N_4112,N_140);
or U6999 (N_6999,N_2611,N_3808);
nor U7000 (N_7000,N_4387,N_4746);
nor U7001 (N_7001,N_4730,N_4681);
xnor U7002 (N_7002,N_3440,N_2249);
nand U7003 (N_7003,N_657,N_1898);
and U7004 (N_7004,N_3122,N_2465);
nand U7005 (N_7005,N_1006,N_288);
xnor U7006 (N_7006,N_4589,N_2055);
nor U7007 (N_7007,N_1928,N_4459);
nor U7008 (N_7008,N_31,N_3133);
nor U7009 (N_7009,N_3793,N_734);
nand U7010 (N_7010,N_1523,N_2133);
and U7011 (N_7011,N_4040,N_3438);
nor U7012 (N_7012,N_3484,N_3799);
nor U7013 (N_7013,N_3313,N_73);
nor U7014 (N_7014,N_678,N_3847);
and U7015 (N_7015,N_610,N_3060);
nor U7016 (N_7016,N_4598,N_4418);
xor U7017 (N_7017,N_3123,N_293);
and U7018 (N_7018,N_4223,N_1043);
and U7019 (N_7019,N_4288,N_4850);
or U7020 (N_7020,N_20,N_1200);
and U7021 (N_7021,N_1427,N_1240);
nand U7022 (N_7022,N_2080,N_3453);
nand U7023 (N_7023,N_374,N_1677);
xnor U7024 (N_7024,N_1467,N_103);
nand U7025 (N_7025,N_1346,N_2316);
nand U7026 (N_7026,N_2186,N_4666);
and U7027 (N_7027,N_2994,N_2383);
nor U7028 (N_7028,N_3663,N_3854);
nor U7029 (N_7029,N_4680,N_2998);
xnor U7030 (N_7030,N_2545,N_1070);
xor U7031 (N_7031,N_3150,N_1448);
or U7032 (N_7032,N_3055,N_4432);
or U7033 (N_7033,N_4196,N_2351);
nor U7034 (N_7034,N_838,N_4153);
xnor U7035 (N_7035,N_4745,N_3467);
nand U7036 (N_7036,N_1426,N_2748);
and U7037 (N_7037,N_545,N_4007);
nand U7038 (N_7038,N_3448,N_3424);
or U7039 (N_7039,N_98,N_404);
and U7040 (N_7040,N_3552,N_109);
nor U7041 (N_7041,N_3425,N_3843);
xor U7042 (N_7042,N_4025,N_4414);
xor U7043 (N_7043,N_3090,N_3826);
or U7044 (N_7044,N_2687,N_767);
and U7045 (N_7045,N_3291,N_4377);
xor U7046 (N_7046,N_4935,N_1905);
nand U7047 (N_7047,N_504,N_3027);
and U7048 (N_7048,N_1751,N_411);
nor U7049 (N_7049,N_2836,N_2529);
nor U7050 (N_7050,N_4725,N_3789);
nand U7051 (N_7051,N_557,N_841);
and U7052 (N_7052,N_2340,N_4624);
xnor U7053 (N_7053,N_2719,N_673);
nand U7054 (N_7054,N_2169,N_619);
or U7055 (N_7055,N_321,N_4345);
nor U7056 (N_7056,N_919,N_4184);
or U7057 (N_7057,N_947,N_441);
or U7058 (N_7058,N_3306,N_4343);
nor U7059 (N_7059,N_4744,N_168);
or U7060 (N_7060,N_2829,N_2929);
or U7061 (N_7061,N_1780,N_4813);
nand U7062 (N_7062,N_2546,N_1163);
nor U7063 (N_7063,N_1249,N_328);
xnor U7064 (N_7064,N_3145,N_1979);
or U7065 (N_7065,N_2603,N_2794);
and U7066 (N_7066,N_4608,N_2910);
and U7067 (N_7067,N_2640,N_4030);
nand U7068 (N_7068,N_2171,N_4767);
xnor U7069 (N_7069,N_1306,N_4519);
nor U7070 (N_7070,N_2323,N_1166);
and U7071 (N_7071,N_886,N_4577);
nand U7072 (N_7072,N_4635,N_4696);
or U7073 (N_7073,N_3581,N_4034);
xor U7074 (N_7074,N_4904,N_495);
and U7075 (N_7075,N_1585,N_3345);
or U7076 (N_7076,N_2021,N_4295);
nor U7077 (N_7077,N_1631,N_3016);
nor U7078 (N_7078,N_4773,N_1506);
and U7079 (N_7079,N_2074,N_331);
nor U7080 (N_7080,N_1827,N_2849);
xnor U7081 (N_7081,N_3601,N_1406);
or U7082 (N_7082,N_241,N_3538);
nor U7083 (N_7083,N_3473,N_2793);
and U7084 (N_7084,N_1157,N_1451);
nand U7085 (N_7085,N_2948,N_1668);
nand U7086 (N_7086,N_515,N_3738);
xor U7087 (N_7087,N_1372,N_3876);
and U7088 (N_7088,N_3430,N_563);
and U7089 (N_7089,N_302,N_3149);
or U7090 (N_7090,N_3403,N_3498);
or U7091 (N_7091,N_1164,N_438);
nand U7092 (N_7092,N_3043,N_3007);
and U7093 (N_7093,N_1729,N_1377);
or U7094 (N_7094,N_2232,N_2706);
or U7095 (N_7095,N_3771,N_4859);
and U7096 (N_7096,N_4149,N_2618);
or U7097 (N_7097,N_3526,N_4331);
and U7098 (N_7098,N_2663,N_3706);
nand U7099 (N_7099,N_3649,N_42);
nor U7100 (N_7100,N_928,N_4092);
nor U7101 (N_7101,N_49,N_4769);
xor U7102 (N_7102,N_999,N_4072);
and U7103 (N_7103,N_1218,N_4808);
xnor U7104 (N_7104,N_4401,N_3971);
xnor U7105 (N_7105,N_740,N_3928);
nand U7106 (N_7106,N_2009,N_1369);
or U7107 (N_7107,N_2377,N_375);
nand U7108 (N_7108,N_2485,N_4236);
nand U7109 (N_7109,N_52,N_1789);
and U7110 (N_7110,N_2450,N_4883);
nor U7111 (N_7111,N_4500,N_4450);
xor U7112 (N_7112,N_4216,N_125);
nor U7113 (N_7113,N_3026,N_656);
or U7114 (N_7114,N_2070,N_1253);
nor U7115 (N_7115,N_4180,N_2573);
or U7116 (N_7116,N_2645,N_468);
xnor U7117 (N_7117,N_1590,N_4966);
and U7118 (N_7118,N_2811,N_4327);
or U7119 (N_7119,N_677,N_167);
or U7120 (N_7120,N_845,N_1398);
nand U7121 (N_7121,N_3089,N_4335);
xnor U7122 (N_7122,N_51,N_475);
xor U7123 (N_7123,N_4493,N_2778);
xor U7124 (N_7124,N_1031,N_134);
or U7125 (N_7125,N_230,N_4140);
nand U7126 (N_7126,N_2885,N_544);
nor U7127 (N_7127,N_3206,N_4835);
nand U7128 (N_7128,N_2597,N_420);
nor U7129 (N_7129,N_682,N_3967);
and U7130 (N_7130,N_1069,N_141);
and U7131 (N_7131,N_902,N_148);
and U7132 (N_7132,N_2531,N_4889);
xnor U7133 (N_7133,N_175,N_2699);
xnor U7134 (N_7134,N_2724,N_3912);
or U7135 (N_7135,N_516,N_794);
xnor U7136 (N_7136,N_1697,N_1699);
and U7137 (N_7137,N_1099,N_1071);
nor U7138 (N_7138,N_1693,N_4342);
and U7139 (N_7139,N_2162,N_4648);
nor U7140 (N_7140,N_1171,N_551);
or U7141 (N_7141,N_1759,N_2449);
or U7142 (N_7142,N_1349,N_3868);
and U7143 (N_7143,N_3569,N_366);
or U7144 (N_7144,N_1713,N_1280);
nor U7145 (N_7145,N_4687,N_3921);
or U7146 (N_7146,N_4479,N_1966);
xor U7147 (N_7147,N_82,N_1129);
or U7148 (N_7148,N_4217,N_1187);
nor U7149 (N_7149,N_4274,N_1421);
and U7150 (N_7150,N_3202,N_4560);
and U7151 (N_7151,N_1931,N_3294);
nand U7152 (N_7152,N_1037,N_827);
or U7153 (N_7153,N_4546,N_1132);
xor U7154 (N_7154,N_4437,N_3890);
xnor U7155 (N_7155,N_2638,N_1851);
nand U7156 (N_7156,N_3278,N_1274);
or U7157 (N_7157,N_107,N_3700);
or U7158 (N_7158,N_4141,N_4968);
xnor U7159 (N_7159,N_2876,N_632);
or U7160 (N_7160,N_3929,N_2010);
or U7161 (N_7161,N_220,N_4097);
xor U7162 (N_7162,N_2857,N_1180);
and U7163 (N_7163,N_3280,N_2503);
nor U7164 (N_7164,N_2636,N_4121);
or U7165 (N_7165,N_2500,N_196);
or U7166 (N_7166,N_2964,N_724);
nand U7167 (N_7167,N_4922,N_1266);
nor U7168 (N_7168,N_2824,N_4127);
nor U7169 (N_7169,N_1828,N_781);
and U7170 (N_7170,N_4302,N_4281);
nand U7171 (N_7171,N_3137,N_2891);
xnor U7172 (N_7172,N_1117,N_3234);
and U7173 (N_7173,N_4535,N_147);
nand U7174 (N_7174,N_1098,N_292);
or U7175 (N_7175,N_1968,N_3433);
xor U7176 (N_7176,N_2452,N_3469);
xnor U7177 (N_7177,N_3065,N_3366);
and U7178 (N_7178,N_1854,N_4312);
and U7179 (N_7179,N_2866,N_2305);
xnor U7180 (N_7180,N_3075,N_2089);
xor U7181 (N_7181,N_415,N_1459);
and U7182 (N_7182,N_2947,N_1839);
nand U7183 (N_7183,N_330,N_346);
xnor U7184 (N_7184,N_492,N_2621);
xnor U7185 (N_7185,N_83,N_2592);
xor U7186 (N_7186,N_3861,N_684);
or U7187 (N_7187,N_2286,N_1796);
xor U7188 (N_7188,N_3012,N_4160);
or U7189 (N_7189,N_3977,N_1929);
nor U7190 (N_7190,N_3892,N_3790);
and U7191 (N_7191,N_3456,N_4963);
or U7192 (N_7192,N_2615,N_1457);
and U7193 (N_7193,N_731,N_4348);
nand U7194 (N_7194,N_1337,N_3186);
nor U7195 (N_7195,N_1461,N_622);
nor U7196 (N_7196,N_3677,N_4176);
or U7197 (N_7197,N_2137,N_3115);
or U7198 (N_7198,N_1047,N_1703);
nand U7199 (N_7199,N_876,N_946);
and U7200 (N_7200,N_2590,N_1599);
and U7201 (N_7201,N_3895,N_4676);
nand U7202 (N_7202,N_942,N_451);
and U7203 (N_7203,N_344,N_2483);
and U7204 (N_7204,N_1511,N_4395);
and U7205 (N_7205,N_3579,N_3982);
nor U7206 (N_7206,N_3004,N_1534);
xnor U7207 (N_7207,N_4364,N_568);
nor U7208 (N_7208,N_2608,N_4117);
or U7209 (N_7209,N_1806,N_75);
nand U7210 (N_7210,N_2668,N_215);
nor U7211 (N_7211,N_1018,N_1734);
and U7212 (N_7212,N_3009,N_3201);
nand U7213 (N_7213,N_2826,N_191);
or U7214 (N_7214,N_1716,N_122);
nand U7215 (N_7215,N_2350,N_665);
and U7216 (N_7216,N_2534,N_3728);
xor U7217 (N_7217,N_548,N_3525);
and U7218 (N_7218,N_2895,N_1216);
nor U7219 (N_7219,N_4978,N_3449);
nor U7220 (N_7220,N_3076,N_1429);
and U7221 (N_7221,N_2652,N_1503);
or U7222 (N_7222,N_3539,N_4558);
nor U7223 (N_7223,N_92,N_2224);
xnor U7224 (N_7224,N_4175,N_3709);
xnor U7225 (N_7225,N_1594,N_1261);
xor U7226 (N_7226,N_3554,N_2937);
xor U7227 (N_7227,N_2728,N_2614);
nor U7228 (N_7228,N_2101,N_2219);
nor U7229 (N_7229,N_189,N_2818);
nand U7230 (N_7230,N_2170,N_1895);
and U7231 (N_7231,N_1685,N_1838);
and U7232 (N_7232,N_3193,N_4351);
nor U7233 (N_7233,N_952,N_3344);
nand U7234 (N_7234,N_4834,N_4105);
nor U7235 (N_7235,N_1350,N_335);
and U7236 (N_7236,N_4555,N_2231);
nand U7237 (N_7237,N_1985,N_1822);
nand U7238 (N_7238,N_1947,N_618);
and U7239 (N_7239,N_2918,N_4845);
xnor U7240 (N_7240,N_126,N_50);
nand U7241 (N_7241,N_726,N_813);
xor U7242 (N_7242,N_1229,N_2902);
or U7243 (N_7243,N_2567,N_3547);
xor U7244 (N_7244,N_4443,N_4042);
or U7245 (N_7245,N_471,N_4485);
xor U7246 (N_7246,N_1097,N_600);
and U7247 (N_7247,N_4708,N_2298);
or U7248 (N_7248,N_3985,N_3431);
nor U7249 (N_7249,N_4611,N_2912);
nor U7250 (N_7250,N_1715,N_4170);
or U7251 (N_7251,N_1969,N_1060);
nor U7252 (N_7252,N_228,N_152);
nand U7253 (N_7253,N_738,N_2915);
nand U7254 (N_7254,N_977,N_388);
xnor U7255 (N_7255,N_2115,N_2601);
or U7256 (N_7256,N_1440,N_1865);
xnor U7257 (N_7257,N_2211,N_695);
and U7258 (N_7258,N_770,N_2521);
xor U7259 (N_7259,N_703,N_1146);
or U7260 (N_7260,N_2908,N_651);
nand U7261 (N_7261,N_3905,N_2207);
or U7262 (N_7262,N_4423,N_3653);
xnor U7263 (N_7263,N_2240,N_4487);
nand U7264 (N_7264,N_1934,N_4091);
xnor U7265 (N_7265,N_4671,N_2571);
nor U7266 (N_7266,N_4009,N_1109);
or U7267 (N_7267,N_808,N_1706);
nand U7268 (N_7268,N_3586,N_1544);
nor U7269 (N_7269,N_4618,N_4181);
nand U7270 (N_7270,N_376,N_3071);
nand U7271 (N_7271,N_1428,N_4258);
and U7272 (N_7272,N_4171,N_3042);
and U7273 (N_7273,N_1562,N_2974);
nand U7274 (N_7274,N_3215,N_4482);
nor U7275 (N_7275,N_1974,N_260);
and U7276 (N_7276,N_268,N_1316);
nor U7277 (N_7277,N_4178,N_3036);
or U7278 (N_7278,N_1379,N_1332);
and U7279 (N_7279,N_1104,N_1617);
and U7280 (N_7280,N_4285,N_4235);
and U7281 (N_7281,N_3051,N_4279);
or U7282 (N_7282,N_614,N_251);
nor U7283 (N_7283,N_1258,N_2242);
xor U7284 (N_7284,N_2409,N_1802);
nor U7285 (N_7285,N_3754,N_1472);
or U7286 (N_7286,N_675,N_178);
or U7287 (N_7287,N_4937,N_4742);
and U7288 (N_7288,N_131,N_1430);
and U7289 (N_7289,N_2669,N_4344);
nor U7290 (N_7290,N_3,N_3978);
or U7291 (N_7291,N_3243,N_4483);
nand U7292 (N_7292,N_1768,N_3660);
and U7293 (N_7293,N_1493,N_1397);
and U7294 (N_7294,N_3816,N_4425);
or U7295 (N_7295,N_1236,N_3117);
or U7296 (N_7296,N_4298,N_1558);
xnor U7297 (N_7297,N_1829,N_3335);
or U7298 (N_7298,N_1067,N_1265);
xnor U7299 (N_7299,N_3933,N_1318);
xnor U7300 (N_7300,N_4440,N_1392);
nor U7301 (N_7301,N_474,N_3158);
nand U7302 (N_7302,N_4514,N_3394);
xnor U7303 (N_7303,N_2487,N_2859);
nor U7304 (N_7304,N_1893,N_839);
nor U7305 (N_7305,N_3196,N_2147);
xnor U7306 (N_7306,N_1014,N_2633);
or U7307 (N_7307,N_4210,N_3749);
or U7308 (N_7308,N_4659,N_4329);
and U7309 (N_7309,N_478,N_3362);
and U7310 (N_7310,N_355,N_401);
xor U7311 (N_7311,N_1436,N_4111);
nand U7312 (N_7312,N_2327,N_428);
or U7313 (N_7313,N_457,N_1361);
or U7314 (N_7314,N_399,N_2585);
nand U7315 (N_7315,N_1625,N_3852);
nor U7316 (N_7316,N_3523,N_3980);
or U7317 (N_7317,N_3088,N_4182);
or U7318 (N_7318,N_151,N_1443);
and U7319 (N_7319,N_1786,N_3595);
nor U7320 (N_7320,N_1811,N_1549);
xnor U7321 (N_7321,N_3908,N_2321);
and U7322 (N_7322,N_3068,N_1490);
nor U7323 (N_7323,N_487,N_931);
xor U7324 (N_7324,N_4166,N_502);
nor U7325 (N_7325,N_1465,N_2425);
and U7326 (N_7326,N_2042,N_4957);
or U7327 (N_7327,N_244,N_3375);
nor U7328 (N_7328,N_3385,N_3063);
and U7329 (N_7329,N_2279,N_2116);
nand U7330 (N_7330,N_2746,N_3052);
nor U7331 (N_7331,N_25,N_1965);
xnor U7332 (N_7332,N_3737,N_3323);
nand U7333 (N_7333,N_2078,N_4826);
or U7334 (N_7334,N_1423,N_93);
nand U7335 (N_7335,N_4305,N_2765);
nand U7336 (N_7336,N_4699,N_2066);
nand U7337 (N_7337,N_562,N_2355);
nor U7338 (N_7338,N_4192,N_821);
and U7339 (N_7339,N_2473,N_491);
nor U7340 (N_7340,N_130,N_3735);
and U7341 (N_7341,N_37,N_2020);
and U7342 (N_7342,N_216,N_2464);
and U7343 (N_7343,N_1808,N_205);
nor U7344 (N_7344,N_2213,N_4586);
or U7345 (N_7345,N_4115,N_3355);
and U7346 (N_7346,N_2838,N_2819);
nor U7347 (N_7347,N_4031,N_2646);
or U7348 (N_7348,N_4065,N_4780);
and U7349 (N_7349,N_4532,N_434);
or U7350 (N_7350,N_3011,N_3670);
nand U7351 (N_7351,N_1543,N_4271);
and U7352 (N_7352,N_4880,N_4126);
or U7353 (N_7353,N_2605,N_3218);
or U7354 (N_7354,N_4723,N_90);
xor U7355 (N_7355,N_1810,N_2306);
xnor U7356 (N_7356,N_4328,N_1912);
and U7357 (N_7357,N_4885,N_4673);
xor U7358 (N_7358,N_3236,N_2148);
nand U7359 (N_7359,N_1593,N_4856);
and U7360 (N_7360,N_2769,N_3522);
xnor U7361 (N_7361,N_4195,N_2707);
nand U7362 (N_7362,N_4574,N_1514);
and U7363 (N_7363,N_4894,N_4133);
and U7364 (N_7364,N_520,N_3634);
nor U7365 (N_7365,N_2139,N_4087);
or U7366 (N_7366,N_3464,N_4958);
and U7367 (N_7367,N_3061,N_3532);
xor U7368 (N_7368,N_3984,N_3159);
or U7369 (N_7369,N_3105,N_3407);
nor U7370 (N_7370,N_1953,N_2557);
and U7371 (N_7371,N_3772,N_2466);
and U7372 (N_7372,N_3248,N_793);
nand U7373 (N_7373,N_3802,N_4755);
nand U7374 (N_7374,N_1310,N_1512);
and U7375 (N_7375,N_3283,N_3081);
nand U7376 (N_7376,N_3914,N_4129);
and U7377 (N_7377,N_2165,N_2684);
and U7378 (N_7378,N_3836,N_2025);
nand U7379 (N_7379,N_1127,N_111);
xor U7380 (N_7380,N_2337,N_735);
and U7381 (N_7381,N_4169,N_4955);
or U7382 (N_7382,N_2505,N_2121);
nand U7383 (N_7383,N_1277,N_1790);
nand U7384 (N_7384,N_4183,N_2081);
nand U7385 (N_7385,N_2244,N_650);
nand U7386 (N_7386,N_2683,N_1577);
and U7387 (N_7387,N_4738,N_2311);
nor U7388 (N_7388,N_3693,N_1330);
and U7389 (N_7389,N_4361,N_2817);
xor U7390 (N_7390,N_1404,N_1742);
and U7391 (N_7391,N_2188,N_4207);
and U7392 (N_7392,N_2797,N_200);
xnor U7393 (N_7393,N_1935,N_4890);
nor U7394 (N_7394,N_4189,N_2210);
or U7395 (N_7395,N_4467,N_725);
nor U7396 (N_7396,N_612,N_2834);
and U7397 (N_7397,N_3489,N_752);
xnor U7398 (N_7398,N_238,N_2537);
nand U7399 (N_7399,N_4113,N_3640);
nand U7400 (N_7400,N_3499,N_4167);
and U7401 (N_7401,N_2860,N_3930);
xor U7402 (N_7402,N_4640,N_3529);
xnor U7403 (N_7403,N_1868,N_423);
nor U7404 (N_7404,N_3814,N_1576);
nand U7405 (N_7405,N_413,N_4524);
and U7406 (N_7406,N_4588,N_2168);
xnor U7407 (N_7407,N_3680,N_686);
or U7408 (N_7408,N_3803,N_3285);
xnor U7409 (N_7409,N_967,N_309);
or U7410 (N_7410,N_322,N_3200);
nand U7411 (N_7411,N_1019,N_1684);
and U7412 (N_7412,N_1529,N_621);
or U7413 (N_7413,N_217,N_1586);
xnor U7414 (N_7414,N_3627,N_2292);
or U7415 (N_7415,N_13,N_186);
nand U7416 (N_7416,N_2897,N_916);
or U7417 (N_7417,N_904,N_1670);
xor U7418 (N_7418,N_4412,N_4722);
or U7419 (N_7419,N_2992,N_1797);
or U7420 (N_7420,N_4473,N_1290);
nand U7421 (N_7421,N_2144,N_295);
nor U7422 (N_7422,N_1884,N_2075);
and U7423 (N_7423,N_2294,N_351);
nand U7424 (N_7424,N_1245,N_1675);
nand U7425 (N_7425,N_2199,N_4469);
nor U7426 (N_7426,N_510,N_2814);
or U7427 (N_7427,N_2788,N_2544);
and U7428 (N_7428,N_2710,N_1296);
xnor U7429 (N_7429,N_3541,N_3164);
and U7430 (N_7430,N_1701,N_4512);
nand U7431 (N_7431,N_2091,N_1926);
or U7432 (N_7432,N_1485,N_3962);
and U7433 (N_7433,N_184,N_2898);
nand U7434 (N_7434,N_45,N_3365);
or U7435 (N_7435,N_1101,N_1110);
or U7436 (N_7436,N_3563,N_4339);
nand U7437 (N_7437,N_2037,N_897);
xor U7438 (N_7438,N_3699,N_2018);
and U7439 (N_7439,N_4930,N_3427);
and U7440 (N_7440,N_2988,N_2695);
or U7441 (N_7441,N_3534,N_69);
nand U7442 (N_7442,N_2777,N_4528);
xor U7443 (N_7443,N_221,N_4431);
nand U7444 (N_7444,N_1391,N_1042);
nor U7445 (N_7445,N_3765,N_1181);
nand U7446 (N_7446,N_1090,N_4902);
xnor U7447 (N_7447,N_812,N_3560);
nor U7448 (N_7448,N_2087,N_1762);
and U7449 (N_7449,N_3587,N_4907);
and U7450 (N_7450,N_3956,N_1885);
nand U7451 (N_7451,N_118,N_1196);
nand U7452 (N_7452,N_2999,N_1402);
and U7453 (N_7453,N_273,N_2558);
and U7454 (N_7454,N_3317,N_3131);
or U7455 (N_7455,N_3400,N_4481);
and U7456 (N_7456,N_996,N_4879);
nor U7457 (N_7457,N_60,N_1174);
nor U7458 (N_7458,N_1817,N_2622);
nand U7459 (N_7459,N_4795,N_921);
nand U7460 (N_7460,N_2302,N_1032);
xor U7461 (N_7461,N_980,N_3095);
nor U7462 (N_7462,N_1049,N_4347);
nand U7463 (N_7463,N_531,N_2097);
nand U7464 (N_7464,N_1646,N_65);
nor U7465 (N_7465,N_3466,N_538);
nor U7466 (N_7466,N_4445,N_685);
and U7467 (N_7467,N_4997,N_2322);
xor U7468 (N_7468,N_48,N_2392);
or U7469 (N_7469,N_1888,N_3559);
nand U7470 (N_7470,N_3661,N_311);
and U7471 (N_7471,N_3839,N_887);
xnor U7472 (N_7472,N_264,N_2205);
nand U7473 (N_7473,N_1217,N_3086);
xnor U7474 (N_7474,N_1710,N_3650);
and U7475 (N_7475,N_145,N_1853);
and U7476 (N_7476,N_4891,N_2124);
and U7477 (N_7477,N_305,N_1170);
nor U7478 (N_7478,N_3686,N_3924);
nand U7479 (N_7479,N_3506,N_315);
or U7480 (N_7480,N_368,N_1481);
nand U7481 (N_7481,N_4270,N_3712);
and U7482 (N_7482,N_3681,N_2041);
and U7483 (N_7483,N_4020,N_2022);
nor U7484 (N_7484,N_1521,N_1875);
and U7485 (N_7485,N_4332,N_4463);
or U7486 (N_7486,N_1113,N_1852);
and U7487 (N_7487,N_1315,N_1403);
xor U7488 (N_7488,N_1681,N_479);
and U7489 (N_7489,N_4010,N_4221);
xnor U7490 (N_7490,N_638,N_4781);
nor U7491 (N_7491,N_511,N_4489);
xor U7492 (N_7492,N_4458,N_535);
nor U7493 (N_7493,N_3846,N_3605);
nand U7494 (N_7494,N_2440,N_3551);
nor U7495 (N_7495,N_3753,N_1328);
and U7496 (N_7496,N_2358,N_755);
xor U7497 (N_7497,N_3170,N_2671);
or U7498 (N_7498,N_2006,N_2660);
and U7499 (N_7499,N_3724,N_3328);
xor U7500 (N_7500,N_3165,N_4816);
xor U7501 (N_7501,N_1377,N_798);
nor U7502 (N_7502,N_1814,N_4864);
nor U7503 (N_7503,N_408,N_363);
or U7504 (N_7504,N_2689,N_4224);
or U7505 (N_7505,N_2117,N_1004);
and U7506 (N_7506,N_3586,N_4041);
and U7507 (N_7507,N_4178,N_907);
xnor U7508 (N_7508,N_2856,N_3500);
or U7509 (N_7509,N_751,N_1185);
or U7510 (N_7510,N_4098,N_195);
or U7511 (N_7511,N_1659,N_1860);
xor U7512 (N_7512,N_1349,N_1810);
nand U7513 (N_7513,N_48,N_2012);
and U7514 (N_7514,N_1623,N_4088);
nand U7515 (N_7515,N_3062,N_3224);
or U7516 (N_7516,N_4160,N_1276);
nand U7517 (N_7517,N_377,N_4256);
xor U7518 (N_7518,N_4029,N_4104);
or U7519 (N_7519,N_3325,N_3018);
or U7520 (N_7520,N_451,N_92);
and U7521 (N_7521,N_2758,N_1459);
xnor U7522 (N_7522,N_3458,N_744);
xnor U7523 (N_7523,N_450,N_323);
nor U7524 (N_7524,N_3401,N_850);
xnor U7525 (N_7525,N_2526,N_3777);
or U7526 (N_7526,N_4049,N_3370);
xor U7527 (N_7527,N_4337,N_4237);
xor U7528 (N_7528,N_1395,N_3035);
and U7529 (N_7529,N_1104,N_3922);
nor U7530 (N_7530,N_4855,N_579);
nand U7531 (N_7531,N_3500,N_3474);
nor U7532 (N_7532,N_2982,N_1294);
nand U7533 (N_7533,N_746,N_4384);
xor U7534 (N_7534,N_2898,N_2022);
nor U7535 (N_7535,N_2588,N_1952);
xor U7536 (N_7536,N_293,N_1318);
nand U7537 (N_7537,N_3424,N_4200);
nor U7538 (N_7538,N_1355,N_2923);
nand U7539 (N_7539,N_3892,N_3969);
xnor U7540 (N_7540,N_1126,N_134);
or U7541 (N_7541,N_3110,N_692);
xnor U7542 (N_7542,N_3445,N_293);
nor U7543 (N_7543,N_1760,N_3824);
and U7544 (N_7544,N_4444,N_277);
or U7545 (N_7545,N_1747,N_973);
and U7546 (N_7546,N_2185,N_2644);
nand U7547 (N_7547,N_56,N_3343);
nand U7548 (N_7548,N_4587,N_618);
nand U7549 (N_7549,N_1678,N_1936);
and U7550 (N_7550,N_785,N_937);
nor U7551 (N_7551,N_1364,N_4793);
and U7552 (N_7552,N_2809,N_3493);
nand U7553 (N_7553,N_160,N_1565);
or U7554 (N_7554,N_1021,N_134);
or U7555 (N_7555,N_508,N_2267);
or U7556 (N_7556,N_1926,N_3025);
and U7557 (N_7557,N_1461,N_3239);
or U7558 (N_7558,N_3484,N_3820);
nor U7559 (N_7559,N_3852,N_220);
nor U7560 (N_7560,N_4860,N_1546);
nor U7561 (N_7561,N_1998,N_4065);
nand U7562 (N_7562,N_4257,N_355);
nor U7563 (N_7563,N_1495,N_4869);
nand U7564 (N_7564,N_2560,N_4654);
xor U7565 (N_7565,N_4085,N_917);
or U7566 (N_7566,N_2050,N_2232);
or U7567 (N_7567,N_3479,N_2676);
and U7568 (N_7568,N_4019,N_1465);
or U7569 (N_7569,N_292,N_2637);
or U7570 (N_7570,N_3774,N_4138);
xor U7571 (N_7571,N_182,N_1175);
or U7572 (N_7572,N_4766,N_1450);
and U7573 (N_7573,N_2350,N_3784);
or U7574 (N_7574,N_723,N_2342);
or U7575 (N_7575,N_1260,N_3325);
nor U7576 (N_7576,N_1830,N_1017);
xor U7577 (N_7577,N_666,N_1093);
nor U7578 (N_7578,N_1047,N_4264);
nor U7579 (N_7579,N_454,N_260);
nand U7580 (N_7580,N_289,N_4670);
or U7581 (N_7581,N_1535,N_165);
or U7582 (N_7582,N_3950,N_3320);
nand U7583 (N_7583,N_4537,N_1782);
nor U7584 (N_7584,N_2047,N_528);
or U7585 (N_7585,N_35,N_3223);
and U7586 (N_7586,N_1585,N_2027);
nor U7587 (N_7587,N_2472,N_4916);
nor U7588 (N_7588,N_1983,N_3182);
or U7589 (N_7589,N_3816,N_2588);
nor U7590 (N_7590,N_1370,N_3609);
and U7591 (N_7591,N_2240,N_43);
nand U7592 (N_7592,N_4170,N_4186);
or U7593 (N_7593,N_1188,N_1292);
and U7594 (N_7594,N_1619,N_1128);
or U7595 (N_7595,N_3187,N_1877);
or U7596 (N_7596,N_3783,N_1752);
or U7597 (N_7597,N_181,N_490);
and U7598 (N_7598,N_3396,N_2622);
nand U7599 (N_7599,N_1974,N_1837);
and U7600 (N_7600,N_160,N_50);
xor U7601 (N_7601,N_4944,N_3159);
and U7602 (N_7602,N_1686,N_3388);
xnor U7603 (N_7603,N_622,N_4558);
xor U7604 (N_7604,N_1359,N_2758);
nand U7605 (N_7605,N_1265,N_162);
or U7606 (N_7606,N_4137,N_4975);
nor U7607 (N_7607,N_3662,N_3145);
nand U7608 (N_7608,N_399,N_3256);
nand U7609 (N_7609,N_4453,N_4346);
xor U7610 (N_7610,N_4978,N_1770);
or U7611 (N_7611,N_3469,N_3266);
xor U7612 (N_7612,N_2276,N_1076);
and U7613 (N_7613,N_1329,N_4718);
and U7614 (N_7614,N_483,N_2107);
nand U7615 (N_7615,N_4851,N_1851);
and U7616 (N_7616,N_3739,N_3507);
xnor U7617 (N_7617,N_1397,N_3676);
xnor U7618 (N_7618,N_1426,N_2474);
nor U7619 (N_7619,N_2846,N_4951);
nand U7620 (N_7620,N_708,N_1801);
or U7621 (N_7621,N_4903,N_894);
or U7622 (N_7622,N_3175,N_2641);
nor U7623 (N_7623,N_1321,N_1702);
or U7624 (N_7624,N_2887,N_2395);
nor U7625 (N_7625,N_3986,N_1035);
xnor U7626 (N_7626,N_715,N_3045);
xnor U7627 (N_7627,N_3385,N_922);
or U7628 (N_7628,N_3348,N_2515);
or U7629 (N_7629,N_3490,N_4732);
nor U7630 (N_7630,N_2798,N_2207);
nand U7631 (N_7631,N_4706,N_3275);
nor U7632 (N_7632,N_2149,N_1709);
xnor U7633 (N_7633,N_3817,N_4627);
nor U7634 (N_7634,N_739,N_488);
nand U7635 (N_7635,N_4158,N_3376);
nand U7636 (N_7636,N_1835,N_2216);
xor U7637 (N_7637,N_3685,N_4310);
nor U7638 (N_7638,N_3364,N_4412);
and U7639 (N_7639,N_3222,N_3092);
nand U7640 (N_7640,N_3091,N_3455);
or U7641 (N_7641,N_92,N_2865);
nand U7642 (N_7642,N_352,N_2901);
nand U7643 (N_7643,N_376,N_3959);
xnor U7644 (N_7644,N_1959,N_616);
xnor U7645 (N_7645,N_1442,N_4209);
and U7646 (N_7646,N_3432,N_4949);
xnor U7647 (N_7647,N_1409,N_1036);
nand U7648 (N_7648,N_4732,N_2839);
nand U7649 (N_7649,N_1314,N_1846);
nor U7650 (N_7650,N_1391,N_4656);
nand U7651 (N_7651,N_4656,N_759);
or U7652 (N_7652,N_3700,N_2879);
or U7653 (N_7653,N_3760,N_1169);
nor U7654 (N_7654,N_3456,N_3799);
and U7655 (N_7655,N_1638,N_4338);
nand U7656 (N_7656,N_4571,N_1155);
nor U7657 (N_7657,N_2232,N_1371);
nor U7658 (N_7658,N_3256,N_1357);
nand U7659 (N_7659,N_2856,N_862);
or U7660 (N_7660,N_2944,N_4212);
xor U7661 (N_7661,N_4704,N_1933);
xnor U7662 (N_7662,N_4037,N_2141);
or U7663 (N_7663,N_2940,N_4844);
or U7664 (N_7664,N_1847,N_3776);
and U7665 (N_7665,N_863,N_910);
and U7666 (N_7666,N_297,N_1102);
or U7667 (N_7667,N_4863,N_2690);
nor U7668 (N_7668,N_1174,N_247);
nand U7669 (N_7669,N_1017,N_3286);
and U7670 (N_7670,N_168,N_2100);
xor U7671 (N_7671,N_4877,N_3303);
nor U7672 (N_7672,N_910,N_3440);
or U7673 (N_7673,N_2509,N_4354);
nor U7674 (N_7674,N_4802,N_308);
nand U7675 (N_7675,N_1235,N_3132);
and U7676 (N_7676,N_3498,N_3122);
xor U7677 (N_7677,N_303,N_876);
nor U7678 (N_7678,N_1122,N_586);
and U7679 (N_7679,N_894,N_4693);
xnor U7680 (N_7680,N_4908,N_4366);
xor U7681 (N_7681,N_73,N_2304);
and U7682 (N_7682,N_4262,N_4064);
nand U7683 (N_7683,N_2558,N_1050);
xor U7684 (N_7684,N_87,N_1643);
xor U7685 (N_7685,N_1647,N_1049);
nand U7686 (N_7686,N_1308,N_3788);
nor U7687 (N_7687,N_2976,N_4007);
nor U7688 (N_7688,N_3032,N_4842);
nand U7689 (N_7689,N_3580,N_3367);
or U7690 (N_7690,N_3886,N_3524);
or U7691 (N_7691,N_4339,N_769);
or U7692 (N_7692,N_1118,N_2314);
or U7693 (N_7693,N_2762,N_2473);
or U7694 (N_7694,N_2335,N_4826);
xnor U7695 (N_7695,N_2731,N_2999);
xnor U7696 (N_7696,N_4252,N_2891);
xnor U7697 (N_7697,N_4896,N_2400);
or U7698 (N_7698,N_4229,N_3161);
nand U7699 (N_7699,N_2297,N_1899);
xor U7700 (N_7700,N_3006,N_1299);
and U7701 (N_7701,N_396,N_4574);
xnor U7702 (N_7702,N_4768,N_3178);
nand U7703 (N_7703,N_4218,N_129);
or U7704 (N_7704,N_3602,N_631);
and U7705 (N_7705,N_676,N_578);
and U7706 (N_7706,N_2599,N_2295);
nand U7707 (N_7707,N_4423,N_1101);
xnor U7708 (N_7708,N_2878,N_3591);
nand U7709 (N_7709,N_4507,N_1826);
nor U7710 (N_7710,N_2428,N_4056);
nand U7711 (N_7711,N_2869,N_203);
or U7712 (N_7712,N_2119,N_922);
and U7713 (N_7713,N_4256,N_1425);
nand U7714 (N_7714,N_2656,N_2285);
and U7715 (N_7715,N_2934,N_1278);
nor U7716 (N_7716,N_83,N_3772);
and U7717 (N_7717,N_4757,N_327);
and U7718 (N_7718,N_2749,N_3726);
nor U7719 (N_7719,N_583,N_369);
nor U7720 (N_7720,N_3651,N_3834);
nand U7721 (N_7721,N_2005,N_3729);
nor U7722 (N_7722,N_4526,N_4973);
or U7723 (N_7723,N_75,N_1687);
and U7724 (N_7724,N_2469,N_1611);
nor U7725 (N_7725,N_3753,N_2480);
xnor U7726 (N_7726,N_4222,N_872);
and U7727 (N_7727,N_1306,N_2403);
and U7728 (N_7728,N_3114,N_1779);
nor U7729 (N_7729,N_4448,N_944);
nor U7730 (N_7730,N_3760,N_3921);
xor U7731 (N_7731,N_2488,N_1474);
or U7732 (N_7732,N_1678,N_3578);
nor U7733 (N_7733,N_4201,N_2868);
and U7734 (N_7734,N_2636,N_791);
nand U7735 (N_7735,N_2616,N_919);
and U7736 (N_7736,N_3873,N_3994);
or U7737 (N_7737,N_3292,N_1461);
nor U7738 (N_7738,N_1670,N_119);
and U7739 (N_7739,N_812,N_4576);
xnor U7740 (N_7740,N_3169,N_4921);
xor U7741 (N_7741,N_1564,N_3608);
nor U7742 (N_7742,N_202,N_2357);
xor U7743 (N_7743,N_1012,N_338);
nor U7744 (N_7744,N_3752,N_1513);
nand U7745 (N_7745,N_986,N_1551);
nor U7746 (N_7746,N_519,N_1978);
or U7747 (N_7747,N_3407,N_920);
and U7748 (N_7748,N_3154,N_850);
and U7749 (N_7749,N_1951,N_800);
or U7750 (N_7750,N_685,N_3516);
xor U7751 (N_7751,N_2550,N_338);
and U7752 (N_7752,N_4944,N_1312);
nand U7753 (N_7753,N_1701,N_1065);
nand U7754 (N_7754,N_4079,N_4508);
nand U7755 (N_7755,N_2214,N_12);
nor U7756 (N_7756,N_3082,N_3066);
or U7757 (N_7757,N_3810,N_2317);
xnor U7758 (N_7758,N_4168,N_1232);
and U7759 (N_7759,N_1985,N_1062);
nor U7760 (N_7760,N_2678,N_991);
xnor U7761 (N_7761,N_4905,N_1855);
nor U7762 (N_7762,N_1991,N_2931);
nor U7763 (N_7763,N_1413,N_2383);
xnor U7764 (N_7764,N_4658,N_61);
xnor U7765 (N_7765,N_527,N_746);
nor U7766 (N_7766,N_2793,N_3555);
nand U7767 (N_7767,N_1961,N_2233);
nand U7768 (N_7768,N_4946,N_506);
nor U7769 (N_7769,N_1002,N_3156);
nor U7770 (N_7770,N_4467,N_2758);
nor U7771 (N_7771,N_3291,N_4846);
nand U7772 (N_7772,N_1370,N_3378);
nand U7773 (N_7773,N_1152,N_3125);
xnor U7774 (N_7774,N_2855,N_3912);
and U7775 (N_7775,N_353,N_2350);
or U7776 (N_7776,N_1506,N_644);
nor U7777 (N_7777,N_1485,N_3885);
xnor U7778 (N_7778,N_230,N_2633);
xnor U7779 (N_7779,N_1619,N_2112);
nor U7780 (N_7780,N_4857,N_842);
nand U7781 (N_7781,N_4823,N_2909);
or U7782 (N_7782,N_3263,N_2511);
nor U7783 (N_7783,N_3032,N_620);
nand U7784 (N_7784,N_4727,N_2532);
and U7785 (N_7785,N_676,N_718);
or U7786 (N_7786,N_4880,N_2654);
nand U7787 (N_7787,N_4711,N_3222);
nand U7788 (N_7788,N_2222,N_4700);
nor U7789 (N_7789,N_2691,N_1371);
xnor U7790 (N_7790,N_4156,N_3325);
or U7791 (N_7791,N_3293,N_4128);
xor U7792 (N_7792,N_1379,N_4586);
xnor U7793 (N_7793,N_44,N_2134);
nand U7794 (N_7794,N_3201,N_3447);
nor U7795 (N_7795,N_622,N_3683);
and U7796 (N_7796,N_4956,N_4597);
nor U7797 (N_7797,N_4007,N_2901);
and U7798 (N_7798,N_378,N_2463);
xnor U7799 (N_7799,N_2004,N_2254);
and U7800 (N_7800,N_1586,N_3051);
or U7801 (N_7801,N_1305,N_1482);
xor U7802 (N_7802,N_4303,N_1390);
nand U7803 (N_7803,N_1041,N_568);
xor U7804 (N_7804,N_1644,N_1242);
and U7805 (N_7805,N_4381,N_4145);
or U7806 (N_7806,N_664,N_862);
xnor U7807 (N_7807,N_3011,N_609);
nand U7808 (N_7808,N_4815,N_3590);
and U7809 (N_7809,N_1707,N_67);
nand U7810 (N_7810,N_1825,N_2718);
xnor U7811 (N_7811,N_4334,N_4495);
nand U7812 (N_7812,N_2327,N_1850);
or U7813 (N_7813,N_3030,N_4387);
nor U7814 (N_7814,N_4267,N_3580);
xor U7815 (N_7815,N_1471,N_2549);
xnor U7816 (N_7816,N_4095,N_4182);
nand U7817 (N_7817,N_1905,N_1151);
xnor U7818 (N_7818,N_463,N_4542);
nor U7819 (N_7819,N_3872,N_2664);
or U7820 (N_7820,N_3253,N_1670);
nor U7821 (N_7821,N_4040,N_3219);
and U7822 (N_7822,N_3329,N_548);
and U7823 (N_7823,N_3005,N_1578);
nand U7824 (N_7824,N_4340,N_4017);
or U7825 (N_7825,N_4141,N_2739);
nand U7826 (N_7826,N_2002,N_76);
xnor U7827 (N_7827,N_1066,N_269);
or U7828 (N_7828,N_3910,N_2798);
or U7829 (N_7829,N_3795,N_683);
or U7830 (N_7830,N_1289,N_644);
xnor U7831 (N_7831,N_2130,N_4328);
nand U7832 (N_7832,N_4760,N_2149);
nor U7833 (N_7833,N_495,N_1402);
nor U7834 (N_7834,N_3705,N_1937);
and U7835 (N_7835,N_3652,N_3993);
xor U7836 (N_7836,N_4366,N_560);
and U7837 (N_7837,N_3123,N_285);
nand U7838 (N_7838,N_1614,N_328);
xnor U7839 (N_7839,N_4760,N_4157);
or U7840 (N_7840,N_1763,N_3396);
xnor U7841 (N_7841,N_76,N_4925);
nand U7842 (N_7842,N_1971,N_3199);
nand U7843 (N_7843,N_3274,N_1941);
nor U7844 (N_7844,N_3667,N_4535);
and U7845 (N_7845,N_1929,N_195);
and U7846 (N_7846,N_3412,N_3404);
nor U7847 (N_7847,N_4426,N_3116);
nor U7848 (N_7848,N_1519,N_4199);
or U7849 (N_7849,N_4627,N_3886);
nor U7850 (N_7850,N_584,N_1244);
xor U7851 (N_7851,N_3468,N_1509);
nand U7852 (N_7852,N_3959,N_4295);
or U7853 (N_7853,N_609,N_3118);
nand U7854 (N_7854,N_882,N_2163);
or U7855 (N_7855,N_2276,N_3408);
xnor U7856 (N_7856,N_3263,N_1283);
nor U7857 (N_7857,N_1944,N_2633);
nand U7858 (N_7858,N_128,N_2425);
nor U7859 (N_7859,N_1489,N_3714);
nand U7860 (N_7860,N_2467,N_624);
or U7861 (N_7861,N_3318,N_1108);
and U7862 (N_7862,N_4684,N_1735);
nor U7863 (N_7863,N_1930,N_2233);
nor U7864 (N_7864,N_2107,N_2786);
nor U7865 (N_7865,N_1691,N_1270);
nor U7866 (N_7866,N_3614,N_4639);
or U7867 (N_7867,N_3057,N_1160);
and U7868 (N_7868,N_4859,N_1677);
nand U7869 (N_7869,N_1722,N_2563);
nand U7870 (N_7870,N_1178,N_3384);
or U7871 (N_7871,N_2243,N_1416);
or U7872 (N_7872,N_3572,N_3224);
nor U7873 (N_7873,N_4576,N_1096);
and U7874 (N_7874,N_2201,N_314);
nor U7875 (N_7875,N_1758,N_1078);
or U7876 (N_7876,N_1009,N_383);
nor U7877 (N_7877,N_2414,N_4948);
or U7878 (N_7878,N_1615,N_2639);
or U7879 (N_7879,N_3488,N_227);
xor U7880 (N_7880,N_3034,N_742);
xnor U7881 (N_7881,N_2791,N_1846);
or U7882 (N_7882,N_754,N_2916);
xnor U7883 (N_7883,N_2938,N_3279);
or U7884 (N_7884,N_3250,N_1466);
xnor U7885 (N_7885,N_3875,N_4118);
nor U7886 (N_7886,N_2914,N_1534);
nand U7887 (N_7887,N_3047,N_1527);
nand U7888 (N_7888,N_3527,N_1788);
nand U7889 (N_7889,N_4879,N_3834);
xor U7890 (N_7890,N_3077,N_924);
nor U7891 (N_7891,N_3998,N_2734);
and U7892 (N_7892,N_1345,N_566);
or U7893 (N_7893,N_855,N_1633);
nand U7894 (N_7894,N_253,N_2620);
or U7895 (N_7895,N_3187,N_158);
and U7896 (N_7896,N_4554,N_3974);
and U7897 (N_7897,N_1220,N_3306);
nand U7898 (N_7898,N_4743,N_3923);
or U7899 (N_7899,N_3426,N_2157);
and U7900 (N_7900,N_4159,N_487);
or U7901 (N_7901,N_4786,N_4899);
and U7902 (N_7902,N_2642,N_671);
or U7903 (N_7903,N_3536,N_4036);
nand U7904 (N_7904,N_281,N_1246);
nor U7905 (N_7905,N_4930,N_2505);
nand U7906 (N_7906,N_3894,N_2752);
xor U7907 (N_7907,N_4859,N_1685);
xnor U7908 (N_7908,N_229,N_1268);
or U7909 (N_7909,N_2333,N_2428);
or U7910 (N_7910,N_2354,N_4804);
nand U7911 (N_7911,N_525,N_376);
or U7912 (N_7912,N_4182,N_857);
xor U7913 (N_7913,N_1257,N_1093);
nor U7914 (N_7914,N_882,N_2373);
nand U7915 (N_7915,N_3121,N_1389);
nor U7916 (N_7916,N_1189,N_2013);
nand U7917 (N_7917,N_2778,N_1782);
xnor U7918 (N_7918,N_2989,N_4098);
nor U7919 (N_7919,N_2098,N_2207);
nor U7920 (N_7920,N_2277,N_2031);
or U7921 (N_7921,N_2511,N_4093);
nand U7922 (N_7922,N_3662,N_2349);
nand U7923 (N_7923,N_1102,N_1976);
xor U7924 (N_7924,N_1377,N_298);
or U7925 (N_7925,N_4758,N_4187);
xnor U7926 (N_7926,N_4888,N_3310);
nand U7927 (N_7927,N_4267,N_3469);
nand U7928 (N_7928,N_1125,N_2423);
nand U7929 (N_7929,N_186,N_3123);
nand U7930 (N_7930,N_2986,N_465);
xor U7931 (N_7931,N_1049,N_3346);
and U7932 (N_7932,N_4665,N_2730);
xnor U7933 (N_7933,N_66,N_1847);
nand U7934 (N_7934,N_385,N_2613);
xor U7935 (N_7935,N_3379,N_638);
nor U7936 (N_7936,N_2526,N_4086);
or U7937 (N_7937,N_741,N_1981);
and U7938 (N_7938,N_4504,N_3195);
and U7939 (N_7939,N_68,N_2546);
nand U7940 (N_7940,N_2639,N_1960);
nand U7941 (N_7941,N_2097,N_2450);
xnor U7942 (N_7942,N_2752,N_3961);
nand U7943 (N_7943,N_2269,N_968);
nand U7944 (N_7944,N_4839,N_3440);
nand U7945 (N_7945,N_704,N_3612);
xnor U7946 (N_7946,N_2863,N_1287);
or U7947 (N_7947,N_3929,N_1984);
nand U7948 (N_7948,N_967,N_4675);
xnor U7949 (N_7949,N_955,N_4484);
nand U7950 (N_7950,N_3980,N_4074);
nor U7951 (N_7951,N_1646,N_3877);
nor U7952 (N_7952,N_4284,N_382);
nor U7953 (N_7953,N_541,N_4275);
nor U7954 (N_7954,N_2996,N_4082);
or U7955 (N_7955,N_4809,N_1245);
nor U7956 (N_7956,N_2981,N_2387);
and U7957 (N_7957,N_3058,N_4645);
nor U7958 (N_7958,N_815,N_3240);
and U7959 (N_7959,N_4795,N_2175);
nor U7960 (N_7960,N_2059,N_2646);
nand U7961 (N_7961,N_1793,N_3914);
nor U7962 (N_7962,N_1586,N_3999);
nor U7963 (N_7963,N_4098,N_3383);
or U7964 (N_7964,N_2705,N_1465);
and U7965 (N_7965,N_1806,N_1499);
or U7966 (N_7966,N_2544,N_2859);
or U7967 (N_7967,N_4051,N_591);
and U7968 (N_7968,N_1234,N_3928);
and U7969 (N_7969,N_1197,N_4707);
xor U7970 (N_7970,N_3585,N_4104);
nand U7971 (N_7971,N_3833,N_768);
or U7972 (N_7972,N_250,N_2977);
xor U7973 (N_7973,N_2450,N_2554);
or U7974 (N_7974,N_375,N_2540);
and U7975 (N_7975,N_3504,N_4082);
or U7976 (N_7976,N_4889,N_4152);
nand U7977 (N_7977,N_2281,N_431);
nor U7978 (N_7978,N_1382,N_3199);
xnor U7979 (N_7979,N_1944,N_979);
xnor U7980 (N_7980,N_682,N_2258);
nand U7981 (N_7981,N_199,N_3153);
nand U7982 (N_7982,N_4341,N_940);
or U7983 (N_7983,N_2602,N_1596);
xnor U7984 (N_7984,N_152,N_270);
xor U7985 (N_7985,N_402,N_116);
and U7986 (N_7986,N_1871,N_4181);
xor U7987 (N_7987,N_1972,N_3215);
and U7988 (N_7988,N_4748,N_4527);
nand U7989 (N_7989,N_1027,N_3224);
nand U7990 (N_7990,N_1135,N_1424);
and U7991 (N_7991,N_3465,N_605);
xor U7992 (N_7992,N_2264,N_709);
and U7993 (N_7993,N_2734,N_3778);
nor U7994 (N_7994,N_593,N_715);
nand U7995 (N_7995,N_1769,N_441);
nor U7996 (N_7996,N_2778,N_3388);
nand U7997 (N_7997,N_2910,N_115);
or U7998 (N_7998,N_1769,N_4750);
xnor U7999 (N_7999,N_1758,N_2597);
or U8000 (N_8000,N_1442,N_2905);
nand U8001 (N_8001,N_2595,N_577);
nand U8002 (N_8002,N_1440,N_1096);
and U8003 (N_8003,N_3844,N_4190);
and U8004 (N_8004,N_1203,N_4625);
nor U8005 (N_8005,N_4938,N_2750);
xnor U8006 (N_8006,N_3764,N_1020);
nor U8007 (N_8007,N_3720,N_1207);
and U8008 (N_8008,N_1997,N_2896);
nand U8009 (N_8009,N_778,N_2521);
xnor U8010 (N_8010,N_2135,N_3003);
or U8011 (N_8011,N_1572,N_389);
or U8012 (N_8012,N_2274,N_166);
nand U8013 (N_8013,N_3764,N_462);
nand U8014 (N_8014,N_3407,N_2287);
or U8015 (N_8015,N_599,N_2007);
nand U8016 (N_8016,N_1255,N_2231);
nor U8017 (N_8017,N_1393,N_465);
or U8018 (N_8018,N_3716,N_4801);
and U8019 (N_8019,N_4641,N_4446);
xor U8020 (N_8020,N_592,N_3074);
and U8021 (N_8021,N_4332,N_3512);
nand U8022 (N_8022,N_4942,N_760);
nand U8023 (N_8023,N_3211,N_2279);
and U8024 (N_8024,N_3933,N_2321);
and U8025 (N_8025,N_1899,N_3450);
xor U8026 (N_8026,N_4734,N_722);
or U8027 (N_8027,N_1042,N_1424);
xnor U8028 (N_8028,N_4000,N_1278);
nor U8029 (N_8029,N_3188,N_4108);
and U8030 (N_8030,N_1277,N_1165);
nand U8031 (N_8031,N_4373,N_370);
and U8032 (N_8032,N_3018,N_3969);
and U8033 (N_8033,N_2715,N_1092);
nor U8034 (N_8034,N_36,N_4725);
nand U8035 (N_8035,N_1373,N_1117);
and U8036 (N_8036,N_2414,N_4118);
nand U8037 (N_8037,N_2180,N_2527);
nand U8038 (N_8038,N_1931,N_1590);
nor U8039 (N_8039,N_2989,N_3985);
or U8040 (N_8040,N_3099,N_3766);
or U8041 (N_8041,N_4890,N_1488);
or U8042 (N_8042,N_2648,N_1520);
nand U8043 (N_8043,N_3623,N_1379);
and U8044 (N_8044,N_4985,N_4624);
xor U8045 (N_8045,N_2120,N_1343);
and U8046 (N_8046,N_4793,N_1690);
or U8047 (N_8047,N_328,N_221);
or U8048 (N_8048,N_2510,N_3625);
nor U8049 (N_8049,N_3617,N_1310);
nor U8050 (N_8050,N_1066,N_408);
nand U8051 (N_8051,N_3116,N_722);
nand U8052 (N_8052,N_3762,N_4507);
nand U8053 (N_8053,N_388,N_4497);
and U8054 (N_8054,N_3684,N_1514);
or U8055 (N_8055,N_4204,N_4935);
xor U8056 (N_8056,N_2662,N_2086);
nand U8057 (N_8057,N_2801,N_1488);
nor U8058 (N_8058,N_3846,N_4409);
nor U8059 (N_8059,N_4445,N_2859);
nor U8060 (N_8060,N_3618,N_2276);
xor U8061 (N_8061,N_3943,N_2710);
or U8062 (N_8062,N_3967,N_2022);
nand U8063 (N_8063,N_4095,N_3717);
nor U8064 (N_8064,N_2575,N_2069);
and U8065 (N_8065,N_1705,N_4062);
and U8066 (N_8066,N_959,N_3951);
xnor U8067 (N_8067,N_422,N_1836);
xnor U8068 (N_8068,N_413,N_4457);
or U8069 (N_8069,N_1982,N_3982);
nand U8070 (N_8070,N_2354,N_699);
and U8071 (N_8071,N_4239,N_278);
and U8072 (N_8072,N_48,N_2621);
and U8073 (N_8073,N_1775,N_444);
or U8074 (N_8074,N_194,N_2854);
and U8075 (N_8075,N_1382,N_2911);
or U8076 (N_8076,N_4415,N_1152);
nand U8077 (N_8077,N_2814,N_4550);
or U8078 (N_8078,N_3521,N_4736);
nor U8079 (N_8079,N_4220,N_1426);
nor U8080 (N_8080,N_1170,N_3547);
nor U8081 (N_8081,N_54,N_1637);
nor U8082 (N_8082,N_2972,N_1732);
and U8083 (N_8083,N_727,N_3714);
nor U8084 (N_8084,N_239,N_3284);
or U8085 (N_8085,N_767,N_3787);
nand U8086 (N_8086,N_1631,N_538);
nand U8087 (N_8087,N_3861,N_3047);
xnor U8088 (N_8088,N_3816,N_3921);
and U8089 (N_8089,N_1107,N_1330);
xor U8090 (N_8090,N_1990,N_1124);
or U8091 (N_8091,N_388,N_1736);
nor U8092 (N_8092,N_2638,N_2366);
or U8093 (N_8093,N_909,N_3298);
and U8094 (N_8094,N_2123,N_952);
or U8095 (N_8095,N_1012,N_2644);
nor U8096 (N_8096,N_61,N_3122);
nand U8097 (N_8097,N_2409,N_1111);
xnor U8098 (N_8098,N_2977,N_152);
nor U8099 (N_8099,N_162,N_3925);
xnor U8100 (N_8100,N_1095,N_2202);
nor U8101 (N_8101,N_1289,N_4108);
nor U8102 (N_8102,N_4822,N_4198);
nand U8103 (N_8103,N_1770,N_242);
nor U8104 (N_8104,N_4573,N_980);
and U8105 (N_8105,N_3478,N_766);
and U8106 (N_8106,N_4795,N_132);
nor U8107 (N_8107,N_2545,N_3449);
nor U8108 (N_8108,N_4690,N_3368);
nor U8109 (N_8109,N_3628,N_2267);
or U8110 (N_8110,N_1277,N_2935);
nand U8111 (N_8111,N_4959,N_2453);
or U8112 (N_8112,N_3861,N_4740);
and U8113 (N_8113,N_3638,N_3671);
or U8114 (N_8114,N_4665,N_517);
and U8115 (N_8115,N_3180,N_678);
nand U8116 (N_8116,N_3097,N_624);
nand U8117 (N_8117,N_4656,N_547);
or U8118 (N_8118,N_2252,N_294);
xnor U8119 (N_8119,N_2802,N_1614);
nand U8120 (N_8120,N_974,N_125);
or U8121 (N_8121,N_3688,N_2699);
nor U8122 (N_8122,N_4735,N_3470);
nor U8123 (N_8123,N_1936,N_3701);
nand U8124 (N_8124,N_278,N_1212);
nor U8125 (N_8125,N_4431,N_1812);
and U8126 (N_8126,N_2455,N_2427);
xnor U8127 (N_8127,N_2101,N_1161);
or U8128 (N_8128,N_3156,N_2407);
or U8129 (N_8129,N_4413,N_3775);
nor U8130 (N_8130,N_102,N_4130);
and U8131 (N_8131,N_3212,N_1892);
and U8132 (N_8132,N_227,N_2326);
and U8133 (N_8133,N_1564,N_2971);
or U8134 (N_8134,N_2948,N_1026);
nor U8135 (N_8135,N_1959,N_59);
and U8136 (N_8136,N_4146,N_5);
and U8137 (N_8137,N_797,N_3133);
xnor U8138 (N_8138,N_2829,N_350);
nor U8139 (N_8139,N_1580,N_1355);
and U8140 (N_8140,N_4258,N_3323);
nor U8141 (N_8141,N_3801,N_4823);
and U8142 (N_8142,N_2861,N_3071);
nand U8143 (N_8143,N_641,N_854);
and U8144 (N_8144,N_3188,N_743);
or U8145 (N_8145,N_2556,N_1663);
or U8146 (N_8146,N_4397,N_2391);
nand U8147 (N_8147,N_412,N_1524);
nand U8148 (N_8148,N_1816,N_3353);
nor U8149 (N_8149,N_2331,N_3037);
and U8150 (N_8150,N_2837,N_941);
nor U8151 (N_8151,N_3531,N_1783);
or U8152 (N_8152,N_2407,N_2375);
or U8153 (N_8153,N_788,N_1349);
or U8154 (N_8154,N_989,N_4785);
or U8155 (N_8155,N_2343,N_3650);
nand U8156 (N_8156,N_1482,N_3528);
xnor U8157 (N_8157,N_2168,N_1525);
nor U8158 (N_8158,N_1559,N_3350);
nor U8159 (N_8159,N_2128,N_924);
or U8160 (N_8160,N_4662,N_2208);
or U8161 (N_8161,N_1694,N_820);
or U8162 (N_8162,N_4553,N_392);
nand U8163 (N_8163,N_2524,N_4423);
xnor U8164 (N_8164,N_3294,N_3164);
xor U8165 (N_8165,N_1856,N_1998);
and U8166 (N_8166,N_1938,N_501);
nor U8167 (N_8167,N_308,N_3165);
nand U8168 (N_8168,N_1094,N_2801);
xnor U8169 (N_8169,N_1129,N_2847);
or U8170 (N_8170,N_186,N_1792);
xor U8171 (N_8171,N_3234,N_3447);
xnor U8172 (N_8172,N_2107,N_401);
and U8173 (N_8173,N_4767,N_2855);
xor U8174 (N_8174,N_876,N_1616);
nand U8175 (N_8175,N_3332,N_4482);
and U8176 (N_8176,N_2057,N_634);
nor U8177 (N_8177,N_2692,N_4283);
or U8178 (N_8178,N_2996,N_1741);
nand U8179 (N_8179,N_1638,N_3294);
and U8180 (N_8180,N_1649,N_771);
nand U8181 (N_8181,N_4464,N_503);
nor U8182 (N_8182,N_2088,N_1159);
or U8183 (N_8183,N_3604,N_536);
nand U8184 (N_8184,N_2837,N_4661);
and U8185 (N_8185,N_311,N_2792);
or U8186 (N_8186,N_4594,N_3793);
and U8187 (N_8187,N_2582,N_780);
nand U8188 (N_8188,N_3332,N_3008);
and U8189 (N_8189,N_1309,N_2712);
xor U8190 (N_8190,N_4683,N_3627);
xnor U8191 (N_8191,N_4077,N_4335);
or U8192 (N_8192,N_2349,N_1252);
and U8193 (N_8193,N_750,N_147);
or U8194 (N_8194,N_2946,N_4042);
nand U8195 (N_8195,N_2619,N_3612);
and U8196 (N_8196,N_4008,N_2049);
xor U8197 (N_8197,N_4912,N_1307);
nor U8198 (N_8198,N_1527,N_3851);
and U8199 (N_8199,N_628,N_1952);
and U8200 (N_8200,N_2723,N_4899);
nor U8201 (N_8201,N_2631,N_1156);
or U8202 (N_8202,N_4062,N_2054);
nor U8203 (N_8203,N_691,N_1265);
xor U8204 (N_8204,N_1808,N_4181);
or U8205 (N_8205,N_2971,N_2826);
xor U8206 (N_8206,N_4033,N_3510);
xor U8207 (N_8207,N_4114,N_4358);
and U8208 (N_8208,N_2779,N_2212);
and U8209 (N_8209,N_2718,N_1667);
and U8210 (N_8210,N_1174,N_2191);
nand U8211 (N_8211,N_4493,N_2327);
nor U8212 (N_8212,N_4622,N_2084);
xnor U8213 (N_8213,N_1671,N_669);
nor U8214 (N_8214,N_2656,N_634);
nand U8215 (N_8215,N_2604,N_2687);
or U8216 (N_8216,N_1200,N_1134);
and U8217 (N_8217,N_3834,N_1195);
or U8218 (N_8218,N_923,N_752);
nor U8219 (N_8219,N_3758,N_4960);
xor U8220 (N_8220,N_3097,N_3370);
nand U8221 (N_8221,N_2874,N_361);
nor U8222 (N_8222,N_2366,N_1809);
or U8223 (N_8223,N_4290,N_679);
and U8224 (N_8224,N_796,N_4534);
and U8225 (N_8225,N_595,N_2889);
nor U8226 (N_8226,N_226,N_2240);
xnor U8227 (N_8227,N_1530,N_4029);
and U8228 (N_8228,N_625,N_4250);
and U8229 (N_8229,N_877,N_2832);
and U8230 (N_8230,N_2353,N_4742);
nor U8231 (N_8231,N_2462,N_81);
and U8232 (N_8232,N_4518,N_1739);
xnor U8233 (N_8233,N_524,N_4704);
nand U8234 (N_8234,N_3999,N_4578);
nand U8235 (N_8235,N_678,N_1604);
xnor U8236 (N_8236,N_1861,N_1676);
nor U8237 (N_8237,N_4236,N_699);
nand U8238 (N_8238,N_651,N_1379);
xor U8239 (N_8239,N_3765,N_3477);
or U8240 (N_8240,N_2425,N_3058);
nand U8241 (N_8241,N_1282,N_3805);
xnor U8242 (N_8242,N_130,N_590);
nand U8243 (N_8243,N_2601,N_3082);
xnor U8244 (N_8244,N_3470,N_2148);
or U8245 (N_8245,N_3814,N_2065);
nand U8246 (N_8246,N_2380,N_162);
and U8247 (N_8247,N_3742,N_652);
xor U8248 (N_8248,N_3475,N_3609);
xnor U8249 (N_8249,N_1256,N_1377);
or U8250 (N_8250,N_859,N_3846);
nand U8251 (N_8251,N_2990,N_4267);
xnor U8252 (N_8252,N_2444,N_2429);
or U8253 (N_8253,N_2213,N_4926);
and U8254 (N_8254,N_3395,N_28);
and U8255 (N_8255,N_2497,N_393);
or U8256 (N_8256,N_2227,N_2868);
or U8257 (N_8257,N_4718,N_1507);
or U8258 (N_8258,N_3512,N_1489);
nand U8259 (N_8259,N_4166,N_1849);
or U8260 (N_8260,N_2009,N_2117);
nor U8261 (N_8261,N_4113,N_1392);
xnor U8262 (N_8262,N_431,N_3642);
nand U8263 (N_8263,N_951,N_3065);
xnor U8264 (N_8264,N_3570,N_4526);
nand U8265 (N_8265,N_3185,N_244);
and U8266 (N_8266,N_1781,N_1149);
nand U8267 (N_8267,N_1509,N_685);
or U8268 (N_8268,N_686,N_4072);
nor U8269 (N_8269,N_1182,N_3562);
nor U8270 (N_8270,N_1680,N_3447);
or U8271 (N_8271,N_441,N_4601);
or U8272 (N_8272,N_4666,N_4872);
and U8273 (N_8273,N_2762,N_405);
or U8274 (N_8274,N_183,N_4168);
and U8275 (N_8275,N_4821,N_3482);
nor U8276 (N_8276,N_379,N_1977);
xnor U8277 (N_8277,N_3243,N_2099);
xor U8278 (N_8278,N_2148,N_425);
xnor U8279 (N_8279,N_1748,N_3058);
xor U8280 (N_8280,N_4139,N_3302);
nand U8281 (N_8281,N_768,N_2473);
or U8282 (N_8282,N_3669,N_4140);
or U8283 (N_8283,N_2378,N_762);
nand U8284 (N_8284,N_1280,N_1770);
nand U8285 (N_8285,N_4507,N_3161);
nand U8286 (N_8286,N_2832,N_2099);
and U8287 (N_8287,N_987,N_4786);
nand U8288 (N_8288,N_943,N_4357);
xnor U8289 (N_8289,N_1029,N_1261);
nor U8290 (N_8290,N_3588,N_4492);
nand U8291 (N_8291,N_3543,N_1465);
and U8292 (N_8292,N_4669,N_245);
nand U8293 (N_8293,N_2345,N_179);
xnor U8294 (N_8294,N_1539,N_4390);
or U8295 (N_8295,N_2137,N_2458);
xor U8296 (N_8296,N_2628,N_3567);
nand U8297 (N_8297,N_4584,N_2701);
nor U8298 (N_8298,N_2216,N_3678);
nor U8299 (N_8299,N_2315,N_3685);
xor U8300 (N_8300,N_4623,N_3611);
and U8301 (N_8301,N_4544,N_2574);
or U8302 (N_8302,N_2824,N_2646);
and U8303 (N_8303,N_3982,N_907);
nor U8304 (N_8304,N_553,N_27);
nor U8305 (N_8305,N_3884,N_2803);
nor U8306 (N_8306,N_3929,N_1028);
and U8307 (N_8307,N_877,N_1584);
and U8308 (N_8308,N_4374,N_444);
nor U8309 (N_8309,N_201,N_2129);
and U8310 (N_8310,N_4213,N_3638);
nand U8311 (N_8311,N_2527,N_3434);
and U8312 (N_8312,N_4329,N_922);
and U8313 (N_8313,N_2725,N_1477);
or U8314 (N_8314,N_3680,N_1383);
nor U8315 (N_8315,N_2983,N_773);
nor U8316 (N_8316,N_2446,N_3881);
nor U8317 (N_8317,N_2532,N_1939);
nand U8318 (N_8318,N_4385,N_4623);
and U8319 (N_8319,N_3529,N_1090);
xnor U8320 (N_8320,N_1518,N_2730);
nor U8321 (N_8321,N_526,N_150);
or U8322 (N_8322,N_3907,N_1249);
nor U8323 (N_8323,N_3089,N_371);
or U8324 (N_8324,N_1890,N_2196);
and U8325 (N_8325,N_2692,N_2158);
nor U8326 (N_8326,N_2810,N_2390);
nor U8327 (N_8327,N_340,N_3330);
nor U8328 (N_8328,N_846,N_4713);
xnor U8329 (N_8329,N_3573,N_661);
nand U8330 (N_8330,N_3633,N_3253);
nand U8331 (N_8331,N_4187,N_362);
and U8332 (N_8332,N_4701,N_2247);
or U8333 (N_8333,N_576,N_3560);
nor U8334 (N_8334,N_1478,N_1861);
and U8335 (N_8335,N_2433,N_2188);
nand U8336 (N_8336,N_2088,N_3785);
nor U8337 (N_8337,N_579,N_2604);
xnor U8338 (N_8338,N_105,N_2750);
nor U8339 (N_8339,N_3340,N_2934);
nor U8340 (N_8340,N_1976,N_395);
and U8341 (N_8341,N_359,N_4362);
nor U8342 (N_8342,N_4072,N_4244);
nor U8343 (N_8343,N_910,N_2114);
or U8344 (N_8344,N_1298,N_3375);
nor U8345 (N_8345,N_1857,N_1171);
nor U8346 (N_8346,N_2295,N_2377);
and U8347 (N_8347,N_416,N_4417);
nor U8348 (N_8348,N_554,N_4138);
or U8349 (N_8349,N_2274,N_4161);
and U8350 (N_8350,N_446,N_2371);
nand U8351 (N_8351,N_4450,N_4494);
or U8352 (N_8352,N_2526,N_2450);
nand U8353 (N_8353,N_391,N_4478);
xnor U8354 (N_8354,N_4818,N_1706);
xnor U8355 (N_8355,N_4144,N_3860);
xnor U8356 (N_8356,N_824,N_3378);
and U8357 (N_8357,N_2655,N_3248);
nand U8358 (N_8358,N_4668,N_3544);
nor U8359 (N_8359,N_1558,N_513);
or U8360 (N_8360,N_2385,N_1891);
or U8361 (N_8361,N_195,N_3138);
and U8362 (N_8362,N_1920,N_1812);
and U8363 (N_8363,N_2354,N_461);
and U8364 (N_8364,N_406,N_3289);
nor U8365 (N_8365,N_2031,N_3175);
xor U8366 (N_8366,N_2038,N_603);
nor U8367 (N_8367,N_1018,N_1597);
nor U8368 (N_8368,N_2191,N_1304);
nand U8369 (N_8369,N_2828,N_321);
nand U8370 (N_8370,N_1588,N_1459);
or U8371 (N_8371,N_687,N_3342);
xnor U8372 (N_8372,N_3546,N_4464);
nor U8373 (N_8373,N_4337,N_4541);
or U8374 (N_8374,N_3881,N_1503);
nand U8375 (N_8375,N_731,N_990);
nand U8376 (N_8376,N_4114,N_2114);
nor U8377 (N_8377,N_2625,N_1687);
and U8378 (N_8378,N_4319,N_4932);
or U8379 (N_8379,N_4230,N_321);
nor U8380 (N_8380,N_2559,N_4444);
nand U8381 (N_8381,N_1527,N_698);
nor U8382 (N_8382,N_1253,N_2000);
nor U8383 (N_8383,N_255,N_1997);
nor U8384 (N_8384,N_2063,N_3083);
and U8385 (N_8385,N_4710,N_1961);
xor U8386 (N_8386,N_4177,N_4122);
or U8387 (N_8387,N_796,N_4036);
or U8388 (N_8388,N_2758,N_213);
or U8389 (N_8389,N_4509,N_55);
and U8390 (N_8390,N_839,N_3082);
and U8391 (N_8391,N_1832,N_1480);
nor U8392 (N_8392,N_4613,N_886);
xor U8393 (N_8393,N_1415,N_4894);
xnor U8394 (N_8394,N_1908,N_3925);
or U8395 (N_8395,N_28,N_3152);
or U8396 (N_8396,N_2891,N_2028);
xor U8397 (N_8397,N_965,N_1429);
xor U8398 (N_8398,N_4311,N_322);
xnor U8399 (N_8399,N_4842,N_1736);
or U8400 (N_8400,N_1983,N_33);
or U8401 (N_8401,N_2829,N_1920);
nor U8402 (N_8402,N_2520,N_1026);
nand U8403 (N_8403,N_2576,N_3978);
and U8404 (N_8404,N_1545,N_3043);
and U8405 (N_8405,N_4235,N_3293);
or U8406 (N_8406,N_1920,N_3870);
nand U8407 (N_8407,N_1463,N_3617);
nor U8408 (N_8408,N_4747,N_994);
or U8409 (N_8409,N_3159,N_3632);
and U8410 (N_8410,N_4954,N_3449);
and U8411 (N_8411,N_4554,N_4549);
nor U8412 (N_8412,N_2890,N_4699);
or U8413 (N_8413,N_3648,N_1604);
nand U8414 (N_8414,N_3900,N_4318);
or U8415 (N_8415,N_1462,N_3031);
nand U8416 (N_8416,N_2604,N_2179);
or U8417 (N_8417,N_90,N_2622);
or U8418 (N_8418,N_1490,N_1205);
or U8419 (N_8419,N_4925,N_4886);
or U8420 (N_8420,N_3020,N_3745);
and U8421 (N_8421,N_1222,N_1421);
nand U8422 (N_8422,N_3480,N_2954);
nand U8423 (N_8423,N_2470,N_2345);
nand U8424 (N_8424,N_1466,N_2560);
nor U8425 (N_8425,N_3612,N_3267);
nor U8426 (N_8426,N_30,N_3199);
or U8427 (N_8427,N_3406,N_350);
nand U8428 (N_8428,N_4081,N_3598);
nand U8429 (N_8429,N_4125,N_1105);
nor U8430 (N_8430,N_1326,N_2974);
or U8431 (N_8431,N_1392,N_2183);
or U8432 (N_8432,N_4370,N_3068);
nand U8433 (N_8433,N_4239,N_2007);
xnor U8434 (N_8434,N_1461,N_2335);
nand U8435 (N_8435,N_4721,N_2952);
nand U8436 (N_8436,N_4601,N_3324);
nor U8437 (N_8437,N_1974,N_3756);
xor U8438 (N_8438,N_1510,N_836);
or U8439 (N_8439,N_819,N_701);
and U8440 (N_8440,N_1792,N_2317);
nor U8441 (N_8441,N_2626,N_4317);
nor U8442 (N_8442,N_2096,N_3284);
xnor U8443 (N_8443,N_995,N_2602);
or U8444 (N_8444,N_4720,N_214);
xor U8445 (N_8445,N_3260,N_452);
nand U8446 (N_8446,N_1706,N_3507);
and U8447 (N_8447,N_335,N_3554);
and U8448 (N_8448,N_3119,N_4289);
or U8449 (N_8449,N_3634,N_4260);
and U8450 (N_8450,N_4225,N_3046);
xnor U8451 (N_8451,N_4772,N_172);
and U8452 (N_8452,N_4221,N_4106);
or U8453 (N_8453,N_2378,N_2603);
or U8454 (N_8454,N_3952,N_3357);
or U8455 (N_8455,N_3784,N_3077);
xor U8456 (N_8456,N_4662,N_4355);
nor U8457 (N_8457,N_2231,N_1049);
xor U8458 (N_8458,N_2978,N_2060);
nor U8459 (N_8459,N_3466,N_4447);
xnor U8460 (N_8460,N_1444,N_2801);
and U8461 (N_8461,N_1593,N_3628);
or U8462 (N_8462,N_3184,N_3098);
nand U8463 (N_8463,N_3867,N_1610);
nand U8464 (N_8464,N_4346,N_4413);
and U8465 (N_8465,N_2368,N_4080);
and U8466 (N_8466,N_1908,N_4027);
xor U8467 (N_8467,N_1917,N_1360);
nand U8468 (N_8468,N_1749,N_4206);
nand U8469 (N_8469,N_2635,N_522);
nor U8470 (N_8470,N_763,N_3688);
and U8471 (N_8471,N_4683,N_2363);
xnor U8472 (N_8472,N_186,N_2128);
xnor U8473 (N_8473,N_1032,N_4776);
or U8474 (N_8474,N_723,N_3452);
or U8475 (N_8475,N_8,N_1242);
nand U8476 (N_8476,N_1176,N_4967);
nor U8477 (N_8477,N_3614,N_989);
and U8478 (N_8478,N_1943,N_1946);
nand U8479 (N_8479,N_3478,N_4358);
or U8480 (N_8480,N_2595,N_2596);
xnor U8481 (N_8481,N_4151,N_1326);
and U8482 (N_8482,N_712,N_4807);
xnor U8483 (N_8483,N_780,N_1197);
xnor U8484 (N_8484,N_2472,N_2328);
or U8485 (N_8485,N_4583,N_1468);
or U8486 (N_8486,N_4325,N_2714);
or U8487 (N_8487,N_1684,N_1941);
xor U8488 (N_8488,N_1743,N_702);
nor U8489 (N_8489,N_995,N_3550);
nand U8490 (N_8490,N_3699,N_4977);
and U8491 (N_8491,N_1070,N_2327);
xnor U8492 (N_8492,N_4854,N_469);
nor U8493 (N_8493,N_2312,N_3332);
nor U8494 (N_8494,N_710,N_752);
nor U8495 (N_8495,N_955,N_4970);
nor U8496 (N_8496,N_3613,N_3909);
xor U8497 (N_8497,N_3112,N_3914);
nand U8498 (N_8498,N_4242,N_1008);
or U8499 (N_8499,N_2487,N_969);
or U8500 (N_8500,N_791,N_3106);
nor U8501 (N_8501,N_3349,N_3779);
nor U8502 (N_8502,N_703,N_4255);
or U8503 (N_8503,N_2795,N_1261);
and U8504 (N_8504,N_87,N_1454);
nand U8505 (N_8505,N_1073,N_4623);
xor U8506 (N_8506,N_4225,N_487);
or U8507 (N_8507,N_4730,N_3444);
nand U8508 (N_8508,N_3696,N_3027);
xor U8509 (N_8509,N_363,N_4827);
nor U8510 (N_8510,N_4178,N_2881);
nor U8511 (N_8511,N_3555,N_218);
xnor U8512 (N_8512,N_4910,N_3487);
and U8513 (N_8513,N_4495,N_2435);
nor U8514 (N_8514,N_72,N_3405);
or U8515 (N_8515,N_379,N_640);
and U8516 (N_8516,N_438,N_211);
nor U8517 (N_8517,N_2795,N_4685);
nor U8518 (N_8518,N_2092,N_4778);
or U8519 (N_8519,N_4815,N_1150);
and U8520 (N_8520,N_2131,N_2178);
xnor U8521 (N_8521,N_2102,N_1370);
or U8522 (N_8522,N_4318,N_4827);
nor U8523 (N_8523,N_1049,N_1205);
nand U8524 (N_8524,N_3236,N_4309);
or U8525 (N_8525,N_3321,N_846);
nor U8526 (N_8526,N_4875,N_2423);
xor U8527 (N_8527,N_2160,N_2171);
nor U8528 (N_8528,N_424,N_4200);
or U8529 (N_8529,N_394,N_4743);
nand U8530 (N_8530,N_4410,N_4234);
nand U8531 (N_8531,N_410,N_2776);
nor U8532 (N_8532,N_1488,N_1521);
nand U8533 (N_8533,N_3732,N_3968);
nand U8534 (N_8534,N_233,N_954);
or U8535 (N_8535,N_2273,N_4936);
xnor U8536 (N_8536,N_1,N_726);
and U8537 (N_8537,N_1826,N_4780);
and U8538 (N_8538,N_2185,N_86);
or U8539 (N_8539,N_1338,N_2489);
and U8540 (N_8540,N_3433,N_4874);
and U8541 (N_8541,N_1350,N_2319);
nor U8542 (N_8542,N_2355,N_3217);
nor U8543 (N_8543,N_1490,N_1038);
nand U8544 (N_8544,N_4354,N_3441);
nor U8545 (N_8545,N_2394,N_4464);
nand U8546 (N_8546,N_402,N_4367);
xnor U8547 (N_8547,N_4510,N_51);
nand U8548 (N_8548,N_2382,N_1974);
xor U8549 (N_8549,N_3019,N_4839);
nand U8550 (N_8550,N_738,N_538);
or U8551 (N_8551,N_178,N_3666);
or U8552 (N_8552,N_1523,N_134);
nor U8553 (N_8553,N_3300,N_4144);
xor U8554 (N_8554,N_3326,N_4859);
and U8555 (N_8555,N_2561,N_2202);
xor U8556 (N_8556,N_4059,N_4409);
nor U8557 (N_8557,N_523,N_592);
nor U8558 (N_8558,N_617,N_1541);
xor U8559 (N_8559,N_542,N_1626);
or U8560 (N_8560,N_2143,N_2808);
nand U8561 (N_8561,N_399,N_4151);
or U8562 (N_8562,N_3514,N_684);
and U8563 (N_8563,N_2068,N_1821);
nand U8564 (N_8564,N_1983,N_1844);
and U8565 (N_8565,N_2260,N_2079);
xnor U8566 (N_8566,N_4946,N_4131);
and U8567 (N_8567,N_2160,N_1867);
nand U8568 (N_8568,N_4203,N_2591);
xnor U8569 (N_8569,N_3978,N_2919);
nor U8570 (N_8570,N_4543,N_2323);
nand U8571 (N_8571,N_3936,N_3579);
nand U8572 (N_8572,N_2097,N_3325);
or U8573 (N_8573,N_3220,N_3312);
and U8574 (N_8574,N_2985,N_856);
or U8575 (N_8575,N_4823,N_1010);
and U8576 (N_8576,N_2795,N_2013);
nor U8577 (N_8577,N_3209,N_3689);
nor U8578 (N_8578,N_880,N_4859);
or U8579 (N_8579,N_496,N_4063);
nand U8580 (N_8580,N_1204,N_2945);
and U8581 (N_8581,N_3010,N_1384);
or U8582 (N_8582,N_524,N_1633);
nand U8583 (N_8583,N_4320,N_3403);
nand U8584 (N_8584,N_4229,N_4464);
nor U8585 (N_8585,N_4221,N_2199);
nor U8586 (N_8586,N_2859,N_1514);
nor U8587 (N_8587,N_4545,N_842);
or U8588 (N_8588,N_457,N_2273);
nor U8589 (N_8589,N_3195,N_2946);
nand U8590 (N_8590,N_4063,N_4507);
or U8591 (N_8591,N_4354,N_1631);
nor U8592 (N_8592,N_1104,N_897);
or U8593 (N_8593,N_932,N_2113);
and U8594 (N_8594,N_3656,N_1745);
nor U8595 (N_8595,N_2584,N_2047);
and U8596 (N_8596,N_1764,N_233);
and U8597 (N_8597,N_3121,N_822);
and U8598 (N_8598,N_4790,N_875);
or U8599 (N_8599,N_4639,N_385);
nor U8600 (N_8600,N_1944,N_661);
nor U8601 (N_8601,N_1505,N_206);
nand U8602 (N_8602,N_782,N_1757);
or U8603 (N_8603,N_4622,N_4996);
xnor U8604 (N_8604,N_2910,N_752);
or U8605 (N_8605,N_4320,N_2296);
nor U8606 (N_8606,N_2961,N_3207);
xor U8607 (N_8607,N_3083,N_3080);
or U8608 (N_8608,N_1383,N_543);
or U8609 (N_8609,N_1742,N_4891);
xnor U8610 (N_8610,N_4384,N_3404);
or U8611 (N_8611,N_3915,N_3731);
xor U8612 (N_8612,N_1601,N_2538);
nor U8613 (N_8613,N_2532,N_2434);
or U8614 (N_8614,N_1430,N_4990);
or U8615 (N_8615,N_3830,N_1107);
nor U8616 (N_8616,N_2919,N_3226);
nor U8617 (N_8617,N_4963,N_2043);
nor U8618 (N_8618,N_316,N_64);
xnor U8619 (N_8619,N_4179,N_4422);
xor U8620 (N_8620,N_4473,N_1281);
or U8621 (N_8621,N_1550,N_3576);
xnor U8622 (N_8622,N_2413,N_4495);
and U8623 (N_8623,N_1940,N_1282);
xor U8624 (N_8624,N_3747,N_3133);
nor U8625 (N_8625,N_4196,N_565);
nor U8626 (N_8626,N_1306,N_3985);
nand U8627 (N_8627,N_4370,N_3658);
nor U8628 (N_8628,N_3122,N_4522);
and U8629 (N_8629,N_2073,N_4081);
or U8630 (N_8630,N_4797,N_657);
xnor U8631 (N_8631,N_3579,N_1406);
and U8632 (N_8632,N_3051,N_4113);
nand U8633 (N_8633,N_4137,N_2293);
or U8634 (N_8634,N_3725,N_3376);
nand U8635 (N_8635,N_4598,N_547);
or U8636 (N_8636,N_3153,N_2028);
and U8637 (N_8637,N_1659,N_1362);
and U8638 (N_8638,N_1753,N_10);
xnor U8639 (N_8639,N_3706,N_519);
and U8640 (N_8640,N_1043,N_2288);
nor U8641 (N_8641,N_4741,N_1423);
or U8642 (N_8642,N_2270,N_1991);
and U8643 (N_8643,N_1637,N_3998);
xor U8644 (N_8644,N_4425,N_3504);
nor U8645 (N_8645,N_499,N_234);
xnor U8646 (N_8646,N_3044,N_3754);
xor U8647 (N_8647,N_4914,N_97);
nor U8648 (N_8648,N_832,N_4809);
and U8649 (N_8649,N_234,N_1488);
xnor U8650 (N_8650,N_2155,N_416);
nor U8651 (N_8651,N_1645,N_1385);
xor U8652 (N_8652,N_3061,N_819);
nor U8653 (N_8653,N_2725,N_1913);
nand U8654 (N_8654,N_587,N_2844);
xor U8655 (N_8655,N_3704,N_1104);
xor U8656 (N_8656,N_3172,N_1480);
xor U8657 (N_8657,N_4689,N_441);
and U8658 (N_8658,N_1829,N_1711);
nand U8659 (N_8659,N_356,N_2995);
or U8660 (N_8660,N_3615,N_357);
or U8661 (N_8661,N_3758,N_1534);
xnor U8662 (N_8662,N_327,N_3476);
and U8663 (N_8663,N_4515,N_314);
and U8664 (N_8664,N_1056,N_3876);
nor U8665 (N_8665,N_85,N_4724);
or U8666 (N_8666,N_322,N_1456);
or U8667 (N_8667,N_3587,N_3227);
xnor U8668 (N_8668,N_3480,N_2394);
or U8669 (N_8669,N_1436,N_1851);
or U8670 (N_8670,N_3736,N_3020);
xor U8671 (N_8671,N_54,N_4098);
and U8672 (N_8672,N_4131,N_1436);
nand U8673 (N_8673,N_4282,N_3321);
nor U8674 (N_8674,N_3335,N_3102);
and U8675 (N_8675,N_4476,N_1372);
nor U8676 (N_8676,N_578,N_1663);
and U8677 (N_8677,N_2135,N_4824);
xor U8678 (N_8678,N_2425,N_2797);
nor U8679 (N_8679,N_2846,N_4652);
xor U8680 (N_8680,N_2443,N_774);
xor U8681 (N_8681,N_2290,N_3997);
or U8682 (N_8682,N_4578,N_3601);
and U8683 (N_8683,N_3000,N_974);
nand U8684 (N_8684,N_3828,N_1920);
or U8685 (N_8685,N_3748,N_2037);
or U8686 (N_8686,N_547,N_4097);
xor U8687 (N_8687,N_1376,N_132);
xnor U8688 (N_8688,N_1073,N_2831);
xnor U8689 (N_8689,N_901,N_2614);
nand U8690 (N_8690,N_881,N_3814);
xnor U8691 (N_8691,N_3614,N_2654);
nand U8692 (N_8692,N_1691,N_3495);
nand U8693 (N_8693,N_4193,N_2205);
nor U8694 (N_8694,N_488,N_2857);
or U8695 (N_8695,N_3202,N_1128);
nor U8696 (N_8696,N_2516,N_838);
xor U8697 (N_8697,N_4653,N_4566);
and U8698 (N_8698,N_314,N_1185);
nor U8699 (N_8699,N_1584,N_3218);
nor U8700 (N_8700,N_3208,N_3054);
nand U8701 (N_8701,N_1112,N_3512);
and U8702 (N_8702,N_2861,N_2375);
xnor U8703 (N_8703,N_1496,N_4619);
nor U8704 (N_8704,N_4328,N_1948);
and U8705 (N_8705,N_3694,N_1387);
nor U8706 (N_8706,N_325,N_2054);
or U8707 (N_8707,N_1603,N_154);
xnor U8708 (N_8708,N_2020,N_4291);
or U8709 (N_8709,N_134,N_51);
nand U8710 (N_8710,N_757,N_1269);
nor U8711 (N_8711,N_2448,N_2790);
xnor U8712 (N_8712,N_2757,N_2633);
or U8713 (N_8713,N_3211,N_902);
nand U8714 (N_8714,N_1158,N_2598);
nand U8715 (N_8715,N_4557,N_2920);
and U8716 (N_8716,N_2147,N_3125);
nor U8717 (N_8717,N_3349,N_721);
nand U8718 (N_8718,N_1343,N_462);
nor U8719 (N_8719,N_3316,N_4968);
nor U8720 (N_8720,N_1924,N_205);
and U8721 (N_8721,N_3427,N_3105);
or U8722 (N_8722,N_433,N_1972);
nand U8723 (N_8723,N_1564,N_609);
or U8724 (N_8724,N_3297,N_4218);
nand U8725 (N_8725,N_2570,N_2404);
and U8726 (N_8726,N_4435,N_2871);
or U8727 (N_8727,N_482,N_2891);
nand U8728 (N_8728,N_4282,N_1058);
and U8729 (N_8729,N_4848,N_3726);
and U8730 (N_8730,N_2518,N_2209);
xnor U8731 (N_8731,N_4523,N_2788);
nand U8732 (N_8732,N_2926,N_3985);
nand U8733 (N_8733,N_3653,N_3416);
or U8734 (N_8734,N_4549,N_3475);
xor U8735 (N_8735,N_3719,N_3031);
or U8736 (N_8736,N_3021,N_645);
and U8737 (N_8737,N_1654,N_948);
nor U8738 (N_8738,N_3477,N_2312);
and U8739 (N_8739,N_4087,N_1694);
xor U8740 (N_8740,N_4464,N_4658);
and U8741 (N_8741,N_1228,N_1608);
xor U8742 (N_8742,N_2232,N_1253);
and U8743 (N_8743,N_1086,N_1285);
and U8744 (N_8744,N_400,N_1699);
nand U8745 (N_8745,N_3358,N_2249);
or U8746 (N_8746,N_4951,N_2975);
nand U8747 (N_8747,N_2996,N_1769);
nor U8748 (N_8748,N_2822,N_4888);
or U8749 (N_8749,N_2109,N_1482);
or U8750 (N_8750,N_4061,N_2512);
nor U8751 (N_8751,N_3270,N_581);
or U8752 (N_8752,N_3682,N_3935);
xnor U8753 (N_8753,N_4375,N_3931);
nand U8754 (N_8754,N_4738,N_4211);
xnor U8755 (N_8755,N_1798,N_2219);
or U8756 (N_8756,N_3201,N_3515);
and U8757 (N_8757,N_140,N_97);
and U8758 (N_8758,N_2546,N_3935);
nand U8759 (N_8759,N_2385,N_2807);
nand U8760 (N_8760,N_884,N_2335);
nor U8761 (N_8761,N_2321,N_4130);
or U8762 (N_8762,N_615,N_3036);
nand U8763 (N_8763,N_4916,N_243);
or U8764 (N_8764,N_2069,N_4602);
nand U8765 (N_8765,N_1337,N_1369);
xnor U8766 (N_8766,N_2189,N_853);
or U8767 (N_8767,N_932,N_150);
xor U8768 (N_8768,N_2112,N_337);
nor U8769 (N_8769,N_6,N_1814);
nor U8770 (N_8770,N_2730,N_4461);
nor U8771 (N_8771,N_3170,N_1307);
nand U8772 (N_8772,N_411,N_1948);
xnor U8773 (N_8773,N_1339,N_341);
nand U8774 (N_8774,N_3327,N_3387);
and U8775 (N_8775,N_1606,N_3230);
and U8776 (N_8776,N_4812,N_440);
and U8777 (N_8777,N_2102,N_3727);
nand U8778 (N_8778,N_2776,N_4310);
nor U8779 (N_8779,N_1270,N_3884);
or U8780 (N_8780,N_1673,N_2010);
and U8781 (N_8781,N_3745,N_1857);
nor U8782 (N_8782,N_733,N_1297);
xor U8783 (N_8783,N_676,N_1455);
or U8784 (N_8784,N_3557,N_4329);
nand U8785 (N_8785,N_3368,N_3176);
nand U8786 (N_8786,N_1675,N_2606);
or U8787 (N_8787,N_742,N_120);
nand U8788 (N_8788,N_38,N_309);
nor U8789 (N_8789,N_632,N_2032);
and U8790 (N_8790,N_845,N_4525);
or U8791 (N_8791,N_1081,N_1185);
nor U8792 (N_8792,N_767,N_1917);
xor U8793 (N_8793,N_548,N_1433);
nand U8794 (N_8794,N_2169,N_1630);
and U8795 (N_8795,N_2123,N_1877);
xor U8796 (N_8796,N_2290,N_768);
or U8797 (N_8797,N_1572,N_1905);
nand U8798 (N_8798,N_1923,N_1603);
and U8799 (N_8799,N_4446,N_2688);
and U8800 (N_8800,N_1458,N_2812);
nor U8801 (N_8801,N_2761,N_2382);
nand U8802 (N_8802,N_2270,N_3848);
nor U8803 (N_8803,N_541,N_143);
nand U8804 (N_8804,N_3151,N_2165);
and U8805 (N_8805,N_928,N_2049);
or U8806 (N_8806,N_3144,N_4618);
xnor U8807 (N_8807,N_1901,N_3788);
nand U8808 (N_8808,N_53,N_4723);
nor U8809 (N_8809,N_3459,N_4122);
nor U8810 (N_8810,N_1346,N_442);
and U8811 (N_8811,N_809,N_4482);
nand U8812 (N_8812,N_4310,N_671);
and U8813 (N_8813,N_1646,N_748);
or U8814 (N_8814,N_789,N_2689);
nand U8815 (N_8815,N_1214,N_4751);
nor U8816 (N_8816,N_4663,N_1214);
and U8817 (N_8817,N_4347,N_515);
nor U8818 (N_8818,N_2642,N_4276);
xnor U8819 (N_8819,N_1092,N_1411);
xor U8820 (N_8820,N_129,N_2001);
xor U8821 (N_8821,N_4078,N_2721);
and U8822 (N_8822,N_2399,N_4946);
xnor U8823 (N_8823,N_2437,N_506);
and U8824 (N_8824,N_3249,N_4602);
and U8825 (N_8825,N_1209,N_3643);
or U8826 (N_8826,N_2876,N_4884);
nor U8827 (N_8827,N_461,N_272);
nor U8828 (N_8828,N_4190,N_4322);
nand U8829 (N_8829,N_579,N_1022);
nand U8830 (N_8830,N_4840,N_4550);
xor U8831 (N_8831,N_3277,N_1383);
nand U8832 (N_8832,N_4669,N_4509);
xnor U8833 (N_8833,N_4878,N_3882);
nor U8834 (N_8834,N_4969,N_765);
or U8835 (N_8835,N_4053,N_1357);
xor U8836 (N_8836,N_96,N_2338);
nor U8837 (N_8837,N_2943,N_1843);
nor U8838 (N_8838,N_4305,N_3569);
nand U8839 (N_8839,N_3663,N_77);
xor U8840 (N_8840,N_2103,N_2245);
nand U8841 (N_8841,N_3025,N_228);
and U8842 (N_8842,N_1969,N_1723);
or U8843 (N_8843,N_4504,N_4273);
nand U8844 (N_8844,N_775,N_4282);
and U8845 (N_8845,N_3001,N_2577);
nor U8846 (N_8846,N_2898,N_4509);
nand U8847 (N_8847,N_3823,N_1152);
nand U8848 (N_8848,N_2994,N_1430);
nor U8849 (N_8849,N_1796,N_3834);
or U8850 (N_8850,N_1060,N_3231);
nor U8851 (N_8851,N_3077,N_1639);
xor U8852 (N_8852,N_555,N_110);
or U8853 (N_8853,N_1986,N_1692);
xor U8854 (N_8854,N_1498,N_3536);
nor U8855 (N_8855,N_4241,N_4082);
nor U8856 (N_8856,N_3014,N_4517);
and U8857 (N_8857,N_3471,N_317);
or U8858 (N_8858,N_3319,N_2528);
or U8859 (N_8859,N_2382,N_187);
nand U8860 (N_8860,N_889,N_4116);
or U8861 (N_8861,N_4400,N_1739);
or U8862 (N_8862,N_3947,N_3977);
nor U8863 (N_8863,N_885,N_2620);
and U8864 (N_8864,N_2499,N_1539);
or U8865 (N_8865,N_780,N_937);
or U8866 (N_8866,N_4361,N_2319);
nand U8867 (N_8867,N_2195,N_4704);
or U8868 (N_8868,N_4075,N_4863);
xnor U8869 (N_8869,N_4049,N_2630);
and U8870 (N_8870,N_3109,N_2324);
nor U8871 (N_8871,N_193,N_4499);
xnor U8872 (N_8872,N_2186,N_4956);
nor U8873 (N_8873,N_75,N_2409);
nand U8874 (N_8874,N_4352,N_3427);
and U8875 (N_8875,N_2584,N_1576);
and U8876 (N_8876,N_2515,N_2374);
and U8877 (N_8877,N_2211,N_2604);
nor U8878 (N_8878,N_1020,N_363);
or U8879 (N_8879,N_4494,N_503);
or U8880 (N_8880,N_2788,N_1296);
nor U8881 (N_8881,N_4515,N_1227);
nand U8882 (N_8882,N_751,N_3374);
or U8883 (N_8883,N_1468,N_2529);
xnor U8884 (N_8884,N_1189,N_1518);
nor U8885 (N_8885,N_533,N_2974);
nand U8886 (N_8886,N_1839,N_1730);
nand U8887 (N_8887,N_4835,N_4071);
nand U8888 (N_8888,N_4758,N_163);
nand U8889 (N_8889,N_1518,N_1153);
xnor U8890 (N_8890,N_4183,N_4482);
and U8891 (N_8891,N_4337,N_2903);
or U8892 (N_8892,N_3584,N_650);
xnor U8893 (N_8893,N_1213,N_3704);
nand U8894 (N_8894,N_343,N_4912);
nand U8895 (N_8895,N_3409,N_2298);
nor U8896 (N_8896,N_2732,N_1392);
nand U8897 (N_8897,N_735,N_2942);
and U8898 (N_8898,N_2973,N_1378);
nand U8899 (N_8899,N_3193,N_390);
xnor U8900 (N_8900,N_2797,N_2779);
nor U8901 (N_8901,N_106,N_4309);
and U8902 (N_8902,N_3284,N_3463);
nor U8903 (N_8903,N_907,N_3269);
or U8904 (N_8904,N_846,N_944);
or U8905 (N_8905,N_4897,N_3493);
nor U8906 (N_8906,N_2071,N_2758);
nor U8907 (N_8907,N_660,N_2968);
or U8908 (N_8908,N_448,N_422);
or U8909 (N_8909,N_4089,N_1967);
or U8910 (N_8910,N_3250,N_3296);
nand U8911 (N_8911,N_2130,N_192);
and U8912 (N_8912,N_4199,N_122);
nor U8913 (N_8913,N_3898,N_107);
xor U8914 (N_8914,N_3708,N_474);
nor U8915 (N_8915,N_3413,N_3978);
nand U8916 (N_8916,N_1007,N_1284);
and U8917 (N_8917,N_1977,N_4023);
nor U8918 (N_8918,N_3148,N_2691);
xor U8919 (N_8919,N_2679,N_2463);
nand U8920 (N_8920,N_2790,N_981);
xnor U8921 (N_8921,N_2396,N_2448);
or U8922 (N_8922,N_2999,N_4248);
or U8923 (N_8923,N_2273,N_1340);
nand U8924 (N_8924,N_3765,N_4512);
or U8925 (N_8925,N_9,N_3484);
xor U8926 (N_8926,N_3707,N_1430);
nor U8927 (N_8927,N_1735,N_324);
or U8928 (N_8928,N_3791,N_2214);
or U8929 (N_8929,N_608,N_1368);
xor U8930 (N_8930,N_2654,N_3378);
nand U8931 (N_8931,N_2893,N_448);
nand U8932 (N_8932,N_649,N_4336);
or U8933 (N_8933,N_1014,N_2853);
xor U8934 (N_8934,N_70,N_2362);
nand U8935 (N_8935,N_4347,N_2349);
and U8936 (N_8936,N_4876,N_3312);
nand U8937 (N_8937,N_1780,N_1943);
and U8938 (N_8938,N_1306,N_221);
and U8939 (N_8939,N_4273,N_3474);
nor U8940 (N_8940,N_4072,N_3247);
or U8941 (N_8941,N_3910,N_276);
xor U8942 (N_8942,N_104,N_885);
nor U8943 (N_8943,N_2250,N_217);
nand U8944 (N_8944,N_524,N_3452);
nor U8945 (N_8945,N_4044,N_4904);
xor U8946 (N_8946,N_1307,N_2871);
xor U8947 (N_8947,N_628,N_3441);
or U8948 (N_8948,N_506,N_4157);
xnor U8949 (N_8949,N_2782,N_3770);
and U8950 (N_8950,N_2605,N_3063);
nand U8951 (N_8951,N_4890,N_3293);
nand U8952 (N_8952,N_1873,N_1670);
or U8953 (N_8953,N_4396,N_2803);
xor U8954 (N_8954,N_2494,N_2848);
nor U8955 (N_8955,N_3613,N_1081);
xnor U8956 (N_8956,N_4319,N_3318);
xnor U8957 (N_8957,N_2324,N_1563);
nor U8958 (N_8958,N_2828,N_4185);
xnor U8959 (N_8959,N_4961,N_431);
and U8960 (N_8960,N_3818,N_3216);
xor U8961 (N_8961,N_3369,N_1013);
nand U8962 (N_8962,N_2566,N_3938);
or U8963 (N_8963,N_1566,N_1229);
or U8964 (N_8964,N_4412,N_3634);
nor U8965 (N_8965,N_1527,N_593);
and U8966 (N_8966,N_2918,N_1242);
and U8967 (N_8967,N_2971,N_57);
or U8968 (N_8968,N_4132,N_2482);
or U8969 (N_8969,N_2165,N_3619);
xor U8970 (N_8970,N_1179,N_47);
nand U8971 (N_8971,N_478,N_4434);
nor U8972 (N_8972,N_2402,N_1224);
nand U8973 (N_8973,N_1267,N_4124);
or U8974 (N_8974,N_185,N_635);
nand U8975 (N_8975,N_1305,N_2681);
and U8976 (N_8976,N_515,N_2663);
nand U8977 (N_8977,N_3190,N_1488);
and U8978 (N_8978,N_2817,N_2964);
or U8979 (N_8979,N_210,N_1676);
and U8980 (N_8980,N_1867,N_723);
and U8981 (N_8981,N_4727,N_1113);
or U8982 (N_8982,N_4598,N_2411);
nand U8983 (N_8983,N_973,N_3554);
and U8984 (N_8984,N_1198,N_4026);
nand U8985 (N_8985,N_2227,N_1467);
or U8986 (N_8986,N_2712,N_1778);
or U8987 (N_8987,N_1722,N_4906);
nand U8988 (N_8988,N_3722,N_4096);
xnor U8989 (N_8989,N_2583,N_3871);
xnor U8990 (N_8990,N_468,N_1595);
and U8991 (N_8991,N_2558,N_966);
and U8992 (N_8992,N_3540,N_621);
nand U8993 (N_8993,N_4720,N_4331);
nor U8994 (N_8994,N_151,N_2567);
and U8995 (N_8995,N_3832,N_3655);
nand U8996 (N_8996,N_4422,N_2121);
xnor U8997 (N_8997,N_2671,N_1371);
nand U8998 (N_8998,N_60,N_4926);
or U8999 (N_8999,N_1910,N_1353);
and U9000 (N_9000,N_288,N_1228);
nor U9001 (N_9001,N_3010,N_957);
or U9002 (N_9002,N_4615,N_4537);
nor U9003 (N_9003,N_3854,N_1908);
or U9004 (N_9004,N_4827,N_1348);
xor U9005 (N_9005,N_4435,N_3169);
nor U9006 (N_9006,N_2280,N_826);
or U9007 (N_9007,N_2183,N_956);
xor U9008 (N_9008,N_876,N_1851);
nor U9009 (N_9009,N_1048,N_1191);
xnor U9010 (N_9010,N_4251,N_383);
xnor U9011 (N_9011,N_1822,N_1122);
nor U9012 (N_9012,N_3802,N_3896);
and U9013 (N_9013,N_3379,N_4802);
xor U9014 (N_9014,N_2214,N_1922);
and U9015 (N_9015,N_2375,N_1799);
nor U9016 (N_9016,N_2753,N_3635);
nand U9017 (N_9017,N_3740,N_2574);
nand U9018 (N_9018,N_204,N_712);
or U9019 (N_9019,N_3251,N_4260);
nor U9020 (N_9020,N_3145,N_3799);
and U9021 (N_9021,N_4176,N_1562);
and U9022 (N_9022,N_1220,N_1110);
nor U9023 (N_9023,N_3743,N_3977);
and U9024 (N_9024,N_4307,N_1560);
and U9025 (N_9025,N_702,N_4585);
xor U9026 (N_9026,N_1917,N_1699);
nor U9027 (N_9027,N_2675,N_3878);
nand U9028 (N_9028,N_1787,N_2613);
nor U9029 (N_9029,N_2828,N_4440);
or U9030 (N_9030,N_95,N_653);
xnor U9031 (N_9031,N_1954,N_619);
nand U9032 (N_9032,N_3291,N_773);
nor U9033 (N_9033,N_221,N_924);
xnor U9034 (N_9034,N_861,N_2765);
nand U9035 (N_9035,N_4786,N_1083);
xor U9036 (N_9036,N_1682,N_1869);
xor U9037 (N_9037,N_4249,N_3723);
nor U9038 (N_9038,N_134,N_2180);
xnor U9039 (N_9039,N_1739,N_1542);
nand U9040 (N_9040,N_4971,N_2341);
xor U9041 (N_9041,N_3702,N_2341);
nand U9042 (N_9042,N_4048,N_551);
and U9043 (N_9043,N_4173,N_2286);
or U9044 (N_9044,N_3686,N_4309);
nand U9045 (N_9045,N_3287,N_4782);
and U9046 (N_9046,N_4972,N_3737);
xnor U9047 (N_9047,N_4026,N_2049);
nand U9048 (N_9048,N_380,N_2481);
and U9049 (N_9049,N_1348,N_3797);
nor U9050 (N_9050,N_3456,N_1426);
nand U9051 (N_9051,N_2385,N_34);
nand U9052 (N_9052,N_2354,N_3620);
nor U9053 (N_9053,N_221,N_2696);
xnor U9054 (N_9054,N_2121,N_882);
and U9055 (N_9055,N_399,N_164);
xor U9056 (N_9056,N_1522,N_1941);
and U9057 (N_9057,N_3932,N_1809);
and U9058 (N_9058,N_3501,N_594);
nand U9059 (N_9059,N_2143,N_2065);
xnor U9060 (N_9060,N_2800,N_4561);
or U9061 (N_9061,N_2525,N_1635);
xnor U9062 (N_9062,N_496,N_1647);
nand U9063 (N_9063,N_4788,N_1429);
or U9064 (N_9064,N_2685,N_2164);
or U9065 (N_9065,N_3667,N_2726);
nor U9066 (N_9066,N_3198,N_326);
nor U9067 (N_9067,N_4356,N_3710);
nand U9068 (N_9068,N_1463,N_3537);
xnor U9069 (N_9069,N_3259,N_4457);
or U9070 (N_9070,N_410,N_3581);
nor U9071 (N_9071,N_686,N_1712);
nor U9072 (N_9072,N_161,N_10);
or U9073 (N_9073,N_1802,N_2012);
nand U9074 (N_9074,N_2309,N_1740);
and U9075 (N_9075,N_2079,N_995);
xnor U9076 (N_9076,N_3658,N_4418);
nand U9077 (N_9077,N_1203,N_444);
nor U9078 (N_9078,N_2037,N_1300);
nand U9079 (N_9079,N_1879,N_2601);
nor U9080 (N_9080,N_2965,N_2228);
nor U9081 (N_9081,N_461,N_1078);
nor U9082 (N_9082,N_3497,N_644);
and U9083 (N_9083,N_108,N_4215);
xor U9084 (N_9084,N_1927,N_3184);
or U9085 (N_9085,N_2121,N_4002);
nor U9086 (N_9086,N_1162,N_3075);
nand U9087 (N_9087,N_2590,N_4495);
xor U9088 (N_9088,N_645,N_4362);
nor U9089 (N_9089,N_3418,N_4393);
nor U9090 (N_9090,N_834,N_4782);
xor U9091 (N_9091,N_888,N_37);
and U9092 (N_9092,N_1393,N_1781);
nor U9093 (N_9093,N_276,N_2775);
nand U9094 (N_9094,N_2055,N_541);
nor U9095 (N_9095,N_4735,N_3734);
and U9096 (N_9096,N_2447,N_4742);
nor U9097 (N_9097,N_2291,N_628);
xnor U9098 (N_9098,N_4156,N_1748);
or U9099 (N_9099,N_1686,N_4248);
nor U9100 (N_9100,N_3744,N_237);
xnor U9101 (N_9101,N_3338,N_3642);
or U9102 (N_9102,N_2487,N_1718);
nand U9103 (N_9103,N_3710,N_4512);
or U9104 (N_9104,N_557,N_2913);
nand U9105 (N_9105,N_2532,N_3234);
and U9106 (N_9106,N_3050,N_1328);
and U9107 (N_9107,N_1757,N_891);
nand U9108 (N_9108,N_2042,N_1553);
nor U9109 (N_9109,N_3317,N_117);
or U9110 (N_9110,N_1773,N_1759);
or U9111 (N_9111,N_3690,N_891);
xor U9112 (N_9112,N_4824,N_2531);
xor U9113 (N_9113,N_3111,N_2554);
and U9114 (N_9114,N_1578,N_3439);
nor U9115 (N_9115,N_233,N_4358);
and U9116 (N_9116,N_3529,N_1998);
nor U9117 (N_9117,N_4504,N_1733);
nand U9118 (N_9118,N_2262,N_1898);
xor U9119 (N_9119,N_1508,N_1314);
and U9120 (N_9120,N_2927,N_3920);
or U9121 (N_9121,N_663,N_2435);
xnor U9122 (N_9122,N_3243,N_3033);
and U9123 (N_9123,N_4204,N_280);
nor U9124 (N_9124,N_4814,N_3895);
or U9125 (N_9125,N_4484,N_325);
and U9126 (N_9126,N_4963,N_1437);
nand U9127 (N_9127,N_3520,N_2018);
xnor U9128 (N_9128,N_4113,N_3137);
xor U9129 (N_9129,N_3360,N_2219);
nor U9130 (N_9130,N_4488,N_3163);
and U9131 (N_9131,N_2627,N_323);
nor U9132 (N_9132,N_480,N_3837);
xnor U9133 (N_9133,N_1085,N_1339);
or U9134 (N_9134,N_387,N_1023);
or U9135 (N_9135,N_2345,N_2056);
nand U9136 (N_9136,N_1553,N_1282);
nand U9137 (N_9137,N_1688,N_778);
nor U9138 (N_9138,N_4879,N_3538);
nand U9139 (N_9139,N_4191,N_3494);
nand U9140 (N_9140,N_1060,N_1246);
nand U9141 (N_9141,N_2561,N_2777);
nand U9142 (N_9142,N_3123,N_2779);
xor U9143 (N_9143,N_1373,N_1467);
or U9144 (N_9144,N_3378,N_2519);
nor U9145 (N_9145,N_3465,N_4671);
xnor U9146 (N_9146,N_4982,N_783);
nand U9147 (N_9147,N_4795,N_1141);
nand U9148 (N_9148,N_1411,N_1890);
xor U9149 (N_9149,N_4577,N_2712);
xnor U9150 (N_9150,N_1182,N_2192);
or U9151 (N_9151,N_3647,N_3645);
xnor U9152 (N_9152,N_3592,N_2022);
nand U9153 (N_9153,N_878,N_764);
nor U9154 (N_9154,N_1663,N_4617);
xor U9155 (N_9155,N_4701,N_2448);
nand U9156 (N_9156,N_1269,N_850);
nor U9157 (N_9157,N_699,N_253);
nor U9158 (N_9158,N_4940,N_4732);
nor U9159 (N_9159,N_2883,N_4850);
or U9160 (N_9160,N_3289,N_2474);
or U9161 (N_9161,N_1602,N_829);
nor U9162 (N_9162,N_683,N_2101);
nor U9163 (N_9163,N_3983,N_803);
and U9164 (N_9164,N_4346,N_4148);
nor U9165 (N_9165,N_912,N_4612);
nand U9166 (N_9166,N_2471,N_1730);
or U9167 (N_9167,N_2047,N_2903);
xor U9168 (N_9168,N_4190,N_1148);
and U9169 (N_9169,N_481,N_33);
or U9170 (N_9170,N_2315,N_3696);
nor U9171 (N_9171,N_3645,N_529);
and U9172 (N_9172,N_4704,N_3759);
nand U9173 (N_9173,N_393,N_1341);
nand U9174 (N_9174,N_1550,N_3150);
and U9175 (N_9175,N_3626,N_3818);
or U9176 (N_9176,N_1175,N_2802);
and U9177 (N_9177,N_3355,N_2857);
nand U9178 (N_9178,N_1681,N_3538);
and U9179 (N_9179,N_4431,N_2642);
xor U9180 (N_9180,N_2207,N_265);
and U9181 (N_9181,N_3754,N_3119);
and U9182 (N_9182,N_1358,N_1749);
and U9183 (N_9183,N_4841,N_3558);
and U9184 (N_9184,N_1203,N_580);
xnor U9185 (N_9185,N_2848,N_195);
or U9186 (N_9186,N_1474,N_4449);
xnor U9187 (N_9187,N_2600,N_587);
nand U9188 (N_9188,N_2436,N_3154);
xor U9189 (N_9189,N_1794,N_4472);
or U9190 (N_9190,N_1893,N_3599);
nand U9191 (N_9191,N_3054,N_1039);
xnor U9192 (N_9192,N_1005,N_98);
or U9193 (N_9193,N_745,N_2875);
nor U9194 (N_9194,N_1689,N_2139);
xnor U9195 (N_9195,N_4840,N_859);
or U9196 (N_9196,N_2853,N_478);
and U9197 (N_9197,N_658,N_4246);
or U9198 (N_9198,N_3825,N_1973);
nor U9199 (N_9199,N_1173,N_1871);
or U9200 (N_9200,N_4421,N_1147);
nand U9201 (N_9201,N_3202,N_762);
or U9202 (N_9202,N_4036,N_2727);
and U9203 (N_9203,N_1371,N_4031);
or U9204 (N_9204,N_1160,N_3096);
and U9205 (N_9205,N_1331,N_4501);
or U9206 (N_9206,N_2998,N_290);
xnor U9207 (N_9207,N_4093,N_149);
nand U9208 (N_9208,N_3946,N_59);
and U9209 (N_9209,N_2511,N_4647);
xor U9210 (N_9210,N_1968,N_3119);
nor U9211 (N_9211,N_1513,N_348);
xor U9212 (N_9212,N_3059,N_4360);
xor U9213 (N_9213,N_4742,N_613);
and U9214 (N_9214,N_2440,N_870);
nor U9215 (N_9215,N_4982,N_4617);
or U9216 (N_9216,N_597,N_4184);
xor U9217 (N_9217,N_2719,N_4694);
nand U9218 (N_9218,N_2728,N_4289);
and U9219 (N_9219,N_1143,N_2937);
or U9220 (N_9220,N_2123,N_1739);
xnor U9221 (N_9221,N_1774,N_2463);
nand U9222 (N_9222,N_1707,N_4243);
xnor U9223 (N_9223,N_4343,N_3020);
xor U9224 (N_9224,N_3329,N_2253);
nor U9225 (N_9225,N_837,N_1831);
and U9226 (N_9226,N_678,N_3666);
xor U9227 (N_9227,N_925,N_1933);
and U9228 (N_9228,N_3691,N_4832);
nor U9229 (N_9229,N_2178,N_162);
nor U9230 (N_9230,N_466,N_4679);
xor U9231 (N_9231,N_531,N_311);
nand U9232 (N_9232,N_951,N_2979);
xor U9233 (N_9233,N_2281,N_4230);
and U9234 (N_9234,N_3525,N_2898);
nand U9235 (N_9235,N_1246,N_1572);
and U9236 (N_9236,N_340,N_3959);
nand U9237 (N_9237,N_3350,N_315);
nand U9238 (N_9238,N_564,N_1131);
or U9239 (N_9239,N_3889,N_1431);
nand U9240 (N_9240,N_2514,N_2344);
nand U9241 (N_9241,N_1111,N_4248);
nor U9242 (N_9242,N_1354,N_314);
and U9243 (N_9243,N_2414,N_4146);
nand U9244 (N_9244,N_1398,N_777);
xnor U9245 (N_9245,N_2975,N_3715);
nand U9246 (N_9246,N_2964,N_840);
and U9247 (N_9247,N_4640,N_2280);
xor U9248 (N_9248,N_4617,N_3968);
and U9249 (N_9249,N_1321,N_3057);
nor U9250 (N_9250,N_1707,N_1298);
or U9251 (N_9251,N_2911,N_281);
nand U9252 (N_9252,N_3231,N_825);
nor U9253 (N_9253,N_1694,N_1267);
xor U9254 (N_9254,N_2415,N_3008);
nor U9255 (N_9255,N_1257,N_1601);
and U9256 (N_9256,N_65,N_3231);
nor U9257 (N_9257,N_1791,N_1507);
and U9258 (N_9258,N_2705,N_4559);
xnor U9259 (N_9259,N_2684,N_2280);
or U9260 (N_9260,N_4084,N_2108);
nand U9261 (N_9261,N_3472,N_1701);
or U9262 (N_9262,N_811,N_1823);
and U9263 (N_9263,N_1267,N_3202);
and U9264 (N_9264,N_3189,N_2002);
or U9265 (N_9265,N_2449,N_2589);
nand U9266 (N_9266,N_2475,N_85);
nand U9267 (N_9267,N_1728,N_3721);
nand U9268 (N_9268,N_4596,N_2654);
and U9269 (N_9269,N_4390,N_2047);
xnor U9270 (N_9270,N_377,N_3544);
nand U9271 (N_9271,N_430,N_2377);
nand U9272 (N_9272,N_3813,N_129);
xnor U9273 (N_9273,N_4869,N_212);
and U9274 (N_9274,N_2798,N_2524);
nand U9275 (N_9275,N_1440,N_2139);
nor U9276 (N_9276,N_620,N_3820);
nand U9277 (N_9277,N_184,N_316);
nor U9278 (N_9278,N_319,N_4402);
or U9279 (N_9279,N_3376,N_3091);
nand U9280 (N_9280,N_4683,N_736);
xor U9281 (N_9281,N_4297,N_3751);
nand U9282 (N_9282,N_4887,N_2552);
nor U9283 (N_9283,N_406,N_1805);
and U9284 (N_9284,N_1730,N_193);
or U9285 (N_9285,N_3563,N_3543);
nand U9286 (N_9286,N_167,N_2935);
nor U9287 (N_9287,N_1586,N_2577);
or U9288 (N_9288,N_788,N_2404);
nor U9289 (N_9289,N_480,N_2895);
nand U9290 (N_9290,N_1067,N_1282);
xnor U9291 (N_9291,N_3149,N_2786);
xnor U9292 (N_9292,N_1596,N_1038);
or U9293 (N_9293,N_1579,N_4116);
and U9294 (N_9294,N_1991,N_2335);
or U9295 (N_9295,N_3839,N_1810);
and U9296 (N_9296,N_1084,N_2638);
and U9297 (N_9297,N_2019,N_1413);
and U9298 (N_9298,N_969,N_3123);
xnor U9299 (N_9299,N_834,N_3658);
nor U9300 (N_9300,N_4534,N_3432);
xor U9301 (N_9301,N_3496,N_4767);
nand U9302 (N_9302,N_2928,N_2611);
xnor U9303 (N_9303,N_4434,N_4674);
nor U9304 (N_9304,N_1251,N_2345);
nand U9305 (N_9305,N_3561,N_2953);
nor U9306 (N_9306,N_2035,N_2985);
nand U9307 (N_9307,N_4504,N_3581);
or U9308 (N_9308,N_4287,N_2274);
or U9309 (N_9309,N_4049,N_3588);
and U9310 (N_9310,N_1128,N_3226);
and U9311 (N_9311,N_4733,N_1389);
xnor U9312 (N_9312,N_3093,N_3848);
xnor U9313 (N_9313,N_4176,N_4609);
xor U9314 (N_9314,N_4683,N_4941);
nor U9315 (N_9315,N_4694,N_1355);
xnor U9316 (N_9316,N_933,N_57);
and U9317 (N_9317,N_3370,N_3569);
nand U9318 (N_9318,N_1520,N_4225);
or U9319 (N_9319,N_4478,N_3051);
nand U9320 (N_9320,N_2379,N_2581);
or U9321 (N_9321,N_3173,N_4427);
xnor U9322 (N_9322,N_3061,N_1809);
or U9323 (N_9323,N_4075,N_149);
nand U9324 (N_9324,N_2757,N_4704);
and U9325 (N_9325,N_1943,N_2733);
xor U9326 (N_9326,N_4832,N_2818);
xor U9327 (N_9327,N_2655,N_2026);
nand U9328 (N_9328,N_4231,N_889);
xnor U9329 (N_9329,N_2987,N_391);
and U9330 (N_9330,N_3602,N_4769);
nor U9331 (N_9331,N_3481,N_2543);
nor U9332 (N_9332,N_4838,N_1096);
nor U9333 (N_9333,N_832,N_2258);
and U9334 (N_9334,N_1349,N_628);
xnor U9335 (N_9335,N_3608,N_1594);
and U9336 (N_9336,N_2841,N_1655);
xnor U9337 (N_9337,N_4679,N_2648);
nor U9338 (N_9338,N_1506,N_1514);
nor U9339 (N_9339,N_2420,N_2809);
or U9340 (N_9340,N_3073,N_4098);
nand U9341 (N_9341,N_4854,N_1788);
xor U9342 (N_9342,N_1229,N_4364);
or U9343 (N_9343,N_4484,N_3527);
nand U9344 (N_9344,N_1342,N_2691);
or U9345 (N_9345,N_2300,N_2147);
nand U9346 (N_9346,N_2945,N_4727);
xor U9347 (N_9347,N_1952,N_3235);
xnor U9348 (N_9348,N_1735,N_4097);
nor U9349 (N_9349,N_1703,N_868);
nand U9350 (N_9350,N_343,N_1570);
nor U9351 (N_9351,N_2159,N_2988);
and U9352 (N_9352,N_1021,N_4824);
or U9353 (N_9353,N_93,N_4551);
and U9354 (N_9354,N_1448,N_3026);
xor U9355 (N_9355,N_2898,N_580);
nand U9356 (N_9356,N_4169,N_923);
and U9357 (N_9357,N_4307,N_856);
xor U9358 (N_9358,N_2499,N_838);
and U9359 (N_9359,N_598,N_4766);
and U9360 (N_9360,N_2593,N_1985);
and U9361 (N_9361,N_2547,N_4230);
xnor U9362 (N_9362,N_3039,N_3892);
nor U9363 (N_9363,N_2171,N_245);
nor U9364 (N_9364,N_3132,N_4252);
nand U9365 (N_9365,N_1091,N_4430);
nor U9366 (N_9366,N_3994,N_713);
nor U9367 (N_9367,N_3361,N_2924);
nand U9368 (N_9368,N_1329,N_1773);
nor U9369 (N_9369,N_378,N_4478);
and U9370 (N_9370,N_2713,N_3231);
nand U9371 (N_9371,N_431,N_1620);
and U9372 (N_9372,N_1217,N_47);
xnor U9373 (N_9373,N_2288,N_4322);
and U9374 (N_9374,N_866,N_775);
and U9375 (N_9375,N_333,N_3971);
and U9376 (N_9376,N_75,N_4534);
or U9377 (N_9377,N_2998,N_764);
xor U9378 (N_9378,N_1404,N_3980);
nor U9379 (N_9379,N_1948,N_1229);
or U9380 (N_9380,N_2179,N_2500);
xor U9381 (N_9381,N_4600,N_592);
and U9382 (N_9382,N_2226,N_1634);
and U9383 (N_9383,N_19,N_3043);
and U9384 (N_9384,N_4515,N_1301);
nor U9385 (N_9385,N_2265,N_165);
and U9386 (N_9386,N_1989,N_2481);
or U9387 (N_9387,N_2384,N_3937);
nor U9388 (N_9388,N_3315,N_105);
xor U9389 (N_9389,N_152,N_1557);
nand U9390 (N_9390,N_4414,N_4102);
and U9391 (N_9391,N_1465,N_4944);
nor U9392 (N_9392,N_4215,N_2365);
nor U9393 (N_9393,N_2690,N_4005);
xnor U9394 (N_9394,N_2266,N_457);
and U9395 (N_9395,N_2381,N_1930);
nor U9396 (N_9396,N_4577,N_1199);
and U9397 (N_9397,N_1423,N_3418);
nor U9398 (N_9398,N_644,N_4038);
or U9399 (N_9399,N_3423,N_3751);
nor U9400 (N_9400,N_3363,N_2573);
nor U9401 (N_9401,N_3779,N_3401);
nand U9402 (N_9402,N_4663,N_1009);
or U9403 (N_9403,N_3335,N_4155);
nor U9404 (N_9404,N_4657,N_2397);
nand U9405 (N_9405,N_3768,N_3501);
or U9406 (N_9406,N_4039,N_4948);
and U9407 (N_9407,N_3855,N_1577);
xnor U9408 (N_9408,N_1973,N_4633);
xor U9409 (N_9409,N_2185,N_169);
nor U9410 (N_9410,N_2902,N_2685);
and U9411 (N_9411,N_3257,N_4854);
nand U9412 (N_9412,N_3342,N_2631);
nand U9413 (N_9413,N_3013,N_231);
nor U9414 (N_9414,N_4733,N_3237);
or U9415 (N_9415,N_3531,N_1051);
and U9416 (N_9416,N_4683,N_4648);
nor U9417 (N_9417,N_1942,N_4936);
and U9418 (N_9418,N_2190,N_3599);
or U9419 (N_9419,N_2399,N_4479);
nor U9420 (N_9420,N_4434,N_3524);
nor U9421 (N_9421,N_4752,N_4392);
or U9422 (N_9422,N_3943,N_2361);
xnor U9423 (N_9423,N_2790,N_1198);
nand U9424 (N_9424,N_2360,N_4617);
and U9425 (N_9425,N_1946,N_3867);
xnor U9426 (N_9426,N_111,N_3166);
nor U9427 (N_9427,N_3972,N_814);
or U9428 (N_9428,N_2394,N_2728);
nand U9429 (N_9429,N_3417,N_4052);
or U9430 (N_9430,N_4435,N_3150);
nor U9431 (N_9431,N_4937,N_4894);
or U9432 (N_9432,N_4223,N_1802);
xor U9433 (N_9433,N_1855,N_3575);
xnor U9434 (N_9434,N_280,N_3512);
nor U9435 (N_9435,N_4512,N_426);
and U9436 (N_9436,N_1247,N_1040);
and U9437 (N_9437,N_4252,N_2013);
or U9438 (N_9438,N_3909,N_3287);
nand U9439 (N_9439,N_155,N_3782);
nor U9440 (N_9440,N_2626,N_858);
and U9441 (N_9441,N_724,N_4133);
and U9442 (N_9442,N_59,N_1762);
and U9443 (N_9443,N_539,N_381);
nor U9444 (N_9444,N_42,N_2268);
and U9445 (N_9445,N_224,N_532);
xnor U9446 (N_9446,N_4538,N_676);
nand U9447 (N_9447,N_283,N_2104);
and U9448 (N_9448,N_3388,N_3001);
xor U9449 (N_9449,N_743,N_3964);
nand U9450 (N_9450,N_1118,N_3739);
or U9451 (N_9451,N_2627,N_2561);
nor U9452 (N_9452,N_2578,N_2991);
nand U9453 (N_9453,N_3867,N_2603);
or U9454 (N_9454,N_2659,N_4668);
or U9455 (N_9455,N_2567,N_2686);
xor U9456 (N_9456,N_4245,N_2701);
xnor U9457 (N_9457,N_3248,N_4739);
nand U9458 (N_9458,N_852,N_45);
nand U9459 (N_9459,N_3766,N_4508);
or U9460 (N_9460,N_1039,N_3520);
xnor U9461 (N_9461,N_642,N_2294);
nor U9462 (N_9462,N_985,N_4741);
nand U9463 (N_9463,N_1991,N_4050);
or U9464 (N_9464,N_2495,N_4013);
and U9465 (N_9465,N_1258,N_1186);
nand U9466 (N_9466,N_4492,N_4852);
xor U9467 (N_9467,N_2932,N_1179);
or U9468 (N_9468,N_3102,N_3851);
and U9469 (N_9469,N_2425,N_1102);
and U9470 (N_9470,N_3419,N_296);
nor U9471 (N_9471,N_4376,N_4897);
nor U9472 (N_9472,N_1863,N_1839);
nand U9473 (N_9473,N_220,N_2383);
and U9474 (N_9474,N_3764,N_1742);
nor U9475 (N_9475,N_4275,N_3574);
xnor U9476 (N_9476,N_4796,N_2918);
xor U9477 (N_9477,N_4062,N_4578);
nand U9478 (N_9478,N_3404,N_3299);
or U9479 (N_9479,N_1952,N_805);
and U9480 (N_9480,N_6,N_3857);
nand U9481 (N_9481,N_74,N_216);
or U9482 (N_9482,N_971,N_1181);
nand U9483 (N_9483,N_1644,N_4637);
or U9484 (N_9484,N_545,N_4963);
or U9485 (N_9485,N_4711,N_4555);
nand U9486 (N_9486,N_3467,N_1989);
or U9487 (N_9487,N_4228,N_2439);
nand U9488 (N_9488,N_2403,N_2706);
xnor U9489 (N_9489,N_4027,N_1708);
or U9490 (N_9490,N_3698,N_389);
nor U9491 (N_9491,N_493,N_1635);
or U9492 (N_9492,N_944,N_4259);
nand U9493 (N_9493,N_2906,N_3962);
nand U9494 (N_9494,N_4727,N_789);
nor U9495 (N_9495,N_1164,N_3211);
xnor U9496 (N_9496,N_41,N_3154);
xor U9497 (N_9497,N_2858,N_174);
nand U9498 (N_9498,N_586,N_2676);
nor U9499 (N_9499,N_628,N_4764);
nand U9500 (N_9500,N_4612,N_1227);
xor U9501 (N_9501,N_116,N_2042);
nand U9502 (N_9502,N_3716,N_638);
nor U9503 (N_9503,N_2581,N_266);
nand U9504 (N_9504,N_1070,N_4237);
and U9505 (N_9505,N_1190,N_1849);
nor U9506 (N_9506,N_3393,N_3543);
nor U9507 (N_9507,N_2779,N_4515);
xor U9508 (N_9508,N_908,N_3616);
or U9509 (N_9509,N_249,N_1665);
nor U9510 (N_9510,N_4410,N_3152);
nand U9511 (N_9511,N_3753,N_2932);
xor U9512 (N_9512,N_4052,N_1638);
nand U9513 (N_9513,N_3679,N_2801);
and U9514 (N_9514,N_2357,N_2482);
xnor U9515 (N_9515,N_2356,N_1392);
nor U9516 (N_9516,N_855,N_207);
or U9517 (N_9517,N_133,N_1658);
nand U9518 (N_9518,N_3799,N_4391);
nand U9519 (N_9519,N_624,N_2820);
nand U9520 (N_9520,N_2157,N_3486);
or U9521 (N_9521,N_3599,N_3347);
nor U9522 (N_9522,N_2804,N_3111);
xor U9523 (N_9523,N_4136,N_1486);
and U9524 (N_9524,N_120,N_3357);
nor U9525 (N_9525,N_759,N_4948);
and U9526 (N_9526,N_541,N_1834);
xnor U9527 (N_9527,N_4212,N_4829);
or U9528 (N_9528,N_4832,N_3341);
and U9529 (N_9529,N_374,N_634);
xnor U9530 (N_9530,N_2254,N_4010);
nand U9531 (N_9531,N_1047,N_1215);
nand U9532 (N_9532,N_3630,N_1680);
nand U9533 (N_9533,N_1720,N_4136);
or U9534 (N_9534,N_1703,N_3681);
and U9535 (N_9535,N_3819,N_2089);
and U9536 (N_9536,N_3474,N_4040);
or U9537 (N_9537,N_1563,N_4449);
or U9538 (N_9538,N_2297,N_3834);
and U9539 (N_9539,N_2898,N_3899);
nor U9540 (N_9540,N_942,N_113);
xnor U9541 (N_9541,N_2825,N_3596);
and U9542 (N_9542,N_2774,N_560);
and U9543 (N_9543,N_3792,N_4216);
nor U9544 (N_9544,N_612,N_4644);
nand U9545 (N_9545,N_216,N_4841);
nor U9546 (N_9546,N_4527,N_2232);
and U9547 (N_9547,N_1822,N_2617);
or U9548 (N_9548,N_3675,N_823);
xor U9549 (N_9549,N_564,N_663);
nand U9550 (N_9550,N_1715,N_3928);
and U9551 (N_9551,N_634,N_300);
xor U9552 (N_9552,N_2670,N_1865);
xnor U9553 (N_9553,N_2345,N_4871);
xnor U9554 (N_9554,N_1961,N_1818);
or U9555 (N_9555,N_134,N_1621);
or U9556 (N_9556,N_3759,N_834);
and U9557 (N_9557,N_654,N_2784);
nand U9558 (N_9558,N_831,N_526);
nor U9559 (N_9559,N_1847,N_197);
or U9560 (N_9560,N_4233,N_2035);
or U9561 (N_9561,N_638,N_198);
or U9562 (N_9562,N_561,N_1487);
nand U9563 (N_9563,N_1511,N_2126);
and U9564 (N_9564,N_3148,N_1063);
nand U9565 (N_9565,N_1594,N_3129);
xor U9566 (N_9566,N_2582,N_4606);
nor U9567 (N_9567,N_3678,N_1540);
and U9568 (N_9568,N_362,N_242);
or U9569 (N_9569,N_1589,N_4473);
nor U9570 (N_9570,N_3019,N_1754);
xor U9571 (N_9571,N_4792,N_203);
nand U9572 (N_9572,N_3254,N_959);
and U9573 (N_9573,N_3398,N_167);
nor U9574 (N_9574,N_962,N_1956);
nor U9575 (N_9575,N_1779,N_2731);
nor U9576 (N_9576,N_2226,N_1720);
nor U9577 (N_9577,N_2990,N_2052);
nand U9578 (N_9578,N_2810,N_4510);
and U9579 (N_9579,N_1363,N_4600);
xor U9580 (N_9580,N_845,N_4558);
xor U9581 (N_9581,N_3600,N_44);
and U9582 (N_9582,N_932,N_992);
nor U9583 (N_9583,N_3962,N_4476);
nor U9584 (N_9584,N_3121,N_3747);
nand U9585 (N_9585,N_2262,N_3815);
and U9586 (N_9586,N_3972,N_4823);
xnor U9587 (N_9587,N_2797,N_4723);
and U9588 (N_9588,N_819,N_2638);
and U9589 (N_9589,N_4394,N_1750);
xnor U9590 (N_9590,N_3687,N_3546);
nor U9591 (N_9591,N_1116,N_3709);
or U9592 (N_9592,N_587,N_2349);
nor U9593 (N_9593,N_662,N_3828);
xor U9594 (N_9594,N_226,N_3825);
and U9595 (N_9595,N_4811,N_3943);
nand U9596 (N_9596,N_3789,N_4568);
and U9597 (N_9597,N_1271,N_2069);
nor U9598 (N_9598,N_4393,N_4740);
nand U9599 (N_9599,N_839,N_613);
xor U9600 (N_9600,N_4359,N_2920);
nor U9601 (N_9601,N_4016,N_2443);
nor U9602 (N_9602,N_1912,N_3374);
nand U9603 (N_9603,N_1225,N_3840);
nor U9604 (N_9604,N_3071,N_1346);
nor U9605 (N_9605,N_2679,N_3538);
nand U9606 (N_9606,N_3475,N_3390);
or U9607 (N_9607,N_4717,N_336);
xor U9608 (N_9608,N_3343,N_398);
nor U9609 (N_9609,N_2600,N_1475);
and U9610 (N_9610,N_1850,N_2935);
or U9611 (N_9611,N_3139,N_1943);
and U9612 (N_9612,N_2673,N_4969);
or U9613 (N_9613,N_4139,N_909);
xnor U9614 (N_9614,N_3560,N_1112);
nand U9615 (N_9615,N_3917,N_156);
or U9616 (N_9616,N_2444,N_1561);
nand U9617 (N_9617,N_469,N_3353);
and U9618 (N_9618,N_3354,N_2571);
xor U9619 (N_9619,N_2612,N_4124);
or U9620 (N_9620,N_4999,N_453);
nor U9621 (N_9621,N_2452,N_136);
xnor U9622 (N_9622,N_1517,N_1292);
or U9623 (N_9623,N_2127,N_4749);
xnor U9624 (N_9624,N_2913,N_4873);
and U9625 (N_9625,N_702,N_1770);
nand U9626 (N_9626,N_2984,N_825);
and U9627 (N_9627,N_1997,N_4573);
xnor U9628 (N_9628,N_1067,N_1982);
xnor U9629 (N_9629,N_1753,N_4539);
nor U9630 (N_9630,N_3604,N_2699);
and U9631 (N_9631,N_3947,N_2211);
or U9632 (N_9632,N_1802,N_4925);
nand U9633 (N_9633,N_3886,N_4254);
or U9634 (N_9634,N_1222,N_787);
or U9635 (N_9635,N_471,N_2939);
nand U9636 (N_9636,N_594,N_889);
and U9637 (N_9637,N_4953,N_3830);
or U9638 (N_9638,N_2092,N_1588);
or U9639 (N_9639,N_3088,N_221);
nand U9640 (N_9640,N_3258,N_944);
nand U9641 (N_9641,N_3201,N_137);
xor U9642 (N_9642,N_4646,N_1564);
and U9643 (N_9643,N_1165,N_1369);
xnor U9644 (N_9644,N_1467,N_1672);
xor U9645 (N_9645,N_2607,N_317);
xor U9646 (N_9646,N_1572,N_1755);
xnor U9647 (N_9647,N_1865,N_689);
and U9648 (N_9648,N_2617,N_4747);
nor U9649 (N_9649,N_3255,N_147);
xnor U9650 (N_9650,N_4404,N_2577);
nor U9651 (N_9651,N_3428,N_3135);
xnor U9652 (N_9652,N_599,N_3197);
or U9653 (N_9653,N_2712,N_4772);
or U9654 (N_9654,N_1746,N_4808);
nand U9655 (N_9655,N_1197,N_95);
or U9656 (N_9656,N_1174,N_995);
nand U9657 (N_9657,N_4290,N_2362);
or U9658 (N_9658,N_463,N_982);
and U9659 (N_9659,N_642,N_973);
nor U9660 (N_9660,N_1707,N_1390);
and U9661 (N_9661,N_4585,N_2262);
or U9662 (N_9662,N_4861,N_4571);
or U9663 (N_9663,N_1270,N_945);
or U9664 (N_9664,N_1106,N_13);
and U9665 (N_9665,N_3568,N_4800);
or U9666 (N_9666,N_2266,N_2885);
nor U9667 (N_9667,N_1395,N_2610);
and U9668 (N_9668,N_3802,N_4303);
nor U9669 (N_9669,N_1667,N_3124);
xnor U9670 (N_9670,N_1356,N_3040);
xor U9671 (N_9671,N_510,N_4892);
and U9672 (N_9672,N_3699,N_3381);
nand U9673 (N_9673,N_1320,N_2041);
nor U9674 (N_9674,N_3044,N_3523);
nor U9675 (N_9675,N_247,N_4356);
xor U9676 (N_9676,N_385,N_352);
nor U9677 (N_9677,N_1920,N_3301);
or U9678 (N_9678,N_3234,N_4849);
or U9679 (N_9679,N_1855,N_3185);
nor U9680 (N_9680,N_374,N_2645);
nand U9681 (N_9681,N_1202,N_4204);
nand U9682 (N_9682,N_3545,N_322);
or U9683 (N_9683,N_4483,N_3999);
or U9684 (N_9684,N_4877,N_4434);
xor U9685 (N_9685,N_530,N_479);
and U9686 (N_9686,N_4009,N_3543);
and U9687 (N_9687,N_1907,N_3386);
xnor U9688 (N_9688,N_3583,N_1562);
or U9689 (N_9689,N_1627,N_2514);
or U9690 (N_9690,N_2440,N_2501);
or U9691 (N_9691,N_4731,N_2866);
nand U9692 (N_9692,N_2471,N_1319);
nand U9693 (N_9693,N_2531,N_1307);
nor U9694 (N_9694,N_1002,N_2243);
xor U9695 (N_9695,N_180,N_2282);
nand U9696 (N_9696,N_3858,N_2421);
or U9697 (N_9697,N_4039,N_4690);
and U9698 (N_9698,N_1686,N_4426);
nor U9699 (N_9699,N_4213,N_4244);
nand U9700 (N_9700,N_2708,N_2531);
and U9701 (N_9701,N_1216,N_2874);
or U9702 (N_9702,N_2972,N_1757);
nor U9703 (N_9703,N_4903,N_1153);
and U9704 (N_9704,N_1540,N_2189);
and U9705 (N_9705,N_3369,N_3177);
xnor U9706 (N_9706,N_2185,N_2468);
and U9707 (N_9707,N_3465,N_1037);
and U9708 (N_9708,N_2162,N_928);
nand U9709 (N_9709,N_4392,N_2845);
or U9710 (N_9710,N_2208,N_4694);
nor U9711 (N_9711,N_3428,N_3375);
xnor U9712 (N_9712,N_4156,N_302);
and U9713 (N_9713,N_1953,N_898);
xor U9714 (N_9714,N_3950,N_306);
xor U9715 (N_9715,N_3400,N_4292);
xnor U9716 (N_9716,N_4269,N_1201);
xor U9717 (N_9717,N_4683,N_526);
and U9718 (N_9718,N_1054,N_3332);
and U9719 (N_9719,N_4739,N_2670);
xor U9720 (N_9720,N_4885,N_4518);
nor U9721 (N_9721,N_2890,N_3497);
xor U9722 (N_9722,N_1687,N_1758);
nor U9723 (N_9723,N_1268,N_4818);
or U9724 (N_9724,N_2722,N_1358);
or U9725 (N_9725,N_2854,N_4231);
or U9726 (N_9726,N_1294,N_2321);
xor U9727 (N_9727,N_1784,N_461);
nor U9728 (N_9728,N_2341,N_1988);
nand U9729 (N_9729,N_1444,N_2114);
nor U9730 (N_9730,N_2044,N_4412);
nand U9731 (N_9731,N_870,N_1841);
nand U9732 (N_9732,N_1693,N_4725);
nor U9733 (N_9733,N_67,N_2868);
nand U9734 (N_9734,N_3908,N_1539);
nor U9735 (N_9735,N_4090,N_2387);
or U9736 (N_9736,N_2720,N_348);
xnor U9737 (N_9737,N_3791,N_2162);
nand U9738 (N_9738,N_2128,N_3073);
or U9739 (N_9739,N_3124,N_2484);
or U9740 (N_9740,N_1037,N_3455);
xnor U9741 (N_9741,N_715,N_1163);
and U9742 (N_9742,N_434,N_3750);
nor U9743 (N_9743,N_1197,N_1225);
nor U9744 (N_9744,N_1735,N_3543);
xor U9745 (N_9745,N_3824,N_4638);
and U9746 (N_9746,N_15,N_4126);
nand U9747 (N_9747,N_2589,N_1320);
and U9748 (N_9748,N_3511,N_1269);
nor U9749 (N_9749,N_1959,N_1875);
or U9750 (N_9750,N_4527,N_3866);
and U9751 (N_9751,N_1339,N_274);
xnor U9752 (N_9752,N_35,N_2842);
nand U9753 (N_9753,N_3294,N_2659);
nor U9754 (N_9754,N_4083,N_495);
nand U9755 (N_9755,N_1929,N_2148);
nand U9756 (N_9756,N_260,N_407);
or U9757 (N_9757,N_3428,N_2062);
and U9758 (N_9758,N_4793,N_3063);
nor U9759 (N_9759,N_4812,N_438);
nand U9760 (N_9760,N_4559,N_4701);
or U9761 (N_9761,N_4796,N_3449);
xor U9762 (N_9762,N_4771,N_4754);
nand U9763 (N_9763,N_1251,N_1107);
and U9764 (N_9764,N_4115,N_4481);
or U9765 (N_9765,N_4303,N_2971);
xor U9766 (N_9766,N_737,N_2431);
xor U9767 (N_9767,N_4224,N_313);
nor U9768 (N_9768,N_1162,N_308);
nor U9769 (N_9769,N_4212,N_4208);
and U9770 (N_9770,N_1509,N_4425);
and U9771 (N_9771,N_3564,N_170);
nor U9772 (N_9772,N_1289,N_1790);
or U9773 (N_9773,N_4886,N_4399);
nor U9774 (N_9774,N_3026,N_1948);
or U9775 (N_9775,N_171,N_4325);
nor U9776 (N_9776,N_2256,N_4296);
xor U9777 (N_9777,N_2525,N_3722);
xor U9778 (N_9778,N_3833,N_1522);
nand U9779 (N_9779,N_3795,N_3157);
xnor U9780 (N_9780,N_4450,N_4153);
or U9781 (N_9781,N_4653,N_861);
and U9782 (N_9782,N_3506,N_3735);
or U9783 (N_9783,N_2763,N_1777);
or U9784 (N_9784,N_155,N_2936);
or U9785 (N_9785,N_3385,N_1093);
nand U9786 (N_9786,N_704,N_1950);
nand U9787 (N_9787,N_4402,N_3023);
or U9788 (N_9788,N_1312,N_2818);
and U9789 (N_9789,N_4401,N_3179);
and U9790 (N_9790,N_2741,N_2024);
and U9791 (N_9791,N_1042,N_3170);
and U9792 (N_9792,N_2311,N_4236);
xor U9793 (N_9793,N_472,N_4665);
nor U9794 (N_9794,N_2191,N_893);
nor U9795 (N_9795,N_2929,N_4378);
and U9796 (N_9796,N_3760,N_4710);
nand U9797 (N_9797,N_4702,N_3704);
and U9798 (N_9798,N_1617,N_2509);
nand U9799 (N_9799,N_1272,N_962);
nand U9800 (N_9800,N_1179,N_3290);
or U9801 (N_9801,N_154,N_3894);
nor U9802 (N_9802,N_4693,N_1511);
or U9803 (N_9803,N_4970,N_1094);
nand U9804 (N_9804,N_70,N_2850);
and U9805 (N_9805,N_105,N_1076);
nor U9806 (N_9806,N_2200,N_4433);
nand U9807 (N_9807,N_2514,N_1465);
xnor U9808 (N_9808,N_4864,N_1774);
or U9809 (N_9809,N_2523,N_3703);
and U9810 (N_9810,N_4318,N_751);
nand U9811 (N_9811,N_3348,N_107);
nand U9812 (N_9812,N_1816,N_264);
and U9813 (N_9813,N_2360,N_637);
or U9814 (N_9814,N_4995,N_1247);
xor U9815 (N_9815,N_2623,N_2219);
nand U9816 (N_9816,N_1493,N_2206);
nand U9817 (N_9817,N_229,N_3222);
or U9818 (N_9818,N_2741,N_3616);
nor U9819 (N_9819,N_342,N_3787);
or U9820 (N_9820,N_1587,N_1974);
nor U9821 (N_9821,N_3030,N_896);
or U9822 (N_9822,N_2298,N_381);
xnor U9823 (N_9823,N_2338,N_2511);
nor U9824 (N_9824,N_4378,N_3978);
and U9825 (N_9825,N_1319,N_4589);
and U9826 (N_9826,N_542,N_1428);
nand U9827 (N_9827,N_1068,N_1170);
and U9828 (N_9828,N_799,N_3206);
xnor U9829 (N_9829,N_3025,N_3176);
and U9830 (N_9830,N_639,N_3775);
nand U9831 (N_9831,N_678,N_2378);
nor U9832 (N_9832,N_3303,N_2761);
nand U9833 (N_9833,N_99,N_4457);
xor U9834 (N_9834,N_1325,N_3381);
and U9835 (N_9835,N_1928,N_1633);
or U9836 (N_9836,N_502,N_577);
nand U9837 (N_9837,N_807,N_4787);
xor U9838 (N_9838,N_2820,N_4153);
nor U9839 (N_9839,N_4625,N_4546);
xor U9840 (N_9840,N_2901,N_1097);
or U9841 (N_9841,N_2871,N_2508);
or U9842 (N_9842,N_2956,N_4122);
and U9843 (N_9843,N_90,N_4790);
xnor U9844 (N_9844,N_3130,N_4700);
nand U9845 (N_9845,N_1933,N_1576);
or U9846 (N_9846,N_2818,N_3996);
xor U9847 (N_9847,N_1216,N_2178);
nand U9848 (N_9848,N_2036,N_3592);
or U9849 (N_9849,N_4511,N_88);
nand U9850 (N_9850,N_2545,N_737);
nand U9851 (N_9851,N_2490,N_1908);
and U9852 (N_9852,N_3280,N_3287);
nor U9853 (N_9853,N_85,N_2048);
xnor U9854 (N_9854,N_481,N_4745);
nor U9855 (N_9855,N_3940,N_4117);
nand U9856 (N_9856,N_1591,N_2188);
xnor U9857 (N_9857,N_1204,N_4651);
nand U9858 (N_9858,N_1275,N_2888);
xor U9859 (N_9859,N_2518,N_2023);
or U9860 (N_9860,N_3763,N_1026);
or U9861 (N_9861,N_2057,N_127);
xor U9862 (N_9862,N_2970,N_4999);
and U9863 (N_9863,N_3867,N_2000);
or U9864 (N_9864,N_2725,N_4349);
nand U9865 (N_9865,N_1038,N_4953);
nor U9866 (N_9866,N_1823,N_4674);
or U9867 (N_9867,N_716,N_4008);
nand U9868 (N_9868,N_4859,N_2936);
nor U9869 (N_9869,N_1322,N_3832);
or U9870 (N_9870,N_3801,N_3740);
and U9871 (N_9871,N_4111,N_4907);
xnor U9872 (N_9872,N_2344,N_3546);
or U9873 (N_9873,N_1439,N_758);
xor U9874 (N_9874,N_4997,N_581);
or U9875 (N_9875,N_3483,N_942);
or U9876 (N_9876,N_1637,N_2590);
xnor U9877 (N_9877,N_2110,N_3163);
and U9878 (N_9878,N_1709,N_4571);
and U9879 (N_9879,N_1485,N_2435);
nand U9880 (N_9880,N_1173,N_2038);
or U9881 (N_9881,N_3980,N_3195);
or U9882 (N_9882,N_122,N_3692);
and U9883 (N_9883,N_2545,N_1658);
nand U9884 (N_9884,N_4875,N_466);
nor U9885 (N_9885,N_1709,N_3400);
and U9886 (N_9886,N_2583,N_2863);
nand U9887 (N_9887,N_25,N_3857);
or U9888 (N_9888,N_3279,N_3306);
and U9889 (N_9889,N_4344,N_3319);
nor U9890 (N_9890,N_2578,N_1034);
nand U9891 (N_9891,N_4447,N_1710);
and U9892 (N_9892,N_4745,N_2180);
or U9893 (N_9893,N_1291,N_2569);
and U9894 (N_9894,N_1531,N_4830);
and U9895 (N_9895,N_1448,N_617);
and U9896 (N_9896,N_1446,N_4426);
nand U9897 (N_9897,N_3798,N_4473);
and U9898 (N_9898,N_1820,N_2724);
or U9899 (N_9899,N_3780,N_1524);
nand U9900 (N_9900,N_1566,N_2852);
nor U9901 (N_9901,N_129,N_355);
xor U9902 (N_9902,N_3707,N_1591);
xnor U9903 (N_9903,N_4726,N_4490);
nand U9904 (N_9904,N_808,N_4238);
and U9905 (N_9905,N_3246,N_2604);
nor U9906 (N_9906,N_748,N_3164);
or U9907 (N_9907,N_3680,N_3466);
nand U9908 (N_9908,N_3268,N_4961);
xor U9909 (N_9909,N_1047,N_4910);
nor U9910 (N_9910,N_447,N_3096);
nand U9911 (N_9911,N_4835,N_4985);
and U9912 (N_9912,N_119,N_231);
nor U9913 (N_9913,N_706,N_284);
or U9914 (N_9914,N_116,N_3118);
and U9915 (N_9915,N_4347,N_3929);
nor U9916 (N_9916,N_4339,N_649);
or U9917 (N_9917,N_1789,N_2106);
and U9918 (N_9918,N_2152,N_799);
nor U9919 (N_9919,N_2789,N_634);
nand U9920 (N_9920,N_487,N_1903);
nand U9921 (N_9921,N_3185,N_4810);
nand U9922 (N_9922,N_2675,N_1144);
nor U9923 (N_9923,N_152,N_1874);
or U9924 (N_9924,N_617,N_2250);
xnor U9925 (N_9925,N_1920,N_1702);
nand U9926 (N_9926,N_3615,N_404);
and U9927 (N_9927,N_4330,N_3996);
or U9928 (N_9928,N_1332,N_2252);
nor U9929 (N_9929,N_2425,N_3337);
xnor U9930 (N_9930,N_4747,N_828);
and U9931 (N_9931,N_1059,N_2845);
and U9932 (N_9932,N_4698,N_1229);
nand U9933 (N_9933,N_3292,N_1508);
xnor U9934 (N_9934,N_1003,N_4952);
or U9935 (N_9935,N_4167,N_402);
nor U9936 (N_9936,N_3876,N_1932);
nor U9937 (N_9937,N_3131,N_2971);
nand U9938 (N_9938,N_2046,N_2378);
or U9939 (N_9939,N_4782,N_3098);
nand U9940 (N_9940,N_1985,N_2867);
and U9941 (N_9941,N_1501,N_353);
nand U9942 (N_9942,N_1384,N_1273);
or U9943 (N_9943,N_3512,N_895);
nand U9944 (N_9944,N_2738,N_3419);
or U9945 (N_9945,N_4224,N_517);
or U9946 (N_9946,N_3659,N_4666);
or U9947 (N_9947,N_319,N_1642);
and U9948 (N_9948,N_3039,N_1018);
xor U9949 (N_9949,N_2329,N_4490);
nor U9950 (N_9950,N_814,N_2442);
nand U9951 (N_9951,N_3939,N_1138);
and U9952 (N_9952,N_2262,N_31);
nand U9953 (N_9953,N_4587,N_4272);
or U9954 (N_9954,N_3865,N_3575);
xnor U9955 (N_9955,N_612,N_3271);
xor U9956 (N_9956,N_166,N_262);
xnor U9957 (N_9957,N_3917,N_3182);
and U9958 (N_9958,N_2955,N_3202);
or U9959 (N_9959,N_4687,N_2758);
or U9960 (N_9960,N_2116,N_3436);
nor U9961 (N_9961,N_3539,N_3002);
nand U9962 (N_9962,N_1487,N_93);
or U9963 (N_9963,N_685,N_1566);
nand U9964 (N_9964,N_1157,N_4981);
nand U9965 (N_9965,N_2809,N_766);
or U9966 (N_9966,N_3241,N_4564);
or U9967 (N_9967,N_1664,N_2106);
xnor U9968 (N_9968,N_1599,N_4125);
nor U9969 (N_9969,N_3467,N_1550);
xor U9970 (N_9970,N_2073,N_3140);
xnor U9971 (N_9971,N_1892,N_3441);
xnor U9972 (N_9972,N_4707,N_1847);
and U9973 (N_9973,N_3104,N_1917);
nor U9974 (N_9974,N_4405,N_4410);
xnor U9975 (N_9975,N_4045,N_2213);
and U9976 (N_9976,N_252,N_4835);
and U9977 (N_9977,N_1145,N_2324);
xor U9978 (N_9978,N_2939,N_76);
xnor U9979 (N_9979,N_1576,N_905);
or U9980 (N_9980,N_1894,N_2402);
and U9981 (N_9981,N_288,N_2598);
nor U9982 (N_9982,N_4844,N_293);
and U9983 (N_9983,N_4475,N_1914);
nor U9984 (N_9984,N_4926,N_644);
or U9985 (N_9985,N_2610,N_2779);
nand U9986 (N_9986,N_122,N_3383);
nand U9987 (N_9987,N_2196,N_1800);
xnor U9988 (N_9988,N_4547,N_2680);
nor U9989 (N_9989,N_3440,N_736);
nand U9990 (N_9990,N_3810,N_3247);
xor U9991 (N_9991,N_1692,N_1275);
nor U9992 (N_9992,N_2801,N_4783);
and U9993 (N_9993,N_2066,N_4009);
or U9994 (N_9994,N_618,N_824);
nand U9995 (N_9995,N_2803,N_3183);
or U9996 (N_9996,N_2881,N_1843);
nand U9997 (N_9997,N_2372,N_3426);
nand U9998 (N_9998,N_2528,N_4388);
nor U9999 (N_9999,N_2999,N_37);
xnor U10000 (N_10000,N_8594,N_5345);
xor U10001 (N_10001,N_6371,N_6335);
nand U10002 (N_10002,N_7462,N_7468);
nor U10003 (N_10003,N_7805,N_6740);
or U10004 (N_10004,N_9606,N_8750);
nor U10005 (N_10005,N_7895,N_7296);
nand U10006 (N_10006,N_6469,N_5021);
xor U10007 (N_10007,N_9103,N_8610);
or U10008 (N_10008,N_6158,N_6035);
nor U10009 (N_10009,N_8154,N_6544);
or U10010 (N_10010,N_6029,N_7672);
nor U10011 (N_10011,N_5362,N_6174);
xor U10012 (N_10012,N_6163,N_6661);
nand U10013 (N_10013,N_8850,N_6139);
or U10014 (N_10014,N_8684,N_7121);
nand U10015 (N_10015,N_6282,N_9706);
and U10016 (N_10016,N_6954,N_8045);
or U10017 (N_10017,N_5924,N_6413);
xor U10018 (N_10018,N_9254,N_8419);
nand U10019 (N_10019,N_7127,N_6470);
nor U10020 (N_10020,N_9758,N_6673);
nand U10021 (N_10021,N_8585,N_7311);
xor U10022 (N_10022,N_7245,N_7486);
or U10023 (N_10023,N_7667,N_9482);
nor U10024 (N_10024,N_7679,N_9846);
xor U10025 (N_10025,N_6758,N_8710);
xnor U10026 (N_10026,N_9666,N_8893);
nand U10027 (N_10027,N_6595,N_8074);
and U10028 (N_10028,N_9720,N_7852);
nand U10029 (N_10029,N_8844,N_9598);
xor U10030 (N_10030,N_9541,N_9984);
nand U10031 (N_10031,N_5286,N_8784);
xnor U10032 (N_10032,N_7971,N_7379);
nand U10033 (N_10033,N_9524,N_7749);
nor U10034 (N_10034,N_8060,N_7936);
and U10035 (N_10035,N_9663,N_8012);
nand U10036 (N_10036,N_5084,N_6564);
and U10037 (N_10037,N_8523,N_9561);
nand U10038 (N_10038,N_6644,N_5927);
and U10039 (N_10039,N_6505,N_6071);
or U10040 (N_10040,N_7859,N_7457);
nand U10041 (N_10041,N_5097,N_6419);
and U10042 (N_10042,N_8270,N_6002);
xor U10043 (N_10043,N_6635,N_7281);
or U10044 (N_10044,N_7785,N_8630);
xnor U10045 (N_10045,N_5184,N_5235);
nand U10046 (N_10046,N_6225,N_6657);
and U10047 (N_10047,N_7878,N_8520);
xnor U10048 (N_10048,N_6884,N_5569);
and U10049 (N_10049,N_6963,N_6379);
nand U10050 (N_10050,N_8998,N_7545);
xnor U10051 (N_10051,N_5769,N_6919);
or U10052 (N_10052,N_7080,N_9430);
or U10053 (N_10053,N_9263,N_7164);
and U10054 (N_10054,N_9310,N_8008);
or U10055 (N_10055,N_7294,N_9415);
or U10056 (N_10056,N_8459,N_9992);
xor U10057 (N_10057,N_7451,N_5478);
and U10058 (N_10058,N_6995,N_6286);
and U10059 (N_10059,N_8628,N_8297);
nor U10060 (N_10060,N_7882,N_7409);
and U10061 (N_10061,N_8526,N_9490);
and U10062 (N_10062,N_9852,N_6345);
or U10063 (N_10063,N_8997,N_6777);
nor U10064 (N_10064,N_8841,N_9968);
or U10065 (N_10065,N_7243,N_9843);
or U10066 (N_10066,N_5009,N_8541);
nand U10067 (N_10067,N_9053,N_5399);
nand U10068 (N_10068,N_6024,N_6079);
or U10069 (N_10069,N_6845,N_5206);
nor U10070 (N_10070,N_5249,N_5827);
nand U10071 (N_10071,N_8747,N_7691);
nand U10072 (N_10072,N_7159,N_9759);
or U10073 (N_10073,N_7980,N_8047);
xnor U10074 (N_10074,N_9258,N_8188);
nor U10075 (N_10075,N_5656,N_6309);
and U10076 (N_10076,N_8957,N_9700);
nand U10077 (N_10077,N_5208,N_5290);
nand U10078 (N_10078,N_7408,N_8615);
nor U10079 (N_10079,N_6625,N_9115);
and U10080 (N_10080,N_9382,N_7982);
and U10081 (N_10081,N_8635,N_7088);
and U10082 (N_10082,N_9776,N_9345);
or U10083 (N_10083,N_5234,N_9256);
or U10084 (N_10084,N_5522,N_8518);
nor U10085 (N_10085,N_5441,N_8253);
nand U10086 (N_10086,N_7270,N_6007);
xnor U10087 (N_10087,N_8268,N_7183);
and U10088 (N_10088,N_7410,N_5634);
or U10089 (N_10089,N_8279,N_5632);
xor U10090 (N_10090,N_6500,N_6528);
or U10091 (N_10091,N_9909,N_8597);
nand U10092 (N_10092,N_8760,N_7232);
xnor U10093 (N_10093,N_9083,N_7189);
nand U10094 (N_10094,N_8796,N_9049);
and U10095 (N_10095,N_5979,N_7222);
or U10096 (N_10096,N_7107,N_7598);
and U10097 (N_10097,N_9161,N_7039);
xor U10098 (N_10098,N_8495,N_7782);
and U10099 (N_10099,N_5390,N_9460);
nor U10100 (N_10100,N_7745,N_6878);
nand U10101 (N_10101,N_7132,N_9965);
nand U10102 (N_10102,N_6868,N_6365);
xnor U10103 (N_10103,N_6981,N_8174);
xor U10104 (N_10104,N_7372,N_7688);
nand U10105 (N_10105,N_5156,N_6367);
nand U10106 (N_10106,N_6811,N_8143);
or U10107 (N_10107,N_9540,N_6802);
nor U10108 (N_10108,N_6630,N_9238);
and U10109 (N_10109,N_6116,N_8579);
xnor U10110 (N_10110,N_7122,N_9546);
nand U10111 (N_10111,N_9592,N_6162);
and U10112 (N_10112,N_5863,N_6111);
nand U10113 (N_10113,N_8129,N_7732);
nor U10114 (N_10114,N_8803,N_6817);
nor U10115 (N_10115,N_7074,N_8073);
nor U10116 (N_10116,N_6858,N_8681);
nand U10117 (N_10117,N_6499,N_6452);
xor U10118 (N_10118,N_5236,N_7970);
xnor U10119 (N_10119,N_5066,N_6570);
nor U10120 (N_10120,N_8137,N_6252);
xnor U10121 (N_10121,N_8554,N_8612);
nor U10122 (N_10122,N_5720,N_9178);
nor U10123 (N_10123,N_8689,N_9383);
nor U10124 (N_10124,N_8500,N_8503);
xor U10125 (N_10125,N_8805,N_5262);
nor U10126 (N_10126,N_5670,N_9569);
and U10127 (N_10127,N_5452,N_7877);
nand U10128 (N_10128,N_9020,N_8015);
or U10129 (N_10129,N_6623,N_8490);
xor U10130 (N_10130,N_5346,N_6479);
and U10131 (N_10131,N_8574,N_8931);
nor U10132 (N_10132,N_6140,N_9389);
or U10133 (N_10133,N_6331,N_8314);
xnor U10134 (N_10134,N_5611,N_8237);
nor U10135 (N_10135,N_9272,N_7856);
nand U10136 (N_10136,N_9227,N_8219);
nand U10137 (N_10137,N_6480,N_5466);
nand U10138 (N_10138,N_6456,N_9275);
or U10139 (N_10139,N_6507,N_5287);
and U10140 (N_10140,N_5157,N_5451);
nor U10141 (N_10141,N_9976,N_6268);
xnor U10142 (N_10142,N_8552,N_9654);
or U10143 (N_10143,N_9499,N_6382);
nor U10144 (N_10144,N_9514,N_8011);
nand U10145 (N_10145,N_8192,N_5059);
xor U10146 (N_10146,N_5558,N_5931);
xor U10147 (N_10147,N_5047,N_5978);
nand U10148 (N_10148,N_9682,N_6068);
xor U10149 (N_10149,N_5505,N_7260);
and U10150 (N_10150,N_7307,N_6596);
xor U10151 (N_10151,N_8470,N_5976);
nand U10152 (N_10152,N_9449,N_6049);
and U10153 (N_10153,N_6267,N_6511);
xnor U10154 (N_10154,N_9420,N_7280);
nor U10155 (N_10155,N_9826,N_6904);
nand U10156 (N_10156,N_9007,N_5412);
nor U10157 (N_10157,N_7276,N_9640);
nand U10158 (N_10158,N_6287,N_8066);
xnor U10159 (N_10159,N_7831,N_8860);
nand U10160 (N_10160,N_9412,N_6491);
xor U10161 (N_10161,N_7933,N_7310);
or U10162 (N_10162,N_8139,N_9403);
and U10163 (N_10163,N_9599,N_9018);
nand U10164 (N_10164,N_9819,N_9211);
nor U10165 (N_10165,N_7459,N_9423);
or U10166 (N_10166,N_8780,N_6149);
nand U10167 (N_10167,N_8598,N_7618);
nor U10168 (N_10168,N_5756,N_7730);
nand U10169 (N_10169,N_9248,N_9804);
xor U10170 (N_10170,N_9332,N_8051);
or U10171 (N_10171,N_8538,N_5594);
or U10172 (N_10172,N_5644,N_5108);
xor U10173 (N_10173,N_7205,N_7670);
and U10174 (N_10174,N_7966,N_9151);
and U10175 (N_10175,N_7113,N_7326);
and U10176 (N_10176,N_5518,N_7776);
nor U10177 (N_10177,N_9709,N_8974);
or U10178 (N_10178,N_6546,N_7028);
xnor U10179 (N_10179,N_7550,N_7577);
nor U10180 (N_10180,N_6654,N_6567);
or U10181 (N_10181,N_5337,N_6349);
and U10182 (N_10182,N_8383,N_8611);
or U10183 (N_10183,N_5414,N_8527);
or U10184 (N_10184,N_8903,N_5155);
xor U10185 (N_10185,N_9989,N_5661);
and U10186 (N_10186,N_9816,N_5483);
and U10187 (N_10187,N_5418,N_6830);
xnor U10188 (N_10188,N_9084,N_5783);
and U10189 (N_10189,N_6683,N_6976);
nand U10190 (N_10190,N_6014,N_5557);
or U10191 (N_10191,N_7511,N_8070);
nand U10192 (N_10192,N_7286,N_8899);
nand U10193 (N_10193,N_6430,N_7634);
or U10194 (N_10194,N_7458,N_9851);
nand U10195 (N_10195,N_7279,N_9455);
and U10196 (N_10196,N_5355,N_8148);
or U10197 (N_10197,N_7325,N_9864);
and U10198 (N_10198,N_5192,N_9690);
or U10199 (N_10199,N_6446,N_7197);
nor U10200 (N_10200,N_6765,N_8214);
nand U10201 (N_10201,N_9557,N_6783);
and U10202 (N_10202,N_7365,N_9260);
nor U10203 (N_10203,N_6501,N_7002);
xor U10204 (N_10204,N_9315,N_5830);
nand U10205 (N_10205,N_7680,N_6509);
and U10206 (N_10206,N_5061,N_8524);
or U10207 (N_10207,N_9408,N_7820);
or U10208 (N_10208,N_6601,N_5387);
nor U10209 (N_10209,N_9250,N_6108);
or U10210 (N_10210,N_9164,N_6649);
and U10211 (N_10211,N_7804,N_5782);
nand U10212 (N_10212,N_5831,N_6561);
and U10213 (N_10213,N_8178,N_6241);
and U10214 (N_10214,N_9707,N_5396);
nand U10215 (N_10215,N_5091,N_5794);
nor U10216 (N_10216,N_8306,N_8382);
nand U10217 (N_10217,N_5460,N_8983);
and U10218 (N_10218,N_8026,N_8591);
and U10219 (N_10219,N_9642,N_5012);
nand U10220 (N_10220,N_9808,N_7777);
nand U10221 (N_10221,N_9177,N_9409);
or U10222 (N_10222,N_7573,N_9450);
or U10223 (N_10223,N_5143,N_5667);
xnor U10224 (N_10224,N_6343,N_5991);
nand U10225 (N_10225,N_9361,N_7125);
nand U10226 (N_10226,N_5673,N_8556);
and U10227 (N_10227,N_5808,N_5544);
nand U10228 (N_10228,N_8986,N_5364);
nand U10229 (N_10229,N_5648,N_5440);
xor U10230 (N_10230,N_9960,N_9346);
nand U10231 (N_10231,N_8406,N_9464);
nor U10232 (N_10232,N_8264,N_7144);
and U10233 (N_10233,N_7789,N_6555);
nand U10234 (N_10234,N_7078,N_8030);
nand U10235 (N_10235,N_9171,N_6016);
or U10236 (N_10236,N_9214,N_5573);
xor U10237 (N_10237,N_8659,N_8711);
xnor U10238 (N_10238,N_6098,N_9981);
nor U10239 (N_10239,N_6619,N_5763);
xnor U10240 (N_10240,N_9442,N_7542);
nand U10241 (N_10241,N_5966,N_5902);
nand U10242 (N_10242,N_6305,N_7721);
or U10243 (N_10243,N_9006,N_6993);
nand U10244 (N_10244,N_8245,N_9107);
nand U10245 (N_10245,N_6097,N_8854);
nor U10246 (N_10246,N_7101,N_6790);
nand U10247 (N_10247,N_9761,N_7910);
nor U10248 (N_10248,N_6171,N_8879);
nor U10249 (N_10249,N_8272,N_8657);
or U10250 (N_10250,N_9590,N_5423);
xnor U10251 (N_10251,N_8818,N_7682);
nor U10252 (N_10252,N_8123,N_5107);
nor U10253 (N_10253,N_7244,N_7689);
nor U10254 (N_10254,N_7665,N_5883);
xnor U10255 (N_10255,N_9046,N_9842);
nand U10256 (N_10256,N_6584,N_6312);
and U10257 (N_10257,N_8894,N_7707);
nor U10258 (N_10258,N_9121,N_7059);
or U10259 (N_10259,N_9193,N_9280);
xor U10260 (N_10260,N_9363,N_9247);
and U10261 (N_10261,N_5868,N_7534);
xor U10262 (N_10262,N_8125,N_5175);
xnor U10263 (N_10263,N_8400,N_7601);
or U10264 (N_10264,N_5899,N_5903);
xor U10265 (N_10265,N_9692,N_7850);
nor U10266 (N_10266,N_7187,N_9052);
xnor U10267 (N_10267,N_5496,N_5067);
nand U10268 (N_10268,N_8863,N_5013);
xnor U10269 (N_10269,N_6231,N_5637);
xor U10270 (N_10270,N_6147,N_7069);
or U10271 (N_10271,N_8592,N_8679);
nor U10272 (N_10272,N_9777,N_9478);
nor U10273 (N_10273,N_7498,N_6871);
and U10274 (N_10274,N_6614,N_9390);
and U10275 (N_10275,N_9696,N_9883);
and U10276 (N_10276,N_8771,N_6733);
nor U10277 (N_10277,N_5566,N_8309);
and U10278 (N_10278,N_7606,N_5260);
xnor U10279 (N_10279,N_9088,N_7212);
nor U10280 (N_10280,N_7677,N_9378);
or U10281 (N_10281,N_8876,N_9518);
nand U10282 (N_10282,N_6086,N_9985);
nor U10283 (N_10283,N_6984,N_5689);
and U10284 (N_10284,N_9385,N_8951);
xor U10285 (N_10285,N_5223,N_8212);
and U10286 (N_10286,N_6234,N_7546);
or U10287 (N_10287,N_7753,N_5560);
and U10288 (N_10288,N_5854,N_7566);
xor U10289 (N_10289,N_5737,N_8791);
or U10290 (N_10290,N_7536,N_5607);
xnor U10291 (N_10291,N_5652,N_8985);
and U10292 (N_10292,N_9319,N_8457);
xor U10293 (N_10293,N_6468,N_9814);
nor U10294 (N_10294,N_7807,N_7399);
and U10295 (N_10295,N_9235,N_7520);
xnor U10296 (N_10296,N_8763,N_6013);
or U10297 (N_10297,N_7156,N_7337);
nor U10298 (N_10298,N_9778,N_5011);
and U10299 (N_10299,N_8878,N_7652);
and U10300 (N_10300,N_5178,N_5385);
or U10301 (N_10301,N_9653,N_7173);
xor U10302 (N_10302,N_6609,N_6730);
nand U10303 (N_10303,N_5666,N_9194);
or U10304 (N_10304,N_9501,N_8277);
xor U10305 (N_10305,N_9135,N_5838);
nand U10306 (N_10306,N_9505,N_7447);
or U10307 (N_10307,N_5153,N_5542);
or U10308 (N_10308,N_6368,N_9217);
or U10309 (N_10309,N_7609,N_8081);
nor U10310 (N_10310,N_8159,N_8901);
xnor U10311 (N_10311,N_6399,N_7622);
xnor U10312 (N_10312,N_6443,N_6893);
nor U10313 (N_10313,N_9497,N_8607);
nand U10314 (N_10314,N_8867,N_5866);
nand U10315 (N_10315,N_7876,N_5056);
xnor U10316 (N_10316,N_7847,N_8057);
xnor U10317 (N_10317,N_6944,N_8732);
or U10318 (N_10318,N_9186,N_7576);
and U10319 (N_10319,N_7258,N_9737);
and U10320 (N_10320,N_7810,N_6914);
nor U10321 (N_10321,N_8472,N_8558);
nor U10322 (N_10322,N_7908,N_5245);
xor U10323 (N_10323,N_8834,N_5599);
nand U10324 (N_10324,N_9069,N_5023);
or U10325 (N_10325,N_5210,N_7434);
xnor U10326 (N_10326,N_7621,N_5041);
and U10327 (N_10327,N_6854,N_8649);
or U10328 (N_10328,N_7729,N_6210);
xnor U10329 (N_10329,N_7502,N_5218);
nand U10330 (N_10330,N_5513,N_7517);
nor U10331 (N_10331,N_7168,N_7111);
and U10332 (N_10332,N_9036,N_6253);
and U10333 (N_10333,N_8157,N_6136);
nor U10334 (N_10334,N_8310,N_7449);
nor U10335 (N_10335,N_7975,N_9352);
xnor U10336 (N_10336,N_7515,N_7196);
xor U10337 (N_10337,N_9948,N_6156);
nand U10338 (N_10338,N_5243,N_6428);
and U10339 (N_10339,N_8151,N_5620);
nand U10340 (N_10340,N_8257,N_7461);
nand U10341 (N_10341,N_8466,N_6762);
or U10342 (N_10342,N_8856,N_9322);
and U10343 (N_10343,N_6977,N_7917);
or U10344 (N_10344,N_6028,N_8748);
nand U10345 (N_10345,N_7705,N_5626);
nand U10346 (N_10346,N_5474,N_7932);
nand U10347 (N_10347,N_6131,N_6226);
nor U10348 (N_10348,N_5029,N_7154);
nor U10349 (N_10349,N_7646,N_8601);
or U10350 (N_10350,N_7623,N_6061);
nand U10351 (N_10351,N_9025,N_5070);
nor U10352 (N_10352,N_7544,N_6994);
nor U10353 (N_10353,N_9773,N_6110);
or U10354 (N_10354,N_8355,N_5182);
nand U10355 (N_10355,N_8966,N_9508);
nor U10356 (N_10356,N_6838,N_5517);
xnor U10357 (N_10357,N_9652,N_7578);
or U10358 (N_10358,N_5616,N_8745);
and U10359 (N_10359,N_5371,N_5617);
nand U10360 (N_10360,N_5468,N_7087);
nand U10361 (N_10361,N_7950,N_9298);
nor U10362 (N_10362,N_9915,N_7809);
nor U10363 (N_10363,N_7851,N_5344);
nor U10364 (N_10364,N_9169,N_7483);
and U10365 (N_10365,N_5915,N_9600);
or U10366 (N_10366,N_8738,N_6196);
or U10367 (N_10367,N_9535,N_5456);
nor U10368 (N_10368,N_8298,N_8980);
nor U10369 (N_10369,N_6451,N_6167);
xnor U10370 (N_10370,N_8839,N_9304);
and U10371 (N_10371,N_6890,N_6193);
xnor U10372 (N_10372,N_8491,N_9243);
and U10373 (N_10373,N_5370,N_7951);
xnor U10374 (N_10374,N_7713,N_7103);
and U10375 (N_10375,N_7999,N_6988);
nand U10376 (N_10376,N_9209,N_6251);
and U10377 (N_10377,N_7097,N_9645);
xor U10378 (N_10378,N_7563,N_6659);
nand U10379 (N_10379,N_5732,N_6771);
nor U10380 (N_10380,N_9101,N_6322);
or U10381 (N_10381,N_9627,N_9399);
nand U10382 (N_10382,N_5824,N_8437);
nor U10383 (N_10383,N_9405,N_7633);
xor U10384 (N_10384,N_6752,N_7822);
and U10385 (N_10385,N_6532,N_5350);
and U10386 (N_10386,N_5189,N_5302);
xnor U10387 (N_10387,N_7055,N_8971);
xnor U10388 (N_10388,N_6788,N_7026);
and U10389 (N_10389,N_7217,N_6690);
or U10390 (N_10390,N_5836,N_8977);
nor U10391 (N_10391,N_9887,N_9647);
xor U10392 (N_10392,N_5610,N_9456);
and U10393 (N_10393,N_5404,N_5685);
nand U10394 (N_10394,N_7538,N_5716);
nand U10395 (N_10395,N_7480,N_7134);
nor U10396 (N_10396,N_6205,N_8956);
nand U10397 (N_10397,N_7118,N_5051);
or U10398 (N_10398,N_5062,N_9753);
nand U10399 (N_10399,N_8058,N_8708);
nor U10400 (N_10400,N_5211,N_9743);
nor U10401 (N_10401,N_8874,N_9017);
and U10402 (N_10402,N_6266,N_7463);
nor U10403 (N_10403,N_9605,N_7991);
and U10404 (N_10404,N_6582,N_9366);
nor U10405 (N_10405,N_9521,N_8654);
nand U10406 (N_10406,N_7869,N_5778);
nand U10407 (N_10407,N_8002,N_9001);
and U10408 (N_10408,N_6834,N_8728);
nand U10409 (N_10409,N_7916,N_7861);
or U10410 (N_10410,N_7763,N_6209);
or U10411 (N_10411,N_5072,N_6172);
xor U10412 (N_10412,N_7959,N_6454);
xnor U10413 (N_10413,N_8937,N_5909);
nand U10414 (N_10414,N_9034,N_7129);
and U10415 (N_10415,N_6153,N_9588);
or U10416 (N_10416,N_5974,N_7549);
nor U10417 (N_10417,N_9585,N_6242);
nor U10418 (N_10418,N_7843,N_5432);
or U10419 (N_10419,N_6724,N_5487);
xor U10420 (N_10420,N_9841,N_8328);
xnor U10421 (N_10421,N_7376,N_6204);
xor U10422 (N_10422,N_9794,N_7067);
and U10423 (N_10423,N_9539,N_8975);
and U10424 (N_10424,N_9307,N_8476);
or U10425 (N_10425,N_5911,N_8845);
xnor U10426 (N_10426,N_5040,N_9413);
nor U10427 (N_10427,N_9106,N_7161);
or U10428 (N_10428,N_5839,N_7455);
xnor U10429 (N_10429,N_9410,N_8388);
nand U10430 (N_10430,N_7760,N_7952);
and U10431 (N_10431,N_7727,N_9990);
xor U10432 (N_10432,N_8294,N_8536);
nor U10433 (N_10433,N_9099,N_8905);
or U10434 (N_10434,N_6581,N_6964);
nor U10435 (N_10435,N_9685,N_9589);
nand U10436 (N_10436,N_8155,N_7758);
xor U10437 (N_10437,N_7465,N_8774);
nand U10438 (N_10438,N_7341,N_6557);
nor U10439 (N_10439,N_9866,N_6285);
nor U10440 (N_10440,N_9172,N_6360);
nand U10441 (N_10441,N_9522,N_8543);
nor U10442 (N_10442,N_8568,N_5845);
xnor U10443 (N_10443,N_6808,N_6534);
nand U10444 (N_10444,N_7360,N_5938);
or U10445 (N_10445,N_5780,N_9215);
nand U10446 (N_10446,N_7522,N_9022);
xnor U10447 (N_10447,N_9580,N_9334);
and U10448 (N_10448,N_6341,N_5219);
and U10449 (N_10449,N_5045,N_6888);
and U10450 (N_10450,N_8701,N_6151);
xnor U10451 (N_10451,N_5576,N_6001);
xor U10452 (N_10452,N_5319,N_5232);
nor U10453 (N_10453,N_7865,N_6179);
and U10454 (N_10454,N_7524,N_8638);
nand U10455 (N_10455,N_7585,N_9959);
and U10456 (N_10456,N_6533,N_8410);
xnor U10457 (N_10457,N_7487,N_6650);
and U10458 (N_10458,N_7570,N_8127);
and U10459 (N_10459,N_7786,N_8823);
xnor U10460 (N_10460,N_9966,N_9453);
nand U10461 (N_10461,N_6085,N_9159);
nand U10462 (N_10462,N_5094,N_9226);
and U10463 (N_10463,N_6810,N_8888);
and U10464 (N_10464,N_5365,N_6812);
and U10465 (N_10465,N_7265,N_9687);
xnor U10466 (N_10466,N_8865,N_5416);
or U10467 (N_10467,N_7482,N_9285);
or U10468 (N_10468,N_9584,N_7031);
and U10469 (N_10469,N_7636,N_8172);
and U10470 (N_10470,N_7233,N_7507);
xor U10471 (N_10471,N_9394,N_5458);
or U10472 (N_10472,N_7762,N_7620);
xor U10473 (N_10473,N_5741,N_5738);
and U10474 (N_10474,N_5101,N_5947);
xnor U10475 (N_10475,N_7060,N_6434);
and U10476 (N_10476,N_5283,N_5612);
nand U10477 (N_10477,N_5395,N_7733);
nor U10478 (N_10478,N_8392,N_7361);
and U10479 (N_10479,N_9122,N_5923);
xnor U10480 (N_10480,N_9509,N_6856);
and U10481 (N_10481,N_6702,N_8673);
nor U10482 (N_10482,N_6148,N_8512);
nor U10483 (N_10483,N_7788,N_6877);
nand U10484 (N_10484,N_5726,N_7997);
nor U10485 (N_10485,N_5424,N_8720);
xor U10486 (N_10486,N_6974,N_7453);
or U10487 (N_10487,N_6235,N_7687);
nor U10488 (N_10488,N_5639,N_7539);
and U10489 (N_10489,N_9344,N_6922);
xor U10490 (N_10490,N_5282,N_8201);
or U10491 (N_10491,N_7826,N_7664);
and U10492 (N_10492,N_6052,N_7095);
and U10493 (N_10493,N_6700,N_6353);
nor U10494 (N_10494,N_6463,N_8622);
nor U10495 (N_10495,N_7630,N_5596);
nand U10496 (N_10496,N_8719,N_8870);
or U10497 (N_10497,N_9467,N_9108);
nor U10498 (N_10498,N_5132,N_6732);
nor U10499 (N_10499,N_8947,N_7704);
xor U10500 (N_10500,N_9803,N_7540);
nor U10501 (N_10501,N_6744,N_9858);
and U10502 (N_10502,N_5724,N_6278);
nand U10503 (N_10503,N_8991,N_8215);
and U10504 (N_10504,N_6270,N_9253);
xor U10505 (N_10505,N_8707,N_8356);
and U10506 (N_10506,N_7089,N_6710);
xnor U10507 (N_10507,N_9722,N_9507);
and U10508 (N_10508,N_5103,N_9899);
and U10509 (N_10509,N_5110,N_7446);
or U10510 (N_10510,N_9324,N_6531);
and U10511 (N_10511,N_9564,N_5315);
nand U10512 (N_10512,N_6768,N_6494);
and U10513 (N_10513,N_8513,N_6938);
or U10514 (N_10514,N_6785,N_7841);
or U10515 (N_10515,N_6407,N_7744);
nand U10516 (N_10516,N_7651,N_6615);
nor U10517 (N_10517,N_5425,N_9531);
and U10518 (N_10518,N_5159,N_9301);
or U10519 (N_10519,N_7560,N_5787);
xor U10520 (N_10520,N_5992,N_5543);
nor U10521 (N_10521,N_7342,N_5746);
and U10522 (N_10522,N_5464,N_5873);
nor U10523 (N_10523,N_7404,N_5860);
nor U10524 (N_10524,N_5985,N_6067);
or U10525 (N_10525,N_8458,N_5882);
nor U10526 (N_10526,N_6437,N_6846);
xor U10527 (N_10527,N_6918,N_6936);
nor U10528 (N_10528,N_7797,N_6417);
nor U10529 (N_10529,N_7362,N_8345);
or U10530 (N_10530,N_5489,N_8254);
and U10531 (N_10531,N_6713,N_5618);
nor U10532 (N_10532,N_8786,N_6796);
nand U10533 (N_10533,N_9922,N_7793);
xor U10534 (N_10534,N_9611,N_5864);
nor U10535 (N_10535,N_7472,N_5681);
and U10536 (N_10536,N_7972,N_7391);
and U10537 (N_10537,N_6138,N_7218);
or U10538 (N_10538,N_7815,N_6741);
nand U10539 (N_10539,N_9244,N_9848);
nand U10540 (N_10540,N_5093,N_9437);
and U10541 (N_10541,N_5377,N_7219);
and U10542 (N_10542,N_9763,N_7421);
or U10543 (N_10543,N_9526,N_5427);
or U10544 (N_10544,N_6329,N_6891);
or U10545 (N_10545,N_7629,N_5682);
nor U10546 (N_10546,N_7037,N_5910);
nand U10547 (N_10547,N_5297,N_6793);
or U10548 (N_10548,N_5248,N_5874);
nor U10549 (N_10549,N_8945,N_7476);
xnor U10550 (N_10550,N_8725,N_9418);
nand U10551 (N_10551,N_5185,N_6749);
xnor U10552 (N_10552,N_5530,N_9748);
nand U10553 (N_10553,N_9398,N_7548);
xnor U10554 (N_10554,N_6429,N_5354);
or U10555 (N_10555,N_9613,N_9212);
xnor U10556 (N_10556,N_8475,N_5823);
nand U10557 (N_10557,N_8925,N_7184);
nand U10558 (N_10558,N_6839,N_6300);
nor U10559 (N_10559,N_6336,N_5028);
xor U10560 (N_10560,N_7690,N_9931);
or U10561 (N_10561,N_9486,N_9735);
nor U10562 (N_10562,N_6861,N_5908);
or U10563 (N_10563,N_7554,N_6950);
xor U10564 (N_10564,N_5240,N_7681);
nand U10565 (N_10565,N_9040,N_6461);
nand U10566 (N_10566,N_9532,N_5848);
xnor U10567 (N_10567,N_6667,N_9447);
xnor U10568 (N_10568,N_6332,N_9134);
or U10569 (N_10569,N_9988,N_6221);
or U10570 (N_10570,N_8346,N_8076);
xor U10571 (N_10571,N_6144,N_8678);
xnor U10572 (N_10572,N_6789,N_7795);
and U10573 (N_10573,N_6009,N_9428);
xnor U10574 (N_10574,N_8350,N_6672);
nor U10575 (N_10575,N_6133,N_9913);
nand U10576 (N_10576,N_7886,N_6441);
nor U10577 (N_10577,N_5890,N_6855);
or U10578 (N_10578,N_6321,N_8113);
nor U10579 (N_10579,N_7523,N_5324);
and U10580 (N_10580,N_9461,N_6873);
nand U10581 (N_10581,N_6462,N_6325);
nand U10582 (N_10582,N_9760,N_6293);
and U10583 (N_10583,N_8533,N_7495);
xnor U10584 (N_10584,N_9621,N_7989);
nor U10585 (N_10585,N_5528,N_8537);
or U10586 (N_10586,N_9658,N_7306);
xnor U10587 (N_10587,N_6645,N_8531);
nand U10588 (N_10588,N_6025,N_9296);
and U10589 (N_10589,N_5251,N_8941);
and U10590 (N_10590,N_5686,N_8781);
nand U10591 (N_10591,N_7354,N_5397);
or U10592 (N_10592,N_7569,N_7769);
nor U10593 (N_10593,N_6633,N_6603);
and U10594 (N_10594,N_9118,N_9143);
nor U10595 (N_10595,N_6638,N_6804);
nand U10596 (N_10596,N_8082,N_7496);
or U10597 (N_10597,N_6522,N_8360);
or U10598 (N_10598,N_8316,N_7017);
nand U10599 (N_10599,N_9853,N_6921);
xor U10600 (N_10600,N_5855,N_9738);
xor U10601 (N_10601,N_6377,N_6677);
nor U10602 (N_10602,N_8872,N_9112);
or U10603 (N_10603,N_8875,N_8608);
xnor U10604 (N_10604,N_8149,N_6042);
nand U10605 (N_10605,N_9294,N_5488);
and U10606 (N_10606,N_9035,N_5982);
and U10607 (N_10607,N_8832,N_9033);
nor U10608 (N_10608,N_7616,N_9047);
nand U10609 (N_10609,N_9786,N_7903);
nand U10610 (N_10610,N_6874,N_9312);
nor U10611 (N_10611,N_9434,N_8404);
or U10612 (N_10612,N_7021,N_6662);
or U10613 (N_10613,N_6647,N_6352);
nor U10614 (N_10614,N_9221,N_8417);
xnor U10615 (N_10615,N_9961,N_9894);
and U10616 (N_10616,N_5629,N_8665);
xor U10617 (N_10617,N_6772,N_8324);
and U10618 (N_10618,N_6255,N_6245);
or U10619 (N_10619,N_8596,N_5482);
xor U10620 (N_10620,N_6545,N_7096);
and U10621 (N_10621,N_6059,N_9463);
nand U10622 (N_10622,N_5106,N_6814);
xnor U10623 (N_10623,N_8121,N_5086);
nand U10624 (N_10624,N_8973,N_6591);
nand U10625 (N_10625,N_8972,N_7930);
and U10626 (N_10626,N_9726,N_6121);
nand U10627 (N_10627,N_6096,N_6637);
xnor U10628 (N_10628,N_5995,N_5342);
xor U10629 (N_10629,N_9572,N_8853);
nor U10630 (N_10630,N_9617,N_5415);
or U10631 (N_10631,N_9755,N_5870);
and U10632 (N_10632,N_8198,N_9341);
xor U10633 (N_10633,N_5552,N_9528);
and U10634 (N_10634,N_8028,N_5984);
nand U10635 (N_10635,N_7284,N_8712);
or U10636 (N_10636,N_7591,N_5520);
nand U10637 (N_10637,N_6194,N_7106);
nand U10638 (N_10638,N_8427,N_6697);
xor U10639 (N_10639,N_5993,N_5406);
nor U10640 (N_10640,N_7202,N_5881);
and U10641 (N_10641,N_7491,N_8027);
nor U10642 (N_10642,N_8072,N_6284);
or U10643 (N_10643,N_5959,N_7438);
nor U10644 (N_10644,N_7909,N_9056);
nor U10645 (N_10645,N_9092,N_7200);
or U10646 (N_10646,N_5796,N_9559);
and U10647 (N_10647,N_7653,N_9009);
and U10648 (N_10648,N_6586,N_5389);
nor U10649 (N_10649,N_9672,N_8938);
xor U10650 (N_10650,N_5770,N_8453);
xor U10651 (N_10651,N_8093,N_6538);
xnor U10652 (N_10652,N_8080,N_8505);
and U10653 (N_10653,N_8077,N_9042);
nor U10654 (N_10654,N_5934,N_5608);
or U10655 (N_10655,N_7559,N_7771);
xor U10656 (N_10656,N_7953,N_5085);
nor U10657 (N_10657,N_5657,N_9769);
xor U10658 (N_10658,N_8798,N_8249);
xnor U10659 (N_10659,N_5334,N_6406);
and U10660 (N_10660,N_9812,N_8811);
xnor U10661 (N_10661,N_8932,N_9003);
nor U10662 (N_10662,N_5294,N_5049);
xor U10663 (N_10663,N_8809,N_5473);
nor U10664 (N_10664,N_6400,N_9469);
and U10665 (N_10665,N_9133,N_5950);
or U10666 (N_10666,N_6142,N_7649);
or U10667 (N_10667,N_6689,N_6769);
nor U10668 (N_10668,N_5000,N_5564);
xnor U10669 (N_10669,N_5529,N_7738);
nand U10670 (N_10670,N_8545,N_6526);
xor U10671 (N_10671,N_5601,N_6442);
and U10672 (N_10672,N_9494,N_6559);
xnor U10673 (N_10673,N_6641,N_5663);
nand U10674 (N_10674,N_7853,N_6592);
xnor U10675 (N_10675,N_7047,N_9462);
nor U10676 (N_10676,N_8041,N_5477);
xor U10677 (N_10677,N_8351,N_8921);
or U10678 (N_10678,N_7094,N_5500);
nand U10679 (N_10679,N_8134,N_7274);
nand U10680 (N_10680,N_7093,N_6906);
nor U10681 (N_10681,N_5321,N_9947);
nor U10682 (N_10682,N_7724,N_5069);
nor U10683 (N_10683,N_5918,N_5151);
nor U10684 (N_10684,N_6975,N_6946);
nor U10685 (N_10685,N_6467,N_9659);
or U10686 (N_10686,N_8705,N_7914);
and U10687 (N_10687,N_7092,N_8373);
nand U10688 (N_10688,N_8022,N_8331);
nand U10689 (N_10689,N_5480,N_5284);
nand U10690 (N_10690,N_8501,N_9750);
xnor U10691 (N_10691,N_6383,N_7439);
nand U10692 (N_10692,N_8243,N_8769);
nand U10693 (N_10693,N_7116,N_7077);
xnor U10694 (N_10694,N_5971,N_8886);
xnor U10695 (N_10695,N_9751,N_7182);
and U10696 (N_10696,N_8486,N_8036);
nor U10697 (N_10697,N_5958,N_8054);
and U10698 (N_10698,N_8367,N_5502);
xor U10699 (N_10699,N_5295,N_5173);
xnor U10700 (N_10700,N_6018,N_5837);
or U10701 (N_10701,N_9905,N_6095);
nand U10702 (N_10702,N_9362,N_6327);
nor U10703 (N_10703,N_5816,N_5904);
and U10704 (N_10704,N_6805,N_8049);
and U10705 (N_10705,N_9480,N_8498);
xnor U10706 (N_10706,N_7614,N_7848);
nand U10707 (N_10707,N_7799,N_6374);
nor U10708 (N_10708,N_9282,N_6809);
nand U10709 (N_10709,N_7198,N_6903);
and U10710 (N_10710,N_9820,N_8758);
and U10711 (N_10711,N_9830,N_7105);
or U10712 (N_10712,N_5754,N_9648);
and U10713 (N_10713,N_9098,N_7488);
or U10714 (N_10714,N_9889,N_9839);
or U10715 (N_10715,N_9665,N_5651);
xnor U10716 (N_10716,N_9504,N_9471);
and U10717 (N_10717,N_9291,N_9348);
nor U10718 (N_10718,N_9881,N_9872);
and U10719 (N_10719,N_5579,N_8824);
nor U10720 (N_10720,N_7993,N_6552);
xnor U10721 (N_10721,N_8004,N_6825);
nand U10722 (N_10722,N_8557,N_6146);
and U10723 (N_10723,N_7774,N_8829);
xnor U10724 (N_10724,N_5690,N_9956);
and U10725 (N_10725,N_8320,N_9129);
and U10726 (N_10726,N_5022,N_9198);
xor U10727 (N_10727,N_7752,N_7710);
or U10728 (N_10728,N_7108,N_5052);
nor U10729 (N_10729,N_5134,N_8098);
or U10730 (N_10730,N_6453,N_7995);
nand U10731 (N_10731,N_8869,N_5174);
and U10732 (N_10732,N_5357,N_7588);
nand U10733 (N_10733,N_5197,N_5120);
or U10734 (N_10734,N_9996,N_9340);
nand U10735 (N_10735,N_7638,N_5340);
or U10736 (N_10736,N_9237,N_7426);
nor U10737 (N_10737,N_8817,N_8590);
xor U10738 (N_10738,N_9372,N_7647);
or U10739 (N_10739,N_5238,N_8090);
and U10740 (N_10740,N_6726,N_7313);
nor U10741 (N_10741,N_6800,N_5186);
or U10742 (N_10742,N_6475,N_7742);
nand U10743 (N_10743,N_7862,N_9201);
and U10744 (N_10744,N_7725,N_5511);
nor U10745 (N_10745,N_7000,N_8180);
nand U10746 (N_10746,N_9303,N_5274);
and U10747 (N_10747,N_6403,N_6998);
nor U10748 (N_10748,N_7935,N_9014);
or U10749 (N_10749,N_5100,N_5835);
nor U10750 (N_10750,N_8735,N_8483);
or U10751 (N_10751,N_7163,N_6177);
and U10752 (N_10752,N_8914,N_8743);
nand U10753 (N_10753,N_7086,N_5745);
and U10754 (N_10754,N_9946,N_7828);
or U10755 (N_10755,N_8964,N_6781);
and U10756 (N_10756,N_8363,N_8386);
xor U10757 (N_10757,N_5574,N_5187);
xnor U10758 (N_10758,N_5703,N_9793);
nor U10759 (N_10759,N_8765,N_5443);
nor U10760 (N_10760,N_9158,N_9718);
nor U10761 (N_10761,N_8516,N_8881);
xnor U10762 (N_10762,N_6674,N_7860);
and U10763 (N_10763,N_5674,N_9677);
and U10764 (N_10764,N_9190,N_8762);
xnor U10765 (N_10765,N_9691,N_9917);
and U10766 (N_10766,N_5900,N_7996);
and U10767 (N_10767,N_9935,N_9369);
xor U10768 (N_10768,N_8043,N_5312);
and U10769 (N_10769,N_8446,N_6562);
or U10770 (N_10770,N_6594,N_5691);
or U10771 (N_10771,N_8770,N_9901);
xor U10772 (N_10772,N_7346,N_7009);
nor U10773 (N_10773,N_6272,N_9037);
nor U10774 (N_10774,N_6553,N_9180);
or U10775 (N_10775,N_7587,N_9583);
xnor U10776 (N_10776,N_8662,N_5853);
or U10777 (N_10777,N_7352,N_6032);
xor U10778 (N_10778,N_8776,N_9940);
nor U10779 (N_10779,N_8525,N_8599);
xor U10780 (N_10780,N_5087,N_9055);
nor U10781 (N_10781,N_9698,N_7902);
xnor U10782 (N_10782,N_9558,N_6543);
and U10783 (N_10783,N_6271,N_8584);
nand U10784 (N_10784,N_9483,N_8833);
or U10785 (N_10785,N_6444,N_7906);
nand U10786 (N_10786,N_8397,N_5523);
xor U10787 (N_10787,N_7209,N_8144);
or U10788 (N_10788,N_6778,N_5930);
xor U10789 (N_10789,N_9587,N_7010);
and U10790 (N_10790,N_8398,N_5242);
nand U10791 (N_10791,N_6669,N_9855);
nand U10792 (N_10792,N_7801,N_8467);
and U10793 (N_10793,N_6598,N_8696);
nor U10794 (N_10794,N_6288,N_5130);
and U10795 (N_10795,N_6763,N_9100);
and U10796 (N_10796,N_5535,N_8960);
nor U10797 (N_10797,N_5841,N_5135);
nor U10798 (N_10798,N_9733,N_8954);
and U10799 (N_10799,N_9358,N_8967);
nor U10800 (N_10800,N_5944,N_9781);
nand U10801 (N_10801,N_9602,N_9929);
nor U10802 (N_10802,N_5800,N_7254);
or U10803 (N_10803,N_8677,N_8855);
and U10804 (N_10804,N_9893,N_6275);
nor U10805 (N_10805,N_9731,N_7148);
and U10806 (N_10806,N_9239,N_9863);
nand U10807 (N_10807,N_6521,N_8616);
xnor U10808 (N_10808,N_9274,N_8871);
or U10809 (N_10809,N_5829,N_5356);
and U10810 (N_10810,N_6743,N_8063);
nand U10811 (N_10811,N_5403,N_8177);
and U10812 (N_10812,N_7358,N_5549);
and U10813 (N_10813,N_5433,N_8037);
nand U10814 (N_10814,N_5002,N_6934);
and U10815 (N_10815,N_8009,N_6021);
xor U10816 (N_10816,N_6363,N_8293);
nand U10817 (N_10817,N_7263,N_7960);
nor U10818 (N_10818,N_5202,N_8566);
nand U10819 (N_10819,N_5289,N_5036);
xnor U10820 (N_10820,N_7675,N_6195);
or U10821 (N_10821,N_5653,N_7251);
xor U10822 (N_10822,N_6291,N_7783);
and U10823 (N_10823,N_7423,N_5074);
or U10824 (N_10824,N_9797,N_5842);
or U10825 (N_10825,N_6351,N_5057);
or U10826 (N_10826,N_7505,N_9032);
and U10827 (N_10827,N_5128,N_7613);
or U10828 (N_10828,N_7485,N_9368);
nor U10829 (N_10829,N_6411,N_6127);
and U10830 (N_10830,N_8281,N_8305);
nor U10831 (N_10831,N_7922,N_9717);
nand U10832 (N_10832,N_7660,N_7889);
nand U10833 (N_10833,N_8141,N_5401);
xnor U10834 (N_10834,N_7065,N_9278);
xor U10835 (N_10835,N_8992,N_7014);
and U10836 (N_10836,N_9941,N_5526);
or U10837 (N_10837,N_9860,N_9869);
xnor U10838 (N_10838,N_6439,N_9771);
nand U10839 (N_10839,N_7130,N_5771);
xnor U10840 (N_10840,N_6484,N_6578);
xnor U10841 (N_10841,N_7929,N_5584);
nand U10842 (N_10842,N_5105,N_8588);
xor U10843 (N_10843,N_7518,N_5430);
or U10844 (N_10844,N_8511,N_6102);
and U10845 (N_10845,N_5307,N_7288);
nand U10846 (N_10846,N_5372,N_8234);
xor U10847 (N_10847,N_7348,N_8484);
nor U10848 (N_10848,N_8736,N_9936);
nand U10849 (N_10849,N_5352,N_7070);
nand U10850 (N_10850,N_8569,N_7394);
or U10851 (N_10851,N_5907,N_8227);
xnor U10852 (N_10852,N_8658,N_5325);
nand U10853 (N_10853,N_9836,N_8439);
or U10854 (N_10854,N_7273,N_5723);
nor U10855 (N_10855,N_6415,N_9850);
xnor U10856 (N_10856,N_6843,N_5527);
nor U10857 (N_10857,N_9441,N_6074);
xnor U10858 (N_10858,N_7965,N_5280);
xnor U10859 (N_10859,N_8207,N_9651);
nor U10860 (N_10860,N_6359,N_8003);
or U10861 (N_10861,N_6754,N_7318);
or U10862 (N_10862,N_7050,N_9071);
nor U10863 (N_10863,N_7479,N_5798);
and U10864 (N_10864,N_9384,N_5285);
xnor U10865 (N_10865,N_9276,N_5200);
nor U10866 (N_10866,N_9754,N_9927);
and U10867 (N_10867,N_8626,N_8904);
nor U10868 (N_10868,N_7879,N_8858);
nor U10869 (N_10869,N_7149,N_9903);
nor U10870 (N_10870,N_6761,N_9149);
or U10871 (N_10871,N_7927,N_7012);
nor U10872 (N_10872,N_7683,N_6181);
and U10873 (N_10873,N_9861,N_6953);
nand U10874 (N_10874,N_8429,N_9353);
nand U10875 (N_10875,N_5327,N_5296);
nand U10876 (N_10876,N_9113,N_6362);
and U10877 (N_10877,N_9789,N_6389);
xnor U10878 (N_10878,N_8364,N_6296);
nor U10879 (N_10879,N_7018,N_6972);
or U10880 (N_10880,N_5898,N_6450);
nand U10881 (N_10881,N_9895,N_5104);
nor U10882 (N_10882,N_6978,N_7102);
and U10883 (N_10883,N_9573,N_5420);
and U10884 (N_10884,N_7640,N_5760);
nand U10885 (N_10885,N_5298,N_9195);
nor U10886 (N_10886,N_7904,N_9785);
nand U10887 (N_10887,N_6840,N_6948);
xnor U10888 (N_10888,N_7351,N_6046);
and U10889 (N_10889,N_6822,N_7146);
nor U10890 (N_10890,N_6213,N_6474);
or U10891 (N_10891,N_6728,N_5475);
nor U10892 (N_10892,N_8734,N_7475);
nand U10893 (N_10893,N_6820,N_6767);
xnor U10894 (N_10894,N_8067,N_6238);
and U10895 (N_10895,N_9821,N_6850);
or U10896 (N_10896,N_5531,N_8808);
xnor U10897 (N_10897,N_9141,N_6880);
nor U10898 (N_10898,N_8989,N_8241);
or U10899 (N_10899,N_8259,N_6425);
nor U10900 (N_10900,N_8979,N_8873);
xnor U10901 (N_10901,N_6387,N_8843);
or U10902 (N_10902,N_9427,N_9974);
or U10903 (N_10903,N_9411,N_6386);
or U10904 (N_10904,N_7627,N_9747);
nand U10905 (N_10905,N_6639,N_6519);
xor U10906 (N_10906,N_6666,N_9550);
nor U10907 (N_10907,N_7514,N_5092);
nand U10908 (N_10908,N_5090,N_7596);
nand U10909 (N_10909,N_8976,N_5696);
xnor U10910 (N_10910,N_5731,N_8445);
xnor U10911 (N_10911,N_9636,N_8349);
nand U10912 (N_10912,N_8197,N_5933);
nand U10913 (N_10913,N_9481,N_7567);
and U10914 (N_10914,N_9379,N_7392);
nand U10915 (N_10915,N_5048,N_6503);
or U10916 (N_10916,N_9065,N_5809);
nor U10917 (N_10917,N_8186,N_8167);
and U10918 (N_10918,N_5428,N_5625);
and U10919 (N_10919,N_7191,N_8050);
nand U10920 (N_10920,N_9674,N_5026);
nor U10921 (N_10921,N_6422,N_5603);
and U10922 (N_10922,N_7583,N_7589);
xor U10923 (N_10923,N_8210,N_7748);
and U10924 (N_10924,N_8939,N_8183);
nand U10925 (N_10925,N_9257,N_7179);
xnor U10926 (N_10926,N_5239,N_9543);
nand U10927 (N_10927,N_7247,N_8448);
xnor U10928 (N_10928,N_6870,N_7635);
or U10929 (N_10929,N_5269,N_6550);
xor U10930 (N_10930,N_6103,N_5509);
nor U10931 (N_10931,N_8804,N_9095);
xnor U10932 (N_10932,N_6915,N_5901);
and U10933 (N_10933,N_9787,N_9575);
and U10934 (N_10934,N_8691,N_6738);
nor U10935 (N_10935,N_5278,N_7048);
nand U10936 (N_10936,N_5642,N_8936);
nor U10937 (N_10937,N_7419,N_6154);
xnor U10938 (N_10938,N_7780,N_8194);
or U10939 (N_10939,N_6207,N_7007);
xor U10940 (N_10940,N_9874,N_8782);
and U10941 (N_10941,N_8548,N_7557);
nand U10942 (N_10942,N_9019,N_5176);
and U10943 (N_10943,N_9952,N_5533);
xor U10944 (N_10944,N_5457,N_9921);
nor U10945 (N_10945,N_7140,N_7385);
and U10946 (N_10946,N_7053,N_9125);
nand U10947 (N_10947,N_8079,N_6299);
xor U10948 (N_10948,N_6008,N_5075);
nand U10949 (N_10949,N_7178,N_8425);
nand U10950 (N_10950,N_5476,N_7378);
and U10951 (N_10951,N_5078,N_6175);
or U10952 (N_10952,N_8646,N_6385);
or U10953 (N_10953,N_8084,N_9667);
nor U10954 (N_10954,N_6112,N_9381);
xnor U10955 (N_10955,N_6525,N_5264);
xor U10956 (N_10956,N_8828,N_9997);
xor U10957 (N_10957,N_9745,N_6378);
xnor U10958 (N_10958,N_6901,N_6283);
and U10959 (N_10959,N_7737,N_5046);
nor U10960 (N_10960,N_8096,N_9224);
and U10961 (N_10961,N_9741,N_9311);
nand U10962 (N_10962,N_5331,N_5668);
nand U10963 (N_10963,N_7015,N_6664);
and U10964 (N_10964,N_8303,N_6780);
xor U10965 (N_10965,N_5300,N_7987);
nor U10966 (N_10966,N_8274,N_7986);
nor U10967 (N_10967,N_8415,N_7881);
or U10968 (N_10968,N_6671,N_9945);
xor U10969 (N_10969,N_8447,N_6648);
or U10970 (N_10970,N_7213,N_7283);
nand U10971 (N_10971,N_9102,N_8244);
nor U10972 (N_10972,N_6440,N_9060);
and U10973 (N_10973,N_9710,N_5980);
and U10974 (N_10974,N_8385,N_9302);
or U10975 (N_10975,N_5570,N_5721);
or U10976 (N_10976,N_9419,N_7708);
xor U10977 (N_10977,N_9416,N_5508);
nor U10978 (N_10978,N_7668,N_9136);
xnor U10979 (N_10979,N_7040,N_9377);
nor U10980 (N_10980,N_5791,N_8357);
and U10981 (N_10981,N_8394,N_6514);
or U10982 (N_10982,N_6211,N_5205);
and U10983 (N_10983,N_9070,N_8928);
and U10984 (N_10984,N_6502,N_5582);
and U10985 (N_10985,N_8642,N_6483);
nor U10986 (N_10986,N_5568,N_8713);
xor U10987 (N_10987,N_8773,N_5997);
xor U10988 (N_10988,N_6576,N_7430);
xor U10989 (N_10989,N_5700,N_9174);
nand U10990 (N_10990,N_9815,N_8999);
and U10991 (N_10991,N_7436,N_7582);
nor U10992 (N_10992,N_9343,N_9716);
or U10993 (N_10993,N_8455,N_8138);
or U10994 (N_10994,N_9970,N_6186);
xnor U10995 (N_10995,N_7100,N_8465);
xor U10996 (N_10996,N_5353,N_6965);
nand U10997 (N_10997,N_7529,N_6745);
or U10998 (N_10998,N_6836,N_6991);
and U10999 (N_10999,N_7300,N_7110);
and U11000 (N_11000,N_5129,N_8255);
nor U11001 (N_11001,N_5419,N_6160);
and U11002 (N_11002,N_7331,N_5516);
nand U11003 (N_11003,N_7152,N_6129);
and U11004 (N_11004,N_7045,N_7694);
or U11005 (N_11005,N_5080,N_8733);
and U11006 (N_11006,N_6011,N_5329);
or U11007 (N_11007,N_8898,N_7381);
nor U11008 (N_11008,N_7330,N_7946);
nor U11009 (N_11009,N_8799,N_5591);
xor U11010 (N_11010,N_8287,N_7816);
nand U11011 (N_11011,N_7574,N_6999);
and U11012 (N_11012,N_7527,N_7370);
or U11013 (N_11013,N_5849,N_9697);
nor U11014 (N_11014,N_9188,N_9184);
nand U11015 (N_11015,N_9775,N_5698);
and U11016 (N_11016,N_9233,N_5761);
xor U11017 (N_11017,N_7701,N_6124);
and U11018 (N_11018,N_7551,N_9612);
nor U11019 (N_11019,N_5421,N_9675);
nor U11020 (N_11020,N_6807,N_5142);
or U11021 (N_11021,N_7355,N_7516);
and U11022 (N_11022,N_8868,N_7314);
and U11023 (N_11023,N_7261,N_5336);
nor U11024 (N_11024,N_8935,N_9729);
xor U11025 (N_11025,N_7528,N_6831);
nor U11026 (N_11026,N_6217,N_7231);
and U11027 (N_11027,N_8247,N_8061);
xnor U11028 (N_11028,N_7023,N_5774);
or U11029 (N_11029,N_6401,N_8494);
or U11030 (N_11030,N_6670,N_5932);
nor U11031 (N_11031,N_6236,N_9807);
or U11032 (N_11032,N_7427,N_6455);
nand U11033 (N_11033,N_8040,N_9796);
nand U11034 (N_11034,N_5374,N_5228);
or U11035 (N_11035,N_7663,N_7619);
xnor U11036 (N_11036,N_5019,N_5341);
nor U11037 (N_11037,N_5224,N_7535);
or U11038 (N_11038,N_8540,N_7195);
and U11039 (N_11039,N_9938,N_8396);
xor U11040 (N_11040,N_8778,N_8692);
and U11041 (N_11041,N_8613,N_5942);
nand U11042 (N_11042,N_8311,N_5008);
or U11043 (N_11043,N_5194,N_9222);
or U11044 (N_11044,N_8267,N_7532);
nand U11045 (N_11045,N_9380,N_8671);
nand U11046 (N_11046,N_9328,N_6123);
or U11047 (N_11047,N_8108,N_5561);
and U11048 (N_11048,N_9273,N_5465);
nand U11049 (N_11049,N_8990,N_5471);
or U11050 (N_11050,N_8085,N_6920);
and U11051 (N_11051,N_6380,N_7594);
nand U11052 (N_11052,N_6135,N_8802);
or U11053 (N_11053,N_5583,N_7973);
and U11054 (N_11054,N_6490,N_9705);
xor U11055 (N_11055,N_8342,N_6169);
nand U11056 (N_11056,N_8631,N_6982);
xor U11057 (N_11057,N_6478,N_9886);
or U11058 (N_11058,N_7918,N_5014);
and U11059 (N_11059,N_8369,N_7641);
and U11060 (N_11060,N_9650,N_8126);
xor U11061 (N_11061,N_9264,N_8837);
nor U11062 (N_11062,N_8088,N_5201);
xnor U11063 (N_11063,N_6080,N_5042);
and U11064 (N_11064,N_5190,N_7291);
nor U11065 (N_11065,N_5996,N_7656);
xnor U11066 (N_11066,N_6339,N_8706);
xor U11067 (N_11067,N_6216,N_6829);
nand U11068 (N_11068,N_7858,N_5955);
xor U11069 (N_11069,N_9765,N_5497);
and U11070 (N_11070,N_5797,N_5384);
or U11071 (N_11071,N_6541,N_7871);
and U11072 (N_11072,N_7150,N_7131);
and U11073 (N_11073,N_8150,N_5894);
nand U11074 (N_11074,N_5752,N_7759);
nand U11075 (N_11075,N_7180,N_9407);
xnor U11076 (N_11076,N_9502,N_8019);
and U11077 (N_11077,N_8083,N_7174);
or U11078 (N_11078,N_8195,N_7661);
xor U11079 (N_11079,N_6818,N_9479);
xor U11080 (N_11080,N_8577,N_7931);
xor U11081 (N_11081,N_6176,N_9867);
or U11082 (N_11082,N_5767,N_6717);
or U11083 (N_11083,N_5633,N_6277);
or U11084 (N_11084,N_6026,N_7402);
nor U11085 (N_11085,N_9991,N_8958);
nor U11086 (N_11086,N_9080,N_5987);
nand U11087 (N_11087,N_8056,N_7181);
xor U11088 (N_11088,N_9325,N_5779);
or U11089 (N_11089,N_6412,N_8086);
and U11090 (N_11090,N_8387,N_7905);
nand U11091 (N_11091,N_7981,N_8934);
nand U11092 (N_11092,N_6088,N_7547);
or U11093 (N_11093,N_8325,N_5550);
nand U11094 (N_11094,N_8438,N_6323);
nor U11095 (N_11095,N_9782,N_7897);
or U11096 (N_11096,N_6530,N_7160);
xnor U11097 (N_11097,N_5728,N_8656);
or U11098 (N_11098,N_6134,N_8655);
xnor U11099 (N_11099,N_9977,N_5572);
nor U11100 (N_11100,N_6506,N_6826);
xor U11101 (N_11101,N_7123,N_8333);
xor U11102 (N_11102,N_7262,N_8731);
nand U11103 (N_11103,N_8847,N_8221);
xor U11104 (N_11104,N_5606,N_5220);
and U11105 (N_11105,N_5299,N_9474);
or U11106 (N_11106,N_9030,N_5861);
and U11107 (N_11107,N_6518,N_9128);
nor U11108 (N_11108,N_6932,N_6599);
xnor U11109 (N_11109,N_9067,N_7628);
and U11110 (N_11110,N_9393,N_9061);
nor U11111 (N_11111,N_9299,N_8561);
xor U11112 (N_11112,N_5832,N_8790);
nor U11113 (N_11113,N_7043,N_5351);
nor U11114 (N_11114,N_8497,N_7746);
xnor U11115 (N_11115,N_5369,N_5311);
and U11116 (N_11116,N_7506,N_8065);
or U11117 (N_11117,N_8147,N_8559);
xor U11118 (N_11118,N_6342,N_8075);
xor U11119 (N_11119,N_8334,N_6276);
and U11120 (N_11120,N_9779,N_5692);
nand U11121 (N_11121,N_6889,N_6563);
nand U11122 (N_11122,N_7063,N_6959);
or U11123 (N_11123,N_5160,N_7625);
nor U11124 (N_11124,N_7454,N_6602);
nor U11125 (N_11125,N_7844,N_9556);
and U11126 (N_11126,N_8452,N_6607);
xnor U11127 (N_11127,N_9329,N_9939);
nand U11128 (N_11128,N_9835,N_9484);
nor U11129 (N_11129,N_7206,N_9266);
nor U11130 (N_11130,N_6844,N_8347);
nand U11131 (N_11131,N_7884,N_5998);
xor U11132 (N_11132,N_8016,N_8271);
nor U11133 (N_11133,N_8815,N_6611);
xnor U11134 (N_11134,N_5655,N_6695);
xnor U11135 (N_11135,N_9609,N_8604);
nor U11136 (N_11136,N_8206,N_9713);
or U11137 (N_11137,N_8623,N_5275);
xnor U11138 (N_11138,N_9912,N_9630);
xnor U11139 (N_11139,N_8422,N_6333);
or U11140 (N_11140,N_8563,N_9027);
and U11141 (N_11141,N_7893,N_5431);
or U11142 (N_11142,N_6517,N_8042);
nor U11143 (N_11143,N_5367,N_6837);
nor U11144 (N_11144,N_6631,N_5679);
nor U11145 (N_11145,N_5649,N_7266);
or U11146 (N_11146,N_7278,N_9197);
or U11147 (N_11147,N_9567,N_7717);
and U11148 (N_11148,N_5578,N_8269);
nand U11149 (N_11149,N_6865,N_8377);
or U11150 (N_11150,N_6753,N_5229);
or U11151 (N_11151,N_6565,N_7432);
xnor U11152 (N_11152,N_6875,N_7969);
and U11153 (N_11153,N_9801,N_6232);
or U11154 (N_11154,N_6787,N_7141);
nand U11155 (N_11155,N_5807,N_9944);
xor U11156 (N_11156,N_7407,N_7728);
nand U11157 (N_11157,N_7655,N_8487);
nor U11158 (N_11158,N_9525,N_7172);
or U11159 (N_11159,N_6384,N_9565);
xnor U11160 (N_11160,N_9683,N_7612);
nand U11161 (N_11161,N_7199,N_8414);
nand U11162 (N_11162,N_7119,N_9271);
and U11163 (N_11163,N_5747,N_6905);
nor U11164 (N_11164,N_5043,N_7349);
nor U11165 (N_11165,N_9476,N_9631);
or U11166 (N_11166,N_8589,N_6979);
or U11167 (N_11167,N_5759,N_9623);
nor U11168 (N_11168,N_6198,N_6064);
nor U11169 (N_11169,N_5073,N_7985);
or U11170 (N_11170,N_5792,N_7503);
nand U11171 (N_11171,N_6189,N_9314);
nand U11172 (N_11172,N_7153,N_9167);
xor U11173 (N_11173,N_7236,N_9681);
and U11174 (N_11174,N_7145,N_9610);
nand U11175 (N_11175,N_8156,N_5010);
nor U11176 (N_11176,N_5138,N_7035);
nand U11177 (N_11177,N_5519,N_5279);
and U11178 (N_11178,N_6547,N_9616);
or U11179 (N_11179,N_6540,N_7246);
xnor U11180 (N_11180,N_5922,N_8101);
nor U11181 (N_11181,N_9818,N_5521);
xnor U11182 (N_11182,N_7992,N_6346);
or U11183 (N_11183,N_6125,N_9044);
nor U11184 (N_11184,N_5316,N_7497);
and U11185 (N_11185,N_7915,N_6060);
or U11186 (N_11186,N_8502,N_6655);
or U11187 (N_11187,N_7894,N_9942);
nand U11188 (N_11188,N_8089,N_6433);
nor U11189 (N_11189,N_8292,N_6912);
or U11190 (N_11190,N_8433,N_7327);
nand U11191 (N_11191,N_5802,N_5869);
nand U11192 (N_11192,N_8515,N_5303);
xor U11193 (N_11193,N_8340,N_6030);
and U11194 (N_11194,N_9967,N_5799);
nand U11195 (N_11195,N_9396,N_6017);
nand U11196 (N_11196,N_6848,N_8005);
or U11197 (N_11197,N_9347,N_7509);
nand U11198 (N_11198,N_8242,N_8924);
and U11199 (N_11199,N_8793,N_5945);
xnor U11200 (N_11200,N_7755,N_8007);
or U11201 (N_11201,N_6083,N_9438);
and U11202 (N_11202,N_5643,N_8091);
and U11203 (N_11203,N_8555,N_5820);
nand U11204 (N_11204,N_8551,N_9452);
and U11205 (N_11205,N_9715,N_6010);
nor U11206 (N_11206,N_6364,N_8754);
and U11207 (N_11207,N_8276,N_7870);
or U11208 (N_11208,N_6962,N_9795);
nor U11209 (N_11209,N_7712,N_8789);
or U11210 (N_11210,N_6315,N_6863);
nand U11211 (N_11211,N_8672,N_6824);
nand U11212 (N_11212,N_6485,N_9117);
xor U11213 (N_11213,N_7230,N_5323);
or U11214 (N_11214,N_8755,N_6908);
and U11215 (N_11215,N_9520,N_5373);
or U11216 (N_11216,N_7833,N_5016);
or U11217 (N_11217,N_9888,N_9231);
xor U11218 (N_11218,N_6699,N_9928);
or U11219 (N_11219,N_7428,N_5137);
nor U11220 (N_11220,N_9139,N_6990);
or U11221 (N_11221,N_5166,N_7369);
xnor U11222 (N_11222,N_8193,N_6955);
or U11223 (N_11223,N_5750,N_9963);
or U11224 (N_11224,N_8851,N_7210);
or U11225 (N_11225,N_5970,N_7773);
and U11226 (N_11226,N_8199,N_5462);
and U11227 (N_11227,N_6152,N_7669);
and U11228 (N_11228,N_5271,N_6720);
or U11229 (N_11229,N_7221,N_9433);
and U11230 (N_11230,N_5231,N_8969);
nand U11231 (N_11231,N_7751,N_8477);
nor U11232 (N_11232,N_8166,N_7513);
and U11233 (N_11233,N_6679,N_5852);
xor U11234 (N_11234,N_8891,N_9766);
nor U11235 (N_11235,N_9477,N_9131);
or U11236 (N_11236,N_8961,N_7339);
and U11237 (N_11237,N_5123,N_7442);
or U11238 (N_11238,N_8650,N_6073);
and U11239 (N_11239,N_6676,N_9356);
nand U11240 (N_11240,N_6015,N_5082);
and U11241 (N_11241,N_9170,N_5102);
nor U11242 (N_11242,N_9138,N_8235);
nor U11243 (N_11243,N_8576,N_6706);
xnor U11244 (N_11244,N_8393,N_5586);
or U11245 (N_11245,N_6044,N_7597);
xor U11246 (N_11246,N_5964,N_6394);
and U11247 (N_11247,N_5951,N_6945);
xnor U11248 (N_11248,N_8884,N_5383);
nor U11249 (N_11249,N_7714,N_5784);
or U11250 (N_11250,N_9132,N_5163);
nor U11251 (N_11251,N_8698,N_9742);
nor U11252 (N_11252,N_8246,N_6819);
nand U11253 (N_11253,N_5459,N_7700);
nor U11254 (N_11254,N_8820,N_8024);
xnor U11255 (N_11255,N_7309,N_6190);
or U11256 (N_11256,N_5554,N_6723);
xnor U11257 (N_11257,N_8683,N_6072);
xnor U11258 (N_11258,N_8950,N_6465);
or U11259 (N_11259,N_9466,N_8669);
nor U11260 (N_11260,N_7874,N_7481);
xnor U11261 (N_11261,N_6486,N_7375);
xnor U11262 (N_11262,N_6432,N_8443);
nor U11263 (N_11263,N_7639,N_9386);
nand U11264 (N_11264,N_8407,N_8020);
and U11265 (N_11265,N_8826,N_7731);
nor U11266 (N_11266,N_9625,N_8783);
and U11267 (N_11267,N_8575,N_8801);
and U11268 (N_11268,N_5267,N_7158);
nand U11269 (N_11269,N_9026,N_8416);
xor U11270 (N_11270,N_8109,N_9828);
nor U11271 (N_11271,N_8361,N_6897);
or U11272 (N_11272,N_6813,N_7308);
or U11273 (N_11273,N_5671,N_8132);
and U11274 (N_11274,N_7526,N_6900);
nand U11275 (N_11275,N_5805,N_7610);
xnor U11276 (N_11276,N_5546,N_9000);
or U11277 (N_11277,N_5604,N_7242);
xor U11278 (N_11278,N_7855,N_6898);
nor U11279 (N_11279,N_6356,N_6851);
and U11280 (N_11280,N_7061,N_6050);
or U11281 (N_11281,N_5333,N_6280);
nand U11282 (N_11282,N_5856,N_5916);
or U11283 (N_11283,N_6106,N_6038);
and U11284 (N_11284,N_6132,N_9005);
nand U11285 (N_11285,N_8812,N_9798);
nor U11286 (N_11286,N_8032,N_8757);
and U11287 (N_11287,N_9045,N_5380);
nor U11288 (N_11288,N_6773,N_7374);
nand U11289 (N_11289,N_9043,N_6168);
xnor U11290 (N_11290,N_5786,N_6684);
nor U11291 (N_11291,N_5115,N_5571);
nand U11292 (N_11292,N_5246,N_7899);
nor U11293 (N_11293,N_9010,N_6000);
nand U11294 (N_11294,N_8676,N_8441);
nand U11295 (N_11295,N_5484,N_7888);
and U11296 (N_11296,N_6718,N_9768);
nor U11297 (N_11297,N_7367,N_9757);
nor U11298 (N_11298,N_8165,N_6971);
nand U11299 (N_11299,N_7382,N_7003);
xor U11300 (N_11300,N_9039,N_9833);
or U11301 (N_11301,N_9620,N_6766);
and U11302 (N_11302,N_9854,N_9306);
nor U11303 (N_11303,N_5887,N_8640);
xor U11304 (N_11304,N_5906,N_5708);
and U11305 (N_11305,N_9614,N_6750);
and U11306 (N_11306,N_5658,N_9297);
nor U11307 (N_11307,N_6926,N_9626);
nand U11308 (N_11308,N_6941,N_6043);
xnor U11309 (N_11309,N_9799,N_8107);
and U11310 (N_11310,N_9727,N_8595);
nor U11311 (N_11311,N_6866,N_8772);
and U11312 (N_11312,N_7042,N_6065);
nor U11313 (N_11313,N_6493,N_7556);
xnor U11314 (N_11314,N_9924,N_6508);
xor U11315 (N_11315,N_9236,N_6847);
nand U11316 (N_11316,N_9510,N_9397);
and U11317 (N_11317,N_8690,N_6675);
and U11318 (N_11318,N_5017,N_8062);
and U11319 (N_11319,N_9391,N_6020);
and U11320 (N_11320,N_8160,N_5426);
and U11321 (N_11321,N_7418,N_6397);
nor U11322 (N_11322,N_9444,N_6997);
nor U11323 (N_11323,N_7673,N_8124);
and U11324 (N_11324,N_8988,N_8440);
and U11325 (N_11325,N_6310,N_8978);
and U11326 (N_11326,N_5534,N_7136);
nand U11327 (N_11327,N_8560,N_7764);
xor U11328 (N_11328,N_8485,N_7812);
nand U11329 (N_11329,N_7787,N_8933);
xnor U11330 (N_11330,N_7800,N_9740);
nand U11331 (N_11331,N_9951,N_7316);
nand U11332 (N_11332,N_5359,N_5893);
nand U11333 (N_11333,N_7388,N_6774);
xor U11334 (N_11334,N_9468,N_8348);
nand U11335 (N_11335,N_7835,N_8984);
xnor U11336 (N_11336,N_9934,N_9911);
and U11337 (N_11337,N_8099,N_8835);
nor U11338 (N_11338,N_8687,N_8694);
xor U11339 (N_11339,N_7165,N_7353);
nor U11340 (N_11340,N_9091,N_6261);
nor U11341 (N_11341,N_5687,N_8571);
or U11342 (N_11342,N_7033,N_6092);
nor U11343 (N_11343,N_5081,N_6294);
nand U11344 (N_11344,N_5695,N_5227);
xnor U11345 (N_11345,N_6913,N_6094);
nand U11346 (N_11346,N_9900,N_7607);
nor U11347 (N_11347,N_6062,N_6402);
and U11348 (N_11348,N_6806,N_8395);
nand U11349 (N_11349,N_6078,N_5920);
nor U11350 (N_11350,N_5735,N_6686);
xor U11351 (N_11351,N_6457,N_6464);
and U11352 (N_11352,N_8806,N_5766);
nor U11353 (N_11353,N_9643,N_8251);
and U11354 (N_11354,N_6958,N_9432);
or U11355 (N_11355,N_9506,N_6696);
xor U11356 (N_11356,N_9290,N_8482);
and U11357 (N_11357,N_7380,N_7249);
nor U11358 (N_11358,N_8384,N_5928);
and U11359 (N_11359,N_8753,N_7676);
xnor U11360 (N_11360,N_8730,N_7814);
xnor U11361 (N_11361,N_6233,N_7940);
nand U11362 (N_11362,N_5917,N_8317);
nor U11363 (N_11363,N_7890,N_7564);
nand U11364 (N_11364,N_5895,N_7873);
and U11365 (N_11365,N_5391,N_7344);
xor U11366 (N_11366,N_7602,N_5715);
or U11367 (N_11367,N_6077,N_8095);
nor U11368 (N_11368,N_9156,N_7098);
or U11369 (N_11369,N_8302,N_8163);
xor U11370 (N_11370,N_7445,N_7919);
nand U11371 (N_11371,N_8970,N_5598);
nand U11372 (N_11372,N_9265,N_9331);
nor U11373 (N_11373,N_6481,N_8944);
and U11374 (N_11374,N_9443,N_7248);
xor U11375 (N_11375,N_9446,N_6577);
or U11376 (N_11376,N_9023,N_5662);
xnor U11377 (N_11377,N_5079,N_5701);
and U11378 (N_11378,N_5790,N_9058);
xnor U11379 (N_11379,N_9679,N_7373);
nand U11380 (N_11380,N_5322,N_5967);
or U11381 (N_11381,N_8624,N_8968);
nor U11382 (N_11382,N_5563,N_7703);
nand U11383 (N_11383,N_8131,N_9498);
or U11384 (N_11384,N_9200,N_7568);
or U11385 (N_11385,N_9414,N_8013);
nor U11386 (N_11386,N_8300,N_8100);
nor U11387 (N_11387,N_6747,N_8895);
and U11388 (N_11388,N_8539,N_9370);
or U11389 (N_11389,N_5254,N_9004);
nand U11390 (N_11390,N_5020,N_7448);
or U11391 (N_11391,N_8344,N_5919);
nand U11392 (N_11392,N_8110,N_9708);
nand U11393 (N_11393,N_5125,N_8670);
and U11394 (N_11394,N_5024,N_6392);
nor U11395 (N_11395,N_8862,N_7335);
and U11396 (N_11396,N_5631,N_8704);
xnor U11397 (N_11397,N_7363,N_8097);
xor U11398 (N_11398,N_9326,N_7898);
and U11399 (N_11399,N_9417,N_9862);
or U11400 (N_11400,N_7143,N_6680);
and U11401 (N_11401,N_8639,N_9649);
xor U11402 (N_11402,N_9639,N_6107);
nor U11403 (N_11403,N_5678,N_8204);
xor U11404 (N_11404,N_8405,N_8819);
xor U11405 (N_11405,N_7734,N_5446);
or U11406 (N_11406,N_7747,N_7954);
and U11407 (N_11407,N_5015,N_7711);
or U11408 (N_11408,N_5449,N_5172);
and U11409 (N_11409,N_5363,N_6307);
or U11410 (N_11410,N_6748,N_6801);
or U11411 (N_11411,N_8228,N_9844);
or U11412 (N_11412,N_6055,N_6708);
or U11413 (N_11413,N_7478,N_9603);
xnor U11414 (N_11414,N_5378,N_5595);
nand U11415 (N_11415,N_5054,N_6201);
nor U11416 (N_11416,N_9849,N_6141);
nor U11417 (N_11417,N_6703,N_5165);
nor U11418 (N_11418,N_8962,N_9788);
or U11419 (N_11419,N_7321,N_8035);
xor U11420 (N_11420,N_6896,N_9436);
and U11421 (N_11421,N_5704,N_6987);
and U11422 (N_11422,N_8549,N_5857);
or U11423 (N_11423,N_8618,N_7433);
xor U11424 (N_11424,N_7285,N_9392);
xor U11425 (N_11425,N_5925,N_8627);
nand U11426 (N_11426,N_7269,N_5941);
nor U11427 (N_11427,N_6986,N_8739);
nand U11428 (N_11428,N_5493,N_9424);
nor U11429 (N_11429,N_7099,N_9096);
or U11430 (N_11430,N_6037,N_5233);
and U11431 (N_11431,N_9548,N_7572);
nand U11432 (N_11432,N_8908,N_7775);
xor U11433 (N_11433,N_9187,N_9066);
and U11434 (N_11434,N_7750,N_7416);
nand U11435 (N_11435,N_7466,N_6473);
nand U11436 (N_11436,N_5935,N_8504);
or U11437 (N_11437,N_7796,N_6223);
nand U11438 (N_11438,N_9059,N_7398);
nor U11439 (N_11439,N_9024,N_5884);
or U11440 (N_11440,N_9756,N_5977);
nor U11441 (N_11441,N_6496,N_7695);
nand U11442 (N_11442,N_9544,N_6164);
and U11443 (N_11443,N_8464,N_5862);
or U11444 (N_11444,N_6274,N_8648);
nor U11445 (N_11445,N_5693,N_8717);
nor U11446 (N_11446,N_8532,N_9130);
xnor U11447 (N_11447,N_7706,N_9725);
xor U11448 (N_11448,N_7637,N_7293);
nand U11449 (N_11449,N_5491,N_8223);
and U11450 (N_11450,N_8225,N_8602);
and U11451 (N_11451,N_9555,N_5058);
and U11452 (N_11452,N_5725,N_6118);
nor U11453 (N_11453,N_9980,N_8278);
xor U11454 (N_11454,N_7976,N_8749);
xor U11455 (N_11455,N_8336,N_7356);
xor U11456 (N_11456,N_7477,N_6418);
xnor U11457 (N_11457,N_5600,N_7580);
nand U11458 (N_11458,N_7234,N_9011);
and U11459 (N_11459,N_7575,N_8890);
or U11460 (N_11460,N_7593,N_6254);
and U11461 (N_11461,N_7854,N_7303);
and U11462 (N_11462,N_9292,N_7767);
nand U11463 (N_11463,N_9728,N_9287);
nand U11464 (N_11464,N_7702,N_7631);
or U11465 (N_11465,N_9536,N_7880);
and U11466 (N_11466,N_6240,N_8759);
nand U11467 (N_11467,N_9289,N_9823);
nor U11468 (N_11468,N_7071,N_7494);
nand U11469 (N_11469,N_9566,N_5755);
xor U11470 (N_11470,N_9087,N_6841);
and U11471 (N_11471,N_5469,N_9216);
nor U11472 (N_11472,N_5313,N_6652);
xnor U11473 (N_11473,N_7301,N_8161);
nand U11474 (N_11474,N_5485,N_5209);
nor U11475 (N_11475,N_7201,N_6967);
nor U11476 (N_11476,N_9487,N_5540);
nand U11477 (N_11477,N_8562,N_9203);
nand U11478 (N_11478,N_8489,N_5499);
or U11479 (N_11479,N_7211,N_5006);
xnor U11480 (N_11480,N_6660,N_6423);
xnor U11481 (N_11481,N_5436,N_5587);
nor U11482 (N_11482,N_8581,N_9051);
nor U11483 (N_11483,N_7076,N_9339);
xor U11484 (N_11484,N_6265,N_7650);
and U11485 (N_11485,N_9387,N_6757);
or U11486 (N_11486,N_7440,N_6688);
and U11487 (N_11487,N_7226,N_8927);
nor U11488 (N_11488,N_9832,N_8078);
and U11489 (N_11489,N_8288,N_8116);
and U11490 (N_11490,N_6128,N_5077);
nor U11491 (N_11491,N_8202,N_9127);
nor U11492 (N_11492,N_7224,N_6497);
or U11493 (N_11493,N_7277,N_7051);
xnor U11494 (N_11494,N_9577,N_5810);
xnor U11495 (N_11495,N_6093,N_6051);
and U11496 (N_11496,N_6867,N_5659);
or U11497 (N_11497,N_9213,N_6636);
nand U11498 (N_11498,N_5635,N_8435);
xnor U11499 (N_11499,N_6627,N_7692);
nand U11500 (N_11500,N_7671,N_9175);
and U11501 (N_11501,N_7838,N_9954);
nand U11502 (N_11502,N_6902,N_5442);
xor U11503 (N_11503,N_5301,N_5492);
nor U11504 (N_11504,N_9085,N_5179);
nor U11505 (N_11505,N_8323,N_7403);
nand U11506 (N_11506,N_7030,N_5225);
or U11507 (N_11507,N_7334,N_5037);
xor U11508 (N_11508,N_7484,N_6558);
or U11509 (N_11509,N_8700,N_8326);
nand U11510 (N_11510,N_5212,N_5765);
nand U11511 (N_11511,N_6782,N_8152);
and U11512 (N_11512,N_8130,N_8339);
and U11513 (N_11513,N_6003,N_6792);
xor U11514 (N_11514,N_8902,N_7437);
nand U11515 (N_11515,N_5429,N_7595);
nand U11516 (N_11516,N_9530,N_5407);
nand U11517 (N_11517,N_6575,N_7287);
nand U11518 (N_11518,N_7685,N_5170);
nor U11519 (N_11519,N_7235,N_8641);
nand U11520 (N_11520,N_6973,N_5486);
nand U11521 (N_11521,N_9770,N_5343);
and U11522 (N_11522,N_6048,N_7386);
and U11523 (N_11523,N_6120,N_7117);
or U11524 (N_11524,N_6087,N_5541);
or U11525 (N_11525,N_7470,N_8068);
xor U11526 (N_11526,N_9723,N_9806);
or U11527 (N_11527,N_7715,N_9791);
or U11528 (N_11528,N_5972,N_7271);
xnor U11529 (N_11529,N_5718,N_8857);
nor U11530 (N_11530,N_9783,N_7501);
nor U11531 (N_11531,N_8693,N_5619);
or U11532 (N_11532,N_9958,N_7963);
and U11533 (N_11533,N_5314,N_5645);
and U11534 (N_11534,N_8519,N_8664);
xnor U11535 (N_11535,N_9489,N_5727);
xnor U11536 (N_11536,N_6739,N_7155);
or U11537 (N_11537,N_8285,N_8621);
or U11538 (N_11538,N_8403,N_6791);
and U11539 (N_11539,N_6727,N_6203);
nand U11540 (N_11540,N_6658,N_6421);
nor U11541 (N_11541,N_6580,N_8033);
and U11542 (N_11542,N_7441,N_7368);
nor U11543 (N_11543,N_6701,N_5361);
nand U11544 (N_11544,N_7171,N_6794);
nand U11545 (N_11545,N_7175,N_5507);
xor U11546 (N_11546,N_6258,N_8115);
nor U11547 (N_11547,N_8740,N_9078);
nand U11548 (N_11548,N_8632,N_5536);
and U11549 (N_11549,N_5388,N_9533);
xor U11550 (N_11550,N_7317,N_7824);
xnor U11551 (N_11551,N_6832,N_5263);
xnor U11552 (N_11552,N_5772,N_8266);
or U11553 (N_11553,N_5753,N_8565);
nand U11554 (N_11554,N_6041,N_8399);
nand U11555 (N_11555,N_7823,N_7414);
nand U11556 (N_11556,N_9576,N_9093);
nand U11557 (N_11557,N_8376,N_8231);
nor U11558 (N_11558,N_8176,N_8714);
nand U11559 (N_11559,N_8462,N_7068);
and U11560 (N_11560,N_9359,N_8963);
xor U11561 (N_11561,N_8332,N_7072);
nor U11562 (N_11562,N_9734,N_9695);
and U11563 (N_11563,N_9166,N_8164);
nand U11564 (N_11564,N_6879,N_6161);
nand U11565 (N_11565,N_6989,N_8838);
nor U11566 (N_11566,N_9810,N_8768);
or U11567 (N_11567,N_6712,N_6426);
and U11568 (N_11568,N_9401,N_8319);
xor U11569 (N_11569,N_6247,N_5035);
nand U11570 (N_11570,N_7450,N_6114);
or U11571 (N_11571,N_7947,N_5775);
and U11572 (N_11572,N_7473,N_9240);
nor U11573 (N_11573,N_9537,N_6218);
xnor U11574 (N_11574,N_9086,N_8644);
nor U11575 (N_11575,N_5126,N_6924);
and U11576 (N_11576,N_9404,N_6527);
and U11577 (N_11577,N_7719,N_9493);
nand U11578 (N_11578,N_6143,N_5310);
and U11579 (N_11579,N_6338,N_9998);
or U11580 (N_11580,N_6100,N_5948);
and U11581 (N_11581,N_9907,N_9908);
and U11582 (N_11582,N_9633,N_6618);
nand U11583 (N_11583,N_8133,N_8046);
nand U11584 (N_11584,N_8913,N_6542);
nand U11585 (N_11585,N_9145,N_6872);
nand U11586 (N_11586,N_6529,N_9082);
and U11587 (N_11587,N_6075,N_9154);
or U11588 (N_11588,N_5688,N_8301);
nand U11589 (N_11589,N_6849,N_6066);
nor U11590 (N_11590,N_8987,N_8094);
nor U11591 (N_11591,N_7697,N_6656);
and U11592 (N_11592,N_6694,N_5071);
nand U11593 (N_11593,N_9618,N_5360);
and U11594 (N_11594,N_9179,N_5514);
xnor U11595 (N_11595,N_5734,N_8069);
and U11596 (N_11596,N_8996,N_9701);
and U11597 (N_11597,N_8402,N_9999);
nor U11598 (N_11598,N_8814,N_9313);
and U11599 (N_11599,N_7599,N_9601);
nor U11600 (N_11600,N_5567,N_7956);
nor U11601 (N_11601,N_9923,N_9364);
or U11602 (N_11602,N_6770,N_8488);
xor U11603 (N_11603,N_8444,N_6588);
or U11604 (N_11604,N_9255,N_9721);
and U11605 (N_11605,N_7943,N_7530);
nand U11606 (N_11606,N_8674,N_9811);
nand U11607 (N_11607,N_6574,N_5879);
and U11608 (N_11608,N_5111,N_9686);
nor U11609 (N_11609,N_7422,N_5237);
xnor U11610 (N_11610,N_8087,N_6961);
nand U11611 (N_11611,N_5819,N_9445);
nand U11612 (N_11612,N_9321,N_6687);
xor U11613 (N_11613,N_8883,N_6960);
xor U11614 (N_11614,N_7204,N_6199);
and U11615 (N_11615,N_9732,N_8059);
xnor U11616 (N_11616,N_7034,N_5422);
and U11617 (N_11617,N_5968,N_5158);
xor U11618 (N_11618,N_9110,N_8145);
nand U11619 (N_11619,N_6249,N_5450);
nor U11620 (N_11620,N_9277,N_7120);
or U11621 (N_11621,N_7323,N_8341);
or U11622 (N_11622,N_5641,N_7431);
xnor U11623 (N_11623,N_9320,N_5145);
or U11624 (N_11624,N_6693,N_8171);
or U11625 (N_11625,N_9930,N_7312);
or U11626 (N_11626,N_5669,N_7723);
xnor U11627 (N_11627,N_8391,N_5545);
xor U11628 (N_11628,N_6828,N_5140);
nor U11629 (N_11629,N_6935,N_5055);
nor U11630 (N_11630,N_6916,N_9890);
nand U11631 (N_11631,N_5986,N_8995);
nand U11632 (N_11632,N_9882,N_8275);
nor U11633 (N_11633,N_6355,N_8327);
nand U11634 (N_11634,N_9028,N_9057);
or U11635 (N_11635,N_8629,N_7044);
xor U11636 (N_11636,N_6566,N_9949);
nor U11637 (N_11637,N_8920,N_8454);
nand U11638 (N_11638,N_9784,N_5147);
or U11639 (N_11639,N_7081,N_5141);
or U11640 (N_11640,N_6350,N_9983);
xor U11641 (N_11641,N_8729,N_9105);
xor U11642 (N_11642,N_5733,N_6876);
xor U11643 (N_11643,N_5438,N_8182);
nand U11644 (N_11644,N_5683,N_6823);
or U11645 (N_11645,N_7057,N_9422);
nor U11646 (N_11646,N_7839,N_8170);
xor U11647 (N_11647,N_9582,N_6709);
and U11648 (N_11648,N_6548,N_9515);
xor U11649 (N_11649,N_9470,N_7521);
or U11650 (N_11650,N_6632,N_9604);
or U11651 (N_11651,N_7648,N_9817);
xor U11652 (N_11652,N_6852,N_5117);
nand U11653 (N_11653,N_9973,N_5003);
xor U11654 (N_11654,N_7984,N_8175);
nor U11655 (N_11655,N_9318,N_8907);
nand U11656 (N_11656,N_6933,N_6391);
nor U11657 (N_11657,N_9622,N_6082);
xnor U11658 (N_11658,N_5844,N_7456);
and U11659 (N_11659,N_6549,N_6510);
and U11660 (N_11660,N_6420,N_5664);
nor U11661 (N_11661,N_5709,N_5241);
nor U11662 (N_11662,N_8761,N_9607);
and U11663 (N_11663,N_7084,N_7698);
nand U11664 (N_11664,N_9774,N_9245);
nand U11665 (N_11665,N_6827,N_9206);
nor U11666 (N_11666,N_5878,N_5556);
nor U11667 (N_11667,N_5758,N_7768);
nand U11668 (N_11668,N_7275,N_5888);
xor U11669 (N_11669,N_8593,N_9330);
and U11670 (N_11670,N_9163,N_8112);
or U11671 (N_11671,N_8943,N_6256);
nand U11672 (N_11672,N_5118,N_9637);
nor U11673 (N_11673,N_8321,N_5850);
xor U11674 (N_11674,N_5525,N_9395);
or U11675 (N_11675,N_6653,N_8442);
nor U11676 (N_11676,N_9225,N_6243);
or U11677 (N_11677,N_5328,N_7091);
or U11678 (N_11678,N_6328,N_7008);
nor U11679 (N_11679,N_6040,N_7741);
and U11680 (N_11680,N_6320,N_7083);
or U11681 (N_11681,N_5547,N_7735);
and U11682 (N_11682,N_7813,N_7803);
xor U11683 (N_11683,N_5088,N_5306);
and U11684 (N_11684,N_9219,N_9978);
and U11685 (N_11685,N_8764,N_8238);
xor U11686 (N_11686,N_5198,N_9668);
or U11687 (N_11687,N_9553,N_7157);
or U11688 (N_11688,N_9554,N_8262);
nand U11689 (N_11689,N_6537,N_8430);
xnor U11690 (N_11690,N_8233,N_6742);
or U11691 (N_11691,N_7332,N_5877);
nor U11692 (N_11692,N_8375,N_7817);
and U11693 (N_11693,N_6886,N_7237);
xnor U11694 (N_11694,N_7808,N_7019);
nand U11695 (N_11695,N_5539,N_7912);
and U11696 (N_11696,N_9563,N_9918);
and U11697 (N_11697,N_6882,N_6319);
and U11698 (N_11698,N_8252,N_7659);
xnor U11699 (N_11699,N_8993,N_9191);
xnor U11700 (N_11700,N_5349,N_8106);
nor U11701 (N_11701,N_7396,N_5148);
xor U11702 (N_11702,N_9431,N_8620);
or U11703 (N_11703,N_8922,N_6308);
nand U11704 (N_11704,N_5926,N_9337);
or U11705 (N_11705,N_9041,N_8044);
or U11706 (N_11706,N_8421,N_9173);
xnor U11707 (N_11707,N_7686,N_7849);
or U11708 (N_11708,N_6711,N_6482);
nor U11709 (N_11709,N_8578,N_8715);
and U11710 (N_11710,N_6646,N_6381);
and U11711 (N_11711,N_8218,N_9702);
xnor U11712 (N_11712,N_6185,N_9473);
nor U11713 (N_11713,N_9916,N_9542);
nand U11714 (N_11714,N_7166,N_6583);
nand U11715 (N_11715,N_7945,N_5448);
nand U11716 (N_11716,N_9503,N_9714);
or U11717 (N_11717,N_8471,N_9910);
and U11718 (N_11718,N_7188,N_7836);
and U11719 (N_11719,N_8103,N_5413);
or U11720 (N_11720,N_9228,N_6682);
nor U11721 (N_11721,N_8680,N_9739);
nand U11722 (N_11722,N_5411,N_7169);
nand U11723 (N_11723,N_9192,N_5504);
or U11724 (N_11724,N_5001,N_9632);
and U11725 (N_11725,N_7772,N_5943);
or U11726 (N_11726,N_9581,N_6313);
nor U11727 (N_11727,N_6388,N_9142);
and U11728 (N_11728,N_9300,N_9809);
or U11729 (N_11729,N_5150,N_5811);
or U11730 (N_11730,N_5654,N_5318);
nand U11731 (N_11731,N_7194,N_9252);
xnor U11732 (N_11732,N_9824,N_6931);
xor U11733 (N_11733,N_6449,N_7863);
and U11734 (N_11734,N_7046,N_7934);
or U11735 (N_11735,N_8140,N_5213);
xor U11736 (N_11736,N_8766,N_7867);
xnor U11737 (N_11737,N_6303,N_9488);
nor U11738 (N_11738,N_7238,N_9904);
xnor U11739 (N_11739,N_7240,N_9825);
nand U11740 (N_11740,N_8230,N_8258);
and U11741 (N_11741,N_5379,N_9628);
nor U11742 (N_11742,N_8614,N_8322);
nor U11743 (N_11743,N_6076,N_9063);
or U11744 (N_11744,N_6069,N_8634);
xor U11745 (N_11745,N_8716,N_5913);
or U11746 (N_11746,N_8105,N_6629);
nand U11747 (N_11747,N_9144,N_7586);
nand U11748 (N_11748,N_6361,N_8889);
and U11749 (N_11749,N_9283,N_8916);
xor U11750 (N_11750,N_7645,N_9669);
or U11751 (N_11751,N_5946,N_9008);
nor U11752 (N_11752,N_7343,N_5622);
xnor U11753 (N_11753,N_7779,N_7054);
nand U11754 (N_11754,N_5277,N_6784);
nor U11755 (N_11755,N_6297,N_8617);
nor U11756 (N_11756,N_6910,N_8216);
nand U11757 (N_11757,N_7654,N_7617);
nor U11758 (N_11758,N_7821,N_5585);
nor U11759 (N_11759,N_9837,N_5293);
and U11760 (N_11760,N_7962,N_5447);
or U11761 (N_11761,N_5940,N_5257);
and U11762 (N_11762,N_6927,N_9932);
or U11763 (N_11763,N_6324,N_9021);
nor U11764 (N_11764,N_9218,N_8282);
or U11765 (N_11765,N_9148,N_6263);
nand U11766 (N_11766,N_8434,N_5776);
nand U11767 (N_11767,N_6472,N_8208);
xor U11768 (N_11768,N_5503,N_5083);
xnor U11769 (N_11769,N_6642,N_9284);
and U11770 (N_11770,N_5697,N_6122);
xnor U11771 (N_11771,N_6622,N_6883);
xor U11772 (N_11772,N_7400,N_5597);
or U11773 (N_11773,N_8709,N_7827);
nand U11774 (N_11774,N_7264,N_5050);
nand U11775 (N_11775,N_7891,N_9772);
nor U11776 (N_11776,N_8236,N_7390);
or U11777 (N_11777,N_8181,N_8637);
and U11778 (N_11778,N_9608,N_8645);
and U11779 (N_11779,N_7798,N_5259);
xnor U11780 (N_11780,N_5510,N_5068);
or U11781 (N_11781,N_7443,N_7029);
nand U11782 (N_11782,N_9838,N_5749);
xor U11783 (N_11783,N_9711,N_6760);
xor U11784 (N_11784,N_5144,N_9937);
nor U11785 (N_11785,N_8685,N_7147);
and U11786 (N_11786,N_8413,N_6159);
or U11787 (N_11787,N_6725,N_8380);
nor U11788 (N_11788,N_5272,N_5096);
nor U11789 (N_11789,N_5099,N_6197);
nor U11790 (N_11790,N_5892,N_5707);
nand U11791 (N_11791,N_7193,N_6746);
xor U11792 (N_11792,N_6678,N_9371);
nor U11793 (N_11793,N_8135,N_8737);
nor U11794 (N_11794,N_5630,N_5309);
xor U11795 (N_11795,N_6759,N_9029);
nor U11796 (N_11796,N_8196,N_8926);
xnor U11797 (N_11797,N_5937,N_8263);
or U11798 (N_11798,N_5777,N_5565);
or U11799 (N_11799,N_8517,N_9552);
xnor U11800 (N_11800,N_6617,N_9207);
nor U11801 (N_11801,N_8468,N_5030);
nand U11802 (N_11802,N_5317,N_6556);
and U11803 (N_11803,N_8122,N_5588);
or U11804 (N_11804,N_6560,N_9374);
xnor U11805 (N_11805,N_6182,N_6393);
or U11806 (N_11806,N_8412,N_8006);
and U11807 (N_11807,N_5027,N_7892);
and U11808 (N_11808,N_7743,N_7328);
nand U11809 (N_11809,N_9655,N_9317);
nor U11810 (N_11810,N_6206,N_7229);
or U11811 (N_11811,N_7611,N_9800);
nor U11812 (N_11812,N_8625,N_6084);
or U11813 (N_11813,N_9684,N_8162);
nand U11814 (N_11814,N_9736,N_8756);
xnor U11815 (N_11815,N_6369,N_9162);
nor U11816 (N_11816,N_8365,N_7802);
nand U11817 (N_11817,N_6302,N_9295);
nor U11818 (N_11818,N_8424,N_5812);
nor U11819 (N_11819,N_9744,N_5730);
and U11820 (N_11820,N_7292,N_6842);
or U11821 (N_11821,N_5381,N_6012);
nand U11822 (N_11822,N_5815,N_5191);
nor U11823 (N_11823,N_6925,N_7025);
and U11824 (N_11824,N_5467,N_9068);
nand U11825 (N_11825,N_9281,N_9090);
and U11826 (N_11826,N_5711,N_5122);
and U11827 (N_11827,N_7938,N_7467);
nor U11828 (N_11828,N_7415,N_5199);
xnor U11829 (N_11829,N_8553,N_7519);
or U11830 (N_11830,N_6705,N_8499);
and U11831 (N_11831,N_8048,N_7064);
or U11832 (N_11832,N_7531,N_9076);
or U11833 (N_11833,N_7020,N_8663);
nand U11834 (N_11834,N_9831,N_8232);
xor U11835 (N_11835,N_6983,N_6053);
and U11836 (N_11836,N_6966,N_7066);
and U11837 (N_11837,N_7192,N_6390);
xnor U11838 (N_11838,N_8564,N_9906);
or U11839 (N_11839,N_5394,N_6269);
xor U11840 (N_11840,N_7624,N_7401);
or U11841 (N_11841,N_9355,N_9513);
nand U11842 (N_11842,N_9079,N_7151);
xor U11843 (N_11843,N_8307,N_5382);
xnor U11844 (N_11844,N_5680,N_7907);
nand U11845 (N_11845,N_7842,N_5444);
xnor U11846 (N_11846,N_7135,N_7592);
or U11847 (N_11847,N_6330,N_7832);
nand U11848 (N_11848,N_5256,N_5956);
nand U11849 (N_11849,N_5859,N_7834);
nand U11850 (N_11850,N_8290,N_9877);
nor U11851 (N_11851,N_9075,N_8409);
or U11852 (N_11852,N_9925,N_6996);
and U11853 (N_11853,N_6512,N_7590);
and U11854 (N_11854,N_5719,N_9641);
xnor U11855 (N_11855,N_6372,N_8660);
xor U11856 (N_11856,N_6273,N_5168);
nor U11857 (N_11857,N_5826,N_6081);
nand U11858 (N_11858,N_5281,N_9119);
nand U11859 (N_11859,N_5445,N_7177);
xor U11860 (N_11860,N_8053,N_9073);
nand U11861 (N_11861,N_9124,N_8647);
xnor U11862 (N_11862,N_5338,N_5063);
and U11863 (N_11863,N_6691,N_6191);
or U11864 (N_11864,N_9549,N_7949);
nor U11865 (N_11865,N_9699,N_8852);
nand U11866 (N_11866,N_5705,N_9223);
nand U11867 (N_11867,N_9562,N_8836);
or U11868 (N_11868,N_7928,N_7845);
and U11869 (N_11869,N_5250,N_6396);
nor U11870 (N_11870,N_5268,N_9547);
and U11871 (N_11871,N_7255,N_5095);
nor U11872 (N_11872,N_6227,N_7267);
or U11873 (N_11873,N_9202,N_7846);
or U11874 (N_11874,N_7338,N_7139);
nand U11875 (N_11875,N_8390,N_5291);
or U11876 (N_11876,N_5463,N_6593);
xnor U11877 (N_11877,N_7866,N_9220);
and U11878 (N_11878,N_5677,N_5961);
nand U11879 (N_11879,N_9365,N_5828);
and U11880 (N_11880,N_8982,N_6923);
nor U11881 (N_11881,N_6513,N_6715);
nand U11882 (N_11882,N_6279,N_9975);
nor U11883 (N_11883,N_9367,N_9568);
or U11884 (N_11884,N_7005,N_5167);
nor U11885 (N_11885,N_5994,N_9993);
nand U11886 (N_11886,N_6714,N_6409);
xor U11887 (N_11887,N_5031,N_5712);
nor U11888 (N_11888,N_6735,N_9062);
xor U11889 (N_11889,N_9902,N_9349);
nand U11890 (N_11890,N_6803,N_8897);
nor U11891 (N_11891,N_8940,N_8358);
nand U11892 (N_11892,N_6612,N_5207);
nand U11893 (N_11893,N_6019,N_9511);
nand U11894 (N_11894,N_9896,N_7790);
and U11895 (N_11895,N_5624,N_5638);
or U11896 (N_11896,N_9357,N_8315);
and U11897 (N_11897,N_7253,N_7124);
and U11898 (N_11898,N_9485,N_7493);
nor U11899 (N_11899,N_5885,N_6090);
and U11900 (N_11900,N_9879,N_9269);
xnor U11901 (N_11901,N_7359,N_8816);
nand U11902 (N_11902,N_8492,N_9878);
xnor U11903 (N_11903,N_6039,N_7268);
or U11904 (N_11904,N_8354,N_8313);
and U11905 (N_11905,N_9012,N_6318);
and U11906 (N_11906,N_7778,N_5740);
nor U11907 (N_11907,N_7371,N_9969);
or U11908 (N_11908,N_6569,N_5538);
nand U11909 (N_11909,N_8296,N_7887);
xor U11910 (N_11910,N_8767,N_9876);
xor U11911 (N_11911,N_5398,N_5053);
xnor U11912 (N_11912,N_6621,N_9926);
nor U11913 (N_11913,N_6786,N_6219);
and U11914 (N_11914,N_6523,N_9689);
xnor U11915 (N_11915,N_7678,N_5472);
nand U11916 (N_11916,N_5273,N_9762);
and U11917 (N_11917,N_6860,N_6608);
and U11918 (N_11918,N_7937,N_7875);
and U11919 (N_11919,N_7900,N_8507);
nand U11920 (N_11920,N_5714,N_6626);
or U11921 (N_11921,N_5803,N_7911);
xnor U11922 (N_11922,N_9661,N_8534);
and U11923 (N_11923,N_8432,N_6600);
nand U11924 (N_11924,N_8211,N_7770);
xnor U11925 (N_11925,N_7552,N_6405);
nand U11926 (N_11926,N_8751,N_6985);
and U11927 (N_11927,N_6899,N_9571);
nor U11928 (N_11928,N_5818,N_8822);
nand U11929 (N_11929,N_9822,N_8741);
nand U11930 (N_11930,N_5806,N_6663);
nor U11931 (N_11931,N_7840,N_9624);
xnor U11932 (N_11932,N_6173,N_6716);
or U11933 (N_11933,N_9031,N_6943);
and U11934 (N_11934,N_7924,N_9155);
nor U11935 (N_11935,N_7921,N_6395);
or U11936 (N_11936,N_6212,N_7794);
and U11937 (N_11937,N_9064,N_5814);
nand U11938 (N_11938,N_8460,N_8001);
xnor U11939 (N_11939,N_6551,N_8378);
and U11940 (N_11940,N_5032,N_8239);
nor U11941 (N_11941,N_7322,N_8071);
nor U11942 (N_11942,N_9054,N_7460);
nor U11943 (N_11943,N_7584,N_9664);
and U11944 (N_11944,N_6166,N_7699);
or U11945 (N_11945,N_7571,N_5793);
xnor U11946 (N_11946,N_5214,N_5461);
or U11947 (N_11947,N_9241,N_9595);
or U11948 (N_11948,N_8666,N_8153);
nor U11949 (N_11949,N_6438,N_6857);
nand U11950 (N_11950,N_9251,N_9673);
xor U11951 (N_11951,N_7825,N_8265);
or U11952 (N_11952,N_5226,N_6056);
and U11953 (N_11953,N_9013,N_9880);
and U11954 (N_11954,N_8718,N_8191);
xor U11955 (N_11955,N_9656,N_9153);
xor U11956 (N_11956,N_8948,N_8064);
and U11957 (N_11957,N_9746,N_5288);
or U11958 (N_11958,N_7176,N_8866);
or U11959 (N_11959,N_6489,N_5332);
xor U11960 (N_11960,N_8260,N_7215);
or U11961 (N_11961,N_5581,N_5555);
or U11962 (N_11962,N_5665,N_9270);
nor U11963 (N_11963,N_9597,N_6184);
xnor U11964 (N_11964,N_9840,N_9865);
nand U11965 (N_11965,N_7366,N_9157);
xor U11966 (N_11966,N_9638,N_6326);
xor U11967 (N_11967,N_9919,N_8479);
nor U11968 (N_11968,N_7142,N_9764);
xor U11969 (N_11969,N_6366,N_7049);
or U11970 (N_11970,N_7162,N_5871);
xor U11971 (N_11971,N_7913,N_5252);
or U11972 (N_11972,N_7112,N_9074);
and U11973 (N_11973,N_7988,N_8092);
nor U11974 (N_11974,N_7336,N_9933);
and U11975 (N_11975,N_7994,N_7252);
or U11976 (N_11976,N_9400,N_5169);
xor U11977 (N_11977,N_5154,N_5757);
nor U11978 (N_11978,N_7027,N_9168);
or U11979 (N_11979,N_7562,N_6524);
and U11980 (N_11980,N_8909,N_8813);
xor U11981 (N_11981,N_9704,N_5124);
and U11982 (N_11982,N_5621,N_6183);
and U11983 (N_11983,N_7644,N_8830);
nand U11984 (N_11984,N_8667,N_5773);
xor U11985 (N_11985,N_9109,N_5867);
and U11986 (N_11986,N_8959,N_5261);
or U11987 (N_11987,N_7420,N_5785);
xnor U11988 (N_11988,N_8912,N_8906);
nor U11989 (N_11989,N_6250,N_6375);
xnor U11990 (N_11990,N_9856,N_7259);
or U11991 (N_11991,N_5221,N_5376);
xnor U11992 (N_11992,N_6917,N_8794);
nand U11993 (N_11993,N_6370,N_5764);
nor U11994 (N_11994,N_7781,N_5889);
nand U11995 (N_11995,N_9421,N_6597);
or U11996 (N_11996,N_6057,N_8119);
xnor U11997 (N_11997,N_9376,N_8777);
or U11998 (N_11998,N_9749,N_7295);
and U11999 (N_11999,N_9081,N_8942);
xor U12000 (N_12000,N_6590,N_9182);
or U12001 (N_12001,N_7241,N_8222);
nand U12002 (N_12002,N_5506,N_9475);
nand U12003 (N_12003,N_9615,N_5358);
xor U12004 (N_12004,N_6058,N_8603);
or U12005 (N_12005,N_6130,N_5817);
nand U12006 (N_12006,N_5408,N_7716);
nor U12007 (N_12007,N_6969,N_7657);
and U12008 (N_12008,N_5702,N_5188);
nand U12009 (N_12009,N_9038,N_5537);
nand U12010 (N_12010,N_5593,N_8535);
xnor U12011 (N_12011,N_5706,N_7006);
xnor U12012 (N_12012,N_6815,N_9920);
xor U12013 (N_12013,N_6504,N_8542);
xor U12014 (N_12014,N_6721,N_7740);
xor U12015 (N_12015,N_5217,N_6119);
and U12016 (N_12016,N_5164,N_7955);
nand U12017 (N_12017,N_5276,N_8431);
and U12018 (N_12018,N_5005,N_9002);
xor U12019 (N_12019,N_7942,N_6316);
xnor U12020 (N_12020,N_7957,N_5392);
nand U12021 (N_12021,N_8029,N_5109);
nand U12022 (N_12022,N_6821,N_6756);
nor U12023 (N_12023,N_8226,N_8522);
or U12024 (N_12024,N_7032,N_9146);
nor U12025 (N_12025,N_8742,N_8953);
nand U12026 (N_12026,N_8023,N_7082);
nor U12027 (N_12027,N_6585,N_6616);
or U12028 (N_12028,N_9570,N_7357);
or U12029 (N_12029,N_7857,N_6109);
or U12030 (N_12030,N_8229,N_8473);
xor U12031 (N_12031,N_6835,N_5575);
nor U12032 (N_12032,N_8372,N_7464);
or U12033 (N_12033,N_5675,N_6337);
or U12034 (N_12034,N_6862,N_8362);
and U12035 (N_12035,N_8582,N_6605);
nor U12036 (N_12036,N_8529,N_5437);
and U12037 (N_12037,N_5684,N_8055);
and U12038 (N_12038,N_6424,N_6495);
nand U12039 (N_12039,N_7968,N_6137);
nor U12040 (N_12040,N_7333,N_9439);
nor U12041 (N_12041,N_6357,N_8136);
and U12042 (N_12042,N_6222,N_8929);
nor U12043 (N_12043,N_5136,N_8283);
and U12044 (N_12044,N_7696,N_5590);
nand U12045 (N_12045,N_9516,N_9440);
nor U12046 (N_12046,N_7709,N_6651);
nor U12047 (N_12047,N_8586,N_5672);
nor U12048 (N_12048,N_6004,N_8521);
and U12049 (N_12049,N_6228,N_7684);
nand U12050 (N_12050,N_7406,N_7948);
xor U12051 (N_12051,N_6520,N_5204);
xnor U12052 (N_12052,N_8117,N_6155);
xnor U12053 (N_12053,N_7766,N_5736);
xnor U12054 (N_12054,N_5795,N_7600);
nor U12055 (N_12055,N_6408,N_8189);
xnor U12056 (N_12056,N_8185,N_8352);
nand U12057 (N_12057,N_7722,N_6992);
or U12058 (N_12058,N_6624,N_5230);
xor U12059 (N_12059,N_9338,N_8653);
xnor U12060 (N_12060,N_6980,N_6797);
nor U12061 (N_12061,N_5434,N_8919);
and U12062 (N_12062,N_5865,N_5330);
nor U12063 (N_12063,N_9914,N_8173);
nand U12064 (N_12064,N_7558,N_7170);
or U12065 (N_12065,N_7452,N_5858);
xnor U12066 (N_12066,N_6187,N_7001);
and U12067 (N_12067,N_9426,N_5742);
xnor U12068 (N_12068,N_7085,N_6005);
and U12069 (N_12069,N_7615,N_5627);
and U12070 (N_12070,N_6229,N_7186);
or U12071 (N_12071,N_6719,N_6476);
and U12072 (N_12072,N_7128,N_8169);
or U12073 (N_12073,N_5161,N_8703);
xnor U12074 (N_12074,N_5181,N_5292);
xor U12075 (N_12075,N_7377,N_7926);
nand U12076 (N_12076,N_5929,N_9406);
xor U12077 (N_12077,N_8449,N_6237);
nor U12078 (N_12078,N_7561,N_5409);
xnor U12079 (N_12079,N_7983,N_7872);
nand U12080 (N_12080,N_5114,N_7492);
xnor U12081 (N_12081,N_7754,N_8142);
nand U12082 (N_12082,N_9111,N_8864);
nand U12083 (N_12083,N_6930,N_6113);
nor U12084 (N_12084,N_8496,N_7920);
nor U12085 (N_12085,N_9847,N_9293);
xnor U12086 (N_12086,N_7718,N_8877);
nor U12087 (N_12087,N_9279,N_9596);
nand U12088 (N_12088,N_5133,N_5936);
nand U12089 (N_12089,N_7389,N_5921);
nand U12090 (N_12090,N_5033,N_5614);
xor U12091 (N_12091,N_9534,N_7350);
or U12092 (N_12092,N_5304,N_5060);
nand U12093 (N_12093,N_5872,N_6295);
or U12094 (N_12094,N_8842,N_6089);
nor U12095 (N_12095,N_6398,N_5640);
nand U12096 (N_12096,N_5896,N_7411);
xor U12097 (N_12097,N_5402,N_6466);
and U12098 (N_12098,N_8480,N_9286);
and U12099 (N_12099,N_5034,N_7508);
nor U12100 (N_12100,N_8547,N_5162);
xnor U12101 (N_12101,N_8190,N_8580);
xor U12102 (N_12102,N_9351,N_8825);
and U12103 (N_12103,N_6259,N_6257);
and U12104 (N_12104,N_5843,N_9342);
nand U12105 (N_12105,N_7469,N_8018);
nand U12106 (N_12106,N_8727,N_7290);
nor U12107 (N_12107,N_7052,N_8510);
nor U12108 (N_12108,N_8184,N_7736);
nand U12109 (N_12109,N_9429,N_8946);
nor U12110 (N_12110,N_8795,N_7058);
and U12111 (N_12111,N_5203,N_8981);
nor U12112 (N_12112,N_6707,N_6516);
nand U12113 (N_12113,N_8682,N_9703);
or U12114 (N_12114,N_5498,N_6620);
nand U12115 (N_12115,N_9199,N_7739);
nand U12116 (N_12116,N_5636,N_5999);
and U12117 (N_12117,N_8930,N_5846);
or U12118 (N_12118,N_5512,N_9249);
xor U12119 (N_12119,N_5646,N_8114);
nand U12120 (N_12120,N_6202,N_9676);
nand U12121 (N_12121,N_8686,N_6640);
or U12122 (N_12122,N_6704,N_5490);
nor U12123 (N_12123,N_8528,N_8187);
nor U12124 (N_12124,N_8379,N_6347);
and U12125 (N_12125,N_8994,N_9435);
or U12126 (N_12126,N_7626,N_9016);
and U12127 (N_12127,N_5781,N_6589);
or U12128 (N_12128,N_8792,N_9591);
or U12129 (N_12129,N_9898,N_6816);
and U12130 (N_12130,N_5455,N_7806);
and U12131 (N_12131,N_5957,N_7608);
xnor U12132 (N_12132,N_7004,N_9327);
nand U12133 (N_12133,N_8918,N_6681);
xor U12134 (N_12134,N_5116,N_8587);
xnor U12135 (N_12135,N_5305,N_6487);
and U12136 (N_12136,N_9496,N_6515);
nor U12137 (N_12137,N_6947,N_9875);
nor U12138 (N_12138,N_9495,N_6460);
xor U12139 (N_12139,N_8775,N_7674);
nor U12140 (N_12140,N_8118,N_5821);
nand U12141 (N_12141,N_6304,N_9350);
xnor U12142 (N_12142,N_6292,N_9971);
nand U12143 (N_12143,N_6215,N_7397);
xor U12144 (N_12144,N_8353,N_5788);
or U12145 (N_12145,N_7227,N_5244);
nand U12146 (N_12146,N_6178,N_6208);
or U12147 (N_12147,N_9517,N_8408);
and U12148 (N_12148,N_5897,N_7967);
xnor U12149 (N_12149,N_7643,N_9519);
nand U12150 (N_12150,N_6942,N_8726);
nand U12151 (N_12151,N_5609,N_7315);
xnor U12152 (N_12152,N_7819,N_9454);
nor U12153 (N_12153,N_5743,N_8544);
and U12154 (N_12154,N_8463,N_5405);
nand U12155 (N_12155,N_8911,N_9072);
nand U12156 (N_12156,N_7961,N_8848);
nor U12157 (N_12157,N_9884,N_7543);
or U12158 (N_12158,N_9834,N_8923);
or U12159 (N_12159,N_5963,N_7257);
and U12160 (N_12160,N_9551,N_7425);
and U12161 (N_12161,N_6885,N_9333);
nor U12162 (N_12162,N_8104,N_5366);
nor U12163 (N_12163,N_7417,N_7137);
nor U12164 (N_12164,N_9140,N_9790);
nand U12165 (N_12165,N_9670,N_6722);
xor U12166 (N_12166,N_9120,N_7282);
or U12167 (N_12167,N_8337,N_5840);
nor U12168 (N_12168,N_6165,N_9165);
and U12169 (N_12169,N_6126,N_8017);
xnor U12170 (N_12170,N_8570,N_7075);
nor U12171 (N_12171,N_6887,N_5410);
and U12172 (N_12172,N_5960,N_8120);
or U12173 (N_12173,N_8450,N_7138);
xor U12174 (N_12174,N_8312,N_9491);
nor U12175 (N_12175,N_5193,N_5121);
and U12176 (N_12176,N_5180,N_6244);
and U12177 (N_12177,N_6376,N_5454);
or U12178 (N_12178,N_6956,N_8343);
xor U12179 (N_12179,N_6579,N_5216);
nor U12180 (N_12180,N_9196,N_8381);
and U12181 (N_12181,N_7864,N_5065);
nor U12182 (N_12182,N_7239,N_7979);
xnor U12183 (N_12183,N_9126,N_6246);
and U12184 (N_12184,N_9373,N_9309);
xnor U12185 (N_12185,N_7974,N_8605);
or U12186 (N_12186,N_8289,N_6604);
xnor U12187 (N_12187,N_9523,N_9586);
or U12188 (N_12188,N_9629,N_8411);
and U12189 (N_12189,N_7413,N_8652);
or U12190 (N_12190,N_9492,N_7062);
nand U12191 (N_12191,N_7605,N_8699);
xor U12192 (N_12192,N_9657,N_9995);
xor U12193 (N_12193,N_7297,N_6968);
or U12194 (N_12194,N_6957,N_5739);
xnor U12195 (N_12195,N_5981,N_6734);
xor U12196 (N_12196,N_5375,N_9160);
and U12197 (N_12197,N_8744,N_7305);
and U12198 (N_12198,N_8493,N_9500);
nand U12199 (N_12199,N_8220,N_7299);
and U12200 (N_12200,N_6737,N_5801);
xnor U12201 (N_12201,N_6939,N_9680);
or U12202 (N_12202,N_6180,N_6951);
or U12203 (N_12203,N_9802,N_8509);
or U12204 (N_12204,N_8788,N_8882);
nand U12205 (N_12205,N_8887,N_5880);
or U12206 (N_12206,N_7581,N_9868);
and U12207 (N_12207,N_6628,N_6260);
xor U12208 (N_12208,N_5183,N_9472);
nor U12209 (N_12209,N_9619,N_7320);
nor U12210 (N_12210,N_6798,N_5623);
or U12211 (N_12211,N_5589,N_5400);
nor U12212 (N_12212,N_6031,N_6937);
xnor U12213 (N_12213,N_9560,N_9336);
xnor U12214 (N_12214,N_9845,N_7784);
and U12215 (N_12215,N_6170,N_9185);
or U12216 (N_12216,N_6536,N_5822);
nand U12217 (N_12217,N_8248,N_9268);
xnor U12218 (N_12218,N_8389,N_5255);
and U12219 (N_12219,N_8827,N_5952);
xor U12220 (N_12220,N_8261,N_7901);
xor U12221 (N_12221,N_9050,N_5602);
or U12222 (N_12222,N_8880,N_5768);
nor U12223 (N_12223,N_8573,N_7500);
or U12224 (N_12224,N_6729,N_5222);
xor U12225 (N_12225,N_9660,N_9015);
nand U12226 (N_12226,N_5914,N_7537);
and U12227 (N_12227,N_6775,N_9048);
and U12228 (N_12228,N_5348,N_5196);
nand U12229 (N_12229,N_7510,N_6157);
xnor U12230 (N_12230,N_5266,N_9077);
nand U12231 (N_12231,N_5386,N_5044);
nor U12232 (N_12232,N_9957,N_8797);
and U12233 (N_12233,N_6776,N_7324);
or U12234 (N_12234,N_7757,N_9512);
or U12235 (N_12235,N_9694,N_8949);
or U12236 (N_12236,N_8643,N_5969);
nand U12237 (N_12237,N_8917,N_7444);
nand U12238 (N_12238,N_7038,N_5813);
nand U12239 (N_12239,N_5562,N_9097);
and U12240 (N_12240,N_5553,N_7541);
xor U12241 (N_12241,N_7250,N_9767);
and U12242 (N_12242,N_9671,N_8724);
and U12243 (N_12243,N_6117,N_6340);
nand U12244 (N_12244,N_5335,N_5326);
xor U12245 (N_12245,N_6358,N_8530);
or U12246 (N_12246,N_7829,N_7208);
xor U12247 (N_12247,N_6188,N_7944);
nor U12248 (N_12248,N_6427,N_5729);
and U12249 (N_12249,N_8418,N_8651);
or U12250 (N_12250,N_6104,N_5592);
nand U12251 (N_12251,N_8213,N_8031);
xor U12252 (N_12252,N_5119,N_7958);
or U12253 (N_12253,N_6006,N_5744);
and U12254 (N_12254,N_8955,N_9305);
nand U12255 (N_12255,N_8810,N_9982);
nor U12256 (N_12256,N_9147,N_5339);
and U12257 (N_12257,N_6023,N_9950);
nor U12258 (N_12258,N_7383,N_9388);
nand U12259 (N_12259,N_5833,N_5949);
nand U12260 (N_12260,N_9246,N_8807);
or U12261 (N_12261,N_8840,N_8010);
nor U12262 (N_12262,N_8420,N_5905);
nor U12263 (N_12263,N_5152,N_6230);
and U12264 (N_12264,N_9593,N_5847);
xnor U12265 (N_12265,N_5577,N_9123);
nor U12266 (N_12266,N_8128,N_8102);
nand U12267 (N_12267,N_7041,N_8831);
xnor U12268 (N_12268,N_8374,N_9719);
xor U12269 (N_12269,N_8335,N_9964);
nand U12270 (N_12270,N_7256,N_9089);
or U12271 (N_12271,N_7013,N_5515);
and U12272 (N_12272,N_6036,N_5875);
and U12273 (N_12273,N_9208,N_5004);
nand U12274 (N_12274,N_5127,N_6606);
or U12275 (N_12275,N_6447,N_7662);
nor U12276 (N_12276,N_9578,N_8702);
xnor U12277 (N_12277,N_8550,N_8508);
nand U12278 (N_12278,N_8846,N_6799);
or U12279 (N_12279,N_6613,N_8240);
nor U12280 (N_12280,N_8474,N_8461);
nor U12281 (N_12281,N_9527,N_5270);
nand U12282 (N_12282,N_9323,N_9805);
or U12283 (N_12283,N_9870,N_7499);
xor U12284 (N_12284,N_7203,N_5548);
or U12285 (N_12285,N_5954,N_9234);
xnor U12286 (N_12286,N_7289,N_9979);
xor U12287 (N_12287,N_7964,N_9813);
xnor U12288 (N_12288,N_8752,N_5886);
or U12289 (N_12289,N_9579,N_5804);
nor U12290 (N_12290,N_6022,N_5939);
nor U12291 (N_12291,N_7016,N_6498);
nand U12292 (N_12292,N_6539,N_8146);
xnor U12293 (N_12293,N_5975,N_6311);
nor U12294 (N_12294,N_6262,N_9752);
or U12295 (N_12295,N_6301,N_8787);
and U12296 (N_12296,N_8304,N_6298);
xor U12297 (N_12297,N_5265,N_6634);
nor U12298 (N_12298,N_9688,N_5762);
xnor U12299 (N_12299,N_6755,N_5435);
or U12300 (N_12300,N_6150,N_6034);
nor U12301 (N_12301,N_9693,N_8014);
and U12302 (N_12302,N_6751,N_8892);
and U12303 (N_12303,N_6192,N_7079);
nor U12304 (N_12304,N_6929,N_8203);
and U12305 (N_12305,N_8695,N_5479);
or U12306 (N_12306,N_7429,N_7603);
and U12307 (N_12307,N_8370,N_9953);
xnor U12308 (N_12308,N_9267,N_9885);
and U12309 (N_12309,N_8583,N_5605);
or U12310 (N_12310,N_8000,N_5876);
nand U12311 (N_12311,N_9116,N_8256);
or U12312 (N_12312,N_6779,N_7489);
xnor U12313 (N_12313,N_9594,N_7632);
nor U12314 (N_12314,N_7329,N_7011);
nand U12315 (N_12315,N_5988,N_8606);
xor U12316 (N_12316,N_5347,N_8111);
and U12317 (N_12317,N_6881,N_9545);
and U12318 (N_12318,N_7553,N_8052);
nor U12319 (N_12319,N_7104,N_9232);
nand U12320 (N_12320,N_7298,N_6054);
nand U12321 (N_12321,N_8514,N_5628);
and U12322 (N_12322,N_5789,N_7405);
nor U12323 (N_12323,N_7364,N_9114);
xor U12324 (N_12324,N_9574,N_7167);
nor U12325 (N_12325,N_7504,N_5025);
or U12326 (N_12326,N_9104,N_8697);
and U12327 (N_12327,N_8636,N_5112);
or U12328 (N_12328,N_9183,N_9242);
nor U12329 (N_12329,N_8849,N_5098);
xor U12330 (N_12330,N_6290,N_6099);
or U12331 (N_12331,N_8318,N_8038);
xor U12332 (N_12332,N_9459,N_5089);
or U12333 (N_12333,N_7512,N_9829);
nand U12334 (N_12334,N_6317,N_8366);
nor U12335 (N_12335,N_6610,N_8299);
or U12336 (N_12336,N_6665,N_8861);
and U12337 (N_12337,N_8224,N_6115);
or U12338 (N_12338,N_5965,N_6952);
xor U12339 (N_12339,N_6145,N_6047);
and U12340 (N_12340,N_5710,N_7090);
or U12341 (N_12341,N_8633,N_5699);
nor U12342 (N_12342,N_6248,N_6535);
nand U12343 (N_12343,N_8426,N_9730);
and U12344 (N_12344,N_5195,N_7818);
and U12345 (N_12345,N_7490,N_6477);
or U12346 (N_12346,N_5962,N_9425);
nand U12347 (N_12347,N_7036,N_8668);
nand U12348 (N_12348,N_8179,N_5076);
or U12349 (N_12349,N_7761,N_9646);
and U12350 (N_12350,N_7340,N_6471);
or U12351 (N_12351,N_6033,N_7022);
or U12352 (N_12352,N_8546,N_6909);
and U12353 (N_12353,N_8785,N_5551);
or U12354 (N_12354,N_7272,N_8572);
nor U12355 (N_12355,N_5018,N_5308);
nand U12356 (N_12356,N_7565,N_7978);
xnor U12357 (N_12357,N_6334,N_7225);
nor U12358 (N_12358,N_9261,N_5953);
nor U12359 (N_12359,N_8859,N_7412);
or U12360 (N_12360,N_9288,N_6869);
nand U12361 (N_12361,N_6572,N_5713);
or U12362 (N_12362,N_7384,N_7304);
nor U12363 (N_12363,N_6214,N_7228);
xnor U12364 (N_12364,N_5171,N_5470);
and U12365 (N_12365,N_6091,N_9662);
and U12366 (N_12366,N_6200,N_8021);
xor U12367 (N_12367,N_8821,N_6833);
nand U12368 (N_12368,N_5039,N_5559);
nor U12369 (N_12369,N_8900,N_6895);
nand U12370 (N_12370,N_6404,N_9987);
and U12371 (N_12371,N_5439,N_8359);
xnor U12372 (N_12372,N_8330,N_8746);
nor U12373 (N_12373,N_7939,N_5660);
and U12374 (N_12374,N_6568,N_9962);
nor U12375 (N_12375,N_8329,N_7990);
or U12376 (N_12376,N_7726,N_9354);
nand U12377 (N_12377,N_6554,N_5253);
xnor U12378 (N_12378,N_7693,N_5722);
xor U12379 (N_12379,N_8451,N_7424);
and U12380 (N_12380,N_8423,N_8965);
nor U12381 (N_12381,N_8250,N_5501);
or U12382 (N_12382,N_7791,N_6928);
nor U12383 (N_12383,N_6264,N_8567);
nand U12384 (N_12384,N_7387,N_6795);
xnor U12385 (N_12385,N_8286,N_8600);
and U12386 (N_12386,N_8158,N_5494);
or U12387 (N_12387,N_7941,N_7756);
nor U12388 (N_12388,N_8506,N_6685);
nor U12389 (N_12389,N_9176,N_5676);
nand U12390 (N_12390,N_6459,N_6410);
or U12391 (N_12391,N_6571,N_6027);
xor U12392 (N_12392,N_8915,N_5524);
nor U12393 (N_12393,N_6431,N_7185);
and U12394 (N_12394,N_8273,N_9538);
nand U12395 (N_12395,N_8217,N_9827);
or U12396 (N_12396,N_5834,N_5038);
xor U12397 (N_12397,N_9635,N_7207);
nand U12398 (N_12398,N_7868,N_6940);
nand U12399 (N_12399,N_6668,N_5247);
nand U12400 (N_12400,N_8401,N_6373);
or U12401 (N_12401,N_6445,N_9308);
nor U12402 (N_12402,N_6344,N_6698);
nand U12403 (N_12403,N_9094,N_8371);
nand U12404 (N_12404,N_9457,N_8779);
or U12405 (N_12405,N_7896,N_6414);
nand U12406 (N_12406,N_9994,N_7056);
nor U12407 (N_12407,N_8481,N_8368);
xnor U12408 (N_12408,N_8723,N_8436);
nand U12409 (N_12409,N_8025,N_7883);
nand U12410 (N_12410,N_9335,N_7533);
and U12411 (N_12411,N_9986,N_5215);
xor U12412 (N_12412,N_5368,N_6306);
xnor U12413 (N_12413,N_7604,N_5113);
nand U12414 (N_12414,N_5481,N_9792);
xnor U12415 (N_12415,N_9262,N_5990);
and U12416 (N_12416,N_9316,N_7073);
xor U12417 (N_12417,N_7214,N_8291);
xor U12418 (N_12418,N_5748,N_6045);
nor U12419 (N_12419,N_8800,N_8952);
nor U12420 (N_12420,N_7347,N_9448);
xnor U12421 (N_12421,N_7126,N_8338);
or U12422 (N_12422,N_5146,N_9871);
nor U12423 (N_12423,N_5647,N_7474);
nor U12424 (N_12424,N_7885,N_7642);
or U12425 (N_12425,N_9678,N_9780);
and U12426 (N_12426,N_9892,N_9189);
nor U12427 (N_12427,N_9451,N_7133);
nand U12428 (N_12428,N_9360,N_7977);
and U12429 (N_12429,N_5891,N_6239);
xnor U12430 (N_12430,N_7555,N_5615);
nand U12431 (N_12431,N_7837,N_7345);
nor U12432 (N_12432,N_9458,N_9891);
nor U12433 (N_12433,N_9955,N_7114);
and U12434 (N_12434,N_6070,N_9712);
nor U12435 (N_12435,N_5320,N_6643);
and U12436 (N_12436,N_5417,N_9465);
xor U12437 (N_12437,N_6348,N_9152);
or U12438 (N_12438,N_6281,N_6573);
xnor U12439 (N_12439,N_5983,N_6436);
nand U12440 (N_12440,N_7109,N_7302);
or U12441 (N_12441,N_7223,N_8205);
nor U12442 (N_12442,N_8722,N_6736);
nand U12443 (N_12443,N_9857,N_5989);
or U12444 (N_12444,N_6458,N_9529);
nor U12445 (N_12445,N_6220,N_5851);
or U12446 (N_12446,N_8284,N_9897);
nand U12447 (N_12447,N_5717,N_6892);
xor U12448 (N_12448,N_8675,N_5258);
nand U12449 (N_12449,N_5495,N_6949);
or U12450 (N_12450,N_5650,N_7220);
nor U12451 (N_12451,N_9205,N_8469);
xnor U12452 (N_12452,N_9402,N_5007);
or U12453 (N_12453,N_7393,N_7925);
xor U12454 (N_12454,N_8034,N_9972);
xor U12455 (N_12455,N_7720,N_9204);
xor U12456 (N_12456,N_6587,N_9375);
and U12457 (N_12457,N_5064,N_7830);
nand U12458 (N_12458,N_5580,N_9230);
nand U12459 (N_12459,N_9210,N_8910);
nand U12460 (N_12460,N_6289,N_6907);
or U12461 (N_12461,N_7471,N_8168);
or U12462 (N_12462,N_6224,N_6764);
or U12463 (N_12463,N_9229,N_5393);
and U12464 (N_12464,N_7923,N_6488);
nand U12465 (N_12465,N_7319,N_8609);
or U12466 (N_12466,N_5177,N_5973);
and U12467 (N_12467,N_8295,N_7435);
nand U12468 (N_12468,N_6692,N_9259);
or U12469 (N_12469,N_5131,N_7216);
xor U12470 (N_12470,N_7525,N_6435);
nor U12471 (N_12471,N_7811,N_6853);
nor U12472 (N_12472,N_5149,N_9150);
or U12473 (N_12473,N_7115,N_6731);
nand U12474 (N_12474,N_8428,N_8896);
nor U12475 (N_12475,N_9634,N_8619);
and U12476 (N_12476,N_6859,N_9724);
nand U12477 (N_12477,N_6314,N_8456);
or U12478 (N_12478,N_7765,N_5825);
or U12479 (N_12479,N_5532,N_7666);
and U12480 (N_12480,N_7190,N_6101);
and U12481 (N_12481,N_5453,N_7395);
or U12482 (N_12482,N_5694,N_9644);
or U12483 (N_12483,N_8039,N_8478);
and U12484 (N_12484,N_6492,N_6864);
or U12485 (N_12485,N_6894,N_7024);
xor U12486 (N_12486,N_8280,N_8661);
xnor U12487 (N_12487,N_7658,N_9943);
or U12488 (N_12488,N_9181,N_8688);
nand U12489 (N_12489,N_6970,N_7998);
xnor U12490 (N_12490,N_5751,N_5613);
or U12491 (N_12491,N_5912,N_7792);
nand U12492 (N_12492,N_8209,N_7579);
and U12493 (N_12493,N_6416,N_6448);
nand U12494 (N_12494,N_8308,N_9873);
nand U12495 (N_12495,N_8721,N_6911);
nor U12496 (N_12496,N_8200,N_9137);
nand U12497 (N_12497,N_6063,N_6354);
or U12498 (N_12498,N_8885,N_6105);
nand U12499 (N_12499,N_5139,N_9859);
or U12500 (N_12500,N_9735,N_5458);
and U12501 (N_12501,N_7672,N_8710);
xor U12502 (N_12502,N_7835,N_6068);
or U12503 (N_12503,N_8419,N_7757);
nand U12504 (N_12504,N_5876,N_5326);
and U12505 (N_12505,N_7330,N_5635);
xor U12506 (N_12506,N_6999,N_6187);
xor U12507 (N_12507,N_8880,N_6703);
and U12508 (N_12508,N_9387,N_6830);
nor U12509 (N_12509,N_6427,N_8321);
nand U12510 (N_12510,N_8537,N_9901);
nor U12511 (N_12511,N_6986,N_6475);
nand U12512 (N_12512,N_5131,N_8096);
xor U12513 (N_12513,N_6632,N_7792);
nor U12514 (N_12514,N_6881,N_7577);
nand U12515 (N_12515,N_7838,N_6656);
or U12516 (N_12516,N_8400,N_9115);
or U12517 (N_12517,N_9790,N_6908);
or U12518 (N_12518,N_9571,N_5826);
xnor U12519 (N_12519,N_7644,N_8972);
xor U12520 (N_12520,N_6696,N_5655);
and U12521 (N_12521,N_8501,N_7485);
and U12522 (N_12522,N_7092,N_6990);
and U12523 (N_12523,N_6635,N_5273);
nand U12524 (N_12524,N_8105,N_9252);
or U12525 (N_12525,N_8580,N_8053);
nand U12526 (N_12526,N_7591,N_8829);
nand U12527 (N_12527,N_9681,N_7950);
nor U12528 (N_12528,N_6299,N_9333);
or U12529 (N_12529,N_8247,N_5280);
or U12530 (N_12530,N_9197,N_5743);
or U12531 (N_12531,N_5355,N_8560);
nand U12532 (N_12532,N_7836,N_6499);
nand U12533 (N_12533,N_9194,N_7411);
or U12534 (N_12534,N_5080,N_9291);
or U12535 (N_12535,N_7576,N_5529);
and U12536 (N_12536,N_8335,N_9409);
or U12537 (N_12537,N_6576,N_6088);
or U12538 (N_12538,N_6000,N_7364);
and U12539 (N_12539,N_8596,N_8228);
nand U12540 (N_12540,N_7011,N_6960);
xor U12541 (N_12541,N_8693,N_7819);
and U12542 (N_12542,N_6502,N_7593);
or U12543 (N_12543,N_6725,N_9333);
or U12544 (N_12544,N_9141,N_8337);
nor U12545 (N_12545,N_9858,N_9614);
nand U12546 (N_12546,N_5163,N_5082);
and U12547 (N_12547,N_7633,N_7678);
and U12548 (N_12548,N_8872,N_7611);
xor U12549 (N_12549,N_6454,N_7659);
and U12550 (N_12550,N_5730,N_9057);
nor U12551 (N_12551,N_7588,N_6548);
or U12552 (N_12552,N_8762,N_7061);
and U12553 (N_12553,N_9484,N_7562);
or U12554 (N_12554,N_6934,N_6540);
nor U12555 (N_12555,N_7212,N_5113);
or U12556 (N_12556,N_7543,N_7851);
nor U12557 (N_12557,N_7471,N_6188);
xor U12558 (N_12558,N_9435,N_8335);
xnor U12559 (N_12559,N_9735,N_9144);
nand U12560 (N_12560,N_7105,N_9112);
and U12561 (N_12561,N_6872,N_7139);
or U12562 (N_12562,N_9866,N_6478);
or U12563 (N_12563,N_8206,N_8538);
xnor U12564 (N_12564,N_5256,N_7317);
and U12565 (N_12565,N_7610,N_8299);
or U12566 (N_12566,N_6524,N_7709);
nand U12567 (N_12567,N_9557,N_6987);
and U12568 (N_12568,N_5786,N_5991);
nor U12569 (N_12569,N_7701,N_7466);
or U12570 (N_12570,N_6579,N_5066);
and U12571 (N_12571,N_7914,N_7971);
nand U12572 (N_12572,N_7227,N_6780);
and U12573 (N_12573,N_8736,N_5741);
and U12574 (N_12574,N_9398,N_8039);
or U12575 (N_12575,N_7577,N_6743);
and U12576 (N_12576,N_5630,N_6483);
and U12577 (N_12577,N_9051,N_5443);
or U12578 (N_12578,N_5340,N_8456);
nor U12579 (N_12579,N_8803,N_9051);
nand U12580 (N_12580,N_5088,N_8117);
nor U12581 (N_12581,N_7583,N_9870);
nand U12582 (N_12582,N_9543,N_8810);
nand U12583 (N_12583,N_5643,N_6571);
nor U12584 (N_12584,N_6279,N_6419);
nor U12585 (N_12585,N_6461,N_9881);
xnor U12586 (N_12586,N_6184,N_9030);
xnor U12587 (N_12587,N_5812,N_5913);
or U12588 (N_12588,N_5821,N_6836);
nor U12589 (N_12589,N_9977,N_7289);
nor U12590 (N_12590,N_8311,N_5367);
xor U12591 (N_12591,N_7965,N_5265);
xnor U12592 (N_12592,N_7888,N_8036);
xnor U12593 (N_12593,N_9914,N_9699);
xnor U12594 (N_12594,N_7319,N_6876);
nor U12595 (N_12595,N_8918,N_5252);
or U12596 (N_12596,N_6564,N_5653);
nor U12597 (N_12597,N_6719,N_5133);
xnor U12598 (N_12598,N_7060,N_8136);
or U12599 (N_12599,N_5746,N_8505);
nand U12600 (N_12600,N_7374,N_8325);
and U12601 (N_12601,N_9039,N_5008);
xnor U12602 (N_12602,N_8821,N_9217);
nand U12603 (N_12603,N_9828,N_7998);
or U12604 (N_12604,N_6204,N_5448);
nand U12605 (N_12605,N_5206,N_6367);
nand U12606 (N_12606,N_8456,N_7719);
and U12607 (N_12607,N_6871,N_5262);
xnor U12608 (N_12608,N_7674,N_8602);
and U12609 (N_12609,N_8764,N_6955);
nand U12610 (N_12610,N_7869,N_9603);
and U12611 (N_12611,N_6393,N_9175);
nor U12612 (N_12612,N_8912,N_9698);
and U12613 (N_12613,N_8026,N_7546);
or U12614 (N_12614,N_8350,N_6543);
nor U12615 (N_12615,N_7333,N_6413);
or U12616 (N_12616,N_9871,N_5592);
nand U12617 (N_12617,N_5987,N_8157);
nor U12618 (N_12618,N_9512,N_5220);
and U12619 (N_12619,N_8864,N_9078);
or U12620 (N_12620,N_8559,N_7633);
and U12621 (N_12621,N_9711,N_7816);
or U12622 (N_12622,N_8446,N_5866);
nor U12623 (N_12623,N_5206,N_6113);
nor U12624 (N_12624,N_6727,N_9658);
nor U12625 (N_12625,N_6241,N_6012);
nand U12626 (N_12626,N_5925,N_6602);
nand U12627 (N_12627,N_6996,N_6976);
nand U12628 (N_12628,N_5363,N_6000);
nand U12629 (N_12629,N_5246,N_5796);
nand U12630 (N_12630,N_5141,N_9603);
nand U12631 (N_12631,N_8935,N_8877);
nor U12632 (N_12632,N_8808,N_8182);
and U12633 (N_12633,N_9708,N_5399);
xnor U12634 (N_12634,N_9196,N_9288);
nand U12635 (N_12635,N_5225,N_7345);
nand U12636 (N_12636,N_6439,N_6039);
nor U12637 (N_12637,N_7158,N_6506);
nor U12638 (N_12638,N_9685,N_8109);
and U12639 (N_12639,N_7159,N_7823);
nor U12640 (N_12640,N_5828,N_8985);
xor U12641 (N_12641,N_9362,N_9180);
or U12642 (N_12642,N_5755,N_5699);
and U12643 (N_12643,N_6101,N_5659);
and U12644 (N_12644,N_9521,N_9917);
and U12645 (N_12645,N_7857,N_9019);
or U12646 (N_12646,N_9516,N_7897);
xor U12647 (N_12647,N_8810,N_7935);
nor U12648 (N_12648,N_9530,N_5433);
xor U12649 (N_12649,N_9632,N_6596);
nand U12650 (N_12650,N_6733,N_8049);
nand U12651 (N_12651,N_8192,N_9362);
xnor U12652 (N_12652,N_9584,N_9815);
nor U12653 (N_12653,N_7949,N_9116);
nand U12654 (N_12654,N_9884,N_8051);
and U12655 (N_12655,N_8307,N_9276);
nand U12656 (N_12656,N_7186,N_6608);
nand U12657 (N_12657,N_5732,N_6024);
xor U12658 (N_12658,N_5496,N_8888);
and U12659 (N_12659,N_6264,N_6707);
and U12660 (N_12660,N_7695,N_7456);
and U12661 (N_12661,N_8518,N_8730);
nand U12662 (N_12662,N_9799,N_8210);
nor U12663 (N_12663,N_8695,N_6457);
nor U12664 (N_12664,N_6928,N_9272);
nor U12665 (N_12665,N_6521,N_7923);
xor U12666 (N_12666,N_7608,N_5711);
xnor U12667 (N_12667,N_9449,N_9466);
or U12668 (N_12668,N_7358,N_9393);
and U12669 (N_12669,N_8665,N_7098);
and U12670 (N_12670,N_6178,N_8405);
xnor U12671 (N_12671,N_7030,N_6967);
or U12672 (N_12672,N_6861,N_7369);
nor U12673 (N_12673,N_7621,N_8734);
nand U12674 (N_12674,N_7825,N_9154);
xor U12675 (N_12675,N_5922,N_7329);
nor U12676 (N_12676,N_7073,N_8543);
or U12677 (N_12677,N_7893,N_8632);
nand U12678 (N_12678,N_5241,N_5234);
xnor U12679 (N_12679,N_8174,N_9390);
nand U12680 (N_12680,N_5043,N_5281);
nor U12681 (N_12681,N_8349,N_8557);
xor U12682 (N_12682,N_7769,N_8141);
or U12683 (N_12683,N_5660,N_7479);
nand U12684 (N_12684,N_9139,N_9310);
xor U12685 (N_12685,N_5226,N_8565);
nor U12686 (N_12686,N_9107,N_5107);
xnor U12687 (N_12687,N_6605,N_7283);
xor U12688 (N_12688,N_8741,N_6520);
xor U12689 (N_12689,N_9593,N_8632);
or U12690 (N_12690,N_8404,N_6655);
nor U12691 (N_12691,N_5188,N_6329);
and U12692 (N_12692,N_8028,N_9116);
nor U12693 (N_12693,N_7997,N_7940);
nor U12694 (N_12694,N_8414,N_5774);
xnor U12695 (N_12695,N_8314,N_5585);
and U12696 (N_12696,N_9413,N_7024);
or U12697 (N_12697,N_8432,N_7307);
xnor U12698 (N_12698,N_8277,N_8827);
nor U12699 (N_12699,N_7303,N_9626);
nor U12700 (N_12700,N_8691,N_5307);
and U12701 (N_12701,N_9800,N_7423);
xor U12702 (N_12702,N_9851,N_5521);
or U12703 (N_12703,N_6032,N_7584);
xnor U12704 (N_12704,N_6026,N_5073);
xnor U12705 (N_12705,N_5594,N_8705);
nand U12706 (N_12706,N_9348,N_8450);
nor U12707 (N_12707,N_6767,N_6117);
nand U12708 (N_12708,N_8191,N_7501);
nand U12709 (N_12709,N_6941,N_6648);
nand U12710 (N_12710,N_8520,N_6739);
xor U12711 (N_12711,N_6250,N_7265);
nor U12712 (N_12712,N_5329,N_7085);
nand U12713 (N_12713,N_6077,N_6053);
xnor U12714 (N_12714,N_6307,N_6031);
xnor U12715 (N_12715,N_8271,N_8900);
and U12716 (N_12716,N_7456,N_7682);
nor U12717 (N_12717,N_8964,N_6113);
and U12718 (N_12718,N_8110,N_5597);
nor U12719 (N_12719,N_8324,N_6516);
or U12720 (N_12720,N_9729,N_9954);
nand U12721 (N_12721,N_5548,N_8288);
nand U12722 (N_12722,N_5186,N_8007);
xor U12723 (N_12723,N_9551,N_5431);
and U12724 (N_12724,N_7220,N_9765);
nor U12725 (N_12725,N_7902,N_6623);
nand U12726 (N_12726,N_7680,N_9928);
nand U12727 (N_12727,N_5525,N_5146);
xor U12728 (N_12728,N_5874,N_6591);
xnor U12729 (N_12729,N_5519,N_7516);
xnor U12730 (N_12730,N_9349,N_6211);
xor U12731 (N_12731,N_6434,N_9100);
xnor U12732 (N_12732,N_8708,N_9154);
nor U12733 (N_12733,N_8080,N_8654);
and U12734 (N_12734,N_5059,N_7684);
and U12735 (N_12735,N_7884,N_9418);
xor U12736 (N_12736,N_5729,N_9364);
or U12737 (N_12737,N_5876,N_8077);
and U12738 (N_12738,N_5751,N_8618);
nand U12739 (N_12739,N_6253,N_5737);
xnor U12740 (N_12740,N_7892,N_6608);
nand U12741 (N_12741,N_7665,N_8955);
or U12742 (N_12742,N_7254,N_5741);
nand U12743 (N_12743,N_5374,N_6681);
xor U12744 (N_12744,N_6907,N_9813);
and U12745 (N_12745,N_8489,N_8735);
xnor U12746 (N_12746,N_6426,N_6087);
nand U12747 (N_12747,N_9981,N_9174);
nand U12748 (N_12748,N_5544,N_7923);
xnor U12749 (N_12749,N_5937,N_9938);
nor U12750 (N_12750,N_8229,N_8315);
xor U12751 (N_12751,N_8252,N_7846);
nand U12752 (N_12752,N_8282,N_6235);
xor U12753 (N_12753,N_9128,N_5631);
and U12754 (N_12754,N_5768,N_5315);
and U12755 (N_12755,N_6696,N_6582);
xor U12756 (N_12756,N_5409,N_5266);
and U12757 (N_12757,N_9846,N_9175);
nor U12758 (N_12758,N_7369,N_6151);
xor U12759 (N_12759,N_9183,N_8766);
nand U12760 (N_12760,N_7691,N_7562);
nand U12761 (N_12761,N_5358,N_8245);
or U12762 (N_12762,N_7496,N_8174);
and U12763 (N_12763,N_6061,N_6710);
nand U12764 (N_12764,N_6567,N_8366);
or U12765 (N_12765,N_5273,N_8254);
xnor U12766 (N_12766,N_7141,N_6055);
xor U12767 (N_12767,N_7009,N_9844);
or U12768 (N_12768,N_6242,N_6415);
nand U12769 (N_12769,N_9874,N_7546);
xor U12770 (N_12770,N_7318,N_6252);
xnor U12771 (N_12771,N_7766,N_8985);
nand U12772 (N_12772,N_8625,N_7102);
and U12773 (N_12773,N_5367,N_6455);
or U12774 (N_12774,N_5260,N_8700);
nand U12775 (N_12775,N_6193,N_6937);
xor U12776 (N_12776,N_7254,N_6009);
and U12777 (N_12777,N_5353,N_7392);
xor U12778 (N_12778,N_6091,N_6555);
xnor U12779 (N_12779,N_8439,N_5704);
or U12780 (N_12780,N_6996,N_7138);
xnor U12781 (N_12781,N_7538,N_7583);
and U12782 (N_12782,N_9437,N_9282);
xor U12783 (N_12783,N_5291,N_7635);
nor U12784 (N_12784,N_7583,N_7200);
and U12785 (N_12785,N_7686,N_7446);
nand U12786 (N_12786,N_7755,N_6093);
nand U12787 (N_12787,N_8067,N_6476);
nand U12788 (N_12788,N_6600,N_8644);
nand U12789 (N_12789,N_6439,N_6675);
or U12790 (N_12790,N_7515,N_6823);
and U12791 (N_12791,N_7874,N_9848);
and U12792 (N_12792,N_9073,N_6559);
and U12793 (N_12793,N_9017,N_6532);
xor U12794 (N_12794,N_6150,N_9294);
or U12795 (N_12795,N_8841,N_7040);
or U12796 (N_12796,N_7858,N_6533);
xnor U12797 (N_12797,N_8803,N_6150);
nand U12798 (N_12798,N_8262,N_9782);
nor U12799 (N_12799,N_7706,N_7447);
and U12800 (N_12800,N_5048,N_6899);
nand U12801 (N_12801,N_9755,N_7678);
nand U12802 (N_12802,N_7852,N_6585);
nor U12803 (N_12803,N_6069,N_5289);
or U12804 (N_12804,N_6518,N_5132);
and U12805 (N_12805,N_6559,N_6675);
or U12806 (N_12806,N_6739,N_8897);
nor U12807 (N_12807,N_8604,N_9493);
xor U12808 (N_12808,N_8758,N_6893);
xnor U12809 (N_12809,N_6114,N_7597);
xor U12810 (N_12810,N_9744,N_9376);
and U12811 (N_12811,N_9211,N_7075);
xor U12812 (N_12812,N_9449,N_7444);
nand U12813 (N_12813,N_5640,N_8764);
nand U12814 (N_12814,N_9004,N_9113);
or U12815 (N_12815,N_9054,N_7042);
or U12816 (N_12816,N_5129,N_9351);
nor U12817 (N_12817,N_8995,N_7428);
and U12818 (N_12818,N_8097,N_6808);
nor U12819 (N_12819,N_7274,N_7642);
and U12820 (N_12820,N_8580,N_7339);
and U12821 (N_12821,N_9683,N_7688);
xnor U12822 (N_12822,N_5411,N_5871);
nor U12823 (N_12823,N_8861,N_5144);
nand U12824 (N_12824,N_9021,N_6542);
xor U12825 (N_12825,N_6482,N_6801);
xnor U12826 (N_12826,N_7816,N_5994);
or U12827 (N_12827,N_7657,N_6525);
xor U12828 (N_12828,N_7785,N_6311);
nor U12829 (N_12829,N_6952,N_5450);
nor U12830 (N_12830,N_6792,N_7671);
or U12831 (N_12831,N_5835,N_8881);
nand U12832 (N_12832,N_7233,N_7897);
nand U12833 (N_12833,N_6824,N_7160);
xnor U12834 (N_12834,N_8268,N_9499);
or U12835 (N_12835,N_6208,N_8339);
and U12836 (N_12836,N_8143,N_5796);
xnor U12837 (N_12837,N_8566,N_7629);
or U12838 (N_12838,N_6686,N_5186);
xor U12839 (N_12839,N_5032,N_9521);
xnor U12840 (N_12840,N_7473,N_9408);
nor U12841 (N_12841,N_5920,N_5772);
or U12842 (N_12842,N_9090,N_5748);
and U12843 (N_12843,N_9998,N_8368);
xnor U12844 (N_12844,N_6730,N_6004);
or U12845 (N_12845,N_5848,N_6195);
xnor U12846 (N_12846,N_7737,N_6623);
xnor U12847 (N_12847,N_7846,N_5006);
nand U12848 (N_12848,N_7231,N_6401);
nand U12849 (N_12849,N_8895,N_5527);
or U12850 (N_12850,N_5319,N_7113);
nor U12851 (N_12851,N_8386,N_8396);
nand U12852 (N_12852,N_7653,N_5576);
and U12853 (N_12853,N_6201,N_8436);
nand U12854 (N_12854,N_5456,N_5191);
xor U12855 (N_12855,N_7748,N_7177);
xnor U12856 (N_12856,N_8852,N_6001);
nor U12857 (N_12857,N_6960,N_9112);
xor U12858 (N_12858,N_6349,N_7306);
or U12859 (N_12859,N_6457,N_6915);
xnor U12860 (N_12860,N_9961,N_7242);
xor U12861 (N_12861,N_9444,N_9417);
nand U12862 (N_12862,N_5149,N_9147);
nor U12863 (N_12863,N_9753,N_5527);
nand U12864 (N_12864,N_5372,N_8025);
and U12865 (N_12865,N_6914,N_7816);
and U12866 (N_12866,N_8769,N_5176);
nor U12867 (N_12867,N_5950,N_5976);
nor U12868 (N_12868,N_7109,N_7748);
or U12869 (N_12869,N_9090,N_7552);
nand U12870 (N_12870,N_6550,N_9389);
xor U12871 (N_12871,N_5919,N_8268);
xnor U12872 (N_12872,N_7794,N_6019);
nand U12873 (N_12873,N_9999,N_5354);
and U12874 (N_12874,N_5060,N_8757);
xnor U12875 (N_12875,N_6556,N_9002);
or U12876 (N_12876,N_9949,N_5028);
nand U12877 (N_12877,N_8072,N_8399);
nor U12878 (N_12878,N_5388,N_9640);
and U12879 (N_12879,N_6773,N_8975);
xor U12880 (N_12880,N_8666,N_8828);
nor U12881 (N_12881,N_9426,N_9583);
nand U12882 (N_12882,N_6761,N_8974);
or U12883 (N_12883,N_8066,N_7670);
xor U12884 (N_12884,N_9389,N_7524);
xor U12885 (N_12885,N_5136,N_7555);
nand U12886 (N_12886,N_8308,N_7466);
and U12887 (N_12887,N_9509,N_8158);
or U12888 (N_12888,N_5193,N_5434);
nor U12889 (N_12889,N_5549,N_7819);
nor U12890 (N_12890,N_9847,N_5350);
nand U12891 (N_12891,N_9479,N_6438);
or U12892 (N_12892,N_5710,N_9783);
or U12893 (N_12893,N_8219,N_8117);
and U12894 (N_12894,N_5528,N_9244);
xnor U12895 (N_12895,N_5108,N_5268);
xnor U12896 (N_12896,N_5850,N_5324);
nand U12897 (N_12897,N_7755,N_5511);
nand U12898 (N_12898,N_9486,N_9251);
and U12899 (N_12899,N_9685,N_8149);
nand U12900 (N_12900,N_7100,N_7053);
nor U12901 (N_12901,N_6018,N_6341);
xor U12902 (N_12902,N_7527,N_9906);
or U12903 (N_12903,N_9160,N_6114);
nand U12904 (N_12904,N_6871,N_7331);
nand U12905 (N_12905,N_8726,N_7261);
nand U12906 (N_12906,N_7832,N_6357);
nor U12907 (N_12907,N_8012,N_5272);
nand U12908 (N_12908,N_6601,N_5924);
nor U12909 (N_12909,N_6956,N_7023);
xnor U12910 (N_12910,N_9252,N_5985);
or U12911 (N_12911,N_7449,N_7917);
nor U12912 (N_12912,N_8067,N_5772);
nor U12913 (N_12913,N_6773,N_5316);
nand U12914 (N_12914,N_9790,N_9554);
nand U12915 (N_12915,N_5876,N_7218);
and U12916 (N_12916,N_8156,N_5609);
nand U12917 (N_12917,N_8695,N_8908);
xnor U12918 (N_12918,N_6360,N_7219);
and U12919 (N_12919,N_5687,N_7427);
nand U12920 (N_12920,N_9155,N_5820);
and U12921 (N_12921,N_9535,N_9739);
and U12922 (N_12922,N_6349,N_5501);
xor U12923 (N_12923,N_9567,N_7809);
or U12924 (N_12924,N_8222,N_9909);
nand U12925 (N_12925,N_7678,N_5072);
nor U12926 (N_12926,N_8887,N_9085);
nand U12927 (N_12927,N_5079,N_8416);
and U12928 (N_12928,N_7993,N_6910);
nand U12929 (N_12929,N_7105,N_5712);
xor U12930 (N_12930,N_7174,N_8736);
or U12931 (N_12931,N_7756,N_8529);
xor U12932 (N_12932,N_8211,N_9806);
nand U12933 (N_12933,N_8630,N_8122);
or U12934 (N_12934,N_8843,N_8940);
or U12935 (N_12935,N_8979,N_9600);
nor U12936 (N_12936,N_5698,N_6825);
nor U12937 (N_12937,N_6154,N_9007);
nor U12938 (N_12938,N_8025,N_8524);
xor U12939 (N_12939,N_6893,N_8498);
nand U12940 (N_12940,N_9920,N_6789);
or U12941 (N_12941,N_6184,N_6008);
nand U12942 (N_12942,N_6793,N_6041);
nand U12943 (N_12943,N_7525,N_5516);
xor U12944 (N_12944,N_6196,N_5510);
nor U12945 (N_12945,N_7267,N_6413);
and U12946 (N_12946,N_7967,N_6612);
nor U12947 (N_12947,N_7821,N_5512);
and U12948 (N_12948,N_9225,N_7959);
xor U12949 (N_12949,N_9220,N_9687);
nor U12950 (N_12950,N_8020,N_9264);
nor U12951 (N_12951,N_7888,N_5756);
or U12952 (N_12952,N_6154,N_8326);
nand U12953 (N_12953,N_6760,N_8876);
nor U12954 (N_12954,N_9335,N_8296);
or U12955 (N_12955,N_6011,N_5403);
nand U12956 (N_12956,N_7440,N_8322);
and U12957 (N_12957,N_7219,N_6692);
nand U12958 (N_12958,N_7002,N_5492);
xnor U12959 (N_12959,N_8159,N_5127);
or U12960 (N_12960,N_9128,N_5926);
or U12961 (N_12961,N_7101,N_7294);
nand U12962 (N_12962,N_7686,N_9291);
nand U12963 (N_12963,N_9193,N_5860);
nand U12964 (N_12964,N_9864,N_8815);
nor U12965 (N_12965,N_7163,N_9728);
and U12966 (N_12966,N_6763,N_8405);
nand U12967 (N_12967,N_9928,N_7637);
nand U12968 (N_12968,N_6454,N_9143);
and U12969 (N_12969,N_7637,N_7433);
or U12970 (N_12970,N_6949,N_5380);
or U12971 (N_12971,N_8468,N_5134);
nand U12972 (N_12972,N_7413,N_7011);
and U12973 (N_12973,N_9412,N_8782);
nor U12974 (N_12974,N_7214,N_8878);
and U12975 (N_12975,N_5454,N_6178);
nor U12976 (N_12976,N_6216,N_8531);
nor U12977 (N_12977,N_8167,N_6380);
and U12978 (N_12978,N_9429,N_8813);
nor U12979 (N_12979,N_6926,N_6289);
nand U12980 (N_12980,N_9986,N_6279);
nor U12981 (N_12981,N_8914,N_8404);
nor U12982 (N_12982,N_8883,N_8583);
nor U12983 (N_12983,N_8425,N_7898);
xnor U12984 (N_12984,N_6399,N_5063);
nor U12985 (N_12985,N_6293,N_9498);
xor U12986 (N_12986,N_7247,N_9875);
nand U12987 (N_12987,N_5082,N_7681);
and U12988 (N_12988,N_9363,N_8284);
nand U12989 (N_12989,N_8018,N_8344);
or U12990 (N_12990,N_9146,N_5580);
nor U12991 (N_12991,N_5266,N_5050);
and U12992 (N_12992,N_8769,N_8719);
nor U12993 (N_12993,N_8102,N_8786);
xor U12994 (N_12994,N_9129,N_7701);
and U12995 (N_12995,N_9827,N_6507);
and U12996 (N_12996,N_8020,N_6188);
or U12997 (N_12997,N_8228,N_5047);
xnor U12998 (N_12998,N_9908,N_7906);
and U12999 (N_12999,N_9282,N_9507);
and U13000 (N_13000,N_5992,N_5656);
nor U13001 (N_13001,N_7858,N_6753);
and U13002 (N_13002,N_7244,N_9876);
nand U13003 (N_13003,N_7451,N_5269);
and U13004 (N_13004,N_7620,N_6257);
and U13005 (N_13005,N_9923,N_9082);
or U13006 (N_13006,N_9185,N_8683);
nand U13007 (N_13007,N_7476,N_5247);
and U13008 (N_13008,N_6596,N_9644);
or U13009 (N_13009,N_5648,N_6207);
nor U13010 (N_13010,N_6825,N_5156);
nor U13011 (N_13011,N_8159,N_9793);
or U13012 (N_13012,N_9767,N_6727);
nand U13013 (N_13013,N_5065,N_7256);
nor U13014 (N_13014,N_9107,N_8219);
or U13015 (N_13015,N_8615,N_6156);
xnor U13016 (N_13016,N_7452,N_8095);
nor U13017 (N_13017,N_6112,N_5952);
and U13018 (N_13018,N_5619,N_7668);
nor U13019 (N_13019,N_6544,N_6905);
xor U13020 (N_13020,N_5847,N_7493);
nor U13021 (N_13021,N_6752,N_8054);
nor U13022 (N_13022,N_6814,N_9899);
and U13023 (N_13023,N_7409,N_6059);
and U13024 (N_13024,N_5917,N_7560);
nand U13025 (N_13025,N_9318,N_9141);
or U13026 (N_13026,N_9626,N_6559);
and U13027 (N_13027,N_9879,N_5197);
nand U13028 (N_13028,N_5219,N_5012);
or U13029 (N_13029,N_5948,N_5301);
nor U13030 (N_13030,N_6030,N_6516);
or U13031 (N_13031,N_7353,N_7743);
and U13032 (N_13032,N_7584,N_5780);
and U13033 (N_13033,N_6797,N_8098);
nor U13034 (N_13034,N_7589,N_6246);
nand U13035 (N_13035,N_7226,N_6181);
nand U13036 (N_13036,N_6689,N_7350);
and U13037 (N_13037,N_9826,N_9231);
xor U13038 (N_13038,N_5938,N_6227);
xnor U13039 (N_13039,N_5397,N_6105);
xnor U13040 (N_13040,N_7639,N_5399);
nor U13041 (N_13041,N_6580,N_5285);
and U13042 (N_13042,N_7441,N_9154);
xor U13043 (N_13043,N_6817,N_5902);
xnor U13044 (N_13044,N_6922,N_7970);
or U13045 (N_13045,N_5820,N_8364);
nand U13046 (N_13046,N_8654,N_6700);
and U13047 (N_13047,N_5600,N_5632);
nand U13048 (N_13048,N_7297,N_5052);
xnor U13049 (N_13049,N_7614,N_6663);
or U13050 (N_13050,N_7365,N_8437);
and U13051 (N_13051,N_8850,N_9537);
nor U13052 (N_13052,N_9184,N_9272);
and U13053 (N_13053,N_7007,N_7779);
nand U13054 (N_13054,N_9067,N_8624);
nand U13055 (N_13055,N_6155,N_9017);
and U13056 (N_13056,N_5880,N_9810);
xor U13057 (N_13057,N_7023,N_9800);
xor U13058 (N_13058,N_5760,N_6003);
xnor U13059 (N_13059,N_6645,N_8835);
or U13060 (N_13060,N_8807,N_6554);
xnor U13061 (N_13061,N_8611,N_5021);
nand U13062 (N_13062,N_9444,N_7441);
and U13063 (N_13063,N_5551,N_8829);
or U13064 (N_13064,N_5262,N_9561);
or U13065 (N_13065,N_6966,N_7845);
and U13066 (N_13066,N_9435,N_6555);
or U13067 (N_13067,N_7168,N_5591);
nor U13068 (N_13068,N_6552,N_5487);
or U13069 (N_13069,N_7963,N_9909);
and U13070 (N_13070,N_7341,N_5165);
nor U13071 (N_13071,N_9712,N_5930);
or U13072 (N_13072,N_5428,N_9168);
or U13073 (N_13073,N_7405,N_7136);
and U13074 (N_13074,N_9640,N_6544);
nor U13075 (N_13075,N_6757,N_9836);
nor U13076 (N_13076,N_5823,N_7133);
or U13077 (N_13077,N_5088,N_5107);
or U13078 (N_13078,N_9918,N_6535);
nor U13079 (N_13079,N_5269,N_8139);
and U13080 (N_13080,N_8448,N_7833);
nand U13081 (N_13081,N_8680,N_8448);
and U13082 (N_13082,N_5253,N_9516);
nor U13083 (N_13083,N_6772,N_7539);
xnor U13084 (N_13084,N_5109,N_6879);
or U13085 (N_13085,N_8808,N_8770);
nand U13086 (N_13086,N_5651,N_7405);
nand U13087 (N_13087,N_9233,N_9906);
or U13088 (N_13088,N_6267,N_7614);
nor U13089 (N_13089,N_7380,N_5425);
nand U13090 (N_13090,N_5236,N_7597);
nor U13091 (N_13091,N_9501,N_8039);
nand U13092 (N_13092,N_5390,N_6061);
and U13093 (N_13093,N_8798,N_5389);
and U13094 (N_13094,N_5276,N_8096);
xor U13095 (N_13095,N_5838,N_6009);
xor U13096 (N_13096,N_8411,N_9892);
and U13097 (N_13097,N_8822,N_6367);
and U13098 (N_13098,N_7005,N_7995);
nand U13099 (N_13099,N_5054,N_9838);
or U13100 (N_13100,N_9132,N_6127);
xnor U13101 (N_13101,N_7425,N_8033);
nand U13102 (N_13102,N_8370,N_6516);
or U13103 (N_13103,N_6726,N_7903);
and U13104 (N_13104,N_6633,N_5172);
nand U13105 (N_13105,N_5843,N_7051);
xnor U13106 (N_13106,N_9845,N_9239);
nand U13107 (N_13107,N_8082,N_7050);
and U13108 (N_13108,N_6920,N_9174);
or U13109 (N_13109,N_7343,N_8005);
nand U13110 (N_13110,N_5886,N_6124);
or U13111 (N_13111,N_8676,N_9170);
nand U13112 (N_13112,N_9450,N_9592);
and U13113 (N_13113,N_6252,N_8692);
or U13114 (N_13114,N_8487,N_7100);
nand U13115 (N_13115,N_8873,N_8935);
nor U13116 (N_13116,N_5526,N_9324);
and U13117 (N_13117,N_9391,N_7586);
xnor U13118 (N_13118,N_6398,N_7026);
nor U13119 (N_13119,N_7117,N_5966);
or U13120 (N_13120,N_7706,N_5454);
and U13121 (N_13121,N_6176,N_8083);
xor U13122 (N_13122,N_6599,N_8698);
and U13123 (N_13123,N_7919,N_7963);
or U13124 (N_13124,N_7023,N_9371);
and U13125 (N_13125,N_7050,N_9273);
xnor U13126 (N_13126,N_5651,N_5750);
nand U13127 (N_13127,N_7879,N_7710);
xor U13128 (N_13128,N_6146,N_6600);
and U13129 (N_13129,N_7911,N_5459);
nand U13130 (N_13130,N_8780,N_7592);
nand U13131 (N_13131,N_8706,N_7914);
or U13132 (N_13132,N_8644,N_6357);
or U13133 (N_13133,N_5639,N_5504);
nor U13134 (N_13134,N_5245,N_5570);
nand U13135 (N_13135,N_7332,N_7471);
nand U13136 (N_13136,N_8431,N_9249);
xnor U13137 (N_13137,N_5424,N_7058);
or U13138 (N_13138,N_8235,N_6589);
or U13139 (N_13139,N_7348,N_8970);
nor U13140 (N_13140,N_7074,N_9282);
xnor U13141 (N_13141,N_5863,N_8968);
nand U13142 (N_13142,N_9560,N_8321);
xor U13143 (N_13143,N_5021,N_6340);
and U13144 (N_13144,N_5380,N_8463);
and U13145 (N_13145,N_8013,N_5908);
xnor U13146 (N_13146,N_9061,N_8575);
and U13147 (N_13147,N_7995,N_8094);
and U13148 (N_13148,N_5059,N_6089);
xor U13149 (N_13149,N_6428,N_7992);
nor U13150 (N_13150,N_7852,N_9859);
nor U13151 (N_13151,N_5391,N_7330);
nor U13152 (N_13152,N_5968,N_5657);
nand U13153 (N_13153,N_7757,N_7024);
and U13154 (N_13154,N_8545,N_6253);
nor U13155 (N_13155,N_8026,N_6607);
or U13156 (N_13156,N_8875,N_7086);
nor U13157 (N_13157,N_7214,N_7874);
and U13158 (N_13158,N_6270,N_5306);
nand U13159 (N_13159,N_8454,N_7929);
xnor U13160 (N_13160,N_6818,N_7371);
and U13161 (N_13161,N_9372,N_5892);
nand U13162 (N_13162,N_5696,N_8643);
nor U13163 (N_13163,N_5104,N_6996);
nor U13164 (N_13164,N_9529,N_8682);
xnor U13165 (N_13165,N_6626,N_9804);
or U13166 (N_13166,N_8297,N_5100);
xor U13167 (N_13167,N_5490,N_6779);
nor U13168 (N_13168,N_9406,N_6585);
xnor U13169 (N_13169,N_9145,N_9111);
or U13170 (N_13170,N_8398,N_6655);
xor U13171 (N_13171,N_5133,N_5058);
and U13172 (N_13172,N_8882,N_9938);
xnor U13173 (N_13173,N_9690,N_9483);
nand U13174 (N_13174,N_6762,N_6832);
or U13175 (N_13175,N_6598,N_7510);
xor U13176 (N_13176,N_7613,N_7551);
xor U13177 (N_13177,N_5911,N_8438);
xor U13178 (N_13178,N_7909,N_9661);
or U13179 (N_13179,N_9345,N_5989);
or U13180 (N_13180,N_8134,N_9457);
nand U13181 (N_13181,N_6007,N_5781);
or U13182 (N_13182,N_5136,N_8073);
and U13183 (N_13183,N_8609,N_6601);
nand U13184 (N_13184,N_8500,N_6662);
or U13185 (N_13185,N_5614,N_7858);
nor U13186 (N_13186,N_5201,N_5732);
nand U13187 (N_13187,N_8485,N_6467);
nand U13188 (N_13188,N_5327,N_9005);
nand U13189 (N_13189,N_6849,N_7289);
nand U13190 (N_13190,N_8779,N_6018);
and U13191 (N_13191,N_6116,N_7361);
or U13192 (N_13192,N_9192,N_8014);
or U13193 (N_13193,N_7961,N_9214);
xor U13194 (N_13194,N_7136,N_5173);
nand U13195 (N_13195,N_8647,N_8905);
and U13196 (N_13196,N_6723,N_9099);
nor U13197 (N_13197,N_9875,N_7073);
nand U13198 (N_13198,N_9354,N_5754);
nor U13199 (N_13199,N_6114,N_6375);
nand U13200 (N_13200,N_9609,N_6777);
and U13201 (N_13201,N_9020,N_6903);
nand U13202 (N_13202,N_5894,N_9776);
xnor U13203 (N_13203,N_9958,N_7389);
xnor U13204 (N_13204,N_6527,N_8777);
or U13205 (N_13205,N_7164,N_7454);
or U13206 (N_13206,N_8902,N_5432);
nor U13207 (N_13207,N_7418,N_5497);
nand U13208 (N_13208,N_9172,N_6366);
nor U13209 (N_13209,N_7671,N_7536);
or U13210 (N_13210,N_8878,N_5376);
nand U13211 (N_13211,N_7933,N_8045);
and U13212 (N_13212,N_6444,N_7911);
nor U13213 (N_13213,N_5537,N_7810);
or U13214 (N_13214,N_9884,N_6870);
xor U13215 (N_13215,N_5737,N_5395);
or U13216 (N_13216,N_5352,N_7538);
xnor U13217 (N_13217,N_9006,N_7829);
xor U13218 (N_13218,N_6097,N_8588);
xnor U13219 (N_13219,N_6150,N_9429);
nand U13220 (N_13220,N_5644,N_9497);
or U13221 (N_13221,N_6234,N_9298);
nand U13222 (N_13222,N_7610,N_6864);
nor U13223 (N_13223,N_6075,N_5911);
and U13224 (N_13224,N_6201,N_5526);
xnor U13225 (N_13225,N_8739,N_6630);
or U13226 (N_13226,N_5139,N_6065);
and U13227 (N_13227,N_6938,N_8381);
nand U13228 (N_13228,N_8721,N_6774);
nor U13229 (N_13229,N_5982,N_8004);
nor U13230 (N_13230,N_6365,N_6379);
xor U13231 (N_13231,N_5751,N_8537);
nand U13232 (N_13232,N_6303,N_8722);
nor U13233 (N_13233,N_6086,N_6835);
xor U13234 (N_13234,N_7684,N_7226);
nor U13235 (N_13235,N_5168,N_5045);
and U13236 (N_13236,N_6979,N_6039);
nand U13237 (N_13237,N_7383,N_8795);
xnor U13238 (N_13238,N_6048,N_6031);
xnor U13239 (N_13239,N_7221,N_9518);
or U13240 (N_13240,N_6083,N_7335);
nor U13241 (N_13241,N_9109,N_5710);
or U13242 (N_13242,N_8839,N_6105);
xnor U13243 (N_13243,N_5864,N_8328);
nand U13244 (N_13244,N_8169,N_7101);
nand U13245 (N_13245,N_7156,N_7832);
nand U13246 (N_13246,N_9877,N_6762);
xnor U13247 (N_13247,N_5653,N_5299);
or U13248 (N_13248,N_6417,N_9395);
nand U13249 (N_13249,N_9627,N_5509);
xor U13250 (N_13250,N_8694,N_9245);
and U13251 (N_13251,N_5811,N_7151);
and U13252 (N_13252,N_9162,N_6865);
xor U13253 (N_13253,N_9144,N_6457);
nor U13254 (N_13254,N_5580,N_5268);
and U13255 (N_13255,N_7082,N_7939);
and U13256 (N_13256,N_7728,N_6899);
and U13257 (N_13257,N_8694,N_6258);
xnor U13258 (N_13258,N_7725,N_6819);
and U13259 (N_13259,N_6456,N_9570);
and U13260 (N_13260,N_6488,N_5304);
nor U13261 (N_13261,N_7249,N_7508);
nand U13262 (N_13262,N_5299,N_8314);
nor U13263 (N_13263,N_5006,N_5286);
nand U13264 (N_13264,N_7569,N_7871);
and U13265 (N_13265,N_7589,N_6748);
and U13266 (N_13266,N_9433,N_9864);
xnor U13267 (N_13267,N_8355,N_7696);
and U13268 (N_13268,N_6859,N_9017);
and U13269 (N_13269,N_9536,N_8916);
or U13270 (N_13270,N_7857,N_5141);
nor U13271 (N_13271,N_8755,N_9571);
or U13272 (N_13272,N_7413,N_5975);
nand U13273 (N_13273,N_7355,N_8486);
nor U13274 (N_13274,N_9704,N_8730);
nand U13275 (N_13275,N_5550,N_9813);
xor U13276 (N_13276,N_6177,N_5836);
nor U13277 (N_13277,N_6709,N_9235);
nand U13278 (N_13278,N_6623,N_5286);
nor U13279 (N_13279,N_7589,N_7893);
or U13280 (N_13280,N_8868,N_6595);
or U13281 (N_13281,N_7439,N_5464);
or U13282 (N_13282,N_6884,N_9579);
nand U13283 (N_13283,N_6505,N_5576);
and U13284 (N_13284,N_8259,N_5362);
nor U13285 (N_13285,N_5280,N_9474);
nand U13286 (N_13286,N_9600,N_6609);
nor U13287 (N_13287,N_5998,N_6340);
or U13288 (N_13288,N_5307,N_6854);
nor U13289 (N_13289,N_5122,N_6399);
or U13290 (N_13290,N_6651,N_6124);
nand U13291 (N_13291,N_7931,N_7485);
nor U13292 (N_13292,N_8124,N_9349);
xnor U13293 (N_13293,N_8793,N_9432);
nor U13294 (N_13294,N_5570,N_7908);
xnor U13295 (N_13295,N_9370,N_5943);
and U13296 (N_13296,N_7522,N_8721);
xnor U13297 (N_13297,N_7056,N_7755);
nor U13298 (N_13298,N_8474,N_5339);
xor U13299 (N_13299,N_9769,N_7867);
and U13300 (N_13300,N_9962,N_6461);
nor U13301 (N_13301,N_8432,N_5779);
xor U13302 (N_13302,N_6500,N_6046);
xnor U13303 (N_13303,N_7870,N_9388);
nor U13304 (N_13304,N_5608,N_7299);
or U13305 (N_13305,N_5382,N_6164);
or U13306 (N_13306,N_9135,N_7162);
nor U13307 (N_13307,N_9569,N_9833);
nor U13308 (N_13308,N_7080,N_9947);
or U13309 (N_13309,N_6995,N_8753);
and U13310 (N_13310,N_5977,N_5499);
nor U13311 (N_13311,N_8947,N_6381);
or U13312 (N_13312,N_8704,N_7637);
nor U13313 (N_13313,N_8077,N_6607);
nand U13314 (N_13314,N_8998,N_9568);
nand U13315 (N_13315,N_8413,N_9201);
and U13316 (N_13316,N_8142,N_8268);
nand U13317 (N_13317,N_7673,N_8747);
and U13318 (N_13318,N_8856,N_9338);
nor U13319 (N_13319,N_8020,N_9064);
nand U13320 (N_13320,N_7471,N_7243);
and U13321 (N_13321,N_7242,N_8544);
and U13322 (N_13322,N_9653,N_7712);
or U13323 (N_13323,N_8897,N_9684);
and U13324 (N_13324,N_8283,N_5116);
xor U13325 (N_13325,N_5275,N_6183);
nor U13326 (N_13326,N_9323,N_6685);
nor U13327 (N_13327,N_9426,N_5255);
nor U13328 (N_13328,N_5724,N_7725);
nand U13329 (N_13329,N_9890,N_7188);
nand U13330 (N_13330,N_5191,N_8178);
nand U13331 (N_13331,N_5656,N_9668);
or U13332 (N_13332,N_5794,N_7591);
xnor U13333 (N_13333,N_5621,N_8541);
nand U13334 (N_13334,N_6956,N_6718);
xor U13335 (N_13335,N_8729,N_6674);
or U13336 (N_13336,N_9601,N_7848);
xor U13337 (N_13337,N_5566,N_8497);
or U13338 (N_13338,N_8961,N_7838);
xnor U13339 (N_13339,N_9415,N_5225);
or U13340 (N_13340,N_6723,N_5271);
and U13341 (N_13341,N_5012,N_5887);
xor U13342 (N_13342,N_9576,N_8883);
or U13343 (N_13343,N_8479,N_6392);
nor U13344 (N_13344,N_9106,N_8680);
nor U13345 (N_13345,N_9063,N_7814);
nand U13346 (N_13346,N_5013,N_9580);
and U13347 (N_13347,N_5550,N_6217);
nor U13348 (N_13348,N_7939,N_9897);
nand U13349 (N_13349,N_8689,N_6330);
nor U13350 (N_13350,N_8237,N_7243);
nand U13351 (N_13351,N_7315,N_6360);
xnor U13352 (N_13352,N_9054,N_7119);
nor U13353 (N_13353,N_8769,N_6323);
xor U13354 (N_13354,N_8189,N_8455);
nor U13355 (N_13355,N_8961,N_9416);
xnor U13356 (N_13356,N_7322,N_5652);
nor U13357 (N_13357,N_6653,N_8181);
or U13358 (N_13358,N_9054,N_6038);
or U13359 (N_13359,N_8426,N_8848);
xor U13360 (N_13360,N_5880,N_6229);
or U13361 (N_13361,N_6599,N_9580);
xnor U13362 (N_13362,N_7905,N_9394);
or U13363 (N_13363,N_8526,N_5166);
nand U13364 (N_13364,N_9599,N_7012);
nor U13365 (N_13365,N_9086,N_6694);
and U13366 (N_13366,N_6539,N_9079);
and U13367 (N_13367,N_8623,N_9132);
xnor U13368 (N_13368,N_6708,N_7388);
or U13369 (N_13369,N_7940,N_9728);
or U13370 (N_13370,N_7076,N_6340);
nand U13371 (N_13371,N_9486,N_5968);
nor U13372 (N_13372,N_6487,N_5461);
and U13373 (N_13373,N_9351,N_9711);
xor U13374 (N_13374,N_8049,N_7611);
xnor U13375 (N_13375,N_5127,N_7172);
xnor U13376 (N_13376,N_7332,N_8875);
or U13377 (N_13377,N_9118,N_9546);
nand U13378 (N_13378,N_8419,N_6082);
xnor U13379 (N_13379,N_9164,N_7351);
and U13380 (N_13380,N_8915,N_9225);
or U13381 (N_13381,N_7423,N_9028);
xor U13382 (N_13382,N_8679,N_7911);
nand U13383 (N_13383,N_6186,N_9207);
and U13384 (N_13384,N_5769,N_7612);
xor U13385 (N_13385,N_5576,N_6012);
and U13386 (N_13386,N_8083,N_9485);
and U13387 (N_13387,N_7301,N_8014);
or U13388 (N_13388,N_6513,N_6406);
nor U13389 (N_13389,N_7139,N_6883);
nand U13390 (N_13390,N_5621,N_5934);
nor U13391 (N_13391,N_6080,N_5840);
nand U13392 (N_13392,N_7613,N_5076);
nor U13393 (N_13393,N_6201,N_5524);
xnor U13394 (N_13394,N_6969,N_9452);
or U13395 (N_13395,N_5165,N_9412);
nand U13396 (N_13396,N_8116,N_8324);
or U13397 (N_13397,N_6165,N_9949);
nand U13398 (N_13398,N_7003,N_6658);
nand U13399 (N_13399,N_7524,N_6181);
nand U13400 (N_13400,N_8044,N_9607);
nand U13401 (N_13401,N_9861,N_5404);
and U13402 (N_13402,N_5129,N_5744);
nor U13403 (N_13403,N_7377,N_6169);
and U13404 (N_13404,N_9147,N_6621);
xor U13405 (N_13405,N_6425,N_5805);
nand U13406 (N_13406,N_5068,N_7636);
xnor U13407 (N_13407,N_5866,N_7695);
xnor U13408 (N_13408,N_9258,N_8497);
or U13409 (N_13409,N_7468,N_9944);
and U13410 (N_13410,N_7801,N_5424);
or U13411 (N_13411,N_9379,N_5982);
nand U13412 (N_13412,N_6734,N_7391);
and U13413 (N_13413,N_7585,N_7160);
and U13414 (N_13414,N_6656,N_6911);
nor U13415 (N_13415,N_5598,N_9650);
or U13416 (N_13416,N_8258,N_5639);
nor U13417 (N_13417,N_6050,N_6195);
nand U13418 (N_13418,N_7051,N_7986);
or U13419 (N_13419,N_5500,N_8544);
nand U13420 (N_13420,N_7045,N_9139);
nand U13421 (N_13421,N_6986,N_7654);
xnor U13422 (N_13422,N_6872,N_9102);
or U13423 (N_13423,N_6136,N_6265);
xor U13424 (N_13424,N_8030,N_9224);
and U13425 (N_13425,N_7331,N_5019);
xor U13426 (N_13426,N_7739,N_9178);
and U13427 (N_13427,N_5817,N_6387);
and U13428 (N_13428,N_7848,N_8825);
nor U13429 (N_13429,N_7843,N_6080);
xnor U13430 (N_13430,N_5000,N_6865);
and U13431 (N_13431,N_7003,N_6024);
nand U13432 (N_13432,N_9568,N_7322);
or U13433 (N_13433,N_6834,N_5721);
or U13434 (N_13434,N_6662,N_8387);
nand U13435 (N_13435,N_9691,N_9035);
nor U13436 (N_13436,N_7324,N_7884);
or U13437 (N_13437,N_6958,N_5731);
nor U13438 (N_13438,N_5808,N_7647);
or U13439 (N_13439,N_7471,N_9488);
xnor U13440 (N_13440,N_8479,N_9860);
or U13441 (N_13441,N_6285,N_8817);
xnor U13442 (N_13442,N_8330,N_9317);
nor U13443 (N_13443,N_5740,N_7269);
nor U13444 (N_13444,N_5958,N_8267);
nand U13445 (N_13445,N_9105,N_9446);
and U13446 (N_13446,N_6172,N_5209);
nand U13447 (N_13447,N_5893,N_5335);
nor U13448 (N_13448,N_8231,N_6244);
and U13449 (N_13449,N_6430,N_5886);
or U13450 (N_13450,N_5847,N_9437);
nor U13451 (N_13451,N_9374,N_7655);
and U13452 (N_13452,N_9775,N_8538);
nand U13453 (N_13453,N_5666,N_5433);
xnor U13454 (N_13454,N_7785,N_7099);
and U13455 (N_13455,N_5659,N_8555);
and U13456 (N_13456,N_8144,N_8457);
nor U13457 (N_13457,N_5898,N_5450);
and U13458 (N_13458,N_5196,N_9112);
and U13459 (N_13459,N_6944,N_9890);
and U13460 (N_13460,N_7539,N_9183);
nor U13461 (N_13461,N_9911,N_7591);
or U13462 (N_13462,N_6939,N_5118);
xnor U13463 (N_13463,N_8190,N_5817);
xor U13464 (N_13464,N_7208,N_7958);
and U13465 (N_13465,N_7402,N_9305);
and U13466 (N_13466,N_5597,N_7684);
xor U13467 (N_13467,N_9044,N_9656);
nor U13468 (N_13468,N_6698,N_6256);
and U13469 (N_13469,N_6859,N_8632);
and U13470 (N_13470,N_7300,N_5469);
or U13471 (N_13471,N_7436,N_5226);
or U13472 (N_13472,N_6621,N_7656);
or U13473 (N_13473,N_7883,N_8458);
nand U13474 (N_13474,N_9822,N_5560);
nand U13475 (N_13475,N_5079,N_5463);
xor U13476 (N_13476,N_6321,N_5468);
nor U13477 (N_13477,N_6774,N_9051);
or U13478 (N_13478,N_9335,N_7870);
nand U13479 (N_13479,N_9567,N_5596);
or U13480 (N_13480,N_6856,N_9230);
nand U13481 (N_13481,N_6447,N_8477);
and U13482 (N_13482,N_7400,N_8244);
or U13483 (N_13483,N_9370,N_9310);
and U13484 (N_13484,N_6193,N_8745);
or U13485 (N_13485,N_5045,N_8043);
and U13486 (N_13486,N_7749,N_7347);
and U13487 (N_13487,N_7068,N_5537);
nor U13488 (N_13488,N_7213,N_7262);
or U13489 (N_13489,N_5620,N_8063);
nor U13490 (N_13490,N_5793,N_6162);
and U13491 (N_13491,N_6302,N_8890);
or U13492 (N_13492,N_7289,N_5394);
or U13493 (N_13493,N_7819,N_9792);
xnor U13494 (N_13494,N_7918,N_7495);
xor U13495 (N_13495,N_9603,N_9451);
xor U13496 (N_13496,N_6646,N_7728);
nand U13497 (N_13497,N_6063,N_6328);
and U13498 (N_13498,N_7278,N_6892);
nor U13499 (N_13499,N_8226,N_7459);
xor U13500 (N_13500,N_7214,N_6053);
xor U13501 (N_13501,N_9528,N_8403);
or U13502 (N_13502,N_5873,N_6171);
xnor U13503 (N_13503,N_7388,N_8986);
nand U13504 (N_13504,N_9066,N_9239);
nor U13505 (N_13505,N_6391,N_9964);
nor U13506 (N_13506,N_9177,N_8857);
and U13507 (N_13507,N_5647,N_9876);
nor U13508 (N_13508,N_9699,N_8224);
xor U13509 (N_13509,N_7262,N_5075);
nor U13510 (N_13510,N_8989,N_9303);
or U13511 (N_13511,N_8585,N_6181);
and U13512 (N_13512,N_9107,N_5385);
and U13513 (N_13513,N_6102,N_9907);
or U13514 (N_13514,N_9739,N_7844);
nand U13515 (N_13515,N_9085,N_9865);
or U13516 (N_13516,N_5007,N_7981);
xor U13517 (N_13517,N_7601,N_9675);
xor U13518 (N_13518,N_5291,N_6821);
or U13519 (N_13519,N_8747,N_8705);
and U13520 (N_13520,N_8282,N_7766);
nand U13521 (N_13521,N_8108,N_6196);
nor U13522 (N_13522,N_7382,N_9646);
nand U13523 (N_13523,N_8660,N_9953);
and U13524 (N_13524,N_5146,N_6884);
and U13525 (N_13525,N_5229,N_5745);
xor U13526 (N_13526,N_9138,N_9712);
and U13527 (N_13527,N_8933,N_8397);
and U13528 (N_13528,N_9371,N_8343);
nand U13529 (N_13529,N_6556,N_8237);
nand U13530 (N_13530,N_6489,N_7224);
or U13531 (N_13531,N_6409,N_5733);
xor U13532 (N_13532,N_6497,N_6518);
nor U13533 (N_13533,N_9203,N_6830);
or U13534 (N_13534,N_7575,N_8565);
nor U13535 (N_13535,N_9637,N_5181);
nor U13536 (N_13536,N_5292,N_6003);
xor U13537 (N_13537,N_5917,N_7783);
nor U13538 (N_13538,N_8107,N_8812);
or U13539 (N_13539,N_8596,N_6089);
nand U13540 (N_13540,N_8506,N_9434);
xor U13541 (N_13541,N_8649,N_6966);
nor U13542 (N_13542,N_5209,N_9827);
and U13543 (N_13543,N_7908,N_6304);
or U13544 (N_13544,N_8998,N_6198);
xor U13545 (N_13545,N_5613,N_7476);
and U13546 (N_13546,N_7897,N_6479);
nand U13547 (N_13547,N_5077,N_5671);
and U13548 (N_13548,N_6174,N_8334);
or U13549 (N_13549,N_7426,N_5559);
nor U13550 (N_13550,N_9793,N_7560);
or U13551 (N_13551,N_9303,N_8858);
and U13552 (N_13552,N_5394,N_7472);
xnor U13553 (N_13553,N_5102,N_8721);
xnor U13554 (N_13554,N_6860,N_8642);
and U13555 (N_13555,N_5706,N_7421);
nand U13556 (N_13556,N_9134,N_8374);
and U13557 (N_13557,N_7469,N_7804);
or U13558 (N_13558,N_9018,N_8264);
nand U13559 (N_13559,N_9467,N_8580);
nand U13560 (N_13560,N_6570,N_7183);
and U13561 (N_13561,N_6074,N_7200);
nor U13562 (N_13562,N_9101,N_8256);
or U13563 (N_13563,N_7772,N_6123);
nor U13564 (N_13564,N_5381,N_7709);
xor U13565 (N_13565,N_8182,N_9452);
and U13566 (N_13566,N_5549,N_9772);
nor U13567 (N_13567,N_6627,N_8516);
nand U13568 (N_13568,N_7284,N_8564);
or U13569 (N_13569,N_9533,N_5086);
nor U13570 (N_13570,N_8061,N_9346);
nand U13571 (N_13571,N_7670,N_7508);
nand U13572 (N_13572,N_9944,N_9395);
and U13573 (N_13573,N_7883,N_6013);
nor U13574 (N_13574,N_7433,N_7494);
and U13575 (N_13575,N_7455,N_8274);
or U13576 (N_13576,N_8868,N_6436);
nor U13577 (N_13577,N_7558,N_7065);
xnor U13578 (N_13578,N_6539,N_9244);
nor U13579 (N_13579,N_6910,N_9255);
nor U13580 (N_13580,N_7353,N_8873);
and U13581 (N_13581,N_8570,N_5305);
nor U13582 (N_13582,N_6785,N_5159);
nand U13583 (N_13583,N_6138,N_6942);
or U13584 (N_13584,N_7874,N_6631);
and U13585 (N_13585,N_7281,N_8911);
and U13586 (N_13586,N_6309,N_8828);
xor U13587 (N_13587,N_6336,N_6395);
and U13588 (N_13588,N_7390,N_5640);
nor U13589 (N_13589,N_6257,N_5529);
and U13590 (N_13590,N_5463,N_6330);
or U13591 (N_13591,N_7548,N_9562);
nand U13592 (N_13592,N_5421,N_6131);
and U13593 (N_13593,N_6429,N_9438);
nor U13594 (N_13594,N_8477,N_7430);
and U13595 (N_13595,N_8742,N_8641);
nand U13596 (N_13596,N_7275,N_6645);
xor U13597 (N_13597,N_8681,N_8231);
nor U13598 (N_13598,N_7032,N_7860);
nor U13599 (N_13599,N_7965,N_9678);
and U13600 (N_13600,N_7552,N_6773);
xnor U13601 (N_13601,N_7297,N_9078);
nand U13602 (N_13602,N_7980,N_8083);
nor U13603 (N_13603,N_5128,N_6899);
xnor U13604 (N_13604,N_5290,N_8913);
nand U13605 (N_13605,N_5945,N_8146);
xnor U13606 (N_13606,N_9960,N_5674);
xor U13607 (N_13607,N_7791,N_6028);
nand U13608 (N_13608,N_6030,N_6539);
or U13609 (N_13609,N_6742,N_6758);
or U13610 (N_13610,N_8976,N_5414);
nand U13611 (N_13611,N_6004,N_8096);
and U13612 (N_13612,N_8145,N_6375);
xor U13613 (N_13613,N_5907,N_8658);
nor U13614 (N_13614,N_8373,N_6886);
nand U13615 (N_13615,N_5484,N_8179);
nor U13616 (N_13616,N_7977,N_5501);
xor U13617 (N_13617,N_5041,N_9338);
and U13618 (N_13618,N_7619,N_6459);
and U13619 (N_13619,N_6608,N_7097);
or U13620 (N_13620,N_8520,N_7817);
and U13621 (N_13621,N_9240,N_7549);
xor U13622 (N_13622,N_5131,N_5308);
and U13623 (N_13623,N_8428,N_8884);
xnor U13624 (N_13624,N_8283,N_6403);
and U13625 (N_13625,N_9075,N_6146);
nand U13626 (N_13626,N_7905,N_5612);
xor U13627 (N_13627,N_7109,N_6034);
nor U13628 (N_13628,N_5510,N_8713);
or U13629 (N_13629,N_5015,N_8426);
and U13630 (N_13630,N_5731,N_8911);
or U13631 (N_13631,N_5954,N_5804);
and U13632 (N_13632,N_6968,N_7737);
nor U13633 (N_13633,N_6845,N_5428);
and U13634 (N_13634,N_8749,N_9488);
nor U13635 (N_13635,N_7200,N_8463);
xnor U13636 (N_13636,N_8682,N_9006);
nand U13637 (N_13637,N_5032,N_6322);
nand U13638 (N_13638,N_6528,N_6424);
and U13639 (N_13639,N_8242,N_5264);
nand U13640 (N_13640,N_9831,N_5529);
or U13641 (N_13641,N_5908,N_8107);
and U13642 (N_13642,N_6806,N_7589);
nand U13643 (N_13643,N_8296,N_9084);
and U13644 (N_13644,N_7943,N_6024);
or U13645 (N_13645,N_6981,N_5014);
xnor U13646 (N_13646,N_6355,N_5590);
and U13647 (N_13647,N_7320,N_8422);
or U13648 (N_13648,N_6594,N_5008);
nor U13649 (N_13649,N_6407,N_7266);
nand U13650 (N_13650,N_9108,N_5965);
or U13651 (N_13651,N_6480,N_5555);
nor U13652 (N_13652,N_6280,N_8953);
nor U13653 (N_13653,N_6848,N_6135);
nor U13654 (N_13654,N_9957,N_6856);
nor U13655 (N_13655,N_6278,N_9205);
nor U13656 (N_13656,N_8357,N_9697);
xnor U13657 (N_13657,N_5142,N_7649);
and U13658 (N_13658,N_7633,N_9995);
nor U13659 (N_13659,N_5871,N_6455);
or U13660 (N_13660,N_7667,N_8440);
or U13661 (N_13661,N_9595,N_7185);
nand U13662 (N_13662,N_8944,N_7315);
nor U13663 (N_13663,N_6937,N_8143);
xnor U13664 (N_13664,N_8014,N_6510);
nor U13665 (N_13665,N_6853,N_5422);
nor U13666 (N_13666,N_6034,N_7694);
nor U13667 (N_13667,N_7205,N_5886);
nand U13668 (N_13668,N_9034,N_8988);
xnor U13669 (N_13669,N_5763,N_9828);
nor U13670 (N_13670,N_8351,N_8945);
and U13671 (N_13671,N_9817,N_5382);
and U13672 (N_13672,N_7285,N_8700);
and U13673 (N_13673,N_6389,N_9965);
nor U13674 (N_13674,N_8173,N_6472);
nand U13675 (N_13675,N_8732,N_8144);
nand U13676 (N_13676,N_9552,N_6379);
xnor U13677 (N_13677,N_8120,N_6881);
or U13678 (N_13678,N_9096,N_6055);
nor U13679 (N_13679,N_7941,N_6847);
nand U13680 (N_13680,N_6740,N_8811);
nor U13681 (N_13681,N_6116,N_9339);
nand U13682 (N_13682,N_9096,N_6698);
nor U13683 (N_13683,N_5960,N_9972);
or U13684 (N_13684,N_7289,N_7302);
and U13685 (N_13685,N_6719,N_7828);
xnor U13686 (N_13686,N_5002,N_8372);
or U13687 (N_13687,N_9561,N_6053);
nor U13688 (N_13688,N_5762,N_5895);
and U13689 (N_13689,N_8212,N_7983);
nor U13690 (N_13690,N_7254,N_8422);
nor U13691 (N_13691,N_7096,N_7063);
nand U13692 (N_13692,N_6798,N_6892);
nand U13693 (N_13693,N_7491,N_7259);
or U13694 (N_13694,N_6886,N_7964);
nor U13695 (N_13695,N_5023,N_8816);
nor U13696 (N_13696,N_5168,N_7749);
nor U13697 (N_13697,N_6992,N_7743);
nand U13698 (N_13698,N_9477,N_9042);
or U13699 (N_13699,N_8758,N_5008);
or U13700 (N_13700,N_9433,N_5866);
nand U13701 (N_13701,N_7908,N_6217);
nand U13702 (N_13702,N_6177,N_8434);
and U13703 (N_13703,N_6696,N_5808);
nor U13704 (N_13704,N_5221,N_6399);
or U13705 (N_13705,N_9916,N_5787);
or U13706 (N_13706,N_7303,N_9297);
or U13707 (N_13707,N_6724,N_9356);
xnor U13708 (N_13708,N_9205,N_7087);
xnor U13709 (N_13709,N_9105,N_9902);
or U13710 (N_13710,N_7960,N_8467);
and U13711 (N_13711,N_6776,N_9492);
and U13712 (N_13712,N_6071,N_7045);
xor U13713 (N_13713,N_6583,N_7101);
nand U13714 (N_13714,N_6793,N_5735);
nand U13715 (N_13715,N_5105,N_5074);
nand U13716 (N_13716,N_9198,N_6461);
nand U13717 (N_13717,N_8735,N_9430);
and U13718 (N_13718,N_5863,N_6118);
xnor U13719 (N_13719,N_9224,N_8730);
nand U13720 (N_13720,N_9675,N_9245);
xnor U13721 (N_13721,N_9215,N_6274);
nand U13722 (N_13722,N_6239,N_8597);
xnor U13723 (N_13723,N_5645,N_6379);
nand U13724 (N_13724,N_7935,N_5384);
xnor U13725 (N_13725,N_7433,N_6452);
and U13726 (N_13726,N_7633,N_6055);
or U13727 (N_13727,N_8723,N_6719);
nor U13728 (N_13728,N_6781,N_7581);
nand U13729 (N_13729,N_5416,N_7264);
nor U13730 (N_13730,N_7631,N_5560);
xnor U13731 (N_13731,N_9361,N_7655);
and U13732 (N_13732,N_9913,N_6961);
or U13733 (N_13733,N_8170,N_7581);
and U13734 (N_13734,N_5918,N_8070);
or U13735 (N_13735,N_8695,N_7338);
and U13736 (N_13736,N_7226,N_9812);
and U13737 (N_13737,N_6820,N_5766);
xor U13738 (N_13738,N_6349,N_7909);
nor U13739 (N_13739,N_8463,N_9537);
and U13740 (N_13740,N_7261,N_7887);
and U13741 (N_13741,N_5078,N_9532);
nor U13742 (N_13742,N_6839,N_5536);
nand U13743 (N_13743,N_5948,N_5455);
xor U13744 (N_13744,N_9620,N_8948);
nor U13745 (N_13745,N_8122,N_9306);
nand U13746 (N_13746,N_7660,N_6544);
and U13747 (N_13747,N_7466,N_5382);
xnor U13748 (N_13748,N_5072,N_8132);
nand U13749 (N_13749,N_9341,N_7774);
nor U13750 (N_13750,N_9509,N_7973);
and U13751 (N_13751,N_5120,N_8366);
or U13752 (N_13752,N_9005,N_5570);
and U13753 (N_13753,N_7526,N_5540);
nor U13754 (N_13754,N_8208,N_7722);
nand U13755 (N_13755,N_7821,N_9320);
nor U13756 (N_13756,N_7249,N_5864);
xor U13757 (N_13757,N_6379,N_5390);
xnor U13758 (N_13758,N_6143,N_6869);
xor U13759 (N_13759,N_6809,N_7562);
xor U13760 (N_13760,N_9379,N_7750);
nor U13761 (N_13761,N_6031,N_5145);
nor U13762 (N_13762,N_6904,N_7038);
xor U13763 (N_13763,N_6476,N_8036);
xor U13764 (N_13764,N_6842,N_6702);
xnor U13765 (N_13765,N_7207,N_7562);
nand U13766 (N_13766,N_7450,N_7070);
or U13767 (N_13767,N_9140,N_5390);
or U13768 (N_13768,N_8496,N_7416);
xnor U13769 (N_13769,N_8511,N_5363);
nand U13770 (N_13770,N_9036,N_6341);
xnor U13771 (N_13771,N_6383,N_9420);
nand U13772 (N_13772,N_5126,N_7631);
nor U13773 (N_13773,N_8581,N_7146);
or U13774 (N_13774,N_7812,N_7820);
xor U13775 (N_13775,N_9351,N_8626);
xor U13776 (N_13776,N_5973,N_6490);
and U13777 (N_13777,N_8872,N_9096);
xor U13778 (N_13778,N_7830,N_9428);
xnor U13779 (N_13779,N_8062,N_6247);
and U13780 (N_13780,N_6897,N_6790);
nor U13781 (N_13781,N_9816,N_7741);
and U13782 (N_13782,N_7913,N_7399);
nand U13783 (N_13783,N_6131,N_5440);
and U13784 (N_13784,N_7272,N_7110);
or U13785 (N_13785,N_9084,N_5229);
xnor U13786 (N_13786,N_7138,N_6658);
and U13787 (N_13787,N_7401,N_7627);
nor U13788 (N_13788,N_6913,N_5337);
xor U13789 (N_13789,N_6155,N_6380);
nand U13790 (N_13790,N_9852,N_6532);
xor U13791 (N_13791,N_9790,N_6636);
xnor U13792 (N_13792,N_5005,N_9553);
nand U13793 (N_13793,N_7025,N_8439);
or U13794 (N_13794,N_7895,N_8357);
nand U13795 (N_13795,N_7348,N_5003);
xor U13796 (N_13796,N_9560,N_7863);
nor U13797 (N_13797,N_7253,N_7390);
xnor U13798 (N_13798,N_6612,N_5415);
nand U13799 (N_13799,N_9472,N_9450);
xor U13800 (N_13800,N_8845,N_5477);
nor U13801 (N_13801,N_5588,N_7707);
and U13802 (N_13802,N_8703,N_8620);
nand U13803 (N_13803,N_5684,N_7890);
or U13804 (N_13804,N_9788,N_6928);
nor U13805 (N_13805,N_8264,N_5265);
and U13806 (N_13806,N_6901,N_8933);
xor U13807 (N_13807,N_6695,N_7189);
and U13808 (N_13808,N_5451,N_7209);
and U13809 (N_13809,N_9795,N_9221);
or U13810 (N_13810,N_9778,N_7870);
xor U13811 (N_13811,N_5310,N_5762);
nor U13812 (N_13812,N_9356,N_5550);
xnor U13813 (N_13813,N_6305,N_9738);
and U13814 (N_13814,N_6122,N_6724);
and U13815 (N_13815,N_7858,N_5528);
or U13816 (N_13816,N_8720,N_8566);
or U13817 (N_13817,N_6878,N_5044);
and U13818 (N_13818,N_6437,N_6711);
nand U13819 (N_13819,N_8241,N_7762);
nand U13820 (N_13820,N_8969,N_9061);
xnor U13821 (N_13821,N_6780,N_7448);
xnor U13822 (N_13822,N_8881,N_9800);
xor U13823 (N_13823,N_8309,N_7535);
nand U13824 (N_13824,N_5134,N_7655);
xor U13825 (N_13825,N_6109,N_5739);
xor U13826 (N_13826,N_8417,N_7983);
and U13827 (N_13827,N_5825,N_9678);
nor U13828 (N_13828,N_8336,N_8811);
nand U13829 (N_13829,N_7705,N_8067);
xor U13830 (N_13830,N_6019,N_5419);
xor U13831 (N_13831,N_7303,N_9091);
or U13832 (N_13832,N_8077,N_9578);
xor U13833 (N_13833,N_9549,N_9869);
xor U13834 (N_13834,N_7570,N_5654);
xnor U13835 (N_13835,N_9816,N_5538);
nand U13836 (N_13836,N_9310,N_6102);
nor U13837 (N_13837,N_9110,N_7342);
and U13838 (N_13838,N_5485,N_5504);
nand U13839 (N_13839,N_6430,N_9779);
and U13840 (N_13840,N_5111,N_5841);
xnor U13841 (N_13841,N_9640,N_5415);
nor U13842 (N_13842,N_5458,N_5820);
and U13843 (N_13843,N_9334,N_7129);
and U13844 (N_13844,N_8253,N_6263);
and U13845 (N_13845,N_5773,N_8562);
or U13846 (N_13846,N_7452,N_8673);
nand U13847 (N_13847,N_5816,N_8778);
and U13848 (N_13848,N_9711,N_5742);
xnor U13849 (N_13849,N_9598,N_8774);
and U13850 (N_13850,N_9798,N_7156);
xnor U13851 (N_13851,N_5763,N_8686);
or U13852 (N_13852,N_8687,N_7380);
nand U13853 (N_13853,N_6941,N_8575);
nor U13854 (N_13854,N_9417,N_6080);
nor U13855 (N_13855,N_7025,N_7854);
or U13856 (N_13856,N_5350,N_6641);
xnor U13857 (N_13857,N_8313,N_8545);
xor U13858 (N_13858,N_6395,N_5409);
or U13859 (N_13859,N_5569,N_7946);
and U13860 (N_13860,N_8621,N_5062);
nor U13861 (N_13861,N_7870,N_8305);
nor U13862 (N_13862,N_7318,N_8315);
or U13863 (N_13863,N_7724,N_8955);
nor U13864 (N_13864,N_5519,N_6265);
nand U13865 (N_13865,N_7843,N_5599);
xor U13866 (N_13866,N_6126,N_9584);
nor U13867 (N_13867,N_5732,N_9436);
and U13868 (N_13868,N_5079,N_5061);
and U13869 (N_13869,N_5040,N_7581);
or U13870 (N_13870,N_6282,N_5162);
xnor U13871 (N_13871,N_7619,N_7498);
nand U13872 (N_13872,N_8037,N_6003);
nand U13873 (N_13873,N_9821,N_6125);
or U13874 (N_13874,N_6096,N_5405);
nor U13875 (N_13875,N_5959,N_6752);
nand U13876 (N_13876,N_8927,N_7168);
or U13877 (N_13877,N_5618,N_7608);
or U13878 (N_13878,N_9811,N_5228);
or U13879 (N_13879,N_7227,N_7112);
or U13880 (N_13880,N_6039,N_9101);
nor U13881 (N_13881,N_6944,N_7350);
and U13882 (N_13882,N_6567,N_7362);
or U13883 (N_13883,N_5685,N_6865);
nor U13884 (N_13884,N_5450,N_6290);
and U13885 (N_13885,N_9570,N_9566);
nor U13886 (N_13886,N_6709,N_9119);
or U13887 (N_13887,N_7654,N_5637);
nor U13888 (N_13888,N_6474,N_7682);
nand U13889 (N_13889,N_9333,N_7025);
xor U13890 (N_13890,N_5847,N_6070);
nor U13891 (N_13891,N_9475,N_8003);
nor U13892 (N_13892,N_7900,N_5114);
or U13893 (N_13893,N_8527,N_8598);
xnor U13894 (N_13894,N_9651,N_9975);
xnor U13895 (N_13895,N_7896,N_9293);
nor U13896 (N_13896,N_9642,N_7048);
and U13897 (N_13897,N_7261,N_7796);
xor U13898 (N_13898,N_8714,N_5260);
xnor U13899 (N_13899,N_6380,N_5513);
nor U13900 (N_13900,N_6412,N_5294);
nor U13901 (N_13901,N_7200,N_5673);
nor U13902 (N_13902,N_8918,N_8551);
xnor U13903 (N_13903,N_5402,N_7071);
nor U13904 (N_13904,N_7142,N_5642);
nor U13905 (N_13905,N_7679,N_6024);
nand U13906 (N_13906,N_9357,N_9874);
and U13907 (N_13907,N_7804,N_8436);
xnor U13908 (N_13908,N_5324,N_7216);
nor U13909 (N_13909,N_9342,N_9013);
and U13910 (N_13910,N_9705,N_9478);
or U13911 (N_13911,N_6868,N_6671);
nor U13912 (N_13912,N_5359,N_8621);
xor U13913 (N_13913,N_7826,N_8774);
nand U13914 (N_13914,N_6322,N_6921);
or U13915 (N_13915,N_7988,N_9661);
nand U13916 (N_13916,N_8969,N_8829);
nor U13917 (N_13917,N_9377,N_7649);
nor U13918 (N_13918,N_7638,N_7903);
or U13919 (N_13919,N_6049,N_9904);
nand U13920 (N_13920,N_9248,N_6832);
xor U13921 (N_13921,N_5788,N_7962);
and U13922 (N_13922,N_5986,N_7819);
nor U13923 (N_13923,N_6143,N_5235);
xor U13924 (N_13924,N_5840,N_5703);
xor U13925 (N_13925,N_6843,N_5732);
nor U13926 (N_13926,N_8360,N_8367);
and U13927 (N_13927,N_9662,N_6080);
or U13928 (N_13928,N_7941,N_7228);
and U13929 (N_13929,N_8936,N_5230);
and U13930 (N_13930,N_9528,N_8252);
nor U13931 (N_13931,N_7855,N_6618);
xor U13932 (N_13932,N_5581,N_6293);
nor U13933 (N_13933,N_5077,N_9202);
or U13934 (N_13934,N_9214,N_9124);
xor U13935 (N_13935,N_6811,N_8358);
xnor U13936 (N_13936,N_6473,N_5265);
and U13937 (N_13937,N_5888,N_7392);
xnor U13938 (N_13938,N_5279,N_5432);
or U13939 (N_13939,N_9547,N_5492);
or U13940 (N_13940,N_7423,N_7220);
xor U13941 (N_13941,N_5462,N_8234);
nor U13942 (N_13942,N_7186,N_8415);
and U13943 (N_13943,N_5747,N_6617);
and U13944 (N_13944,N_9470,N_5265);
or U13945 (N_13945,N_8202,N_8779);
xor U13946 (N_13946,N_7455,N_5018);
nand U13947 (N_13947,N_7495,N_8917);
and U13948 (N_13948,N_9638,N_6701);
nor U13949 (N_13949,N_8092,N_8067);
nor U13950 (N_13950,N_6392,N_9488);
and U13951 (N_13951,N_5371,N_9450);
xor U13952 (N_13952,N_9845,N_9461);
nand U13953 (N_13953,N_5298,N_7696);
and U13954 (N_13954,N_8844,N_8476);
and U13955 (N_13955,N_9032,N_8167);
nand U13956 (N_13956,N_9200,N_6968);
xor U13957 (N_13957,N_7675,N_9997);
and U13958 (N_13958,N_9932,N_9830);
or U13959 (N_13959,N_8168,N_9222);
xor U13960 (N_13960,N_6580,N_8287);
nor U13961 (N_13961,N_7453,N_6027);
or U13962 (N_13962,N_8634,N_5057);
or U13963 (N_13963,N_7189,N_7406);
nand U13964 (N_13964,N_7476,N_6939);
nand U13965 (N_13965,N_7240,N_6393);
nand U13966 (N_13966,N_7653,N_7603);
or U13967 (N_13967,N_7842,N_7176);
or U13968 (N_13968,N_8392,N_6797);
xor U13969 (N_13969,N_6109,N_8476);
or U13970 (N_13970,N_7230,N_5010);
or U13971 (N_13971,N_7809,N_9022);
nor U13972 (N_13972,N_5567,N_5920);
nor U13973 (N_13973,N_8804,N_8492);
nor U13974 (N_13974,N_7609,N_6749);
xnor U13975 (N_13975,N_7727,N_6131);
nor U13976 (N_13976,N_8548,N_6152);
and U13977 (N_13977,N_6899,N_8824);
xnor U13978 (N_13978,N_6687,N_9037);
nor U13979 (N_13979,N_5736,N_9826);
nor U13980 (N_13980,N_7121,N_6451);
xor U13981 (N_13981,N_6797,N_9475);
nand U13982 (N_13982,N_5565,N_6894);
xnor U13983 (N_13983,N_5180,N_7204);
or U13984 (N_13984,N_8695,N_9450);
nand U13985 (N_13985,N_7336,N_9461);
and U13986 (N_13986,N_9017,N_6060);
or U13987 (N_13987,N_5705,N_5228);
nor U13988 (N_13988,N_5847,N_6444);
xor U13989 (N_13989,N_8583,N_5391);
nor U13990 (N_13990,N_9478,N_7087);
nor U13991 (N_13991,N_5236,N_8221);
xor U13992 (N_13992,N_9904,N_9656);
or U13993 (N_13993,N_7178,N_7536);
or U13994 (N_13994,N_9506,N_8830);
nand U13995 (N_13995,N_9649,N_9549);
and U13996 (N_13996,N_9334,N_9534);
or U13997 (N_13997,N_6652,N_5470);
or U13998 (N_13998,N_5630,N_7443);
xnor U13999 (N_13999,N_8561,N_5038);
or U14000 (N_14000,N_7395,N_6441);
or U14001 (N_14001,N_7303,N_6093);
xor U14002 (N_14002,N_8604,N_8422);
nand U14003 (N_14003,N_5751,N_9361);
nand U14004 (N_14004,N_6959,N_9762);
nor U14005 (N_14005,N_9759,N_9950);
or U14006 (N_14006,N_6639,N_6676);
nand U14007 (N_14007,N_8359,N_8914);
xor U14008 (N_14008,N_6030,N_7510);
or U14009 (N_14009,N_6852,N_7513);
or U14010 (N_14010,N_5700,N_6151);
or U14011 (N_14011,N_5179,N_7778);
or U14012 (N_14012,N_5183,N_9964);
xor U14013 (N_14013,N_9982,N_7694);
and U14014 (N_14014,N_6158,N_7634);
or U14015 (N_14015,N_9451,N_9717);
and U14016 (N_14016,N_5273,N_5516);
nor U14017 (N_14017,N_6659,N_6486);
xor U14018 (N_14018,N_7830,N_6693);
or U14019 (N_14019,N_7050,N_9623);
xor U14020 (N_14020,N_5267,N_5144);
nand U14021 (N_14021,N_5508,N_9995);
or U14022 (N_14022,N_5834,N_5543);
nand U14023 (N_14023,N_6852,N_7786);
nand U14024 (N_14024,N_6271,N_6058);
nand U14025 (N_14025,N_9044,N_5388);
nand U14026 (N_14026,N_5731,N_7182);
or U14027 (N_14027,N_8696,N_7393);
xor U14028 (N_14028,N_9241,N_6477);
xnor U14029 (N_14029,N_9097,N_8439);
xor U14030 (N_14030,N_6525,N_5418);
nand U14031 (N_14031,N_6259,N_9451);
or U14032 (N_14032,N_8647,N_7161);
and U14033 (N_14033,N_6493,N_9822);
xor U14034 (N_14034,N_8629,N_5987);
nand U14035 (N_14035,N_9519,N_9366);
xnor U14036 (N_14036,N_8470,N_6946);
nand U14037 (N_14037,N_7657,N_7899);
and U14038 (N_14038,N_9208,N_5333);
or U14039 (N_14039,N_8233,N_9752);
or U14040 (N_14040,N_5143,N_6631);
or U14041 (N_14041,N_8008,N_6630);
and U14042 (N_14042,N_6995,N_5603);
or U14043 (N_14043,N_7837,N_9759);
or U14044 (N_14044,N_5043,N_7794);
xor U14045 (N_14045,N_5968,N_9436);
or U14046 (N_14046,N_6400,N_6744);
or U14047 (N_14047,N_8042,N_8645);
and U14048 (N_14048,N_5338,N_6384);
nor U14049 (N_14049,N_5606,N_8695);
nor U14050 (N_14050,N_9846,N_6083);
xnor U14051 (N_14051,N_8769,N_7947);
nand U14052 (N_14052,N_8474,N_7231);
xor U14053 (N_14053,N_9890,N_8986);
xnor U14054 (N_14054,N_7451,N_7532);
nand U14055 (N_14055,N_8803,N_7855);
nand U14056 (N_14056,N_9080,N_8946);
and U14057 (N_14057,N_9831,N_6934);
nand U14058 (N_14058,N_9126,N_9521);
xor U14059 (N_14059,N_9453,N_8845);
and U14060 (N_14060,N_7355,N_7661);
xnor U14061 (N_14061,N_6938,N_8473);
nor U14062 (N_14062,N_6039,N_6541);
or U14063 (N_14063,N_5983,N_6835);
nand U14064 (N_14064,N_7923,N_5065);
nor U14065 (N_14065,N_6284,N_7538);
xnor U14066 (N_14066,N_6297,N_6145);
nand U14067 (N_14067,N_9115,N_6871);
nor U14068 (N_14068,N_6115,N_9679);
and U14069 (N_14069,N_6240,N_5685);
nor U14070 (N_14070,N_5873,N_5486);
nor U14071 (N_14071,N_5861,N_7978);
xnor U14072 (N_14072,N_9040,N_6793);
nand U14073 (N_14073,N_8384,N_6814);
nor U14074 (N_14074,N_9133,N_5197);
or U14075 (N_14075,N_7117,N_9545);
and U14076 (N_14076,N_9607,N_5297);
nand U14077 (N_14077,N_5996,N_5607);
nor U14078 (N_14078,N_8856,N_7214);
nor U14079 (N_14079,N_7703,N_7800);
nand U14080 (N_14080,N_7082,N_9213);
nor U14081 (N_14081,N_6251,N_5045);
and U14082 (N_14082,N_8613,N_9189);
or U14083 (N_14083,N_6328,N_9193);
and U14084 (N_14084,N_9911,N_8992);
nor U14085 (N_14085,N_8571,N_6631);
and U14086 (N_14086,N_7532,N_6725);
or U14087 (N_14087,N_7723,N_6730);
nor U14088 (N_14088,N_9397,N_5982);
or U14089 (N_14089,N_7252,N_8013);
xnor U14090 (N_14090,N_5564,N_7323);
nor U14091 (N_14091,N_8865,N_7363);
and U14092 (N_14092,N_8589,N_6253);
nand U14093 (N_14093,N_5409,N_9366);
and U14094 (N_14094,N_9928,N_9044);
nor U14095 (N_14095,N_5628,N_9791);
nand U14096 (N_14096,N_9906,N_8166);
nor U14097 (N_14097,N_5876,N_9140);
or U14098 (N_14098,N_8048,N_7686);
or U14099 (N_14099,N_7074,N_7144);
nor U14100 (N_14100,N_9706,N_5545);
xnor U14101 (N_14101,N_6854,N_9999);
nor U14102 (N_14102,N_6347,N_5119);
nand U14103 (N_14103,N_9062,N_7472);
xnor U14104 (N_14104,N_9369,N_7154);
and U14105 (N_14105,N_8562,N_7558);
or U14106 (N_14106,N_8860,N_7527);
or U14107 (N_14107,N_5025,N_9035);
and U14108 (N_14108,N_9278,N_7694);
nor U14109 (N_14109,N_7225,N_7030);
xor U14110 (N_14110,N_6651,N_9433);
xor U14111 (N_14111,N_9420,N_6203);
nor U14112 (N_14112,N_9873,N_8278);
and U14113 (N_14113,N_9607,N_7753);
and U14114 (N_14114,N_5342,N_7347);
or U14115 (N_14115,N_8968,N_8111);
and U14116 (N_14116,N_6925,N_9091);
xor U14117 (N_14117,N_5127,N_5953);
xor U14118 (N_14118,N_8094,N_6246);
or U14119 (N_14119,N_9963,N_6103);
and U14120 (N_14120,N_7809,N_7591);
nand U14121 (N_14121,N_9272,N_7993);
or U14122 (N_14122,N_5967,N_7702);
nor U14123 (N_14123,N_9316,N_7120);
nand U14124 (N_14124,N_5357,N_7192);
xor U14125 (N_14125,N_5667,N_9953);
nor U14126 (N_14126,N_9310,N_5927);
nor U14127 (N_14127,N_7484,N_6430);
and U14128 (N_14128,N_9993,N_8299);
xor U14129 (N_14129,N_8084,N_6155);
nand U14130 (N_14130,N_7866,N_8639);
nor U14131 (N_14131,N_9662,N_6394);
xor U14132 (N_14132,N_8974,N_7223);
or U14133 (N_14133,N_9671,N_6688);
xnor U14134 (N_14134,N_9910,N_8333);
or U14135 (N_14135,N_7609,N_5925);
nand U14136 (N_14136,N_5116,N_6042);
nor U14137 (N_14137,N_8935,N_5383);
xnor U14138 (N_14138,N_8058,N_9496);
and U14139 (N_14139,N_7558,N_8183);
or U14140 (N_14140,N_7320,N_6639);
nand U14141 (N_14141,N_5380,N_9715);
or U14142 (N_14142,N_7016,N_6044);
nand U14143 (N_14143,N_6485,N_5548);
nand U14144 (N_14144,N_8006,N_5352);
and U14145 (N_14145,N_7171,N_7200);
nand U14146 (N_14146,N_5957,N_9554);
nor U14147 (N_14147,N_5020,N_5558);
xor U14148 (N_14148,N_5026,N_8254);
nor U14149 (N_14149,N_7931,N_7250);
nor U14150 (N_14150,N_6289,N_6160);
and U14151 (N_14151,N_8686,N_6934);
nor U14152 (N_14152,N_7093,N_7594);
or U14153 (N_14153,N_9243,N_8367);
or U14154 (N_14154,N_6642,N_7331);
nor U14155 (N_14155,N_5221,N_7745);
nor U14156 (N_14156,N_5559,N_6949);
xnor U14157 (N_14157,N_8820,N_9640);
nand U14158 (N_14158,N_9649,N_8439);
nor U14159 (N_14159,N_9492,N_6152);
nor U14160 (N_14160,N_9038,N_5727);
nor U14161 (N_14161,N_7102,N_5585);
or U14162 (N_14162,N_7476,N_7449);
xor U14163 (N_14163,N_8544,N_9614);
or U14164 (N_14164,N_9785,N_9493);
or U14165 (N_14165,N_9508,N_7042);
nor U14166 (N_14166,N_9678,N_9677);
nand U14167 (N_14167,N_7658,N_5816);
or U14168 (N_14168,N_9819,N_9781);
nor U14169 (N_14169,N_8535,N_9674);
and U14170 (N_14170,N_7162,N_7741);
xnor U14171 (N_14171,N_6450,N_7766);
or U14172 (N_14172,N_6983,N_5504);
nor U14173 (N_14173,N_6518,N_5527);
and U14174 (N_14174,N_8026,N_8283);
or U14175 (N_14175,N_6351,N_8421);
or U14176 (N_14176,N_5630,N_8032);
and U14177 (N_14177,N_5089,N_8313);
nor U14178 (N_14178,N_8933,N_5918);
nand U14179 (N_14179,N_9580,N_6554);
and U14180 (N_14180,N_5821,N_6915);
nor U14181 (N_14181,N_7205,N_8580);
nor U14182 (N_14182,N_9559,N_9861);
nor U14183 (N_14183,N_9522,N_6572);
or U14184 (N_14184,N_7753,N_8785);
xnor U14185 (N_14185,N_5811,N_9743);
and U14186 (N_14186,N_8584,N_8496);
nand U14187 (N_14187,N_6123,N_5514);
xnor U14188 (N_14188,N_8689,N_9576);
or U14189 (N_14189,N_7580,N_8969);
xor U14190 (N_14190,N_8403,N_6960);
nand U14191 (N_14191,N_6261,N_7055);
xnor U14192 (N_14192,N_9831,N_9080);
and U14193 (N_14193,N_8408,N_9675);
nand U14194 (N_14194,N_8065,N_8750);
nand U14195 (N_14195,N_8347,N_7444);
or U14196 (N_14196,N_9855,N_9653);
xor U14197 (N_14197,N_5994,N_5777);
nor U14198 (N_14198,N_9453,N_8584);
nor U14199 (N_14199,N_7779,N_6549);
nand U14200 (N_14200,N_8371,N_7917);
nor U14201 (N_14201,N_9642,N_6165);
nand U14202 (N_14202,N_6427,N_7113);
xor U14203 (N_14203,N_9531,N_6591);
nand U14204 (N_14204,N_6293,N_9474);
nor U14205 (N_14205,N_5635,N_5603);
nand U14206 (N_14206,N_9246,N_5944);
nor U14207 (N_14207,N_7513,N_5488);
and U14208 (N_14208,N_9626,N_9268);
xnor U14209 (N_14209,N_6438,N_7976);
nor U14210 (N_14210,N_9577,N_5837);
xnor U14211 (N_14211,N_7256,N_9847);
xnor U14212 (N_14212,N_6521,N_7742);
xnor U14213 (N_14213,N_7256,N_7968);
and U14214 (N_14214,N_6454,N_6590);
and U14215 (N_14215,N_6332,N_5033);
and U14216 (N_14216,N_9805,N_5581);
nor U14217 (N_14217,N_7707,N_7987);
and U14218 (N_14218,N_5196,N_6425);
nor U14219 (N_14219,N_9391,N_5981);
or U14220 (N_14220,N_6500,N_9944);
and U14221 (N_14221,N_6885,N_6653);
nand U14222 (N_14222,N_5823,N_7728);
nand U14223 (N_14223,N_6576,N_5133);
nand U14224 (N_14224,N_5562,N_8384);
nand U14225 (N_14225,N_9845,N_8637);
xnor U14226 (N_14226,N_5790,N_6266);
nand U14227 (N_14227,N_8025,N_7077);
or U14228 (N_14228,N_8914,N_7811);
nand U14229 (N_14229,N_9702,N_5220);
nand U14230 (N_14230,N_6801,N_6607);
nand U14231 (N_14231,N_6496,N_9665);
nor U14232 (N_14232,N_8610,N_7464);
xnor U14233 (N_14233,N_5728,N_9386);
or U14234 (N_14234,N_9177,N_5186);
and U14235 (N_14235,N_6207,N_7572);
nand U14236 (N_14236,N_6349,N_8063);
nor U14237 (N_14237,N_8446,N_7063);
nand U14238 (N_14238,N_6010,N_8963);
and U14239 (N_14239,N_7161,N_7152);
and U14240 (N_14240,N_7589,N_9968);
nand U14241 (N_14241,N_6766,N_7202);
nor U14242 (N_14242,N_8777,N_5123);
nand U14243 (N_14243,N_7031,N_9744);
or U14244 (N_14244,N_7893,N_5883);
or U14245 (N_14245,N_8831,N_9217);
xor U14246 (N_14246,N_6861,N_5518);
nor U14247 (N_14247,N_5540,N_9241);
xor U14248 (N_14248,N_7789,N_6850);
nand U14249 (N_14249,N_6596,N_6708);
nand U14250 (N_14250,N_9430,N_8847);
or U14251 (N_14251,N_7746,N_5310);
and U14252 (N_14252,N_8908,N_9455);
or U14253 (N_14253,N_7506,N_7728);
and U14254 (N_14254,N_6652,N_5863);
and U14255 (N_14255,N_5204,N_5681);
and U14256 (N_14256,N_8313,N_9654);
and U14257 (N_14257,N_8867,N_7571);
nand U14258 (N_14258,N_6313,N_6239);
nor U14259 (N_14259,N_5607,N_9275);
nor U14260 (N_14260,N_6133,N_8363);
and U14261 (N_14261,N_8179,N_7036);
and U14262 (N_14262,N_6327,N_9182);
xor U14263 (N_14263,N_6135,N_5387);
or U14264 (N_14264,N_6348,N_7385);
nor U14265 (N_14265,N_9838,N_7015);
and U14266 (N_14266,N_7620,N_6819);
xnor U14267 (N_14267,N_8501,N_5715);
and U14268 (N_14268,N_8962,N_7707);
or U14269 (N_14269,N_7725,N_6604);
or U14270 (N_14270,N_7703,N_7682);
nor U14271 (N_14271,N_6562,N_8340);
and U14272 (N_14272,N_5581,N_7727);
nand U14273 (N_14273,N_9711,N_6272);
and U14274 (N_14274,N_5549,N_7371);
and U14275 (N_14275,N_8303,N_7189);
or U14276 (N_14276,N_9976,N_5347);
or U14277 (N_14277,N_9805,N_9015);
xor U14278 (N_14278,N_7685,N_9956);
nand U14279 (N_14279,N_6471,N_5420);
nand U14280 (N_14280,N_6384,N_7400);
xnor U14281 (N_14281,N_7325,N_6960);
nor U14282 (N_14282,N_8336,N_7505);
xnor U14283 (N_14283,N_7820,N_6995);
and U14284 (N_14284,N_6824,N_7497);
nor U14285 (N_14285,N_5787,N_9796);
xor U14286 (N_14286,N_9550,N_9653);
and U14287 (N_14287,N_5590,N_5220);
nor U14288 (N_14288,N_8180,N_8715);
or U14289 (N_14289,N_6809,N_6761);
xnor U14290 (N_14290,N_5943,N_6339);
or U14291 (N_14291,N_8543,N_9286);
or U14292 (N_14292,N_7001,N_8847);
nor U14293 (N_14293,N_5663,N_5321);
nand U14294 (N_14294,N_5472,N_5347);
nand U14295 (N_14295,N_5484,N_5314);
xor U14296 (N_14296,N_7847,N_6168);
and U14297 (N_14297,N_9530,N_6565);
nand U14298 (N_14298,N_7097,N_9933);
nor U14299 (N_14299,N_9376,N_6319);
nor U14300 (N_14300,N_9242,N_9763);
or U14301 (N_14301,N_8201,N_9702);
nand U14302 (N_14302,N_7940,N_9795);
nand U14303 (N_14303,N_9605,N_5465);
xnor U14304 (N_14304,N_9705,N_8873);
xnor U14305 (N_14305,N_7945,N_9507);
xor U14306 (N_14306,N_5927,N_5701);
and U14307 (N_14307,N_8445,N_5798);
or U14308 (N_14308,N_7393,N_9224);
nor U14309 (N_14309,N_6716,N_5075);
or U14310 (N_14310,N_8160,N_5111);
nor U14311 (N_14311,N_7499,N_8285);
or U14312 (N_14312,N_6633,N_6018);
xnor U14313 (N_14313,N_8495,N_9321);
nand U14314 (N_14314,N_7343,N_9768);
and U14315 (N_14315,N_5303,N_9516);
and U14316 (N_14316,N_6266,N_8038);
or U14317 (N_14317,N_6557,N_8756);
nor U14318 (N_14318,N_5412,N_7496);
and U14319 (N_14319,N_9881,N_7226);
or U14320 (N_14320,N_7778,N_6057);
nor U14321 (N_14321,N_5478,N_7628);
and U14322 (N_14322,N_5306,N_9060);
xor U14323 (N_14323,N_7742,N_9759);
or U14324 (N_14324,N_5061,N_7338);
and U14325 (N_14325,N_8837,N_9352);
nand U14326 (N_14326,N_5394,N_5104);
nand U14327 (N_14327,N_5204,N_8215);
xor U14328 (N_14328,N_6404,N_7882);
xnor U14329 (N_14329,N_9317,N_5554);
nand U14330 (N_14330,N_6867,N_6498);
or U14331 (N_14331,N_7100,N_9848);
nor U14332 (N_14332,N_9628,N_6649);
xor U14333 (N_14333,N_9236,N_6885);
or U14334 (N_14334,N_6383,N_9976);
xnor U14335 (N_14335,N_7392,N_7976);
or U14336 (N_14336,N_9745,N_8401);
nand U14337 (N_14337,N_9243,N_9020);
nand U14338 (N_14338,N_8059,N_9733);
nand U14339 (N_14339,N_6020,N_9812);
and U14340 (N_14340,N_8679,N_8335);
xnor U14341 (N_14341,N_9040,N_6130);
nand U14342 (N_14342,N_8494,N_7381);
nand U14343 (N_14343,N_9803,N_5447);
nand U14344 (N_14344,N_7911,N_9262);
nor U14345 (N_14345,N_8350,N_8325);
nor U14346 (N_14346,N_8881,N_7890);
nor U14347 (N_14347,N_6054,N_8553);
xor U14348 (N_14348,N_8527,N_8081);
and U14349 (N_14349,N_5567,N_9144);
nand U14350 (N_14350,N_8685,N_5393);
or U14351 (N_14351,N_7850,N_9134);
nor U14352 (N_14352,N_9414,N_9915);
xnor U14353 (N_14353,N_9901,N_9422);
or U14354 (N_14354,N_8034,N_9862);
nor U14355 (N_14355,N_6037,N_9588);
xor U14356 (N_14356,N_9078,N_9758);
and U14357 (N_14357,N_7574,N_8695);
and U14358 (N_14358,N_9330,N_5345);
and U14359 (N_14359,N_6595,N_8629);
xor U14360 (N_14360,N_7898,N_6766);
and U14361 (N_14361,N_6325,N_6640);
xnor U14362 (N_14362,N_8886,N_5032);
xor U14363 (N_14363,N_6731,N_5656);
xnor U14364 (N_14364,N_6550,N_5296);
or U14365 (N_14365,N_9149,N_9516);
nor U14366 (N_14366,N_5275,N_7657);
nor U14367 (N_14367,N_8636,N_6911);
and U14368 (N_14368,N_8714,N_9602);
xor U14369 (N_14369,N_6592,N_8514);
or U14370 (N_14370,N_5054,N_5023);
nor U14371 (N_14371,N_8463,N_9294);
and U14372 (N_14372,N_6636,N_6599);
and U14373 (N_14373,N_7863,N_6275);
xnor U14374 (N_14374,N_6634,N_9536);
nand U14375 (N_14375,N_6907,N_7199);
xnor U14376 (N_14376,N_8408,N_9202);
xnor U14377 (N_14377,N_9604,N_7604);
nor U14378 (N_14378,N_5472,N_7223);
or U14379 (N_14379,N_7065,N_7710);
nand U14380 (N_14380,N_9693,N_6369);
nand U14381 (N_14381,N_7123,N_8119);
nand U14382 (N_14382,N_7922,N_6013);
nand U14383 (N_14383,N_6859,N_7843);
or U14384 (N_14384,N_7412,N_5099);
nor U14385 (N_14385,N_6012,N_5560);
or U14386 (N_14386,N_9064,N_7877);
nand U14387 (N_14387,N_8816,N_7522);
or U14388 (N_14388,N_8660,N_5271);
or U14389 (N_14389,N_8699,N_9229);
and U14390 (N_14390,N_6636,N_8223);
and U14391 (N_14391,N_8889,N_7375);
xnor U14392 (N_14392,N_8390,N_8743);
and U14393 (N_14393,N_5471,N_5861);
or U14394 (N_14394,N_7673,N_6288);
nor U14395 (N_14395,N_6687,N_9816);
nor U14396 (N_14396,N_6771,N_9243);
nor U14397 (N_14397,N_6756,N_9592);
and U14398 (N_14398,N_8169,N_9290);
and U14399 (N_14399,N_7210,N_9918);
or U14400 (N_14400,N_6576,N_6056);
and U14401 (N_14401,N_5506,N_7798);
or U14402 (N_14402,N_9801,N_9559);
nor U14403 (N_14403,N_8268,N_8026);
xor U14404 (N_14404,N_6062,N_5718);
nor U14405 (N_14405,N_7141,N_5049);
nor U14406 (N_14406,N_5912,N_7563);
and U14407 (N_14407,N_5855,N_5132);
nand U14408 (N_14408,N_8948,N_6835);
nor U14409 (N_14409,N_6560,N_7443);
nor U14410 (N_14410,N_7750,N_5163);
or U14411 (N_14411,N_5861,N_7424);
and U14412 (N_14412,N_8477,N_5725);
xor U14413 (N_14413,N_7822,N_6052);
nor U14414 (N_14414,N_6674,N_8376);
xnor U14415 (N_14415,N_7466,N_7934);
nor U14416 (N_14416,N_7395,N_8464);
nand U14417 (N_14417,N_7419,N_8916);
or U14418 (N_14418,N_6801,N_5942);
or U14419 (N_14419,N_7450,N_7831);
and U14420 (N_14420,N_5303,N_6268);
or U14421 (N_14421,N_8188,N_9094);
xnor U14422 (N_14422,N_5165,N_5646);
or U14423 (N_14423,N_6154,N_9843);
or U14424 (N_14424,N_9979,N_5184);
xnor U14425 (N_14425,N_6836,N_6654);
and U14426 (N_14426,N_6458,N_8450);
and U14427 (N_14427,N_6650,N_8073);
nand U14428 (N_14428,N_9189,N_5801);
and U14429 (N_14429,N_5314,N_9961);
xor U14430 (N_14430,N_5362,N_9670);
and U14431 (N_14431,N_5026,N_7776);
xnor U14432 (N_14432,N_9669,N_7246);
nor U14433 (N_14433,N_6265,N_5283);
nand U14434 (N_14434,N_5151,N_5435);
and U14435 (N_14435,N_5381,N_7942);
or U14436 (N_14436,N_6632,N_5617);
xor U14437 (N_14437,N_6668,N_8339);
nor U14438 (N_14438,N_6208,N_9227);
xnor U14439 (N_14439,N_5433,N_7024);
nand U14440 (N_14440,N_6799,N_8842);
nor U14441 (N_14441,N_7503,N_8777);
nor U14442 (N_14442,N_7356,N_9687);
nor U14443 (N_14443,N_5443,N_8421);
and U14444 (N_14444,N_9227,N_9670);
and U14445 (N_14445,N_9463,N_7867);
xor U14446 (N_14446,N_7198,N_8088);
and U14447 (N_14447,N_8837,N_6472);
and U14448 (N_14448,N_8310,N_8289);
nor U14449 (N_14449,N_7006,N_6615);
nand U14450 (N_14450,N_9513,N_9156);
nand U14451 (N_14451,N_6123,N_5454);
and U14452 (N_14452,N_6756,N_7527);
and U14453 (N_14453,N_5351,N_7590);
and U14454 (N_14454,N_5295,N_9977);
xor U14455 (N_14455,N_9133,N_7974);
or U14456 (N_14456,N_5861,N_9465);
nor U14457 (N_14457,N_7314,N_7652);
and U14458 (N_14458,N_7100,N_8721);
nor U14459 (N_14459,N_8819,N_5739);
nor U14460 (N_14460,N_6635,N_9453);
nand U14461 (N_14461,N_9395,N_5039);
xnor U14462 (N_14462,N_8681,N_6908);
or U14463 (N_14463,N_6706,N_8983);
nor U14464 (N_14464,N_5606,N_5212);
or U14465 (N_14465,N_8090,N_7491);
and U14466 (N_14466,N_5137,N_5340);
nand U14467 (N_14467,N_5596,N_5252);
or U14468 (N_14468,N_9147,N_6460);
xor U14469 (N_14469,N_5760,N_6835);
nand U14470 (N_14470,N_5362,N_5804);
nor U14471 (N_14471,N_7628,N_6509);
xnor U14472 (N_14472,N_9186,N_6866);
or U14473 (N_14473,N_5727,N_5422);
or U14474 (N_14474,N_6292,N_7015);
xnor U14475 (N_14475,N_6689,N_9252);
nor U14476 (N_14476,N_7931,N_7665);
nor U14477 (N_14477,N_9122,N_6194);
nor U14478 (N_14478,N_5946,N_7155);
and U14479 (N_14479,N_7317,N_5467);
xor U14480 (N_14480,N_6709,N_7793);
nand U14481 (N_14481,N_9411,N_7151);
nand U14482 (N_14482,N_5589,N_9508);
and U14483 (N_14483,N_6905,N_7617);
nand U14484 (N_14484,N_7163,N_7448);
or U14485 (N_14485,N_7164,N_6498);
and U14486 (N_14486,N_9152,N_6707);
or U14487 (N_14487,N_6491,N_9910);
nand U14488 (N_14488,N_7888,N_6048);
or U14489 (N_14489,N_9539,N_6387);
nor U14490 (N_14490,N_5107,N_6958);
nand U14491 (N_14491,N_7100,N_7862);
nand U14492 (N_14492,N_8006,N_6092);
and U14493 (N_14493,N_9264,N_8419);
and U14494 (N_14494,N_9091,N_9884);
and U14495 (N_14495,N_8700,N_5504);
and U14496 (N_14496,N_5595,N_5152);
nand U14497 (N_14497,N_6166,N_8191);
xor U14498 (N_14498,N_7558,N_6299);
and U14499 (N_14499,N_6938,N_6073);
xor U14500 (N_14500,N_8236,N_8322);
or U14501 (N_14501,N_5850,N_7654);
nor U14502 (N_14502,N_7834,N_7246);
xor U14503 (N_14503,N_5965,N_7839);
xnor U14504 (N_14504,N_7691,N_7807);
xor U14505 (N_14505,N_6292,N_7056);
and U14506 (N_14506,N_5299,N_6914);
nand U14507 (N_14507,N_9155,N_6200);
nand U14508 (N_14508,N_8879,N_6993);
and U14509 (N_14509,N_5912,N_8988);
nand U14510 (N_14510,N_6440,N_6336);
and U14511 (N_14511,N_5074,N_8439);
or U14512 (N_14512,N_7435,N_6183);
xor U14513 (N_14513,N_7993,N_8796);
and U14514 (N_14514,N_6259,N_5915);
nand U14515 (N_14515,N_6716,N_5541);
nand U14516 (N_14516,N_5327,N_9064);
or U14517 (N_14517,N_8594,N_9914);
or U14518 (N_14518,N_9468,N_5951);
and U14519 (N_14519,N_9737,N_7413);
nor U14520 (N_14520,N_9166,N_7832);
and U14521 (N_14521,N_6795,N_8651);
nor U14522 (N_14522,N_7131,N_9277);
nand U14523 (N_14523,N_6951,N_7227);
and U14524 (N_14524,N_5079,N_9429);
and U14525 (N_14525,N_5195,N_6704);
nor U14526 (N_14526,N_8787,N_9720);
xnor U14527 (N_14527,N_9768,N_5385);
nor U14528 (N_14528,N_5795,N_9704);
xor U14529 (N_14529,N_8963,N_9908);
nand U14530 (N_14530,N_7636,N_5252);
xnor U14531 (N_14531,N_8954,N_7166);
nor U14532 (N_14532,N_9062,N_8435);
and U14533 (N_14533,N_7737,N_6279);
nand U14534 (N_14534,N_8698,N_7753);
or U14535 (N_14535,N_8675,N_7296);
or U14536 (N_14536,N_6410,N_9740);
nand U14537 (N_14537,N_7448,N_6299);
nor U14538 (N_14538,N_7680,N_6378);
nor U14539 (N_14539,N_8921,N_5797);
nor U14540 (N_14540,N_5804,N_9533);
nand U14541 (N_14541,N_9983,N_5745);
or U14542 (N_14542,N_5214,N_7304);
nand U14543 (N_14543,N_5172,N_5596);
nand U14544 (N_14544,N_8954,N_6908);
nand U14545 (N_14545,N_7949,N_7479);
nand U14546 (N_14546,N_5499,N_8894);
and U14547 (N_14547,N_6639,N_5782);
and U14548 (N_14548,N_7230,N_7293);
or U14549 (N_14549,N_9069,N_7588);
nor U14550 (N_14550,N_5328,N_7780);
nand U14551 (N_14551,N_9055,N_5211);
nand U14552 (N_14552,N_9491,N_5969);
xnor U14553 (N_14553,N_7057,N_5273);
xor U14554 (N_14554,N_6012,N_6544);
nand U14555 (N_14555,N_6620,N_9311);
nor U14556 (N_14556,N_9545,N_9265);
xnor U14557 (N_14557,N_8620,N_9783);
nor U14558 (N_14558,N_7861,N_7526);
and U14559 (N_14559,N_8163,N_5215);
nor U14560 (N_14560,N_6971,N_8014);
nor U14561 (N_14561,N_9598,N_6706);
or U14562 (N_14562,N_7235,N_7849);
or U14563 (N_14563,N_5231,N_6041);
nor U14564 (N_14564,N_6349,N_9568);
nand U14565 (N_14565,N_7974,N_6225);
nand U14566 (N_14566,N_8401,N_5463);
xnor U14567 (N_14567,N_8848,N_9915);
and U14568 (N_14568,N_9717,N_8196);
or U14569 (N_14569,N_7642,N_6037);
or U14570 (N_14570,N_8454,N_8778);
nand U14571 (N_14571,N_6545,N_7959);
or U14572 (N_14572,N_5351,N_9783);
xnor U14573 (N_14573,N_6130,N_5262);
or U14574 (N_14574,N_8916,N_5233);
and U14575 (N_14575,N_6957,N_9611);
and U14576 (N_14576,N_5531,N_5235);
or U14577 (N_14577,N_7315,N_7842);
nand U14578 (N_14578,N_8309,N_8620);
nor U14579 (N_14579,N_7212,N_5531);
or U14580 (N_14580,N_8496,N_9326);
or U14581 (N_14581,N_6162,N_7125);
and U14582 (N_14582,N_7321,N_5680);
nand U14583 (N_14583,N_8470,N_7372);
xnor U14584 (N_14584,N_9517,N_5920);
nor U14585 (N_14585,N_5015,N_7253);
nor U14586 (N_14586,N_6468,N_8695);
xor U14587 (N_14587,N_5471,N_7833);
xnor U14588 (N_14588,N_7484,N_5073);
xor U14589 (N_14589,N_5574,N_6303);
nor U14590 (N_14590,N_9574,N_5526);
xor U14591 (N_14591,N_7500,N_9401);
or U14592 (N_14592,N_8426,N_6669);
nand U14593 (N_14593,N_9532,N_6457);
or U14594 (N_14594,N_8203,N_5013);
nand U14595 (N_14595,N_5295,N_6222);
nand U14596 (N_14596,N_8084,N_5472);
and U14597 (N_14597,N_6086,N_8992);
nand U14598 (N_14598,N_7164,N_8881);
xor U14599 (N_14599,N_5532,N_6577);
xnor U14600 (N_14600,N_7819,N_7585);
and U14601 (N_14601,N_8234,N_6489);
nor U14602 (N_14602,N_6588,N_8777);
xnor U14603 (N_14603,N_9841,N_6170);
xor U14604 (N_14604,N_5390,N_8004);
nand U14605 (N_14605,N_8167,N_5265);
and U14606 (N_14606,N_5080,N_8128);
or U14607 (N_14607,N_8174,N_7576);
and U14608 (N_14608,N_8518,N_8456);
nand U14609 (N_14609,N_9630,N_6874);
xnor U14610 (N_14610,N_8148,N_9996);
nand U14611 (N_14611,N_7892,N_5718);
xor U14612 (N_14612,N_9378,N_8708);
nand U14613 (N_14613,N_7192,N_7403);
xor U14614 (N_14614,N_9713,N_6220);
and U14615 (N_14615,N_9941,N_6754);
or U14616 (N_14616,N_6150,N_9412);
and U14617 (N_14617,N_8455,N_8888);
nand U14618 (N_14618,N_5539,N_5273);
or U14619 (N_14619,N_6302,N_9959);
nor U14620 (N_14620,N_6020,N_9497);
xnor U14621 (N_14621,N_8462,N_7122);
and U14622 (N_14622,N_7445,N_9781);
nand U14623 (N_14623,N_8539,N_5154);
nand U14624 (N_14624,N_8749,N_5707);
xor U14625 (N_14625,N_5462,N_9781);
nand U14626 (N_14626,N_8280,N_9932);
and U14627 (N_14627,N_6432,N_6280);
and U14628 (N_14628,N_5525,N_6657);
nand U14629 (N_14629,N_6678,N_5166);
nor U14630 (N_14630,N_6895,N_7889);
and U14631 (N_14631,N_8840,N_8634);
nor U14632 (N_14632,N_7046,N_9308);
and U14633 (N_14633,N_6959,N_9996);
nor U14634 (N_14634,N_8108,N_5208);
and U14635 (N_14635,N_6233,N_7906);
xnor U14636 (N_14636,N_7021,N_7029);
nand U14637 (N_14637,N_6471,N_9202);
or U14638 (N_14638,N_5832,N_9203);
xnor U14639 (N_14639,N_6518,N_6180);
or U14640 (N_14640,N_6530,N_7269);
nand U14641 (N_14641,N_5656,N_8953);
xor U14642 (N_14642,N_7685,N_6417);
or U14643 (N_14643,N_5686,N_7274);
nand U14644 (N_14644,N_7175,N_9824);
xor U14645 (N_14645,N_9059,N_7081);
and U14646 (N_14646,N_6002,N_6554);
or U14647 (N_14647,N_7227,N_6101);
nand U14648 (N_14648,N_7908,N_8183);
and U14649 (N_14649,N_8454,N_6289);
nor U14650 (N_14650,N_8780,N_5253);
nand U14651 (N_14651,N_5525,N_5283);
nor U14652 (N_14652,N_8528,N_9101);
nand U14653 (N_14653,N_9083,N_7715);
nor U14654 (N_14654,N_8932,N_7359);
nor U14655 (N_14655,N_5020,N_7185);
or U14656 (N_14656,N_6422,N_8563);
or U14657 (N_14657,N_9414,N_9090);
xnor U14658 (N_14658,N_5565,N_5352);
nor U14659 (N_14659,N_9744,N_6223);
nand U14660 (N_14660,N_6089,N_5219);
nand U14661 (N_14661,N_7654,N_8536);
nand U14662 (N_14662,N_7508,N_9316);
or U14663 (N_14663,N_6302,N_6732);
or U14664 (N_14664,N_5707,N_6384);
nor U14665 (N_14665,N_7158,N_6617);
xor U14666 (N_14666,N_6734,N_5020);
and U14667 (N_14667,N_7016,N_5121);
xor U14668 (N_14668,N_5658,N_8483);
and U14669 (N_14669,N_6866,N_7214);
or U14670 (N_14670,N_5654,N_9289);
nor U14671 (N_14671,N_8163,N_7961);
nor U14672 (N_14672,N_6793,N_6651);
nand U14673 (N_14673,N_8856,N_6069);
nor U14674 (N_14674,N_6837,N_8819);
nand U14675 (N_14675,N_7908,N_8965);
nor U14676 (N_14676,N_9618,N_6397);
or U14677 (N_14677,N_5063,N_9536);
nand U14678 (N_14678,N_7139,N_7985);
and U14679 (N_14679,N_7379,N_7925);
xor U14680 (N_14680,N_5565,N_9100);
nor U14681 (N_14681,N_8056,N_9172);
nor U14682 (N_14682,N_7795,N_7146);
or U14683 (N_14683,N_9389,N_9353);
nand U14684 (N_14684,N_7188,N_6158);
nor U14685 (N_14685,N_7644,N_9681);
nand U14686 (N_14686,N_7548,N_7389);
xnor U14687 (N_14687,N_5555,N_5575);
nor U14688 (N_14688,N_6367,N_8142);
nand U14689 (N_14689,N_7439,N_8437);
and U14690 (N_14690,N_6328,N_6450);
xnor U14691 (N_14691,N_8416,N_8366);
nor U14692 (N_14692,N_6057,N_9678);
xor U14693 (N_14693,N_8637,N_9057);
nand U14694 (N_14694,N_9463,N_5428);
xor U14695 (N_14695,N_9694,N_9624);
nor U14696 (N_14696,N_8916,N_7713);
nor U14697 (N_14697,N_9928,N_8114);
or U14698 (N_14698,N_6230,N_6338);
nor U14699 (N_14699,N_9920,N_5403);
xor U14700 (N_14700,N_5361,N_8721);
xor U14701 (N_14701,N_6113,N_9847);
and U14702 (N_14702,N_6511,N_8905);
nand U14703 (N_14703,N_6270,N_7083);
xor U14704 (N_14704,N_8972,N_8425);
or U14705 (N_14705,N_7345,N_5721);
and U14706 (N_14706,N_5481,N_9098);
nor U14707 (N_14707,N_5935,N_8538);
and U14708 (N_14708,N_9643,N_5076);
or U14709 (N_14709,N_6913,N_6650);
nor U14710 (N_14710,N_6640,N_5548);
or U14711 (N_14711,N_5056,N_9542);
nor U14712 (N_14712,N_8397,N_6548);
nand U14713 (N_14713,N_9763,N_6621);
or U14714 (N_14714,N_7373,N_8563);
or U14715 (N_14715,N_7112,N_9901);
xnor U14716 (N_14716,N_5048,N_8387);
nor U14717 (N_14717,N_6863,N_8444);
xor U14718 (N_14718,N_8181,N_8221);
or U14719 (N_14719,N_5080,N_7624);
nand U14720 (N_14720,N_8697,N_6275);
nand U14721 (N_14721,N_9384,N_8290);
nor U14722 (N_14722,N_7063,N_5026);
and U14723 (N_14723,N_9006,N_6242);
xnor U14724 (N_14724,N_7323,N_8623);
xnor U14725 (N_14725,N_6196,N_9787);
and U14726 (N_14726,N_7404,N_5668);
and U14727 (N_14727,N_6428,N_5730);
or U14728 (N_14728,N_5489,N_7917);
xnor U14729 (N_14729,N_6242,N_6534);
xnor U14730 (N_14730,N_6894,N_8408);
and U14731 (N_14731,N_6172,N_7660);
nor U14732 (N_14732,N_9504,N_9327);
nor U14733 (N_14733,N_7832,N_9543);
xnor U14734 (N_14734,N_8301,N_7206);
nand U14735 (N_14735,N_9163,N_7831);
and U14736 (N_14736,N_9731,N_6148);
or U14737 (N_14737,N_8494,N_6427);
xor U14738 (N_14738,N_9453,N_5238);
nor U14739 (N_14739,N_8259,N_8222);
xnor U14740 (N_14740,N_7426,N_9538);
and U14741 (N_14741,N_9827,N_7475);
or U14742 (N_14742,N_9452,N_5884);
nor U14743 (N_14743,N_8268,N_8173);
and U14744 (N_14744,N_6350,N_9048);
or U14745 (N_14745,N_7345,N_8207);
xor U14746 (N_14746,N_5787,N_7888);
and U14747 (N_14747,N_5136,N_7351);
xnor U14748 (N_14748,N_7206,N_9238);
nor U14749 (N_14749,N_9763,N_8210);
nor U14750 (N_14750,N_6294,N_9063);
nand U14751 (N_14751,N_8699,N_7565);
nand U14752 (N_14752,N_8551,N_8840);
nor U14753 (N_14753,N_7743,N_8375);
and U14754 (N_14754,N_9053,N_7862);
nand U14755 (N_14755,N_5877,N_9765);
and U14756 (N_14756,N_9206,N_7739);
nand U14757 (N_14757,N_9752,N_9674);
nand U14758 (N_14758,N_8373,N_8196);
nor U14759 (N_14759,N_7604,N_5553);
and U14760 (N_14760,N_5911,N_8827);
xnor U14761 (N_14761,N_7465,N_7343);
and U14762 (N_14762,N_7025,N_5399);
xnor U14763 (N_14763,N_6541,N_7024);
nand U14764 (N_14764,N_6250,N_9787);
or U14765 (N_14765,N_7839,N_8132);
nand U14766 (N_14766,N_6891,N_9305);
nand U14767 (N_14767,N_5959,N_9086);
nand U14768 (N_14768,N_6193,N_6620);
nor U14769 (N_14769,N_6553,N_5752);
nand U14770 (N_14770,N_9867,N_7423);
xnor U14771 (N_14771,N_9449,N_8786);
nor U14772 (N_14772,N_8738,N_7626);
xnor U14773 (N_14773,N_8005,N_5668);
nor U14774 (N_14774,N_7064,N_8954);
and U14775 (N_14775,N_7670,N_6718);
nand U14776 (N_14776,N_7465,N_7155);
nor U14777 (N_14777,N_6708,N_7173);
xnor U14778 (N_14778,N_6517,N_5126);
or U14779 (N_14779,N_5629,N_9745);
xor U14780 (N_14780,N_8679,N_5041);
and U14781 (N_14781,N_8542,N_5693);
and U14782 (N_14782,N_8739,N_8106);
or U14783 (N_14783,N_5755,N_9464);
or U14784 (N_14784,N_6697,N_6420);
nand U14785 (N_14785,N_6564,N_8477);
and U14786 (N_14786,N_6755,N_9474);
xor U14787 (N_14787,N_7289,N_9090);
nor U14788 (N_14788,N_8314,N_8676);
nand U14789 (N_14789,N_7591,N_8751);
nor U14790 (N_14790,N_7739,N_6135);
xnor U14791 (N_14791,N_7989,N_9296);
xor U14792 (N_14792,N_9909,N_8923);
nor U14793 (N_14793,N_9723,N_6772);
and U14794 (N_14794,N_8752,N_6364);
or U14795 (N_14795,N_6230,N_7751);
or U14796 (N_14796,N_8225,N_6277);
nor U14797 (N_14797,N_6632,N_5140);
and U14798 (N_14798,N_9400,N_5083);
and U14799 (N_14799,N_7105,N_9263);
nor U14800 (N_14800,N_5516,N_7280);
or U14801 (N_14801,N_5510,N_8952);
nor U14802 (N_14802,N_8964,N_7244);
nor U14803 (N_14803,N_9227,N_5351);
nand U14804 (N_14804,N_7133,N_9426);
nand U14805 (N_14805,N_6102,N_8610);
nand U14806 (N_14806,N_5821,N_7729);
xnor U14807 (N_14807,N_6102,N_5430);
xnor U14808 (N_14808,N_7929,N_7652);
or U14809 (N_14809,N_8868,N_7132);
and U14810 (N_14810,N_8505,N_6395);
nand U14811 (N_14811,N_7216,N_7320);
nand U14812 (N_14812,N_8856,N_5089);
or U14813 (N_14813,N_7980,N_6561);
and U14814 (N_14814,N_9239,N_9754);
nand U14815 (N_14815,N_8017,N_7449);
or U14816 (N_14816,N_9590,N_9515);
xor U14817 (N_14817,N_9576,N_8552);
nand U14818 (N_14818,N_8824,N_8532);
or U14819 (N_14819,N_5054,N_7180);
xor U14820 (N_14820,N_5270,N_8193);
xor U14821 (N_14821,N_9524,N_7356);
nor U14822 (N_14822,N_9524,N_6910);
nand U14823 (N_14823,N_7885,N_8040);
nor U14824 (N_14824,N_7373,N_9195);
nor U14825 (N_14825,N_6033,N_5769);
or U14826 (N_14826,N_8046,N_6247);
nand U14827 (N_14827,N_7360,N_7228);
and U14828 (N_14828,N_5337,N_5252);
or U14829 (N_14829,N_8721,N_7256);
and U14830 (N_14830,N_5442,N_5716);
xnor U14831 (N_14831,N_8255,N_7844);
or U14832 (N_14832,N_5591,N_9461);
nand U14833 (N_14833,N_9832,N_6298);
xnor U14834 (N_14834,N_8519,N_5856);
or U14835 (N_14835,N_5288,N_7910);
nand U14836 (N_14836,N_6016,N_8168);
or U14837 (N_14837,N_8646,N_8224);
and U14838 (N_14838,N_7086,N_6077);
and U14839 (N_14839,N_9597,N_7900);
nand U14840 (N_14840,N_7546,N_6692);
nand U14841 (N_14841,N_7963,N_7666);
or U14842 (N_14842,N_5244,N_8830);
or U14843 (N_14843,N_9774,N_5605);
xor U14844 (N_14844,N_8998,N_6736);
and U14845 (N_14845,N_8068,N_7330);
or U14846 (N_14846,N_9204,N_7252);
or U14847 (N_14847,N_8552,N_5070);
xnor U14848 (N_14848,N_5962,N_6056);
and U14849 (N_14849,N_8316,N_9684);
nor U14850 (N_14850,N_5237,N_5762);
xor U14851 (N_14851,N_9506,N_8655);
xnor U14852 (N_14852,N_7784,N_7528);
or U14853 (N_14853,N_8995,N_7547);
xnor U14854 (N_14854,N_8652,N_8445);
xor U14855 (N_14855,N_7935,N_6413);
and U14856 (N_14856,N_8305,N_5965);
xnor U14857 (N_14857,N_7539,N_6257);
or U14858 (N_14858,N_6933,N_6445);
nand U14859 (N_14859,N_7406,N_5058);
and U14860 (N_14860,N_5293,N_6783);
xnor U14861 (N_14861,N_9718,N_7971);
nor U14862 (N_14862,N_5104,N_6766);
or U14863 (N_14863,N_6606,N_7136);
or U14864 (N_14864,N_9186,N_7927);
nand U14865 (N_14865,N_9384,N_8712);
nor U14866 (N_14866,N_5127,N_7308);
nand U14867 (N_14867,N_8484,N_8521);
or U14868 (N_14868,N_5567,N_7429);
nand U14869 (N_14869,N_7136,N_7800);
nand U14870 (N_14870,N_7751,N_7217);
xor U14871 (N_14871,N_6895,N_6789);
nand U14872 (N_14872,N_9930,N_5878);
or U14873 (N_14873,N_9276,N_9923);
xnor U14874 (N_14874,N_7159,N_8909);
nor U14875 (N_14875,N_7716,N_5530);
nand U14876 (N_14876,N_9746,N_5866);
nand U14877 (N_14877,N_8599,N_5074);
nand U14878 (N_14878,N_9142,N_8477);
nor U14879 (N_14879,N_9837,N_7784);
xnor U14880 (N_14880,N_7646,N_6920);
nor U14881 (N_14881,N_7048,N_9057);
nand U14882 (N_14882,N_5801,N_8382);
nor U14883 (N_14883,N_5846,N_7724);
or U14884 (N_14884,N_8296,N_9148);
and U14885 (N_14885,N_7666,N_9946);
xor U14886 (N_14886,N_7160,N_5206);
or U14887 (N_14887,N_5415,N_8504);
or U14888 (N_14888,N_7846,N_8761);
nand U14889 (N_14889,N_6494,N_6557);
nor U14890 (N_14890,N_8183,N_9359);
and U14891 (N_14891,N_5201,N_7371);
nor U14892 (N_14892,N_7371,N_9235);
or U14893 (N_14893,N_5960,N_6769);
nand U14894 (N_14894,N_7410,N_8440);
nor U14895 (N_14895,N_6838,N_9076);
nor U14896 (N_14896,N_6231,N_8567);
and U14897 (N_14897,N_6100,N_6479);
xor U14898 (N_14898,N_8544,N_8580);
nand U14899 (N_14899,N_5141,N_5195);
or U14900 (N_14900,N_5219,N_9046);
or U14901 (N_14901,N_7305,N_7333);
nor U14902 (N_14902,N_8735,N_6760);
nor U14903 (N_14903,N_9065,N_9990);
nor U14904 (N_14904,N_5651,N_9579);
or U14905 (N_14905,N_8751,N_6743);
and U14906 (N_14906,N_7873,N_9157);
xor U14907 (N_14907,N_8177,N_9685);
xor U14908 (N_14908,N_7434,N_9154);
xnor U14909 (N_14909,N_9044,N_9026);
and U14910 (N_14910,N_8157,N_9827);
xnor U14911 (N_14911,N_8719,N_5911);
nor U14912 (N_14912,N_8317,N_9377);
or U14913 (N_14913,N_5434,N_5849);
xor U14914 (N_14914,N_7229,N_7926);
and U14915 (N_14915,N_6295,N_8350);
and U14916 (N_14916,N_8377,N_6664);
or U14917 (N_14917,N_5075,N_6931);
and U14918 (N_14918,N_6438,N_8968);
nor U14919 (N_14919,N_5229,N_7984);
nor U14920 (N_14920,N_5207,N_9920);
or U14921 (N_14921,N_5069,N_9758);
and U14922 (N_14922,N_7496,N_7730);
and U14923 (N_14923,N_6253,N_6374);
and U14924 (N_14924,N_6016,N_6391);
and U14925 (N_14925,N_7880,N_8445);
nand U14926 (N_14926,N_8230,N_5007);
xnor U14927 (N_14927,N_7159,N_6091);
or U14928 (N_14928,N_7348,N_6708);
and U14929 (N_14929,N_6438,N_8199);
and U14930 (N_14930,N_7419,N_5459);
xnor U14931 (N_14931,N_7878,N_9143);
nand U14932 (N_14932,N_6816,N_6795);
or U14933 (N_14933,N_9743,N_9290);
xor U14934 (N_14934,N_6812,N_7243);
nor U14935 (N_14935,N_9420,N_8941);
xor U14936 (N_14936,N_9924,N_5362);
nor U14937 (N_14937,N_5189,N_7738);
xor U14938 (N_14938,N_8723,N_9777);
nor U14939 (N_14939,N_7901,N_5214);
or U14940 (N_14940,N_6512,N_5514);
or U14941 (N_14941,N_7415,N_9194);
or U14942 (N_14942,N_9886,N_9363);
nor U14943 (N_14943,N_8509,N_5481);
xnor U14944 (N_14944,N_6378,N_5699);
or U14945 (N_14945,N_7678,N_6288);
nand U14946 (N_14946,N_8749,N_8618);
and U14947 (N_14947,N_7793,N_9016);
or U14948 (N_14948,N_9359,N_7055);
nand U14949 (N_14949,N_8042,N_5734);
xor U14950 (N_14950,N_7629,N_6897);
xnor U14951 (N_14951,N_5919,N_5020);
or U14952 (N_14952,N_6839,N_6214);
and U14953 (N_14953,N_5632,N_7999);
xnor U14954 (N_14954,N_9559,N_5408);
and U14955 (N_14955,N_5727,N_9923);
and U14956 (N_14956,N_9501,N_6580);
xnor U14957 (N_14957,N_6747,N_5529);
nand U14958 (N_14958,N_7969,N_7821);
or U14959 (N_14959,N_9531,N_6628);
xnor U14960 (N_14960,N_8259,N_7239);
xnor U14961 (N_14961,N_9370,N_7268);
or U14962 (N_14962,N_6226,N_8214);
xor U14963 (N_14963,N_7639,N_8139);
and U14964 (N_14964,N_8080,N_6053);
or U14965 (N_14965,N_7198,N_9809);
nand U14966 (N_14966,N_8073,N_8864);
nand U14967 (N_14967,N_6642,N_8220);
nand U14968 (N_14968,N_8868,N_5410);
nor U14969 (N_14969,N_5865,N_5792);
and U14970 (N_14970,N_5613,N_9331);
xor U14971 (N_14971,N_6163,N_6840);
or U14972 (N_14972,N_5645,N_9438);
nor U14973 (N_14973,N_8735,N_5273);
and U14974 (N_14974,N_8791,N_7921);
and U14975 (N_14975,N_7921,N_5280);
and U14976 (N_14976,N_5347,N_5688);
nor U14977 (N_14977,N_8017,N_7211);
nand U14978 (N_14978,N_7524,N_8773);
nor U14979 (N_14979,N_5630,N_9823);
nand U14980 (N_14980,N_9189,N_9648);
nor U14981 (N_14981,N_7262,N_5318);
xor U14982 (N_14982,N_6148,N_7108);
xnor U14983 (N_14983,N_9625,N_6683);
xor U14984 (N_14984,N_8835,N_8176);
or U14985 (N_14985,N_5217,N_5573);
nor U14986 (N_14986,N_6694,N_8582);
and U14987 (N_14987,N_5759,N_5905);
and U14988 (N_14988,N_7030,N_7881);
and U14989 (N_14989,N_8393,N_6787);
or U14990 (N_14990,N_6802,N_6180);
nand U14991 (N_14991,N_7781,N_9958);
nand U14992 (N_14992,N_8537,N_9541);
or U14993 (N_14993,N_7750,N_5147);
nor U14994 (N_14994,N_5345,N_9511);
nand U14995 (N_14995,N_6194,N_5625);
nand U14996 (N_14996,N_7895,N_7172);
or U14997 (N_14997,N_5092,N_6363);
and U14998 (N_14998,N_9186,N_9571);
nand U14999 (N_14999,N_8529,N_7668);
nand U15000 (N_15000,N_12375,N_12537);
xor U15001 (N_15001,N_12414,N_13056);
and U15002 (N_15002,N_14741,N_11624);
nand U15003 (N_15003,N_12271,N_12387);
nor U15004 (N_15004,N_12397,N_13214);
or U15005 (N_15005,N_10154,N_10688);
nand U15006 (N_15006,N_13844,N_14394);
and U15007 (N_15007,N_14171,N_13209);
or U15008 (N_15008,N_10027,N_13494);
and U15009 (N_15009,N_10560,N_11321);
and U15010 (N_15010,N_12383,N_14249);
or U15011 (N_15011,N_13632,N_12662);
xor U15012 (N_15012,N_14871,N_11623);
nand U15013 (N_15013,N_10801,N_13597);
nand U15014 (N_15014,N_13359,N_12869);
nor U15015 (N_15015,N_11074,N_10327);
nor U15016 (N_15016,N_14144,N_11785);
xor U15017 (N_15017,N_11763,N_10996);
nand U15018 (N_15018,N_11508,N_13477);
and U15019 (N_15019,N_12098,N_12436);
xnor U15020 (N_15020,N_11073,N_14983);
xnor U15021 (N_15021,N_12756,N_11903);
and U15022 (N_15022,N_11323,N_11496);
nor U15023 (N_15023,N_13231,N_13652);
nor U15024 (N_15024,N_10828,N_10180);
nor U15025 (N_15025,N_10293,N_11909);
and U15026 (N_15026,N_12648,N_11856);
nand U15027 (N_15027,N_13598,N_10537);
nand U15028 (N_15028,N_13470,N_13460);
nor U15029 (N_15029,N_13305,N_12054);
or U15030 (N_15030,N_11382,N_10173);
xor U15031 (N_15031,N_11373,N_13116);
nor U15032 (N_15032,N_13979,N_14486);
or U15033 (N_15033,N_11503,N_12325);
or U15034 (N_15034,N_11448,N_14867);
nor U15035 (N_15035,N_11228,N_12020);
and U15036 (N_15036,N_10695,N_10418);
nand U15037 (N_15037,N_13747,N_10858);
xor U15038 (N_15038,N_11134,N_11020);
or U15039 (N_15039,N_12295,N_10124);
nor U15040 (N_15040,N_12453,N_13081);
xor U15041 (N_15041,N_10726,N_14930);
xnor U15042 (N_15042,N_11002,N_10047);
and U15043 (N_15043,N_14580,N_10482);
nand U15044 (N_15044,N_14328,N_14095);
nor U15045 (N_15045,N_13294,N_14522);
nor U15046 (N_15046,N_14287,N_12493);
xnor U15047 (N_15047,N_13548,N_10244);
or U15048 (N_15048,N_14788,N_12310);
xnor U15049 (N_15049,N_12723,N_11702);
or U15050 (N_15050,N_13031,N_14977);
xor U15051 (N_15051,N_10110,N_14664);
nand U15052 (N_15052,N_13828,N_12289);
or U15053 (N_15053,N_11263,N_11286);
nor U15054 (N_15054,N_14431,N_14904);
and U15055 (N_15055,N_14107,N_11842);
nand U15056 (N_15056,N_13017,N_14634);
nor U15057 (N_15057,N_13790,N_10582);
xor U15058 (N_15058,N_13211,N_12277);
or U15059 (N_15059,N_12423,N_12591);
or U15060 (N_15060,N_13076,N_10501);
nand U15061 (N_15061,N_14742,N_10126);
nand U15062 (N_15062,N_14678,N_10837);
nor U15063 (N_15063,N_14417,N_14818);
or U15064 (N_15064,N_10646,N_14419);
and U15065 (N_15065,N_13707,N_12055);
nor U15066 (N_15066,N_11684,N_10343);
nor U15067 (N_15067,N_14336,N_10937);
and U15068 (N_15068,N_12534,N_10385);
and U15069 (N_15069,N_12180,N_11621);
and U15070 (N_15070,N_11556,N_11719);
nand U15071 (N_15071,N_12092,N_11867);
or U15072 (N_15072,N_13126,N_13408);
nor U15073 (N_15073,N_12175,N_12068);
nor U15074 (N_15074,N_10079,N_13662);
and U15075 (N_15075,N_10383,N_12316);
and U15076 (N_15076,N_11056,N_11462);
or U15077 (N_15077,N_14143,N_14497);
nor U15078 (N_15078,N_10734,N_13190);
and U15079 (N_15079,N_11067,N_12240);
or U15080 (N_15080,N_10861,N_11232);
nand U15081 (N_15081,N_10532,N_11054);
xor U15082 (N_15082,N_14375,N_11670);
nand U15083 (N_15083,N_11326,N_10622);
or U15084 (N_15084,N_10497,N_12206);
and U15085 (N_15085,N_14811,N_13400);
xor U15086 (N_15086,N_14412,N_13133);
nor U15087 (N_15087,N_10502,N_11590);
nor U15088 (N_15088,N_14384,N_13634);
xnor U15089 (N_15089,N_11728,N_10149);
xor U15090 (N_15090,N_11827,N_10849);
nor U15091 (N_15091,N_13881,N_10403);
nand U15092 (N_15092,N_12368,N_14797);
xnor U15093 (N_15093,N_13394,N_14764);
and U15094 (N_15094,N_10061,N_10478);
or U15095 (N_15095,N_10146,N_13735);
and U15096 (N_15096,N_12774,N_14714);
nor U15097 (N_15097,N_14146,N_12053);
nor U15098 (N_15098,N_14573,N_10966);
nand U15099 (N_15099,N_12629,N_10670);
nor U15100 (N_15100,N_11769,N_11596);
xnor U15101 (N_15101,N_14832,N_10657);
xor U15102 (N_15102,N_13462,N_10183);
and U15103 (N_15103,N_10971,N_11970);
or U15104 (N_15104,N_14790,N_10404);
and U15105 (N_15105,N_10323,N_10813);
nor U15106 (N_15106,N_10266,N_14594);
xor U15107 (N_15107,N_12740,N_12279);
nand U15108 (N_15108,N_14033,N_14680);
nor U15109 (N_15109,N_10766,N_11519);
nand U15110 (N_15110,N_11172,N_14861);
or U15111 (N_15111,N_10460,N_14553);
nor U15112 (N_15112,N_14032,N_10083);
or U15113 (N_15113,N_14214,N_13086);
xnor U15114 (N_15114,N_11136,N_13576);
and U15115 (N_15115,N_10211,N_14174);
or U15116 (N_15116,N_12655,N_11145);
or U15117 (N_15117,N_10210,N_10239);
or U15118 (N_15118,N_11929,N_10200);
or U15119 (N_15119,N_12589,N_13677);
nor U15120 (N_15120,N_14109,N_14383);
xor U15121 (N_15121,N_13474,N_14135);
or U15122 (N_15122,N_14975,N_12699);
nand U15123 (N_15123,N_10246,N_11546);
nor U15124 (N_15124,N_10227,N_10958);
nor U15125 (N_15125,N_10367,N_10171);
nor U15126 (N_15126,N_12808,N_10155);
xor U15127 (N_15127,N_10267,N_11413);
nand U15128 (N_15128,N_12272,N_14645);
and U15129 (N_15129,N_14476,N_12964);
nor U15130 (N_15130,N_13299,N_14963);
and U15131 (N_15131,N_10402,N_11425);
nand U15132 (N_15132,N_12799,N_14087);
xor U15133 (N_15133,N_13645,N_13401);
nand U15134 (N_15134,N_12566,N_13393);
xor U15135 (N_15135,N_13637,N_11376);
nor U15136 (N_15136,N_11848,N_13430);
and U15137 (N_15137,N_11191,N_11348);
and U15138 (N_15138,N_14882,N_12709);
nand U15139 (N_15139,N_10922,N_12601);
xor U15140 (N_15140,N_12538,N_13475);
xnor U15141 (N_15141,N_12299,N_12812);
and U15142 (N_15142,N_12760,N_12646);
nor U15143 (N_15143,N_10477,N_13314);
or U15144 (N_15144,N_14863,N_13850);
nand U15145 (N_15145,N_13010,N_10811);
and U15146 (N_15146,N_13951,N_14083);
nand U15147 (N_15147,N_12650,N_12425);
xor U15148 (N_15148,N_11154,N_11133);
or U15149 (N_15149,N_10053,N_14381);
or U15150 (N_15150,N_14006,N_11488);
nand U15151 (N_15151,N_12035,N_10365);
xnor U15152 (N_15152,N_10559,N_13628);
or U15153 (N_15153,N_12486,N_12926);
xnor U15154 (N_15154,N_12849,N_12746);
nor U15155 (N_15155,N_13286,N_11241);
and U15156 (N_15156,N_12111,N_12074);
xnor U15157 (N_15157,N_11226,N_10744);
and U15158 (N_15158,N_14539,N_12977);
xor U15159 (N_15159,N_14926,N_10091);
nand U15160 (N_15160,N_14357,N_12136);
or U15161 (N_15161,N_12701,N_11548);
nand U15162 (N_15162,N_10767,N_11040);
nand U15163 (N_15163,N_12750,N_13627);
or U15164 (N_15164,N_12044,N_13738);
xnor U15165 (N_15165,N_11042,N_13817);
nand U15166 (N_15166,N_10702,N_14869);
or U15167 (N_15167,N_13841,N_13437);
xnor U15168 (N_15168,N_10097,N_12941);
nand U15169 (N_15169,N_13660,N_13778);
or U15170 (N_15170,N_12007,N_12541);
and U15171 (N_15171,N_14778,N_13102);
nand U15172 (N_15172,N_12787,N_13216);
or U15173 (N_15173,N_11721,N_10757);
or U15174 (N_15174,N_11212,N_14886);
or U15175 (N_15175,N_10997,N_12003);
nand U15176 (N_15176,N_12531,N_14212);
or U15177 (N_15177,N_12927,N_10212);
nand U15178 (N_15178,N_12885,N_13283);
nor U15179 (N_15179,N_12820,N_10369);
and U15180 (N_15180,N_14331,N_11317);
and U15181 (N_15181,N_13878,N_14880);
and U15182 (N_15182,N_13343,N_11638);
and U15183 (N_15183,N_14663,N_14755);
or U15184 (N_15184,N_11540,N_14183);
nand U15185 (N_15185,N_12796,N_11277);
or U15186 (N_15186,N_10269,N_14531);
nor U15187 (N_15187,N_12004,N_10534);
nand U15188 (N_15188,N_13332,N_14614);
and U15189 (N_15189,N_13171,N_13119);
and U15190 (N_15190,N_11731,N_10204);
nor U15191 (N_15191,N_10144,N_13834);
nand U15192 (N_15192,N_10678,N_11756);
or U15193 (N_15193,N_12382,N_10468);
nor U15194 (N_15194,N_10209,N_14814);
xnor U15195 (N_15195,N_12899,N_13501);
and U15196 (N_15196,N_13921,N_12973);
or U15197 (N_15197,N_12568,N_13906);
or U15198 (N_15198,N_14668,N_12022);
nor U15199 (N_15199,N_14765,N_11696);
nand U15200 (N_15200,N_11676,N_14411);
nand U15201 (N_15201,N_11126,N_13302);
and U15202 (N_15202,N_11423,N_14825);
and U15203 (N_15203,N_13520,N_12608);
nor U15204 (N_15204,N_10805,N_10127);
nor U15205 (N_15205,N_13202,N_10007);
xnor U15206 (N_15206,N_11507,N_12547);
or U15207 (N_15207,N_12117,N_12611);
nand U15208 (N_15208,N_10281,N_10846);
nor U15209 (N_15209,N_14468,N_12904);
nand U15210 (N_15210,N_13155,N_12737);
and U15211 (N_15211,N_12887,N_14513);
and U15212 (N_15212,N_13080,N_13972);
or U15213 (N_15213,N_10684,N_13710);
or U15214 (N_15214,N_10274,N_14442);
or U15215 (N_15215,N_14072,N_12417);
nor U15216 (N_15216,N_11475,N_11659);
and U15217 (N_15217,N_12783,N_14872);
xor U15218 (N_15218,N_10668,N_11818);
xor U15219 (N_15219,N_12489,N_13952);
nand U15220 (N_15220,N_13390,N_14337);
or U15221 (N_15221,N_14622,N_12613);
or U15222 (N_15222,N_14820,N_13529);
nand U15223 (N_15223,N_11222,N_11890);
nor U15224 (N_15224,N_13585,N_11589);
and U15225 (N_15225,N_10205,N_12094);
or U15226 (N_15226,N_11467,N_14474);
nand U15227 (N_15227,N_13625,N_11965);
or U15228 (N_15228,N_13543,N_13024);
nand U15229 (N_15229,N_14687,N_14216);
nand U15230 (N_15230,N_13239,N_11761);
and U15231 (N_15231,N_13362,N_12890);
or U15232 (N_15232,N_11754,N_12922);
nand U15233 (N_15233,N_14967,N_11248);
and U15234 (N_15234,N_13331,N_14488);
or U15235 (N_15235,N_11278,N_14435);
nand U15236 (N_15236,N_13916,N_14739);
xnor U15237 (N_15237,N_12731,N_10930);
and U15238 (N_15238,N_13059,N_11967);
or U15239 (N_15239,N_12286,N_14280);
nand U15240 (N_15240,N_12641,N_12355);
nand U15241 (N_15241,N_11129,N_13780);
nor U15242 (N_15242,N_11863,N_14639);
nor U15243 (N_15243,N_14180,N_12880);
xor U15244 (N_15244,N_13499,N_10021);
and U15245 (N_15245,N_13422,N_12738);
xor U15246 (N_15246,N_14877,N_13657);
nand U15247 (N_15247,N_14315,N_12025);
xor U15248 (N_15248,N_14079,N_14247);
or U15249 (N_15249,N_14686,N_14062);
and U15250 (N_15250,N_11982,N_14641);
xnor U15251 (N_15251,N_12642,N_14376);
nor U15252 (N_15252,N_11435,N_12771);
nor U15253 (N_15253,N_11406,N_13669);
and U15254 (N_15254,N_14708,N_10890);
nand U15255 (N_15255,N_13129,N_11440);
and U15256 (N_15256,N_13630,N_12418);
nand U15257 (N_15257,N_12378,N_12315);
nand U15258 (N_15258,N_10391,N_11672);
nor U15259 (N_15259,N_11678,N_13933);
nor U15260 (N_15260,N_11987,N_11267);
nand U15261 (N_15261,N_13125,N_12115);
or U15262 (N_15262,N_10243,N_14746);
or U15263 (N_15263,N_11718,N_12125);
and U15264 (N_15264,N_10794,N_14467);
xor U15265 (N_15265,N_13176,N_10341);
or U15266 (N_15266,N_13733,N_12882);
or U15267 (N_15267,N_12599,N_11030);
and U15268 (N_15268,N_13504,N_11036);
and U15269 (N_15269,N_12146,N_13227);
xnor U15270 (N_15270,N_13293,N_10119);
and U15271 (N_15271,N_10078,N_11788);
and U15272 (N_15272,N_13347,N_12574);
xnor U15273 (N_15273,N_11377,N_12216);
and U15274 (N_15274,N_12249,N_13606);
nand U15275 (N_15275,N_12472,N_11904);
or U15276 (N_15276,N_11549,N_14172);
xnor U15277 (N_15277,N_10040,N_13215);
nor U15278 (N_15278,N_12631,N_13686);
xor U15279 (N_15279,N_12525,N_14374);
xnor U15280 (N_15280,N_12988,N_12294);
xnor U15281 (N_15281,N_13737,N_14723);
nor U15282 (N_15282,N_12260,N_10314);
and U15283 (N_15283,N_10557,N_14182);
and U15284 (N_15284,N_11434,N_11415);
or U15285 (N_15285,N_12238,N_11114);
or U15286 (N_15286,N_12958,N_12516);
nand U15287 (N_15287,N_10218,N_13654);
nand U15288 (N_15288,N_13030,N_10038);
nand U15289 (N_15289,N_12246,N_14995);
nand U15290 (N_15290,N_10492,N_13050);
nand U15291 (N_15291,N_14367,N_13111);
and U15292 (N_15292,N_10228,N_10015);
or U15293 (N_15293,N_10229,N_12154);
xor U15294 (N_15294,N_13755,N_14969);
and U15295 (N_15295,N_14155,N_11269);
nor U15296 (N_15296,N_14430,N_12652);
and U15297 (N_15297,N_12282,N_10595);
or U15298 (N_15298,N_14703,N_12030);
nand U15299 (N_15299,N_12886,N_11260);
and U15300 (N_15300,N_14695,N_13500);
xnor U15301 (N_15301,N_13058,N_11685);
nand U15302 (N_15302,N_13693,N_12497);
xnor U15303 (N_15303,N_14193,N_11561);
or U15304 (N_15304,N_13229,N_12466);
or U15305 (N_15305,N_10261,N_12093);
xnor U15306 (N_15306,N_10238,N_12056);
xor U15307 (N_15307,N_10134,N_12350);
or U15308 (N_15308,N_13262,N_12976);
and U15309 (N_15309,N_10615,N_13451);
nor U15310 (N_15310,N_12214,N_11041);
nor U15311 (N_15311,N_13827,N_12815);
nand U15312 (N_15312,N_11622,N_10320);
xor U15313 (N_15313,N_12586,N_11487);
nor U15314 (N_15314,N_14436,N_10700);
and U15315 (N_15315,N_12256,N_10270);
xnor U15316 (N_15316,N_13484,N_11257);
and U15317 (N_15317,N_11931,N_11880);
nor U15318 (N_15318,N_13511,N_11290);
nand U15319 (N_15319,N_13406,N_13869);
and U15320 (N_15320,N_12580,N_12097);
or U15321 (N_15321,N_11905,N_13592);
or U15322 (N_15322,N_12012,N_12506);
nor U15323 (N_15323,N_11521,N_12433);
or U15324 (N_15324,N_14769,N_13498);
and U15325 (N_15325,N_13246,N_11109);
and U15326 (N_15326,N_14660,N_10712);
nor U15327 (N_15327,N_13704,N_10125);
xor U15328 (N_15328,N_13091,N_13144);
nand U15329 (N_15329,N_12048,N_14541);
nand U15330 (N_15330,N_12575,N_14473);
or U15331 (N_15331,N_13649,N_11439);
or U15332 (N_15332,N_12703,N_10226);
nand U15333 (N_15333,N_10392,N_10498);
nand U15334 (N_15334,N_10372,N_11968);
nor U15335 (N_15335,N_10536,N_13757);
or U15336 (N_15336,N_10533,N_13789);
xnor U15337 (N_15337,N_13276,N_12535);
nand U15338 (N_15338,N_10311,N_12780);
nand U15339 (N_15339,N_10245,N_11059);
nor U15340 (N_15340,N_11108,N_12908);
xnor U15341 (N_15341,N_14899,N_14750);
nand U15342 (N_15342,N_10606,N_13333);
and U15343 (N_15343,N_14190,N_14941);
and U15344 (N_15344,N_14233,N_14237);
and U15345 (N_15345,N_10408,N_13694);
or U15346 (N_15346,N_12412,N_10535);
or U15347 (N_15347,N_12929,N_12847);
xor U15348 (N_15348,N_10612,N_13535);
nor U15349 (N_15349,N_14834,N_14051);
nor U15350 (N_15350,N_11595,N_14728);
nand U15351 (N_15351,N_10647,N_14824);
xnor U15352 (N_15352,N_11796,N_11554);
xnor U15353 (N_15353,N_12266,N_13913);
or U15354 (N_15354,N_14391,N_14276);
nor U15355 (N_15355,N_13388,N_11520);
or U15356 (N_15356,N_10593,N_13919);
nand U15357 (N_15357,N_13425,N_14757);
or U15358 (N_15358,N_10529,N_11255);
xor U15359 (N_15359,N_11906,N_11803);
and U15360 (N_15360,N_13665,N_11452);
nor U15361 (N_15361,N_11760,N_12223);
nand U15362 (N_15362,N_11292,N_11274);
nand U15363 (N_15363,N_14662,N_14923);
nand U15364 (N_15364,N_10452,N_10998);
or U15365 (N_15365,N_14627,N_12131);
and U15366 (N_15366,N_14506,N_10499);
nand U15367 (N_15367,N_14241,N_14866);
xor U15368 (N_15368,N_10605,N_13413);
nand U15369 (N_15369,N_10708,N_13719);
nand U15370 (N_15370,N_10783,N_14425);
nand U15371 (N_15371,N_10494,N_11409);
or U15372 (N_15372,N_11747,N_11745);
and U15373 (N_15373,N_13655,N_11646);
and U15374 (N_15374,N_14992,N_14002);
nor U15375 (N_15375,N_14630,N_11865);
nor U15376 (N_15376,N_10627,N_14158);
or U15377 (N_15377,N_13263,N_14218);
nand U15378 (N_15378,N_14418,N_14000);
nand U15379 (N_15379,N_12868,N_12894);
nand U15380 (N_15380,N_10043,N_12720);
nand U15381 (N_15381,N_12957,N_10661);
xnor U15382 (N_15382,N_10891,N_13376);
xor U15383 (N_15383,N_11221,N_10654);
nand U15384 (N_15384,N_11217,N_12563);
or U15385 (N_15385,N_14857,N_12215);
nand U15386 (N_15386,N_11220,N_13788);
nand U15387 (N_15387,N_11280,N_10067);
nand U15388 (N_15388,N_10064,N_14369);
and U15389 (N_15389,N_13999,N_11077);
nand U15390 (N_15390,N_10962,N_12590);
xor U15391 (N_15391,N_13743,N_11422);
xnor U15392 (N_15392,N_10014,N_14323);
and U15393 (N_15393,N_10729,N_10221);
or U15394 (N_15394,N_14701,N_11273);
nand U15395 (N_15395,N_11876,N_13567);
nand U15396 (N_15396,N_11509,N_14716);
nor U15397 (N_15397,N_13415,N_11601);
or U15398 (N_15398,N_12500,N_13014);
xnor U15399 (N_15399,N_12311,N_13853);
nand U15400 (N_15400,N_10546,N_12269);
and U15401 (N_15401,N_11988,N_14745);
xor U15402 (N_15402,N_11330,N_10165);
nor U15403 (N_15403,N_11797,N_10363);
or U15404 (N_15404,N_12191,N_13929);
nand U15405 (N_15405,N_10103,N_12764);
and U15406 (N_15406,N_10225,N_11083);
nand U15407 (N_15407,N_14300,N_11935);
or U15408 (N_15408,N_10822,N_12679);
nand U15409 (N_15409,N_11016,N_13366);
nor U15410 (N_15410,N_14542,N_10268);
nor U15411 (N_15411,N_12519,N_12852);
or U15412 (N_15412,N_12715,N_11699);
nor U15413 (N_15413,N_10252,N_11304);
nor U15414 (N_15414,N_14868,N_13615);
nand U15415 (N_15415,N_12782,N_10434);
and U15416 (N_15416,N_13479,N_14173);
or U15417 (N_15417,N_13717,N_10470);
nor U15418 (N_15418,N_10387,N_13443);
or U15419 (N_15419,N_11265,N_13901);
and U15420 (N_15420,N_12651,N_14958);
or U15421 (N_15421,N_10574,N_12234);
nand U15422 (N_15422,N_10297,N_13638);
xnor U15423 (N_15423,N_14591,N_13983);
nor U15424 (N_15424,N_12265,N_12807);
xnor U15425 (N_15425,N_11098,N_14564);
nor U15426 (N_15426,N_10711,N_10604);
nand U15427 (N_15427,N_11944,N_13029);
nor U15428 (N_15428,N_13731,N_10806);
nor U15429 (N_15429,N_10682,N_10706);
nor U15430 (N_15430,N_12933,N_13960);
or U15431 (N_15431,N_13426,N_14700);
xor U15432 (N_15432,N_14905,N_12443);
xor U15433 (N_15433,N_14134,N_10417);
or U15434 (N_15434,N_14165,N_14084);
and U15435 (N_15435,N_12354,N_11147);
and U15436 (N_15436,N_14264,N_10800);
or U15437 (N_15437,N_13631,N_14556);
nor U15438 (N_15438,N_13466,N_11878);
xnor U15439 (N_15439,N_13402,N_14342);
nor U15440 (N_15440,N_14243,N_13832);
nor U15441 (N_15441,N_10659,N_13911);
and U15442 (N_15442,N_12626,N_12730);
nand U15443 (N_15443,N_13387,N_14458);
nor U15444 (N_15444,N_10300,N_13196);
and U15445 (N_15445,N_10915,N_12322);
nor U15446 (N_15446,N_12967,N_14791);
nor U15447 (N_15447,N_12167,N_10396);
nor U15448 (N_15448,N_10899,N_12747);
and U15449 (N_15449,N_14160,N_13022);
xor U15450 (N_15450,N_11531,N_10056);
and U15451 (N_15451,N_11347,N_14719);
nor U15452 (N_15452,N_13275,N_11091);
or U15453 (N_15453,N_11851,N_14934);
and U15454 (N_15454,N_14253,N_14485);
and U15455 (N_15455,N_13165,N_12842);
xor U15456 (N_15456,N_13830,N_13090);
nand U15457 (N_15457,N_12106,N_10773);
and U15458 (N_15458,N_13551,N_10032);
nor U15459 (N_15459,N_12491,N_10852);
nor U15460 (N_15460,N_14067,N_14349);
nor U15461 (N_15461,N_13106,N_14782);
nor U15462 (N_15462,N_13871,N_14546);
or U15463 (N_15463,N_14149,N_11463);
nor U15464 (N_15464,N_11875,N_12853);
xor U15465 (N_15465,N_10992,N_13962);
nand U15466 (N_15466,N_14988,N_12145);
nand U15467 (N_15467,N_13702,N_10919);
nor U15468 (N_15468,N_12381,N_11334);
nand U15469 (N_15469,N_12911,N_13265);
nor U15470 (N_15470,N_10414,N_12729);
nor U15471 (N_15471,N_14942,N_10756);
or U15472 (N_15472,N_10410,N_11571);
nor U15473 (N_15473,N_12577,N_12036);
nor U15474 (N_15474,N_14515,N_11236);
xor U15475 (N_15475,N_12494,N_10948);
or U15476 (N_15476,N_14895,N_11655);
and U15477 (N_15477,N_13556,N_11533);
xnor U15478 (N_15478,N_11526,N_11853);
xor U15479 (N_15479,N_10095,N_14944);
xnor U15480 (N_15480,N_10462,N_10985);
nand U15481 (N_15481,N_12384,N_11163);
nand U15482 (N_15482,N_13664,N_11682);
nand U15483 (N_15483,N_11949,N_10916);
nor U15484 (N_15484,N_13851,N_10959);
nand U15485 (N_15485,N_13483,N_13213);
and U15486 (N_15486,N_10954,N_11169);
and U15487 (N_15487,N_12011,N_10359);
nor U15488 (N_15488,N_10636,N_10104);
or U15489 (N_15489,N_12187,N_13714);
and U15490 (N_15490,N_14758,N_14952);
nand U15491 (N_15491,N_11062,N_12252);
nand U15492 (N_15492,N_14061,N_11183);
and U15493 (N_15493,N_10505,N_11698);
nor U15494 (N_15494,N_13754,N_11179);
and U15495 (N_15495,N_13025,N_14685);
nor U15496 (N_15496,N_10895,N_12785);
xor U15497 (N_15497,N_13341,N_14015);
or U15498 (N_15498,N_13491,N_11502);
and U15499 (N_15499,N_10545,N_13800);
nand U15500 (N_15500,N_12840,N_14837);
and U15501 (N_15501,N_11639,N_12018);
nor U15502 (N_15502,N_12776,N_14206);
and U15503 (N_15503,N_11264,N_10185);
or U15504 (N_15504,N_13903,N_11835);
and U15505 (N_15505,N_14535,N_14520);
nor U15506 (N_15506,N_12464,N_13021);
xnor U15507 (N_15507,N_13922,N_10669);
nand U15508 (N_15508,N_11097,N_14840);
or U15509 (N_15509,N_13750,N_14512);
nand U15510 (N_15510,N_11444,N_11581);
and U15511 (N_15511,N_12901,N_10247);
nand U15512 (N_15512,N_10672,N_11063);
nor U15513 (N_15513,N_11732,N_12965);
nor U15514 (N_15514,N_12085,N_10237);
nor U15515 (N_15515,N_12201,N_14672);
and U15516 (N_15516,N_12546,N_13968);
and U15517 (N_15517,N_14354,N_12656);
or U15518 (N_15518,N_14235,N_11087);
nor U15519 (N_15519,N_10106,N_14221);
or U15520 (N_15520,N_11375,N_10292);
and U15521 (N_15521,N_13748,N_12471);
or U15522 (N_15522,N_14377,N_11606);
nor U15523 (N_15523,N_12826,N_10330);
and U15524 (N_15524,N_12700,N_10306);
nor U15525 (N_15525,N_14492,N_13875);
and U15526 (N_15526,N_13744,N_13724);
nand U15527 (N_15527,N_10288,N_13218);
and U15528 (N_15528,N_12033,N_11146);
and U15529 (N_15529,N_14976,N_11660);
nand U15530 (N_15530,N_14536,N_10942);
or U15531 (N_15531,N_10749,N_12837);
or U15532 (N_15532,N_11588,N_12517);
xnor U15533 (N_15533,N_13296,N_13020);
or U15534 (N_15534,N_13109,N_11846);
xor U15535 (N_15535,N_12757,N_10881);
nand U15536 (N_15536,N_13146,N_12806);
xnor U15537 (N_15537,N_11626,N_12076);
nor U15538 (N_15538,N_12609,N_14073);
nor U15539 (N_15539,N_14655,N_11722);
or U15540 (N_15540,N_14484,N_12619);
nand U15541 (N_15541,N_10164,N_11208);
and U15542 (N_15542,N_12571,N_10401);
xor U15543 (N_15543,N_10145,N_11838);
nor U15544 (N_15544,N_10511,N_11344);
nand U15545 (N_15545,N_13530,N_12241);
nand U15546 (N_15546,N_14609,N_11188);
nand U15547 (N_15547,N_11930,N_11389);
nand U15548 (N_15548,N_14897,N_12006);
xnor U15549 (N_15549,N_13382,N_11957);
xor U15550 (N_15550,N_11726,N_11362);
nor U15551 (N_15551,N_14978,N_10380);
xor U15552 (N_15552,N_10563,N_10010);
nand U15553 (N_15553,N_11092,N_10405);
xnor U15554 (N_15554,N_11336,N_14296);
xnor U15555 (N_15555,N_10474,N_12428);
nor U15556 (N_15556,N_12504,N_13545);
xnor U15557 (N_15557,N_11959,N_10873);
or U15558 (N_15558,N_13516,N_14178);
nand U15559 (N_15559,N_10662,N_13943);
or U15560 (N_15560,N_10847,N_13170);
nor U15561 (N_15561,N_12258,N_11920);
or U15562 (N_15562,N_12440,N_12588);
and U15563 (N_15563,N_12480,N_10045);
nor U15564 (N_15564,N_12181,N_10825);
xor U15565 (N_15565,N_12724,N_13222);
nor U15566 (N_15566,N_12770,N_12308);
and U15567 (N_15567,N_12912,N_13775);
or U15568 (N_15568,N_14465,N_14379);
xor U15569 (N_15569,N_11008,N_13000);
xor U15570 (N_15570,N_14950,N_11513);
nor U15571 (N_15571,N_13135,N_10926);
nand U15572 (N_15572,N_13340,N_14157);
or U15573 (N_15573,N_14702,N_11195);
or U15574 (N_15574,N_12259,N_14581);
xor U15575 (N_15575,N_10680,N_10035);
nor U15576 (N_15576,N_12073,N_13346);
xnor U15577 (N_15577,N_13978,N_13114);
nor U15578 (N_15578,N_12474,N_13473);
or U15579 (N_15579,N_10877,N_13923);
xnor U15580 (N_15580,N_13891,N_10500);
xor U15581 (N_15581,N_13235,N_11945);
nor U15582 (N_15582,N_11155,N_11913);
or U15583 (N_15583,N_10547,N_14656);
nor U15584 (N_15584,N_12114,N_13280);
xor U15585 (N_15585,N_14128,N_11579);
nor U15586 (N_15586,N_13446,N_10579);
nor U15587 (N_15587,N_11771,N_10133);
nor U15588 (N_15588,N_11393,N_10746);
nor U15589 (N_15589,N_12910,N_14912);
nand U15590 (N_15590,N_14756,N_12891);
and U15591 (N_15591,N_10109,N_11268);
or U15592 (N_15592,N_11033,N_10153);
xnor U15593 (N_15593,N_14023,N_14439);
nor U15594 (N_15594,N_12400,N_11039);
xnor U15595 (N_15595,N_11667,N_14998);
and U15596 (N_15596,N_12907,N_11096);
or U15597 (N_15597,N_14652,N_13110);
or U15598 (N_15598,N_10660,N_11498);
nand U15599 (N_15599,N_10335,N_12671);
nor U15600 (N_15600,N_13712,N_13643);
xor U15601 (N_15601,N_13253,N_11256);
xnor U15602 (N_15602,N_10970,N_14804);
nand U15603 (N_15603,N_12824,N_12705);
nand U15604 (N_15604,N_13525,N_11289);
or U15605 (N_15605,N_11332,N_11327);
nor U15606 (N_15606,N_14105,N_11517);
nand U15607 (N_15607,N_13191,N_14705);
nor U15608 (N_15608,N_11105,N_11557);
or U15609 (N_15609,N_14048,N_13703);
nand U15610 (N_15610,N_12567,N_13187);
and U15611 (N_15611,N_10028,N_14754);
and U15612 (N_15612,N_12745,N_13992);
nor U15613 (N_15613,N_10331,N_12430);
nand U15614 (N_15614,N_14673,N_11736);
nand U15615 (N_15615,N_13452,N_11266);
nand U15616 (N_15616,N_11072,N_12463);
nor U15617 (N_15617,N_13699,N_13060);
xor U15618 (N_15618,N_11777,N_14021);
or U15619 (N_15619,N_14838,N_11947);
nand U15620 (N_15620,N_12884,N_13095);
xor U15621 (N_15621,N_10074,N_11907);
xor U15622 (N_15622,N_12520,N_13345);
and U15623 (N_15623,N_14078,N_13204);
and U15624 (N_15624,N_14808,N_12208);
or U15625 (N_15625,N_12478,N_10561);
nand U15626 (N_15626,N_12318,N_14334);
xnor U15627 (N_15627,N_10360,N_10233);
or U15628 (N_15628,N_14316,N_11564);
xor U15629 (N_15629,N_11697,N_12391);
and U15630 (N_15630,N_10493,N_14452);
or U15631 (N_15631,N_13831,N_11132);
nand U15632 (N_15632,N_10329,N_13131);
nand U15633 (N_15633,N_10257,N_13688);
xnor U15634 (N_15634,N_10213,N_10602);
or U15635 (N_15635,N_12835,N_14288);
and U15636 (N_15636,N_11230,N_10943);
xor U15637 (N_15637,N_10503,N_11385);
xnor U15638 (N_15638,N_14091,N_10620);
and U15639 (N_15639,N_11864,N_11175);
nand U15640 (N_15640,N_13077,N_12219);
and U15641 (N_15641,N_11538,N_10886);
or U15642 (N_15642,N_14565,N_10515);
nor U15643 (N_15643,N_13635,N_11421);
or U15644 (N_15644,N_13228,N_10192);
nor U15645 (N_15645,N_10305,N_11692);
xor U15646 (N_15646,N_11166,N_14055);
xnor U15647 (N_15647,N_14118,N_14244);
or U15648 (N_15648,N_10117,N_12481);
xnor U15649 (N_15649,N_10302,N_14226);
and U15650 (N_15650,N_11821,N_14986);
or U15651 (N_15651,N_11370,N_13149);
and U15652 (N_15652,N_11461,N_14606);
nor U15653 (N_15653,N_14050,N_13433);
and U15654 (N_15654,N_11159,N_12692);
xnor U15655 (N_15655,N_13961,N_12057);
nand U15656 (N_15656,N_13350,N_14027);
xor U15657 (N_15657,N_11110,N_10214);
nand U15658 (N_15658,N_14052,N_12292);
or U15659 (N_15659,N_14677,N_11356);
nand U15660 (N_15660,N_10169,N_13485);
xor U15661 (N_15661,N_13399,N_13320);
xor U15662 (N_15662,N_10619,N_11238);
and U15663 (N_15663,N_12263,N_13998);
nand U15664 (N_15664,N_13271,N_13445);
xnor U15665 (N_15665,N_14187,N_10947);
or U15666 (N_15666,N_10005,N_12328);
and U15667 (N_15667,N_11443,N_13016);
and U15668 (N_15668,N_10339,N_10793);
nand U15669 (N_15669,N_11657,N_10910);
xor U15670 (N_15670,N_11032,N_13609);
nor U15671 (N_15671,N_11076,N_12333);
or U15672 (N_15672,N_11333,N_12037);
nor U15673 (N_15673,N_10691,N_11198);
or U15674 (N_15674,N_14371,N_13863);
or U15675 (N_15675,N_14928,N_11691);
nand U15676 (N_15676,N_10698,N_11176);
xnor U15677 (N_15677,N_14968,N_10093);
nor U15678 (N_15678,N_12276,N_11820);
nand U15679 (N_15679,N_13206,N_11734);
or U15680 (N_15680,N_11542,N_14329);
or U15681 (N_15681,N_10356,N_11814);
and U15682 (N_15682,N_14625,N_14166);
and U15683 (N_15683,N_13104,N_12992);
and U15684 (N_15684,N_10921,N_13752);
and U15685 (N_15685,N_10696,N_11598);
xor U15686 (N_15686,N_13794,N_13338);
nor U15687 (N_15687,N_12281,N_13618);
nand U15688 (N_15688,N_11367,N_10473);
or U15689 (N_15689,N_13722,N_11600);
xor U15690 (N_15690,N_11161,N_11384);
xnor U15691 (N_15691,N_11429,N_14773);
xor U15692 (N_15692,N_11537,N_13461);
or U15693 (N_15693,N_12804,N_10362);
or U15694 (N_15694,N_12177,N_13771);
nor U15695 (N_15695,N_10046,N_14610);
or U15696 (N_15696,N_12370,N_12961);
xnor U15697 (N_15697,N_11934,N_14338);
nand U15698 (N_15698,N_11998,N_14242);
nand U15699 (N_15699,N_14984,N_12512);
and U15700 (N_15700,N_14326,N_12936);
or U15701 (N_15701,N_13591,N_11164);
xor U15702 (N_15702,N_11897,N_11453);
nor U15703 (N_15703,N_14286,N_10963);
and U15704 (N_15704,N_11778,N_13061);
or U15705 (N_15705,N_14993,N_14441);
xnor U15706 (N_15706,N_10542,N_13138);
xor U15707 (N_15707,N_11449,N_12818);
nand U15708 (N_15708,N_12702,N_10928);
nor U15709 (N_15709,N_14164,N_14860);
and U15710 (N_15710,N_10905,N_11632);
nand U15711 (N_15711,N_11148,N_11790);
nand U15712 (N_15712,N_12230,N_14878);
nand U15713 (N_15713,N_14313,N_10342);
and U15714 (N_15714,N_13193,N_14198);
nor U15715 (N_15715,N_12775,N_14859);
nor U15716 (N_15716,N_13282,N_14628);
or U15717 (N_15717,N_10406,N_14036);
or U15718 (N_15718,N_14302,N_13661);
or U15719 (N_15719,N_14711,N_14698);
and U15720 (N_15720,N_10319,N_14282);
and U15721 (N_15721,N_12064,N_10186);
and U15722 (N_15722,N_11404,N_14281);
nor U15723 (N_15723,N_14731,N_12711);
nand U15724 (N_15724,N_11528,N_14846);
nor U15725 (N_15725,N_12051,N_10114);
or U15726 (N_15726,N_10643,N_12137);
and U15727 (N_15727,N_13469,N_11550);
or U15728 (N_15728,N_14661,N_10148);
or U15729 (N_15729,N_14684,N_13565);
and U15730 (N_15730,N_13259,N_10710);
or U15731 (N_15731,N_12188,N_13860);
nand U15732 (N_15732,N_10866,N_12970);
nor U15733 (N_15733,N_11186,N_11471);
and U15734 (N_15734,N_12149,N_13113);
nand U15735 (N_15735,N_11490,N_10562);
and U15736 (N_15736,N_12624,N_10840);
and U15737 (N_15737,N_11117,N_12606);
and U15738 (N_15738,N_12222,N_14308);
nor U15739 (N_15739,N_13118,N_14767);
and U15740 (N_15740,N_10976,N_12421);
nor U15741 (N_15741,N_14059,N_12706);
and U15742 (N_15742,N_11952,N_12644);
and U15743 (N_15743,N_14478,N_14642);
nand U15744 (N_15744,N_13588,N_11679);
or U15745 (N_15745,N_10350,N_11368);
or U15746 (N_15746,N_12953,N_11364);
xor U15747 (N_15747,N_12742,N_10697);
and U15748 (N_15748,N_13398,N_10423);
or U15749 (N_15749,N_10689,N_14472);
nand U15750 (N_15750,N_11031,N_10263);
nor U15751 (N_15751,N_11113,N_11402);
xor U15752 (N_15752,N_12233,N_11954);
xnor U15753 (N_15753,N_14451,N_11740);
and U15754 (N_15754,N_14736,N_10370);
xnor U15755 (N_15755,N_13666,N_10573);
and U15756 (N_15756,N_13602,N_10220);
nand U15757 (N_15757,N_14768,N_13804);
and U15758 (N_15758,N_13453,N_10885);
or U15759 (N_15759,N_11341,N_10514);
nand U15760 (N_15760,N_13158,N_10459);
nand U15761 (N_15761,N_10174,N_13488);
nand U15762 (N_15762,N_12089,N_11832);
nand U15763 (N_15763,N_12593,N_12189);
xor U15764 (N_15764,N_13808,N_14130);
or U15765 (N_15765,N_12625,N_12183);
nand U15766 (N_15766,N_12620,N_13153);
and U15767 (N_15767,N_13995,N_11958);
nand U15768 (N_15768,N_14393,N_12784);
nand U15769 (N_15769,N_12304,N_10716);
or U15770 (N_15770,N_13036,N_11674);
nor U15771 (N_15771,N_14508,N_10581);
xnor U15772 (N_15772,N_11530,N_11963);
xor U15773 (N_15773,N_14240,N_10379);
nor U15774 (N_15774,N_12539,N_13233);
nor U15775 (N_15775,N_14262,N_14312);
and U15776 (N_15776,N_14805,N_11671);
and U15777 (N_15777,N_14030,N_10737);
or U15778 (N_15778,N_10249,N_13300);
or U15779 (N_15779,N_10495,N_12598);
and U15780 (N_15780,N_14910,N_10309);
and U15781 (N_15781,N_11350,N_13254);
nand U15782 (N_15782,N_10166,N_14121);
and U15783 (N_15783,N_14856,N_10610);
and U15784 (N_15784,N_14509,N_12264);
xnor U15785 (N_15785,N_10904,N_12113);
or U15786 (N_15786,N_11465,N_12467);
nor U15787 (N_15787,N_12455,N_14285);
xnor U15788 (N_15788,N_12897,N_10743);
and U15789 (N_15789,N_11279,N_10395);
xnor U15790 (N_15790,N_11891,N_13934);
xor U15791 (N_15791,N_11854,N_14629);
and U15792 (N_15792,N_11902,N_12150);
or U15793 (N_15793,N_12811,N_14156);
nand U15794 (N_15794,N_14007,N_10821);
and U15795 (N_15795,N_14191,N_14848);
or U15796 (N_15796,N_11942,N_12821);
nor U15797 (N_15797,N_12323,N_12663);
and U15798 (N_15798,N_10554,N_12274);
xnor U15799 (N_15799,N_10455,N_10446);
or U15800 (N_15800,N_11544,N_12059);
or U15801 (N_15801,N_12697,N_14386);
xnor U15802 (N_15802,N_14258,N_13019);
xor U15803 (N_15803,N_13521,N_12950);
or U15804 (N_15804,N_11197,N_12915);
nand U15805 (N_15805,N_12565,N_10287);
and U15806 (N_15806,N_14385,N_13910);
and U15807 (N_15807,N_11120,N_14291);
nand U15808 (N_15808,N_14487,N_12573);
nand U15809 (N_15809,N_13247,N_11553);
nor U15810 (N_15810,N_11516,N_10872);
xnor U15811 (N_15811,N_11663,N_13045);
and U15812 (N_15812,N_14077,N_13006);
nand U15813 (N_15813,N_10967,N_14955);
and U15814 (N_15814,N_12343,N_12217);
nor U15815 (N_15815,N_13732,N_12377);
and U15816 (N_15816,N_12134,N_14945);
nand U15817 (N_15817,N_10484,N_11061);
and U15818 (N_15818,N_10789,N_10940);
and U15819 (N_15819,N_12712,N_12190);
and U15820 (N_15820,N_12162,N_11203);
and U15821 (N_15821,N_11099,N_11603);
nor U15822 (N_15822,N_13990,N_12348);
or U15823 (N_15823,N_11335,N_11824);
nor U15824 (N_15824,N_13578,N_14793);
nor U15825 (N_15825,N_11787,N_11594);
nor U15826 (N_15826,N_11565,N_13596);
nor U15827 (N_15827,N_11190,N_12017);
and U15828 (N_15828,N_12193,N_13243);
and U15829 (N_15829,N_10107,N_13955);
nand U15830 (N_15830,N_14605,N_13695);
nor U15831 (N_15831,N_10553,N_14408);
and U15832 (N_15832,N_11653,N_14819);
and U15833 (N_15833,N_13378,N_10193);
and U15834 (N_15834,N_12503,N_14823);
xor U15835 (N_15835,N_10276,N_10303);
and U15836 (N_15836,N_13156,N_11995);
nor U15837 (N_15837,N_13074,N_11157);
and U15838 (N_15838,N_11149,N_12127);
or U15839 (N_15839,N_13539,N_12822);
or U15840 (N_15840,N_11437,N_10296);
and U15841 (N_15841,N_11447,N_14595);
nor U15842 (N_15842,N_13419,N_11456);
nor U15843 (N_15843,N_11312,N_12101);
xnor U15844 (N_15844,N_11980,N_14047);
nor U15845 (N_15845,N_14398,N_11433);
and U15846 (N_15846,N_14545,N_10603);
or U15847 (N_15847,N_10784,N_11640);
xnor U15848 (N_15848,N_10809,N_13801);
nand U15849 (N_15849,N_14674,N_11458);
nand U15850 (N_15850,N_13797,N_12227);
and U15851 (N_15851,N_12778,N_13167);
nor U15852 (N_15852,N_14318,N_11070);
nor U15853 (N_15853,N_13985,N_10223);
xor U15854 (N_15854,N_13745,N_13278);
nand U15855 (N_15855,N_14068,N_14481);
and U15856 (N_15856,N_10111,N_14268);
nand U15857 (N_15857,N_12921,N_13379);
nand U15858 (N_15858,N_12415,N_14401);
or U15859 (N_15859,N_11536,N_11580);
nor U15860 (N_15860,N_11202,N_10065);
nand U15861 (N_15861,N_12597,N_10988);
nor U15862 (N_15862,N_10686,N_13611);
xnor U15863 (N_15863,N_12411,N_12530);
or U15864 (N_15864,N_10259,N_12447);
xor U15865 (N_15865,N_11881,N_10447);
xnor U15866 (N_15866,N_10576,N_14136);
nand U15867 (N_15867,N_10424,N_10803);
nand U15868 (N_15868,N_13147,N_10933);
or U15869 (N_15869,N_14632,N_11215);
xor U15870 (N_15870,N_11857,N_14251);
nor U15871 (N_15871,N_14994,N_10176);
xnor U15872 (N_15872,N_12148,N_10020);
nand U15873 (N_15873,N_13367,N_14884);
nor U15874 (N_15874,N_14462,N_10941);
nor U15875 (N_15875,N_10714,N_13982);
nor U15876 (N_15876,N_14689,N_12435);
and U15877 (N_15877,N_12969,N_12509);
and U15878 (N_15878,N_11205,N_13041);
or U15879 (N_15879,N_14697,N_14813);
nor U15880 (N_15880,N_14220,N_11313);
nor U15881 (N_15881,N_12643,N_12751);
xor U15882 (N_15882,N_12498,N_13826);
nand U15883 (N_15883,N_13793,N_12477);
nor U15884 (N_15884,N_14448,N_14370);
nand U15885 (N_15885,N_10731,N_13481);
or U15886 (N_15886,N_11446,N_12242);
nand U15887 (N_15887,N_11689,N_13183);
and U15888 (N_15888,N_14637,N_14012);
nor U15889 (N_15889,N_12889,N_14681);
nor U15890 (N_15890,N_14651,N_12527);
nand U15891 (N_15891,N_11359,N_13427);
or U15892 (N_15892,N_12357,N_10747);
nor U15893 (N_15893,N_13486,N_13988);
and U15894 (N_15894,N_14097,N_10179);
nor U15895 (N_15895,N_14310,N_13577);
or U15896 (N_15896,N_12528,N_12513);
nor U15897 (N_15897,N_11106,N_14675);
xnor U15898 (N_15898,N_13964,N_11972);
and U15899 (N_15899,N_13351,N_13079);
xor U15900 (N_15900,N_12465,N_10431);
xnor U15901 (N_15901,N_12532,N_12027);
xnor U15902 (N_15902,N_13904,N_13679);
nor U15903 (N_15903,N_11261,N_13309);
or U15904 (N_15904,N_13786,N_13335);
or U15905 (N_15905,N_13524,N_13550);
and U15906 (N_15906,N_10848,N_13391);
xnor U15907 (N_15907,N_10857,N_11866);
or U15908 (N_15908,N_13123,N_12855);
nor U15909 (N_15909,N_13084,N_10428);
xnor U15910 (N_15910,N_10798,N_13356);
nor U15911 (N_15911,N_14192,N_12133);
or U15912 (N_15912,N_11104,N_14426);
or U15913 (N_15913,N_14885,N_11329);
nor U15914 (N_15914,N_14602,N_14650);
nor U15915 (N_15915,N_14779,N_11293);
and U15916 (N_15916,N_14579,N_13644);
and U15917 (N_15917,N_13471,N_10411);
nor U15918 (N_15918,N_11620,N_14227);
and U15919 (N_15919,N_11505,N_12896);
xnor U15920 (N_15920,N_14219,N_13092);
nand U15921 (N_15921,N_10024,N_13064);
xor U15922 (N_15922,N_12502,N_11704);
xor U15923 (N_15923,N_10867,N_11355);
xor U15924 (N_15924,N_12424,N_12353);
nor U15925 (N_15925,N_11703,N_13617);
or U15926 (N_15926,N_12002,N_11028);
and U15927 (N_15927,N_11977,N_14405);
nor U15928 (N_15928,N_12075,N_11245);
and U15929 (N_15929,N_13971,N_11024);
xnor U15930 (N_15930,N_12451,N_10308);
or U15931 (N_15931,N_13692,N_12329);
nor U15932 (N_15932,N_10600,N_14707);
or U15933 (N_15933,N_13112,N_11939);
nor U15934 (N_15934,N_13468,N_10632);
and U15935 (N_15935,N_13032,N_10236);
nor U15936 (N_15936,N_10975,N_10555);
xnor U15937 (N_15937,N_10983,N_10086);
nand U15938 (N_15938,N_14543,N_12584);
and U15939 (N_15939,N_14889,N_14572);
nand U15940 (N_15940,N_14841,N_14892);
and U15941 (N_15941,N_10354,N_14167);
or U15942 (N_15942,N_14918,N_11428);
nor U15943 (N_15943,N_12255,N_10195);
xnor U15944 (N_15944,N_11272,N_12324);
and U15945 (N_15945,N_11879,N_12934);
or U15946 (N_15946,N_11739,N_13647);
nand U15947 (N_15947,N_12696,N_12398);
or U15948 (N_15948,N_11572,N_12218);
and U15949 (N_15949,N_12086,N_10250);
nand U15950 (N_15950,N_14333,N_10264);
and U15951 (N_15951,N_13464,N_13781);
nor U15952 (N_15952,N_14902,N_11207);
or U15953 (N_15953,N_14549,N_14259);
or U15954 (N_15954,N_14350,N_14090);
or U15955 (N_15955,N_10089,N_14987);
xnor U15956 (N_15956,N_11921,N_14306);
nand U15957 (N_15957,N_14387,N_11884);
nand U15958 (N_15958,N_13478,N_12199);
nor U15959 (N_15959,N_11353,N_12066);
xor U15960 (N_15960,N_13528,N_14403);
nor U15961 (N_15961,N_13802,N_14850);
nor U15962 (N_15962,N_10640,N_14284);
nor U15963 (N_15963,N_13736,N_13444);
and U15964 (N_15964,N_12873,N_11567);
nand U15965 (N_15965,N_11345,N_12736);
and U15966 (N_15966,N_10859,N_13787);
nand U15967 (N_15967,N_13944,N_10050);
and U15968 (N_15968,N_13418,N_13221);
nor U15969 (N_15969,N_11253,N_10285);
nor U15970 (N_15970,N_10217,N_11403);
and U15971 (N_15971,N_11843,N_14017);
nand U15972 (N_15972,N_12572,N_13825);
and U15973 (N_15973,N_13034,N_13482);
nor U15974 (N_15974,N_12684,N_13220);
xor U15975 (N_15975,N_10644,N_11758);
or U15976 (N_15976,N_14345,N_11781);
or U15977 (N_15977,N_11064,N_11927);
xor U15978 (N_15978,N_11140,N_11573);
nand U15979 (N_15979,N_13353,N_14438);
nor U15980 (N_15980,N_14990,N_13765);
xor U15981 (N_15981,N_13819,N_12351);
or U15982 (N_15982,N_12406,N_12112);
nor U15983 (N_15983,N_13456,N_13872);
nor U15984 (N_15984,N_14903,N_12155);
nor U15985 (N_15985,N_11473,N_13762);
or U15986 (N_15986,N_10031,N_14638);
nand U15987 (N_15987,N_14608,N_13536);
nand U15988 (N_15988,N_14359,N_11081);
or U15989 (N_15989,N_11116,N_11616);
xnor U15990 (N_15990,N_10159,N_12676);
xnor U15991 (N_15991,N_13926,N_14320);
nor U15992 (N_15992,N_10758,N_10286);
xnor U15993 (N_15993,N_14598,N_14301);
or U15994 (N_15994,N_14640,N_13509);
or U15995 (N_15995,N_13414,N_14997);
and U15996 (N_15996,N_14706,N_10733);
and U15997 (N_15997,N_11025,N_14098);
nand U15998 (N_15998,N_13848,N_11770);
nor U15999 (N_15999,N_14503,N_13514);
and U16000 (N_16000,N_13768,N_13435);
nand U16001 (N_16001,N_13866,N_10075);
xor U16002 (N_16002,N_14266,N_12618);
nor U16003 (N_16003,N_13798,N_12082);
or U16004 (N_16004,N_11683,N_14343);
nand U16005 (N_16005,N_14898,N_12332);
xnor U16006 (N_16006,N_12553,N_14185);
nor U16007 (N_16007,N_10902,N_14340);
nand U16008 (N_16008,N_13354,N_13839);
nor U16009 (N_16009,N_14232,N_12392);
nand U16010 (N_16010,N_12470,N_10824);
nand U16011 (N_16011,N_12989,N_10390);
xnor U16012 (N_16012,N_10202,N_12753);
nand U16013 (N_16013,N_14445,N_11844);
xor U16014 (N_16014,N_12856,N_11476);
nor U16015 (N_16015,N_11816,N_14844);
nor U16016 (N_16016,N_12996,N_12878);
nor U16017 (N_16017,N_10393,N_10977);
and U16018 (N_16018,N_14330,N_14114);
xor U16019 (N_16019,N_10384,N_11871);
xor U16020 (N_16020,N_10944,N_12236);
nor U16021 (N_16021,N_14527,N_14854);
xor U16022 (N_16022,N_14532,N_11361);
or U16023 (N_16023,N_13925,N_12293);
nor U16024 (N_16024,N_13534,N_14116);
xnor U16025 (N_16025,N_10140,N_11174);
or U16026 (N_16026,N_12096,N_12576);
and U16027 (N_16027,N_11379,N_14875);
nor U16028 (N_16028,N_13103,N_13610);
nand U16029 (N_16029,N_10589,N_10909);
xnor U16030 (N_16030,N_11713,N_14906);
or U16031 (N_16031,N_12968,N_10538);
and U16032 (N_16032,N_12860,N_10738);
xor U16033 (N_16033,N_10430,N_14704);
and U16034 (N_16034,N_13552,N_12072);
and U16035 (N_16035,N_10623,N_12848);
xor U16036 (N_16036,N_11765,N_13917);
and U16037 (N_16037,N_12001,N_14303);
nand U16038 (N_16038,N_11644,N_12198);
and U16039 (N_16039,N_12071,N_12169);
nand U16040 (N_16040,N_13884,N_11706);
nand U16041 (N_16041,N_13763,N_10071);
nand U16042 (N_16042,N_14935,N_13380);
and U16043 (N_16043,N_10649,N_10123);
xor U16044 (N_16044,N_13465,N_13377);
nand U16045 (N_16045,N_10699,N_14948);
xor U16046 (N_16046,N_14225,N_10456);
xnor U16047 (N_16047,N_10713,N_12416);
xor U16048 (N_16048,N_10625,N_13590);
nand U16049 (N_16049,N_13531,N_14635);
nand U16050 (N_16050,N_14437,N_13048);
or U16051 (N_16051,N_10139,N_14346);
nand U16052 (N_16052,N_14272,N_12253);
nor U16053 (N_16053,N_11123,N_10098);
and U16054 (N_16054,N_11566,N_10466);
or U16055 (N_16055,N_14683,N_10352);
xnor U16056 (N_16056,N_10725,N_14537);
xnor U16057 (N_16057,N_10762,N_12069);
nand U16058 (N_16058,N_11225,N_13527);
xnor U16059 (N_16059,N_13751,N_12850);
xor U16060 (N_16060,N_11325,N_10791);
nor U16061 (N_16061,N_12061,N_11119);
nand U16062 (N_16062,N_11141,N_11585);
nand U16063 (N_16063,N_12000,N_14283);
nand U16064 (N_16064,N_11497,N_11525);
nor U16065 (N_16065,N_12906,N_12251);
xnor U16066 (N_16066,N_10077,N_12021);
or U16067 (N_16067,N_14290,N_10049);
nor U16068 (N_16068,N_14873,N_13855);
nand U16069 (N_16069,N_12226,N_13143);
xor U16070 (N_16070,N_12419,N_10135);
and U16071 (N_16071,N_11975,N_10066);
nand U16072 (N_16072,N_12371,N_11427);
nand U16073 (N_16073,N_10621,N_12388);
and U16074 (N_16074,N_10340,N_13049);
nand U16075 (N_16075,N_14574,N_11284);
or U16076 (N_16076,N_14382,N_13316);
and U16077 (N_16077,N_14800,N_14321);
and U16078 (N_16078,N_10147,N_13234);
and U16079 (N_16079,N_12956,N_14748);
nor U16080 (N_16080,N_13436,N_13434);
nand U16081 (N_16081,N_11424,N_10770);
nand U16082 (N_16082,N_11784,N_12100);
or U16083 (N_16083,N_11237,N_13162);
nor U16084 (N_16084,N_14028,N_14245);
or U16085 (N_16085,N_10652,N_11239);
xnor U16086 (N_16086,N_12334,N_13023);
xor U16087 (N_16087,N_14938,N_11586);
nor U16088 (N_16088,N_11575,N_10917);
nor U16089 (N_16089,N_10616,N_11811);
nor U16090 (N_16090,N_11649,N_13796);
nor U16091 (N_16091,N_11137,N_13257);
nor U16092 (N_16092,N_11068,N_13767);
and U16093 (N_16093,N_11650,N_10690);
xor U16094 (N_16094,N_11082,N_10069);
nor U16095 (N_16095,N_12658,N_10337);
nor U16096 (N_16096,N_10463,N_12615);
nand U16097 (N_16097,N_12026,N_11932);
nand U16098 (N_16098,N_10635,N_14829);
or U16099 (N_16099,N_14372,N_11985);
and U16100 (N_16100,N_10251,N_12938);
or U16101 (N_16101,N_13364,N_14131);
xor U16102 (N_16102,N_11319,N_12213);
nand U16103 (N_16103,N_13947,N_10832);
nor U16104 (N_16104,N_12667,N_12763);
nor U16105 (N_16105,N_14188,N_13766);
nor U16106 (N_16106,N_14682,N_11861);
and U16107 (N_16107,N_11071,N_14217);
nand U16108 (N_16108,N_12221,N_14529);
nor U16109 (N_16109,N_12024,N_11457);
or U16110 (N_16110,N_14177,N_13810);
nor U16111 (N_16111,N_12781,N_14516);
xnor U16112 (N_16112,N_12758,N_11837);
xnor U16113 (N_16113,N_10033,N_13681);
xor U16114 (N_16114,N_10701,N_10761);
and U16115 (N_16115,N_12543,N_11800);
nor U16116 (N_16116,N_10122,N_13896);
or U16117 (N_16117,N_10448,N_12691);
nor U16118 (N_16118,N_13770,N_11743);
xor U16119 (N_16119,N_12935,N_12617);
xor U16120 (N_16120,N_11642,N_12065);
and U16121 (N_16121,N_11715,N_11914);
nor U16122 (N_16122,N_14295,N_12990);
nor U16123 (N_16123,N_13900,N_12374);
and U16124 (N_16124,N_13683,N_14142);
nor U16125 (N_16125,N_12482,N_13843);
nand U16126 (N_16126,N_14929,N_11895);
nor U16127 (N_16127,N_13685,N_13001);
nand U16128 (N_16128,N_13942,N_13223);
nor U16129 (N_16129,N_12245,N_11558);
nor U16130 (N_16130,N_14876,N_14289);
xor U16131 (N_16131,N_11858,N_12444);
xnor U16132 (N_16132,N_10345,N_10626);
and U16133 (N_16133,N_13684,N_10255);
nand U16134 (N_16134,N_14559,N_11121);
nor U16135 (N_16135,N_13893,N_11631);
xnor U16136 (N_16136,N_11470,N_14957);
xnor U16137 (N_16137,N_12621,N_14890);
nor U16138 (N_16138,N_12858,N_14106);
or U16139 (N_16139,N_10076,N_13861);
nor U16140 (N_16140,N_13967,N_14058);
or U16141 (N_16141,N_10219,N_14801);
nand U16142 (N_16142,N_10639,N_10687);
xor U16143 (N_16143,N_12476,N_12828);
nand U16144 (N_16144,N_10371,N_11964);
or U16145 (N_16145,N_11252,N_10995);
or U16146 (N_16146,N_11545,N_11937);
nor U16147 (N_16147,N_10333,N_14368);
nor U16148 (N_16148,N_12717,N_10704);
and U16149 (N_16149,N_11792,N_11569);
nand U16150 (N_16150,N_11680,N_11511);
nand U16151 (N_16151,N_13409,N_11287);
xnor U16152 (N_16152,N_13873,N_14511);
xnor U16153 (N_16153,N_14946,N_11608);
nand U16154 (N_16154,N_13842,N_13011);
nor U16155 (N_16155,N_11366,N_10527);
or U16156 (N_16156,N_10433,N_13740);
and U16157 (N_16157,N_12951,N_10018);
nor U16158 (N_16158,N_10577,N_10248);
nand U16159 (N_16159,N_10057,N_13883);
and U16160 (N_16160,N_14936,N_11044);
nand U16161 (N_16161,N_11494,N_10907);
nor U16162 (N_16162,N_12019,N_13369);
xor U16163 (N_16163,N_14649,N_14195);
and U16164 (N_16164,N_11180,N_12600);
nand U16165 (N_16165,N_10063,N_10539);
or U16166 (N_16166,N_10778,N_11417);
nor U16167 (N_16167,N_12462,N_13038);
xnor U16168 (N_16168,N_11026,N_12805);
nor U16169 (N_16169,N_12228,N_13163);
or U16170 (N_16170,N_11607,N_13241);
nor U16171 (N_16171,N_12511,N_11675);
xor U16172 (N_16172,N_14352,N_10449);
xnor U16173 (N_16173,N_11751,N_10518);
or U16174 (N_16174,N_10278,N_13849);
nor U16175 (N_16175,N_10000,N_12713);
xnor U16176 (N_16176,N_13914,N_13141);
or U16177 (N_16177,N_14231,N_14737);
or U16178 (N_16178,N_10628,N_10400);
and U16179 (N_16179,N_13868,N_12309);
xor U16180 (N_16180,N_10802,N_12319);
xnor U16181 (N_16181,N_11047,N_11003);
or U16182 (N_16182,N_12604,N_12034);
or U16183 (N_16183,N_10750,N_14964);
xnor U16184 (N_16184,N_13807,N_10901);
and U16185 (N_16185,N_11669,N_12558);
xnor U16186 (N_16186,N_11641,N_10509);
or U16187 (N_16187,N_10189,N_14413);
nor U16188 (N_16188,N_14464,N_10614);
or U16189 (N_16189,N_11662,N_11755);
and U16190 (N_16190,N_10570,N_11602);
or U16191 (N_16191,N_10151,N_13833);
nand U16192 (N_16192,N_10273,N_10294);
nor U16193 (N_16193,N_12743,N_10580);
or U16194 (N_16194,N_13687,N_14339);
nor U16195 (N_16195,N_14896,N_14234);
nand U16196 (N_16196,N_11111,N_10011);
and U16197 (N_16197,N_13073,N_11085);
nand U16198 (N_16198,N_11744,N_10458);
xor U16199 (N_16199,N_10897,N_13572);
or U16200 (N_16200,N_13417,N_10476);
and U16201 (N_16201,N_13670,N_13492);
nand U16202 (N_16202,N_14569,N_10705);
xnor U16203 (N_16203,N_12210,N_13088);
nand U16204 (N_16204,N_12280,N_10982);
and U16205 (N_16205,N_13071,N_14454);
or U16206 (N_16206,N_10637,N_13518);
xnor U16207 (N_16207,N_13795,N_10472);
or U16208 (N_16208,N_13777,N_12438);
or U16209 (N_16209,N_12683,N_14100);
or U16210 (N_16210,N_10030,N_11075);
xor U16211 (N_16211,N_12321,N_12829);
and U16212 (N_16212,N_12431,N_10986);
and U16213 (N_16213,N_10519,N_11532);
xnor U16214 (N_16214,N_13935,N_14842);
nor U16215 (N_16215,N_13026,N_13502);
nand U16216 (N_16216,N_10012,N_14294);
and U16217 (N_16217,N_12903,N_11125);
nand U16218 (N_16218,N_13252,N_11618);
xor U16219 (N_16219,N_10993,N_13134);
xnor U16220 (N_16220,N_13973,N_14210);
nor U16221 (N_16221,N_14179,N_14623);
xnor U16222 (N_16222,N_11664,N_10755);
xnor U16223 (N_16223,N_12859,N_13820);
or U16224 (N_16224,N_10892,N_12360);
or U16225 (N_16225,N_14388,N_13874);
nor U16226 (N_16226,N_11103,N_11307);
or U16227 (N_16227,N_14795,N_14489);
and U16228 (N_16228,N_13392,N_11981);
nor U16229 (N_16229,N_14273,N_13936);
and U16230 (N_16230,N_13784,N_12268);
nor U16231 (N_16231,N_14132,N_10804);
xnor U16232 (N_16232,N_11892,N_12121);
and U16233 (N_16233,N_12337,N_12182);
nand U16234 (N_16234,N_13575,N_13846);
nor U16235 (N_16235,N_10279,N_10207);
nor U16236 (N_16236,N_13864,N_13301);
nand U16237 (N_16237,N_11338,N_13937);
xor U16238 (N_16238,N_11701,N_13974);
nor U16239 (N_16239,N_14909,N_14517);
or U16240 (N_16240,N_10194,N_10681);
and U16241 (N_16241,N_12338,N_10782);
xnor U16242 (N_16242,N_11250,N_14631);
or U16243 (N_16243,N_10131,N_11251);
nand U16244 (N_16244,N_12960,N_13272);
nor U16245 (N_16245,N_12851,N_13344);
nand U16246 (N_16246,N_11860,N_12515);
and U16247 (N_16247,N_13523,N_11102);
nor U16248 (N_16248,N_11518,N_13441);
xnor U16249 (N_16249,N_14852,N_10587);
nand U16250 (N_16250,N_14921,N_11127);
nor U16251 (N_16251,N_11629,N_14031);
nand U16252 (N_16252,N_11305,N_11150);
xnor U16253 (N_16253,N_13312,N_12505);
nand U16254 (N_16254,N_14922,N_10152);
xnor U16255 (N_16255,N_13885,N_13603);
nor U16256 (N_16256,N_13431,N_10461);
nand U16257 (N_16257,N_13671,N_14491);
and U16258 (N_16258,N_10949,N_14169);
nand U16259 (N_16259,N_10754,N_13329);
xnor U16260 (N_16260,N_10648,N_10510);
nor U16261 (N_16261,N_14726,N_13258);
xor U16262 (N_16262,N_12902,N_12983);
or U16263 (N_16263,N_10080,N_14747);
nand U16264 (N_16264,N_11563,N_11007);
xnor U16265 (N_16265,N_10280,N_10346);
or U16266 (N_16266,N_14186,N_14777);
nor U16267 (N_16267,N_14309,N_14831);
and U16268 (N_16268,N_11767,N_11303);
or U16269 (N_16269,N_13352,N_11151);
xor U16270 (N_16270,N_13148,N_11365);
nand U16271 (N_16271,N_13004,N_12344);
nand U16272 (N_16272,N_13159,N_14752);
nor U16273 (N_16273,N_11216,N_11080);
nor U16274 (N_16274,N_14676,N_14730);
nand U16275 (N_16275,N_14324,N_10785);
nand U16276 (N_16276,N_10709,N_12254);
nor U16277 (N_16277,N_10290,N_13238);
nor U16278 (N_16278,N_14395,N_12165);
and U16279 (N_16279,N_11027,N_10029);
or U16280 (N_16280,N_14263,N_14415);
and U16281 (N_16281,N_10034,N_14471);
nand U16282 (N_16282,N_11351,N_14200);
and U16283 (N_16283,N_14126,N_14344);
and U16284 (N_16284,N_14616,N_12930);
xnor U16285 (N_16285,N_11665,N_10638);
nand U16286 (N_16286,N_11898,N_14432);
or U16287 (N_16287,N_13396,N_14004);
xnor U16288 (N_16288,N_10889,N_11107);
xnor U16289 (N_16289,N_10552,N_11634);
xor U16290 (N_16290,N_12562,N_12229);
nand U16291 (N_16291,N_11766,N_12985);
xnor U16292 (N_16292,N_13963,N_11962);
or U16293 (N_16293,N_10116,N_12861);
nand U16294 (N_16294,N_12434,N_14181);
xor U16295 (N_16295,N_10364,N_11442);
xnor U16296 (N_16296,N_11584,N_14647);
nor U16297 (N_16297,N_10508,N_10160);
or U16298 (N_16298,N_12678,N_10835);
or U16299 (N_16299,N_13506,N_10017);
nor U16300 (N_16300,N_12346,N_12102);
and U16301 (N_16301,N_10436,N_14865);
nand U16302 (N_16302,N_11052,N_14085);
and U16303 (N_16303,N_11057,N_12220);
nor U16304 (N_16304,N_14996,N_13311);
nand U16305 (N_16305,N_13816,N_11153);
or U16306 (N_16306,N_11648,N_12039);
and U16307 (N_16307,N_14960,N_11454);
or U16308 (N_16308,N_12164,N_11491);
nor U16309 (N_16309,N_14720,N_13337);
nand U16310 (N_16310,N_10019,N_13604);
xor U16311 (N_16311,N_12725,N_12982);
nor U16312 (N_16312,N_13207,N_13145);
nor U16313 (N_16313,N_12794,N_13663);
nand U16314 (N_16314,N_14648,N_12157);
and U16315 (N_16315,N_14455,N_12105);
or U16316 (N_16316,N_14392,N_14453);
and U16317 (N_16317,N_13093,N_11534);
xor U16318 (N_16318,N_10347,N_13760);
xnor U16319 (N_16319,N_12645,N_14070);
nand U16320 (N_16320,N_12015,N_10879);
nand U16321 (N_16321,N_14981,N_14916);
and U16322 (N_16322,N_14881,N_10999);
xor U16323 (N_16323,N_13624,N_13496);
nand U16324 (N_16324,N_13698,N_13432);
and U16325 (N_16325,N_13224,N_10272);
xor U16326 (N_16326,N_11688,N_10717);
nor U16327 (N_16327,N_14851,N_10863);
and U16328 (N_16328,N_13416,N_12083);
xor U16329 (N_16329,N_11050,N_14999);
and U16330 (N_16330,N_10765,N_14699);
nand U16331 (N_16331,N_11922,N_12402);
nor U16332 (N_16332,N_12363,N_14989);
nor U16333 (N_16333,N_13696,N_13008);
and U16334 (N_16334,N_13641,N_13166);
nand U16335 (N_16335,N_10344,N_14299);
or U16336 (N_16336,N_12031,N_13812);
or U16337 (N_16337,N_12122,N_10586);
xor U16338 (N_16338,N_11727,N_11555);
and U16339 (N_16339,N_14712,N_10851);
nor U16340 (N_16340,N_12762,N_13673);
and U16341 (N_16341,N_10679,N_10068);
nand U16342 (N_16342,N_12284,N_11574);
nor U16343 (N_16343,N_12561,N_14099);
xnor U16344 (N_16344,N_12305,N_10601);
and U16345 (N_16345,N_10388,N_10834);
nor U16346 (N_16346,N_11928,N_13447);
nor U16347 (N_16347,N_14830,N_10197);
nor U16348 (N_16348,N_14045,N_14802);
and U16349 (N_16349,N_10820,N_13361);
and U16350 (N_16350,N_13705,N_13099);
or U16351 (N_16351,N_12636,N_11048);
xnor U16352 (N_16352,N_14422,N_14949);
or U16353 (N_16353,N_12283,N_14400);
nand U16354 (N_16354,N_14738,N_12336);
nand U16355 (N_16355,N_14498,N_12099);
xnor U16356 (N_16356,N_13273,N_11053);
nor U16357 (N_16357,N_14414,N_13847);
and U16358 (N_16358,N_14900,N_14760);
or U16359 (N_16359,N_13385,N_14104);
or U16360 (N_16360,N_11576,N_12179);
and U16361 (N_16361,N_11708,N_10351);
nor U16362 (N_16362,N_14406,N_13288);
nand U16363 (N_16363,N_11276,N_14693);
and U16364 (N_16364,N_12987,N_13132);
xnor U16365 (N_16365,N_14786,N_10719);
or U16366 (N_16366,N_11477,N_13039);
and U16367 (N_16367,N_12163,N_10980);
or U16368 (N_16368,N_10471,N_13454);
xor U16369 (N_16369,N_10520,N_12765);
nor U16370 (N_16370,N_12361,N_14194);
nor U16371 (N_16371,N_14424,N_14460);
and U16372 (N_16372,N_11259,N_11432);
nor U16373 (N_16373,N_12270,N_13085);
and U16374 (N_16374,N_13619,N_11291);
or U16375 (N_16375,N_10003,N_13908);
nand U16376 (N_16376,N_13659,N_13161);
and U16377 (N_16377,N_13291,N_14011);
or U16378 (N_16378,N_14626,N_14913);
nor U16379 (N_16379,N_14018,N_10175);
nand U16380 (N_16380,N_11400,N_10234);
xor U16381 (N_16381,N_11181,N_13449);
nand U16382 (N_16382,N_13949,N_13546);
or U16383 (N_16383,N_12359,N_13899);
nand U16384 (N_16384,N_10673,N_13185);
and U16385 (N_16385,N_11339,N_12521);
xnor U16386 (N_16386,N_12107,N_13098);
nand U16387 (N_16387,N_12298,N_12612);
nor U16388 (N_16388,N_12817,N_12457);
xnor U16389 (N_16389,N_12800,N_12442);
nor U16390 (N_16390,N_10584,N_13867);
xnor U16391 (N_16391,N_11006,N_11515);
nor U16392 (N_16392,N_14924,N_14447);
or U16393 (N_16393,N_14499,N_14965);
or U16394 (N_16394,N_12178,N_12287);
and U16395 (N_16395,N_14117,N_13330);
and U16396 (N_16396,N_14583,N_13018);
nand U16397 (N_16397,N_14086,N_12224);
or U16398 (N_16398,N_12714,N_14064);
nor U16399 (N_16399,N_14440,N_13612);
nor U16400 (N_16400,N_12540,N_12132);
xnor U16401 (N_16401,N_10906,N_13862);
nor U16402 (N_16402,N_12623,N_10486);
and U16403 (N_16403,N_11786,N_12441);
xnor U16404 (N_16404,N_13182,N_10389);
and U16405 (N_16405,N_14080,N_14361);
nor U16406 (N_16406,N_12943,N_12735);
and U16407 (N_16407,N_10753,N_10797);
or U16408 (N_16408,N_11822,N_13574);
xnor U16409 (N_16409,N_13542,N_14129);
nor U16410 (N_16410,N_12330,N_13746);
or U16411 (N_16411,N_13595,N_14257);
xnor U16412 (N_16412,N_13653,N_10720);
nor U16413 (N_16413,N_11630,N_12898);
and U16414 (N_16414,N_14101,N_12825);
and U16415 (N_16415,N_11094,N_12660);
or U16416 (N_16416,N_14552,N_11430);
xor U16417 (N_16417,N_10887,N_11829);
nor U16418 (N_16418,N_13012,N_11249);
and U16419 (N_16419,N_13837,N_12686);
nor U16420 (N_16420,N_13573,N_13226);
and U16421 (N_16421,N_10262,N_12917);
xor U16422 (N_16422,N_10469,N_14821);
xnor U16423 (N_16423,N_11978,N_13313);
xnor U16424 (N_16424,N_11955,N_11862);
and U16425 (N_16425,N_14843,N_11604);
and U16426 (N_16426,N_11723,N_12991);
nor U16427 (N_16427,N_12196,N_11445);
or U16428 (N_16428,N_10634,N_10265);
or U16429 (N_16429,N_14966,N_13310);
or U16430 (N_16430,N_13298,N_10368);
xnor U16431 (N_16431,N_14908,N_14271);
and U16432 (N_16432,N_11714,N_12931);
or U16433 (N_16433,N_13729,N_11656);
nor U16434 (N_16434,N_12940,N_13623);
and U16435 (N_16435,N_11951,N_14919);
xnor U16436 (N_16436,N_10936,N_13541);
nor U16437 (N_16437,N_14557,N_11804);
and U16438 (N_16438,N_12347,N_11483);
nand U16439 (N_16439,N_10908,N_10591);
nand U16440 (N_16440,N_11158,N_12634);
or U16441 (N_16441,N_10934,N_11143);
nand U16442 (N_16442,N_12830,N_13650);
or U16443 (N_16443,N_12579,N_13160);
and U16444 (N_16444,N_11194,N_13726);
nand U16445 (N_16445,N_14665,N_14269);
nand U16446 (N_16446,N_12173,N_10301);
or U16447 (N_16447,N_11772,N_14524);
nand U16448 (N_16448,N_11014,N_11100);
nand U16449 (N_16449,N_11746,N_14721);
or U16450 (N_16450,N_14568,N_14043);
and U16451 (N_16451,N_10548,N_14355);
and U16452 (N_16452,N_14150,N_14140);
nand U16453 (N_16453,N_14615,N_11610);
and U16454 (N_16454,N_13836,N_12408);
or U16455 (N_16455,N_13895,N_10763);
or U16456 (N_16456,N_12843,N_14940);
nor U16457 (N_16457,N_11311,N_12302);
nand U16458 (N_16458,N_13987,N_12687);
xnor U16459 (N_16459,N_14003,N_10191);
or U16460 (N_16460,N_11383,N_14325);
and U16461 (N_16461,N_14014,N_10376);
xor U16462 (N_16462,N_14607,N_11724);
nand U16463 (N_16463,N_13608,N_12016);
and U16464 (N_16464,N_12427,N_14362);
nand U16465 (N_16465,N_11472,N_12448);
nand U16466 (N_16466,N_13357,N_10671);
nor U16467 (N_16467,N_13219,N_10583);
nand U16468 (N_16468,N_11464,N_14666);
or U16469 (N_16469,N_10138,N_10884);
and U16470 (N_16470,N_10850,N_12194);
nand U16471 (N_16471,N_12306,N_13890);
xor U16472 (N_16472,N_10375,N_14776);
nand U16473 (N_16473,N_11035,N_13805);
or U16474 (N_16474,N_14785,N_10952);
nand U16475 (N_16475,N_13256,N_12139);
and U16476 (N_16476,N_13537,N_11112);
and U16477 (N_16477,N_12326,N_10924);
and U16478 (N_16478,N_14151,N_12045);
nand U16479 (N_16479,N_14236,N_10407);
and U16480 (N_16480,N_11331,N_11414);
xor U16481 (N_16481,N_10799,N_13622);
and U16482 (N_16482,N_11218,N_12551);
nand U16483 (N_16483,N_13442,N_13175);
nand U16484 (N_16484,N_13561,N_11948);
xnor U16485 (N_16485,N_13680,N_11748);
xnor U16486 (N_16486,N_13912,N_14239);
xor U16487 (N_16487,N_13562,N_10981);
xnor U16488 (N_16488,N_11295,N_13194);
and U16489 (N_16489,N_11635,N_12109);
nor U16490 (N_16490,N_11340,N_13097);
nand U16491 (N_16491,N_10613,N_12726);
or U16492 (N_16492,N_13931,N_10170);
nand U16493 (N_16493,N_13601,N_11046);
xnor U16494 (N_16494,N_13706,N_14961);
and U16495 (N_16495,N_11789,N_13181);
xor U16496 (N_16496,N_14298,N_13117);
or U16497 (N_16497,N_11227,N_12666);
xnor U16498 (N_16498,N_12909,N_12358);
or U16499 (N_16499,N_10838,N_12108);
or U16500 (N_16500,N_11940,N_13087);
xor U16501 (N_16501,N_12622,N_13381);
nand U16502 (N_16502,N_11043,N_12831);
nor U16503 (N_16503,N_12994,N_14544);
or U16504 (N_16504,N_10780,N_12862);
and U16505 (N_16505,N_11015,N_13584);
or U16506 (N_16506,N_11299,N_13813);
nor U16507 (N_16507,N_13811,N_13723);
or U16508 (N_16508,N_13656,N_12959);
nor U16509 (N_16509,N_13068,N_13051);
nor U16510 (N_16510,N_12810,N_12673);
nand U16511 (N_16511,N_11209,N_13101);
nand U16512 (N_16512,N_11885,N_13489);
or U16513 (N_16513,N_10677,N_13365);
nand U16514 (N_16514,N_12404,N_11078);
or U16515 (N_16515,N_12468,N_10215);
or U16516 (N_16516,N_10865,N_11431);
nor U16517 (N_16517,N_11420,N_13996);
xnor U16518 (N_16518,N_12952,N_12595);
xnor U16519 (N_16519,N_13835,N_13728);
or U16520 (N_16520,N_11651,N_14798);
xor U16521 (N_16521,N_11661,N_10491);
xor U16522 (N_16522,N_13336,N_10490);
or U16523 (N_16523,N_14456,N_13814);
and U16524 (N_16524,N_12014,N_10883);
and U16525 (N_16525,N_10868,N_13142);
or U16526 (N_16526,N_10201,N_12469);
xnor U16527 (N_16527,N_14479,N_10568);
and U16528 (N_16528,N_12060,N_13856);
xor U16529 (N_16529,N_11037,N_10445);
nor U16530 (N_16530,N_14575,N_13066);
or U16531 (N_16531,N_11369,N_14428);
nand U16532 (N_16532,N_13100,N_10525);
nor U16533 (N_16533,N_10036,N_11742);
and U16534 (N_16534,N_11234,N_10956);
xor U16535 (N_16535,N_12090,N_11956);
xor U16536 (N_16536,N_10240,N_14327);
nor U16537 (N_16537,N_12212,N_10496);
nand U16538 (N_16538,N_10334,N_10196);
and U16539 (N_16539,N_14555,N_14088);
and U16540 (N_16540,N_11826,N_13774);
or U16541 (N_16541,N_11841,N_12529);
xor U16542 (N_16542,N_10304,N_11213);
and U16543 (N_16543,N_14709,N_12032);
nor U16544 (N_16544,N_14710,N_10745);
xor U16545 (N_16545,N_12995,N_13373);
or U16546 (N_16546,N_12103,N_13718);
nor U16547 (N_16547,N_10062,N_14123);
or U16548 (N_16548,N_14596,N_12999);
and U16549 (N_16549,N_13065,N_12616);
nand U16550 (N_16550,N_14103,N_10382);
xnor U16551 (N_16551,N_10105,N_13005);
xor U16552 (N_16552,N_12170,N_12549);
xor U16553 (N_16553,N_14404,N_11391);
nand U16554 (N_16554,N_13880,N_12569);
or U16555 (N_16555,N_14547,N_11156);
xor U16556 (N_16556,N_14035,N_14599);
and U16557 (N_16557,N_14466,N_10972);
nand U16558 (N_16558,N_11258,N_13560);
nor U16559 (N_16559,N_12802,N_11309);
xnor U16560 (N_16560,N_14679,N_13579);
or U16561 (N_16561,N_12197,N_12413);
xor U16562 (N_16562,N_11991,N_13172);
and U16563 (N_16563,N_10101,N_11681);
or U16564 (N_16564,N_14576,N_11243);
and U16565 (N_16565,N_11349,N_12564);
and U16566 (N_16566,N_10397,N_10932);
or U16567 (N_16567,N_11419,N_13858);
xnor U16568 (N_16568,N_12130,N_10723);
and U16569 (N_16569,N_13002,N_11484);
nand U16570 (N_16570,N_14558,N_14203);
or U16571 (N_16571,N_14567,N_13976);
nand U16572 (N_16572,N_11460,N_14620);
and U16573 (N_16573,N_14658,N_12809);
and U16574 (N_16574,N_10230,N_12545);
nor U16575 (N_16575,N_12801,N_14175);
nand U16576 (N_16576,N_10994,N_11318);
nor U16577 (N_16577,N_10172,N_12420);
nor U16578 (N_16578,N_14836,N_13428);
xor U16579 (N_16579,N_11013,N_13563);
xor U16580 (N_16580,N_12475,N_12123);
nor U16581 (N_16581,N_14482,N_13094);
nor U16582 (N_16582,N_14076,N_11122);
and U16583 (N_16583,N_10087,N_12925);
nand U16584 (N_16584,N_12023,N_13674);
and U16585 (N_16585,N_14020,N_11060);
nor U16586 (N_16586,N_11069,N_13179);
and U16587 (N_16587,N_14612,N_12554);
nand U16588 (N_16588,N_12390,N_11162);
xnor U16589 (N_16589,N_14560,N_12141);
and U16590 (N_16590,N_13640,N_11481);
and U16591 (N_16591,N_11973,N_12078);
nor U16592 (N_16592,N_11830,N_13818);
nand U16593 (N_16593,N_10398,N_14827);
or U16594 (N_16594,N_14353,N_11168);
xor U16595 (N_16595,N_13042,N_12161);
xor U16596 (N_16596,N_10483,N_10938);
nand U16597 (N_16597,N_12962,N_13395);
xor U16598 (N_16598,N_12041,N_11741);
or U16599 (N_16599,N_14010,N_12285);
or U16600 (N_16600,N_10911,N_11633);
and U16601 (N_16601,N_10437,N_14127);
xor U16602 (N_16602,N_14696,N_14416);
xnor U16603 (N_16603,N_11936,N_10439);
nand U16604 (N_16604,N_13823,N_14571);
or U16605 (N_16605,N_10258,N_12345);
nor U16606 (N_16606,N_14619,N_11597);
nor U16607 (N_16607,N_13137,N_13371);
and U16608 (N_16608,N_13028,N_14292);
nor U16609 (N_16609,N_10569,N_12649);
xnor U16610 (N_16610,N_11559,N_11275);
and U16611 (N_16611,N_13410,N_13930);
xnor U16612 (N_16612,N_14835,N_14444);
or U16613 (N_16613,N_10313,N_10025);
or U16614 (N_16614,N_12156,N_11324);
nand U16615 (N_16615,N_11058,N_14246);
xnor U16616 (N_16616,N_14019,N_13195);
or U16617 (N_16617,N_12047,N_14533);
nand U16618 (N_16618,N_12733,N_12607);
xor U16619 (N_16619,N_12749,N_10184);
nor U16620 (N_16620,N_12449,N_10058);
or U16621 (N_16621,N_13009,N_12640);
nor U16622 (N_16622,N_12526,N_14907);
nand U16623 (N_16623,N_11617,N_10683);
nor U16624 (N_16624,N_13522,N_13907);
nor U16625 (N_16625,N_14407,N_12557);
nor U16626 (N_16626,N_11782,N_10946);
xor U16627 (N_16627,N_10129,N_10108);
nand U16628 (N_16628,N_10427,N_12128);
and U16629 (N_16629,N_12841,N_13375);
xor U16630 (N_16630,N_13761,N_14915);
nor U16631 (N_16631,N_14125,N_13629);
or U16632 (N_16632,N_11686,N_12814);
or U16633 (N_16633,N_10121,N_10203);
and U16634 (N_16634,N_12452,N_14254);
xnor U16635 (N_16635,N_10318,N_14548);
or U16636 (N_16636,N_10854,N_12362);
xnor U16637 (N_16637,N_14816,N_11357);
nor U16638 (N_16638,N_14657,N_10052);
or U16639 (N_16639,N_10599,N_14780);
xor U16640 (N_16640,N_10598,N_13458);
nor U16641 (N_16641,N_12195,N_11886);
and U16642 (N_16642,N_12587,N_11224);
nand U16643 (N_16643,N_13636,N_11666);
or U16644 (N_16644,N_12603,N_12581);
nor U16645 (N_16645,N_12380,N_10142);
xnor U16646 (N_16646,N_12186,N_12971);
nor U16647 (N_16647,N_11705,N_12079);
xor U16648 (N_16648,N_12479,N_11986);
and U16649 (N_16649,N_13759,N_12536);
nor U16650 (N_16650,N_10054,N_11810);
or U16651 (N_16651,N_11643,N_11390);
nor U16652 (N_16652,N_12734,N_13957);
nand U16653 (N_16653,N_12159,N_10777);
xnor U16654 (N_16654,N_13057,N_14624);
xnor U16655 (N_16655,N_10457,N_10438);
xnor U16656 (N_16656,N_11302,N_11799);
xnor U16657 (N_16657,N_10504,N_12998);
nand U16658 (N_16658,N_14874,N_12585);
and U16659 (N_16659,N_10042,N_13267);
and U16660 (N_16660,N_13083,N_14617);
and U16661 (N_16661,N_14008,N_14762);
or U16662 (N_16662,N_12313,N_10451);
nand U16663 (N_16663,N_12839,N_11780);
xor U16664 (N_16664,N_11499,N_14526);
and U16665 (N_16665,N_12437,N_13303);
and U16666 (N_16666,N_13096,N_12394);
nor U16667 (N_16667,N_14771,N_12533);
xor U16668 (N_16668,N_14025,N_12439);
xnor U16669 (N_16669,N_12046,N_10231);
and U16670 (N_16670,N_10663,N_11774);
or U16671 (N_16671,N_11889,N_10807);
or U16672 (N_16672,N_13150,N_11004);
or U16673 (N_16673,N_11380,N_11819);
xnor U16674 (N_16674,N_13067,N_10984);
xor U16675 (N_16675,N_10001,N_12657);
xor U16676 (N_16676,N_13037,N_12372);
and U16677 (N_16677,N_13322,N_14774);
or U16678 (N_16678,N_13127,N_12088);
xnor U16679 (N_16679,N_13003,N_11877);
nor U16680 (N_16680,N_13513,N_13386);
and U16681 (N_16681,N_10918,N_13697);
nand U16682 (N_16682,N_12635,N_12296);
xnor U16683 (N_16683,N_12495,N_11372);
and U16684 (N_16684,N_13898,N_11360);
xor U16685 (N_16685,N_13672,N_13977);
xor U16686 (N_16686,N_12203,N_14590);
nand U16687 (N_16687,N_11783,N_10955);
nand U16688 (N_16688,N_13749,N_14530);
or U16689 (N_16689,N_10008,N_12993);
xnor U16690 (N_16690,N_10592,N_10059);
nor U16691 (N_16691,N_13505,N_14311);
nor U16692 (N_16692,N_11451,N_12682);
xnor U16693 (N_16693,N_14783,N_10658);
nand U16694 (N_16694,N_14153,N_12632);
nor U16695 (N_16695,N_13756,N_14038);
nor U16696 (N_16696,N_11189,N_12710);
and U16697 (N_16697,N_10727,N_10291);
nor U16698 (N_16698,N_14147,N_10894);
and U16699 (N_16699,N_13701,N_14016);
and U16700 (N_16700,N_13423,N_12454);
or U16701 (N_16701,N_12879,N_13532);
nand U16702 (N_16702,N_11647,N_11996);
or U16703 (N_16703,N_10645,N_13173);
and U16704 (N_16704,N_14009,N_10115);
xnor U16705 (N_16705,N_13325,N_11314);
nand U16706 (N_16706,N_10487,N_12654);
and U16707 (N_16707,N_12664,N_12050);
and U16708 (N_16708,N_11753,N_13709);
nor U16709 (N_16709,N_11011,N_12202);
xor U16710 (N_16710,N_14613,N_13420);
xor U16711 (N_16711,N_10112,N_10310);
xor U16712 (N_16712,N_11813,N_14184);
xor U16713 (N_16713,N_13776,N_12834);
nand U16714 (N_16714,N_11316,N_12116);
and U16715 (N_16715,N_12250,N_13994);
nand U16716 (N_16716,N_14991,N_12916);
xor U16717 (N_16717,N_13107,N_11710);
nand U16718 (N_16718,N_14399,N_10522);
nor U16719 (N_16719,N_14853,N_12754);
or U16720 (N_16720,N_13941,N_13720);
nand U16721 (N_16721,N_10158,N_10355);
or U16722 (N_16722,N_13403,N_13852);
xnor U16723 (N_16723,N_10845,N_11712);
nand U16724 (N_16724,N_12473,N_11240);
or U16725 (N_16725,N_12312,N_10676);
xor U16726 (N_16726,N_11412,N_11000);
nor U16727 (N_16727,N_14973,N_10748);
xnor U16728 (N_16728,N_10585,N_11918);
nor U16729 (N_16729,N_13711,N_14715);
and U16730 (N_16730,N_13405,N_10181);
nor U16731 (N_16731,N_10435,N_12459);
and U16732 (N_16732,N_11281,N_13348);
nand U16733 (N_16733,N_12144,N_12845);
nor U16734 (N_16734,N_14740,N_14586);
nand U16735 (N_16735,N_14954,N_14604);
nor U16736 (N_16736,N_14718,N_10277);
and U16737 (N_16737,N_13950,N_12739);
nand U16738 (N_16738,N_10633,N_10722);
or U16739 (N_16739,N_13323,N_11990);
xor U16740 (N_16740,N_14402,N_13621);
nand U16741 (N_16741,N_12875,N_14633);
or U16742 (N_16742,N_11387,N_12232);
xnor U16743 (N_16743,N_10328,N_12768);
xnor U16744 (N_16744,N_14621,N_12548);
nor U16745 (N_16745,N_14920,N_11636);
and U16746 (N_16746,N_12870,N_10815);
nand U16747 (N_16747,N_13198,N_13981);
or U16748 (N_16748,N_14893,N_11135);
nor U16749 (N_16749,N_10991,N_14792);
or U16750 (N_16750,N_13480,N_14956);
or U16751 (N_16751,N_11668,N_12707);
nor U16752 (N_16752,N_12211,N_12307);
nand U16753 (N_16753,N_12009,N_11847);
or U16754 (N_16754,N_11352,N_13783);
xor U16755 (N_16755,N_10516,N_11808);
nand U16756 (N_16756,N_10816,N_10092);
and U16757 (N_16757,N_14980,N_14161);
xor U16758 (N_16758,N_10039,N_10506);
xnor U16759 (N_16759,N_12407,N_11926);
nor U16760 (N_16760,N_10465,N_14734);
nand U16761 (N_16761,N_11578,N_10253);
and U16762 (N_16762,N_12492,N_12923);
xor U16763 (N_16763,N_14039,N_11223);
or U16764 (N_16764,N_14277,N_12487);
nor U16765 (N_16765,N_14196,N_10099);
or U16766 (N_16766,N_13526,N_14826);
or U16767 (N_16767,N_14275,N_10667);
and U16768 (N_16768,N_11887,N_13809);
or U16769 (N_16769,N_14189,N_12063);
nand U16770 (N_16770,N_10084,N_13876);
xnor U16771 (N_16771,N_11405,N_13324);
nor U16772 (N_16772,N_13927,N_10692);
nor U16773 (N_16773,N_10735,N_14817);
or U16774 (N_16774,N_10880,N_14347);
nor U16775 (N_16775,N_14611,N_10666);
and U16776 (N_16776,N_13180,N_13360);
nand U16777 (N_16777,N_14380,N_14223);
xor U16778 (N_16778,N_11079,N_12301);
xor U16779 (N_16779,N_10951,N_10556);
or U16780 (N_16780,N_14041,N_14037);
or U16781 (N_16781,N_11859,N_14199);
nand U16782 (N_16782,N_13055,N_10454);
or U16783 (N_16783,N_14145,N_10558);
nand U16784 (N_16784,N_12680,N_14159);
and U16785 (N_16785,N_11090,N_11809);
nand U16786 (N_16786,N_13730,N_12661);
and U16787 (N_16787,N_12932,N_13969);
nand U16788 (N_16788,N_14833,N_10831);
or U16789 (N_16789,N_13547,N_13236);
nand U16790 (N_16790,N_14618,N_11677);
or U16791 (N_16791,N_12077,N_10674);
nand U16792 (N_16792,N_13888,N_10023);
nand U16793 (N_16793,N_11852,N_13013);
and U16794 (N_16794,N_13383,N_13157);
nand U16795 (N_16795,N_14034,N_10732);
or U16796 (N_16796,N_14205,N_14659);
nor U16797 (N_16797,N_10651,N_10254);
or U16798 (N_16798,N_12883,N_14951);
nand U16799 (N_16799,N_14519,N_10381);
nor U16800 (N_16800,N_11831,N_12876);
and U16801 (N_16801,N_11707,N_11900);
or U16802 (N_16802,N_12741,N_13459);
or U16803 (N_16803,N_12867,N_11337);
nand U16804 (N_16804,N_13915,N_11812);
nor U16805 (N_16805,N_12129,N_10386);
xor U16806 (N_16806,N_12158,N_13169);
nand U16807 (N_16807,N_12275,N_13865);
or U16808 (N_16808,N_10594,N_11401);
nor U16809 (N_16809,N_10326,N_14446);
and U16810 (N_16810,N_11308,N_13564);
xnor U16811 (N_16811,N_11320,N_10156);
nor U16812 (N_16812,N_11687,N_13295);
nor U16813 (N_16813,N_11310,N_11394);
nor U16814 (N_16814,N_11214,N_11983);
xor U16815 (N_16815,N_12596,N_13741);
nand U16816 (N_16816,N_11802,N_14770);
and U16817 (N_16817,N_10760,N_12507);
and U16818 (N_16818,N_12042,N_12522);
xnor U16819 (N_16819,N_10282,N_14260);
or U16820 (N_16820,N_13902,N_12409);
and U16821 (N_16821,N_12823,N_12892);
or U16822 (N_16822,N_11086,N_12335);
xnor U16823 (N_16823,N_11645,N_12385);
xor U16824 (N_16824,N_12365,N_11562);
xor U16825 (N_16825,N_10409,N_11358);
nand U16826 (N_16826,N_12225,N_13178);
nor U16827 (N_16827,N_10833,N_11034);
and U16828 (N_16828,N_14049,N_12084);
or U16829 (N_16829,N_13130,N_13307);
nor U16830 (N_16830,N_13339,N_11192);
xor U16831 (N_16831,N_11654,N_10315);
nand U16832 (N_16832,N_14870,N_12393);
nand U16833 (N_16833,N_10322,N_13716);
nand U16834 (N_16834,N_12857,N_10242);
or U16835 (N_16835,N_11495,N_10235);
or U16836 (N_16836,N_10566,N_11523);
nor U16837 (N_16837,N_14154,N_14694);
xor U16838 (N_16838,N_13384,N_14554);
nor U16839 (N_16839,N_10818,N_11806);
xnor U16840 (N_16840,N_10374,N_12185);
nand U16841 (N_16841,N_11775,N_13251);
or U16842 (N_16842,N_10113,N_12231);
and U16843 (N_16843,N_12777,N_12140);
nand U16844 (N_16844,N_12237,N_12460);
and U16845 (N_16845,N_13667,N_13821);
nand U16846 (N_16846,N_14601,N_12772);
or U16847 (N_16847,N_11527,N_11486);
nand U16848 (N_16848,N_12997,N_13177);
or U16849 (N_16849,N_11298,N_10990);
xnor U16850 (N_16850,N_10945,N_11984);
nor U16851 (N_16851,N_14914,N_11839);
xnor U16852 (N_16852,N_14119,N_13108);
or U16853 (N_16853,N_10070,N_12816);
xor U16854 (N_16854,N_11794,N_11160);
xnor U16855 (N_16855,N_12582,N_12389);
nand U16856 (N_16856,N_12592,N_10312);
nor U16857 (N_16857,N_13782,N_11833);
nor U16858 (N_16858,N_13217,N_14255);
nand U16859 (N_16859,N_11593,N_10544);
xor U16860 (N_16860,N_14858,N_13205);
or U16861 (N_16861,N_10874,N_14278);
nand U16862 (N_16862,N_12677,N_13613);
xor U16863 (N_16863,N_12151,N_10128);
nor U16864 (N_16864,N_14518,N_13370);
and U16865 (N_16865,N_13739,N_13614);
and U16866 (N_16866,N_14562,N_11201);
xor U16867 (N_16867,N_14265,N_12120);
or U16868 (N_16868,N_10819,N_11199);
nand U16869 (N_16869,N_10752,N_12978);
nor U16870 (N_16870,N_11468,N_10222);
nor U16871 (N_16871,N_13208,N_11328);
and U16872 (N_16872,N_12638,N_11953);
nor U16873 (N_16873,N_12773,N_12864);
xor U16874 (N_16874,N_10137,N_11894);
xnor U16875 (N_16875,N_13658,N_10256);
xor U16876 (N_16876,N_14042,N_14985);
nor U16877 (N_16877,N_10844,N_13675);
nor U16878 (N_16878,N_13287,N_12948);
nand U16879 (N_16879,N_11924,N_12866);
nor U16880 (N_16880,N_12247,N_12594);
nand U16881 (N_16881,N_12152,N_14654);
or U16882 (N_16882,N_14427,N_11535);
and U16883 (N_16883,N_10578,N_11095);
xnor U16884 (N_16884,N_13566,N_13882);
and U16885 (N_16885,N_11306,N_13455);
nor U16886 (N_16886,N_12244,N_10856);
or U16887 (N_16887,N_12396,N_10617);
nand U16888 (N_16888,N_12905,N_14585);
or U16889 (N_16889,N_13517,N_12445);
nand U16890 (N_16890,N_14507,N_10157);
nand U16891 (N_16891,N_13870,N_14753);
nor U16892 (N_16892,N_14307,N_12628);
nand U16893 (N_16893,N_10898,N_11798);
nand U16894 (N_16894,N_14879,N_14122);
nand U16895 (N_16895,N_13358,N_13289);
or U16896 (N_16896,N_10284,N_12508);
nor U16897 (N_16897,N_12827,N_13269);
or U16898 (N_16898,N_13894,N_13424);
xnor U16899 (N_16899,N_13089,N_12888);
xnor U16900 (N_16900,N_12659,N_11051);
nor U16901 (N_16901,N_11694,N_11612);
and U16902 (N_16902,N_10190,N_13154);
and U16903 (N_16903,N_12570,N_10199);
and U16904 (N_16904,N_13245,N_12789);
or U16905 (N_16905,N_11211,N_10893);
and U16906 (N_16906,N_10715,N_11738);
nor U16907 (N_16907,N_10467,N_11049);
nor U16908 (N_16908,N_10317,N_12104);
and U16909 (N_16909,N_12366,N_10072);
and U16910 (N_16910,N_14799,N_13633);
nand U16911 (N_16911,N_14577,N_14643);
nor U16912 (N_16912,N_13857,N_10664);
xnor U16913 (N_16913,N_14044,N_13407);
xnor U16914 (N_16914,N_12979,N_12610);
and U16915 (N_16915,N_10526,N_12544);
and U16916 (N_16916,N_14933,N_12766);
and U16917 (N_16917,N_11466,N_14713);
nor U16918 (N_16918,N_12670,N_11315);
nand U16919 (N_16919,N_10608,N_11395);
nand U16920 (N_16920,N_14433,N_13152);
or U16921 (N_16921,N_14069,N_14366);
xor U16922 (N_16922,N_14093,N_14250);
and U16923 (N_16923,N_12945,N_14722);
or U16924 (N_16924,N_11711,N_11480);
and U16925 (N_16925,N_13607,N_13570);
nand U16926 (N_16926,N_13909,N_13457);
xnor U16927 (N_16927,N_11716,N_13583);
xnor U16928 (N_16928,N_11184,N_14947);
xnor U16929 (N_16929,N_11652,N_11045);
nor U16930 (N_16930,N_11979,N_10090);
or U16931 (N_16931,N_13040,N_11599);
nand U16932 (N_16932,N_14775,N_11725);
nand U16933 (N_16933,N_12708,N_14138);
xnor U16934 (N_16934,N_11807,N_13815);
xor U16935 (N_16935,N_14670,N_14410);
or U16936 (N_16936,N_12160,N_10241);
xor U16937 (N_16937,N_12405,N_12013);
nand U16938 (N_16938,N_11171,N_14071);
or U16939 (N_16939,N_11019,N_10935);
nor U16940 (N_16940,N_10609,N_11029);
and U16941 (N_16941,N_12204,N_13682);
and U16942 (N_16942,N_10521,N_10524);
nand U16943 (N_16943,N_11693,N_11619);
xnor U16944 (N_16944,N_13497,N_12043);
nor U16945 (N_16945,N_10630,N_12138);
nor U16946 (N_16946,N_13557,N_12748);
nand U16947 (N_16947,N_14213,N_10096);
xor U16948 (N_16948,N_11504,N_11012);
nor U16949 (N_16949,N_11118,N_11908);
nor U16950 (N_16950,N_12403,N_13063);
nor U16951 (N_16951,N_11773,N_14551);
nor U16952 (N_16952,N_14332,N_10774);
xor U16953 (N_16953,N_10549,N_14894);
xor U16954 (N_16954,N_12980,N_12356);
xnor U16955 (N_16955,N_10441,N_13046);
xor U16956 (N_16956,N_14815,N_13124);
or U16957 (N_16957,N_14163,N_11115);
nand U16958 (N_16958,N_10624,N_14060);
xnor U16959 (N_16959,N_12119,N_13773);
or U16960 (N_16960,N_12895,N_13281);
xor U16961 (N_16961,N_12633,N_13648);
xnor U16962 (N_16962,N_14901,N_12918);
or U16963 (N_16963,N_10596,N_11717);
nand U16964 (N_16964,N_13189,N_13297);
nand U16965 (N_16965,N_13859,N_10703);
nand U16966 (N_16966,N_12556,N_12665);
and U16967 (N_16967,N_13970,N_10541);
and U16968 (N_16968,N_10316,N_12483);
nor U16969 (N_16969,N_12171,N_14761);
xor U16970 (N_16970,N_13069,N_11896);
nand U16971 (N_16971,N_10876,N_13803);
xnor U16972 (N_16972,N_10826,N_14669);
xor U16973 (N_16973,N_10823,N_13540);
or U16974 (N_16974,N_11919,N_12080);
nand U16975 (N_16975,N_14806,N_10060);
nor U16976 (N_16976,N_11605,N_10037);
or U16977 (N_16977,N_11474,N_10485);
or U16978 (N_16978,N_13975,N_11779);
nor U16979 (N_16979,N_10741,N_11410);
or U16980 (N_16980,N_10855,N_13700);
nand U16981 (N_16981,N_11868,N_12488);
nor U16982 (N_16982,N_14584,N_11547);
and U16983 (N_16983,N_14725,N_12320);
nor U16984 (N_16984,N_13879,N_11764);
nand U16985 (N_16985,N_12846,N_12728);
nand U16986 (N_16986,N_11793,N_13806);
or U16987 (N_16987,N_12399,N_13587);
nor U16988 (N_16988,N_14911,N_10786);
nand U16989 (N_16989,N_14749,N_10540);
and U16990 (N_16990,N_13232,N_14883);
nand U16991 (N_16991,N_10419,N_13487);
nand U16992 (N_16992,N_10571,N_14211);
nand U16993 (N_16993,N_11193,N_14849);
xnor U16994 (N_16994,N_10450,N_10953);
or U16995 (N_16995,N_11165,N_11582);
and U16996 (N_16996,N_11915,N_11392);
nand U16997 (N_16997,N_11177,N_12422);
xnor U16998 (N_16998,N_12704,N_10132);
and U16999 (N_16999,N_14514,N_12668);
nor U17000 (N_17000,N_12881,N_14053);
or U17001 (N_17001,N_11729,N_11855);
nor U17002 (N_17002,N_13959,N_12135);
and U17003 (N_17003,N_10871,N_14459);
xnor U17004 (N_17004,N_14566,N_12235);
or U17005 (N_17005,N_11294,N_14690);
or U17006 (N_17006,N_10480,N_13792);
xor U17007 (N_17007,N_10781,N_13274);
nor U17008 (N_17008,N_13708,N_13580);
xnor U17009 (N_17009,N_14046,N_11614);
and U17010 (N_17010,N_12458,N_13105);
or U17011 (N_17011,N_10208,N_11971);
nor U17012 (N_17012,N_14862,N_14743);
nor U17013 (N_17013,N_14348,N_10378);
and U17014 (N_17014,N_13668,N_12779);
and U17015 (N_17015,N_13264,N_14931);
nor U17016 (N_17016,N_14470,N_10073);
nor U17017 (N_17017,N_13582,N_11200);
or U17018 (N_17018,N_11492,N_11101);
nand U17019 (N_17019,N_12560,N_10853);
and U17020 (N_17020,N_11730,N_11371);
and U17021 (N_17021,N_13758,N_11233);
xnor U17022 (N_17022,N_10987,N_12954);
xnor U17023 (N_17023,N_12364,N_14056);
and U17024 (N_17024,N_14925,N_13203);
and U17025 (N_17025,N_12142,N_10442);
or U17026 (N_17026,N_10082,N_10421);
and U17027 (N_17027,N_13958,N_10973);
xnor U17028 (N_17028,N_10923,N_13555);
nor U17029 (N_17029,N_12865,N_14653);
nor U17030 (N_17030,N_11690,N_10724);
or U17031 (N_17031,N_14510,N_11009);
and U17032 (N_17032,N_10790,N_14495);
xnor U17033 (N_17033,N_10827,N_10769);
and U17034 (N_17034,N_11438,N_12813);
xnor U17035 (N_17035,N_12550,N_13838);
nand U17036 (N_17036,N_10167,N_14528);
xnor U17037 (N_17037,N_10507,N_14953);
and U17038 (N_17038,N_10336,N_12349);
or U17039 (N_17039,N_14113,N_12793);
nor U17040 (N_17040,N_10841,N_13954);
or U17041 (N_17041,N_10929,N_14096);
and U17042 (N_17042,N_10551,N_10022);
or U17043 (N_17043,N_14358,N_13250);
nand U17044 (N_17044,N_13230,N_10759);
or U17045 (N_17045,N_13953,N_11173);
and U17046 (N_17046,N_14229,N_10721);
or U17047 (N_17047,N_11791,N_14409);
nand U17048 (N_17048,N_13490,N_13317);
or U17049 (N_17049,N_14168,N_10216);
or U17050 (N_17050,N_13581,N_14588);
nor U17051 (N_17051,N_12914,N_14252);
nand U17052 (N_17052,N_12317,N_14207);
or U17053 (N_17053,N_10048,N_10864);
nor U17054 (N_17054,N_13503,N_11943);
xor U17055 (N_17055,N_12379,N_14457);
and U17056 (N_17056,N_14504,N_14534);
and U17057 (N_17057,N_13508,N_11658);
nand U17058 (N_17058,N_12719,N_10041);
nor U17059 (N_17059,N_13920,N_11750);
xnor U17060 (N_17060,N_12893,N_10888);
or U17061 (N_17061,N_13689,N_10182);
xnor U17062 (N_17062,N_13600,N_11196);
and U17063 (N_17063,N_12552,N_10878);
xor U17064 (N_17064,N_14932,N_11001);
and U17065 (N_17065,N_12461,N_11543);
and U17066 (N_17066,N_13734,N_14373);
xnor U17067 (N_17067,N_13997,N_14162);
xor U17068 (N_17068,N_10324,N_12192);
nand U17069 (N_17069,N_14197,N_14603);
or U17070 (N_17070,N_13948,N_14727);
xor U17071 (N_17071,N_14201,N_14075);
and U17072 (N_17072,N_11300,N_13559);
nand U17073 (N_17073,N_13946,N_11363);
or U17074 (N_17074,N_11994,N_13268);
or U17075 (N_17075,N_12038,N_14054);
or U17076 (N_17076,N_10348,N_12342);
or U17077 (N_17077,N_13476,N_14962);
or U17078 (N_17078,N_14490,N_10307);
xnor U17079 (N_17079,N_12209,N_12832);
nor U17080 (N_17080,N_11823,N_13197);
or U17081 (N_17081,N_10120,N_10177);
xor U17082 (N_17082,N_12854,N_13412);
or U17083 (N_17083,N_10055,N_14839);
xor U17084 (N_17084,N_11560,N_14493);
nand U17085 (N_17085,N_10464,N_13121);
nand U17086 (N_17086,N_10168,N_12630);
and U17087 (N_17087,N_14397,N_13549);
xor U17088 (N_17088,N_10914,N_14111);
and U17089 (N_17089,N_10295,N_14692);
nand U17090 (N_17090,N_11552,N_12010);
and U17091 (N_17091,N_12524,N_11933);
and U17092 (N_17092,N_13075,N_14887);
xor U17093 (N_17093,N_13799,N_13715);
nor U17094 (N_17094,N_10550,N_13840);
or U17095 (N_17095,N_12070,N_13440);
xnor U17096 (N_17096,N_11489,N_12166);
and U17097 (N_17097,N_14390,N_12675);
xor U17098 (N_17098,N_13033,N_14724);
nor U17099 (N_17099,N_13186,N_11815);
xor U17100 (N_17100,N_12205,N_10590);
nand U17101 (N_17101,N_10044,N_11992);
or U17102 (N_17102,N_14972,N_14137);
nor U17103 (N_17103,N_10289,N_11229);
nor U17104 (N_17104,N_11178,N_13467);
or U17105 (N_17105,N_11911,N_11450);
xor U17106 (N_17106,N_11297,N_11426);
xnor U17107 (N_17107,N_11021,N_13463);
nand U17108 (N_17108,N_12947,N_10543);
nand U17109 (N_17109,N_13120,N_12386);
and U17110 (N_17110,N_13355,N_13984);
xnor U17111 (N_17111,N_10655,N_10523);
nand U17112 (N_17112,N_10373,N_10772);
nand U17113 (N_17113,N_11244,N_11997);
nor U17114 (N_17114,N_10085,N_13128);
and U17115 (N_17115,N_11946,N_10575);
and U17116 (N_17116,N_12872,N_14688);
nor U17117 (N_17117,N_13905,N_14364);
nand U17118 (N_17118,N_14847,N_14796);
and U17119 (N_17119,N_13225,N_11828);
xor U17120 (N_17120,N_10013,N_13939);
xor U17121 (N_17121,N_11418,N_11873);
or U17122 (N_17122,N_12174,N_14477);
or U17123 (N_17123,N_13605,N_14502);
xor U17124 (N_17124,N_10353,N_10141);
or U17125 (N_17125,N_10513,N_11018);
nand U17126 (N_17126,N_10051,N_10728);
and U17127 (N_17127,N_12290,N_12490);
and U17128 (N_17128,N_12732,N_14322);
nand U17129 (N_17129,N_11204,N_14646);
and U17130 (N_17130,N_14525,N_13237);
nor U17131 (N_17131,N_11733,N_13139);
nand U17132 (N_17132,N_11737,N_12605);
xnor U17133 (N_17133,N_11673,N_13308);
or U17134 (N_17134,N_14029,N_13242);
and U17135 (N_17135,N_11872,N_11296);
xor U17136 (N_17136,N_12955,N_14001);
xor U17137 (N_17137,N_12450,N_12972);
and U17138 (N_17138,N_10642,N_11506);
or U17139 (N_17139,N_13742,N_11938);
xor U17140 (N_17140,N_10796,N_10118);
or U17141 (N_17141,N_11628,N_14202);
nor U17142 (N_17142,N_14483,N_10843);
xor U17143 (N_17143,N_14351,N_10150);
xnor U17144 (N_17144,N_10961,N_13342);
xnor U17145 (N_17145,N_11762,N_10775);
nor U17146 (N_17146,N_10730,N_10361);
xnor U17147 (N_17147,N_13519,N_10338);
or U17148 (N_17148,N_10377,N_10842);
xor U17149 (N_17149,N_14589,N_12790);
and U17150 (N_17150,N_12067,N_11961);
xor U17151 (N_17151,N_10453,N_12798);
and U17152 (N_17152,N_12695,N_12614);
or U17153 (N_17153,N_12456,N_13199);
and U17154 (N_17154,N_13620,N_13822);
and U17155 (N_17155,N_10974,N_12752);
nand U17156 (N_17156,N_11801,N_12485);
or U17157 (N_17157,N_10656,N_11759);
nor U17158 (N_17158,N_11478,N_13188);
nor U17159 (N_17159,N_12499,N_11888);
xnor U17160 (N_17160,N_14891,N_11916);
nand U17161 (N_17161,N_11501,N_14505);
nor U17162 (N_17162,N_11976,N_14341);
nand U17163 (N_17163,N_12653,N_14772);
nand U17164 (N_17164,N_12518,N_11541);
nor U17165 (N_17165,N_12273,N_10088);
xor U17166 (N_17166,N_12087,N_10950);
nor U17167 (N_17167,N_10565,N_10611);
or U17168 (N_17168,N_11142,N_10399);
and U17169 (N_17169,N_11583,N_12920);
and U17170 (N_17170,N_10178,N_10862);
and U17171 (N_17171,N_13713,N_14365);
xnor U17172 (N_17172,N_10653,N_10026);
xor U17173 (N_17173,N_14784,N_11235);
or U17174 (N_17174,N_10002,N_11874);
xor U17175 (N_17175,N_12352,N_10232);
nand U17176 (N_17176,N_10869,N_10479);
nand U17177 (N_17177,N_14040,N_13646);
nor U17178 (N_17178,N_12819,N_11941);
nor U17179 (N_17179,N_14074,N_12432);
or U17180 (N_17180,N_13319,N_14766);
nand U17181 (N_17181,N_12426,N_11170);
or U17182 (N_17182,N_14864,N_10130);
and U17183 (N_17183,N_13639,N_12429);
xor U17184 (N_17184,N_13421,N_11301);
nand U17185 (N_17185,N_14789,N_11131);
or U17186 (N_17186,N_10420,N_12176);
or U17187 (N_17187,N_14297,N_12744);
and U17188 (N_17188,N_13507,N_13889);
or U17189 (N_17189,N_10425,N_10512);
nor U17190 (N_17190,N_14102,N_13886);
nand U17191 (N_17191,N_10787,N_14215);
nand U17192 (N_17192,N_13569,N_12126);
xor U17193 (N_17193,N_13326,N_11022);
and U17194 (N_17194,N_11152,N_10771);
nor U17195 (N_17195,N_11514,N_10875);
nor U17196 (N_17196,N_14671,N_13240);
xor U17197 (N_17197,N_11834,N_13568);
or U17198 (N_17198,N_10641,N_14644);
xor U17199 (N_17199,N_10358,N_13986);
nor U17200 (N_17200,N_10675,N_14475);
and U17201 (N_17201,N_12555,N_13007);
or U17202 (N_17202,N_11849,N_14763);
nor U17203 (N_17203,N_11343,N_13928);
or U17204 (N_17204,N_11322,N_10693);
or U17205 (N_17205,N_14959,N_10739);
nand U17206 (N_17206,N_14521,N_11539);
xor U17207 (N_17207,N_10694,N_11139);
nor U17208 (N_17208,N_12143,N_10224);
xor U17209 (N_17209,N_13824,N_10162);
nor U17210 (N_17210,N_13945,N_10882);
or U17211 (N_17211,N_13328,N_14081);
and U17212 (N_17212,N_10443,N_14845);
and U17213 (N_17213,N_13072,N_11700);
nor U17214 (N_17214,N_10416,N_12339);
nor U17215 (N_17215,N_14781,N_12168);
nor U17216 (N_17216,N_13397,N_10444);
nor U17217 (N_17217,N_14691,N_12984);
xnor U17218 (N_17218,N_10957,N_12583);
nor U17219 (N_17219,N_12341,N_13593);
xnor U17220 (N_17220,N_13495,N_11455);
xor U17221 (N_17221,N_13938,N_14822);
xnor U17222 (N_17222,N_10275,N_12028);
xnor U17223 (N_17223,N_10978,N_10764);
or U17224 (N_17224,N_11482,N_14461);
and U17225 (N_17225,N_13261,N_12755);
nor U17226 (N_17226,N_12863,N_12803);
nand U17227 (N_17227,N_11993,N_14421);
and U17228 (N_17228,N_11354,N_10740);
nor U17229 (N_17229,N_13212,N_12410);
and U17230 (N_17230,N_13429,N_12681);
and U17231 (N_17231,N_10965,N_12792);
and U17232 (N_17232,N_14094,N_10572);
nor U17233 (N_17233,N_10163,N_12698);
or U17234 (N_17234,N_14717,N_10808);
nand U17235 (N_17235,N_11757,N_12716);
or U17236 (N_17236,N_10665,N_12510);
xor U17237 (N_17237,N_14170,N_14356);
xnor U17238 (N_17238,N_14443,N_14152);
nand U17239 (N_17239,N_11568,N_11017);
or U17240 (N_17240,N_10768,N_14317);
and U17241 (N_17241,N_14855,N_10814);
xnor U17242 (N_17242,N_12147,N_14267);
and U17243 (N_17243,N_13290,N_13626);
and U17244 (N_17244,N_11206,N_13285);
and U17245 (N_17245,N_13558,N_14450);
nor U17246 (N_17246,N_14812,N_14082);
and U17247 (N_17247,N_10912,N_10896);
or U17248 (N_17248,N_10736,N_12963);
and U17249 (N_17249,N_11436,N_13753);
xor U17250 (N_17250,N_12257,N_12769);
or U17251 (N_17251,N_12091,N_12248);
xor U17252 (N_17252,N_11138,N_11381);
xor U17253 (N_17253,N_14013,N_11577);
xor U17254 (N_17254,N_13327,N_13174);
nand U17255 (N_17255,N_13279,N_12838);
or U17256 (N_17256,N_11500,N_12095);
nand U17257 (N_17257,N_12974,N_11805);
xnor U17258 (N_17258,N_14563,N_14176);
nor U17259 (N_17259,N_12672,N_14256);
and U17260 (N_17260,N_14120,N_11825);
nand U17261 (N_17261,N_11870,N_13277);
nor U17262 (N_17262,N_10751,N_12559);
nor U17263 (N_17263,N_11950,N_12373);
nor U17264 (N_17264,N_14208,N_14807);
or U17265 (N_17265,N_14110,N_11023);
xor U17266 (N_17266,N_14501,N_14733);
nor U17267 (N_17267,N_13115,N_12331);
or U17268 (N_17268,N_12110,N_13599);
nand U17269 (N_17269,N_12008,N_10016);
xnor U17270 (N_17270,N_10394,N_14423);
nand U17271 (N_17271,N_10528,N_10650);
nor U17272 (N_17272,N_13493,N_14293);
or U17273 (N_17273,N_13553,N_13829);
nand U17274 (N_17274,N_10795,N_14597);
nor U17275 (N_17275,N_13349,N_12939);
or U17276 (N_17276,N_13200,N_13052);
xor U17277 (N_17277,N_14335,N_10413);
nor U17278 (N_17278,N_12200,N_10187);
or U17279 (N_17279,N_14494,N_14115);
and U17280 (N_17280,N_14022,N_10979);
or U17281 (N_17281,N_12913,N_10081);
xor U17282 (N_17282,N_13727,N_14523);
xor U17283 (N_17283,N_10742,N_10332);
nand U17284 (N_17284,N_12239,N_10903);
or U17285 (N_17285,N_13047,N_12542);
or U17286 (N_17286,N_10618,N_10900);
nand U17287 (N_17287,N_12267,N_10531);
nor U17288 (N_17288,N_11989,N_11609);
or U17289 (N_17289,N_10931,N_10349);
or U17290 (N_17290,N_11399,N_13965);
and U17291 (N_17291,N_14744,N_14314);
or U17292 (N_17292,N_11167,N_10830);
nor U17293 (N_17293,N_14279,N_11246);
nand U17294 (N_17294,N_13571,N_13044);
nand U17295 (N_17295,N_12767,N_13151);
xor U17296 (N_17296,N_14270,N_11270);
nor U17297 (N_17297,N_13854,N_11512);
and U17298 (N_17298,N_10776,N_14592);
nor U17299 (N_17299,N_11378,N_12058);
and U17300 (N_17300,N_11551,N_13270);
and U17301 (N_17301,N_11910,N_13266);
nand U17302 (N_17302,N_12946,N_14230);
nand U17303 (N_17303,N_14970,N_12049);
and U17304 (N_17304,N_12124,N_12688);
or U17305 (N_17305,N_14570,N_13991);
nand U17306 (N_17306,N_13439,N_13791);
and U17307 (N_17307,N_13510,N_10325);
and U17308 (N_17308,N_11613,N_14224);
or U17309 (N_17309,N_12795,N_11901);
and U17310 (N_17310,N_13260,N_11969);
xnor U17311 (N_17311,N_14305,N_11899);
nor U17312 (N_17312,N_13054,N_13450);
nor U17313 (N_17313,N_12786,N_13769);
nand U17314 (N_17314,N_13249,N_13255);
xnor U17315 (N_17315,N_10788,N_14939);
nand U17316 (N_17316,N_13404,N_13070);
xor U17317 (N_17317,N_11960,N_14434);
and U17318 (N_17318,N_13015,N_11396);
or U17319 (N_17319,N_10588,N_10475);
xor U17320 (N_17320,N_11124,N_13053);
nor U17321 (N_17321,N_14057,N_14636);
and U17322 (N_17322,N_14593,N_14065);
nor U17323 (N_17323,N_10685,N_10707);
xor U17324 (N_17324,N_12797,N_11752);
nand U17325 (N_17325,N_12395,N_11912);
xnor U17326 (N_17326,N_12788,N_14787);
nand U17327 (N_17327,N_11407,N_14667);
or U17328 (N_17328,N_13184,N_11342);
and U17329 (N_17329,N_12727,N_10968);
nor U17330 (N_17330,N_11084,N_10143);
nand U17331 (N_17331,N_10422,N_12501);
or U17332 (N_17332,N_12297,N_14141);
nor U17333 (N_17333,N_10836,N_10357);
nand U17334 (N_17334,N_11479,N_12986);
and U17335 (N_17335,N_14026,N_12314);
xnor U17336 (N_17336,N_11695,N_10188);
and U17337 (N_17337,N_12340,N_14204);
and U17338 (N_17338,N_11869,N_13690);
nand U17339 (N_17339,N_10260,N_14587);
and U17340 (N_17340,N_12261,N_13244);
nor U17341 (N_17341,N_11262,N_11282);
nor U17342 (N_17342,N_10567,N_11271);
and U17343 (N_17343,N_11923,N_14809);
xor U17344 (N_17344,N_12924,N_10839);
nand U17345 (N_17345,N_13472,N_14024);
and U17346 (N_17346,N_10964,N_12300);
nand U17347 (N_17347,N_10564,N_10860);
xnor U17348 (N_17348,N_11625,N_12602);
nand U17349 (N_17349,N_13764,N_12052);
xor U17350 (N_17350,N_13168,N_12900);
or U17351 (N_17351,N_10607,N_14943);
nor U17352 (N_17352,N_11182,N_13642);
nand U17353 (N_17353,N_12685,N_10597);
xor U17354 (N_17354,N_10481,N_10927);
xnor U17355 (N_17355,N_12759,N_13725);
and U17356 (N_17356,N_10009,N_10792);
nor U17357 (N_17357,N_12184,N_13892);
or U17358 (N_17358,N_14089,N_10517);
nand U17359 (N_17359,N_11720,N_13122);
and U17360 (N_17360,N_11288,N_10298);
xor U17361 (N_17361,N_12966,N_14066);
nor U17362 (N_17362,N_13363,N_12874);
nand U17363 (N_17363,N_10299,N_12836);
or U17364 (N_17364,N_12761,N_14360);
nor U17365 (N_17365,N_13897,N_11285);
xor U17366 (N_17366,N_11768,N_11709);
and U17367 (N_17367,N_10960,N_10161);
nand U17368 (N_17368,N_11038,N_11883);
xnor U17369 (N_17369,N_12005,N_10939);
nand U17370 (N_17370,N_14496,N_12721);
or U17371 (N_17371,N_13544,N_10432);
or U17372 (N_17372,N_14538,N_11346);
nand U17373 (N_17373,N_13721,N_10631);
nand U17374 (N_17374,N_11749,N_12401);
and U17375 (N_17375,N_13651,N_10102);
nand U17376 (N_17376,N_14378,N_11840);
or U17377 (N_17377,N_10870,N_13140);
nor U17378 (N_17378,N_10283,N_11611);
or U17379 (N_17379,N_12647,N_14092);
xnor U17380 (N_17380,N_12278,N_11459);
nor U17381 (N_17381,N_14578,N_10366);
nor U17382 (N_17382,N_11128,N_14480);
nor U17383 (N_17383,N_13284,N_11254);
nand U17384 (N_17384,N_12981,N_13924);
xnor U17385 (N_17385,N_10321,N_11398);
xnor U17386 (N_17386,N_11845,N_13594);
nand U17387 (N_17387,N_13887,N_14222);
or U17388 (N_17388,N_14751,N_12367);
xor U17389 (N_17389,N_12243,N_13448);
or U17390 (N_17390,N_14828,N_11510);
xnor U17391 (N_17391,N_13877,N_13533);
and U17392 (N_17392,N_12722,N_13372);
nor U17393 (N_17393,N_13993,N_12627);
or U17394 (N_17394,N_12303,N_13554);
and U17395 (N_17395,N_10206,N_14389);
and U17396 (N_17396,N_14261,N_11210);
nor U17397 (N_17397,N_12081,N_13772);
or U17398 (N_17398,N_13966,N_12376);
nand U17399 (N_17399,N_14735,N_12514);
xor U17400 (N_17400,N_12669,N_11005);
or U17401 (N_17401,N_12153,N_14449);
nor U17402 (N_17402,N_12062,N_11185);
xnor U17403 (N_17403,N_14238,N_11219);
and U17404 (N_17404,N_12637,N_11795);
or U17405 (N_17405,N_13691,N_10489);
nand U17406 (N_17406,N_13918,N_10989);
and U17407 (N_17407,N_13845,N_13779);
or U17408 (N_17408,N_10920,N_10779);
and U17409 (N_17409,N_13210,N_11529);
nor U17410 (N_17410,N_14209,N_13374);
and U17411 (N_17411,N_11242,N_13956);
and U17412 (N_17412,N_12578,N_13334);
nand U17413 (N_17413,N_13164,N_14108);
and U17414 (N_17414,N_12639,N_10812);
and U17415 (N_17415,N_12674,N_14063);
nand U17416 (N_17416,N_11441,N_11817);
or U17417 (N_17417,N_13538,N_10429);
xnor U17418 (N_17418,N_14500,N_12928);
nand U17419 (N_17419,N_13989,N_14463);
nor U17420 (N_17420,N_14888,N_11130);
nand U17421 (N_17421,N_12262,N_13201);
xor U17422 (N_17422,N_11010,N_12791);
or U17423 (N_17423,N_13292,N_13616);
xor U17424 (N_17424,N_13438,N_11966);
nand U17425 (N_17425,N_12937,N_14794);
and U17426 (N_17426,N_14937,N_11592);
and U17427 (N_17427,N_13062,N_12844);
nor U17428 (N_17428,N_10829,N_11587);
nor U17429 (N_17429,N_14982,N_11591);
and U17430 (N_17430,N_14979,N_14917);
nand U17431 (N_17431,N_11088,N_12919);
or U17432 (N_17432,N_14228,N_13932);
nand U17433 (N_17433,N_11247,N_11386);
and U17434 (N_17434,N_10969,N_11144);
nor U17435 (N_17435,N_14582,N_10271);
nand U17436 (N_17436,N_14274,N_11522);
xor U17437 (N_17437,N_11735,N_13043);
or U17438 (N_17438,N_14429,N_13589);
xnor U17439 (N_17439,N_10488,N_12944);
nand U17440 (N_17440,N_12446,N_10412);
xor U17441 (N_17441,N_13676,N_11776);
or U17442 (N_17442,N_11093,N_14561);
and U17443 (N_17443,N_11836,N_10094);
or U17444 (N_17444,N_12694,N_11893);
xor U17445 (N_17445,N_13368,N_11283);
or U17446 (N_17446,N_13678,N_14112);
xnor U17447 (N_17447,N_12942,N_14363);
or U17448 (N_17448,N_11374,N_11089);
and U17449 (N_17449,N_12172,N_10198);
or U17450 (N_17450,N_14148,N_13940);
nor U17451 (N_17451,N_13389,N_14550);
xor U17452 (N_17452,N_12690,N_13515);
nor U17453 (N_17453,N_14396,N_11408);
and U17454 (N_17454,N_13315,N_11411);
and U17455 (N_17455,N_11627,N_14540);
or U17456 (N_17456,N_12029,N_14005);
nand U17457 (N_17457,N_12207,N_14803);
xnor U17458 (N_17458,N_10415,N_13980);
or U17459 (N_17459,N_11850,N_11469);
nand U17460 (N_17460,N_11917,N_12871);
xor U17461 (N_17461,N_13248,N_11999);
or U17462 (N_17462,N_12040,N_12693);
and U17463 (N_17463,N_13304,N_14974);
and U17464 (N_17464,N_13136,N_10004);
nand U17465 (N_17465,N_13306,N_12975);
and U17466 (N_17466,N_10913,N_10136);
xnor U17467 (N_17467,N_14319,N_11882);
xnor U17468 (N_17468,N_13785,N_12718);
and U17469 (N_17469,N_12288,N_10100);
xor U17470 (N_17470,N_13082,N_11493);
and U17471 (N_17471,N_11974,N_13318);
or U17472 (N_17472,N_14600,N_10440);
and U17473 (N_17473,N_12484,N_13078);
nand U17474 (N_17474,N_11925,N_10925);
nor U17475 (N_17475,N_10810,N_12949);
nand U17476 (N_17476,N_13586,N_13321);
or U17477 (N_17477,N_13027,N_11065);
and U17478 (N_17478,N_11397,N_14810);
nand U17479 (N_17479,N_12496,N_14759);
or U17480 (N_17480,N_11524,N_12833);
nor U17481 (N_17481,N_14139,N_14133);
or U17482 (N_17482,N_12369,N_11485);
or U17483 (N_17483,N_11066,N_10718);
or U17484 (N_17484,N_12877,N_10817);
nor U17485 (N_17485,N_14304,N_11055);
or U17486 (N_17486,N_14971,N_12523);
and U17487 (N_17487,N_12118,N_11231);
nand U17488 (N_17488,N_13192,N_12291);
nor U17489 (N_17489,N_11637,N_14729);
or U17490 (N_17490,N_14732,N_14469);
or U17491 (N_17491,N_11570,N_10629);
nor U17492 (N_17492,N_13035,N_13411);
nor U17493 (N_17493,N_10426,N_11615);
or U17494 (N_17494,N_12327,N_12689);
or U17495 (N_17495,N_14248,N_11388);
or U17496 (N_17496,N_13512,N_10530);
nand U17497 (N_17497,N_14420,N_14927);
or U17498 (N_17498,N_14124,N_10006);
and U17499 (N_17499,N_11187,N_11416);
and U17500 (N_17500,N_11125,N_12040);
or U17501 (N_17501,N_13670,N_12850);
nand U17502 (N_17502,N_14036,N_11581);
xnor U17503 (N_17503,N_13118,N_10986);
nand U17504 (N_17504,N_10491,N_12938);
and U17505 (N_17505,N_10726,N_10332);
and U17506 (N_17506,N_12755,N_13473);
xor U17507 (N_17507,N_10386,N_10510);
xnor U17508 (N_17508,N_10491,N_10958);
and U17509 (N_17509,N_12120,N_10507);
nor U17510 (N_17510,N_11751,N_14550);
nor U17511 (N_17511,N_13958,N_10752);
or U17512 (N_17512,N_14141,N_13710);
or U17513 (N_17513,N_14107,N_11334);
and U17514 (N_17514,N_11605,N_13622);
nand U17515 (N_17515,N_12968,N_14369);
nor U17516 (N_17516,N_14536,N_14946);
or U17517 (N_17517,N_12394,N_10192);
and U17518 (N_17518,N_10996,N_11919);
nand U17519 (N_17519,N_10442,N_11881);
xor U17520 (N_17520,N_13378,N_10135);
and U17521 (N_17521,N_12838,N_14916);
nand U17522 (N_17522,N_12463,N_13276);
or U17523 (N_17523,N_11809,N_13824);
and U17524 (N_17524,N_10995,N_13161);
or U17525 (N_17525,N_10531,N_10025);
and U17526 (N_17526,N_14728,N_12587);
xor U17527 (N_17527,N_10775,N_14764);
or U17528 (N_17528,N_14936,N_13987);
nand U17529 (N_17529,N_14911,N_11871);
xor U17530 (N_17530,N_13084,N_10955);
or U17531 (N_17531,N_10006,N_12176);
and U17532 (N_17532,N_10797,N_10648);
nand U17533 (N_17533,N_11715,N_12926);
or U17534 (N_17534,N_12263,N_14498);
xnor U17535 (N_17535,N_14900,N_13651);
xor U17536 (N_17536,N_14988,N_13314);
and U17537 (N_17537,N_13056,N_13692);
or U17538 (N_17538,N_11931,N_14025);
nand U17539 (N_17539,N_13123,N_11608);
or U17540 (N_17540,N_10908,N_14798);
xor U17541 (N_17541,N_12294,N_11027);
nor U17542 (N_17542,N_12909,N_12168);
nor U17543 (N_17543,N_10433,N_10519);
and U17544 (N_17544,N_14944,N_12927);
nand U17545 (N_17545,N_14004,N_12060);
nand U17546 (N_17546,N_13439,N_11656);
or U17547 (N_17547,N_14129,N_13451);
nand U17548 (N_17548,N_10290,N_13358);
nand U17549 (N_17549,N_14021,N_11943);
and U17550 (N_17550,N_14415,N_10616);
or U17551 (N_17551,N_13094,N_10035);
and U17552 (N_17552,N_13431,N_10665);
and U17553 (N_17553,N_12816,N_14474);
or U17554 (N_17554,N_11997,N_11118);
xor U17555 (N_17555,N_14515,N_14691);
nand U17556 (N_17556,N_12116,N_11824);
xor U17557 (N_17557,N_12807,N_11425);
nor U17558 (N_17558,N_13669,N_13328);
or U17559 (N_17559,N_14976,N_14181);
and U17560 (N_17560,N_13346,N_12787);
xor U17561 (N_17561,N_12569,N_11709);
nand U17562 (N_17562,N_14058,N_11555);
nor U17563 (N_17563,N_14605,N_12455);
or U17564 (N_17564,N_11301,N_13295);
or U17565 (N_17565,N_12609,N_13706);
xor U17566 (N_17566,N_12519,N_11126);
nor U17567 (N_17567,N_10212,N_10419);
nor U17568 (N_17568,N_14345,N_10687);
or U17569 (N_17569,N_11843,N_12428);
or U17570 (N_17570,N_11934,N_10032);
nor U17571 (N_17571,N_11486,N_14742);
and U17572 (N_17572,N_13531,N_11476);
xnor U17573 (N_17573,N_14824,N_10164);
nand U17574 (N_17574,N_14802,N_14172);
xnor U17575 (N_17575,N_14369,N_10712);
xnor U17576 (N_17576,N_14010,N_13971);
and U17577 (N_17577,N_11275,N_13235);
nor U17578 (N_17578,N_11013,N_10692);
nand U17579 (N_17579,N_10195,N_10522);
nand U17580 (N_17580,N_14755,N_10852);
or U17581 (N_17581,N_10288,N_13646);
and U17582 (N_17582,N_14957,N_14650);
or U17583 (N_17583,N_10072,N_13393);
and U17584 (N_17584,N_14874,N_11081);
and U17585 (N_17585,N_12212,N_13349);
nor U17586 (N_17586,N_13904,N_12882);
or U17587 (N_17587,N_11830,N_12594);
xnor U17588 (N_17588,N_14563,N_12137);
and U17589 (N_17589,N_12899,N_13913);
nor U17590 (N_17590,N_11714,N_13967);
xor U17591 (N_17591,N_12447,N_14482);
xor U17592 (N_17592,N_12428,N_12703);
xnor U17593 (N_17593,N_14972,N_13660);
xnor U17594 (N_17594,N_13533,N_13856);
and U17595 (N_17595,N_10497,N_10631);
and U17596 (N_17596,N_12269,N_14098);
or U17597 (N_17597,N_11791,N_10592);
or U17598 (N_17598,N_13421,N_13878);
nand U17599 (N_17599,N_12141,N_13201);
and U17600 (N_17600,N_10476,N_12529);
xor U17601 (N_17601,N_11389,N_12237);
xnor U17602 (N_17602,N_11895,N_10419);
or U17603 (N_17603,N_14172,N_14982);
xor U17604 (N_17604,N_11759,N_12953);
xor U17605 (N_17605,N_11925,N_10030);
or U17606 (N_17606,N_12966,N_13863);
nor U17607 (N_17607,N_12009,N_14877);
nand U17608 (N_17608,N_13670,N_13967);
xnor U17609 (N_17609,N_12717,N_12585);
nor U17610 (N_17610,N_14851,N_11258);
xor U17611 (N_17611,N_12716,N_12550);
and U17612 (N_17612,N_12778,N_14555);
nor U17613 (N_17613,N_12452,N_11105);
and U17614 (N_17614,N_14662,N_12546);
nor U17615 (N_17615,N_14534,N_10948);
nor U17616 (N_17616,N_10588,N_14088);
xnor U17617 (N_17617,N_12410,N_13284);
nand U17618 (N_17618,N_11083,N_12507);
nand U17619 (N_17619,N_10285,N_10782);
xor U17620 (N_17620,N_13222,N_11923);
and U17621 (N_17621,N_11967,N_12481);
xnor U17622 (N_17622,N_13012,N_12084);
or U17623 (N_17623,N_11309,N_14022);
nand U17624 (N_17624,N_14487,N_11089);
nor U17625 (N_17625,N_10673,N_11725);
or U17626 (N_17626,N_13252,N_11275);
xor U17627 (N_17627,N_11675,N_14322);
nand U17628 (N_17628,N_12952,N_10540);
and U17629 (N_17629,N_10806,N_14278);
xnor U17630 (N_17630,N_13589,N_11732);
xor U17631 (N_17631,N_12293,N_14513);
or U17632 (N_17632,N_13690,N_14261);
nor U17633 (N_17633,N_14807,N_13517);
nand U17634 (N_17634,N_13089,N_14248);
nand U17635 (N_17635,N_13519,N_11235);
nor U17636 (N_17636,N_14031,N_10343);
and U17637 (N_17637,N_14659,N_13210);
or U17638 (N_17638,N_11048,N_13496);
and U17639 (N_17639,N_11415,N_14221);
or U17640 (N_17640,N_13483,N_14905);
nand U17641 (N_17641,N_10305,N_14024);
nand U17642 (N_17642,N_10569,N_10692);
xor U17643 (N_17643,N_10967,N_14257);
and U17644 (N_17644,N_13441,N_13279);
nor U17645 (N_17645,N_14203,N_14382);
nor U17646 (N_17646,N_12394,N_11833);
xnor U17647 (N_17647,N_10027,N_10137);
nor U17648 (N_17648,N_14204,N_12969);
or U17649 (N_17649,N_14681,N_13837);
and U17650 (N_17650,N_14415,N_10267);
nand U17651 (N_17651,N_12681,N_11342);
nor U17652 (N_17652,N_14866,N_14693);
and U17653 (N_17653,N_14248,N_11140);
xnor U17654 (N_17654,N_11067,N_11299);
xor U17655 (N_17655,N_12966,N_11305);
xnor U17656 (N_17656,N_12605,N_12523);
nor U17657 (N_17657,N_11207,N_11655);
nand U17658 (N_17658,N_14184,N_10275);
and U17659 (N_17659,N_11548,N_13907);
nand U17660 (N_17660,N_10926,N_14542);
and U17661 (N_17661,N_10033,N_13811);
xor U17662 (N_17662,N_13319,N_12145);
and U17663 (N_17663,N_14435,N_10629);
or U17664 (N_17664,N_13266,N_12310);
nor U17665 (N_17665,N_13747,N_10876);
and U17666 (N_17666,N_10838,N_13147);
nand U17667 (N_17667,N_10283,N_12284);
and U17668 (N_17668,N_13844,N_13462);
nand U17669 (N_17669,N_14595,N_14810);
or U17670 (N_17670,N_14796,N_11410);
xor U17671 (N_17671,N_11894,N_12195);
nand U17672 (N_17672,N_12525,N_14942);
xor U17673 (N_17673,N_14475,N_13746);
nand U17674 (N_17674,N_11291,N_10326);
or U17675 (N_17675,N_13083,N_14939);
xor U17676 (N_17676,N_10910,N_12274);
or U17677 (N_17677,N_11860,N_11652);
nand U17678 (N_17678,N_13426,N_14870);
xor U17679 (N_17679,N_11850,N_14145);
xnor U17680 (N_17680,N_10157,N_12588);
nand U17681 (N_17681,N_10247,N_11463);
nor U17682 (N_17682,N_11955,N_10291);
xor U17683 (N_17683,N_14261,N_10815);
nand U17684 (N_17684,N_13261,N_13486);
xor U17685 (N_17685,N_14333,N_11289);
nand U17686 (N_17686,N_11918,N_12419);
and U17687 (N_17687,N_12230,N_12642);
or U17688 (N_17688,N_13896,N_10798);
nand U17689 (N_17689,N_13910,N_12543);
xor U17690 (N_17690,N_11474,N_13295);
xor U17691 (N_17691,N_12346,N_10202);
nor U17692 (N_17692,N_14320,N_13815);
and U17693 (N_17693,N_10183,N_10573);
or U17694 (N_17694,N_12405,N_13471);
or U17695 (N_17695,N_14054,N_11411);
xnor U17696 (N_17696,N_14177,N_14969);
or U17697 (N_17697,N_14540,N_13696);
and U17698 (N_17698,N_10814,N_12174);
nor U17699 (N_17699,N_11580,N_10793);
nand U17700 (N_17700,N_11528,N_14689);
nand U17701 (N_17701,N_12198,N_10207);
nor U17702 (N_17702,N_10531,N_10057);
xor U17703 (N_17703,N_10703,N_11497);
nand U17704 (N_17704,N_10905,N_13336);
xnor U17705 (N_17705,N_10903,N_12000);
nor U17706 (N_17706,N_14625,N_12165);
and U17707 (N_17707,N_12923,N_12293);
xnor U17708 (N_17708,N_13958,N_10382);
nand U17709 (N_17709,N_14004,N_11166);
and U17710 (N_17710,N_11718,N_14435);
xnor U17711 (N_17711,N_14506,N_10246);
nor U17712 (N_17712,N_11236,N_13180);
nand U17713 (N_17713,N_14749,N_12808);
or U17714 (N_17714,N_12559,N_10808);
nor U17715 (N_17715,N_11213,N_10390);
nand U17716 (N_17716,N_13932,N_10356);
or U17717 (N_17717,N_10229,N_10189);
xor U17718 (N_17718,N_11460,N_11022);
xor U17719 (N_17719,N_12596,N_12108);
xor U17720 (N_17720,N_14729,N_11438);
and U17721 (N_17721,N_10708,N_14274);
and U17722 (N_17722,N_12389,N_13306);
nand U17723 (N_17723,N_14816,N_10149);
xor U17724 (N_17724,N_11303,N_12688);
and U17725 (N_17725,N_14199,N_10922);
or U17726 (N_17726,N_12854,N_13708);
nor U17727 (N_17727,N_11136,N_11436);
nand U17728 (N_17728,N_12801,N_13184);
or U17729 (N_17729,N_14472,N_11361);
or U17730 (N_17730,N_10036,N_11787);
or U17731 (N_17731,N_14501,N_14626);
nand U17732 (N_17732,N_13131,N_10823);
and U17733 (N_17733,N_12048,N_12358);
nand U17734 (N_17734,N_11671,N_11101);
or U17735 (N_17735,N_12780,N_10297);
xor U17736 (N_17736,N_12091,N_10322);
and U17737 (N_17737,N_14017,N_11288);
xor U17738 (N_17738,N_12342,N_13733);
xor U17739 (N_17739,N_11617,N_10722);
xor U17740 (N_17740,N_13152,N_13250);
nand U17741 (N_17741,N_11961,N_11393);
nor U17742 (N_17742,N_11507,N_14186);
and U17743 (N_17743,N_10572,N_11338);
and U17744 (N_17744,N_13885,N_10550);
nor U17745 (N_17745,N_11626,N_14566);
nor U17746 (N_17746,N_13711,N_14779);
nor U17747 (N_17747,N_14603,N_11075);
nand U17748 (N_17748,N_14578,N_14115);
nor U17749 (N_17749,N_11868,N_10240);
nand U17750 (N_17750,N_12087,N_11765);
xnor U17751 (N_17751,N_11077,N_10170);
nor U17752 (N_17752,N_13521,N_12656);
nor U17753 (N_17753,N_11805,N_10395);
nor U17754 (N_17754,N_12944,N_10317);
and U17755 (N_17755,N_14145,N_11677);
xnor U17756 (N_17756,N_10832,N_11295);
nand U17757 (N_17757,N_12950,N_13590);
and U17758 (N_17758,N_14054,N_11494);
nand U17759 (N_17759,N_10755,N_10683);
and U17760 (N_17760,N_14977,N_11274);
xnor U17761 (N_17761,N_10876,N_12867);
xnor U17762 (N_17762,N_11104,N_14203);
xnor U17763 (N_17763,N_10437,N_13206);
and U17764 (N_17764,N_12486,N_11654);
nor U17765 (N_17765,N_14649,N_12707);
xnor U17766 (N_17766,N_12063,N_12184);
xnor U17767 (N_17767,N_11098,N_14472);
nand U17768 (N_17768,N_11334,N_12101);
nand U17769 (N_17769,N_10113,N_11975);
and U17770 (N_17770,N_11237,N_14745);
xor U17771 (N_17771,N_11960,N_10903);
nand U17772 (N_17772,N_11038,N_14858);
or U17773 (N_17773,N_11410,N_14458);
and U17774 (N_17774,N_14689,N_14407);
or U17775 (N_17775,N_14285,N_14235);
nor U17776 (N_17776,N_12537,N_14221);
nor U17777 (N_17777,N_14664,N_12020);
nand U17778 (N_17778,N_13938,N_11068);
or U17779 (N_17779,N_13320,N_14096);
and U17780 (N_17780,N_11267,N_14674);
nand U17781 (N_17781,N_13177,N_12952);
nand U17782 (N_17782,N_10136,N_10675);
xnor U17783 (N_17783,N_10332,N_12762);
and U17784 (N_17784,N_11259,N_10596);
and U17785 (N_17785,N_13997,N_12711);
xor U17786 (N_17786,N_11179,N_13134);
or U17787 (N_17787,N_12435,N_13436);
nor U17788 (N_17788,N_10651,N_14809);
xnor U17789 (N_17789,N_14054,N_11382);
and U17790 (N_17790,N_11929,N_14050);
nor U17791 (N_17791,N_10234,N_10133);
or U17792 (N_17792,N_13604,N_14054);
nand U17793 (N_17793,N_12076,N_13219);
xnor U17794 (N_17794,N_14694,N_14159);
xnor U17795 (N_17795,N_13555,N_12570);
and U17796 (N_17796,N_10711,N_13477);
nor U17797 (N_17797,N_12343,N_13544);
xnor U17798 (N_17798,N_10168,N_11276);
nand U17799 (N_17799,N_13477,N_11312);
or U17800 (N_17800,N_12253,N_12526);
nand U17801 (N_17801,N_13500,N_11799);
and U17802 (N_17802,N_10153,N_14539);
xor U17803 (N_17803,N_12184,N_10627);
or U17804 (N_17804,N_11822,N_14102);
xnor U17805 (N_17805,N_10917,N_11563);
nand U17806 (N_17806,N_11865,N_12184);
xor U17807 (N_17807,N_13708,N_10720);
nor U17808 (N_17808,N_10604,N_13454);
xor U17809 (N_17809,N_10714,N_11309);
xnor U17810 (N_17810,N_13528,N_10259);
and U17811 (N_17811,N_13553,N_10140);
or U17812 (N_17812,N_11051,N_10596);
nand U17813 (N_17813,N_11689,N_11717);
or U17814 (N_17814,N_12616,N_11730);
or U17815 (N_17815,N_10202,N_14012);
xor U17816 (N_17816,N_11897,N_11254);
nand U17817 (N_17817,N_13495,N_10029);
and U17818 (N_17818,N_10419,N_12514);
nand U17819 (N_17819,N_12351,N_12846);
and U17820 (N_17820,N_12425,N_14582);
nand U17821 (N_17821,N_10892,N_13485);
or U17822 (N_17822,N_10470,N_14980);
nor U17823 (N_17823,N_13827,N_11073);
nor U17824 (N_17824,N_10182,N_13387);
nand U17825 (N_17825,N_11759,N_14826);
xor U17826 (N_17826,N_10272,N_14729);
and U17827 (N_17827,N_13294,N_14523);
or U17828 (N_17828,N_10029,N_14960);
and U17829 (N_17829,N_10620,N_12919);
and U17830 (N_17830,N_10001,N_13257);
or U17831 (N_17831,N_14706,N_14967);
nor U17832 (N_17832,N_10308,N_12416);
or U17833 (N_17833,N_10582,N_11689);
xor U17834 (N_17834,N_13666,N_13750);
xor U17835 (N_17835,N_10197,N_10353);
nand U17836 (N_17836,N_13003,N_12109);
or U17837 (N_17837,N_11035,N_14928);
or U17838 (N_17838,N_10941,N_10431);
or U17839 (N_17839,N_12579,N_11431);
nor U17840 (N_17840,N_13294,N_10892);
xor U17841 (N_17841,N_11391,N_12327);
xnor U17842 (N_17842,N_10930,N_12848);
or U17843 (N_17843,N_12935,N_10245);
and U17844 (N_17844,N_11924,N_12343);
xor U17845 (N_17845,N_10769,N_13434);
xor U17846 (N_17846,N_10107,N_14890);
nand U17847 (N_17847,N_14591,N_14242);
or U17848 (N_17848,N_13507,N_12438);
nand U17849 (N_17849,N_11190,N_10335);
nor U17850 (N_17850,N_11629,N_14583);
nand U17851 (N_17851,N_10339,N_14069);
nor U17852 (N_17852,N_12518,N_10092);
and U17853 (N_17853,N_12709,N_10799);
and U17854 (N_17854,N_10677,N_11756);
or U17855 (N_17855,N_12444,N_14121);
or U17856 (N_17856,N_11584,N_14731);
or U17857 (N_17857,N_12156,N_14529);
nor U17858 (N_17858,N_12335,N_13149);
xor U17859 (N_17859,N_11785,N_14435);
or U17860 (N_17860,N_12300,N_11367);
and U17861 (N_17861,N_14761,N_10196);
nand U17862 (N_17862,N_14476,N_11752);
nand U17863 (N_17863,N_14436,N_11073);
and U17864 (N_17864,N_13043,N_11869);
nor U17865 (N_17865,N_13883,N_13158);
xnor U17866 (N_17866,N_11982,N_13974);
nor U17867 (N_17867,N_14713,N_10687);
nor U17868 (N_17868,N_14662,N_14496);
or U17869 (N_17869,N_14352,N_13037);
nor U17870 (N_17870,N_12939,N_13614);
nor U17871 (N_17871,N_13205,N_10056);
xor U17872 (N_17872,N_12574,N_13128);
xnor U17873 (N_17873,N_10704,N_13918);
nor U17874 (N_17874,N_14072,N_14261);
or U17875 (N_17875,N_13136,N_12904);
xnor U17876 (N_17876,N_10880,N_12481);
xor U17877 (N_17877,N_14010,N_11829);
and U17878 (N_17878,N_11682,N_14010);
nor U17879 (N_17879,N_12425,N_11376);
nor U17880 (N_17880,N_11419,N_11518);
and U17881 (N_17881,N_12777,N_14614);
xnor U17882 (N_17882,N_10134,N_13004);
xnor U17883 (N_17883,N_11293,N_14061);
nor U17884 (N_17884,N_13941,N_11764);
nor U17885 (N_17885,N_14176,N_12309);
xor U17886 (N_17886,N_14111,N_14975);
and U17887 (N_17887,N_13401,N_13342);
or U17888 (N_17888,N_12392,N_12848);
xnor U17889 (N_17889,N_13408,N_14467);
xnor U17890 (N_17890,N_12770,N_12938);
and U17891 (N_17891,N_12752,N_10740);
nor U17892 (N_17892,N_11673,N_10307);
or U17893 (N_17893,N_12521,N_10653);
nor U17894 (N_17894,N_13333,N_14210);
xor U17895 (N_17895,N_11640,N_12677);
xor U17896 (N_17896,N_14037,N_12673);
and U17897 (N_17897,N_10912,N_11218);
nand U17898 (N_17898,N_10561,N_14458);
nand U17899 (N_17899,N_10721,N_11657);
nor U17900 (N_17900,N_11426,N_11285);
nand U17901 (N_17901,N_14796,N_13090);
nand U17902 (N_17902,N_11036,N_10031);
or U17903 (N_17903,N_12232,N_11484);
nor U17904 (N_17904,N_11149,N_12101);
and U17905 (N_17905,N_10836,N_11765);
xnor U17906 (N_17906,N_14999,N_10232);
xor U17907 (N_17907,N_14429,N_12261);
nand U17908 (N_17908,N_10901,N_10241);
xnor U17909 (N_17909,N_10016,N_10943);
and U17910 (N_17910,N_13932,N_13545);
xor U17911 (N_17911,N_13341,N_11893);
or U17912 (N_17912,N_13425,N_10583);
xor U17913 (N_17913,N_13026,N_10952);
or U17914 (N_17914,N_14957,N_13607);
xor U17915 (N_17915,N_10130,N_10913);
or U17916 (N_17916,N_10073,N_13588);
nand U17917 (N_17917,N_10643,N_13736);
nor U17918 (N_17918,N_14754,N_10653);
nor U17919 (N_17919,N_13602,N_11037);
nand U17920 (N_17920,N_13289,N_11576);
nor U17921 (N_17921,N_14234,N_14449);
and U17922 (N_17922,N_11518,N_11358);
nand U17923 (N_17923,N_12539,N_14923);
nand U17924 (N_17924,N_13595,N_13228);
xnor U17925 (N_17925,N_11142,N_12667);
or U17926 (N_17926,N_13289,N_10452);
nand U17927 (N_17927,N_11919,N_11945);
xnor U17928 (N_17928,N_10932,N_12184);
or U17929 (N_17929,N_13099,N_12363);
nand U17930 (N_17930,N_11456,N_13369);
and U17931 (N_17931,N_14159,N_12718);
nor U17932 (N_17932,N_10783,N_10175);
and U17933 (N_17933,N_10197,N_10545);
or U17934 (N_17934,N_14021,N_12143);
and U17935 (N_17935,N_12476,N_11743);
and U17936 (N_17936,N_11897,N_10725);
xor U17937 (N_17937,N_12357,N_12479);
nand U17938 (N_17938,N_14096,N_10218);
or U17939 (N_17939,N_10950,N_14194);
nor U17940 (N_17940,N_11904,N_10983);
xnor U17941 (N_17941,N_13953,N_13521);
nor U17942 (N_17942,N_11595,N_14746);
xor U17943 (N_17943,N_10332,N_14301);
nor U17944 (N_17944,N_13969,N_12271);
xor U17945 (N_17945,N_12836,N_14681);
nand U17946 (N_17946,N_13322,N_13513);
nor U17947 (N_17947,N_13198,N_11360);
nand U17948 (N_17948,N_12242,N_13342);
and U17949 (N_17949,N_10386,N_13248);
xnor U17950 (N_17950,N_14650,N_12622);
nand U17951 (N_17951,N_12562,N_10445);
nor U17952 (N_17952,N_12706,N_11357);
and U17953 (N_17953,N_13275,N_10438);
xor U17954 (N_17954,N_14974,N_13998);
nand U17955 (N_17955,N_13554,N_14855);
xor U17956 (N_17956,N_14286,N_10886);
nor U17957 (N_17957,N_12626,N_11196);
xnor U17958 (N_17958,N_11329,N_13542);
xnor U17959 (N_17959,N_13434,N_12172);
and U17960 (N_17960,N_12065,N_13296);
nand U17961 (N_17961,N_12527,N_13301);
nor U17962 (N_17962,N_10730,N_12030);
xnor U17963 (N_17963,N_12788,N_10402);
xor U17964 (N_17964,N_11031,N_12382);
xor U17965 (N_17965,N_10459,N_12288);
nand U17966 (N_17966,N_13133,N_13875);
xnor U17967 (N_17967,N_13366,N_13873);
and U17968 (N_17968,N_12820,N_12883);
and U17969 (N_17969,N_12182,N_11716);
nor U17970 (N_17970,N_11064,N_13679);
and U17971 (N_17971,N_11461,N_10182);
or U17972 (N_17972,N_11172,N_10219);
nor U17973 (N_17973,N_11615,N_14592);
xor U17974 (N_17974,N_14713,N_10853);
or U17975 (N_17975,N_13342,N_13695);
nand U17976 (N_17976,N_10200,N_11915);
and U17977 (N_17977,N_13427,N_14578);
xnor U17978 (N_17978,N_13590,N_12587);
xor U17979 (N_17979,N_14755,N_11854);
or U17980 (N_17980,N_10094,N_10379);
xor U17981 (N_17981,N_14792,N_13532);
nor U17982 (N_17982,N_14998,N_12533);
xor U17983 (N_17983,N_10476,N_11336);
xor U17984 (N_17984,N_14446,N_10409);
and U17985 (N_17985,N_13122,N_12916);
or U17986 (N_17986,N_11488,N_12638);
and U17987 (N_17987,N_10138,N_13317);
nor U17988 (N_17988,N_14608,N_14828);
or U17989 (N_17989,N_10365,N_10446);
and U17990 (N_17990,N_10059,N_12994);
xor U17991 (N_17991,N_14058,N_10742);
nor U17992 (N_17992,N_10635,N_11703);
or U17993 (N_17993,N_13914,N_13026);
and U17994 (N_17994,N_11590,N_13750);
and U17995 (N_17995,N_12955,N_13874);
nor U17996 (N_17996,N_10087,N_11312);
xnor U17997 (N_17997,N_12774,N_12714);
and U17998 (N_17998,N_12581,N_12561);
nor U17999 (N_17999,N_12388,N_11988);
and U18000 (N_18000,N_10627,N_12580);
nand U18001 (N_18001,N_11550,N_13100);
nand U18002 (N_18002,N_14921,N_14606);
nor U18003 (N_18003,N_12851,N_13927);
nand U18004 (N_18004,N_13808,N_11564);
xor U18005 (N_18005,N_11557,N_11882);
nand U18006 (N_18006,N_10998,N_12548);
nand U18007 (N_18007,N_14406,N_10011);
or U18008 (N_18008,N_12545,N_11937);
nand U18009 (N_18009,N_11834,N_12988);
or U18010 (N_18010,N_14259,N_14850);
nand U18011 (N_18011,N_14039,N_14229);
nor U18012 (N_18012,N_12471,N_12270);
nor U18013 (N_18013,N_10904,N_13879);
nor U18014 (N_18014,N_13298,N_14184);
and U18015 (N_18015,N_10194,N_10450);
and U18016 (N_18016,N_14451,N_13597);
or U18017 (N_18017,N_11442,N_12897);
and U18018 (N_18018,N_14646,N_10367);
or U18019 (N_18019,N_11335,N_11232);
or U18020 (N_18020,N_12289,N_12797);
nor U18021 (N_18021,N_10011,N_14530);
nor U18022 (N_18022,N_14213,N_14682);
nand U18023 (N_18023,N_14000,N_11238);
xor U18024 (N_18024,N_10933,N_11366);
and U18025 (N_18025,N_11770,N_10818);
nor U18026 (N_18026,N_13073,N_13648);
nand U18027 (N_18027,N_12685,N_14190);
or U18028 (N_18028,N_10882,N_12269);
nor U18029 (N_18029,N_10620,N_13581);
nand U18030 (N_18030,N_14259,N_12010);
or U18031 (N_18031,N_14169,N_11610);
xor U18032 (N_18032,N_12087,N_11186);
nor U18033 (N_18033,N_13167,N_10128);
and U18034 (N_18034,N_10142,N_12965);
and U18035 (N_18035,N_14625,N_11445);
or U18036 (N_18036,N_14183,N_14537);
and U18037 (N_18037,N_13566,N_12091);
or U18038 (N_18038,N_11922,N_13955);
nand U18039 (N_18039,N_11040,N_13049);
or U18040 (N_18040,N_14873,N_13604);
xor U18041 (N_18041,N_14222,N_11107);
or U18042 (N_18042,N_13750,N_14250);
and U18043 (N_18043,N_12758,N_11418);
or U18044 (N_18044,N_11225,N_11712);
and U18045 (N_18045,N_13884,N_13130);
xnor U18046 (N_18046,N_13640,N_12020);
nand U18047 (N_18047,N_13348,N_11331);
nor U18048 (N_18048,N_11221,N_11305);
nor U18049 (N_18049,N_12125,N_12083);
xor U18050 (N_18050,N_11094,N_14499);
nand U18051 (N_18051,N_13742,N_11417);
or U18052 (N_18052,N_10571,N_13340);
and U18053 (N_18053,N_10202,N_14881);
or U18054 (N_18054,N_12033,N_12250);
xnor U18055 (N_18055,N_13077,N_12737);
nand U18056 (N_18056,N_12559,N_10393);
nor U18057 (N_18057,N_11618,N_10303);
nor U18058 (N_18058,N_13136,N_10413);
xor U18059 (N_18059,N_11938,N_14976);
or U18060 (N_18060,N_13491,N_12377);
xor U18061 (N_18061,N_11151,N_13217);
xor U18062 (N_18062,N_13173,N_10909);
nor U18063 (N_18063,N_12460,N_12771);
or U18064 (N_18064,N_10027,N_11835);
nor U18065 (N_18065,N_11897,N_11995);
and U18066 (N_18066,N_13069,N_10106);
or U18067 (N_18067,N_10538,N_10413);
nor U18068 (N_18068,N_13260,N_13858);
nand U18069 (N_18069,N_12483,N_11131);
or U18070 (N_18070,N_10425,N_12487);
nor U18071 (N_18071,N_10590,N_12823);
xor U18072 (N_18072,N_10137,N_12245);
xor U18073 (N_18073,N_12611,N_14327);
xor U18074 (N_18074,N_11531,N_12162);
xnor U18075 (N_18075,N_11325,N_13047);
and U18076 (N_18076,N_12638,N_11082);
nor U18077 (N_18077,N_14016,N_12035);
or U18078 (N_18078,N_10274,N_10734);
nor U18079 (N_18079,N_11437,N_12001);
or U18080 (N_18080,N_14696,N_13164);
or U18081 (N_18081,N_11536,N_11376);
nor U18082 (N_18082,N_14133,N_12668);
or U18083 (N_18083,N_13804,N_11573);
nor U18084 (N_18084,N_14969,N_11055);
nand U18085 (N_18085,N_14716,N_14974);
and U18086 (N_18086,N_13079,N_11076);
xnor U18087 (N_18087,N_12282,N_12082);
nand U18088 (N_18088,N_12984,N_14894);
nand U18089 (N_18089,N_11376,N_14713);
xnor U18090 (N_18090,N_10570,N_14883);
nor U18091 (N_18091,N_13318,N_10220);
or U18092 (N_18092,N_13814,N_13441);
or U18093 (N_18093,N_12497,N_12771);
or U18094 (N_18094,N_14541,N_13651);
nand U18095 (N_18095,N_10721,N_10192);
and U18096 (N_18096,N_13525,N_14209);
nor U18097 (N_18097,N_12945,N_11524);
nand U18098 (N_18098,N_13063,N_12821);
or U18099 (N_18099,N_13902,N_13711);
xor U18100 (N_18100,N_10720,N_13255);
and U18101 (N_18101,N_11830,N_11395);
or U18102 (N_18102,N_10288,N_12708);
nor U18103 (N_18103,N_14825,N_13084);
nor U18104 (N_18104,N_12760,N_13983);
nor U18105 (N_18105,N_12221,N_11361);
and U18106 (N_18106,N_11049,N_12000);
xnor U18107 (N_18107,N_10570,N_11140);
and U18108 (N_18108,N_10028,N_10897);
nand U18109 (N_18109,N_12374,N_11903);
nor U18110 (N_18110,N_14213,N_14729);
and U18111 (N_18111,N_13160,N_11630);
nand U18112 (N_18112,N_14090,N_14078);
nor U18113 (N_18113,N_14342,N_10910);
nor U18114 (N_18114,N_14106,N_14690);
xnor U18115 (N_18115,N_10596,N_13784);
or U18116 (N_18116,N_10938,N_14045);
xnor U18117 (N_18117,N_10864,N_10419);
nand U18118 (N_18118,N_14514,N_11739);
xnor U18119 (N_18119,N_10559,N_11023);
nand U18120 (N_18120,N_14821,N_10737);
or U18121 (N_18121,N_10533,N_14811);
nor U18122 (N_18122,N_11463,N_10473);
xnor U18123 (N_18123,N_12073,N_11157);
nor U18124 (N_18124,N_11311,N_12649);
and U18125 (N_18125,N_11959,N_10368);
xor U18126 (N_18126,N_10622,N_11513);
nand U18127 (N_18127,N_14838,N_14421);
nor U18128 (N_18128,N_13105,N_11514);
and U18129 (N_18129,N_13717,N_10275);
or U18130 (N_18130,N_13877,N_11731);
xnor U18131 (N_18131,N_10239,N_11331);
nand U18132 (N_18132,N_12034,N_14489);
or U18133 (N_18133,N_10102,N_12189);
nor U18134 (N_18134,N_13653,N_14811);
nand U18135 (N_18135,N_14682,N_14745);
xnor U18136 (N_18136,N_10500,N_12459);
xnor U18137 (N_18137,N_14242,N_12379);
nor U18138 (N_18138,N_13714,N_12699);
xnor U18139 (N_18139,N_12623,N_12578);
and U18140 (N_18140,N_13414,N_12084);
or U18141 (N_18141,N_12896,N_13510);
and U18142 (N_18142,N_12558,N_13577);
xor U18143 (N_18143,N_10066,N_10032);
and U18144 (N_18144,N_14596,N_12318);
nor U18145 (N_18145,N_11168,N_14168);
nor U18146 (N_18146,N_11770,N_13516);
nor U18147 (N_18147,N_13672,N_14068);
or U18148 (N_18148,N_13875,N_10022);
xnor U18149 (N_18149,N_13245,N_12127);
or U18150 (N_18150,N_11217,N_12166);
or U18151 (N_18151,N_13075,N_11101);
and U18152 (N_18152,N_11119,N_10762);
nor U18153 (N_18153,N_14700,N_14841);
and U18154 (N_18154,N_14808,N_10988);
nor U18155 (N_18155,N_13147,N_11947);
xor U18156 (N_18156,N_10949,N_11024);
xnor U18157 (N_18157,N_12860,N_14027);
and U18158 (N_18158,N_14849,N_11633);
and U18159 (N_18159,N_12409,N_13050);
nor U18160 (N_18160,N_12429,N_10767);
nand U18161 (N_18161,N_10009,N_10431);
or U18162 (N_18162,N_13734,N_11916);
nand U18163 (N_18163,N_13013,N_14956);
nor U18164 (N_18164,N_12048,N_12682);
xnor U18165 (N_18165,N_12351,N_14097);
xor U18166 (N_18166,N_13401,N_11019);
xnor U18167 (N_18167,N_14741,N_12124);
xor U18168 (N_18168,N_12084,N_10487);
or U18169 (N_18169,N_12203,N_13120);
and U18170 (N_18170,N_12013,N_13128);
xnor U18171 (N_18171,N_12807,N_11774);
nand U18172 (N_18172,N_10216,N_12974);
nor U18173 (N_18173,N_12784,N_14929);
and U18174 (N_18174,N_12618,N_12090);
xor U18175 (N_18175,N_10406,N_13321);
and U18176 (N_18176,N_14658,N_11255);
nor U18177 (N_18177,N_10652,N_11928);
xor U18178 (N_18178,N_12782,N_13672);
nand U18179 (N_18179,N_13733,N_13073);
xor U18180 (N_18180,N_12505,N_12318);
xnor U18181 (N_18181,N_10509,N_11381);
and U18182 (N_18182,N_13674,N_11139);
xor U18183 (N_18183,N_12489,N_14827);
or U18184 (N_18184,N_11332,N_10980);
nand U18185 (N_18185,N_10645,N_11527);
nor U18186 (N_18186,N_11962,N_11807);
nor U18187 (N_18187,N_13351,N_10917);
nand U18188 (N_18188,N_10114,N_13826);
and U18189 (N_18189,N_12175,N_11701);
and U18190 (N_18190,N_10336,N_10139);
nand U18191 (N_18191,N_13090,N_13125);
or U18192 (N_18192,N_12303,N_10147);
or U18193 (N_18193,N_11568,N_14073);
or U18194 (N_18194,N_14761,N_13559);
or U18195 (N_18195,N_13906,N_10782);
nand U18196 (N_18196,N_14843,N_12384);
nor U18197 (N_18197,N_13135,N_14996);
nand U18198 (N_18198,N_12943,N_12646);
nor U18199 (N_18199,N_14856,N_12736);
xnor U18200 (N_18200,N_14936,N_11316);
nor U18201 (N_18201,N_10965,N_13035);
nor U18202 (N_18202,N_14281,N_13857);
and U18203 (N_18203,N_14682,N_11784);
xnor U18204 (N_18204,N_10910,N_13006);
or U18205 (N_18205,N_11162,N_12799);
xor U18206 (N_18206,N_10356,N_11824);
xnor U18207 (N_18207,N_14734,N_14044);
xnor U18208 (N_18208,N_10625,N_13237);
nand U18209 (N_18209,N_14617,N_13190);
nand U18210 (N_18210,N_14995,N_12264);
nand U18211 (N_18211,N_12365,N_10887);
xnor U18212 (N_18212,N_10976,N_14590);
and U18213 (N_18213,N_10449,N_10923);
and U18214 (N_18214,N_14821,N_12372);
nand U18215 (N_18215,N_14616,N_11412);
xor U18216 (N_18216,N_11848,N_12904);
nand U18217 (N_18217,N_12628,N_12266);
and U18218 (N_18218,N_13324,N_12089);
nor U18219 (N_18219,N_14257,N_10689);
xor U18220 (N_18220,N_12365,N_14592);
nor U18221 (N_18221,N_10589,N_14105);
nor U18222 (N_18222,N_12827,N_14313);
xor U18223 (N_18223,N_11889,N_13967);
nor U18224 (N_18224,N_10336,N_10982);
and U18225 (N_18225,N_13219,N_13674);
nor U18226 (N_18226,N_14918,N_12896);
or U18227 (N_18227,N_14071,N_13393);
nand U18228 (N_18228,N_13340,N_13839);
or U18229 (N_18229,N_11315,N_11514);
or U18230 (N_18230,N_13575,N_13795);
or U18231 (N_18231,N_13365,N_12518);
nor U18232 (N_18232,N_14715,N_12964);
xor U18233 (N_18233,N_13317,N_14395);
or U18234 (N_18234,N_10848,N_10023);
nand U18235 (N_18235,N_12567,N_13739);
xor U18236 (N_18236,N_11136,N_12917);
xor U18237 (N_18237,N_11867,N_10189);
nor U18238 (N_18238,N_11394,N_12438);
nand U18239 (N_18239,N_10519,N_11494);
xor U18240 (N_18240,N_12066,N_10657);
or U18241 (N_18241,N_14645,N_12462);
nor U18242 (N_18242,N_10969,N_11073);
or U18243 (N_18243,N_13316,N_11976);
and U18244 (N_18244,N_11904,N_13691);
nand U18245 (N_18245,N_11634,N_13693);
or U18246 (N_18246,N_10770,N_12964);
or U18247 (N_18247,N_10817,N_12439);
nor U18248 (N_18248,N_12951,N_11388);
xnor U18249 (N_18249,N_11790,N_12392);
and U18250 (N_18250,N_13813,N_14905);
and U18251 (N_18251,N_13194,N_12312);
xnor U18252 (N_18252,N_11523,N_10701);
or U18253 (N_18253,N_13001,N_14759);
xnor U18254 (N_18254,N_10860,N_13333);
or U18255 (N_18255,N_13621,N_12856);
nand U18256 (N_18256,N_12729,N_10574);
and U18257 (N_18257,N_14448,N_14201);
xor U18258 (N_18258,N_12672,N_12947);
xnor U18259 (N_18259,N_12311,N_12739);
or U18260 (N_18260,N_10473,N_12991);
nor U18261 (N_18261,N_11864,N_11575);
and U18262 (N_18262,N_14665,N_11737);
nor U18263 (N_18263,N_11679,N_14459);
nor U18264 (N_18264,N_11034,N_10968);
xor U18265 (N_18265,N_14119,N_10414);
and U18266 (N_18266,N_14703,N_12805);
and U18267 (N_18267,N_11572,N_10755);
xor U18268 (N_18268,N_12203,N_13616);
and U18269 (N_18269,N_14591,N_10507);
and U18270 (N_18270,N_10889,N_10553);
nand U18271 (N_18271,N_13381,N_14664);
nor U18272 (N_18272,N_10806,N_14353);
or U18273 (N_18273,N_12180,N_12929);
nor U18274 (N_18274,N_11305,N_11386);
nand U18275 (N_18275,N_13794,N_11349);
xor U18276 (N_18276,N_12699,N_12624);
nand U18277 (N_18277,N_10888,N_14487);
and U18278 (N_18278,N_13864,N_12041);
xnor U18279 (N_18279,N_10522,N_13105);
xnor U18280 (N_18280,N_14720,N_12121);
nand U18281 (N_18281,N_10743,N_11501);
and U18282 (N_18282,N_13935,N_14220);
xor U18283 (N_18283,N_14368,N_10580);
or U18284 (N_18284,N_13160,N_11758);
and U18285 (N_18285,N_11704,N_13574);
nand U18286 (N_18286,N_11387,N_10425);
or U18287 (N_18287,N_14426,N_12968);
or U18288 (N_18288,N_10654,N_13840);
or U18289 (N_18289,N_12300,N_13500);
nand U18290 (N_18290,N_14532,N_11463);
xor U18291 (N_18291,N_13001,N_10902);
or U18292 (N_18292,N_14106,N_14651);
or U18293 (N_18293,N_11494,N_11600);
xnor U18294 (N_18294,N_11263,N_10449);
or U18295 (N_18295,N_14976,N_12334);
or U18296 (N_18296,N_10783,N_13155);
xnor U18297 (N_18297,N_12931,N_14102);
or U18298 (N_18298,N_10018,N_14106);
xnor U18299 (N_18299,N_14657,N_10907);
or U18300 (N_18300,N_12049,N_13764);
or U18301 (N_18301,N_14450,N_12486);
nor U18302 (N_18302,N_14116,N_11324);
and U18303 (N_18303,N_10113,N_10403);
nor U18304 (N_18304,N_12115,N_13490);
and U18305 (N_18305,N_13300,N_12054);
and U18306 (N_18306,N_10825,N_13981);
and U18307 (N_18307,N_10014,N_11927);
nand U18308 (N_18308,N_13195,N_14753);
nor U18309 (N_18309,N_14502,N_14555);
nor U18310 (N_18310,N_14450,N_10251);
nor U18311 (N_18311,N_11704,N_12139);
nor U18312 (N_18312,N_13523,N_12920);
xor U18313 (N_18313,N_13096,N_11479);
nor U18314 (N_18314,N_10143,N_13134);
or U18315 (N_18315,N_11891,N_11844);
nand U18316 (N_18316,N_10649,N_13609);
and U18317 (N_18317,N_14720,N_14920);
nor U18318 (N_18318,N_13261,N_10981);
xnor U18319 (N_18319,N_12385,N_11317);
or U18320 (N_18320,N_10935,N_10616);
and U18321 (N_18321,N_10569,N_11289);
and U18322 (N_18322,N_11054,N_12670);
xnor U18323 (N_18323,N_10570,N_12959);
and U18324 (N_18324,N_10733,N_13138);
xnor U18325 (N_18325,N_11531,N_12245);
and U18326 (N_18326,N_13844,N_13204);
nor U18327 (N_18327,N_12549,N_11573);
nor U18328 (N_18328,N_13004,N_12348);
and U18329 (N_18329,N_12222,N_10873);
xor U18330 (N_18330,N_11048,N_12983);
and U18331 (N_18331,N_11158,N_11884);
xnor U18332 (N_18332,N_13604,N_12735);
and U18333 (N_18333,N_12127,N_13717);
nand U18334 (N_18334,N_10427,N_14635);
and U18335 (N_18335,N_14631,N_12415);
nand U18336 (N_18336,N_12976,N_10126);
xor U18337 (N_18337,N_11361,N_10148);
nor U18338 (N_18338,N_12112,N_14449);
or U18339 (N_18339,N_10414,N_10590);
nand U18340 (N_18340,N_12116,N_13847);
nor U18341 (N_18341,N_14553,N_13834);
and U18342 (N_18342,N_13859,N_10991);
nand U18343 (N_18343,N_13868,N_10852);
nand U18344 (N_18344,N_10935,N_12342);
and U18345 (N_18345,N_14263,N_11415);
xnor U18346 (N_18346,N_13607,N_10427);
nor U18347 (N_18347,N_10058,N_11607);
and U18348 (N_18348,N_14138,N_11973);
and U18349 (N_18349,N_13680,N_14623);
or U18350 (N_18350,N_11757,N_14474);
or U18351 (N_18351,N_13994,N_13690);
or U18352 (N_18352,N_11487,N_14906);
and U18353 (N_18353,N_11811,N_11870);
or U18354 (N_18354,N_11055,N_10389);
or U18355 (N_18355,N_11491,N_13730);
or U18356 (N_18356,N_13946,N_13746);
nand U18357 (N_18357,N_12254,N_14415);
or U18358 (N_18358,N_11344,N_14406);
nor U18359 (N_18359,N_13993,N_12566);
nand U18360 (N_18360,N_13185,N_10493);
nor U18361 (N_18361,N_13361,N_11008);
nand U18362 (N_18362,N_14934,N_14619);
nor U18363 (N_18363,N_11582,N_12785);
nor U18364 (N_18364,N_14859,N_14561);
and U18365 (N_18365,N_11748,N_14442);
and U18366 (N_18366,N_11941,N_14905);
nand U18367 (N_18367,N_13012,N_12088);
and U18368 (N_18368,N_10268,N_10638);
xnor U18369 (N_18369,N_10623,N_12629);
xor U18370 (N_18370,N_14756,N_14333);
xnor U18371 (N_18371,N_10021,N_12563);
nand U18372 (N_18372,N_14897,N_13740);
nand U18373 (N_18373,N_10725,N_10480);
and U18374 (N_18374,N_12399,N_14436);
xnor U18375 (N_18375,N_14369,N_13136);
or U18376 (N_18376,N_11492,N_12790);
or U18377 (N_18377,N_10952,N_12463);
and U18378 (N_18378,N_12707,N_13513);
xnor U18379 (N_18379,N_14064,N_12263);
or U18380 (N_18380,N_14439,N_13597);
and U18381 (N_18381,N_13183,N_10872);
nor U18382 (N_18382,N_12810,N_13119);
and U18383 (N_18383,N_13967,N_14738);
xnor U18384 (N_18384,N_10434,N_10894);
or U18385 (N_18385,N_14140,N_10742);
and U18386 (N_18386,N_14078,N_12466);
nor U18387 (N_18387,N_13094,N_10591);
xnor U18388 (N_18388,N_14187,N_14527);
and U18389 (N_18389,N_11382,N_14305);
xor U18390 (N_18390,N_14578,N_11959);
nor U18391 (N_18391,N_11015,N_12641);
nor U18392 (N_18392,N_12119,N_14765);
nand U18393 (N_18393,N_14671,N_12378);
and U18394 (N_18394,N_11119,N_11089);
and U18395 (N_18395,N_13815,N_13046);
xnor U18396 (N_18396,N_13008,N_10539);
and U18397 (N_18397,N_11858,N_12828);
xor U18398 (N_18398,N_11154,N_14748);
or U18399 (N_18399,N_12447,N_13533);
xnor U18400 (N_18400,N_13246,N_10940);
xor U18401 (N_18401,N_10708,N_13885);
or U18402 (N_18402,N_10597,N_10440);
and U18403 (N_18403,N_12588,N_14950);
nor U18404 (N_18404,N_11309,N_10364);
or U18405 (N_18405,N_13263,N_10936);
nand U18406 (N_18406,N_10234,N_14281);
nor U18407 (N_18407,N_12765,N_10588);
xnor U18408 (N_18408,N_14229,N_12142);
or U18409 (N_18409,N_13847,N_11931);
nand U18410 (N_18410,N_12451,N_11745);
nor U18411 (N_18411,N_13237,N_12752);
or U18412 (N_18412,N_11830,N_14517);
or U18413 (N_18413,N_14512,N_11327);
nor U18414 (N_18414,N_12826,N_10157);
and U18415 (N_18415,N_10089,N_14633);
xnor U18416 (N_18416,N_12554,N_13069);
or U18417 (N_18417,N_11763,N_10488);
and U18418 (N_18418,N_14446,N_12015);
nor U18419 (N_18419,N_14356,N_13973);
nor U18420 (N_18420,N_12858,N_13301);
and U18421 (N_18421,N_14645,N_11303);
xnor U18422 (N_18422,N_13301,N_11417);
xnor U18423 (N_18423,N_12875,N_13379);
xnor U18424 (N_18424,N_11317,N_12960);
xor U18425 (N_18425,N_12619,N_13097);
xor U18426 (N_18426,N_11109,N_13021);
nor U18427 (N_18427,N_14967,N_10290);
or U18428 (N_18428,N_13947,N_10393);
nand U18429 (N_18429,N_11161,N_13614);
xor U18430 (N_18430,N_13435,N_13288);
xor U18431 (N_18431,N_10374,N_12272);
and U18432 (N_18432,N_12806,N_13216);
nand U18433 (N_18433,N_12587,N_10502);
and U18434 (N_18434,N_13355,N_10791);
nand U18435 (N_18435,N_11655,N_11469);
and U18436 (N_18436,N_14456,N_13399);
nand U18437 (N_18437,N_11572,N_10280);
nor U18438 (N_18438,N_13936,N_14457);
or U18439 (N_18439,N_13834,N_13986);
nand U18440 (N_18440,N_10206,N_12530);
and U18441 (N_18441,N_11589,N_11643);
nand U18442 (N_18442,N_12235,N_10750);
nor U18443 (N_18443,N_11625,N_10804);
nor U18444 (N_18444,N_10880,N_12434);
nand U18445 (N_18445,N_11457,N_13853);
or U18446 (N_18446,N_13027,N_10178);
nor U18447 (N_18447,N_11192,N_12646);
and U18448 (N_18448,N_13250,N_13510);
nor U18449 (N_18449,N_14747,N_13970);
xor U18450 (N_18450,N_14304,N_12239);
and U18451 (N_18451,N_11597,N_13917);
nor U18452 (N_18452,N_12248,N_12786);
nor U18453 (N_18453,N_14327,N_13022);
and U18454 (N_18454,N_10823,N_10585);
nor U18455 (N_18455,N_10425,N_10475);
xor U18456 (N_18456,N_14389,N_13792);
nand U18457 (N_18457,N_10274,N_13894);
nor U18458 (N_18458,N_10636,N_13464);
xor U18459 (N_18459,N_14672,N_13192);
and U18460 (N_18460,N_11605,N_14846);
and U18461 (N_18461,N_10742,N_11869);
or U18462 (N_18462,N_13989,N_13100);
or U18463 (N_18463,N_10468,N_11277);
nand U18464 (N_18464,N_11241,N_10588);
xor U18465 (N_18465,N_11504,N_13550);
or U18466 (N_18466,N_11020,N_11343);
nand U18467 (N_18467,N_11336,N_13449);
or U18468 (N_18468,N_12695,N_14159);
xnor U18469 (N_18469,N_13988,N_13803);
and U18470 (N_18470,N_13104,N_10326);
or U18471 (N_18471,N_14354,N_14634);
and U18472 (N_18472,N_11862,N_13539);
and U18473 (N_18473,N_10141,N_12397);
nor U18474 (N_18474,N_14788,N_13086);
xor U18475 (N_18475,N_10926,N_12873);
xor U18476 (N_18476,N_14383,N_14026);
nor U18477 (N_18477,N_10834,N_13502);
nor U18478 (N_18478,N_12383,N_12777);
and U18479 (N_18479,N_11649,N_10220);
xor U18480 (N_18480,N_14595,N_12122);
and U18481 (N_18481,N_10785,N_13028);
nor U18482 (N_18482,N_14865,N_10317);
xor U18483 (N_18483,N_14261,N_11425);
and U18484 (N_18484,N_12999,N_12358);
xor U18485 (N_18485,N_14879,N_14537);
nor U18486 (N_18486,N_10011,N_12518);
or U18487 (N_18487,N_13799,N_14122);
and U18488 (N_18488,N_12358,N_11830);
nand U18489 (N_18489,N_14434,N_11050);
or U18490 (N_18490,N_14873,N_12976);
xnor U18491 (N_18491,N_12152,N_13733);
and U18492 (N_18492,N_14851,N_11387);
nand U18493 (N_18493,N_14547,N_13214);
or U18494 (N_18494,N_10085,N_10552);
or U18495 (N_18495,N_10695,N_12268);
or U18496 (N_18496,N_14887,N_10725);
xnor U18497 (N_18497,N_13192,N_10241);
nand U18498 (N_18498,N_13172,N_10107);
nand U18499 (N_18499,N_12031,N_11622);
nor U18500 (N_18500,N_13599,N_11461);
nor U18501 (N_18501,N_11308,N_10233);
xor U18502 (N_18502,N_11150,N_11749);
and U18503 (N_18503,N_13409,N_13582);
or U18504 (N_18504,N_12526,N_10167);
nand U18505 (N_18505,N_14861,N_10667);
xor U18506 (N_18506,N_10937,N_14724);
nand U18507 (N_18507,N_12130,N_11047);
xnor U18508 (N_18508,N_14181,N_11598);
and U18509 (N_18509,N_11672,N_10902);
nand U18510 (N_18510,N_10374,N_12515);
nand U18511 (N_18511,N_10320,N_14674);
nand U18512 (N_18512,N_14960,N_14520);
xor U18513 (N_18513,N_14991,N_13199);
nand U18514 (N_18514,N_11685,N_11551);
nand U18515 (N_18515,N_11883,N_10886);
or U18516 (N_18516,N_12219,N_12056);
nor U18517 (N_18517,N_12217,N_14177);
nand U18518 (N_18518,N_12182,N_10132);
or U18519 (N_18519,N_14557,N_10372);
nand U18520 (N_18520,N_12203,N_11795);
nand U18521 (N_18521,N_13158,N_13575);
or U18522 (N_18522,N_10545,N_13204);
or U18523 (N_18523,N_10344,N_10215);
or U18524 (N_18524,N_14641,N_10264);
xnor U18525 (N_18525,N_12362,N_14627);
nor U18526 (N_18526,N_12641,N_11610);
xor U18527 (N_18527,N_10566,N_14188);
and U18528 (N_18528,N_13644,N_14159);
and U18529 (N_18529,N_13104,N_14276);
and U18530 (N_18530,N_11976,N_13192);
nor U18531 (N_18531,N_14966,N_11816);
or U18532 (N_18532,N_12269,N_11848);
nand U18533 (N_18533,N_10083,N_14609);
and U18534 (N_18534,N_10645,N_12634);
or U18535 (N_18535,N_10400,N_12879);
nor U18536 (N_18536,N_10739,N_13802);
and U18537 (N_18537,N_12809,N_13254);
nor U18538 (N_18538,N_12389,N_11481);
xnor U18539 (N_18539,N_11236,N_12754);
nand U18540 (N_18540,N_11043,N_10922);
or U18541 (N_18541,N_11102,N_13248);
or U18542 (N_18542,N_14286,N_11426);
xnor U18543 (N_18543,N_10279,N_10540);
nand U18544 (N_18544,N_14567,N_10991);
nand U18545 (N_18545,N_12169,N_12498);
nor U18546 (N_18546,N_12862,N_11414);
and U18547 (N_18547,N_11010,N_10139);
and U18548 (N_18548,N_12325,N_13314);
xnor U18549 (N_18549,N_10451,N_14785);
nand U18550 (N_18550,N_14659,N_10793);
xnor U18551 (N_18551,N_13423,N_10826);
nor U18552 (N_18552,N_13528,N_11725);
nand U18553 (N_18553,N_13629,N_13989);
and U18554 (N_18554,N_12558,N_14635);
or U18555 (N_18555,N_14995,N_13516);
and U18556 (N_18556,N_12910,N_13435);
or U18557 (N_18557,N_10857,N_12434);
nor U18558 (N_18558,N_13541,N_10625);
or U18559 (N_18559,N_14720,N_12725);
nand U18560 (N_18560,N_12064,N_14846);
and U18561 (N_18561,N_10988,N_10629);
nand U18562 (N_18562,N_11369,N_14002);
nand U18563 (N_18563,N_11580,N_13581);
nand U18564 (N_18564,N_10131,N_12362);
or U18565 (N_18565,N_13816,N_10943);
nand U18566 (N_18566,N_14421,N_14916);
nor U18567 (N_18567,N_10739,N_14866);
nand U18568 (N_18568,N_11929,N_10346);
nand U18569 (N_18569,N_14805,N_14032);
xnor U18570 (N_18570,N_11016,N_10053);
or U18571 (N_18571,N_14675,N_13774);
xnor U18572 (N_18572,N_14944,N_13877);
xor U18573 (N_18573,N_14553,N_14311);
nand U18574 (N_18574,N_11012,N_12286);
nor U18575 (N_18575,N_12516,N_12164);
nand U18576 (N_18576,N_13603,N_12291);
nor U18577 (N_18577,N_12893,N_14168);
or U18578 (N_18578,N_14737,N_12778);
nor U18579 (N_18579,N_14880,N_13422);
xnor U18580 (N_18580,N_14765,N_14365);
nand U18581 (N_18581,N_13436,N_13470);
nand U18582 (N_18582,N_12498,N_11933);
nor U18583 (N_18583,N_12285,N_14103);
and U18584 (N_18584,N_11571,N_13551);
nor U18585 (N_18585,N_11232,N_13818);
or U18586 (N_18586,N_12872,N_12095);
and U18587 (N_18587,N_12049,N_13840);
xnor U18588 (N_18588,N_13593,N_14397);
and U18589 (N_18589,N_11125,N_12813);
and U18590 (N_18590,N_10339,N_14855);
or U18591 (N_18591,N_12737,N_14062);
nand U18592 (N_18592,N_10741,N_10029);
or U18593 (N_18593,N_10405,N_13907);
nand U18594 (N_18594,N_12216,N_11491);
nor U18595 (N_18595,N_11102,N_11133);
xnor U18596 (N_18596,N_13304,N_10423);
nor U18597 (N_18597,N_11508,N_12661);
xnor U18598 (N_18598,N_11651,N_10993);
nor U18599 (N_18599,N_14071,N_14709);
nor U18600 (N_18600,N_12005,N_13766);
or U18601 (N_18601,N_14703,N_12268);
and U18602 (N_18602,N_10597,N_13157);
and U18603 (N_18603,N_14590,N_14448);
nand U18604 (N_18604,N_13000,N_14783);
and U18605 (N_18605,N_11824,N_14592);
and U18606 (N_18606,N_11122,N_10938);
and U18607 (N_18607,N_12864,N_12675);
and U18608 (N_18608,N_14557,N_14157);
or U18609 (N_18609,N_13434,N_11547);
nand U18610 (N_18610,N_14997,N_14803);
and U18611 (N_18611,N_10499,N_10909);
and U18612 (N_18612,N_11844,N_10972);
nor U18613 (N_18613,N_11168,N_14174);
nor U18614 (N_18614,N_11716,N_14117);
nor U18615 (N_18615,N_12583,N_13101);
and U18616 (N_18616,N_11375,N_14843);
nand U18617 (N_18617,N_10415,N_10273);
xor U18618 (N_18618,N_12281,N_14270);
nand U18619 (N_18619,N_10718,N_11797);
or U18620 (N_18620,N_14590,N_13614);
and U18621 (N_18621,N_14983,N_10817);
and U18622 (N_18622,N_12679,N_13894);
or U18623 (N_18623,N_12474,N_11936);
nor U18624 (N_18624,N_14990,N_12170);
nor U18625 (N_18625,N_10323,N_13731);
nor U18626 (N_18626,N_12111,N_13620);
nor U18627 (N_18627,N_14790,N_10345);
xnor U18628 (N_18628,N_11441,N_13418);
or U18629 (N_18629,N_10737,N_11175);
xnor U18630 (N_18630,N_11117,N_12146);
xor U18631 (N_18631,N_14007,N_11014);
xor U18632 (N_18632,N_12304,N_13373);
nor U18633 (N_18633,N_10910,N_14538);
nor U18634 (N_18634,N_14164,N_10272);
nor U18635 (N_18635,N_10504,N_14901);
or U18636 (N_18636,N_10812,N_12153);
nor U18637 (N_18637,N_13726,N_10748);
nand U18638 (N_18638,N_13356,N_12222);
xnor U18639 (N_18639,N_13399,N_12390);
nand U18640 (N_18640,N_10211,N_14829);
and U18641 (N_18641,N_13172,N_11386);
or U18642 (N_18642,N_11182,N_12968);
or U18643 (N_18643,N_10473,N_11703);
nand U18644 (N_18644,N_12613,N_10509);
nand U18645 (N_18645,N_12877,N_10935);
and U18646 (N_18646,N_10541,N_11334);
nand U18647 (N_18647,N_12312,N_14399);
nand U18648 (N_18648,N_13958,N_11171);
nand U18649 (N_18649,N_13573,N_14301);
and U18650 (N_18650,N_13163,N_11464);
nor U18651 (N_18651,N_14886,N_13876);
and U18652 (N_18652,N_11493,N_11764);
and U18653 (N_18653,N_10739,N_12886);
nand U18654 (N_18654,N_14152,N_13116);
xnor U18655 (N_18655,N_13602,N_10451);
or U18656 (N_18656,N_11338,N_13787);
nand U18657 (N_18657,N_12584,N_14149);
and U18658 (N_18658,N_11443,N_12730);
and U18659 (N_18659,N_13665,N_10285);
nand U18660 (N_18660,N_11025,N_13358);
nor U18661 (N_18661,N_12223,N_13817);
nor U18662 (N_18662,N_13616,N_14313);
nand U18663 (N_18663,N_14447,N_10058);
and U18664 (N_18664,N_11426,N_11350);
nand U18665 (N_18665,N_13218,N_14777);
nor U18666 (N_18666,N_12057,N_13836);
xnor U18667 (N_18667,N_13274,N_10308);
and U18668 (N_18668,N_10587,N_14749);
nand U18669 (N_18669,N_11782,N_13741);
nand U18670 (N_18670,N_11219,N_11553);
xnor U18671 (N_18671,N_12159,N_12585);
or U18672 (N_18672,N_11084,N_12787);
xor U18673 (N_18673,N_14349,N_10667);
nand U18674 (N_18674,N_12374,N_12707);
and U18675 (N_18675,N_11650,N_14047);
and U18676 (N_18676,N_14223,N_10871);
nor U18677 (N_18677,N_12761,N_13388);
nand U18678 (N_18678,N_11378,N_12315);
xnor U18679 (N_18679,N_12203,N_11602);
xor U18680 (N_18680,N_11421,N_14925);
and U18681 (N_18681,N_12213,N_14797);
nor U18682 (N_18682,N_10322,N_14351);
or U18683 (N_18683,N_13642,N_14117);
nor U18684 (N_18684,N_14244,N_11890);
nor U18685 (N_18685,N_13199,N_11515);
nor U18686 (N_18686,N_13571,N_13369);
nand U18687 (N_18687,N_14644,N_13059);
nor U18688 (N_18688,N_12670,N_10661);
and U18689 (N_18689,N_11265,N_11217);
nand U18690 (N_18690,N_10682,N_14882);
or U18691 (N_18691,N_10720,N_11275);
nor U18692 (N_18692,N_11289,N_10097);
nor U18693 (N_18693,N_13495,N_11305);
xnor U18694 (N_18694,N_10377,N_12186);
nand U18695 (N_18695,N_11603,N_14866);
xor U18696 (N_18696,N_14768,N_12264);
nand U18697 (N_18697,N_12399,N_10293);
xor U18698 (N_18698,N_12492,N_13944);
and U18699 (N_18699,N_10275,N_14172);
and U18700 (N_18700,N_14390,N_13177);
nor U18701 (N_18701,N_13443,N_13154);
and U18702 (N_18702,N_14723,N_10777);
or U18703 (N_18703,N_10946,N_10298);
nand U18704 (N_18704,N_10820,N_10805);
or U18705 (N_18705,N_10472,N_12287);
and U18706 (N_18706,N_14324,N_10615);
nand U18707 (N_18707,N_14900,N_12338);
nand U18708 (N_18708,N_10836,N_10725);
and U18709 (N_18709,N_11158,N_14673);
nor U18710 (N_18710,N_14021,N_14507);
nand U18711 (N_18711,N_10716,N_14335);
and U18712 (N_18712,N_13404,N_10856);
nand U18713 (N_18713,N_14374,N_13631);
nand U18714 (N_18714,N_14081,N_10865);
and U18715 (N_18715,N_14449,N_14907);
or U18716 (N_18716,N_13988,N_12611);
and U18717 (N_18717,N_14427,N_11192);
or U18718 (N_18718,N_11702,N_12442);
and U18719 (N_18719,N_11044,N_14192);
and U18720 (N_18720,N_13594,N_14768);
nor U18721 (N_18721,N_11617,N_10765);
nor U18722 (N_18722,N_10678,N_14229);
nand U18723 (N_18723,N_13004,N_14407);
and U18724 (N_18724,N_12857,N_11185);
or U18725 (N_18725,N_10247,N_12176);
xnor U18726 (N_18726,N_14754,N_11995);
or U18727 (N_18727,N_10703,N_14934);
xor U18728 (N_18728,N_12448,N_10025);
and U18729 (N_18729,N_14969,N_11214);
or U18730 (N_18730,N_13848,N_14269);
and U18731 (N_18731,N_11307,N_10061);
or U18732 (N_18732,N_10340,N_12572);
nor U18733 (N_18733,N_14600,N_14813);
or U18734 (N_18734,N_12085,N_11088);
or U18735 (N_18735,N_12609,N_13264);
and U18736 (N_18736,N_13128,N_13546);
nor U18737 (N_18737,N_11392,N_10288);
nor U18738 (N_18738,N_10189,N_13595);
nand U18739 (N_18739,N_13334,N_13845);
nor U18740 (N_18740,N_13724,N_13163);
nand U18741 (N_18741,N_12149,N_10342);
and U18742 (N_18742,N_12403,N_12450);
or U18743 (N_18743,N_13702,N_14277);
and U18744 (N_18744,N_14324,N_10880);
nand U18745 (N_18745,N_13840,N_10939);
nand U18746 (N_18746,N_13233,N_10330);
nand U18747 (N_18747,N_14920,N_11764);
xnor U18748 (N_18748,N_12039,N_10286);
xor U18749 (N_18749,N_10529,N_13859);
xor U18750 (N_18750,N_11159,N_12994);
or U18751 (N_18751,N_11121,N_10461);
xnor U18752 (N_18752,N_11441,N_10944);
nor U18753 (N_18753,N_10383,N_12635);
or U18754 (N_18754,N_11378,N_13930);
and U18755 (N_18755,N_13518,N_13954);
nand U18756 (N_18756,N_12684,N_14991);
nor U18757 (N_18757,N_11746,N_13978);
xnor U18758 (N_18758,N_11732,N_14191);
nand U18759 (N_18759,N_11741,N_12219);
or U18760 (N_18760,N_13654,N_13079);
xnor U18761 (N_18761,N_13828,N_12754);
nand U18762 (N_18762,N_10394,N_13016);
or U18763 (N_18763,N_12278,N_11956);
nand U18764 (N_18764,N_13939,N_12472);
nand U18765 (N_18765,N_14669,N_14272);
nor U18766 (N_18766,N_11418,N_12144);
or U18767 (N_18767,N_12460,N_13326);
nor U18768 (N_18768,N_12020,N_14051);
nand U18769 (N_18769,N_12001,N_14058);
xor U18770 (N_18770,N_13198,N_10680);
or U18771 (N_18771,N_12554,N_14478);
and U18772 (N_18772,N_11691,N_10617);
or U18773 (N_18773,N_11211,N_14357);
nand U18774 (N_18774,N_10411,N_14503);
nor U18775 (N_18775,N_13928,N_13087);
and U18776 (N_18776,N_11023,N_10215);
nor U18777 (N_18777,N_12975,N_12804);
nand U18778 (N_18778,N_12483,N_13152);
and U18779 (N_18779,N_13523,N_12438);
or U18780 (N_18780,N_13609,N_13489);
nand U18781 (N_18781,N_11081,N_13466);
or U18782 (N_18782,N_12476,N_11838);
xnor U18783 (N_18783,N_14428,N_14015);
nand U18784 (N_18784,N_14512,N_13751);
and U18785 (N_18785,N_11252,N_14432);
or U18786 (N_18786,N_10294,N_10431);
or U18787 (N_18787,N_10892,N_14268);
and U18788 (N_18788,N_13296,N_13727);
xor U18789 (N_18789,N_14775,N_14732);
nand U18790 (N_18790,N_11498,N_11976);
nor U18791 (N_18791,N_13398,N_14598);
and U18792 (N_18792,N_13803,N_14839);
or U18793 (N_18793,N_11462,N_12445);
nor U18794 (N_18794,N_10897,N_13253);
xor U18795 (N_18795,N_14302,N_13692);
or U18796 (N_18796,N_11099,N_10308);
nor U18797 (N_18797,N_12357,N_11757);
nand U18798 (N_18798,N_12429,N_12981);
and U18799 (N_18799,N_12682,N_12937);
nand U18800 (N_18800,N_13300,N_13317);
xor U18801 (N_18801,N_14327,N_13766);
xor U18802 (N_18802,N_10407,N_14686);
nor U18803 (N_18803,N_14275,N_14368);
nand U18804 (N_18804,N_14899,N_11479);
nand U18805 (N_18805,N_14262,N_12159);
nand U18806 (N_18806,N_13899,N_13831);
nand U18807 (N_18807,N_11147,N_11203);
xnor U18808 (N_18808,N_12226,N_13343);
xor U18809 (N_18809,N_10011,N_10906);
or U18810 (N_18810,N_12414,N_13780);
xnor U18811 (N_18811,N_14944,N_12041);
nor U18812 (N_18812,N_14041,N_13271);
and U18813 (N_18813,N_11123,N_12909);
and U18814 (N_18814,N_12774,N_13438);
or U18815 (N_18815,N_10620,N_13534);
and U18816 (N_18816,N_14717,N_13011);
nand U18817 (N_18817,N_14647,N_13550);
xnor U18818 (N_18818,N_13933,N_14109);
or U18819 (N_18819,N_11051,N_11211);
xor U18820 (N_18820,N_13224,N_10525);
xnor U18821 (N_18821,N_14902,N_10877);
nor U18822 (N_18822,N_11587,N_12826);
xor U18823 (N_18823,N_12339,N_11513);
and U18824 (N_18824,N_11839,N_14524);
and U18825 (N_18825,N_12301,N_14569);
or U18826 (N_18826,N_12052,N_12935);
xor U18827 (N_18827,N_10415,N_14062);
nor U18828 (N_18828,N_13555,N_11246);
and U18829 (N_18829,N_12891,N_10321);
or U18830 (N_18830,N_12758,N_13903);
or U18831 (N_18831,N_11975,N_11063);
xor U18832 (N_18832,N_13436,N_13208);
xor U18833 (N_18833,N_11296,N_13859);
xnor U18834 (N_18834,N_12104,N_10448);
and U18835 (N_18835,N_14228,N_13099);
and U18836 (N_18836,N_10366,N_13498);
and U18837 (N_18837,N_12293,N_13958);
nand U18838 (N_18838,N_14573,N_11615);
nand U18839 (N_18839,N_10290,N_11010);
nand U18840 (N_18840,N_12095,N_10824);
nand U18841 (N_18841,N_13671,N_14107);
xnor U18842 (N_18842,N_14846,N_11054);
nor U18843 (N_18843,N_13905,N_10538);
or U18844 (N_18844,N_14429,N_12017);
xor U18845 (N_18845,N_12764,N_10401);
or U18846 (N_18846,N_13194,N_14685);
nor U18847 (N_18847,N_12249,N_13471);
nor U18848 (N_18848,N_13861,N_13134);
nand U18849 (N_18849,N_13819,N_14592);
nand U18850 (N_18850,N_11027,N_10706);
xor U18851 (N_18851,N_12587,N_14864);
nand U18852 (N_18852,N_10326,N_10923);
and U18853 (N_18853,N_14499,N_14218);
xor U18854 (N_18854,N_14709,N_11782);
xnor U18855 (N_18855,N_10207,N_11935);
and U18856 (N_18856,N_14117,N_12872);
nand U18857 (N_18857,N_10526,N_10752);
nor U18858 (N_18858,N_13843,N_11835);
and U18859 (N_18859,N_10023,N_14507);
nor U18860 (N_18860,N_13890,N_11572);
nor U18861 (N_18861,N_12695,N_12105);
nor U18862 (N_18862,N_10453,N_12357);
nand U18863 (N_18863,N_14034,N_14226);
and U18864 (N_18864,N_14049,N_12748);
nand U18865 (N_18865,N_14628,N_13780);
or U18866 (N_18866,N_12305,N_10347);
and U18867 (N_18867,N_14223,N_14925);
xnor U18868 (N_18868,N_14631,N_11546);
or U18869 (N_18869,N_10731,N_13060);
xnor U18870 (N_18870,N_13574,N_12315);
nor U18871 (N_18871,N_12518,N_14779);
or U18872 (N_18872,N_12389,N_10753);
xnor U18873 (N_18873,N_12350,N_12019);
and U18874 (N_18874,N_13325,N_10469);
or U18875 (N_18875,N_10812,N_10781);
nor U18876 (N_18876,N_14451,N_10051);
or U18877 (N_18877,N_11049,N_12678);
and U18878 (N_18878,N_12710,N_10417);
xor U18879 (N_18879,N_12470,N_14199);
or U18880 (N_18880,N_11295,N_11504);
nand U18881 (N_18881,N_13627,N_11426);
and U18882 (N_18882,N_10881,N_10720);
nand U18883 (N_18883,N_11150,N_13054);
nor U18884 (N_18884,N_13492,N_14348);
xnor U18885 (N_18885,N_11843,N_11490);
and U18886 (N_18886,N_13231,N_10316);
or U18887 (N_18887,N_12735,N_12233);
and U18888 (N_18888,N_11360,N_12732);
nor U18889 (N_18889,N_11343,N_11932);
nor U18890 (N_18890,N_13129,N_11966);
nor U18891 (N_18891,N_14510,N_12454);
nor U18892 (N_18892,N_11687,N_12341);
and U18893 (N_18893,N_11037,N_10587);
and U18894 (N_18894,N_11467,N_11144);
and U18895 (N_18895,N_14636,N_10228);
xor U18896 (N_18896,N_10384,N_10078);
xor U18897 (N_18897,N_11095,N_14010);
nand U18898 (N_18898,N_12384,N_14948);
nand U18899 (N_18899,N_11078,N_11937);
or U18900 (N_18900,N_14889,N_12558);
and U18901 (N_18901,N_11681,N_13159);
or U18902 (N_18902,N_14599,N_11164);
and U18903 (N_18903,N_12516,N_10267);
nand U18904 (N_18904,N_13674,N_12878);
xor U18905 (N_18905,N_11677,N_10312);
nand U18906 (N_18906,N_11461,N_14794);
or U18907 (N_18907,N_11999,N_10192);
and U18908 (N_18908,N_13117,N_13126);
xor U18909 (N_18909,N_10542,N_13800);
nand U18910 (N_18910,N_12126,N_13764);
and U18911 (N_18911,N_10958,N_11744);
xor U18912 (N_18912,N_11591,N_10842);
or U18913 (N_18913,N_12943,N_10722);
or U18914 (N_18914,N_11691,N_13941);
and U18915 (N_18915,N_10645,N_10330);
and U18916 (N_18916,N_13134,N_11879);
xor U18917 (N_18917,N_14507,N_12611);
or U18918 (N_18918,N_11823,N_11498);
xor U18919 (N_18919,N_11988,N_11238);
nand U18920 (N_18920,N_14177,N_12831);
nand U18921 (N_18921,N_11662,N_12307);
or U18922 (N_18922,N_12511,N_13992);
or U18923 (N_18923,N_10172,N_13254);
and U18924 (N_18924,N_10566,N_10501);
xnor U18925 (N_18925,N_12680,N_13195);
and U18926 (N_18926,N_13325,N_14846);
or U18927 (N_18927,N_11230,N_11116);
nand U18928 (N_18928,N_12401,N_14198);
and U18929 (N_18929,N_10726,N_13045);
or U18930 (N_18930,N_10115,N_14243);
nand U18931 (N_18931,N_13348,N_11606);
xor U18932 (N_18932,N_10748,N_11810);
nand U18933 (N_18933,N_12728,N_13100);
and U18934 (N_18934,N_10293,N_10278);
nor U18935 (N_18935,N_12679,N_13248);
nand U18936 (N_18936,N_12702,N_13212);
or U18937 (N_18937,N_12015,N_13095);
nor U18938 (N_18938,N_10150,N_12583);
nand U18939 (N_18939,N_13378,N_11711);
nand U18940 (N_18940,N_10822,N_14763);
and U18941 (N_18941,N_14461,N_10670);
and U18942 (N_18942,N_10898,N_11306);
or U18943 (N_18943,N_10347,N_11601);
and U18944 (N_18944,N_14989,N_12039);
or U18945 (N_18945,N_14748,N_13488);
xnor U18946 (N_18946,N_13746,N_13433);
nor U18947 (N_18947,N_14427,N_10577);
nor U18948 (N_18948,N_14569,N_13514);
nand U18949 (N_18949,N_12054,N_10865);
nor U18950 (N_18950,N_11425,N_14340);
or U18951 (N_18951,N_11578,N_11834);
nand U18952 (N_18952,N_13276,N_11323);
and U18953 (N_18953,N_10097,N_10190);
and U18954 (N_18954,N_14022,N_11926);
or U18955 (N_18955,N_12309,N_12386);
or U18956 (N_18956,N_12164,N_14830);
and U18957 (N_18957,N_13511,N_14375);
or U18958 (N_18958,N_11739,N_12147);
xnor U18959 (N_18959,N_13080,N_14328);
or U18960 (N_18960,N_13333,N_13864);
and U18961 (N_18961,N_12099,N_12959);
nand U18962 (N_18962,N_13486,N_13254);
nor U18963 (N_18963,N_12817,N_10429);
or U18964 (N_18964,N_12698,N_10349);
xor U18965 (N_18965,N_11822,N_13713);
nor U18966 (N_18966,N_14113,N_14700);
and U18967 (N_18967,N_13711,N_14784);
xnor U18968 (N_18968,N_12997,N_12844);
and U18969 (N_18969,N_14388,N_14718);
xnor U18970 (N_18970,N_11049,N_13565);
nor U18971 (N_18971,N_11784,N_11111);
nor U18972 (N_18972,N_14060,N_13577);
xnor U18973 (N_18973,N_12176,N_12105);
xnor U18974 (N_18974,N_13019,N_13528);
nand U18975 (N_18975,N_12508,N_13599);
and U18976 (N_18976,N_14253,N_14013);
nand U18977 (N_18977,N_14994,N_10363);
xor U18978 (N_18978,N_14271,N_13800);
nand U18979 (N_18979,N_13436,N_14647);
and U18980 (N_18980,N_13441,N_12192);
nor U18981 (N_18981,N_12038,N_10400);
or U18982 (N_18982,N_13330,N_12451);
and U18983 (N_18983,N_13273,N_11363);
nor U18984 (N_18984,N_13060,N_13093);
xor U18985 (N_18985,N_13262,N_14848);
or U18986 (N_18986,N_14962,N_10822);
nor U18987 (N_18987,N_10987,N_12109);
xnor U18988 (N_18988,N_11764,N_12663);
or U18989 (N_18989,N_11623,N_10366);
xor U18990 (N_18990,N_11502,N_11748);
and U18991 (N_18991,N_10692,N_12761);
and U18992 (N_18992,N_13436,N_11315);
nand U18993 (N_18993,N_10037,N_12230);
nand U18994 (N_18994,N_11470,N_13321);
and U18995 (N_18995,N_11406,N_12002);
nand U18996 (N_18996,N_11293,N_13967);
nand U18997 (N_18997,N_12725,N_12108);
xor U18998 (N_18998,N_10809,N_14061);
nor U18999 (N_18999,N_14173,N_11378);
nor U19000 (N_19000,N_11249,N_12048);
xnor U19001 (N_19001,N_14087,N_12941);
nand U19002 (N_19002,N_10440,N_14302);
xnor U19003 (N_19003,N_13837,N_11446);
nor U19004 (N_19004,N_11959,N_11387);
or U19005 (N_19005,N_13824,N_13734);
xor U19006 (N_19006,N_14274,N_10161);
or U19007 (N_19007,N_13625,N_13070);
xnor U19008 (N_19008,N_14224,N_13647);
or U19009 (N_19009,N_13314,N_14659);
xnor U19010 (N_19010,N_12431,N_11899);
or U19011 (N_19011,N_12830,N_11300);
and U19012 (N_19012,N_11191,N_13746);
xnor U19013 (N_19013,N_11164,N_12220);
nor U19014 (N_19014,N_10384,N_11987);
and U19015 (N_19015,N_11337,N_10957);
and U19016 (N_19016,N_14552,N_10845);
nor U19017 (N_19017,N_11136,N_14048);
xnor U19018 (N_19018,N_11038,N_14998);
and U19019 (N_19019,N_11083,N_13803);
or U19020 (N_19020,N_13562,N_10049);
nand U19021 (N_19021,N_10875,N_10712);
or U19022 (N_19022,N_14800,N_14079);
and U19023 (N_19023,N_12149,N_12725);
xnor U19024 (N_19024,N_14607,N_14253);
xnor U19025 (N_19025,N_13626,N_11679);
or U19026 (N_19026,N_13725,N_10224);
and U19027 (N_19027,N_14296,N_14563);
nand U19028 (N_19028,N_13423,N_12926);
nand U19029 (N_19029,N_12213,N_12635);
xnor U19030 (N_19030,N_10698,N_11145);
nand U19031 (N_19031,N_14661,N_11209);
and U19032 (N_19032,N_14991,N_13678);
xnor U19033 (N_19033,N_12094,N_10505);
nor U19034 (N_19034,N_11111,N_12040);
nand U19035 (N_19035,N_11947,N_13861);
xor U19036 (N_19036,N_12256,N_11147);
nor U19037 (N_19037,N_14844,N_12058);
xnor U19038 (N_19038,N_11755,N_13085);
nand U19039 (N_19039,N_10602,N_13306);
and U19040 (N_19040,N_13670,N_12077);
or U19041 (N_19041,N_13402,N_11794);
and U19042 (N_19042,N_12916,N_13275);
nor U19043 (N_19043,N_12567,N_12234);
or U19044 (N_19044,N_11032,N_12963);
or U19045 (N_19045,N_12656,N_11410);
and U19046 (N_19046,N_11617,N_14974);
nor U19047 (N_19047,N_13465,N_10704);
and U19048 (N_19048,N_13382,N_11068);
nand U19049 (N_19049,N_10460,N_10041);
nor U19050 (N_19050,N_10339,N_10445);
and U19051 (N_19051,N_14387,N_12600);
or U19052 (N_19052,N_14180,N_13051);
and U19053 (N_19053,N_13440,N_10711);
nand U19054 (N_19054,N_11709,N_11234);
nand U19055 (N_19055,N_13549,N_12269);
or U19056 (N_19056,N_10125,N_14035);
or U19057 (N_19057,N_13479,N_12262);
nand U19058 (N_19058,N_12209,N_13919);
nor U19059 (N_19059,N_13284,N_12171);
nand U19060 (N_19060,N_12963,N_14940);
nand U19061 (N_19061,N_13737,N_10001);
nand U19062 (N_19062,N_11907,N_14550);
nand U19063 (N_19063,N_11372,N_11882);
nand U19064 (N_19064,N_11548,N_11937);
nand U19065 (N_19065,N_11758,N_10010);
or U19066 (N_19066,N_14263,N_14390);
and U19067 (N_19067,N_11318,N_14331);
nor U19068 (N_19068,N_10461,N_14040);
nor U19069 (N_19069,N_10641,N_13183);
or U19070 (N_19070,N_10635,N_12029);
xor U19071 (N_19071,N_13573,N_14145);
nor U19072 (N_19072,N_12110,N_10059);
and U19073 (N_19073,N_12703,N_11067);
nand U19074 (N_19074,N_11724,N_13215);
nand U19075 (N_19075,N_12183,N_11522);
xnor U19076 (N_19076,N_13404,N_13792);
and U19077 (N_19077,N_14843,N_13415);
and U19078 (N_19078,N_14142,N_14970);
and U19079 (N_19079,N_13973,N_14943);
nor U19080 (N_19080,N_14632,N_10301);
nand U19081 (N_19081,N_13712,N_11796);
nor U19082 (N_19082,N_11790,N_12875);
xor U19083 (N_19083,N_13569,N_14784);
and U19084 (N_19084,N_12726,N_13532);
nor U19085 (N_19085,N_10985,N_14300);
nor U19086 (N_19086,N_10493,N_10602);
and U19087 (N_19087,N_14709,N_10768);
nand U19088 (N_19088,N_11831,N_10489);
and U19089 (N_19089,N_13466,N_14987);
and U19090 (N_19090,N_14796,N_10857);
or U19091 (N_19091,N_11456,N_12231);
and U19092 (N_19092,N_13309,N_13880);
and U19093 (N_19093,N_10080,N_13121);
or U19094 (N_19094,N_12071,N_12533);
nand U19095 (N_19095,N_11842,N_11148);
or U19096 (N_19096,N_14476,N_12577);
xnor U19097 (N_19097,N_14792,N_10511);
and U19098 (N_19098,N_13340,N_11070);
or U19099 (N_19099,N_14568,N_11870);
xor U19100 (N_19100,N_11706,N_10515);
xor U19101 (N_19101,N_14278,N_11973);
xor U19102 (N_19102,N_14336,N_13182);
nor U19103 (N_19103,N_11669,N_12528);
and U19104 (N_19104,N_12786,N_11611);
nor U19105 (N_19105,N_13327,N_13964);
or U19106 (N_19106,N_12539,N_12310);
and U19107 (N_19107,N_10093,N_12863);
or U19108 (N_19108,N_13277,N_13531);
nand U19109 (N_19109,N_10910,N_12314);
or U19110 (N_19110,N_14088,N_14809);
nor U19111 (N_19111,N_10583,N_14531);
nor U19112 (N_19112,N_10634,N_14335);
and U19113 (N_19113,N_10146,N_11333);
or U19114 (N_19114,N_11595,N_12818);
nand U19115 (N_19115,N_11024,N_12013);
xor U19116 (N_19116,N_10715,N_10087);
or U19117 (N_19117,N_14279,N_14874);
or U19118 (N_19118,N_11175,N_14868);
nor U19119 (N_19119,N_12323,N_13531);
and U19120 (N_19120,N_12334,N_11807);
nand U19121 (N_19121,N_11886,N_11026);
xor U19122 (N_19122,N_14751,N_14990);
nand U19123 (N_19123,N_12985,N_11580);
xor U19124 (N_19124,N_14583,N_14358);
and U19125 (N_19125,N_13822,N_13131);
or U19126 (N_19126,N_10424,N_10344);
or U19127 (N_19127,N_13007,N_14614);
nor U19128 (N_19128,N_13680,N_11791);
or U19129 (N_19129,N_11128,N_14553);
xnor U19130 (N_19130,N_11046,N_10203);
nor U19131 (N_19131,N_12418,N_14891);
xor U19132 (N_19132,N_13055,N_10304);
nor U19133 (N_19133,N_11579,N_13762);
xor U19134 (N_19134,N_14126,N_14295);
or U19135 (N_19135,N_11741,N_12123);
and U19136 (N_19136,N_14554,N_13602);
xnor U19137 (N_19137,N_14891,N_12685);
xor U19138 (N_19138,N_11190,N_13773);
nand U19139 (N_19139,N_10328,N_13099);
xnor U19140 (N_19140,N_11027,N_14487);
xnor U19141 (N_19141,N_10629,N_13475);
nand U19142 (N_19142,N_10998,N_14709);
nand U19143 (N_19143,N_14141,N_12584);
nor U19144 (N_19144,N_12016,N_13745);
and U19145 (N_19145,N_14607,N_11439);
nand U19146 (N_19146,N_14339,N_14075);
nand U19147 (N_19147,N_13599,N_12090);
xnor U19148 (N_19148,N_14212,N_14941);
or U19149 (N_19149,N_12483,N_11230);
or U19150 (N_19150,N_11023,N_13340);
or U19151 (N_19151,N_13233,N_10157);
or U19152 (N_19152,N_10369,N_10581);
or U19153 (N_19153,N_11525,N_13768);
or U19154 (N_19154,N_11664,N_14535);
nor U19155 (N_19155,N_13723,N_12583);
nor U19156 (N_19156,N_10470,N_14398);
and U19157 (N_19157,N_10480,N_14414);
nand U19158 (N_19158,N_12084,N_14829);
or U19159 (N_19159,N_11624,N_14762);
and U19160 (N_19160,N_13459,N_11471);
nand U19161 (N_19161,N_14420,N_12537);
nor U19162 (N_19162,N_13278,N_10397);
nor U19163 (N_19163,N_14856,N_11642);
and U19164 (N_19164,N_12146,N_12465);
nand U19165 (N_19165,N_14156,N_14296);
nor U19166 (N_19166,N_10163,N_10487);
nor U19167 (N_19167,N_11250,N_12239);
and U19168 (N_19168,N_11442,N_13184);
nand U19169 (N_19169,N_12879,N_12521);
or U19170 (N_19170,N_13572,N_10255);
nand U19171 (N_19171,N_10806,N_12264);
nor U19172 (N_19172,N_12833,N_12976);
or U19173 (N_19173,N_12297,N_12063);
or U19174 (N_19174,N_12746,N_12353);
nor U19175 (N_19175,N_12036,N_13498);
or U19176 (N_19176,N_11263,N_13926);
nor U19177 (N_19177,N_11331,N_14130);
xnor U19178 (N_19178,N_12711,N_13236);
xor U19179 (N_19179,N_10327,N_10599);
xnor U19180 (N_19180,N_11399,N_12071);
and U19181 (N_19181,N_13351,N_13985);
or U19182 (N_19182,N_10644,N_11221);
nand U19183 (N_19183,N_10405,N_11742);
nand U19184 (N_19184,N_14797,N_13666);
or U19185 (N_19185,N_10144,N_12700);
or U19186 (N_19186,N_12357,N_13831);
nor U19187 (N_19187,N_11698,N_10003);
and U19188 (N_19188,N_14100,N_13470);
or U19189 (N_19189,N_14988,N_12762);
nand U19190 (N_19190,N_14148,N_14521);
nand U19191 (N_19191,N_11093,N_14358);
or U19192 (N_19192,N_10329,N_10038);
xnor U19193 (N_19193,N_11279,N_11821);
and U19194 (N_19194,N_13844,N_10600);
or U19195 (N_19195,N_11576,N_11192);
nor U19196 (N_19196,N_10365,N_14321);
and U19197 (N_19197,N_11960,N_11921);
and U19198 (N_19198,N_14902,N_14621);
nand U19199 (N_19199,N_14907,N_13480);
and U19200 (N_19200,N_14426,N_10354);
nand U19201 (N_19201,N_11784,N_12965);
nor U19202 (N_19202,N_13939,N_13772);
or U19203 (N_19203,N_14071,N_14592);
nand U19204 (N_19204,N_14913,N_12023);
or U19205 (N_19205,N_14856,N_13382);
and U19206 (N_19206,N_13145,N_13946);
nand U19207 (N_19207,N_14099,N_13201);
nand U19208 (N_19208,N_13950,N_13670);
or U19209 (N_19209,N_13356,N_12703);
nor U19210 (N_19210,N_10812,N_11886);
or U19211 (N_19211,N_14021,N_12687);
or U19212 (N_19212,N_14599,N_12747);
or U19213 (N_19213,N_13521,N_13338);
and U19214 (N_19214,N_12724,N_11618);
nor U19215 (N_19215,N_11702,N_14914);
and U19216 (N_19216,N_12498,N_10198);
nor U19217 (N_19217,N_14009,N_12927);
xor U19218 (N_19218,N_10236,N_13684);
nor U19219 (N_19219,N_10219,N_12912);
nand U19220 (N_19220,N_11000,N_14458);
or U19221 (N_19221,N_12365,N_11255);
nand U19222 (N_19222,N_10623,N_14462);
nand U19223 (N_19223,N_14832,N_12131);
and U19224 (N_19224,N_13366,N_14886);
nor U19225 (N_19225,N_13339,N_10942);
xnor U19226 (N_19226,N_14390,N_14477);
and U19227 (N_19227,N_11677,N_11696);
nor U19228 (N_19228,N_12341,N_14102);
or U19229 (N_19229,N_10761,N_12696);
or U19230 (N_19230,N_11207,N_14551);
nor U19231 (N_19231,N_12209,N_11525);
and U19232 (N_19232,N_11677,N_14111);
nor U19233 (N_19233,N_11997,N_12022);
xnor U19234 (N_19234,N_10456,N_14656);
or U19235 (N_19235,N_12303,N_10034);
xor U19236 (N_19236,N_12541,N_10245);
nor U19237 (N_19237,N_13522,N_13266);
nand U19238 (N_19238,N_11042,N_13622);
nor U19239 (N_19239,N_12982,N_14938);
and U19240 (N_19240,N_10700,N_12420);
xnor U19241 (N_19241,N_10210,N_14300);
nand U19242 (N_19242,N_12215,N_10475);
xnor U19243 (N_19243,N_14190,N_14853);
nor U19244 (N_19244,N_13832,N_14039);
or U19245 (N_19245,N_11332,N_14564);
xor U19246 (N_19246,N_14719,N_12696);
xor U19247 (N_19247,N_10371,N_14650);
and U19248 (N_19248,N_10891,N_11326);
nor U19249 (N_19249,N_12181,N_13314);
xor U19250 (N_19250,N_10367,N_14978);
and U19251 (N_19251,N_13024,N_12719);
or U19252 (N_19252,N_12239,N_11766);
and U19253 (N_19253,N_10868,N_10841);
and U19254 (N_19254,N_14448,N_14338);
and U19255 (N_19255,N_14285,N_12367);
and U19256 (N_19256,N_10988,N_11445);
and U19257 (N_19257,N_14261,N_14880);
or U19258 (N_19258,N_10825,N_13349);
nor U19259 (N_19259,N_11462,N_10345);
or U19260 (N_19260,N_12259,N_10258);
and U19261 (N_19261,N_13457,N_11744);
and U19262 (N_19262,N_12959,N_14777);
xor U19263 (N_19263,N_11647,N_12208);
xnor U19264 (N_19264,N_13071,N_11363);
or U19265 (N_19265,N_12280,N_11845);
or U19266 (N_19266,N_14754,N_14048);
and U19267 (N_19267,N_13181,N_11589);
nor U19268 (N_19268,N_11688,N_12841);
and U19269 (N_19269,N_10796,N_10737);
and U19270 (N_19270,N_13295,N_13613);
nand U19271 (N_19271,N_14262,N_12991);
and U19272 (N_19272,N_12775,N_14259);
nand U19273 (N_19273,N_13255,N_13000);
and U19274 (N_19274,N_14090,N_11209);
nand U19275 (N_19275,N_11571,N_12651);
nand U19276 (N_19276,N_14405,N_12817);
or U19277 (N_19277,N_13789,N_11964);
or U19278 (N_19278,N_11239,N_14680);
or U19279 (N_19279,N_10748,N_14840);
nand U19280 (N_19280,N_14686,N_12376);
and U19281 (N_19281,N_13311,N_11317);
and U19282 (N_19282,N_13598,N_12365);
nor U19283 (N_19283,N_12632,N_12528);
or U19284 (N_19284,N_13524,N_13478);
nand U19285 (N_19285,N_14574,N_14348);
or U19286 (N_19286,N_14650,N_14505);
and U19287 (N_19287,N_11546,N_12814);
nor U19288 (N_19288,N_12718,N_10511);
and U19289 (N_19289,N_13641,N_10699);
nand U19290 (N_19290,N_10134,N_11297);
and U19291 (N_19291,N_11741,N_12448);
and U19292 (N_19292,N_11168,N_14560);
or U19293 (N_19293,N_14811,N_14661);
nand U19294 (N_19294,N_11144,N_13164);
xnor U19295 (N_19295,N_10850,N_12332);
or U19296 (N_19296,N_12364,N_13241);
xnor U19297 (N_19297,N_10818,N_14514);
and U19298 (N_19298,N_13182,N_11388);
nor U19299 (N_19299,N_13365,N_13034);
or U19300 (N_19300,N_10545,N_12551);
or U19301 (N_19301,N_10922,N_12099);
and U19302 (N_19302,N_10248,N_11363);
nor U19303 (N_19303,N_11408,N_10948);
nand U19304 (N_19304,N_11498,N_14658);
and U19305 (N_19305,N_11619,N_14187);
nand U19306 (N_19306,N_10408,N_11784);
xnor U19307 (N_19307,N_11117,N_10581);
and U19308 (N_19308,N_13671,N_11635);
nand U19309 (N_19309,N_14196,N_13182);
nand U19310 (N_19310,N_10402,N_12272);
nor U19311 (N_19311,N_12759,N_12226);
nor U19312 (N_19312,N_11098,N_12689);
or U19313 (N_19313,N_12267,N_14972);
or U19314 (N_19314,N_11607,N_10199);
nor U19315 (N_19315,N_11005,N_10055);
nand U19316 (N_19316,N_10970,N_14310);
nor U19317 (N_19317,N_10027,N_13635);
xor U19318 (N_19318,N_12969,N_10814);
and U19319 (N_19319,N_11200,N_12869);
nor U19320 (N_19320,N_11731,N_14518);
nor U19321 (N_19321,N_12759,N_10325);
or U19322 (N_19322,N_13557,N_10679);
xnor U19323 (N_19323,N_12655,N_13277);
and U19324 (N_19324,N_14359,N_12086);
or U19325 (N_19325,N_12364,N_13546);
nand U19326 (N_19326,N_12006,N_14792);
nor U19327 (N_19327,N_11794,N_10356);
or U19328 (N_19328,N_14250,N_11207);
and U19329 (N_19329,N_11636,N_12470);
nand U19330 (N_19330,N_12014,N_13552);
and U19331 (N_19331,N_10185,N_10697);
or U19332 (N_19332,N_14248,N_14440);
and U19333 (N_19333,N_13466,N_11953);
nand U19334 (N_19334,N_13514,N_10406);
xnor U19335 (N_19335,N_10251,N_11331);
nor U19336 (N_19336,N_12664,N_11477);
or U19337 (N_19337,N_12038,N_13679);
or U19338 (N_19338,N_11932,N_13649);
nor U19339 (N_19339,N_13085,N_11851);
xor U19340 (N_19340,N_14046,N_10227);
or U19341 (N_19341,N_10739,N_14538);
nand U19342 (N_19342,N_12575,N_11011);
xor U19343 (N_19343,N_10435,N_11297);
nand U19344 (N_19344,N_10856,N_12359);
nand U19345 (N_19345,N_10720,N_14178);
or U19346 (N_19346,N_12101,N_14840);
nor U19347 (N_19347,N_13990,N_11202);
nor U19348 (N_19348,N_10452,N_14835);
nor U19349 (N_19349,N_11042,N_11339);
nor U19350 (N_19350,N_12808,N_11075);
nor U19351 (N_19351,N_12626,N_10478);
nor U19352 (N_19352,N_13185,N_11734);
nor U19353 (N_19353,N_12003,N_13732);
and U19354 (N_19354,N_10584,N_10052);
nor U19355 (N_19355,N_12311,N_13202);
nor U19356 (N_19356,N_14847,N_11764);
xnor U19357 (N_19357,N_14489,N_14043);
xor U19358 (N_19358,N_14388,N_14082);
nand U19359 (N_19359,N_12202,N_11982);
nor U19360 (N_19360,N_10387,N_13788);
nand U19361 (N_19361,N_14057,N_13372);
nand U19362 (N_19362,N_11186,N_11393);
or U19363 (N_19363,N_14002,N_14768);
nand U19364 (N_19364,N_10759,N_11812);
nand U19365 (N_19365,N_12186,N_14426);
or U19366 (N_19366,N_10134,N_10215);
nand U19367 (N_19367,N_10096,N_12837);
nand U19368 (N_19368,N_13206,N_10447);
nor U19369 (N_19369,N_13153,N_10135);
or U19370 (N_19370,N_11930,N_13182);
and U19371 (N_19371,N_11463,N_14982);
nor U19372 (N_19372,N_12311,N_13616);
nand U19373 (N_19373,N_11904,N_11110);
xor U19374 (N_19374,N_10444,N_12021);
xnor U19375 (N_19375,N_10597,N_12266);
or U19376 (N_19376,N_11207,N_14221);
or U19377 (N_19377,N_13616,N_10146);
nor U19378 (N_19378,N_11667,N_12024);
xnor U19379 (N_19379,N_10714,N_13238);
and U19380 (N_19380,N_10465,N_13671);
and U19381 (N_19381,N_14208,N_13491);
nor U19382 (N_19382,N_10938,N_14172);
nor U19383 (N_19383,N_14522,N_10876);
and U19384 (N_19384,N_10449,N_12295);
and U19385 (N_19385,N_12873,N_11370);
nand U19386 (N_19386,N_11349,N_12634);
nor U19387 (N_19387,N_14633,N_12359);
nor U19388 (N_19388,N_13393,N_14525);
xor U19389 (N_19389,N_12698,N_11829);
and U19390 (N_19390,N_12477,N_14277);
or U19391 (N_19391,N_13442,N_12432);
nor U19392 (N_19392,N_11739,N_12725);
nor U19393 (N_19393,N_12503,N_13092);
nor U19394 (N_19394,N_10678,N_13365);
nor U19395 (N_19395,N_14056,N_10220);
and U19396 (N_19396,N_12758,N_13266);
or U19397 (N_19397,N_10265,N_11418);
and U19398 (N_19398,N_14489,N_13318);
nor U19399 (N_19399,N_13058,N_14230);
xnor U19400 (N_19400,N_13536,N_14611);
and U19401 (N_19401,N_14097,N_13994);
xor U19402 (N_19402,N_12176,N_12131);
and U19403 (N_19403,N_10518,N_12094);
nand U19404 (N_19404,N_12410,N_11305);
xnor U19405 (N_19405,N_10319,N_11005);
or U19406 (N_19406,N_12779,N_10903);
xnor U19407 (N_19407,N_12812,N_10264);
and U19408 (N_19408,N_14937,N_11223);
xor U19409 (N_19409,N_12718,N_10611);
nand U19410 (N_19410,N_14490,N_14141);
xnor U19411 (N_19411,N_12286,N_14541);
or U19412 (N_19412,N_14765,N_11784);
nor U19413 (N_19413,N_14522,N_12728);
or U19414 (N_19414,N_10556,N_11476);
and U19415 (N_19415,N_11994,N_12187);
xor U19416 (N_19416,N_11772,N_12581);
nor U19417 (N_19417,N_12163,N_12770);
xnor U19418 (N_19418,N_14101,N_10555);
or U19419 (N_19419,N_13651,N_10089);
nor U19420 (N_19420,N_14900,N_12311);
and U19421 (N_19421,N_13109,N_14247);
nand U19422 (N_19422,N_10145,N_10996);
xnor U19423 (N_19423,N_10522,N_12426);
xnor U19424 (N_19424,N_12771,N_11612);
or U19425 (N_19425,N_12412,N_14538);
nand U19426 (N_19426,N_12074,N_10678);
or U19427 (N_19427,N_14472,N_10474);
and U19428 (N_19428,N_13902,N_11568);
or U19429 (N_19429,N_13996,N_12330);
and U19430 (N_19430,N_13870,N_11785);
or U19431 (N_19431,N_10772,N_12840);
nand U19432 (N_19432,N_11260,N_10513);
nor U19433 (N_19433,N_11189,N_13234);
or U19434 (N_19434,N_11866,N_13713);
or U19435 (N_19435,N_12157,N_14888);
nor U19436 (N_19436,N_14574,N_14295);
nor U19437 (N_19437,N_12975,N_13109);
nand U19438 (N_19438,N_13549,N_10087);
or U19439 (N_19439,N_10614,N_11489);
xor U19440 (N_19440,N_10922,N_13385);
and U19441 (N_19441,N_11309,N_14564);
nor U19442 (N_19442,N_14198,N_10835);
nor U19443 (N_19443,N_11029,N_13443);
xnor U19444 (N_19444,N_11825,N_12773);
or U19445 (N_19445,N_13972,N_14720);
or U19446 (N_19446,N_14218,N_14019);
nor U19447 (N_19447,N_11209,N_13771);
or U19448 (N_19448,N_10066,N_13404);
or U19449 (N_19449,N_13001,N_11577);
and U19450 (N_19450,N_13892,N_11519);
nand U19451 (N_19451,N_14816,N_14429);
and U19452 (N_19452,N_12916,N_11034);
xnor U19453 (N_19453,N_13567,N_12371);
xor U19454 (N_19454,N_11767,N_14885);
and U19455 (N_19455,N_13988,N_12950);
nor U19456 (N_19456,N_14496,N_11672);
xor U19457 (N_19457,N_12298,N_13535);
xor U19458 (N_19458,N_10417,N_10916);
or U19459 (N_19459,N_13045,N_12266);
and U19460 (N_19460,N_12934,N_12194);
xor U19461 (N_19461,N_13141,N_10606);
and U19462 (N_19462,N_12636,N_13663);
xnor U19463 (N_19463,N_12214,N_13565);
and U19464 (N_19464,N_10298,N_10077);
and U19465 (N_19465,N_11022,N_12686);
nand U19466 (N_19466,N_11091,N_12097);
and U19467 (N_19467,N_12866,N_11016);
xor U19468 (N_19468,N_12256,N_14174);
nand U19469 (N_19469,N_14906,N_11406);
and U19470 (N_19470,N_13337,N_13894);
and U19471 (N_19471,N_12758,N_10034);
nor U19472 (N_19472,N_10027,N_10473);
xnor U19473 (N_19473,N_10402,N_13399);
nor U19474 (N_19474,N_11063,N_14328);
or U19475 (N_19475,N_14276,N_12082);
xor U19476 (N_19476,N_11733,N_14516);
nor U19477 (N_19477,N_13252,N_10469);
or U19478 (N_19478,N_10336,N_12442);
nand U19479 (N_19479,N_11664,N_13756);
xnor U19480 (N_19480,N_14763,N_11920);
xor U19481 (N_19481,N_12975,N_11231);
and U19482 (N_19482,N_11572,N_11074);
nand U19483 (N_19483,N_11060,N_13817);
nand U19484 (N_19484,N_13951,N_10743);
nor U19485 (N_19485,N_11371,N_12366);
and U19486 (N_19486,N_11282,N_11181);
and U19487 (N_19487,N_12570,N_11959);
xor U19488 (N_19488,N_11885,N_13856);
nor U19489 (N_19489,N_10657,N_14756);
nor U19490 (N_19490,N_13184,N_11015);
or U19491 (N_19491,N_12178,N_12528);
nor U19492 (N_19492,N_13158,N_13319);
and U19493 (N_19493,N_13580,N_12305);
and U19494 (N_19494,N_13524,N_12005);
nor U19495 (N_19495,N_12101,N_14006);
nand U19496 (N_19496,N_10402,N_12951);
nor U19497 (N_19497,N_14159,N_10618);
or U19498 (N_19498,N_12517,N_10902);
nor U19499 (N_19499,N_14780,N_10387);
or U19500 (N_19500,N_12795,N_14823);
nand U19501 (N_19501,N_13245,N_11931);
xnor U19502 (N_19502,N_11245,N_14134);
and U19503 (N_19503,N_10639,N_14642);
xnor U19504 (N_19504,N_13693,N_11412);
nand U19505 (N_19505,N_12879,N_11928);
nand U19506 (N_19506,N_14662,N_14401);
xnor U19507 (N_19507,N_12371,N_11867);
xnor U19508 (N_19508,N_11600,N_14546);
or U19509 (N_19509,N_13667,N_11060);
nor U19510 (N_19510,N_11149,N_10141);
nand U19511 (N_19511,N_11702,N_14407);
and U19512 (N_19512,N_11295,N_14781);
nor U19513 (N_19513,N_13567,N_10669);
or U19514 (N_19514,N_12950,N_10735);
and U19515 (N_19515,N_12721,N_12987);
and U19516 (N_19516,N_13003,N_13385);
nand U19517 (N_19517,N_13662,N_13764);
and U19518 (N_19518,N_11922,N_14953);
or U19519 (N_19519,N_10185,N_11565);
or U19520 (N_19520,N_13252,N_11889);
nor U19521 (N_19521,N_12365,N_12726);
and U19522 (N_19522,N_12468,N_12789);
or U19523 (N_19523,N_13983,N_10245);
and U19524 (N_19524,N_14153,N_10104);
nor U19525 (N_19525,N_10420,N_11999);
nand U19526 (N_19526,N_12806,N_10799);
nor U19527 (N_19527,N_12885,N_14956);
nor U19528 (N_19528,N_14571,N_13272);
xor U19529 (N_19529,N_13897,N_13668);
nand U19530 (N_19530,N_14755,N_11593);
xnor U19531 (N_19531,N_13746,N_10089);
nand U19532 (N_19532,N_11928,N_10515);
xnor U19533 (N_19533,N_14052,N_13599);
nor U19534 (N_19534,N_13637,N_10006);
and U19535 (N_19535,N_11248,N_14899);
or U19536 (N_19536,N_13125,N_14898);
or U19537 (N_19537,N_14903,N_11999);
or U19538 (N_19538,N_13769,N_11205);
nand U19539 (N_19539,N_10592,N_13384);
or U19540 (N_19540,N_13259,N_14642);
nand U19541 (N_19541,N_10756,N_12523);
xor U19542 (N_19542,N_13829,N_11773);
nand U19543 (N_19543,N_12124,N_12244);
and U19544 (N_19544,N_10739,N_10518);
or U19545 (N_19545,N_14584,N_10425);
and U19546 (N_19546,N_10315,N_12403);
or U19547 (N_19547,N_12312,N_12203);
or U19548 (N_19548,N_13638,N_14263);
nand U19549 (N_19549,N_10036,N_10620);
nand U19550 (N_19550,N_13198,N_10863);
and U19551 (N_19551,N_11926,N_13466);
xnor U19552 (N_19552,N_11131,N_12896);
xnor U19553 (N_19553,N_11155,N_11943);
or U19554 (N_19554,N_10405,N_10972);
and U19555 (N_19555,N_11817,N_10973);
nand U19556 (N_19556,N_13805,N_12082);
or U19557 (N_19557,N_12298,N_10615);
nand U19558 (N_19558,N_10550,N_12599);
and U19559 (N_19559,N_11480,N_11825);
and U19560 (N_19560,N_10220,N_12539);
or U19561 (N_19561,N_11417,N_10209);
or U19562 (N_19562,N_12905,N_13234);
nand U19563 (N_19563,N_12202,N_14608);
or U19564 (N_19564,N_14150,N_10462);
or U19565 (N_19565,N_12494,N_11390);
or U19566 (N_19566,N_14586,N_12162);
and U19567 (N_19567,N_11552,N_12611);
or U19568 (N_19568,N_13379,N_13394);
nand U19569 (N_19569,N_13866,N_13194);
xnor U19570 (N_19570,N_14712,N_12342);
nor U19571 (N_19571,N_10279,N_11277);
and U19572 (N_19572,N_12934,N_12072);
nor U19573 (N_19573,N_13562,N_11095);
nor U19574 (N_19574,N_11351,N_13547);
nor U19575 (N_19575,N_11682,N_14828);
and U19576 (N_19576,N_13806,N_11662);
or U19577 (N_19577,N_11632,N_11712);
and U19578 (N_19578,N_12821,N_12995);
and U19579 (N_19579,N_14101,N_13597);
and U19580 (N_19580,N_14383,N_14246);
nor U19581 (N_19581,N_11829,N_12097);
and U19582 (N_19582,N_11907,N_13680);
nor U19583 (N_19583,N_14459,N_10107);
and U19584 (N_19584,N_11590,N_11778);
xnor U19585 (N_19585,N_14487,N_10895);
nor U19586 (N_19586,N_12268,N_12142);
nand U19587 (N_19587,N_10231,N_13912);
nor U19588 (N_19588,N_14159,N_11516);
or U19589 (N_19589,N_12116,N_12511);
nor U19590 (N_19590,N_11525,N_13696);
or U19591 (N_19591,N_13794,N_14487);
nor U19592 (N_19592,N_12469,N_13045);
xnor U19593 (N_19593,N_13873,N_11856);
and U19594 (N_19594,N_14095,N_11246);
nand U19595 (N_19595,N_11343,N_11920);
nor U19596 (N_19596,N_13756,N_14315);
or U19597 (N_19597,N_10089,N_14252);
nor U19598 (N_19598,N_14776,N_13337);
and U19599 (N_19599,N_14069,N_12992);
nor U19600 (N_19600,N_14429,N_10553);
nand U19601 (N_19601,N_14852,N_13656);
nor U19602 (N_19602,N_13065,N_13077);
xor U19603 (N_19603,N_10157,N_14296);
and U19604 (N_19604,N_12524,N_11692);
and U19605 (N_19605,N_13474,N_14399);
xor U19606 (N_19606,N_13367,N_14585);
nor U19607 (N_19607,N_13890,N_12290);
and U19608 (N_19608,N_10919,N_14486);
and U19609 (N_19609,N_12050,N_13523);
or U19610 (N_19610,N_12489,N_13958);
or U19611 (N_19611,N_13364,N_14739);
and U19612 (N_19612,N_13247,N_13456);
or U19613 (N_19613,N_11355,N_13578);
and U19614 (N_19614,N_11409,N_13760);
and U19615 (N_19615,N_12429,N_10035);
and U19616 (N_19616,N_12215,N_10009);
and U19617 (N_19617,N_14603,N_14101);
and U19618 (N_19618,N_10196,N_11367);
and U19619 (N_19619,N_11765,N_12022);
nand U19620 (N_19620,N_11428,N_13967);
nor U19621 (N_19621,N_12813,N_14144);
xor U19622 (N_19622,N_11505,N_10406);
or U19623 (N_19623,N_10794,N_14742);
nor U19624 (N_19624,N_14130,N_14277);
or U19625 (N_19625,N_10739,N_12993);
nor U19626 (N_19626,N_12670,N_12027);
xnor U19627 (N_19627,N_13879,N_14877);
or U19628 (N_19628,N_10007,N_12663);
nor U19629 (N_19629,N_12163,N_12703);
or U19630 (N_19630,N_11661,N_14156);
nor U19631 (N_19631,N_11473,N_12338);
or U19632 (N_19632,N_13315,N_10485);
or U19633 (N_19633,N_14692,N_10685);
nand U19634 (N_19634,N_13469,N_14162);
or U19635 (N_19635,N_11288,N_13456);
nand U19636 (N_19636,N_11122,N_10751);
and U19637 (N_19637,N_10379,N_10461);
nand U19638 (N_19638,N_10587,N_14603);
or U19639 (N_19639,N_13529,N_12135);
xor U19640 (N_19640,N_14665,N_12224);
and U19641 (N_19641,N_11200,N_10810);
nor U19642 (N_19642,N_14979,N_11554);
or U19643 (N_19643,N_10747,N_10418);
nand U19644 (N_19644,N_12329,N_12432);
and U19645 (N_19645,N_10083,N_10689);
xnor U19646 (N_19646,N_14925,N_10850);
xnor U19647 (N_19647,N_12594,N_12036);
or U19648 (N_19648,N_11293,N_12825);
nor U19649 (N_19649,N_13365,N_13803);
nor U19650 (N_19650,N_13638,N_11166);
nor U19651 (N_19651,N_14426,N_11469);
or U19652 (N_19652,N_13747,N_12599);
nand U19653 (N_19653,N_11556,N_12113);
nor U19654 (N_19654,N_14115,N_14622);
xor U19655 (N_19655,N_10271,N_13966);
xor U19656 (N_19656,N_10771,N_14984);
xor U19657 (N_19657,N_14113,N_10580);
nand U19658 (N_19658,N_11446,N_12434);
and U19659 (N_19659,N_10766,N_12709);
nor U19660 (N_19660,N_12657,N_14587);
or U19661 (N_19661,N_11139,N_11125);
nor U19662 (N_19662,N_10792,N_14958);
xnor U19663 (N_19663,N_14922,N_12656);
nor U19664 (N_19664,N_11990,N_13535);
nor U19665 (N_19665,N_13569,N_14158);
or U19666 (N_19666,N_13569,N_12362);
and U19667 (N_19667,N_10691,N_10104);
nor U19668 (N_19668,N_13988,N_10795);
and U19669 (N_19669,N_12080,N_13338);
nor U19670 (N_19670,N_14388,N_10960);
nor U19671 (N_19671,N_13066,N_10370);
or U19672 (N_19672,N_10655,N_12534);
or U19673 (N_19673,N_14314,N_10221);
nand U19674 (N_19674,N_11355,N_10989);
xnor U19675 (N_19675,N_13224,N_13032);
or U19676 (N_19676,N_13822,N_11881);
nor U19677 (N_19677,N_11738,N_13462);
nor U19678 (N_19678,N_11695,N_13651);
or U19679 (N_19679,N_11675,N_11235);
xnor U19680 (N_19680,N_12603,N_12169);
xor U19681 (N_19681,N_12655,N_14458);
and U19682 (N_19682,N_10845,N_10663);
nand U19683 (N_19683,N_14993,N_10547);
xor U19684 (N_19684,N_13131,N_14503);
or U19685 (N_19685,N_10414,N_10712);
nand U19686 (N_19686,N_13648,N_14223);
nand U19687 (N_19687,N_13520,N_10173);
xnor U19688 (N_19688,N_12427,N_13962);
xor U19689 (N_19689,N_13446,N_14242);
xnor U19690 (N_19690,N_10510,N_13361);
nor U19691 (N_19691,N_13093,N_13561);
nor U19692 (N_19692,N_12117,N_12990);
nand U19693 (N_19693,N_11315,N_11481);
or U19694 (N_19694,N_13064,N_12813);
xnor U19695 (N_19695,N_12913,N_12801);
and U19696 (N_19696,N_11470,N_11433);
nor U19697 (N_19697,N_10176,N_11420);
xnor U19698 (N_19698,N_10284,N_12708);
xor U19699 (N_19699,N_11172,N_10825);
nand U19700 (N_19700,N_10396,N_12043);
and U19701 (N_19701,N_11359,N_14941);
or U19702 (N_19702,N_13824,N_10567);
or U19703 (N_19703,N_13504,N_13231);
nand U19704 (N_19704,N_12351,N_14128);
and U19705 (N_19705,N_13450,N_10433);
nand U19706 (N_19706,N_10763,N_11898);
or U19707 (N_19707,N_11548,N_10966);
nand U19708 (N_19708,N_10781,N_13717);
xnor U19709 (N_19709,N_12218,N_13646);
xor U19710 (N_19710,N_12048,N_11622);
nand U19711 (N_19711,N_10219,N_11349);
nor U19712 (N_19712,N_11427,N_14146);
nand U19713 (N_19713,N_10908,N_11642);
or U19714 (N_19714,N_10958,N_10332);
and U19715 (N_19715,N_11435,N_13354);
xnor U19716 (N_19716,N_12462,N_11189);
and U19717 (N_19717,N_13023,N_14131);
nor U19718 (N_19718,N_10581,N_13014);
nor U19719 (N_19719,N_10671,N_10490);
nor U19720 (N_19720,N_13625,N_13298);
and U19721 (N_19721,N_13188,N_13633);
xnor U19722 (N_19722,N_14210,N_13071);
xor U19723 (N_19723,N_14901,N_13492);
or U19724 (N_19724,N_14153,N_12990);
and U19725 (N_19725,N_13287,N_12074);
nor U19726 (N_19726,N_12548,N_11778);
and U19727 (N_19727,N_12811,N_13398);
and U19728 (N_19728,N_11530,N_11423);
nor U19729 (N_19729,N_11319,N_13106);
or U19730 (N_19730,N_12056,N_14486);
nand U19731 (N_19731,N_12708,N_11324);
and U19732 (N_19732,N_13035,N_13360);
or U19733 (N_19733,N_11977,N_11236);
and U19734 (N_19734,N_12566,N_14875);
or U19735 (N_19735,N_12323,N_12035);
xnor U19736 (N_19736,N_13694,N_10754);
or U19737 (N_19737,N_11197,N_12229);
xor U19738 (N_19738,N_14533,N_13858);
nand U19739 (N_19739,N_14511,N_10859);
nor U19740 (N_19740,N_11900,N_11723);
xnor U19741 (N_19741,N_12875,N_12372);
and U19742 (N_19742,N_10971,N_11102);
or U19743 (N_19743,N_12836,N_12417);
xnor U19744 (N_19744,N_14083,N_14356);
or U19745 (N_19745,N_14465,N_11808);
and U19746 (N_19746,N_13168,N_10336);
nand U19747 (N_19747,N_10815,N_11569);
nor U19748 (N_19748,N_12838,N_12710);
xor U19749 (N_19749,N_10052,N_12259);
and U19750 (N_19750,N_12670,N_13290);
or U19751 (N_19751,N_11850,N_13689);
nor U19752 (N_19752,N_12717,N_10310);
or U19753 (N_19753,N_13074,N_10209);
and U19754 (N_19754,N_14145,N_11957);
nand U19755 (N_19755,N_13902,N_10313);
nor U19756 (N_19756,N_13402,N_10450);
or U19757 (N_19757,N_13408,N_11589);
nor U19758 (N_19758,N_10348,N_10941);
xor U19759 (N_19759,N_12952,N_12357);
and U19760 (N_19760,N_14216,N_12449);
or U19761 (N_19761,N_14138,N_11531);
nand U19762 (N_19762,N_14315,N_14058);
xnor U19763 (N_19763,N_14277,N_14176);
and U19764 (N_19764,N_14287,N_14219);
nor U19765 (N_19765,N_11278,N_11821);
nand U19766 (N_19766,N_12269,N_11134);
xnor U19767 (N_19767,N_14648,N_11178);
xor U19768 (N_19768,N_11467,N_12408);
and U19769 (N_19769,N_10922,N_11457);
and U19770 (N_19770,N_10261,N_10676);
or U19771 (N_19771,N_10080,N_11888);
and U19772 (N_19772,N_12220,N_14572);
and U19773 (N_19773,N_13122,N_10048);
nor U19774 (N_19774,N_10718,N_13343);
nor U19775 (N_19775,N_10594,N_12640);
nor U19776 (N_19776,N_10510,N_11931);
xor U19777 (N_19777,N_11022,N_10569);
and U19778 (N_19778,N_10198,N_11788);
nor U19779 (N_19779,N_13731,N_12326);
nand U19780 (N_19780,N_12016,N_14619);
and U19781 (N_19781,N_13926,N_10510);
nor U19782 (N_19782,N_14468,N_14457);
or U19783 (N_19783,N_10449,N_13281);
and U19784 (N_19784,N_12576,N_14216);
xor U19785 (N_19785,N_12714,N_11452);
nor U19786 (N_19786,N_12384,N_10035);
or U19787 (N_19787,N_14833,N_13935);
or U19788 (N_19788,N_13704,N_11830);
or U19789 (N_19789,N_10665,N_13127);
xor U19790 (N_19790,N_11554,N_12659);
nand U19791 (N_19791,N_11503,N_11855);
nor U19792 (N_19792,N_11314,N_12271);
nor U19793 (N_19793,N_14089,N_12804);
nor U19794 (N_19794,N_10197,N_10902);
and U19795 (N_19795,N_13343,N_10933);
nor U19796 (N_19796,N_10020,N_12764);
nor U19797 (N_19797,N_10093,N_10453);
and U19798 (N_19798,N_13569,N_12387);
nand U19799 (N_19799,N_14156,N_13695);
nor U19800 (N_19800,N_10405,N_11171);
and U19801 (N_19801,N_11097,N_12811);
nor U19802 (N_19802,N_12067,N_13400);
or U19803 (N_19803,N_10809,N_12179);
nor U19804 (N_19804,N_13641,N_12816);
or U19805 (N_19805,N_10994,N_13368);
nand U19806 (N_19806,N_12421,N_13353);
nor U19807 (N_19807,N_13516,N_12892);
nor U19808 (N_19808,N_13161,N_13220);
nor U19809 (N_19809,N_10541,N_12083);
nand U19810 (N_19810,N_11444,N_12423);
or U19811 (N_19811,N_11144,N_10224);
nand U19812 (N_19812,N_14734,N_14721);
nand U19813 (N_19813,N_12186,N_14711);
or U19814 (N_19814,N_14738,N_14644);
nor U19815 (N_19815,N_14581,N_12268);
nor U19816 (N_19816,N_14875,N_12113);
or U19817 (N_19817,N_13551,N_12750);
and U19818 (N_19818,N_12119,N_10830);
nor U19819 (N_19819,N_13549,N_11443);
and U19820 (N_19820,N_12665,N_14685);
or U19821 (N_19821,N_12374,N_12787);
nand U19822 (N_19822,N_14605,N_12098);
nor U19823 (N_19823,N_11664,N_10207);
nand U19824 (N_19824,N_11289,N_13411);
or U19825 (N_19825,N_10114,N_11074);
xor U19826 (N_19826,N_11524,N_14785);
xnor U19827 (N_19827,N_12405,N_13473);
or U19828 (N_19828,N_12036,N_13957);
nor U19829 (N_19829,N_14444,N_10977);
xnor U19830 (N_19830,N_14316,N_11764);
or U19831 (N_19831,N_13503,N_12554);
xnor U19832 (N_19832,N_11579,N_11378);
or U19833 (N_19833,N_13125,N_14508);
nor U19834 (N_19834,N_12257,N_11619);
nor U19835 (N_19835,N_14412,N_10065);
and U19836 (N_19836,N_12829,N_14132);
and U19837 (N_19837,N_12132,N_14281);
and U19838 (N_19838,N_11785,N_10614);
nor U19839 (N_19839,N_12201,N_12029);
and U19840 (N_19840,N_11028,N_11362);
or U19841 (N_19841,N_13228,N_11177);
xnor U19842 (N_19842,N_10552,N_14259);
nor U19843 (N_19843,N_13849,N_12750);
or U19844 (N_19844,N_10102,N_13363);
and U19845 (N_19845,N_13304,N_11253);
xor U19846 (N_19846,N_12501,N_14999);
or U19847 (N_19847,N_14972,N_13940);
xor U19848 (N_19848,N_11748,N_13869);
nand U19849 (N_19849,N_10830,N_10626);
nand U19850 (N_19850,N_10852,N_12917);
nor U19851 (N_19851,N_11411,N_14086);
nor U19852 (N_19852,N_11517,N_12692);
nor U19853 (N_19853,N_13307,N_13126);
and U19854 (N_19854,N_14855,N_10782);
and U19855 (N_19855,N_14470,N_10133);
nor U19856 (N_19856,N_12193,N_14724);
nand U19857 (N_19857,N_11362,N_11602);
or U19858 (N_19858,N_11992,N_14280);
or U19859 (N_19859,N_11273,N_12496);
nor U19860 (N_19860,N_13546,N_10461);
and U19861 (N_19861,N_11479,N_14494);
and U19862 (N_19862,N_14039,N_14603);
or U19863 (N_19863,N_10064,N_10833);
xnor U19864 (N_19864,N_14773,N_10898);
and U19865 (N_19865,N_11095,N_10520);
xnor U19866 (N_19866,N_13322,N_14703);
and U19867 (N_19867,N_11305,N_11747);
nor U19868 (N_19868,N_11888,N_14503);
nor U19869 (N_19869,N_14225,N_14970);
or U19870 (N_19870,N_13986,N_13583);
nand U19871 (N_19871,N_11103,N_10053);
xor U19872 (N_19872,N_11096,N_11171);
xnor U19873 (N_19873,N_12659,N_13550);
nor U19874 (N_19874,N_11944,N_14421);
xor U19875 (N_19875,N_11869,N_14972);
or U19876 (N_19876,N_12347,N_10559);
or U19877 (N_19877,N_13401,N_13720);
xor U19878 (N_19878,N_14990,N_11460);
or U19879 (N_19879,N_12951,N_10101);
nor U19880 (N_19880,N_10697,N_11563);
or U19881 (N_19881,N_14685,N_11760);
or U19882 (N_19882,N_10443,N_14155);
xnor U19883 (N_19883,N_12410,N_11872);
nand U19884 (N_19884,N_12262,N_10039);
nand U19885 (N_19885,N_11968,N_13603);
xnor U19886 (N_19886,N_10004,N_14177);
xor U19887 (N_19887,N_13875,N_12227);
and U19888 (N_19888,N_11576,N_10805);
nor U19889 (N_19889,N_12778,N_10325);
nand U19890 (N_19890,N_11987,N_12451);
nor U19891 (N_19891,N_14832,N_11352);
or U19892 (N_19892,N_11570,N_10608);
xnor U19893 (N_19893,N_14540,N_14353);
or U19894 (N_19894,N_12537,N_11375);
nor U19895 (N_19895,N_14639,N_14414);
or U19896 (N_19896,N_10079,N_13758);
nand U19897 (N_19897,N_11855,N_12260);
nand U19898 (N_19898,N_14193,N_11675);
xnor U19899 (N_19899,N_13259,N_12152);
and U19900 (N_19900,N_11867,N_14409);
and U19901 (N_19901,N_14911,N_10706);
and U19902 (N_19902,N_11557,N_14563);
xor U19903 (N_19903,N_10472,N_12412);
nand U19904 (N_19904,N_14255,N_11468);
nor U19905 (N_19905,N_13310,N_13320);
and U19906 (N_19906,N_12100,N_13366);
or U19907 (N_19907,N_13815,N_13371);
or U19908 (N_19908,N_11832,N_11655);
xnor U19909 (N_19909,N_14843,N_14205);
or U19910 (N_19910,N_12458,N_14184);
nand U19911 (N_19911,N_11051,N_13387);
or U19912 (N_19912,N_10585,N_14130);
and U19913 (N_19913,N_11925,N_13021);
and U19914 (N_19914,N_11333,N_10919);
xnor U19915 (N_19915,N_14212,N_11092);
nand U19916 (N_19916,N_11427,N_10055);
and U19917 (N_19917,N_11519,N_13266);
or U19918 (N_19918,N_10166,N_11709);
nor U19919 (N_19919,N_11470,N_10794);
nand U19920 (N_19920,N_11672,N_11191);
and U19921 (N_19921,N_12787,N_11741);
nand U19922 (N_19922,N_13050,N_13204);
xnor U19923 (N_19923,N_14089,N_11678);
xor U19924 (N_19924,N_12521,N_12970);
xnor U19925 (N_19925,N_13791,N_11768);
nand U19926 (N_19926,N_12738,N_11509);
or U19927 (N_19927,N_14954,N_14343);
and U19928 (N_19928,N_13372,N_11330);
and U19929 (N_19929,N_11440,N_10828);
or U19930 (N_19930,N_10863,N_10323);
nor U19931 (N_19931,N_14777,N_10821);
and U19932 (N_19932,N_13448,N_14026);
nor U19933 (N_19933,N_14411,N_11912);
nor U19934 (N_19934,N_13488,N_11953);
or U19935 (N_19935,N_11816,N_14695);
nor U19936 (N_19936,N_11012,N_10364);
or U19937 (N_19937,N_14282,N_10010);
and U19938 (N_19938,N_13863,N_10233);
or U19939 (N_19939,N_14765,N_11781);
nor U19940 (N_19940,N_12527,N_10792);
nand U19941 (N_19941,N_14763,N_14938);
or U19942 (N_19942,N_14495,N_10125);
or U19943 (N_19943,N_13867,N_14083);
or U19944 (N_19944,N_13654,N_13052);
nand U19945 (N_19945,N_11327,N_13714);
or U19946 (N_19946,N_10092,N_11125);
and U19947 (N_19947,N_14592,N_10558);
nor U19948 (N_19948,N_13268,N_11996);
nor U19949 (N_19949,N_11221,N_10081);
nor U19950 (N_19950,N_12237,N_14304);
nor U19951 (N_19951,N_10099,N_12911);
and U19952 (N_19952,N_11423,N_10310);
xnor U19953 (N_19953,N_12690,N_10813);
and U19954 (N_19954,N_11154,N_12897);
nand U19955 (N_19955,N_11398,N_12929);
and U19956 (N_19956,N_10899,N_12874);
nor U19957 (N_19957,N_12351,N_13988);
nand U19958 (N_19958,N_11211,N_10423);
or U19959 (N_19959,N_10390,N_12800);
nand U19960 (N_19960,N_11835,N_12409);
or U19961 (N_19961,N_11086,N_11561);
nand U19962 (N_19962,N_12805,N_12477);
nor U19963 (N_19963,N_14205,N_12618);
xnor U19964 (N_19964,N_10386,N_10466);
or U19965 (N_19965,N_12978,N_14042);
or U19966 (N_19966,N_11376,N_10771);
nor U19967 (N_19967,N_12392,N_14086);
or U19968 (N_19968,N_11322,N_11218);
or U19969 (N_19969,N_11118,N_10393);
and U19970 (N_19970,N_11258,N_14153);
xnor U19971 (N_19971,N_12229,N_11483);
and U19972 (N_19972,N_14521,N_10422);
nor U19973 (N_19973,N_11197,N_12556);
and U19974 (N_19974,N_14988,N_14768);
nand U19975 (N_19975,N_13939,N_14278);
or U19976 (N_19976,N_14445,N_14370);
xor U19977 (N_19977,N_11926,N_13207);
xor U19978 (N_19978,N_11150,N_12902);
xnor U19979 (N_19979,N_14210,N_13125);
nor U19980 (N_19980,N_13934,N_14598);
xor U19981 (N_19981,N_14582,N_13886);
nand U19982 (N_19982,N_14497,N_14606);
xor U19983 (N_19983,N_11885,N_14272);
xor U19984 (N_19984,N_12705,N_12869);
xor U19985 (N_19985,N_11861,N_10695);
or U19986 (N_19986,N_12028,N_10464);
and U19987 (N_19987,N_11348,N_14389);
nor U19988 (N_19988,N_13737,N_13581);
nor U19989 (N_19989,N_12459,N_12110);
and U19990 (N_19990,N_12088,N_13559);
nand U19991 (N_19991,N_11406,N_13474);
and U19992 (N_19992,N_10356,N_10842);
nand U19993 (N_19993,N_11520,N_14687);
nor U19994 (N_19994,N_11145,N_13368);
or U19995 (N_19995,N_14052,N_13104);
and U19996 (N_19996,N_14125,N_12393);
nor U19997 (N_19997,N_13627,N_12188);
nand U19998 (N_19998,N_14283,N_11966);
xor U19999 (N_19999,N_10523,N_10650);
and U20000 (N_20000,N_15273,N_17324);
nand U20001 (N_20001,N_18319,N_15869);
nor U20002 (N_20002,N_17530,N_17197);
or U20003 (N_20003,N_17274,N_17719);
nor U20004 (N_20004,N_19922,N_15089);
and U20005 (N_20005,N_18255,N_15978);
xor U20006 (N_20006,N_15636,N_16676);
and U20007 (N_20007,N_16782,N_18538);
nand U20008 (N_20008,N_15593,N_15909);
xor U20009 (N_20009,N_15166,N_16649);
nor U20010 (N_20010,N_19394,N_17373);
xnor U20011 (N_20011,N_16071,N_19968);
and U20012 (N_20012,N_17567,N_15729);
nor U20013 (N_20013,N_17890,N_16586);
or U20014 (N_20014,N_17370,N_19767);
or U20015 (N_20015,N_18049,N_18887);
nor U20016 (N_20016,N_16047,N_15497);
and U20017 (N_20017,N_17407,N_16240);
or U20018 (N_20018,N_18335,N_18279);
or U20019 (N_20019,N_17309,N_18326);
nand U20020 (N_20020,N_19954,N_17690);
or U20021 (N_20021,N_16791,N_17691);
xor U20022 (N_20022,N_19865,N_19761);
nor U20023 (N_20023,N_16143,N_18671);
nor U20024 (N_20024,N_16572,N_19817);
and U20025 (N_20025,N_18123,N_19385);
or U20026 (N_20026,N_17327,N_17910);
nor U20027 (N_20027,N_18657,N_15478);
xnor U20028 (N_20028,N_18509,N_18805);
nor U20029 (N_20029,N_15738,N_19484);
nor U20030 (N_20030,N_15227,N_18659);
nor U20031 (N_20031,N_19001,N_15706);
and U20032 (N_20032,N_16999,N_19542);
xor U20033 (N_20033,N_19032,N_15225);
xor U20034 (N_20034,N_15361,N_17047);
xnor U20035 (N_20035,N_19605,N_18185);
or U20036 (N_20036,N_18354,N_18639);
or U20037 (N_20037,N_18433,N_19552);
nor U20038 (N_20038,N_16723,N_16697);
nor U20039 (N_20039,N_18179,N_16687);
nand U20040 (N_20040,N_18737,N_17437);
xor U20041 (N_20041,N_15150,N_19169);
nor U20042 (N_20042,N_16952,N_18467);
and U20043 (N_20043,N_15237,N_17640);
xnor U20044 (N_20044,N_18209,N_18690);
nand U20045 (N_20045,N_17516,N_19438);
nand U20046 (N_20046,N_18940,N_15112);
and U20047 (N_20047,N_17716,N_17617);
nand U20048 (N_20048,N_16118,N_19979);
nand U20049 (N_20049,N_17646,N_18637);
or U20050 (N_20050,N_17702,N_19435);
xnor U20051 (N_20051,N_16756,N_15968);
xnor U20052 (N_20052,N_15580,N_19614);
or U20053 (N_20053,N_15291,N_18083);
nand U20054 (N_20054,N_17715,N_18833);
and U20055 (N_20055,N_16076,N_18660);
or U20056 (N_20056,N_19617,N_18807);
and U20057 (N_20057,N_15412,N_19720);
xnor U20058 (N_20058,N_16223,N_19769);
xnor U20059 (N_20059,N_16208,N_16961);
and U20060 (N_20060,N_19084,N_16006);
nor U20061 (N_20061,N_18156,N_19238);
nor U20062 (N_20062,N_17221,N_17749);
and U20063 (N_20063,N_19127,N_19983);
nand U20064 (N_20064,N_19192,N_15976);
nor U20065 (N_20065,N_16986,N_15325);
nor U20066 (N_20066,N_16082,N_16693);
xnor U20067 (N_20067,N_16979,N_18447);
and U20068 (N_20068,N_16144,N_15234);
xor U20069 (N_20069,N_17934,N_16343);
nand U20070 (N_20070,N_15376,N_16477);
or U20071 (N_20071,N_18563,N_16902);
and U20072 (N_20072,N_16413,N_15422);
or U20073 (N_20073,N_18856,N_17031);
or U20074 (N_20074,N_19715,N_16500);
or U20075 (N_20075,N_16157,N_18720);
xor U20076 (N_20076,N_16885,N_15456);
xor U20077 (N_20077,N_18851,N_15604);
nand U20078 (N_20078,N_19877,N_18970);
and U20079 (N_20079,N_17310,N_16179);
nor U20080 (N_20080,N_18625,N_15681);
xor U20081 (N_20081,N_15695,N_18468);
or U20082 (N_20082,N_17552,N_15193);
nor U20083 (N_20083,N_19670,N_15365);
nor U20084 (N_20084,N_15268,N_15929);
nand U20085 (N_20085,N_18967,N_19912);
and U20086 (N_20086,N_18161,N_17559);
or U20087 (N_20087,N_17081,N_18537);
or U20088 (N_20088,N_17494,N_17770);
and U20089 (N_20089,N_16570,N_15616);
nor U20090 (N_20090,N_19228,N_16142);
xnor U20091 (N_20091,N_17644,N_18489);
nand U20092 (N_20092,N_15798,N_16848);
or U20093 (N_20093,N_16169,N_18982);
xnor U20094 (N_20094,N_17215,N_18705);
or U20095 (N_20095,N_17829,N_15508);
xor U20096 (N_20096,N_18448,N_17103);
nand U20097 (N_20097,N_18608,N_18697);
and U20098 (N_20098,N_15094,N_16865);
xor U20099 (N_20099,N_15264,N_16149);
xor U20100 (N_20100,N_15534,N_17160);
nor U20101 (N_20101,N_18526,N_19258);
nand U20102 (N_20102,N_19647,N_18842);
xnor U20103 (N_20103,N_18175,N_18748);
xnor U20104 (N_20104,N_18847,N_17677);
xnor U20105 (N_20105,N_15667,N_19500);
and U20106 (N_20106,N_18614,N_15151);
nand U20107 (N_20107,N_18277,N_17734);
and U20108 (N_20108,N_17481,N_16613);
xor U20109 (N_20109,N_19694,N_17224);
nor U20110 (N_20110,N_18182,N_18774);
nand U20111 (N_20111,N_15334,N_16763);
and U20112 (N_20112,N_19994,N_15866);
or U20113 (N_20113,N_16721,N_15691);
xor U20114 (N_20114,N_18581,N_18871);
or U20115 (N_20115,N_16129,N_19477);
xnor U20116 (N_20116,N_19463,N_15028);
nor U20117 (N_20117,N_18477,N_17956);
nand U20118 (N_20118,N_15039,N_19990);
xor U20119 (N_20119,N_16573,N_15648);
nor U20120 (N_20120,N_19023,N_18337);
nor U20121 (N_20121,N_17433,N_19250);
xor U20122 (N_20122,N_16259,N_16060);
nor U20123 (N_20123,N_15609,N_18088);
or U20124 (N_20124,N_17245,N_16673);
nand U20125 (N_20125,N_17429,N_17882);
nand U20126 (N_20126,N_19585,N_19848);
nand U20127 (N_20127,N_15188,N_17776);
xor U20128 (N_20128,N_15296,N_16686);
nand U20129 (N_20129,N_15374,N_18595);
xnor U20130 (N_20130,N_18864,N_18997);
or U20131 (N_20131,N_19696,N_19285);
xnor U20132 (N_20132,N_17030,N_15625);
and U20133 (N_20133,N_19684,N_17460);
and U20134 (N_20134,N_16102,N_18874);
nor U20135 (N_20135,N_19952,N_19995);
and U20136 (N_20136,N_16376,N_18691);
and U20137 (N_20137,N_18663,N_19443);
nand U20138 (N_20138,N_17416,N_18907);
nand U20139 (N_20139,N_17326,N_16733);
nand U20140 (N_20140,N_18206,N_16631);
nand U20141 (N_20141,N_17529,N_18760);
and U20142 (N_20142,N_18305,N_15505);
nand U20143 (N_20143,N_16176,N_19150);
xnor U20144 (N_20144,N_16226,N_16850);
and U20145 (N_20145,N_16031,N_18309);
xor U20146 (N_20146,N_19704,N_15134);
xnor U20147 (N_20147,N_18945,N_16893);
and U20148 (N_20148,N_16725,N_18218);
xor U20149 (N_20149,N_15895,N_19388);
or U20150 (N_20150,N_15977,N_16053);
xor U20151 (N_20151,N_19945,N_18485);
and U20152 (N_20152,N_17408,N_19346);
xor U20153 (N_20153,N_15049,N_19279);
xor U20154 (N_20154,N_18293,N_17984);
nor U20155 (N_20155,N_16526,N_18572);
xor U20156 (N_20156,N_17780,N_17787);
xnor U20157 (N_20157,N_16136,N_16314);
or U20158 (N_20158,N_15198,N_17930);
nand U20159 (N_20159,N_18999,N_19075);
or U20160 (N_20160,N_17966,N_17392);
xnor U20161 (N_20161,N_17333,N_17187);
nand U20162 (N_20162,N_17152,N_16416);
or U20163 (N_20163,N_15860,N_15630);
or U20164 (N_20164,N_18883,N_18230);
or U20165 (N_20165,N_18109,N_19277);
and U20166 (N_20166,N_15520,N_15675);
and U20167 (N_20167,N_16451,N_15103);
and U20168 (N_20168,N_17122,N_18543);
and U20169 (N_20169,N_16207,N_15404);
nor U20170 (N_20170,N_19038,N_17551);
or U20171 (N_20171,N_17534,N_16213);
nand U20172 (N_20172,N_19368,N_17786);
or U20173 (N_20173,N_18002,N_16625);
xnor U20174 (N_20174,N_19008,N_18127);
or U20175 (N_20175,N_17410,N_18938);
or U20176 (N_20176,N_19861,N_17842);
and U20177 (N_20177,N_15913,N_18222);
xnor U20178 (N_20178,N_16010,N_18056);
nor U20179 (N_20179,N_15160,N_16701);
nand U20180 (N_20180,N_18456,N_18393);
nor U20181 (N_20181,N_17827,N_16890);
xnor U20182 (N_20182,N_17070,N_15135);
nand U20183 (N_20183,N_16985,N_18446);
nor U20184 (N_20184,N_17233,N_17057);
and U20185 (N_20185,N_19918,N_16998);
or U20186 (N_20186,N_17112,N_15360);
or U20187 (N_20187,N_17538,N_17574);
xor U20188 (N_20188,N_18895,N_15006);
xnor U20189 (N_20189,N_16846,N_19327);
nand U20190 (N_20190,N_19989,N_19702);
and U20191 (N_20191,N_18976,N_19188);
xor U20192 (N_20192,N_19129,N_18414);
nor U20193 (N_20193,N_15726,N_15770);
or U20194 (N_20194,N_15725,N_19022);
or U20195 (N_20195,N_17687,N_19316);
nor U20196 (N_20196,N_15889,N_17346);
nand U20197 (N_20197,N_19882,N_17709);
xnor U20198 (N_20198,N_19657,N_15692);
nor U20199 (N_20199,N_18269,N_19752);
or U20200 (N_20200,N_19849,N_15104);
and U20201 (N_20201,N_15437,N_15917);
or U20202 (N_20202,N_19413,N_19459);
nor U20203 (N_20203,N_18181,N_16228);
nor U20204 (N_20204,N_19935,N_16840);
nor U20205 (N_20205,N_17980,N_19747);
xnor U20206 (N_20206,N_16962,N_19690);
xnor U20207 (N_20207,N_17150,N_15179);
and U20208 (N_20208,N_16080,N_18108);
xnor U20209 (N_20209,N_17027,N_16069);
xor U20210 (N_20210,N_16964,N_19875);
xnor U20211 (N_20211,N_15776,N_19859);
or U20212 (N_20212,N_19183,N_16540);
xnor U20213 (N_20213,N_15984,N_16175);
nor U20214 (N_20214,N_17501,N_15221);
or U20215 (N_20215,N_17015,N_18324);
nor U20216 (N_20216,N_19687,N_18570);
or U20217 (N_20217,N_18115,N_17514);
and U20218 (N_20218,N_19019,N_19921);
and U20219 (N_20219,N_17847,N_18121);
nand U20220 (N_20220,N_17263,N_19399);
or U20221 (N_20221,N_15495,N_17158);
or U20222 (N_20222,N_19522,N_18104);
xnor U20223 (N_20223,N_19259,N_18102);
and U20224 (N_20224,N_15091,N_19051);
nor U20225 (N_20225,N_16162,N_16700);
xor U20226 (N_20226,N_15546,N_16014);
xnor U20227 (N_20227,N_16828,N_15473);
nor U20228 (N_20228,N_18184,N_16012);
xor U20229 (N_20229,N_16922,N_18942);
nand U20230 (N_20230,N_15285,N_18371);
and U20231 (N_20231,N_17859,N_19535);
xor U20232 (N_20232,N_15341,N_16432);
and U20233 (N_20233,N_15014,N_19158);
or U20234 (N_20234,N_18922,N_19886);
nor U20235 (N_20235,N_19932,N_19504);
nor U20236 (N_20236,N_18212,N_18726);
xor U20237 (N_20237,N_17051,N_15176);
and U20238 (N_20238,N_18172,N_18832);
xnor U20239 (N_20239,N_15849,N_18404);
nand U20240 (N_20240,N_16263,N_19637);
and U20241 (N_20241,N_16125,N_19962);
xor U20242 (N_20242,N_15346,N_15088);
or U20243 (N_20243,N_15133,N_19306);
nor U20244 (N_20244,N_19488,N_18521);
nand U20245 (N_20245,N_18149,N_16295);
xnor U20246 (N_20246,N_15541,N_19312);
nor U20247 (N_20247,N_16741,N_15059);
or U20248 (N_20248,N_19709,N_19205);
nor U20249 (N_20249,N_17190,N_16242);
and U20250 (N_20250,N_15253,N_16891);
xor U20251 (N_20251,N_19430,N_15511);
and U20252 (N_20252,N_17819,N_19703);
or U20253 (N_20253,N_17178,N_17121);
xor U20254 (N_20254,N_18954,N_18520);
xor U20255 (N_20255,N_18809,N_18263);
and U20256 (N_20256,N_16418,N_15287);
nor U20257 (N_20257,N_18507,N_19988);
nor U20258 (N_20258,N_17176,N_16659);
xor U20259 (N_20259,N_19831,N_17194);
xor U20260 (N_20260,N_16027,N_18364);
nand U20261 (N_20261,N_17356,N_16100);
nand U20262 (N_20262,N_18294,N_15572);
xor U20263 (N_20263,N_17174,N_16904);
xor U20264 (N_20264,N_17772,N_16220);
and U20265 (N_20265,N_18913,N_19785);
nor U20266 (N_20266,N_16443,N_18806);
nor U20267 (N_20267,N_17142,N_19380);
and U20268 (N_20268,N_19787,N_16735);
xnor U20269 (N_20269,N_19708,N_18965);
and U20270 (N_20270,N_18289,N_18267);
nor U20271 (N_20271,N_15766,N_19778);
and U20272 (N_20272,N_17556,N_18870);
and U20273 (N_20273,N_15836,N_16232);
or U20274 (N_20274,N_19819,N_17712);
nor U20275 (N_20275,N_15768,N_18486);
nor U20276 (N_20276,N_16488,N_15197);
nand U20277 (N_20277,N_17428,N_15174);
xor U20278 (N_20278,N_18273,N_19230);
nor U20279 (N_20279,N_15584,N_16387);
and U20280 (N_20280,N_19593,N_18139);
or U20281 (N_20281,N_18252,N_15010);
nor U20282 (N_20282,N_19378,N_15202);
nor U20283 (N_20283,N_17633,N_19403);
nor U20284 (N_20284,N_19701,N_16260);
or U20285 (N_20285,N_16534,N_17475);
and U20286 (N_20286,N_17541,N_19288);
or U20287 (N_20287,N_17074,N_19537);
or U20288 (N_20288,N_18441,N_15666);
nor U20289 (N_20289,N_18541,N_15207);
nor U20290 (N_20290,N_16678,N_19402);
or U20291 (N_20291,N_15102,N_15178);
or U20292 (N_20292,N_19664,N_16868);
xnor U20293 (N_20293,N_19253,N_18544);
nor U20294 (N_20294,N_16675,N_18710);
or U20295 (N_20295,N_15213,N_16373);
and U20296 (N_20296,N_18300,N_19397);
or U20297 (N_20297,N_15694,N_15704);
nand U20298 (N_20298,N_15186,N_18312);
nor U20299 (N_20299,N_16287,N_16899);
nor U20300 (N_20300,N_19634,N_19674);
and U20301 (N_20301,N_16331,N_19298);
nor U20302 (N_20302,N_17685,N_17650);
or U20303 (N_20303,N_18349,N_15639);
or U20304 (N_20304,N_17296,N_15382);
xor U20305 (N_20305,N_19592,N_19247);
and U20306 (N_20306,N_17595,N_17752);
and U20307 (N_20307,N_18491,N_16085);
nand U20308 (N_20308,N_19746,N_16078);
nor U20309 (N_20309,N_15079,N_16230);
or U20310 (N_20310,N_18611,N_16056);
and U20311 (N_20311,N_18196,N_15333);
xnor U20312 (N_20312,N_18885,N_19324);
and U20313 (N_20313,N_17608,N_19226);
or U20314 (N_20314,N_18037,N_15272);
and U20315 (N_20315,N_16005,N_17542);
or U20316 (N_20316,N_19748,N_17155);
or U20317 (N_20317,N_16249,N_16720);
nand U20318 (N_20318,N_15525,N_15923);
or U20319 (N_20319,N_15959,N_16235);
and U20320 (N_20320,N_19612,N_15757);
nand U20321 (N_20321,N_18063,N_16928);
nor U20322 (N_20322,N_17273,N_16475);
nor U20323 (N_20323,N_16320,N_16271);
nand U20324 (N_20324,N_17406,N_16640);
nor U20325 (N_20325,N_19619,N_19263);
or U20326 (N_20326,N_18910,N_17383);
and U20327 (N_20327,N_18615,N_16583);
xnor U20328 (N_20328,N_19879,N_18858);
nand U20329 (N_20329,N_17730,N_15395);
nand U20330 (N_20330,N_16087,N_16317);
nor U20331 (N_20331,N_18899,N_16728);
nor U20332 (N_20332,N_16272,N_18794);
nor U20333 (N_20333,N_18183,N_15689);
nor U20334 (N_20334,N_18060,N_16536);
nand U20335 (N_20335,N_19797,N_17483);
nor U20336 (N_20336,N_19853,N_17722);
nor U20337 (N_20337,N_17762,N_18952);
xor U20338 (N_20338,N_17200,N_19591);
nor U20339 (N_20339,N_18989,N_17396);
and U20340 (N_20340,N_19965,N_17974);
or U20341 (N_20341,N_15660,N_15850);
or U20342 (N_20342,N_18015,N_16576);
and U20343 (N_20343,N_18223,N_15686);
nand U20344 (N_20344,N_17331,N_18192);
xnor U20345 (N_20345,N_15925,N_17670);
nor U20346 (N_20346,N_15792,N_19362);
and U20347 (N_20347,N_17821,N_16760);
nor U20348 (N_20348,N_18853,N_19464);
nand U20349 (N_20349,N_15423,N_17905);
and U20350 (N_20350,N_19731,N_16296);
or U20351 (N_20351,N_17211,N_15516);
nor U20352 (N_20352,N_15979,N_16812);
and U20353 (N_20353,N_18042,N_17116);
and U20354 (N_20354,N_17012,N_19889);
nand U20355 (N_20355,N_18918,N_18709);
or U20356 (N_20356,N_17320,N_15410);
nand U20357 (N_20357,N_18167,N_16533);
nand U20358 (N_20358,N_18716,N_19085);
xor U20359 (N_20359,N_16286,N_17196);
xnor U20360 (N_20360,N_19901,N_18158);
and U20361 (N_20361,N_17700,N_16140);
nand U20362 (N_20362,N_17618,N_18009);
xor U20363 (N_20363,N_15489,N_15524);
or U20364 (N_20364,N_18022,N_18400);
or U20365 (N_20365,N_15779,N_18694);
and U20366 (N_20366,N_16004,N_16439);
xnor U20367 (N_20367,N_16363,N_15282);
or U20368 (N_20368,N_17886,N_18771);
and U20369 (N_20369,N_19110,N_17159);
xor U20370 (N_20370,N_17765,N_18376);
xor U20371 (N_20371,N_19938,N_18857);
xnor U20372 (N_20372,N_15761,N_19248);
xor U20373 (N_20373,N_16658,N_15783);
nor U20374 (N_20374,N_16344,N_15249);
or U20375 (N_20375,N_18189,N_19256);
xor U20376 (N_20376,N_17052,N_18490);
and U20377 (N_20377,N_15201,N_18873);
and U20378 (N_20378,N_17991,N_18107);
or U20379 (N_20379,N_17004,N_19622);
nor U20380 (N_20380,N_15055,N_17874);
or U20381 (N_20381,N_15989,N_15062);
or U20382 (N_20382,N_18266,N_16497);
and U20383 (N_20383,N_16975,N_17203);
or U20384 (N_20384,N_16983,N_19349);
or U20385 (N_20385,N_18262,N_18692);
or U20386 (N_20386,N_17405,N_18069);
or U20387 (N_20387,N_17896,N_15475);
nor U20388 (N_20388,N_19723,N_19620);
or U20389 (N_20389,N_16872,N_15309);
nand U20390 (N_20390,N_15125,N_18131);
and U20391 (N_20391,N_19265,N_19329);
nand U20392 (N_20392,N_15279,N_15311);
nor U20393 (N_20393,N_15357,N_17117);
or U20394 (N_20394,N_16245,N_16114);
xnor U20395 (N_20395,N_16467,N_17621);
nand U20396 (N_20396,N_19598,N_17773);
and U20397 (N_20397,N_17841,N_17627);
nor U20398 (N_20398,N_15522,N_19314);
xnor U20399 (N_20399,N_19341,N_18631);
or U20400 (N_20400,N_19013,N_18078);
and U20401 (N_20401,N_17989,N_18401);
nor U20402 (N_20402,N_17334,N_15251);
and U20403 (N_20403,N_15269,N_18213);
and U20404 (N_20404,N_18367,N_19271);
xnor U20405 (N_20405,N_16219,N_16178);
nor U20406 (N_20406,N_16771,N_16474);
nor U20407 (N_20407,N_16730,N_19146);
or U20408 (N_20408,N_15023,N_15187);
and U20409 (N_20409,N_16943,N_18318);
xnor U20410 (N_20410,N_17885,N_15741);
xor U20411 (N_20411,N_17347,N_16861);
or U20412 (N_20412,N_19303,N_16106);
nor U20413 (N_20413,N_15631,N_18817);
nor U20414 (N_20414,N_16332,N_16486);
and U20415 (N_20415,N_18351,N_18203);
nand U20416 (N_20416,N_18238,N_19232);
or U20417 (N_20417,N_17492,N_16581);
or U20418 (N_20418,N_15915,N_16281);
xnor U20419 (N_20419,N_16426,N_16601);
nor U20420 (N_20420,N_18087,N_17319);
nand U20421 (N_20421,N_16553,N_19427);
and U20422 (N_20422,N_18609,N_19959);
or U20423 (N_20423,N_15995,N_18540);
xnor U20424 (N_20424,N_19212,N_15370);
xor U20425 (N_20425,N_19342,N_15470);
and U20426 (N_20426,N_19676,N_18068);
and U20427 (N_20427,N_15229,N_15068);
or U20428 (N_20428,N_18464,N_19523);
nand U20429 (N_20429,N_17413,N_19718);
nor U20430 (N_20430,N_17115,N_18141);
nor U20431 (N_20431,N_16339,N_19320);
xnor U20432 (N_20432,N_16966,N_17629);
and U20433 (N_20433,N_19958,N_17335);
xnor U20434 (N_20434,N_15332,N_18610);
nor U20435 (N_20435,N_19642,N_16137);
and U20436 (N_20436,N_16304,N_17948);
and U20437 (N_20437,N_19097,N_15687);
nor U20438 (N_20438,N_18408,N_15673);
nor U20439 (N_20439,N_15244,N_16099);
or U20440 (N_20440,N_15956,N_15228);
or U20441 (N_20441,N_15057,N_16013);
xor U20442 (N_20442,N_18834,N_18778);
xnor U20443 (N_20443,N_18018,N_16973);
and U20444 (N_20444,N_17459,N_15420);
nor U20445 (N_20445,N_18453,N_18148);
and U20446 (N_20446,N_16982,N_17915);
nand U20447 (N_20447,N_15809,N_18302);
xnor U20448 (N_20448,N_17083,N_18484);
and U20449 (N_20449,N_15999,N_17997);
or U20450 (N_20450,N_15339,N_19207);
nor U20451 (N_20451,N_19616,N_18850);
and U20452 (N_20452,N_15937,N_18765);
nor U20453 (N_20453,N_17435,N_15119);
nand U20454 (N_20454,N_17132,N_15363);
nand U20455 (N_20455,N_19832,N_19297);
or U20456 (N_20456,N_16022,N_15231);
nand U20457 (N_20457,N_18035,N_18514);
nand U20458 (N_20458,N_19509,N_18536);
and U20459 (N_20459,N_15621,N_18390);
nand U20460 (N_20460,N_19025,N_19291);
xnor U20461 (N_20461,N_16935,N_16117);
nor U20462 (N_20462,N_19469,N_17880);
xnor U20463 (N_20463,N_19215,N_15303);
or U20464 (N_20464,N_19375,N_19643);
and U20465 (N_20465,N_19119,N_19090);
and U20466 (N_20466,N_17402,N_18398);
and U20467 (N_20467,N_16411,N_15814);
nand U20468 (N_20468,N_17258,N_19417);
xnor U20469 (N_20469,N_16103,N_17018);
and U20470 (N_20470,N_16268,N_17314);
or U20471 (N_20471,N_16064,N_16374);
and U20472 (N_20472,N_18144,N_19573);
xnor U20473 (N_20473,N_17614,N_19360);
nand U20474 (N_20474,N_16378,N_17119);
or U20475 (N_20475,N_19985,N_16769);
nor U20476 (N_20476,N_15901,N_15816);
or U20477 (N_20477,N_16968,N_17423);
and U20478 (N_20478,N_18225,N_16599);
xnor U20479 (N_20479,N_17144,N_15192);
nor U20480 (N_20480,N_17707,N_16616);
xor U20481 (N_20481,N_17511,N_16299);
or U20482 (N_20482,N_19186,N_19982);
nor U20483 (N_20483,N_17533,N_16476);
or U20484 (N_20484,N_16446,N_16264);
and U20485 (N_20485,N_17041,N_15787);
nand U20486 (N_20486,N_19412,N_17486);
nand U20487 (N_20487,N_19784,N_17342);
or U20488 (N_20488,N_18126,N_17061);
nor U20489 (N_20489,N_16662,N_18296);
and U20490 (N_20490,N_19911,N_18641);
nand U20491 (N_20491,N_19757,N_17705);
and U20492 (N_20492,N_18437,N_15784);
xor U20493 (N_20493,N_17313,N_18622);
and U20494 (N_20494,N_18689,N_15204);
nor U20495 (N_20495,N_19623,N_16250);
or U20496 (N_20496,N_19960,N_17751);
xor U20497 (N_20497,N_15718,N_17971);
and U20498 (N_20498,N_15419,N_15550);
nor U20499 (N_20499,N_18169,N_16712);
nand U20500 (N_20500,N_17942,N_16550);
xor U20501 (N_20501,N_17286,N_19914);
nand U20502 (N_20502,N_16200,N_15946);
nor U20503 (N_20503,N_18800,N_18191);
nand U20504 (N_20504,N_17240,N_19781);
nor U20505 (N_20505,N_15751,N_19017);
and U20506 (N_20506,N_17815,N_19028);
xor U20507 (N_20507,N_18784,N_18308);
or U20508 (N_20508,N_17937,N_19024);
nand U20509 (N_20509,N_17875,N_17728);
nand U20510 (N_20510,N_17293,N_15808);
xor U20511 (N_20511,N_17171,N_19147);
and U20512 (N_20512,N_15483,N_19373);
or U20513 (N_20513,N_16822,N_17732);
xnor U20514 (N_20514,N_18943,N_18812);
xor U20515 (N_20515,N_16564,N_17639);
nor U20516 (N_20516,N_15206,N_18996);
and U20517 (N_20517,N_19118,N_18506);
nor U20518 (N_20518,N_18772,N_16774);
nand U20519 (N_20519,N_17778,N_18380);
nor U20520 (N_20520,N_17305,N_19162);
or U20521 (N_20521,N_19045,N_16753);
xnor U20522 (N_20522,N_15371,N_17596);
and U20523 (N_20523,N_19707,N_18993);
or U20524 (N_20524,N_15566,N_15459);
or U20525 (N_20525,N_16750,N_16894);
nand U20526 (N_20526,N_18823,N_18450);
and U20527 (N_20527,N_15945,N_18487);
or U20528 (N_20528,N_15000,N_18915);
nor U20529 (N_20529,N_17104,N_17216);
nor U20530 (N_20530,N_16306,N_15713);
xor U20531 (N_20531,N_17065,N_16514);
and U20532 (N_20532,N_16650,N_15313);
or U20533 (N_20533,N_19937,N_18808);
nand U20534 (N_20534,N_18299,N_16496);
nand U20535 (N_20535,N_15843,N_16450);
xor U20536 (N_20536,N_17816,N_15782);
nor U20537 (N_20537,N_18329,N_15343);
xor U20538 (N_20538,N_17445,N_15355);
nand U20539 (N_20539,N_15677,N_18966);
nand U20540 (N_20540,N_15185,N_19734);
and U20541 (N_20541,N_17040,N_18884);
nand U20542 (N_20542,N_18419,N_15710);
xor U20543 (N_20543,N_19340,N_16185);
nor U20544 (N_20544,N_15805,N_18229);
xnor U20545 (N_20545,N_18596,N_15997);
nand U20546 (N_20546,N_18640,N_16410);
or U20547 (N_20547,N_15868,N_16766);
and U20548 (N_20548,N_18136,N_17118);
and U20549 (N_20549,N_15015,N_17105);
xor U20550 (N_20550,N_18143,N_18457);
nor U20551 (N_20551,N_18178,N_16291);
or U20552 (N_20552,N_17427,N_17080);
nor U20553 (N_20553,N_16748,N_17518);
nor U20554 (N_20554,N_19421,N_15467);
and U20555 (N_20555,N_16180,N_17175);
xnor U20556 (N_20556,N_18407,N_19943);
or U20557 (N_20557,N_15670,N_16194);
and U20558 (N_20558,N_17059,N_16008);
nor U20559 (N_20559,N_18561,N_18846);
and U20560 (N_20560,N_16941,N_15693);
xnor U20561 (N_20561,N_19508,N_17055);
nand U20562 (N_20562,N_15013,N_18438);
nand U20563 (N_20563,N_15607,N_17350);
or U20564 (N_20564,N_17126,N_16987);
xnor U20565 (N_20565,N_17557,N_16847);
nand U20566 (N_20566,N_17724,N_17382);
nor U20567 (N_20567,N_19538,N_15862);
and U20568 (N_20568,N_16120,N_19763);
nand U20569 (N_20569,N_19867,N_15340);
nor U20570 (N_20570,N_17733,N_16279);
xnor U20571 (N_20571,N_15987,N_17237);
or U20572 (N_20572,N_17035,N_15480);
nand U20573 (N_20573,N_19191,N_16124);
nor U20574 (N_20574,N_19174,N_16589);
and U20575 (N_20575,N_15994,N_15629);
nand U20576 (N_20576,N_16566,N_19857);
nand U20577 (N_20577,N_17001,N_15400);
or U20578 (N_20578,N_17999,N_16772);
and U20579 (N_20579,N_19574,N_15304);
or U20580 (N_20580,N_18227,N_18950);
xor U20581 (N_20581,N_16646,N_19244);
xnor U20582 (N_20582,N_19292,N_15708);
and U20583 (N_20583,N_18499,N_17688);
and U20584 (N_20584,N_19583,N_17811);
xnor U20585 (N_20585,N_17218,N_18958);
nand U20586 (N_20586,N_15884,N_19142);
nor U20587 (N_20587,N_17862,N_19126);
or U20588 (N_20588,N_15139,N_17545);
nand U20589 (N_20589,N_17301,N_18416);
xnor U20590 (N_20590,N_19406,N_17050);
or U20591 (N_20591,N_17214,N_17272);
nor U20592 (N_20592,N_17371,N_16866);
and U20593 (N_20593,N_15444,N_15705);
xor U20594 (N_20594,N_15832,N_19262);
and U20595 (N_20595,N_17806,N_19020);
xnor U20596 (N_20596,N_15157,N_19284);
or U20597 (N_20597,N_15763,N_17694);
nand U20598 (N_20598,N_15949,N_15634);
nand U20599 (N_20599,N_17863,N_15403);
nor U20600 (N_20600,N_15449,N_18937);
and U20601 (N_20601,N_16019,N_19980);
nand U20602 (N_20602,N_17894,N_16995);
xnor U20603 (N_20603,N_19845,N_16384);
xnor U20604 (N_20604,N_15942,N_17513);
nor U20605 (N_20605,N_18236,N_16335);
or U20606 (N_20606,N_16382,N_15839);
or U20607 (N_20607,N_19227,N_15211);
nor U20608 (N_20608,N_15671,N_16542);
or U20609 (N_20609,N_17978,N_19776);
or U20610 (N_20610,N_18550,N_16171);
xor U20611 (N_20611,N_18916,N_19495);
or U20612 (N_20612,N_17758,N_17208);
or U20613 (N_20613,N_15690,N_19479);
nand U20614 (N_20614,N_16844,N_15031);
nand U20615 (N_20615,N_18723,N_15430);
and U20616 (N_20616,N_19554,N_18429);
nor U20617 (N_20617,N_18936,N_18759);
nand U20618 (N_20618,N_18946,N_17610);
nand U20619 (N_20619,N_15684,N_16367);
nor U20620 (N_20620,N_16048,N_15672);
nand U20621 (N_20621,N_15822,N_15728);
nand U20622 (N_20622,N_19821,N_18796);
nor U20623 (N_20623,N_17161,N_16541);
nor U20624 (N_20624,N_19041,N_15820);
xnor U20625 (N_20625,N_15171,N_15337);
or U20626 (N_20626,N_16420,N_16632);
nor U20627 (N_20627,N_19499,N_17498);
xnor U20628 (N_20628,N_18677,N_17926);
nand U20629 (N_20629,N_18046,N_17876);
nand U20630 (N_20630,N_18524,N_15804);
xor U20631 (N_20631,N_15683,N_18281);
xnor U20632 (N_20632,N_17704,N_16234);
nand U20633 (N_20633,N_19468,N_17790);
or U20634 (N_20634,N_16801,N_17870);
nand U20635 (N_20635,N_17357,N_16127);
or U20636 (N_20636,N_15571,N_18552);
nor U20637 (N_20637,N_16342,N_19446);
or U20638 (N_20638,N_18177,N_19266);
or U20639 (N_20639,N_15394,N_17663);
and U20640 (N_20640,N_17101,N_16372);
or U20641 (N_20641,N_19765,N_15443);
nor U20642 (N_20642,N_19482,N_19740);
xor U20643 (N_20643,N_16447,N_19996);
nor U20644 (N_20644,N_18297,N_16907);
and U20645 (N_20645,N_17284,N_16293);
and U20646 (N_20646,N_18330,N_15754);
and U20647 (N_20647,N_18105,N_16824);
xor U20648 (N_20648,N_19947,N_19418);
xnor U20649 (N_20649,N_15238,N_19700);
and U20650 (N_20650,N_19059,N_17927);
and U20651 (N_20651,N_17450,N_15380);
and U20652 (N_20652,N_18317,N_19037);
nand U20653 (N_20653,N_16364,N_15071);
and U20654 (N_20654,N_17365,N_17631);
or U20655 (N_20655,N_16088,N_19206);
nor U20656 (N_20656,N_16729,N_17395);
xor U20657 (N_20657,N_16752,N_16857);
nand U20658 (N_20658,N_19473,N_15111);
nor U20659 (N_20659,N_18815,N_16449);
nor U20660 (N_20660,N_16284,N_19425);
or U20661 (N_20661,N_19931,N_16579);
nor U20662 (N_20662,N_15299,N_15105);
nor U20663 (N_20663,N_19693,N_18355);
or U20664 (N_20664,N_19128,N_18522);
or U20665 (N_20665,N_15722,N_15848);
or U20666 (N_20666,N_17093,N_18855);
nand U20667 (N_20667,N_18642,N_15256);
and U20668 (N_20668,N_19739,N_19987);
xnor U20669 (N_20669,N_19946,N_19728);
nand U20670 (N_20670,N_15329,N_16626);
xor U20671 (N_20671,N_16635,N_16380);
xor U20672 (N_20672,N_19727,N_15938);
nor U20673 (N_20673,N_16531,N_19040);
nor U20674 (N_20674,N_16133,N_16517);
nand U20675 (N_20675,N_18341,N_17389);
xnor U20676 (N_20676,N_17199,N_17021);
or U20677 (N_20677,N_17680,N_19280);
xnor U20678 (N_20678,N_18844,N_18980);
nor U20679 (N_20679,N_19168,N_18264);
nand U20680 (N_20680,N_18712,N_16130);
and U20681 (N_20681,N_19208,N_16487);
xor U20682 (N_20682,N_15696,N_19249);
or U20683 (N_20683,N_18542,N_19109);
or U20684 (N_20684,N_19138,N_15554);
and U20685 (N_20685,N_15418,N_16222);
xor U20686 (N_20686,N_17456,N_18841);
xnor U20687 (N_20687,N_18298,N_16933);
and U20688 (N_20688,N_15501,N_16164);
or U20689 (N_20689,N_17329,N_16183);
nor U20690 (N_20690,N_15876,N_16406);
xor U20691 (N_20691,N_15196,N_16537);
and U20692 (N_20692,N_19511,N_19007);
xor U20693 (N_20693,N_16978,N_19636);
xor U20694 (N_20694,N_19540,N_15599);
and U20695 (N_20695,N_19078,N_18579);
and U20696 (N_20696,N_19758,N_17801);
xnor U20697 (N_20697,N_15819,N_19762);
nor U20698 (N_20698,N_18512,N_16093);
or U20699 (N_20699,N_16307,N_17693);
nor U20700 (N_20700,N_15426,N_18322);
and U20701 (N_20701,N_16837,N_17539);
or U20702 (N_20702,N_17796,N_18280);
and U20703 (N_20703,N_19915,N_17332);
nand U20704 (N_20704,N_19582,N_18556);
nand U20705 (N_20705,N_16021,N_18460);
and U20706 (N_20706,N_18919,N_17911);
and U20707 (N_20707,N_16838,N_17441);
nor U20708 (N_20708,N_16726,N_18802);
nor U20709 (N_20709,N_19489,N_16211);
xnor U20710 (N_20710,N_18199,N_18578);
xor U20711 (N_20711,N_16815,N_17028);
or U20712 (N_20712,N_17289,N_19252);
nor U20713 (N_20713,N_19193,N_18242);
nand U20714 (N_20714,N_17519,N_16009);
nand U20715 (N_20715,N_19649,N_19677);
xor U20716 (N_20716,N_15411,N_17570);
or U20717 (N_20717,N_16956,N_15985);
nand U20718 (N_20718,N_16161,N_18819);
and U20719 (N_20719,N_18670,N_17607);
xor U20720 (N_20720,N_16876,N_16490);
nand U20721 (N_20721,N_19596,N_19374);
and U20722 (N_20722,N_19555,N_19201);
and U20723 (N_20723,N_17579,N_15128);
or U20724 (N_20724,N_19426,N_18866);
xor U20725 (N_20725,N_16839,N_15391);
xor U20726 (N_20726,N_19351,N_16043);
or U20727 (N_20727,N_17897,N_17944);
nor U20728 (N_20728,N_16833,N_17785);
nor U20729 (N_20729,N_18652,N_18811);
and U20730 (N_20730,N_17271,N_19184);
or U20731 (N_20731,N_17869,N_17189);
nor U20732 (N_20732,N_16593,N_18669);
or U20733 (N_20733,N_19928,N_17461);
nor U20734 (N_20734,N_16094,N_15762);
or U20735 (N_20735,N_18674,N_19895);
nor U20736 (N_20736,N_16755,N_15887);
nand U20737 (N_20737,N_16623,N_17630);
nand U20738 (N_20738,N_19029,N_17647);
or U20739 (N_20739,N_15081,N_19348);
nor U20740 (N_20740,N_15998,N_16860);
nand U20741 (N_20741,N_16600,N_16045);
nand U20742 (N_20742,N_18052,N_19369);
xnor U20743 (N_20743,N_16911,N_15295);
xor U20744 (N_20744,N_17771,N_16917);
nand U20745 (N_20745,N_17452,N_17544);
or U20746 (N_20746,N_16595,N_18385);
or U20747 (N_20747,N_15297,N_19107);
nor U20748 (N_20748,N_16414,N_18868);
or U20749 (N_20749,N_16942,N_19630);
nand U20750 (N_20750,N_18743,N_18459);
and U20751 (N_20751,N_19153,N_17959);
nand U20752 (N_20752,N_15930,N_18244);
and U20753 (N_20753,N_19713,N_18635);
or U20754 (N_20754,N_19423,N_17537);
or U20755 (N_20755,N_17257,N_15858);
and U20756 (N_20756,N_18010,N_16381);
xnor U20757 (N_20757,N_16326,N_18738);
nor U20758 (N_20758,N_16854,N_19735);
nor U20759 (N_20759,N_17602,N_16571);
and U20760 (N_20760,N_17140,N_17170);
or U20761 (N_20761,N_15800,N_19833);
xor U20762 (N_20762,N_15723,N_18029);
and U20763 (N_20763,N_16400,N_17718);
nand U20764 (N_20764,N_16377,N_15632);
or U20765 (N_20765,N_15935,N_15336);
or U20766 (N_20766,N_18623,N_18496);
nor U20767 (N_20767,N_18575,N_17916);
nand U20768 (N_20768,N_18031,N_17086);
nor U20769 (N_20769,N_15320,N_16867);
xnor U20770 (N_20770,N_17855,N_18732);
or U20771 (N_20771,N_18041,N_18064);
xnor U20772 (N_20772,N_18565,N_17184);
or U20773 (N_20773,N_17804,N_19214);
or U20774 (N_20774,N_15903,N_16493);
xor U20775 (N_20775,N_16025,N_18903);
and U20776 (N_20776,N_16327,N_19419);
and U20777 (N_20777,N_19217,N_17128);
and U20778 (N_20778,N_18605,N_16328);
xnor U20779 (N_20779,N_15236,N_19775);
and U20780 (N_20780,N_15540,N_17699);
nor U20781 (N_20781,N_15921,N_16813);
nor U20782 (N_20782,N_16802,N_18933);
and U20783 (N_20783,N_16218,N_15659);
or U20784 (N_20784,N_18198,N_17753);
and U20785 (N_20785,N_18113,N_19662);
and U20786 (N_20786,N_18948,N_19866);
nor U20787 (N_20787,N_16453,N_16912);
and U20788 (N_20788,N_17735,N_19345);
and U20789 (N_20789,N_16777,N_17438);
nor U20790 (N_20790,N_19669,N_19382);
or U20791 (N_20791,N_17750,N_16465);
and U20792 (N_20792,N_19149,N_15349);
nand U20793 (N_20793,N_15398,N_19561);
nand U20794 (N_20794,N_18099,N_18384);
nor U20795 (N_20795,N_17078,N_17512);
nand U20796 (N_20796,N_15442,N_17562);
nor U20797 (N_20797,N_16324,N_19810);
nor U20798 (N_20798,N_18742,N_19828);
and U20799 (N_20799,N_17102,N_17737);
nand U20800 (N_20800,N_18831,N_19898);
or U20801 (N_20801,N_19520,N_18114);
or U20802 (N_20802,N_15771,N_19944);
nor U20803 (N_20803,N_16612,N_17060);
nor U20804 (N_20804,N_16680,N_15812);
or U20805 (N_20805,N_16804,N_15864);
nand U20806 (N_20806,N_18981,N_18436);
nor U20807 (N_20807,N_18430,N_17943);
nand U20808 (N_20808,N_16026,N_18892);
nand U20809 (N_20809,N_18119,N_16724);
xnor U20810 (N_20810,N_16582,N_16544);
xor U20811 (N_20811,N_17739,N_19251);
and U20812 (N_20812,N_15758,N_15920);
nor U20813 (N_20813,N_15801,N_16641);
or U20814 (N_20814,N_17649,N_18247);
nand U20815 (N_20815,N_18173,N_18788);
and U20816 (N_20816,N_15981,N_17443);
and U20817 (N_20817,N_17604,N_17269);
nor U20818 (N_20818,N_18128,N_16530);
or U20819 (N_20819,N_17763,N_15290);
xor U20820 (N_20820,N_15538,N_17246);
or U20821 (N_20821,N_16483,N_15928);
or U20822 (N_20822,N_15595,N_16858);
nor U20823 (N_20823,N_15248,N_18235);
nor U20824 (N_20824,N_19387,N_15138);
nand U20825 (N_20825,N_15388,N_15589);
or U20826 (N_20826,N_19571,N_16492);
or U20827 (N_20827,N_16528,N_18232);
nand U20828 (N_20828,N_19347,N_15975);
or U20829 (N_20829,N_17823,N_18271);
nand U20830 (N_20830,N_16826,N_15200);
xnor U20831 (N_20831,N_15092,N_18444);
or U20832 (N_20832,N_17798,N_17419);
nor U20833 (N_20833,N_15471,N_17540);
and U20834 (N_20834,N_18908,N_16892);
nor U20835 (N_20835,N_16189,N_18389);
nand U20836 (N_20836,N_18483,N_17384);
nand U20837 (N_20837,N_16809,N_17368);
or U20838 (N_20838,N_17839,N_19551);
and U20839 (N_20839,N_18515,N_16206);
or U20840 (N_20840,N_19553,N_17738);
nor U20841 (N_20841,N_18339,N_19840);
xor U20842 (N_20842,N_19286,N_19680);
and U20843 (N_20843,N_17830,N_18224);
nor U20844 (N_20844,N_15328,N_17954);
nand U20845 (N_20845,N_19719,N_16193);
xor U20846 (N_20846,N_19530,N_18804);
or U20847 (N_20847,N_15402,N_16166);
xnor U20848 (N_20848,N_17345,N_19472);
nor U20849 (N_20849,N_19160,N_15326);
and U20850 (N_20850,N_18685,N_19926);
xor U20851 (N_20851,N_17799,N_19152);
xnor U20852 (N_20852,N_16525,N_15306);
or U20853 (N_20853,N_15399,N_18315);
or U20854 (N_20854,N_15011,N_19454);
and U20855 (N_20855,N_16661,N_15778);
or U20856 (N_20856,N_19282,N_18566);
nor U20857 (N_20857,N_17376,N_18435);
and U20858 (N_20858,N_18684,N_18208);
and U20859 (N_20859,N_17442,N_18643);
nand U20860 (N_20860,N_18180,N_18654);
xnor U20861 (N_20861,N_18399,N_18835);
or U20862 (N_20862,N_19624,N_18551);
xor U20863 (N_20863,N_19940,N_15324);
nand U20864 (N_20864,N_19744,N_15646);
and U20865 (N_20865,N_16415,N_17462);
and U20866 (N_20866,N_17125,N_18379);
xor U20867 (N_20867,N_16276,N_18062);
or U20868 (N_20868,N_17044,N_19791);
and U20869 (N_20869,N_19350,N_17071);
and U20870 (N_20870,N_17403,N_15226);
or U20871 (N_20871,N_19120,N_19948);
and U20872 (N_20872,N_19311,N_15067);
nand U20873 (N_20873,N_15026,N_15739);
xnor U20874 (N_20874,N_18363,N_16970);
and U20875 (N_20875,N_19145,N_15955);
nor U20876 (N_20876,N_17163,N_17351);
nand U20877 (N_20877,N_16174,N_15153);
nor U20878 (N_20878,N_16785,N_16398);
and U20879 (N_20879,N_15844,N_15093);
nand U20880 (N_20880,N_15257,N_18053);
xnor U20881 (N_20881,N_18043,N_16895);
and U20882 (N_20882,N_17094,N_19475);
nand U20883 (N_20883,N_15058,N_17096);
or U20884 (N_20884,N_17803,N_18769);
xor U20885 (N_20885,N_17660,N_18795);
xor U20886 (N_20886,N_17560,N_18134);
or U20887 (N_20887,N_15649,N_16805);
nor U20888 (N_20888,N_18207,N_15029);
nand U20889 (N_20889,N_17409,N_15002);
or U20890 (N_20890,N_15742,N_19722);
nor U20891 (N_20891,N_18651,N_16743);
xor U20892 (N_20892,N_18095,N_18854);
xor U20893 (N_20893,N_15679,N_15702);
xor U20894 (N_20894,N_17777,N_16329);
or U20895 (N_20895,N_17168,N_15856);
xor U20896 (N_20896,N_16011,N_18987);
nor U20897 (N_20897,N_18734,N_15733);
and U20898 (N_20898,N_17487,N_17290);
xnor U20899 (N_20899,N_18012,N_17504);
or U20900 (N_20900,N_19269,N_18394);
or U20901 (N_20901,N_17259,N_16835);
and U20902 (N_20902,N_17895,N_18116);
nor U20903 (N_20903,N_19759,N_19491);
and U20904 (N_20904,N_16141,N_15549);
nand U20905 (N_20905,N_16421,N_19487);
or U20906 (N_20906,N_15662,N_16796);
nor U20907 (N_20907,N_16560,N_18036);
nand U20908 (N_20908,N_19505,N_16736);
xnor U20909 (N_20909,N_19313,N_19939);
nand U20910 (N_20910,N_17490,N_18386);
nor U20911 (N_20911,N_16302,N_17756);
or U20912 (N_20912,N_17935,N_16460);
xnor U20913 (N_20913,N_17056,N_19756);
nor U20914 (N_20914,N_16303,N_19294);
and U20915 (N_20915,N_19272,N_18562);
or U20916 (N_20916,N_17338,N_16003);
nand U20917 (N_20917,N_17131,N_16879);
nor U20918 (N_20918,N_19173,N_19907);
and U20919 (N_20919,N_17861,N_17588);
nor U20920 (N_20920,N_16489,N_16637);
and U20921 (N_20921,N_15130,N_15218);
xor U20922 (N_20922,N_17281,N_15818);
and U20923 (N_20923,N_15281,N_17020);
nor U20924 (N_20924,N_19497,N_15190);
and U20925 (N_20925,N_18097,N_17039);
nand U20926 (N_20926,N_18140,N_16549);
xnor U20927 (N_20927,N_17820,N_19971);
and U20928 (N_20928,N_18476,N_19981);
and U20929 (N_20929,N_18701,N_15265);
and U20930 (N_20930,N_17976,N_19543);
nand U20931 (N_20931,N_17098,N_19239);
xnor U20932 (N_20932,N_16734,N_18889);
nor U20933 (N_20933,N_17181,N_17264);
nand U20934 (N_20934,N_18995,N_18574);
xor U20935 (N_20935,N_17521,N_19321);
xor U20936 (N_20936,N_17774,N_16934);
or U20937 (N_20937,N_17814,N_15933);
xor U20938 (N_20938,N_19531,N_15740);
nor U20939 (N_20939,N_18226,N_18055);
nand U20940 (N_20940,N_16630,N_18332);
xor U20941 (N_20941,N_16706,N_18632);
nand U20942 (N_20942,N_18445,N_17953);
nand U20943 (N_20943,N_18194,N_15548);
and U20944 (N_20944,N_15642,N_19692);
nand U20945 (N_20945,N_17397,N_17465);
or U20946 (N_20946,N_15474,N_15472);
nor U20947 (N_20947,N_19381,N_18347);
nand U20948 (N_20948,N_19799,N_17067);
nand U20949 (N_20949,N_17575,N_19261);
or U20950 (N_20950,N_18843,N_16024);
nand U20951 (N_20951,N_18424,N_18681);
xor U20952 (N_20952,N_16265,N_17252);
and U20953 (N_20953,N_19071,N_18118);
nor U20954 (N_20954,N_16318,N_18284);
xnor U20955 (N_20955,N_19629,N_17477);
nand U20956 (N_20956,N_18786,N_18975);
xnor U20957 (N_20957,N_15170,N_19235);
or U20958 (N_20958,N_16927,N_16574);
xnor U20959 (N_20959,N_18333,N_16463);
or U20960 (N_20960,N_16471,N_18849);
nor U20961 (N_20961,N_19519,N_19366);
and U20962 (N_20962,N_19367,N_18142);
or U20963 (N_20963,N_16681,N_16016);
xnor U20964 (N_20964,N_16385,N_18790);
nand U20965 (N_20965,N_18528,N_17697);
or U20966 (N_20966,N_19453,N_16058);
and U20967 (N_20967,N_15943,N_15359);
xnor U20968 (N_20968,N_16561,N_15352);
or U20969 (N_20969,N_19114,N_19827);
and U20970 (N_20970,N_16028,N_19782);
or U20971 (N_20971,N_17362,N_16588);
nand U20972 (N_20972,N_16154,N_16798);
and U20973 (N_20973,N_16762,N_18612);
xnor U20974 (N_20974,N_17550,N_15567);
nor U20975 (N_20975,N_19372,N_18073);
nand U20976 (N_20976,N_17328,N_16587);
or U20977 (N_20977,N_15040,N_15840);
nand U20978 (N_20978,N_16437,N_15066);
nand U20979 (N_20979,N_18100,N_18250);
and U20980 (N_20980,N_15647,N_19796);
xnor U20981 (N_20981,N_18733,N_17077);
or U20982 (N_20982,N_15537,N_15498);
xnor U20983 (N_20983,N_18470,N_16862);
or U20984 (N_20984,N_17303,N_18342);
or U20985 (N_20985,N_18545,N_19117);
nor U20986 (N_20986,N_17717,N_17589);
and U20987 (N_20987,N_19950,N_17451);
nand U20988 (N_20988,N_16300,N_16072);
and U20989 (N_20989,N_18529,N_18050);
nand U20990 (N_20990,N_19695,N_16543);
nor U20991 (N_20991,N_19673,N_15137);
xnor U20992 (N_20992,N_18629,N_18890);
xnor U20993 (N_20993,N_15601,N_17932);
nor U20994 (N_20994,N_18475,N_17755);
nor U20995 (N_20995,N_19414,N_15278);
or U20996 (N_20996,N_18969,N_17768);
nand U20997 (N_20997,N_17587,N_15753);
nand U20998 (N_20998,N_16823,N_17635);
and U20999 (N_20999,N_15970,N_17287);
xnor U21000 (N_21000,N_15148,N_15069);
or U21001 (N_21001,N_17185,N_16551);
or U21002 (N_21002,N_18439,N_18283);
nand U21003 (N_21003,N_18549,N_18863);
and U21004 (N_21004,N_15891,N_18508);
nor U21005 (N_21005,N_15877,N_15076);
nand U21006 (N_21006,N_16217,N_15330);
xnor U21007 (N_21007,N_17023,N_17641);
xnor U21008 (N_21008,N_19565,N_19501);
nand U21009 (N_21009,N_16032,N_18523);
xnor U21010 (N_21010,N_19726,N_19604);
and U21011 (N_21011,N_18789,N_16951);
or U21012 (N_21012,N_19344,N_17234);
or U21013 (N_21013,N_19302,N_15875);
nor U21014 (N_21014,N_15857,N_19481);
or U21015 (N_21015,N_17068,N_19595);
nor U21016 (N_21016,N_19904,N_15532);
nand U21017 (N_21017,N_18725,N_16945);
and U21018 (N_21018,N_18160,N_19976);
or U21019 (N_21019,N_17291,N_15050);
nand U21020 (N_21020,N_16539,N_17133);
nor U21021 (N_21021,N_18034,N_19264);
nand U21022 (N_21022,N_19813,N_17134);
nor U21023 (N_21023,N_16212,N_19104);
nor U21024 (N_21024,N_15254,N_16417);
nor U21025 (N_21025,N_17464,N_15208);
nand U21026 (N_21026,N_17476,N_19668);
nand U21027 (N_21027,N_15791,N_17495);
or U21028 (N_21028,N_18164,N_15276);
xor U21029 (N_21029,N_18584,N_15060);
or U21030 (N_21030,N_19255,N_16221);
nand U21031 (N_21031,N_18696,N_15199);
nand U21032 (N_21032,N_15181,N_17833);
nand U21033 (N_21033,N_17344,N_16994);
xor U21034 (N_21034,N_16900,N_18288);
nand U21035 (N_21035,N_19838,N_16989);
and U21036 (N_21036,N_15308,N_16007);
nand U21037 (N_21037,N_18735,N_16282);
or U21038 (N_21038,N_17270,N_17256);
or U21039 (N_21039,N_15707,N_16065);
nor U21040 (N_21040,N_16992,N_19590);
xnor U21041 (N_21041,N_19790,N_16191);
nand U21042 (N_21042,N_19854,N_16225);
nor U21043 (N_21043,N_16135,N_18214);
and U21044 (N_21044,N_18443,N_16814);
or U21045 (N_21045,N_15957,N_19030);
nand U21046 (N_21046,N_18481,N_19766);
xor U21047 (N_21047,N_17312,N_16074);
or U21048 (N_21048,N_16897,N_17340);
or U21049 (N_21049,N_17527,N_16580);
nor U21050 (N_21050,N_15774,N_16116);
or U21051 (N_21051,N_17123,N_19156);
or U21052 (N_21052,N_18604,N_19563);
and U21053 (N_21053,N_19607,N_18350);
nand U21054 (N_21054,N_16333,N_17167);
xnor U21055 (N_21055,N_16555,N_18274);
and U21056 (N_21056,N_19897,N_17526);
and U21057 (N_21057,N_16097,N_19179);
and U21058 (N_21058,N_15597,N_16508);
xnor U21059 (N_21059,N_19716,N_19383);
nand U21060 (N_21060,N_17446,N_17138);
nand U21061 (N_21061,N_15656,N_17970);
or U21062 (N_21062,N_16851,N_16972);
and U21063 (N_21063,N_15083,N_18675);
and U21064 (N_21064,N_16464,N_17455);
xor U21065 (N_21065,N_16527,N_17235);
nand U21066 (N_21066,N_16128,N_18471);
and U21067 (N_21067,N_16310,N_17166);
nor U21068 (N_21068,N_18220,N_17090);
nor U21069 (N_21069,N_18075,N_19697);
xor U21070 (N_21070,N_16253,N_16829);
xnor U21071 (N_21071,N_15298,N_19474);
or U21072 (N_21072,N_19871,N_18900);
nor U21073 (N_21073,N_15543,N_19492);
and U21074 (N_21074,N_19997,N_18962);
and U21075 (N_21075,N_16841,N_15396);
or U21076 (N_21076,N_15793,N_18146);
xor U21077 (N_21077,N_17729,N_19236);
or U21078 (N_21078,N_19768,N_18941);
nor U21079 (N_21079,N_18947,N_15841);
nand U21080 (N_21080,N_17924,N_16170);
nor U21081 (N_21081,N_18886,N_15961);
and U21082 (N_21082,N_17157,N_17673);
xnor U21083 (N_21083,N_18821,N_15633);
and U21084 (N_21084,N_18362,N_16988);
nor U21085 (N_21085,N_16611,N_18106);
or U21086 (N_21086,N_16388,N_17149);
or U21087 (N_21087,N_19199,N_17708);
nor U21088 (N_21088,N_19141,N_16251);
or U21089 (N_21089,N_18497,N_18994);
or U21090 (N_21090,N_18111,N_19197);
nor U21091 (N_21091,N_19287,N_19356);
and U21092 (N_21092,N_15143,N_18103);
or U21093 (N_21093,N_19627,N_19920);
nand U21094 (N_21094,N_19820,N_18020);
xnor U21095 (N_21095,N_18934,N_18649);
xnor U21096 (N_21096,N_15477,N_16205);
xnor U21097 (N_21097,N_18781,N_16050);
nor U21098 (N_21098,N_18211,N_17469);
nor U21099 (N_21099,N_15678,N_19850);
nor U21100 (N_21100,N_19073,N_15056);
nor U21101 (N_21101,N_16598,N_19518);
nand U21102 (N_21102,N_18585,N_18559);
nand U21103 (N_21103,N_18708,N_18613);
and U21104 (N_21104,N_17262,N_19364);
nor U21105 (N_21105,N_18797,N_16757);
and U21106 (N_21106,N_16916,N_19749);
or U21107 (N_21107,N_18766,N_19672);
or U21108 (N_21108,N_17720,N_18421);
or U21109 (N_21109,N_16552,N_16423);
xnor U21110 (N_21110,N_18602,N_18534);
or U21111 (N_21111,N_17436,N_16355);
and U21112 (N_21112,N_15453,N_19541);
nand U21113 (N_21113,N_17424,N_18260);
and U21114 (N_21114,N_15246,N_18495);
nand U21115 (N_21115,N_16821,N_16605);
xor U21116 (N_21116,N_16946,N_17912);
xnor U21117 (N_21117,N_19974,N_19410);
nor U21118 (N_21118,N_16375,N_15338);
nor U21119 (N_21119,N_17108,N_18894);
nor U21120 (N_21120,N_18661,N_16903);
nor U21121 (N_21121,N_16156,N_16789);
nor U21122 (N_21122,N_19774,N_17871);
nor U21123 (N_21123,N_17899,N_16369);
nand U21124 (N_21124,N_17917,N_15073);
or U21125 (N_21125,N_18348,N_19633);
or U21126 (N_21126,N_17993,N_16122);
xnor U21127 (N_21127,N_16499,N_15815);
nand U21128 (N_21128,N_19490,N_19586);
xor U21129 (N_21129,N_15893,N_15061);
nor U21130 (N_21130,N_17212,N_16518);
xor U21131 (N_21131,N_19163,N_19587);
xor U21132 (N_21132,N_19476,N_16620);
nor U21133 (N_21133,N_16955,N_17921);
nand U21134 (N_21134,N_15168,N_19076);
xor U21135 (N_21135,N_17981,N_17619);
nor U21136 (N_21136,N_15233,N_19486);
nor U21137 (N_21137,N_16412,N_18749);
xor U21138 (N_21138,N_19112,N_16930);
or U21139 (N_21139,N_16285,N_18747);
and U21140 (N_21140,N_17606,N_18406);
and U21141 (N_21141,N_15379,N_19194);
nor U21142 (N_21142,N_19103,N_17580);
and U21143 (N_21143,N_19441,N_18321);
and U21144 (N_21144,N_16925,N_18906);
or U21145 (N_21145,N_16652,N_18730);
or U21146 (N_21146,N_18278,N_15159);
xor U21147 (N_21147,N_16288,N_15947);
nand U21148 (N_21148,N_15585,N_18422);
nor U21149 (N_21149,N_19798,N_19743);
xor U21150 (N_21150,N_15986,N_19326);
or U21151 (N_21151,N_18129,N_19113);
or U21152 (N_21152,N_19539,N_19074);
nor U21153 (N_21153,N_17219,N_18065);
xnor U21154 (N_21154,N_17792,N_17714);
or U21155 (N_21155,N_19337,N_16231);
and U21156 (N_21156,N_16991,N_17229);
nand U21157 (N_21157,N_19544,N_15243);
nor U21158 (N_21158,N_17592,N_15223);
or U21159 (N_21159,N_18428,N_19283);
nand U21160 (N_21160,N_19639,N_19658);
and U21161 (N_21161,N_18479,N_16356);
nand U21162 (N_21162,N_19391,N_19400);
and U21163 (N_21163,N_15885,N_17813);
or U21164 (N_21164,N_16081,N_19532);
nand U21165 (N_21165,N_15164,N_19396);
nand U21166 (N_21166,N_16323,N_15775);
nand U21167 (N_21167,N_18673,N_17339);
and U21168 (N_21168,N_17110,N_17034);
and U21169 (N_21169,N_17584,N_19231);
or U21170 (N_21170,N_18683,N_18546);
nand U21171 (N_21171,N_15063,N_15096);
xor U21172 (N_21172,N_15115,N_16196);
xor U21173 (N_21173,N_15517,N_15777);
xnor U21174 (N_21174,N_17076,N_19290);
or U21175 (N_21175,N_19220,N_17986);
nand U21176 (N_21176,N_19884,N_15267);
nor U21177 (N_21177,N_18130,N_18243);
xor U21178 (N_21178,N_18353,N_16657);
and U21179 (N_21179,N_17919,N_19824);
nand U21180 (N_21180,N_18869,N_18826);
or U21181 (N_21181,N_17945,N_15375);
or U21182 (N_21182,N_17951,N_16722);
or U21183 (N_21183,N_19547,N_17434);
and U21184 (N_21184,N_15644,N_19072);
or U21185 (N_21185,N_15911,N_19336);
nand U21186 (N_21186,N_17892,N_19986);
nand U21187 (N_21187,N_17522,N_17359);
and U21188 (N_21188,N_19467,N_17835);
and U21189 (N_21189,N_19930,N_18058);
nand U21190 (N_21190,N_16929,N_16096);
and U21191 (N_21191,N_19485,N_15491);
and U21192 (N_21192,N_16622,N_18261);
nand U21193 (N_21193,N_16873,N_19641);
or U21194 (N_21194,N_15027,N_19144);
nor U21195 (N_21195,N_16864,N_18314);
nor U21196 (N_21196,N_17854,N_18228);
xnor U21197 (N_21197,N_16308,N_18717);
xnor U21198 (N_21198,N_15606,N_18216);
and U21199 (N_21199,N_19010,N_17849);
and U21200 (N_21200,N_17482,N_16454);
xor U21201 (N_21201,N_19771,N_18646);
xnor U21202 (N_21202,N_16280,N_19353);
nand U21203 (N_21203,N_15515,N_15241);
nand U21204 (N_21204,N_18193,N_16997);
nor U21205 (N_21205,N_15824,N_16820);
nor U21206 (N_21206,N_15965,N_18992);
nand U21207 (N_21207,N_16690,N_16091);
or U21208 (N_21208,N_19730,N_15559);
nor U21209 (N_21209,N_15888,N_19745);
nor U21210 (N_21210,N_15465,N_17220);
xor U21211 (N_21211,N_18162,N_17524);
nor U21212 (N_21212,N_16430,N_15496);
xor U21213 (N_21213,N_18233,N_17995);
xor U21214 (N_21214,N_15528,N_18902);
nand U21215 (N_21215,N_18047,N_17038);
or U21216 (N_21216,N_16448,N_19046);
or U21217 (N_21217,N_18859,N_17568);
and U21218 (N_21218,N_16799,N_18656);
nand U21219 (N_21219,N_16698,N_16111);
xor U21220 (N_21220,N_15542,N_16442);
nand U21221 (N_21221,N_19788,N_18827);
nor U21222 (N_21222,N_16098,N_16294);
nand U21223 (N_21223,N_16949,N_17360);
or U21224 (N_21224,N_18814,N_15788);
nor U21225 (N_21225,N_19416,N_15372);
or U21226 (N_21226,N_18359,N_18626);
nand U21227 (N_21227,N_18955,N_19480);
or U21228 (N_21228,N_17298,N_16685);
or U21229 (N_21229,N_15007,N_15640);
xor U21230 (N_21230,N_19031,N_17472);
and U21231 (N_21231,N_18017,N_16792);
or U21232 (N_21232,N_15810,N_16113);
nand U21233 (N_21233,N_17931,N_15535);
nor U21234 (N_21234,N_18564,N_15764);
xnor U21235 (N_21235,N_19742,N_17572);
xor U21236 (N_21236,N_16313,N_16940);
and U21237 (N_21237,N_19067,N_16779);
or U21238 (N_21238,N_16428,N_16609);
nor U21239 (N_21239,N_17420,N_18893);
and U21240 (N_21240,N_15924,N_18171);
and U21241 (N_21241,N_18555,N_19011);
or U21242 (N_21242,N_19237,N_17883);
and U21243 (N_21243,N_19737,N_15993);
xnor U21244 (N_21244,N_16749,N_16434);
nor U21245 (N_21245,N_15736,N_18676);
or U21246 (N_21246,N_18027,N_19653);
or U21247 (N_21247,N_18929,N_17058);
xnor U21248 (N_21248,N_17788,N_19036);
nand U21249 (N_21249,N_16563,N_17085);
xor U21250 (N_21250,N_15122,N_18200);
xor U21251 (N_21251,N_17887,N_18603);
xnor U21252 (N_21252,N_18449,N_19826);
xor U21253 (N_21253,N_18357,N_16195);
or U21254 (N_21254,N_18124,N_17581);
nand U21255 (N_21255,N_19999,N_15136);
nand U21256 (N_21256,N_18245,N_15712);
nor U21257 (N_21257,N_16073,N_17769);
nand U21258 (N_21258,N_17665,N_19594);
nand U21259 (N_21259,N_17754,N_15799);
or U21260 (N_21260,N_18852,N_17253);
nand U21261 (N_21261,N_19896,N_18248);
xor U21262 (N_21262,N_15413,N_16654);
and U21263 (N_21263,N_16107,N_16554);
nand U21264 (N_21264,N_19015,N_17097);
xor U21265 (N_21265,N_17226,N_19754);
xnor U21266 (N_21266,N_16974,N_16651);
nand U21267 (N_21267,N_16371,N_17900);
nand U21268 (N_21268,N_17748,N_15610);
nor U21269 (N_21269,N_19056,N_16029);
and U21270 (N_21270,N_18588,N_15499);
nand U21271 (N_21271,N_19415,N_18860);
and U21272 (N_21272,N_16341,N_16038);
or U21273 (N_21273,N_16719,N_17440);
nor U21274 (N_21274,N_18715,N_18829);
and U21275 (N_21275,N_19780,N_15141);
nand U21276 (N_21276,N_19568,N_19328);
xnor U21277 (N_21277,N_19562,N_17766);
or U21278 (N_21278,N_15882,N_15446);
xor U21279 (N_21279,N_18822,N_19978);
nor U21280 (N_21280,N_17994,N_16515);
xor U21281 (N_21281,N_16520,N_19471);
nand U21282 (N_21282,N_16139,N_15397);
nor U21283 (N_21283,N_19267,N_19837);
nor U21284 (N_21284,N_17497,N_16151);
and U21285 (N_21285,N_16472,N_15389);
and U21286 (N_21286,N_18077,N_15932);
or U21287 (N_21287,N_18197,N_16389);
nand U21288 (N_21288,N_15912,N_19923);
xnor U21289 (N_21289,N_15663,N_19082);
xnor U21290 (N_21290,N_19517,N_17369);
xnor U21291 (N_21291,N_18480,N_15556);
and U21292 (N_21292,N_15428,N_16309);
nand U21293 (N_21293,N_18039,N_18310);
nand U21294 (N_21294,N_15558,N_19445);
nand U21295 (N_21295,N_19154,N_17198);
nor U21296 (N_21296,N_18093,N_16738);
and U21297 (N_21297,N_18008,N_17757);
nand U21298 (N_21298,N_16513,N_17449);
nand U21299 (N_21299,N_19172,N_17913);
and U21300 (N_21300,N_19166,N_16519);
nor U21301 (N_21301,N_16731,N_17669);
and U21302 (N_21302,N_18478,N_19829);
or U21303 (N_21303,N_17620,N_19710);
nand U21304 (N_21304,N_19420,N_15482);
nor U21305 (N_21305,N_15036,N_17278);
nor U21306 (N_21306,N_15126,N_19100);
and U21307 (N_21307,N_16672,N_16386);
nor U21308 (N_21308,N_19157,N_16123);
or U21309 (N_21309,N_18465,N_19209);
or U21310 (N_21310,N_19159,N_16322);
or U21311 (N_21311,N_17439,N_19164);
nand U21312 (N_21312,N_18383,N_18425);
nor U21313 (N_21313,N_17826,N_17597);
nand U21314 (N_21314,N_16184,N_19524);
xnor U21315 (N_21315,N_18770,N_19009);
xnor U21316 (N_21316,N_18589,N_15401);
nand U21317 (N_21317,N_17130,N_16419);
nand U21318 (N_21318,N_17844,N_17251);
and U21319 (N_21319,N_17230,N_16505);
nand U21320 (N_21320,N_16521,N_19610);
nor U21321 (N_21321,N_17622,N_19601);
xor U21322 (N_21322,N_15020,N_16037);
or U21323 (N_21323,N_16764,N_16522);
and U21324 (N_21324,N_17531,N_16504);
or U21325 (N_21325,N_18378,N_16905);
or U21326 (N_21326,N_15469,N_15385);
xor U21327 (N_21327,N_17283,N_15072);
xor U21328 (N_21328,N_16849,N_15090);
or U21329 (N_21329,N_17232,N_15051);
nand U21330 (N_21330,N_18998,N_15033);
and U21331 (N_21331,N_17013,N_16391);
nand U21332 (N_21332,N_15878,N_16896);
nand U21333 (N_21333,N_19021,N_17210);
nand U21334 (N_21334,N_17037,N_16436);
nand U21335 (N_21335,N_17300,N_19318);
nand U21336 (N_21336,N_18074,N_18875);
xor U21337 (N_21337,N_16379,N_18678);
xor U21338 (N_21338,N_16671,N_18331);
nand U21339 (N_21339,N_18944,N_19807);
nor U21340 (N_21340,N_15175,N_19578);
xnor U21341 (N_21341,N_18375,N_17285);
nor U21342 (N_21342,N_18358,N_18092);
nand U21343 (N_21343,N_17805,N_19844);
or U21344 (N_21344,N_17664,N_15087);
and U21345 (N_21345,N_16901,N_19223);
xor U21346 (N_21346,N_18234,N_17740);
nand U21347 (N_21347,N_17600,N_15106);
nand U21348 (N_21348,N_18427,N_19855);
xor U21349 (N_21349,N_16797,N_15927);
nor U21350 (N_21350,N_18724,N_15132);
xor U21351 (N_21351,N_16708,N_15255);
nor U21352 (N_21352,N_15991,N_15655);
xnor U21353 (N_21353,N_16350,N_17394);
and U21354 (N_21354,N_16146,N_15124);
xor U21355 (N_21355,N_17393,N_17025);
xnor U21356 (N_21356,N_17636,N_19814);
nand U21357 (N_21357,N_17277,N_19068);
xor U21358 (N_21358,N_17398,N_16485);
nor U21359 (N_21359,N_18023,N_17679);
or U21360 (N_21360,N_19770,N_15650);
nand U21361 (N_21361,N_16887,N_16262);
or U21362 (N_21362,N_18527,N_17352);
xor U21363 (N_21363,N_19094,N_18066);
nor U21364 (N_21364,N_19494,N_15828);
and U21365 (N_21365,N_18410,N_18911);
xor U21366 (N_21366,N_17426,N_17092);
xnor U21367 (N_21367,N_18072,N_16906);
nand U21368 (N_21368,N_15874,N_16051);
or U21369 (N_21369,N_16404,N_19825);
or U21370 (N_21370,N_17488,N_15366);
or U21371 (N_21371,N_18006,N_18256);
nor U21372 (N_21372,N_15462,N_17611);
xnor U21373 (N_21373,N_15351,N_17571);
xor U21374 (N_21374,N_17207,N_18241);
xnor U21375 (N_21375,N_18361,N_19873);
nand U21376 (N_21376,N_18474,N_18828);
xnor U21377 (N_21377,N_16699,N_16248);
or U21378 (N_21378,N_15509,N_19361);
nand U21379 (N_21379,N_15075,N_17379);
nand U21380 (N_21380,N_19786,N_18699);
nor U21381 (N_21381,N_15466,N_16607);
nor U21382 (N_21382,N_16246,N_15641);
xor U21383 (N_21383,N_19870,N_18620);
nand U21384 (N_21384,N_18577,N_16158);
nor U21385 (N_21385,N_15427,N_16878);
and U21386 (N_21386,N_16182,N_17960);
xnor U21387 (N_21387,N_18598,N_15526);
nor U21388 (N_21388,N_17793,N_16855);
xor U21389 (N_21389,N_19878,N_18098);
nor U21390 (N_21390,N_16237,N_19012);
nor U21391 (N_21391,N_19370,N_18094);
and U21392 (N_21392,N_17601,N_19992);
and U21393 (N_21393,N_15685,N_16845);
xnor U21394 (N_21394,N_16075,N_15668);
nor U21395 (N_21395,N_19755,N_15969);
xnor U21396 (N_21396,N_17202,N_18702);
xor U21397 (N_21397,N_18753,N_15645);
nand U21398 (N_21398,N_17241,N_19908);
xnor U21399 (N_21399,N_18714,N_17165);
or U21400 (N_21400,N_17837,N_18345);
nand U21401 (N_21401,N_17553,N_16963);
or U21402 (N_21402,N_17651,N_19613);
nor U21403 (N_21403,N_15046,N_16819);
and U21404 (N_21404,N_16244,N_16834);
nor U21405 (N_21405,N_17616,N_16863);
nand U21406 (N_21406,N_18594,N_17907);
xnor U21407 (N_21407,N_18897,N_19970);
nand U21408 (N_21408,N_17247,N_15582);
xnor U21409 (N_21409,N_19305,N_19432);
and U21410 (N_21410,N_15345,N_17191);
and U21411 (N_21411,N_19964,N_16629);
and U21412 (N_21412,N_15082,N_16269);
and U21413 (N_21413,N_15883,N_19052);
or U21414 (N_21414,N_17248,N_17817);
nand U21415 (N_21415,N_17789,N_17390);
nand U21416 (N_21416,N_18369,N_15951);
xor U21417 (N_21417,N_16888,N_16759);
or U21418 (N_21418,N_16319,N_15676);
or U21419 (N_21419,N_16660,N_18905);
or U21420 (N_21420,N_15865,N_17517);
xnor U21421 (N_21421,N_17010,N_16298);
and U21422 (N_21422,N_18086,N_16340);
nand U21423 (N_21423,N_17479,N_15658);
nand U21424 (N_21424,N_19683,N_18306);
or U21425 (N_21425,N_18925,N_16780);
and U21426 (N_21426,N_16954,N_19204);
nor U21427 (N_21427,N_16702,N_17139);
nand U21428 (N_21428,N_19513,N_17846);
and U21429 (N_21429,N_19424,N_16215);
nor U21430 (N_21430,N_17032,N_16252);
xor U21431 (N_21431,N_16063,N_16209);
or U21432 (N_21432,N_17583,N_18038);
nor U21433 (N_21433,N_17852,N_18040);
and U21434 (N_21434,N_17447,N_15384);
xnor U21435 (N_21435,N_18431,N_19392);
nand U21436 (N_21436,N_16913,N_19338);
nor U21437 (N_21437,N_16575,N_18728);
xnor U21438 (N_21438,N_19106,N_19606);
nor U21439 (N_21439,N_15619,N_17988);
and U21440 (N_21440,N_16615,N_15806);
xnor U21441 (N_21441,N_17355,N_16131);
nand U21442 (N_21442,N_18792,N_17471);
nor U21443 (N_21443,N_17593,N_16761);
or U21444 (N_21444,N_18466,N_18328);
or U21445 (N_21445,N_18210,N_16811);
or U21446 (N_21446,N_18653,N_15488);
xor U21447 (N_21447,N_16345,N_19431);
and U21448 (N_21448,N_18787,N_15854);
nor U21449 (N_21449,N_17710,N_18879);
or U21450 (N_21450,N_19175,N_15765);
nor U21451 (N_21451,N_19408,N_16089);
xor U21452 (N_21452,N_19116,N_19567);
xor U21453 (N_21453,N_16957,N_19450);
xor U21454 (N_21454,N_15250,N_18510);
or U21455 (N_21455,N_15025,N_16273);
and U21456 (N_21456,N_19760,N_18985);
or U21457 (N_21457,N_17146,N_18202);
nand U21458 (N_21458,N_16810,N_16938);
or U21459 (N_21459,N_16643,N_18352);
and U21460 (N_21460,N_17064,N_16795);
nor U21461 (N_21461,N_17063,N_19088);
xnor U21462 (N_21462,N_17418,N_16301);
nor U21463 (N_21463,N_15414,N_16482);
or U21464 (N_21464,N_18001,N_18991);
xnor U21465 (N_21465,N_17642,N_16441);
and U21466 (N_21466,N_15724,N_19065);
nor U21467 (N_21467,N_18259,N_15457);
and U21468 (N_21468,N_15169,N_16751);
nor U21469 (N_21469,N_18307,N_19688);
xnor U21470 (N_21470,N_16173,N_16034);
nand U21471 (N_21471,N_18695,N_18591);
xnor U21472 (N_21472,N_19377,N_16177);
and U21473 (N_21473,N_16617,N_15919);
nor U21474 (N_21474,N_17491,N_16592);
xor U21475 (N_21475,N_19883,N_16204);
or U21476 (N_21476,N_19625,N_19608);
or U21477 (N_21477,N_17682,N_17043);
nor U21478 (N_21478,N_18569,N_16667);
and U21479 (N_21479,N_18513,N_17742);
and U21480 (N_21480,N_19458,N_16603);
xor U21481 (N_21481,N_18548,N_16466);
nor U21482 (N_21482,N_19478,N_16030);
nand U21483 (N_21483,N_18700,N_18170);
xnor U21484 (N_21484,N_16110,N_19039);
and U21485 (N_21485,N_19393,N_17547);
and U21486 (N_21486,N_19246,N_17510);
nand U21487 (N_21487,N_18026,N_17091);
xnor U21488 (N_21488,N_19101,N_17005);
nor U21489 (N_21489,N_17908,N_17850);
nor U21490 (N_21490,N_15870,N_15431);
nand U21491 (N_21491,N_18346,N_17213);
and U21492 (N_21492,N_17188,N_18432);
nor U21493 (N_21493,N_18275,N_15966);
nor U21494 (N_21494,N_19685,N_17007);
or U21495 (N_21495,N_19219,N_16353);
and U21496 (N_21496,N_17949,N_19717);
nand U21497 (N_21497,N_15561,N_18462);
nand U21498 (N_21498,N_17925,N_15147);
or U21499 (N_21499,N_18775,N_16694);
nand U21500 (N_21500,N_17414,N_16842);
nand U21501 (N_21501,N_18750,N_18593);
or U21502 (N_21502,N_15626,N_18557);
xnor U21503 (N_21503,N_16095,N_15172);
and U21504 (N_21504,N_17979,N_19631);
or U21505 (N_21505,N_19584,N_16608);
nor U21506 (N_21506,N_19442,N_19182);
and U21507 (N_21507,N_16656,N_17502);
nor U21508 (N_21508,N_17000,N_17901);
nand U21509 (N_21509,N_19779,N_15405);
xor U21510 (N_21510,N_19890,N_19880);
or U21511 (N_21511,N_19894,N_16800);
nand U21512 (N_21512,N_17145,N_16444);
or U21513 (N_21513,N_19661,N_16236);
or U21514 (N_21514,N_15004,N_15703);
nor U21515 (N_21515,N_16104,N_16150);
nor U21516 (N_21516,N_18320,N_17380);
or U21517 (N_21517,N_17661,N_18744);
or U21518 (N_21518,N_16545,N_18000);
nor U21519 (N_21519,N_16257,N_16624);
and U21520 (N_21520,N_15510,N_15117);
xnor U21521 (N_21521,N_19270,N_15409);
nand U21522 (N_21522,N_15583,N_19176);
nor U21523 (N_21523,N_19016,N_15972);
xnor U21524 (N_21524,N_19864,N_18370);
or U21525 (N_21525,N_19556,N_17676);
nand U21526 (N_21526,N_15415,N_19243);
nor U21527 (N_21527,N_17828,N_17569);
xor U21528 (N_21528,N_15831,N_18163);
and U21529 (N_21529,N_15258,N_19900);
nand U21530 (N_21530,N_15240,N_17865);
and U21531 (N_21531,N_17453,N_18081);
nand U21532 (N_21532,N_18024,N_16258);
or U21533 (N_21533,N_16562,N_16397);
and U21534 (N_21534,N_15527,N_16547);
nor U21535 (N_21535,N_17135,N_17458);
nor U21536 (N_21536,N_16931,N_19437);
or U21537 (N_21537,N_18898,N_18968);
and U21538 (N_21538,N_16939,N_15195);
nor U21539 (N_21539,N_16655,N_18877);
and U21540 (N_21540,N_17888,N_15588);
and U21541 (N_21541,N_15441,N_19404);
and U21542 (N_21542,N_15570,N_18839);
and U21543 (N_21543,N_19333,N_15813);
nor U21544 (N_21544,N_17808,N_18336);
nand U21545 (N_21545,N_18838,N_18014);
xnor U21546 (N_21546,N_16703,N_15288);
nand U21547 (N_21547,N_18762,N_16510);
nand U21548 (N_21548,N_18567,N_19398);
and U21549 (N_21549,N_15900,N_17902);
nand U21550 (N_21550,N_19211,N_15845);
xor U21551 (N_21551,N_18862,N_15358);
and U21552 (N_21552,N_18773,N_19502);
and U21553 (N_21553,N_19365,N_17615);
or U21554 (N_21554,N_16480,N_19632);
nor U21555 (N_21555,N_18469,N_18951);
xor U21556 (N_21556,N_17268,N_17546);
xor U21557 (N_21557,N_19822,N_19738);
xor U21558 (N_21558,N_15086,N_19549);
or U21559 (N_21559,N_15605,N_19165);
nand U21560 (N_21560,N_15458,N_16790);
nand U21561 (N_21561,N_16677,N_16875);
and U21562 (N_21562,N_15194,N_19171);
nor U21563 (N_21563,N_19801,N_19783);
and U21564 (N_21564,N_15454,N_19626);
xnor U21565 (N_21565,N_16882,N_18295);
and U21566 (N_21566,N_17325,N_19576);
nand U21567 (N_21567,N_17599,N_18721);
nand U21568 (N_21568,N_16886,N_18756);
and U21569 (N_21569,N_15078,N_16337);
nand U21570 (N_21570,N_18888,N_19200);
xor U21571 (N_21571,N_16165,N_15100);
nand U21572 (N_21572,N_18599,N_19339);
nand U21573 (N_21573,N_19679,N_15180);
nand U21574 (N_21574,N_19609,N_17818);
nand U21575 (N_21575,N_17940,N_18286);
or U21576 (N_21576,N_15730,N_19916);
or U21577 (N_21577,N_19648,N_16105);
or U21578 (N_21578,N_17689,N_18583);
nor U21579 (N_21579,N_15688,N_15224);
and U21580 (N_21580,N_18201,N_19714);
nand U21581 (N_21581,N_16077,N_17467);
xnor U21582 (N_21582,N_17594,N_16704);
nor U21583 (N_21583,N_15035,N_15144);
nand U21584 (N_21584,N_18500,N_19917);
nor U21585 (N_21585,N_17543,N_19275);
and U21586 (N_21586,N_17415,N_17425);
or U21587 (N_21587,N_19611,N_17147);
or U21588 (N_21588,N_18215,N_15613);
nor U21589 (N_21589,N_18867,N_15097);
nand U21590 (N_21590,N_17977,N_16057);
and U21591 (N_21591,N_16336,N_15377);
xor U21592 (N_21592,N_19027,N_15165);
nor U21593 (N_21593,N_18865,N_16843);
nor U21594 (N_21594,N_19122,N_18882);
and U21595 (N_21595,N_18494,N_16948);
or U21596 (N_21596,N_18921,N_18204);
nor U21597 (N_21597,N_17653,N_15344);
nand U21598 (N_21598,N_16457,N_17612);
or U21599 (N_21599,N_19803,N_18059);
xor U21600 (N_21600,N_17723,N_17950);
and U21601 (N_21601,N_19102,N_18780);
nand U21602 (N_21602,N_16002,N_18754);
nand U21603 (N_21603,N_15881,N_17323);
nand U21604 (N_21604,N_16684,N_18272);
xor U21605 (N_21605,N_18876,N_16108);
xor U21606 (N_21606,N_17444,N_18782);
xnor U21607 (N_21607,N_19615,N_16424);
xnor U21608 (N_21608,N_15958,N_16818);
nor U21609 (N_21609,N_16977,N_15873);
nor U21610 (N_21610,N_18688,N_19891);
nor U21611 (N_21611,N_17288,N_17082);
or U21612 (N_21612,N_18667,N_15608);
and U21613 (N_21613,N_17231,N_16768);
or U21614 (N_21614,N_16524,N_15432);
nand U21615 (N_21615,N_15120,N_15189);
or U21616 (N_21616,N_19210,N_18645);
and U21617 (N_21617,N_18374,N_19973);
or U21618 (N_21618,N_19315,N_18757);
and U21619 (N_21619,N_15564,N_19293);
nor U21620 (N_21620,N_15417,N_19452);
xnor U21621 (N_21621,N_19706,N_18745);
xnor U21622 (N_21622,N_19195,N_15833);
nor U21623 (N_21623,N_17656,N_16924);
nor U21624 (N_21624,N_19793,N_18628);
or U21625 (N_21625,N_15053,N_19132);
nor U21626 (N_21626,N_17582,N_16578);
or U21627 (N_21627,N_15755,N_17872);
xnor U21628 (N_21628,N_15954,N_15988);
nor U21629 (N_21629,N_16495,N_17049);
nor U21630 (N_21630,N_19588,N_18698);
nor U21631 (N_21631,N_16691,N_17686);
and U21632 (N_21632,N_15210,N_18418);
xnor U21633 (N_21633,N_16365,N_18151);
and U21634 (N_21634,N_17564,N_17317);
and U21635 (N_21635,N_18680,N_19906);
or U21636 (N_21636,N_15963,N_17162);
and U21637 (N_21637,N_15962,N_18682);
nand U21638 (N_21638,N_16767,N_15219);
and U21639 (N_21639,N_15781,N_19057);
nor U21640 (N_21640,N_17701,N_17367);
xnor U21641 (N_21641,N_19550,N_19580);
nor U21642 (N_21642,N_19317,N_17914);
xnor U21643 (N_21643,N_19818,N_19181);
xor U21644 (N_21644,N_15182,N_16023);
xnor U21645 (N_21645,N_15245,N_18630);
nor U21646 (N_21646,N_15183,N_18138);
nor U21647 (N_21647,N_15902,N_15746);
nand U21648 (N_21648,N_18155,N_15019);
nor U21649 (N_21649,N_19233,N_18923);
and U21650 (N_21650,N_17695,N_15916);
nor U21651 (N_21651,N_15743,N_18532);
nand U21652 (N_21652,N_18731,N_15654);
or U21653 (N_21653,N_19440,N_15772);
nand U21654 (N_21654,N_19638,N_16584);
nand U21655 (N_21655,N_16403,N_15596);
or U21656 (N_21656,N_18392,N_19654);
and U21657 (N_21657,N_16503,N_16529);
or U21658 (N_21658,N_16614,N_16292);
or U21659 (N_21659,N_15335,N_19069);
nand U21660 (N_21660,N_17576,N_15952);
and U21661 (N_21661,N_15439,N_16134);
and U21662 (N_21662,N_18703,N_15908);
and U21663 (N_21663,N_19357,N_15941);
or U21664 (N_21664,N_15894,N_17634);
and U21665 (N_21665,N_16647,N_15008);
nand U21666 (N_21666,N_18617,N_19802);
and U21667 (N_21667,N_19483,N_15110);
xor U21668 (N_21668,N_18388,N_17667);
nor U21669 (N_21669,N_19081,N_16479);
nor U21670 (N_21670,N_18964,N_15024);
or U21671 (N_21671,N_17017,N_17069);
or U21672 (N_21672,N_15262,N_16068);
nand U21673 (N_21673,N_18265,N_19635);
xnor U21674 (N_21674,N_16338,N_19663);
and U21675 (N_21675,N_16055,N_17761);
xnor U21676 (N_21676,N_15323,N_15408);
or U21677 (N_21677,N_19811,N_18076);
nand U21678 (N_21678,N_15045,N_17304);
and U21679 (N_21679,N_18848,N_16132);
or U21680 (N_21680,N_15579,N_17987);
and U21681 (N_21681,N_18547,N_19656);
and U21682 (N_21682,N_19808,N_16683);
nor U21683 (N_21683,N_15817,N_17554);
or U21684 (N_21684,N_19839,N_16168);
or U21685 (N_21685,N_16653,N_18417);
nand U21686 (N_21686,N_17386,N_17628);
nand U21687 (N_21687,N_18881,N_15123);
or U21688 (N_21688,N_15301,N_18251);
nand U21689 (N_21689,N_19577,N_16409);
or U21690 (N_21690,N_19705,N_15512);
nand U21691 (N_21691,N_18618,N_16203);
and U21692 (N_21692,N_18019,N_16971);
xnor U21693 (N_21693,N_17741,N_18048);
xor U21694 (N_21694,N_19942,N_19681);
nand U21695 (N_21695,N_15786,N_17363);
and U21696 (N_21696,N_15461,N_15154);
and U21697 (N_21697,N_17008,N_17499);
nand U21698 (N_21698,N_16565,N_17655);
xnor U21699 (N_21699,N_18662,N_19395);
xor U21700 (N_21700,N_16776,N_17294);
and U21701 (N_21701,N_18327,N_19371);
nand U21702 (N_21702,N_16101,N_16688);
and U21703 (N_21703,N_18658,N_17851);
or U21704 (N_21704,N_15576,N_15047);
nor U21705 (N_21705,N_16425,N_19570);
and U21706 (N_21706,N_18147,N_18054);
nand U21707 (N_21707,N_17029,N_16083);
and U21708 (N_21708,N_15697,N_19148);
xor U21709 (N_21709,N_19307,N_18979);
or U21710 (N_21710,N_16990,N_15369);
xnor U21711 (N_21711,N_17764,N_16775);
xnor U21712 (N_21712,N_19047,N_16947);
nor U21713 (N_21713,N_15811,N_15261);
xor U21714 (N_21714,N_18498,N_18249);
and U21715 (N_21715,N_15906,N_17860);
nand U21716 (N_21716,N_19533,N_18101);
nand U21717 (N_21717,N_19856,N_19053);
nand U21718 (N_21718,N_15661,N_17884);
or U21719 (N_21719,N_15149,N_19300);
or U21720 (N_21720,N_15996,N_15042);
xnor U21721 (N_21721,N_17684,N_17053);
xnor U21722 (N_21722,N_18755,N_18693);
and U21723 (N_21723,N_15794,N_15305);
nand U21724 (N_21724,N_15627,N_15682);
nand U21725 (N_21725,N_16783,N_15539);
and U21726 (N_21726,N_18666,N_15614);
or U21727 (N_21727,N_16921,N_18412);
and U21728 (N_21728,N_16498,N_18159);
and U21729 (N_21729,N_18463,N_18553);
nor U21730 (N_21730,N_18668,N_18268);
or U21731 (N_21731,N_19095,N_15967);
nor U21732 (N_21732,N_17856,N_16462);
nand U21733 (N_21733,N_18313,N_16770);
and U21734 (N_21734,N_17703,N_19086);
or U21735 (N_21735,N_18157,N_16692);
nand U21736 (N_21736,N_19026,N_18112);
nand U21737 (N_21737,N_16502,N_16358);
xor U21738 (N_21738,N_16594,N_18067);
and U21739 (N_21739,N_19034,N_18030);
xnor U21740 (N_21740,N_19225,N_15214);
nand U21741 (N_21741,N_16445,N_17003);
nor U21742 (N_21742,N_19881,N_18799);
and U21743 (N_21743,N_17399,N_19448);
and U21744 (N_21744,N_18366,N_15551);
nor U21745 (N_21745,N_16061,N_19682);
nor U21746 (N_21746,N_17361,N_16084);
nor U21747 (N_21747,N_17958,N_15452);
or U21748 (N_21748,N_18219,N_17099);
and U21749 (N_21749,N_16255,N_16199);
nor U21750 (N_21750,N_18003,N_15904);
xnor U21751 (N_21751,N_18096,N_17024);
nand U21752 (N_21752,N_18285,N_17046);
and U21753 (N_21753,N_19887,N_16915);
nor U21754 (N_21754,N_15835,N_17217);
and U21755 (N_21755,N_17322,N_19525);
or U21756 (N_21756,N_19689,N_16243);
nor U21757 (N_21757,N_18282,N_19750);
or U21758 (N_21758,N_17857,N_15674);
and U21759 (N_21759,N_19334,N_19245);
nand U21760 (N_21760,N_18530,N_18291);
or U21761 (N_21761,N_15140,N_15292);
nand U21762 (N_21762,N_19961,N_19851);
nor U21763 (N_21763,N_15890,N_19925);
xor U21764 (N_21764,N_15623,N_16597);
nor U21765 (N_21765,N_15886,N_19892);
nand U21766 (N_21766,N_17299,N_17825);
or U21767 (N_21767,N_15834,N_18028);
and U21768 (N_21768,N_18783,N_15364);
nand U21769 (N_21769,N_18719,N_18810);
and U21770 (N_21770,N_19189,N_18896);
nand U21771 (N_21771,N_19401,N_19503);
nand U21772 (N_21772,N_16758,N_19963);
nor U21773 (N_21773,N_15709,N_18005);
xor U21774 (N_21774,N_19241,N_16394);
nand U21775 (N_21775,N_17666,N_19407);
and U21776 (N_21776,N_17473,N_15435);
or U21777 (N_21777,N_16746,N_15048);
and U21778 (N_21778,N_16908,N_17968);
or U21779 (N_21779,N_15350,N_17306);
and U21780 (N_21780,N_17343,N_19876);
or U21781 (N_21781,N_15624,N_16516);
nor U21782 (N_21782,N_19033,N_16254);
xor U21783 (N_21783,N_16044,N_17223);
nand U21784 (N_21784,N_17775,N_19035);
nand U21785 (N_21785,N_17100,N_18971);
nand U21786 (N_21786,N_19331,N_16393);
or U21787 (N_21787,N_17391,N_15552);
or U21788 (N_21788,N_15203,N_19956);
xor U21789 (N_21789,N_19004,N_19510);
xnor U21790 (N_21790,N_16670,N_16877);
nand U21791 (N_21791,N_15950,N_15012);
and U21792 (N_21792,N_19131,N_18377);
nand U21793 (N_21793,N_15863,N_18025);
nand U21794 (N_21794,N_16192,N_16435);
or U21795 (N_21795,N_17624,N_16627);
nand U21796 (N_21796,N_18825,N_15760);
and U21797 (N_21797,N_15796,N_15158);
nor U21798 (N_21798,N_18516,N_17941);
nand U21799 (N_21799,N_15530,N_17555);
xnor U21800 (N_21800,N_15037,N_15460);
nor U21801 (N_21801,N_18776,N_17014);
nor U21802 (N_21802,N_19953,N_17939);
nand U21803 (N_21803,N_18718,N_15383);
and U21804 (N_21804,N_19885,N_16556);
and U21805 (N_21805,N_17848,N_16399);
or U21806 (N_21806,N_19969,N_15563);
xor U21807 (N_21807,N_16305,N_18935);
or U21808 (N_21808,N_15851,N_15533);
and U21809 (N_21809,N_17836,N_19496);
and U21810 (N_21810,N_16368,N_15280);
xnor U21811 (N_21811,N_19773,N_17006);
nor U21812 (N_21812,N_15926,N_19125);
xnor U21813 (N_21813,N_17957,N_16461);
xnor U21814 (N_21814,N_18791,N_19558);
xnor U21815 (N_21815,N_17493,N_19161);
nor U21816 (N_21816,N_17965,N_15373);
and U21817 (N_21817,N_16786,N_15184);
and U21818 (N_21818,N_15406,N_18912);
and U21819 (N_21819,N_15494,N_17736);
xnor U21820 (N_21820,N_17591,N_15507);
nand U21821 (N_21821,N_18303,N_15637);
xnor U21822 (N_21822,N_16709,N_15568);
and U21823 (N_21823,N_15899,N_18633);
xnor U21824 (N_21824,N_19343,N_15438);
nand U21825 (N_21825,N_16227,N_16747);
or U21826 (N_21826,N_17866,N_17388);
or U21827 (N_21827,N_15547,N_15085);
nor U21828 (N_21828,N_16187,N_15744);
nor U21829 (N_21829,N_16808,N_15504);
or U21830 (N_21830,N_17421,N_16247);
nor U21831 (N_21831,N_15252,N_17470);
nand U21832 (N_21832,N_18706,N_15838);
nor U21833 (N_21833,N_18365,N_15523);
nor U21834 (N_21834,N_18195,N_17909);
or U21835 (N_21835,N_16773,N_16402);
or U21836 (N_21836,N_15953,N_16396);
nand U21837 (N_21837,N_16825,N_18004);
or U21838 (N_21838,N_19054,N_15407);
xnor U21839 (N_21839,N_16664,N_19640);
xor U21840 (N_21840,N_15578,N_17042);
nand U21841 (N_21841,N_19098,N_15980);
nor U21842 (N_21842,N_16067,N_18082);
or U21843 (N_21843,N_16548,N_16642);
or U21844 (N_21844,N_16883,N_15052);
or U21845 (N_21845,N_16713,N_19581);
nor U21846 (N_21846,N_19058,N_18511);
or U21847 (N_21847,N_19998,N_18387);
and U21848 (N_21848,N_18914,N_16330);
nand U21849 (N_21849,N_16360,N_16806);
nor U21850 (N_21850,N_18240,N_17840);
and U21851 (N_21851,N_15905,N_17831);
or U21852 (N_21852,N_17558,N_17563);
xnor U21853 (N_21853,N_19276,N_15592);
nand U21854 (N_21854,N_19087,N_19281);
and U21855 (N_21855,N_17195,N_17084);
or U21856 (N_21856,N_17261,N_19061);
or U21857 (N_21857,N_19600,N_18953);
or U21858 (N_21858,N_18021,N_16718);
nand U21859 (N_21859,N_18153,N_17795);
nor U21860 (N_21860,N_17192,N_17377);
and U21861 (N_21861,N_16362,N_17276);
or U21862 (N_21862,N_19470,N_18403);
and U21863 (N_21863,N_16311,N_15293);
nand U21864 (N_21864,N_18785,N_15481);
nand U21865 (N_21865,N_18007,N_17585);
xnor U21866 (N_21866,N_15294,N_18568);
nand U21867 (N_21867,N_17983,N_15711);
nor U21868 (N_21868,N_15826,N_17430);
nand U21869 (N_21869,N_15821,N_18258);
nor U21870 (N_21870,N_18768,N_15455);
xor U21871 (N_21871,N_18137,N_19559);
nand U21872 (N_21872,N_19724,N_17938);
and U21873 (N_21873,N_19698,N_16062);
or U21874 (N_21874,N_16816,N_16568);
nor U21875 (N_21875,N_17431,N_18070);
nand U21876 (N_21876,N_17933,N_16668);
or U21877 (N_21877,N_18334,N_17164);
nor U21878 (N_21878,N_19934,N_15600);
and U21879 (N_21879,N_18013,N_17992);
nor U21880 (N_21880,N_18301,N_15657);
nand U21881 (N_21881,N_19134,N_16370);
and U21882 (N_21882,N_15871,N_19794);
xor U21883 (N_21883,N_16715,N_19905);
and U21884 (N_21884,N_16705,N_16267);
xnor U21885 (N_21885,N_17186,N_16732);
or U21886 (N_21886,N_18758,N_19049);
nor U21887 (N_21887,N_18767,N_16923);
nand U21888 (N_21888,N_19913,N_16880);
or U21889 (N_21889,N_19274,N_17868);
xnor U21890 (N_21890,N_16401,N_18091);
nor U21891 (N_21891,N_16197,N_19572);
xor U21892 (N_21892,N_16481,N_15156);
or U21893 (N_21893,N_16408,N_18861);
or U21894 (N_21894,N_17662,N_19359);
or U21895 (N_21895,N_18426,N_16509);
nand U21896 (N_21896,N_15003,N_19079);
or U21897 (N_21897,N_19221,N_19309);
or U21898 (N_21898,N_15506,N_19652);
and U21899 (N_21899,N_17002,N_16159);
nor U21900 (N_21900,N_16261,N_17985);
xnor U21901 (N_21901,N_17812,N_19847);
or U21902 (N_21902,N_19268,N_16754);
nor U21903 (N_21903,N_17964,N_15565);
xnor U21904 (N_21904,N_19725,N_15602);
and U21905 (N_21905,N_15232,N_16976);
nor U21906 (N_21906,N_19733,N_15322);
nand U21907 (N_21907,N_15348,N_19003);
nor U21908 (N_21908,N_17054,N_16040);
nor U21909 (N_21909,N_16644,N_17578);
or U21910 (N_21910,N_16427,N_15513);
nor U21911 (N_21911,N_17485,N_19678);
and U21912 (N_21912,N_15041,N_15664);
or U21913 (N_21913,N_15362,N_18125);
nand U21914 (N_21914,N_17998,N_16277);
nor U21915 (N_21915,N_16163,N_19449);
nand U21916 (N_21916,N_16052,N_17509);
and U21917 (N_21917,N_15767,N_15464);
nand U21918 (N_21918,N_18501,N_19666);
nand U21919 (N_21919,N_19466,N_15586);
nand U21920 (N_21920,N_17658,N_17454);
and U21921 (N_21921,N_18554,N_16852);
nand U21922 (N_21922,N_17349,N_16395);
xnor U21923 (N_21923,N_15493,N_17638);
or U21924 (N_21924,N_19888,N_16494);
or U21925 (N_21925,N_16621,N_19534);
and U21926 (N_21926,N_17412,N_15001);
xor U21927 (N_21927,N_15098,N_15043);
nor U21928 (N_21928,N_17744,N_18956);
or U21929 (N_21929,N_15145,N_15009);
nor U21930 (N_21930,N_18576,N_17652);
or U21931 (N_21931,N_16636,N_16739);
nor U21932 (N_21932,N_17169,N_16126);
nand U21933 (N_21933,N_17967,N_18830);
nand U21934 (N_21934,N_16316,N_19751);
and U21935 (N_21935,N_19093,N_16803);
or U21936 (N_21936,N_17066,N_17791);
and U21937 (N_21937,N_16538,N_19254);
and U21938 (N_21938,N_17009,N_19843);
nor U21939 (N_21939,N_15017,N_15315);
nand U21940 (N_21940,N_16256,N_19456);
nand U21941 (N_21941,N_17062,N_16266);
or U21942 (N_21942,N_18707,N_17904);
or U21943 (N_21943,N_19736,N_19602);
and U21944 (N_21944,N_18186,N_16349);
nand U21945 (N_21945,N_17898,N_16969);
nor U21946 (N_21946,N_16717,N_17075);
nand U21947 (N_21947,N_15121,N_19816);
nand U21948 (N_21948,N_17520,N_18672);
xor U21949 (N_21949,N_18764,N_19295);
xor U21950 (N_21950,N_18343,N_19836);
or U21951 (N_21951,N_18636,N_15490);
nor U21952 (N_21952,N_15209,N_18237);
xnor U21953 (N_21953,N_18257,N_18150);
nor U21954 (N_21954,N_15146,N_19332);
nand U21955 (N_21955,N_18926,N_16993);
or U21956 (N_21956,N_18761,N_19659);
and U21957 (N_21957,N_19080,N_17809);
or U21958 (N_21958,N_15242,N_18818);
and U21959 (N_21959,N_15569,N_15514);
xnor U21960 (N_21960,N_16869,N_19444);
nand U21961 (N_21961,N_18217,N_16351);
and U21962 (N_21962,N_15853,N_15756);
and U21963 (N_21963,N_15191,N_18837);
nand U21964 (N_21964,N_18751,N_18722);
nor U21965 (N_21965,N_15099,N_19108);
nor U21966 (N_21966,N_16950,N_18535);
nand U21967 (N_21967,N_16359,N_17401);
or U21968 (N_21968,N_17236,N_19006);
nor U21969 (N_21969,N_17129,N_15867);
xnor U21970 (N_21970,N_15440,N_17466);
nor U21971 (N_21971,N_19941,N_18959);
nand U21972 (N_21972,N_15463,N_17782);
xor U21973 (N_21973,N_17713,N_17227);
nand U21974 (N_21974,N_15167,N_18472);
and U21975 (N_21975,N_15717,N_19465);
or U21976 (N_21976,N_19299,N_19042);
xnor U21977 (N_21977,N_15734,N_19711);
xnor U21978 (N_21978,N_15368,N_19957);
xnor U21979 (N_21979,N_19862,N_16714);
and U21980 (N_21980,N_15378,N_17311);
nand U21981 (N_21981,N_15347,N_15701);
nand U21982 (N_21982,N_17127,N_19196);
nand U21983 (N_21983,N_17623,N_18679);
and U21984 (N_21984,N_15577,N_16602);
nand U21985 (N_21985,N_15317,N_15108);
xnor U21986 (N_21986,N_19439,N_17249);
nor U21987 (N_21987,N_18648,N_19805);
nand U21988 (N_21988,N_16980,N_15021);
or U21989 (N_21989,N_15429,N_16079);
xor U21990 (N_21990,N_17381,N_17505);
and U21991 (N_21991,N_15177,N_19273);
nor U21992 (N_21992,N_17404,N_15748);
xor U21993 (N_21993,N_17448,N_15286);
xor U21994 (N_21994,N_17706,N_15284);
nand U21995 (N_21995,N_18777,N_18395);
and U21996 (N_21996,N_19376,N_18110);
or U21997 (N_21997,N_17478,N_18356);
xnor U21998 (N_21998,N_16039,N_19660);
xor U21999 (N_21999,N_17955,N_15574);
nor U22000 (N_22000,N_15331,N_18120);
or U22001 (N_22001,N_17721,N_15635);
and U22002 (N_22002,N_16506,N_15152);
or U22003 (N_22003,N_17881,N_16000);
xor U22004 (N_22004,N_18176,N_16468);
or U22005 (N_22005,N_16944,N_17243);
xnor U22006 (N_22006,N_15855,N_17936);
or U22007 (N_22007,N_19545,N_16645);
or U22008 (N_22008,N_16201,N_18798);
nor U22009 (N_22009,N_19411,N_19322);
nor U22010 (N_22010,N_19966,N_18011);
nor U22011 (N_22011,N_17975,N_19043);
or U22012 (N_22012,N_19869,N_16033);
and U22013 (N_22013,N_17095,N_19048);
and U22014 (N_22014,N_16567,N_18560);
nand U22015 (N_22015,N_19841,N_17797);
and U22016 (N_22016,N_15643,N_16155);
or U22017 (N_22017,N_18752,N_17238);
and U22018 (N_22018,N_15263,N_19130);
and U22019 (N_22019,N_18686,N_17973);
or U22020 (N_22020,N_17659,N_16511);
and U22021 (N_22021,N_18580,N_15216);
nand U22022 (N_22022,N_16422,N_15038);
nor U22023 (N_22023,N_19646,N_15555);
and U22024 (N_22024,N_19927,N_15109);
or U22025 (N_22025,N_17341,N_18397);
nand U22026 (N_22026,N_17422,N_18988);
nand U22027 (N_22027,N_17019,N_15314);
and U22028 (N_22028,N_16046,N_15318);
or U22029 (N_22029,N_17503,N_18381);
and U22030 (N_22030,N_17784,N_18174);
or U22031 (N_22031,N_19457,N_16473);
or U22032 (N_22032,N_19234,N_17508);
xnor U22033 (N_22033,N_16881,N_16383);
nand U22034 (N_22034,N_17225,N_15790);
nand U22035 (N_22035,N_18391,N_17632);
or U22036 (N_22036,N_15720,N_15598);
xnor U22037 (N_22037,N_17206,N_17725);
and U22038 (N_22038,N_16910,N_18816);
or U22039 (N_22039,N_19218,N_16871);
or U22040 (N_22040,N_15553,N_18840);
and U22041 (N_22041,N_19203,N_15319);
nor U22042 (N_22042,N_18793,N_16210);
or U22043 (N_22043,N_15897,N_15651);
xor U22044 (N_22044,N_19044,N_16478);
nand U22045 (N_22045,N_15259,N_16639);
nor U22046 (N_22046,N_16035,N_19178);
or U22047 (N_22047,N_16238,N_19451);
nand U22048 (N_22048,N_16347,N_16784);
xor U22049 (N_22049,N_17111,N_19060);
or U22050 (N_22050,N_16610,N_17182);
or U22051 (N_22051,N_17297,N_15392);
xnor U22052 (N_22052,N_19301,N_19644);
or U22053 (N_22053,N_16239,N_18909);
or U22054 (N_22054,N_15982,N_18650);
and U22055 (N_22055,N_17154,N_17204);
nor U22056 (N_22056,N_17523,N_18239);
and U22057 (N_22057,N_15898,N_16361);
and U22058 (N_22058,N_18763,N_19955);
xor U22059 (N_22059,N_15107,N_18032);
xnor U22060 (N_22060,N_17282,N_16831);
nor U22061 (N_22061,N_19536,N_18901);
nor U22062 (N_22062,N_16224,N_18836);
and U22063 (N_22063,N_18187,N_19240);
and U22064 (N_22064,N_17743,N_15721);
xnor U22065 (N_22065,N_16440,N_18634);
and U22066 (N_22066,N_17275,N_19077);
nor U22067 (N_22067,N_15620,N_15101);
or U22068 (N_22068,N_19564,N_16633);
or U22069 (N_22069,N_16160,N_16334);
and U22070 (N_22070,N_17033,N_15113);
nand U22071 (N_22071,N_16042,N_16870);
nor U22072 (N_22072,N_15653,N_17675);
xor U22073 (N_22073,N_15698,N_16433);
or U22074 (N_22074,N_19091,N_19721);
and U22075 (N_22075,N_19111,N_19213);
nor U22076 (N_22076,N_18246,N_19187);
xor U22077 (N_22077,N_17834,N_15879);
nand U22078 (N_22078,N_15173,N_17671);
nor U22079 (N_22079,N_17822,N_16707);
xnor U22080 (N_22080,N_16959,N_15536);
nor U22081 (N_22081,N_16967,N_15795);
nor U22082 (N_22082,N_15573,N_19506);
nand U22083 (N_22083,N_17946,N_19795);
or U22084 (N_22084,N_18168,N_17173);
nor U22085 (N_22085,N_16455,N_19806);
or U22086 (N_22086,N_18961,N_15699);
or U22087 (N_22087,N_15936,N_15591);
nand U22088 (N_22088,N_17088,N_17180);
nand U22089 (N_22089,N_17302,N_19834);
nand U22090 (N_22090,N_18221,N_18084);
nand U22091 (N_22091,N_19190,N_18442);
or U22092 (N_22092,N_16619,N_19597);
xnor U22093 (N_22093,N_16315,N_16459);
xor U22094 (N_22094,N_16470,N_17906);
xor U22095 (N_22095,N_16145,N_16737);
xnor U22096 (N_22096,N_16577,N_18824);
xnor U22097 (N_22097,N_18963,N_19177);
nand U22098 (N_22098,N_17681,N_16109);
nor U22099 (N_22099,N_17891,N_16874);
nor U22100 (N_22100,N_15492,N_17114);
xnor U22101 (N_22101,N_18927,N_17364);
and U22102 (N_22102,N_18891,N_17141);
nand U22103 (N_22103,N_18323,N_16765);
nor U22104 (N_22104,N_17106,N_18647);
xor U22105 (N_22105,N_15992,N_16405);
nor U22106 (N_22106,N_16148,N_17457);
nand U22107 (N_22107,N_15803,N_18045);
nand U22108 (N_22108,N_19460,N_19650);
or U22109 (N_22109,N_15521,N_16832);
xnor U22110 (N_22110,N_15847,N_18089);
or U22111 (N_22111,N_19089,N_19222);
nand U22112 (N_22112,N_19667,N_17308);
nand U22113 (N_22113,N_17496,N_15129);
and U22114 (N_22114,N_17878,N_19139);
or U22115 (N_22115,N_15964,N_18704);
nor U22116 (N_22116,N_16740,N_19655);
xor U22117 (N_22117,N_17873,N_17474);
nand U22118 (N_22118,N_17337,N_16918);
or U22119 (N_22119,N_17668,N_19115);
or U22120 (N_22120,N_15557,N_15638);
or U22121 (N_22121,N_16312,N_18711);
nand U22122 (N_22122,N_18373,N_19167);
or U22123 (N_22123,N_15715,N_19860);
or U22124 (N_22124,N_18739,N_18344);
and U22125 (N_22125,N_17156,N_17637);
and U22126 (N_22126,N_15727,N_19354);
and U22127 (N_22127,N_18607,N_15587);
xor U22128 (N_22128,N_17678,N_19330);
nor U22129 (N_22129,N_15032,N_17148);
or U22130 (N_22130,N_15581,N_18061);
and U22131 (N_22131,N_16241,N_17265);
xor U22132 (N_22132,N_15436,N_18254);
nor U22133 (N_22133,N_18423,N_16682);
nand U22134 (N_22134,N_15737,N_18638);
and U22135 (N_22135,N_17800,N_17996);
or U22136 (N_22136,N_19804,N_16015);
nor U22137 (N_22137,N_19363,N_15827);
nor U22138 (N_22138,N_16695,N_19789);
nor U22139 (N_22139,N_15780,N_19699);
xnor U22140 (N_22140,N_19135,N_18957);
nand U22141 (N_22141,N_16606,N_15386);
nor U22142 (N_22142,N_17432,N_18488);
nor U22143 (N_22143,N_16788,N_19096);
nor U22144 (N_22144,N_15829,N_17645);
or U22145 (N_22145,N_19830,N_18270);
nor U22146 (N_22146,N_15797,N_19984);
nor U22147 (N_22147,N_15239,N_19386);
and U22148 (N_22148,N_17295,N_15217);
and U22149 (N_22149,N_16546,N_19260);
or U22150 (N_22150,N_17036,N_19772);
xor U22151 (N_22151,N_18917,N_19712);
and U22152 (N_22152,N_16634,N_16559);
nand U22153 (N_22153,N_18801,N_19977);
xor U22154 (N_22154,N_18978,N_16710);
and U22155 (N_22155,N_19066,N_19121);
nand U22156 (N_22156,N_16352,N_19815);
or U22157 (N_22157,N_17193,N_15054);
or U22158 (N_22158,N_17838,N_18531);
xor U22159 (N_22159,N_18590,N_15769);
and U22160 (N_22160,N_17500,N_15939);
or U22161 (N_22161,N_15880,N_16390);
and U22162 (N_22162,N_17929,N_16112);
nor U22163 (N_22163,N_16202,N_16689);
or U22164 (N_22164,N_15747,N_15283);
nand U22165 (N_22165,N_16456,N_19526);
xor U22166 (N_22166,N_19991,N_18973);
and U22167 (N_22167,N_19902,N_19428);
nand U22168 (N_22168,N_19809,N_19546);
xnor U22169 (N_22169,N_15447,N_17864);
or U22170 (N_22170,N_18492,N_15700);
nor U22171 (N_22171,N_15070,N_17573);
or U22172 (N_22172,N_15018,N_19070);
and U22173 (N_22173,N_17022,N_17613);
and U22174 (N_22174,N_19143,N_16960);
xnor U22175 (N_22175,N_17267,N_18276);
nand U22176 (N_22176,N_15759,N_18741);
nand U22177 (N_22177,N_15116,N_19579);
or U22178 (N_22178,N_15934,N_19185);
xnor U22179 (N_22179,N_15590,N_15944);
xor U22180 (N_22180,N_18304,N_15390);
and U22181 (N_22181,N_19764,N_17260);
nand U22182 (N_22182,N_18924,N_15823);
and U22183 (N_22183,N_17183,N_19352);
and U22184 (N_22184,N_17824,N_15562);
nand U22185 (N_22185,N_18736,N_18949);
nor U22186 (N_22186,N_15274,N_15594);
xnor U22187 (N_22187,N_15560,N_16984);
xor U22188 (N_22188,N_19289,N_15307);
nor U22189 (N_22189,N_16523,N_17366);
xor U22190 (N_22190,N_18311,N_19951);
nor U22191 (N_22191,N_16596,N_15387);
and U22192 (N_22192,N_17315,N_17228);
or U22193 (N_22193,N_15940,N_18803);
or U22194 (N_22194,N_16787,N_17385);
and U22195 (N_22195,N_18558,N_18904);
nor U22196 (N_22196,N_16152,N_19515);
or U22197 (N_22197,N_16501,N_15487);
or U22198 (N_22198,N_19198,N_17280);
and U22199 (N_22199,N_15846,N_18325);
nand U22200 (N_22200,N_18597,N_16198);
xor U22201 (N_22201,N_19140,N_15859);
xor U22202 (N_22202,N_18316,N_15393);
xor U22203 (N_22203,N_18878,N_16325);
nor U22204 (N_22204,N_16817,N_16429);
nand U22205 (N_22205,N_15484,N_17598);
nor U22206 (N_22206,N_15852,N_16512);
or U22207 (N_22207,N_15618,N_17903);
xnor U22208 (N_22208,N_19308,N_18601);
xnor U22209 (N_22209,N_18845,N_19105);
nand U22210 (N_22210,N_16889,N_17696);
xnor U22211 (N_22211,N_18451,N_18977);
xor U22212 (N_22212,N_17120,N_17683);
nand U22213 (N_22213,N_16407,N_17731);
and U22214 (N_22214,N_17292,N_17136);
xor U22215 (N_22215,N_17372,N_18505);
or U22216 (N_22216,N_15773,N_17528);
and U22217 (N_22217,N_19429,N_17073);
and U22218 (N_22218,N_18872,N_19893);
and U22219 (N_22219,N_15044,N_17089);
xor U22220 (N_22220,N_16321,N_15266);
xor U22221 (N_22221,N_15931,N_18624);
and U22222 (N_22222,N_16348,N_18592);
or U22223 (N_22223,N_19842,N_16932);
nand U22224 (N_22224,N_17672,N_15425);
nor U22225 (N_22225,N_16590,N_16936);
nand U22226 (N_22226,N_15448,N_18458);
nor U22227 (N_22227,N_16059,N_15485);
nor U22228 (N_22228,N_15302,N_15896);
and U22229 (N_22229,N_15034,N_19224);
nand U22230 (N_22230,N_16121,N_17205);
nand U22231 (N_22231,N_15802,N_17561);
and U22232 (N_22232,N_15131,N_15892);
xor U22233 (N_22233,N_16086,N_17648);
or U22234 (N_22234,N_15342,N_17177);
nor U22235 (N_22235,N_19936,N_19621);
nand U22236 (N_22236,N_19557,N_16036);
nand U22237 (N_22237,N_18455,N_19686);
nand U22238 (N_22238,N_18454,N_16346);
nor U22239 (N_22239,N_17747,N_16452);
nand U22240 (N_22240,N_18253,N_18493);
nand U22241 (N_22241,N_17879,N_18434);
xor U22242 (N_22242,N_19422,N_19319);
and U22243 (N_22243,N_17549,N_19355);
nand U22244 (N_22244,N_16827,N_15785);
or U22245 (N_22245,N_15247,N_16070);
xnor U22246 (N_22246,N_17745,N_19628);
and U22247 (N_22247,N_15910,N_15321);
nand U22248 (N_22248,N_17746,N_18920);
or U22249 (N_22249,N_17536,N_16778);
xor U22250 (N_22250,N_15842,N_15434);
and U22251 (N_22251,N_16458,N_16017);
nor U22252 (N_22252,N_15519,N_17506);
or U22253 (N_22253,N_19133,N_17087);
xor U22254 (N_22254,N_16742,N_18960);
xnor U22255 (N_22255,N_19384,N_15205);
nor U22256 (N_22256,N_15327,N_18974);
and U22257 (N_22257,N_18482,N_16188);
xor U22258 (N_22258,N_18813,N_18600);
and U22259 (N_22259,N_15356,N_19933);
or U22260 (N_22260,N_19812,N_16054);
and U22261 (N_22261,N_19137,N_19014);
xnor U22262 (N_22262,N_15433,N_15716);
or U22263 (N_22263,N_17952,N_17307);
xnor U22264 (N_22264,N_18932,N_16119);
or U22265 (N_22265,N_15665,N_19528);
and U22266 (N_22266,N_18452,N_15479);
nor U22267 (N_22267,N_17124,N_17316);
or U22268 (N_22268,N_15531,N_19461);
or U22269 (N_22269,N_18287,N_19527);
and U22270 (N_22270,N_15300,N_16172);
nor U22271 (N_22271,N_19323,N_18396);
nor U22272 (N_22272,N_17353,N_18085);
or U22273 (N_22273,N_19874,N_18627);
or U22274 (N_22274,N_16138,N_19529);
and U22275 (N_22275,N_15652,N_18133);
and U22276 (N_22276,N_17242,N_18166);
nor U22277 (N_22277,N_17026,N_17209);
and U22278 (N_22278,N_17480,N_18746);
nand U22279 (N_22279,N_18145,N_17760);
and U22280 (N_22280,N_16696,N_17779);
xnor U22281 (N_22281,N_16115,N_17759);
nand U22282 (N_22282,N_17417,N_15669);
nor U22283 (N_22283,N_19846,N_15127);
or U22284 (N_22284,N_16066,N_15731);
nand U22285 (N_22285,N_17463,N_17489);
or U22286 (N_22286,N_18533,N_16283);
xnor U22287 (N_22287,N_17525,N_17515);
or U22288 (N_22288,N_15476,N_16354);
nand U22289 (N_22289,N_19455,N_16716);
or U22290 (N_22290,N_16431,N_15735);
nand U22291 (N_22291,N_17843,N_16853);
nor U22292 (N_22292,N_15212,N_15354);
nand U22293 (N_22293,N_18820,N_19064);
xor U22294 (N_22294,N_17113,N_16147);
and U22295 (N_22295,N_16018,N_19863);
nand U22296 (N_22296,N_16937,N_17532);
nand U22297 (N_22297,N_18090,N_15486);
nor U22298 (N_22298,N_16919,N_17279);
nand U22299 (N_22299,N_18503,N_16665);
xor U22300 (N_22300,N_16628,N_15424);
and U22301 (N_22301,N_18368,N_16830);
xnor U22302 (N_22302,N_15450,N_15544);
nor U22303 (N_22303,N_15421,N_17889);
and U22304 (N_22304,N_18621,N_16049);
nand U22305 (N_22305,N_16679,N_18071);
or U22306 (N_22306,N_18117,N_16020);
nand U22307 (N_22307,N_17698,N_15750);
nand U22308 (N_22308,N_15277,N_19304);
or U22309 (N_22309,N_19514,N_16532);
and U22310 (N_22310,N_17577,N_17011);
and U22311 (N_22311,N_16920,N_19180);
nand U22312 (N_22312,N_15065,N_16569);
nand U22313 (N_22313,N_16591,N_18713);
nand U22314 (N_22314,N_16366,N_16669);
and U22315 (N_22315,N_17626,N_15615);
nand U22316 (N_22316,N_16290,N_16638);
or U22317 (N_22317,N_17411,N_18729);
nor U22318 (N_22318,N_15617,N_18440);
nor U22319 (N_22319,N_15235,N_19018);
nand U22320 (N_22320,N_17961,N_18152);
or U22321 (N_22321,N_17468,N_15502);
xnor U22322 (N_22322,N_19868,N_18727);
xnor U22323 (N_22323,N_19823,N_16781);
and U22324 (N_22324,N_15948,N_17990);
or U22325 (N_22325,N_18606,N_19447);
nor U22326 (N_22326,N_17107,N_15161);
and U22327 (N_22327,N_18880,N_19310);
and U22328 (N_22328,N_17969,N_17565);
and U22329 (N_22329,N_18986,N_19548);
nand U22330 (N_22330,N_15381,N_15732);
xnor U22331 (N_22331,N_19151,N_16214);
xor U22332 (N_22332,N_16794,N_16958);
nand U22333 (N_22333,N_19335,N_19436);
and U22334 (N_22334,N_15222,N_18405);
and U22335 (N_22335,N_18360,N_15451);
or U22336 (N_22336,N_17867,N_19379);
nor U22337 (N_22337,N_17920,N_15789);
and U22338 (N_22338,N_15163,N_19498);
nand U22339 (N_22339,N_19005,N_18573);
nor U22340 (N_22340,N_19405,N_17674);
nand U22341 (N_22341,N_17783,N_16167);
and U22342 (N_22342,N_18033,N_16744);
xor U22343 (N_22343,N_15367,N_19645);
nand U22344 (N_22344,N_16663,N_19083);
or U22345 (N_22345,N_15316,N_18205);
nor U22346 (N_22346,N_18154,N_17922);
nor U22347 (N_22347,N_19507,N_19924);
nor U22348 (N_22348,N_17153,N_17923);
or U22349 (N_22349,N_15022,N_17625);
nand U22350 (N_22350,N_18587,N_15575);
xor U22351 (N_22351,N_18984,N_16507);
and U22352 (N_22352,N_17845,N_18519);
nand U22353 (N_22353,N_16190,N_17239);
nor U22354 (N_22354,N_19296,N_17586);
xnor U22355 (N_22355,N_18983,N_17781);
nand U22356 (N_22356,N_16914,N_15603);
or U22357 (N_22357,N_17201,N_18972);
nor U22358 (N_22358,N_16186,N_17348);
xor U22359 (N_22359,N_17400,N_17318);
nand U22360 (N_22360,N_16727,N_16965);
nand U22361 (N_22361,N_16807,N_15095);
nand U22362 (N_22362,N_17374,N_18372);
or U22363 (N_22363,N_18939,N_19575);
and U22364 (N_22364,N_16884,N_15837);
and U22365 (N_22365,N_15230,N_19462);
nor U22366 (N_22366,N_15612,N_15114);
xor U22367 (N_22367,N_19434,N_17918);
or U22368 (N_22368,N_15118,N_18411);
or U22369 (N_22369,N_16618,N_18502);
nor U22370 (N_22370,N_16092,N_16297);
and U22371 (N_22371,N_17072,N_15503);
or U22372 (N_22372,N_19800,N_15353);
and U22373 (N_22373,N_15611,N_17358);
and U22374 (N_22374,N_16711,N_18473);
xor U22375 (N_22375,N_19651,N_17048);
and U22376 (N_22376,N_19691,N_19899);
xor U22377 (N_22377,N_16216,N_18231);
or U22378 (N_22378,N_19777,N_18382);
and U22379 (N_22379,N_19202,N_17179);
and U22380 (N_22380,N_19521,N_17387);
nor U22381 (N_22381,N_17657,N_19325);
xor U22382 (N_22382,N_15529,N_16270);
nor U22383 (N_22383,N_17079,N_18619);
and U22384 (N_22384,N_19618,N_15922);
or U22385 (N_22385,N_16484,N_18188);
and U22386 (N_22386,N_15500,N_16229);
and U22387 (N_22387,N_15310,N_17244);
nor U22388 (N_22388,N_17877,N_19569);
nand U22389 (N_22389,N_17548,N_19732);
and U22390 (N_22390,N_17266,N_16898);
nor U22391 (N_22391,N_18016,N_19872);
xnor U22392 (N_22392,N_15545,N_18044);
and U22393 (N_22393,N_17692,N_19433);
xor U22394 (N_22394,N_15971,N_16604);
xnor U22395 (N_22395,N_17378,N_19216);
xnor U22396 (N_22396,N_15271,N_19852);
xnor U22397 (N_22397,N_18409,N_18415);
nand U22398 (N_22398,N_16836,N_15714);
and U22399 (N_22399,N_19919,N_16793);
xor U22400 (N_22400,N_18504,N_16557);
nand U22401 (N_22401,N_15752,N_19099);
or U22402 (N_22402,N_15084,N_17590);
xnor U22403 (N_22403,N_15312,N_17928);
nand U22404 (N_22404,N_17711,N_19753);
nand U22405 (N_22405,N_17963,N_17947);
and U22406 (N_22406,N_18779,N_19603);
xnor U22407 (N_22407,N_15030,N_19062);
or U22408 (N_22408,N_18665,N_15275);
xnor U22409 (N_22409,N_19055,N_18135);
nor U22410 (N_22410,N_16953,N_16491);
or U22411 (N_22411,N_19063,N_15719);
nor U22412 (N_22412,N_19792,N_18290);
nor U22413 (N_22413,N_15215,N_18616);
nor U22414 (N_22414,N_15445,N_19910);
or U22415 (N_22415,N_15830,N_19972);
and U22416 (N_22416,N_19409,N_15260);
or U22417 (N_22417,N_16275,N_15622);
and U22418 (N_22418,N_18292,N_19155);
nand U22419 (N_22419,N_18420,N_16181);
and U22420 (N_22420,N_19002,N_16981);
nand U22421 (N_22421,N_18122,N_16090);
xnor U22422 (N_22422,N_15825,N_17045);
nand U22423 (N_22423,N_15628,N_16233);
nand U22424 (N_22424,N_18687,N_15155);
xor U22425 (N_22425,N_19671,N_16558);
and U22426 (N_22426,N_18990,N_19993);
xnor U22427 (N_22427,N_17962,N_18190);
nor U22428 (N_22428,N_18338,N_15074);
nand U22429 (N_22429,N_17375,N_19566);
nor U22430 (N_22430,N_18402,N_19000);
nor U22431 (N_22431,N_18165,N_19123);
or U22432 (N_22432,N_18571,N_15745);
and U22433 (N_22433,N_16535,N_18928);
and U22434 (N_22434,N_15973,N_18340);
nand U22435 (N_22435,N_19278,N_18079);
or U22436 (N_22436,N_17535,N_17137);
or U22437 (N_22437,N_18461,N_15468);
or U22438 (N_22438,N_15990,N_17982);
xnor U22439 (N_22439,N_17609,N_18586);
xnor U22440 (N_22440,N_15807,N_15016);
and U22441 (N_22441,N_15080,N_17972);
xor U22442 (N_22442,N_16666,N_16856);
nor U22443 (N_22443,N_17605,N_18051);
xor U22444 (N_22444,N_19516,N_19136);
or U22445 (N_22445,N_19903,N_19493);
nand U22446 (N_22446,N_16648,N_17853);
nor U22447 (N_22447,N_16289,N_19242);
and U22448 (N_22448,N_19665,N_15974);
xnor U22449 (N_22449,N_18740,N_15005);
xor U22450 (N_22450,N_16392,N_18517);
xor U22451 (N_22451,N_17336,N_16909);
nand U22452 (N_22452,N_15749,N_17254);
xor U22453 (N_22453,N_18644,N_18582);
or U22454 (N_22454,N_17109,N_15220);
or U22455 (N_22455,N_15907,N_19835);
nand U22456 (N_22456,N_19589,N_17654);
xnor U22457 (N_22457,N_17250,N_19124);
or U22458 (N_22458,N_17794,N_16001);
or U22459 (N_22459,N_15983,N_17484);
nor U22460 (N_22460,N_19512,N_15064);
nand U22461 (N_22461,N_17330,N_16274);
and U22462 (N_22462,N_15914,N_19389);
nor U22463 (N_22463,N_16674,N_15289);
and U22464 (N_22464,N_15270,N_15960);
xnor U22465 (N_22465,N_19599,N_16469);
nand U22466 (N_22466,N_15918,N_18539);
nand U22467 (N_22467,N_19050,N_19967);
or U22468 (N_22468,N_16859,N_17566);
xnor U22469 (N_22469,N_15416,N_17726);
or U22470 (N_22470,N_16357,N_16153);
nor U22471 (N_22471,N_17727,N_16041);
nand U22472 (N_22472,N_19358,N_18413);
and U22473 (N_22473,N_18655,N_19092);
or U22474 (N_22474,N_18525,N_17143);
nand U22475 (N_22475,N_18080,N_17767);
xnor U22476 (N_22476,N_17222,N_18664);
xnor U22477 (N_22477,N_17354,N_17172);
nor U22478 (N_22478,N_19675,N_17255);
or U22479 (N_22479,N_19975,N_15872);
nor U22480 (N_22480,N_15680,N_18132);
nor U22481 (N_22481,N_17603,N_16278);
or U22482 (N_22482,N_19929,N_18930);
nand U22483 (N_22483,N_17832,N_19390);
and U22484 (N_22484,N_16745,N_17802);
nor U22485 (N_22485,N_17507,N_16585);
and U22486 (N_22486,N_18057,N_17807);
xnor U22487 (N_22487,N_19741,N_17858);
nand U22488 (N_22488,N_15077,N_19949);
nor U22489 (N_22489,N_15861,N_17810);
and U22490 (N_22490,N_19560,N_17893);
nor U22491 (N_22491,N_19170,N_17151);
and U22492 (N_22492,N_16996,N_18518);
nand U22493 (N_22493,N_19257,N_17321);
nand U22494 (N_22494,N_15142,N_19858);
or U22495 (N_22495,N_15162,N_15518);
or U22496 (N_22496,N_16926,N_17643);
xor U22497 (N_22497,N_18931,N_19909);
and U22498 (N_22498,N_17016,N_19229);
nand U22499 (N_22499,N_19729,N_16438);
xor U22500 (N_22500,N_19431,N_18143);
nand U22501 (N_22501,N_16556,N_15444);
or U22502 (N_22502,N_19348,N_17653);
nor U22503 (N_22503,N_15002,N_18761);
nor U22504 (N_22504,N_15255,N_19893);
nor U22505 (N_22505,N_18348,N_17336);
xnor U22506 (N_22506,N_19171,N_16696);
nor U22507 (N_22507,N_16751,N_18354);
nand U22508 (N_22508,N_15862,N_17598);
xnor U22509 (N_22509,N_15435,N_18725);
and U22510 (N_22510,N_15155,N_16519);
nand U22511 (N_22511,N_18948,N_16266);
and U22512 (N_22512,N_15336,N_15882);
xnor U22513 (N_22513,N_16055,N_18202);
nor U22514 (N_22514,N_19311,N_15592);
xor U22515 (N_22515,N_15214,N_16828);
xor U22516 (N_22516,N_17851,N_15932);
and U22517 (N_22517,N_17751,N_16091);
nand U22518 (N_22518,N_15927,N_19037);
xnor U22519 (N_22519,N_17462,N_18298);
nand U22520 (N_22520,N_16555,N_15743);
nand U22521 (N_22521,N_17766,N_18600);
nor U22522 (N_22522,N_17352,N_17326);
nand U22523 (N_22523,N_17573,N_17385);
xnor U22524 (N_22524,N_19545,N_16089);
nor U22525 (N_22525,N_17214,N_18213);
and U22526 (N_22526,N_18805,N_19250);
xor U22527 (N_22527,N_15977,N_16913);
nand U22528 (N_22528,N_15550,N_15908);
nor U22529 (N_22529,N_15887,N_19958);
and U22530 (N_22530,N_19080,N_16779);
and U22531 (N_22531,N_18889,N_17732);
nor U22532 (N_22532,N_18837,N_15869);
nor U22533 (N_22533,N_15712,N_18010);
nor U22534 (N_22534,N_16995,N_18216);
xor U22535 (N_22535,N_19457,N_19242);
nor U22536 (N_22536,N_19540,N_16308);
xor U22537 (N_22537,N_16252,N_17888);
and U22538 (N_22538,N_19371,N_18536);
nor U22539 (N_22539,N_19838,N_18730);
nand U22540 (N_22540,N_15607,N_18348);
xor U22541 (N_22541,N_18363,N_15387);
nor U22542 (N_22542,N_15208,N_18088);
nand U22543 (N_22543,N_16614,N_16243);
or U22544 (N_22544,N_16561,N_17805);
nand U22545 (N_22545,N_15662,N_19841);
nor U22546 (N_22546,N_15612,N_15131);
or U22547 (N_22547,N_19087,N_17408);
nor U22548 (N_22548,N_15550,N_18272);
xor U22549 (N_22549,N_15378,N_19450);
xor U22550 (N_22550,N_19451,N_15301);
nand U22551 (N_22551,N_17968,N_19889);
nand U22552 (N_22552,N_19616,N_17039);
and U22553 (N_22553,N_17097,N_16048);
and U22554 (N_22554,N_18838,N_16800);
nor U22555 (N_22555,N_18333,N_19779);
nor U22556 (N_22556,N_18510,N_15642);
or U22557 (N_22557,N_19861,N_19357);
or U22558 (N_22558,N_15713,N_18241);
nand U22559 (N_22559,N_15476,N_19533);
nand U22560 (N_22560,N_15223,N_18299);
nor U22561 (N_22561,N_18699,N_19950);
nand U22562 (N_22562,N_17389,N_15958);
or U22563 (N_22563,N_17632,N_16838);
or U22564 (N_22564,N_17930,N_18958);
or U22565 (N_22565,N_17061,N_18668);
and U22566 (N_22566,N_15043,N_17538);
or U22567 (N_22567,N_19952,N_15087);
and U22568 (N_22568,N_17573,N_17193);
or U22569 (N_22569,N_16899,N_15304);
and U22570 (N_22570,N_16316,N_19731);
nand U22571 (N_22571,N_16185,N_19905);
or U22572 (N_22572,N_19566,N_18442);
or U22573 (N_22573,N_17723,N_15205);
or U22574 (N_22574,N_15789,N_18022);
or U22575 (N_22575,N_15587,N_16313);
nand U22576 (N_22576,N_16825,N_15980);
nor U22577 (N_22577,N_16147,N_16790);
nor U22578 (N_22578,N_19569,N_16455);
and U22579 (N_22579,N_16809,N_19189);
xnor U22580 (N_22580,N_19036,N_19462);
or U22581 (N_22581,N_16970,N_15927);
or U22582 (N_22582,N_16346,N_15508);
nand U22583 (N_22583,N_16641,N_19351);
xor U22584 (N_22584,N_19115,N_18118);
and U22585 (N_22585,N_19255,N_19665);
and U22586 (N_22586,N_15657,N_17102);
xor U22587 (N_22587,N_18749,N_19924);
xor U22588 (N_22588,N_15120,N_19195);
nor U22589 (N_22589,N_19257,N_18796);
and U22590 (N_22590,N_15632,N_17599);
nor U22591 (N_22591,N_19851,N_19139);
and U22592 (N_22592,N_15180,N_16275);
or U22593 (N_22593,N_16562,N_17457);
or U22594 (N_22594,N_17387,N_15850);
or U22595 (N_22595,N_16995,N_17938);
xnor U22596 (N_22596,N_15952,N_16399);
or U22597 (N_22597,N_16579,N_16342);
xnor U22598 (N_22598,N_15577,N_17688);
and U22599 (N_22599,N_19743,N_15329);
and U22600 (N_22600,N_19857,N_16525);
nor U22601 (N_22601,N_19360,N_18275);
and U22602 (N_22602,N_16862,N_19522);
or U22603 (N_22603,N_19882,N_15933);
nor U22604 (N_22604,N_16929,N_19556);
nor U22605 (N_22605,N_18832,N_18025);
nand U22606 (N_22606,N_17902,N_16286);
nor U22607 (N_22607,N_15783,N_15073);
nor U22608 (N_22608,N_19124,N_16111);
nor U22609 (N_22609,N_18578,N_15702);
xnor U22610 (N_22610,N_17008,N_18887);
nand U22611 (N_22611,N_19976,N_17116);
or U22612 (N_22612,N_15757,N_19685);
xnor U22613 (N_22613,N_19537,N_17202);
xor U22614 (N_22614,N_15472,N_18511);
and U22615 (N_22615,N_19821,N_18019);
xnor U22616 (N_22616,N_17607,N_17790);
xor U22617 (N_22617,N_16524,N_19383);
or U22618 (N_22618,N_16677,N_19727);
nor U22619 (N_22619,N_19587,N_18547);
nand U22620 (N_22620,N_19838,N_16953);
or U22621 (N_22621,N_18660,N_16029);
xnor U22622 (N_22622,N_18760,N_19704);
nor U22623 (N_22623,N_18122,N_19167);
or U22624 (N_22624,N_15498,N_16630);
xnor U22625 (N_22625,N_15415,N_15496);
nand U22626 (N_22626,N_15651,N_18711);
xor U22627 (N_22627,N_17271,N_19693);
and U22628 (N_22628,N_18411,N_18126);
or U22629 (N_22629,N_18846,N_15639);
and U22630 (N_22630,N_15310,N_15665);
nand U22631 (N_22631,N_19132,N_18273);
nand U22632 (N_22632,N_17255,N_18462);
or U22633 (N_22633,N_15809,N_18741);
or U22634 (N_22634,N_18730,N_19295);
xnor U22635 (N_22635,N_19868,N_16545);
nand U22636 (N_22636,N_15653,N_17513);
xor U22637 (N_22637,N_18458,N_15024);
xor U22638 (N_22638,N_18527,N_16845);
nand U22639 (N_22639,N_15137,N_17528);
or U22640 (N_22640,N_18410,N_16613);
nor U22641 (N_22641,N_15539,N_17362);
xor U22642 (N_22642,N_16908,N_19282);
and U22643 (N_22643,N_15757,N_15943);
and U22644 (N_22644,N_19379,N_18408);
xor U22645 (N_22645,N_17205,N_15995);
xor U22646 (N_22646,N_18246,N_18039);
or U22647 (N_22647,N_18325,N_19196);
xnor U22648 (N_22648,N_19900,N_17459);
xor U22649 (N_22649,N_17973,N_19604);
and U22650 (N_22650,N_19173,N_15407);
nor U22651 (N_22651,N_16121,N_16300);
nand U22652 (N_22652,N_15129,N_16358);
nor U22653 (N_22653,N_16902,N_18607);
nor U22654 (N_22654,N_15964,N_15573);
xnor U22655 (N_22655,N_15625,N_16947);
and U22656 (N_22656,N_19520,N_19832);
or U22657 (N_22657,N_15644,N_19456);
and U22658 (N_22658,N_16373,N_15399);
and U22659 (N_22659,N_17179,N_19061);
nor U22660 (N_22660,N_18969,N_18680);
nand U22661 (N_22661,N_15361,N_16212);
or U22662 (N_22662,N_16974,N_19235);
and U22663 (N_22663,N_18199,N_19860);
nand U22664 (N_22664,N_15680,N_15497);
and U22665 (N_22665,N_16185,N_15095);
nor U22666 (N_22666,N_15896,N_19236);
nor U22667 (N_22667,N_18925,N_18773);
or U22668 (N_22668,N_19985,N_16901);
nor U22669 (N_22669,N_17059,N_15510);
or U22670 (N_22670,N_16223,N_18216);
xor U22671 (N_22671,N_15181,N_18069);
xnor U22672 (N_22672,N_17539,N_18079);
xor U22673 (N_22673,N_18214,N_15481);
nor U22674 (N_22674,N_17397,N_19521);
nor U22675 (N_22675,N_19227,N_19911);
nand U22676 (N_22676,N_16998,N_15029);
xor U22677 (N_22677,N_17310,N_15899);
and U22678 (N_22678,N_18664,N_16472);
or U22679 (N_22679,N_19614,N_17116);
nand U22680 (N_22680,N_19611,N_15616);
or U22681 (N_22681,N_18329,N_16903);
xor U22682 (N_22682,N_17389,N_17018);
xor U22683 (N_22683,N_16755,N_15041);
nand U22684 (N_22684,N_18418,N_17573);
nor U22685 (N_22685,N_16162,N_19039);
nor U22686 (N_22686,N_15698,N_18663);
nand U22687 (N_22687,N_15266,N_17879);
or U22688 (N_22688,N_18658,N_17810);
or U22689 (N_22689,N_17951,N_15336);
nor U22690 (N_22690,N_18269,N_19358);
xor U22691 (N_22691,N_15884,N_16440);
nor U22692 (N_22692,N_15651,N_18462);
or U22693 (N_22693,N_16012,N_19671);
or U22694 (N_22694,N_15075,N_17132);
xnor U22695 (N_22695,N_16151,N_19628);
or U22696 (N_22696,N_15348,N_16486);
xnor U22697 (N_22697,N_19574,N_19315);
and U22698 (N_22698,N_16780,N_19349);
xor U22699 (N_22699,N_16414,N_16203);
xor U22700 (N_22700,N_16800,N_18825);
nand U22701 (N_22701,N_15900,N_16898);
and U22702 (N_22702,N_17352,N_15339);
and U22703 (N_22703,N_17250,N_19187);
or U22704 (N_22704,N_16206,N_17203);
xor U22705 (N_22705,N_18255,N_18953);
nor U22706 (N_22706,N_19811,N_16470);
xnor U22707 (N_22707,N_18596,N_15265);
or U22708 (N_22708,N_19868,N_16941);
nor U22709 (N_22709,N_18616,N_17675);
or U22710 (N_22710,N_16595,N_18258);
nand U22711 (N_22711,N_17350,N_15639);
nor U22712 (N_22712,N_16121,N_19709);
nor U22713 (N_22713,N_15949,N_19284);
nor U22714 (N_22714,N_16262,N_15624);
or U22715 (N_22715,N_17345,N_16041);
and U22716 (N_22716,N_16934,N_16089);
nor U22717 (N_22717,N_15362,N_19859);
or U22718 (N_22718,N_17372,N_16881);
xor U22719 (N_22719,N_16874,N_19724);
or U22720 (N_22720,N_19376,N_16694);
nor U22721 (N_22721,N_16173,N_17360);
xor U22722 (N_22722,N_19147,N_19836);
or U22723 (N_22723,N_15758,N_19766);
or U22724 (N_22724,N_15402,N_15186);
and U22725 (N_22725,N_19410,N_17713);
nand U22726 (N_22726,N_19338,N_16144);
or U22727 (N_22727,N_19981,N_18179);
or U22728 (N_22728,N_17868,N_17418);
xnor U22729 (N_22729,N_17567,N_16796);
nand U22730 (N_22730,N_18628,N_15818);
or U22731 (N_22731,N_16998,N_16560);
nand U22732 (N_22732,N_19448,N_17572);
nor U22733 (N_22733,N_16073,N_17315);
nor U22734 (N_22734,N_19548,N_15254);
nor U22735 (N_22735,N_19062,N_16692);
and U22736 (N_22736,N_16949,N_15127);
or U22737 (N_22737,N_18186,N_19118);
nor U22738 (N_22738,N_19911,N_17941);
xnor U22739 (N_22739,N_18886,N_17378);
xor U22740 (N_22740,N_15229,N_16577);
nand U22741 (N_22741,N_16304,N_18012);
and U22742 (N_22742,N_18015,N_16459);
nand U22743 (N_22743,N_18470,N_19961);
nand U22744 (N_22744,N_19392,N_19293);
xor U22745 (N_22745,N_19718,N_19054);
nor U22746 (N_22746,N_18606,N_18679);
nor U22747 (N_22747,N_18594,N_15633);
and U22748 (N_22748,N_19303,N_15892);
and U22749 (N_22749,N_16982,N_18616);
and U22750 (N_22750,N_18002,N_17030);
and U22751 (N_22751,N_16391,N_18940);
or U22752 (N_22752,N_15015,N_17505);
or U22753 (N_22753,N_17617,N_15001);
nand U22754 (N_22754,N_19792,N_17670);
and U22755 (N_22755,N_19525,N_15063);
or U22756 (N_22756,N_18912,N_19848);
or U22757 (N_22757,N_18441,N_16355);
nor U22758 (N_22758,N_19002,N_16264);
nand U22759 (N_22759,N_19384,N_15295);
nor U22760 (N_22760,N_15791,N_18026);
and U22761 (N_22761,N_15289,N_16229);
xor U22762 (N_22762,N_19695,N_19550);
nor U22763 (N_22763,N_17179,N_19438);
or U22764 (N_22764,N_16058,N_15322);
xnor U22765 (N_22765,N_17096,N_16918);
xor U22766 (N_22766,N_17138,N_19273);
xor U22767 (N_22767,N_19939,N_15957);
nand U22768 (N_22768,N_18021,N_15794);
xor U22769 (N_22769,N_16230,N_18434);
and U22770 (N_22770,N_15279,N_18776);
and U22771 (N_22771,N_15818,N_16897);
or U22772 (N_22772,N_18916,N_19385);
and U22773 (N_22773,N_18897,N_19647);
nor U22774 (N_22774,N_18760,N_19203);
nand U22775 (N_22775,N_16735,N_18292);
nand U22776 (N_22776,N_18920,N_16745);
or U22777 (N_22777,N_19420,N_15481);
xnor U22778 (N_22778,N_15069,N_17945);
or U22779 (N_22779,N_16042,N_19707);
xor U22780 (N_22780,N_15497,N_16798);
nor U22781 (N_22781,N_15414,N_15406);
nor U22782 (N_22782,N_17263,N_16388);
nor U22783 (N_22783,N_19133,N_16814);
xor U22784 (N_22784,N_17929,N_18700);
or U22785 (N_22785,N_15978,N_18414);
and U22786 (N_22786,N_15360,N_17836);
nor U22787 (N_22787,N_18212,N_18695);
and U22788 (N_22788,N_19506,N_18617);
xnor U22789 (N_22789,N_17345,N_16930);
nand U22790 (N_22790,N_18796,N_15725);
xor U22791 (N_22791,N_19944,N_15181);
nand U22792 (N_22792,N_16110,N_17464);
or U22793 (N_22793,N_15111,N_16056);
or U22794 (N_22794,N_18730,N_18667);
xor U22795 (N_22795,N_18349,N_18838);
and U22796 (N_22796,N_19919,N_19248);
xor U22797 (N_22797,N_19138,N_19421);
or U22798 (N_22798,N_16827,N_15047);
nand U22799 (N_22799,N_19431,N_17824);
xnor U22800 (N_22800,N_18331,N_15430);
or U22801 (N_22801,N_15562,N_19686);
nand U22802 (N_22802,N_15975,N_18489);
xor U22803 (N_22803,N_18720,N_18402);
xor U22804 (N_22804,N_15924,N_17429);
nor U22805 (N_22805,N_19875,N_17736);
xor U22806 (N_22806,N_16504,N_18944);
nor U22807 (N_22807,N_19003,N_15640);
and U22808 (N_22808,N_16259,N_15821);
nor U22809 (N_22809,N_18057,N_19429);
xnor U22810 (N_22810,N_16565,N_15393);
and U22811 (N_22811,N_19011,N_19783);
or U22812 (N_22812,N_16931,N_18490);
nand U22813 (N_22813,N_17873,N_15497);
nor U22814 (N_22814,N_17318,N_17881);
nand U22815 (N_22815,N_16810,N_15540);
nand U22816 (N_22816,N_16487,N_17319);
nor U22817 (N_22817,N_15256,N_16741);
and U22818 (N_22818,N_16595,N_19008);
or U22819 (N_22819,N_15452,N_18644);
nor U22820 (N_22820,N_15656,N_15032);
nand U22821 (N_22821,N_15329,N_16660);
or U22822 (N_22822,N_17929,N_16453);
nor U22823 (N_22823,N_19266,N_15877);
xnor U22824 (N_22824,N_16867,N_17911);
nor U22825 (N_22825,N_17233,N_15348);
or U22826 (N_22826,N_17534,N_19993);
or U22827 (N_22827,N_17458,N_16127);
and U22828 (N_22828,N_19745,N_18715);
nand U22829 (N_22829,N_17047,N_19332);
or U22830 (N_22830,N_16830,N_17879);
or U22831 (N_22831,N_17817,N_18799);
nand U22832 (N_22832,N_15420,N_16006);
or U22833 (N_22833,N_17690,N_15057);
or U22834 (N_22834,N_17449,N_15609);
and U22835 (N_22835,N_15082,N_17186);
xor U22836 (N_22836,N_19685,N_15502);
nand U22837 (N_22837,N_16886,N_19319);
nand U22838 (N_22838,N_15719,N_16345);
xnor U22839 (N_22839,N_15841,N_19040);
xnor U22840 (N_22840,N_18918,N_18930);
nor U22841 (N_22841,N_19323,N_15649);
and U22842 (N_22842,N_19256,N_17104);
or U22843 (N_22843,N_16030,N_18975);
xnor U22844 (N_22844,N_18065,N_18080);
nand U22845 (N_22845,N_15995,N_19401);
and U22846 (N_22846,N_16394,N_19399);
xnor U22847 (N_22847,N_19303,N_18757);
or U22848 (N_22848,N_18294,N_18314);
or U22849 (N_22849,N_15637,N_18544);
or U22850 (N_22850,N_15453,N_18359);
nand U22851 (N_22851,N_19028,N_18092);
or U22852 (N_22852,N_16639,N_19774);
and U22853 (N_22853,N_16556,N_19077);
or U22854 (N_22854,N_18326,N_16934);
and U22855 (N_22855,N_16357,N_19491);
nand U22856 (N_22856,N_17300,N_18171);
nand U22857 (N_22857,N_15943,N_19662);
nand U22858 (N_22858,N_19176,N_15903);
nor U22859 (N_22859,N_18316,N_16334);
and U22860 (N_22860,N_16424,N_18306);
nand U22861 (N_22861,N_18766,N_18161);
or U22862 (N_22862,N_18333,N_16181);
and U22863 (N_22863,N_15292,N_19066);
xor U22864 (N_22864,N_15398,N_18597);
and U22865 (N_22865,N_17668,N_18074);
xor U22866 (N_22866,N_15057,N_18847);
nand U22867 (N_22867,N_15752,N_18575);
nand U22868 (N_22868,N_19696,N_15018);
xnor U22869 (N_22869,N_15503,N_16668);
nor U22870 (N_22870,N_19360,N_16049);
xor U22871 (N_22871,N_19765,N_16001);
nand U22872 (N_22872,N_17234,N_15467);
and U22873 (N_22873,N_15569,N_16079);
nand U22874 (N_22874,N_19053,N_16596);
and U22875 (N_22875,N_19984,N_19864);
nand U22876 (N_22876,N_19313,N_19102);
nand U22877 (N_22877,N_15287,N_18251);
nand U22878 (N_22878,N_17403,N_15310);
nor U22879 (N_22879,N_16157,N_17148);
xnor U22880 (N_22880,N_16784,N_17864);
or U22881 (N_22881,N_19249,N_15231);
xor U22882 (N_22882,N_19051,N_16133);
and U22883 (N_22883,N_17356,N_19758);
or U22884 (N_22884,N_16122,N_15720);
or U22885 (N_22885,N_16299,N_17609);
nor U22886 (N_22886,N_16517,N_15333);
or U22887 (N_22887,N_15129,N_15533);
nor U22888 (N_22888,N_17637,N_15958);
xnor U22889 (N_22889,N_17588,N_18825);
or U22890 (N_22890,N_16114,N_19359);
and U22891 (N_22891,N_19536,N_17426);
or U22892 (N_22892,N_17328,N_15514);
or U22893 (N_22893,N_18103,N_15269);
or U22894 (N_22894,N_18249,N_17633);
xor U22895 (N_22895,N_19368,N_18359);
or U22896 (N_22896,N_16555,N_19035);
xor U22897 (N_22897,N_16117,N_15087);
or U22898 (N_22898,N_15225,N_17959);
xnor U22899 (N_22899,N_18272,N_15023);
nand U22900 (N_22900,N_18049,N_17402);
xor U22901 (N_22901,N_19526,N_17504);
nor U22902 (N_22902,N_15217,N_19103);
nor U22903 (N_22903,N_16750,N_16823);
xnor U22904 (N_22904,N_18771,N_15606);
xnor U22905 (N_22905,N_16287,N_19831);
nor U22906 (N_22906,N_15260,N_18562);
nor U22907 (N_22907,N_16848,N_18570);
or U22908 (N_22908,N_17623,N_15515);
xnor U22909 (N_22909,N_18744,N_18802);
and U22910 (N_22910,N_19907,N_19246);
nand U22911 (N_22911,N_18651,N_17202);
xor U22912 (N_22912,N_16616,N_17748);
nor U22913 (N_22913,N_16324,N_15878);
nand U22914 (N_22914,N_17049,N_16468);
nand U22915 (N_22915,N_16906,N_18046);
or U22916 (N_22916,N_17388,N_15629);
and U22917 (N_22917,N_17765,N_17209);
and U22918 (N_22918,N_19104,N_17183);
nand U22919 (N_22919,N_16041,N_16061);
and U22920 (N_22920,N_16649,N_18315);
xor U22921 (N_22921,N_19142,N_18283);
and U22922 (N_22922,N_18033,N_17620);
and U22923 (N_22923,N_19196,N_17807);
nand U22924 (N_22924,N_17780,N_16074);
nand U22925 (N_22925,N_15368,N_19259);
and U22926 (N_22926,N_17541,N_19190);
or U22927 (N_22927,N_18486,N_17232);
and U22928 (N_22928,N_17083,N_15903);
nor U22929 (N_22929,N_16025,N_16728);
or U22930 (N_22930,N_16411,N_19867);
and U22931 (N_22931,N_18243,N_15769);
nand U22932 (N_22932,N_15786,N_19278);
or U22933 (N_22933,N_17028,N_17896);
xnor U22934 (N_22934,N_18076,N_15034);
nand U22935 (N_22935,N_18929,N_18846);
and U22936 (N_22936,N_18379,N_16474);
or U22937 (N_22937,N_18083,N_15503);
xor U22938 (N_22938,N_17876,N_18777);
nor U22939 (N_22939,N_16683,N_16484);
nor U22940 (N_22940,N_16675,N_18437);
or U22941 (N_22941,N_19012,N_16632);
and U22942 (N_22942,N_18088,N_17675);
xnor U22943 (N_22943,N_18019,N_17567);
nand U22944 (N_22944,N_18714,N_16104);
xor U22945 (N_22945,N_18573,N_17940);
xor U22946 (N_22946,N_15808,N_19235);
xor U22947 (N_22947,N_18282,N_16466);
nand U22948 (N_22948,N_18392,N_16195);
or U22949 (N_22949,N_19643,N_17264);
nor U22950 (N_22950,N_15880,N_18377);
and U22951 (N_22951,N_19250,N_15122);
xnor U22952 (N_22952,N_15905,N_16004);
xor U22953 (N_22953,N_18278,N_19712);
nand U22954 (N_22954,N_19700,N_15759);
and U22955 (N_22955,N_19807,N_19274);
nand U22956 (N_22956,N_18447,N_18141);
nand U22957 (N_22957,N_16993,N_17850);
nand U22958 (N_22958,N_17908,N_15364);
nor U22959 (N_22959,N_18349,N_18650);
nand U22960 (N_22960,N_19801,N_17342);
and U22961 (N_22961,N_16162,N_19086);
nand U22962 (N_22962,N_18051,N_19649);
xor U22963 (N_22963,N_17781,N_17114);
nor U22964 (N_22964,N_16021,N_15759);
or U22965 (N_22965,N_19069,N_18919);
nor U22966 (N_22966,N_16359,N_18139);
or U22967 (N_22967,N_16405,N_16606);
and U22968 (N_22968,N_18766,N_19821);
nor U22969 (N_22969,N_19497,N_18256);
and U22970 (N_22970,N_18876,N_18067);
nand U22971 (N_22971,N_17581,N_18047);
nand U22972 (N_22972,N_16638,N_17819);
and U22973 (N_22973,N_15185,N_18218);
nand U22974 (N_22974,N_17266,N_18174);
or U22975 (N_22975,N_17125,N_17527);
nand U22976 (N_22976,N_19557,N_18686);
nor U22977 (N_22977,N_17114,N_16991);
or U22978 (N_22978,N_15565,N_15883);
or U22979 (N_22979,N_17981,N_15928);
and U22980 (N_22980,N_17399,N_15011);
and U22981 (N_22981,N_19441,N_16862);
nand U22982 (N_22982,N_18588,N_18069);
nand U22983 (N_22983,N_17723,N_15746);
and U22984 (N_22984,N_18009,N_15599);
and U22985 (N_22985,N_15253,N_18202);
or U22986 (N_22986,N_19281,N_19132);
or U22987 (N_22987,N_16152,N_19776);
and U22988 (N_22988,N_16572,N_16044);
or U22989 (N_22989,N_18151,N_17904);
or U22990 (N_22990,N_17771,N_17026);
xor U22991 (N_22991,N_15074,N_17704);
and U22992 (N_22992,N_17068,N_18649);
and U22993 (N_22993,N_15272,N_16169);
nor U22994 (N_22994,N_17664,N_17595);
or U22995 (N_22995,N_18213,N_15217);
xor U22996 (N_22996,N_19563,N_17774);
or U22997 (N_22997,N_17766,N_15025);
or U22998 (N_22998,N_18390,N_17777);
or U22999 (N_22999,N_17443,N_18222);
xor U23000 (N_23000,N_17457,N_19632);
nor U23001 (N_23001,N_15754,N_17469);
nor U23002 (N_23002,N_15113,N_18483);
or U23003 (N_23003,N_16913,N_18086);
nand U23004 (N_23004,N_16856,N_15900);
nor U23005 (N_23005,N_17521,N_16758);
and U23006 (N_23006,N_16640,N_15292);
nand U23007 (N_23007,N_19423,N_16167);
xnor U23008 (N_23008,N_17410,N_16786);
nor U23009 (N_23009,N_19226,N_15136);
or U23010 (N_23010,N_17998,N_17850);
nor U23011 (N_23011,N_15920,N_17313);
nand U23012 (N_23012,N_19417,N_16007);
nor U23013 (N_23013,N_15527,N_15051);
xnor U23014 (N_23014,N_17829,N_18762);
nor U23015 (N_23015,N_16192,N_18423);
xnor U23016 (N_23016,N_16589,N_18760);
and U23017 (N_23017,N_17019,N_18555);
and U23018 (N_23018,N_17138,N_19319);
nand U23019 (N_23019,N_15259,N_18761);
or U23020 (N_23020,N_18849,N_19914);
and U23021 (N_23021,N_18818,N_19382);
nand U23022 (N_23022,N_17625,N_16029);
and U23023 (N_23023,N_17221,N_17484);
nand U23024 (N_23024,N_19848,N_16635);
nor U23025 (N_23025,N_16944,N_19982);
nand U23026 (N_23026,N_18653,N_18598);
xnor U23027 (N_23027,N_17883,N_18515);
nand U23028 (N_23028,N_18946,N_16362);
nor U23029 (N_23029,N_15079,N_19995);
and U23030 (N_23030,N_15913,N_15524);
or U23031 (N_23031,N_16372,N_15726);
or U23032 (N_23032,N_19300,N_17728);
or U23033 (N_23033,N_18724,N_15697);
nor U23034 (N_23034,N_15991,N_19650);
nand U23035 (N_23035,N_19414,N_16797);
nand U23036 (N_23036,N_16599,N_19710);
nand U23037 (N_23037,N_17722,N_18526);
and U23038 (N_23038,N_17387,N_17350);
xnor U23039 (N_23039,N_15183,N_17077);
nor U23040 (N_23040,N_15263,N_17185);
and U23041 (N_23041,N_15084,N_15773);
and U23042 (N_23042,N_18128,N_17389);
xor U23043 (N_23043,N_17170,N_16208);
or U23044 (N_23044,N_16963,N_18298);
nor U23045 (N_23045,N_19245,N_15570);
xnor U23046 (N_23046,N_15660,N_17858);
xor U23047 (N_23047,N_15574,N_17133);
xnor U23048 (N_23048,N_18255,N_16192);
or U23049 (N_23049,N_19921,N_17154);
or U23050 (N_23050,N_19958,N_17219);
xor U23051 (N_23051,N_17157,N_17610);
or U23052 (N_23052,N_18789,N_19996);
nand U23053 (N_23053,N_19493,N_16999);
and U23054 (N_23054,N_17527,N_17138);
nand U23055 (N_23055,N_18693,N_16456);
nor U23056 (N_23056,N_18513,N_17872);
xnor U23057 (N_23057,N_15484,N_18322);
xnor U23058 (N_23058,N_18516,N_17091);
nand U23059 (N_23059,N_19778,N_17622);
nand U23060 (N_23060,N_19511,N_15094);
nand U23061 (N_23061,N_17279,N_15008);
nor U23062 (N_23062,N_19207,N_18087);
or U23063 (N_23063,N_17490,N_17069);
nand U23064 (N_23064,N_18052,N_18856);
nand U23065 (N_23065,N_16624,N_19883);
or U23066 (N_23066,N_18314,N_19729);
and U23067 (N_23067,N_15614,N_17494);
or U23068 (N_23068,N_17381,N_15113);
xor U23069 (N_23069,N_18838,N_16471);
and U23070 (N_23070,N_19427,N_15687);
xnor U23071 (N_23071,N_18163,N_17211);
nand U23072 (N_23072,N_17042,N_17041);
xor U23073 (N_23073,N_17256,N_18231);
or U23074 (N_23074,N_15378,N_15929);
nor U23075 (N_23075,N_19015,N_18294);
xor U23076 (N_23076,N_19711,N_16888);
xor U23077 (N_23077,N_18099,N_18058);
nor U23078 (N_23078,N_15685,N_16643);
xnor U23079 (N_23079,N_15895,N_16891);
nor U23080 (N_23080,N_18133,N_17849);
and U23081 (N_23081,N_17730,N_18969);
nor U23082 (N_23082,N_15891,N_19907);
xor U23083 (N_23083,N_16836,N_15810);
or U23084 (N_23084,N_15459,N_18770);
or U23085 (N_23085,N_18322,N_16410);
or U23086 (N_23086,N_16815,N_19848);
xor U23087 (N_23087,N_19823,N_16908);
nand U23088 (N_23088,N_18727,N_15491);
xor U23089 (N_23089,N_16086,N_17973);
xor U23090 (N_23090,N_19234,N_18614);
nor U23091 (N_23091,N_18385,N_19810);
nand U23092 (N_23092,N_16094,N_17323);
nor U23093 (N_23093,N_16374,N_16435);
and U23094 (N_23094,N_17495,N_15192);
nor U23095 (N_23095,N_18644,N_15670);
nor U23096 (N_23096,N_16587,N_16830);
nand U23097 (N_23097,N_16045,N_16065);
or U23098 (N_23098,N_18107,N_16891);
nor U23099 (N_23099,N_15531,N_15121);
or U23100 (N_23100,N_15955,N_18750);
or U23101 (N_23101,N_16664,N_15972);
and U23102 (N_23102,N_18550,N_15752);
or U23103 (N_23103,N_16634,N_19684);
xor U23104 (N_23104,N_19392,N_17735);
xor U23105 (N_23105,N_18353,N_18147);
xor U23106 (N_23106,N_19095,N_16418);
nor U23107 (N_23107,N_16831,N_18516);
nor U23108 (N_23108,N_19665,N_17729);
and U23109 (N_23109,N_15851,N_16173);
xnor U23110 (N_23110,N_15708,N_16158);
and U23111 (N_23111,N_17772,N_17661);
nand U23112 (N_23112,N_19867,N_19160);
or U23113 (N_23113,N_15226,N_15027);
nor U23114 (N_23114,N_17581,N_16302);
nor U23115 (N_23115,N_17224,N_18082);
and U23116 (N_23116,N_18122,N_15657);
xor U23117 (N_23117,N_15089,N_19750);
nor U23118 (N_23118,N_19079,N_18682);
and U23119 (N_23119,N_16429,N_19799);
and U23120 (N_23120,N_19763,N_16339);
nor U23121 (N_23121,N_19354,N_15961);
nand U23122 (N_23122,N_17552,N_18454);
xor U23123 (N_23123,N_16464,N_18361);
and U23124 (N_23124,N_16809,N_19199);
xnor U23125 (N_23125,N_16926,N_16303);
nor U23126 (N_23126,N_16831,N_15706);
or U23127 (N_23127,N_18781,N_18896);
and U23128 (N_23128,N_17596,N_17366);
or U23129 (N_23129,N_16381,N_16577);
nor U23130 (N_23130,N_17815,N_18843);
xor U23131 (N_23131,N_18074,N_15289);
xor U23132 (N_23132,N_17323,N_16719);
xor U23133 (N_23133,N_16078,N_17645);
xor U23134 (N_23134,N_18890,N_15642);
or U23135 (N_23135,N_19642,N_16126);
and U23136 (N_23136,N_18957,N_18063);
and U23137 (N_23137,N_18981,N_19552);
xnor U23138 (N_23138,N_16289,N_15754);
or U23139 (N_23139,N_16519,N_15109);
nor U23140 (N_23140,N_17725,N_17842);
and U23141 (N_23141,N_15870,N_18778);
and U23142 (N_23142,N_19558,N_19427);
nor U23143 (N_23143,N_15924,N_15551);
or U23144 (N_23144,N_17347,N_17282);
xnor U23145 (N_23145,N_19752,N_18324);
nand U23146 (N_23146,N_15915,N_19674);
xor U23147 (N_23147,N_17515,N_16574);
xnor U23148 (N_23148,N_18211,N_17224);
xor U23149 (N_23149,N_15920,N_17056);
and U23150 (N_23150,N_17253,N_19662);
or U23151 (N_23151,N_16824,N_19398);
xor U23152 (N_23152,N_15998,N_16820);
nor U23153 (N_23153,N_15395,N_16568);
or U23154 (N_23154,N_16310,N_18061);
nor U23155 (N_23155,N_15985,N_15186);
nor U23156 (N_23156,N_19860,N_16035);
xnor U23157 (N_23157,N_17176,N_15526);
xor U23158 (N_23158,N_19648,N_16918);
and U23159 (N_23159,N_18907,N_17479);
nor U23160 (N_23160,N_15633,N_18496);
nand U23161 (N_23161,N_17846,N_19365);
nor U23162 (N_23162,N_18200,N_15078);
or U23163 (N_23163,N_17472,N_18371);
nand U23164 (N_23164,N_15120,N_15499);
xor U23165 (N_23165,N_16837,N_15421);
xor U23166 (N_23166,N_18921,N_15939);
nor U23167 (N_23167,N_19892,N_16264);
nor U23168 (N_23168,N_17607,N_16719);
and U23169 (N_23169,N_15697,N_15173);
nand U23170 (N_23170,N_15130,N_17369);
and U23171 (N_23171,N_15475,N_18592);
xnor U23172 (N_23172,N_19361,N_17920);
and U23173 (N_23173,N_18761,N_18629);
xnor U23174 (N_23174,N_18503,N_16177);
and U23175 (N_23175,N_19631,N_15651);
nor U23176 (N_23176,N_18852,N_16976);
xor U23177 (N_23177,N_17142,N_15840);
or U23178 (N_23178,N_15179,N_18345);
xnor U23179 (N_23179,N_16280,N_16165);
or U23180 (N_23180,N_18651,N_17748);
or U23181 (N_23181,N_19239,N_16137);
nor U23182 (N_23182,N_16186,N_18202);
nor U23183 (N_23183,N_19966,N_15827);
or U23184 (N_23184,N_15884,N_15341);
or U23185 (N_23185,N_15566,N_19197);
xor U23186 (N_23186,N_15349,N_19951);
nand U23187 (N_23187,N_18084,N_17673);
nand U23188 (N_23188,N_18457,N_18294);
or U23189 (N_23189,N_17186,N_15323);
xor U23190 (N_23190,N_15290,N_15867);
and U23191 (N_23191,N_16330,N_17968);
or U23192 (N_23192,N_15027,N_17820);
nand U23193 (N_23193,N_18185,N_15753);
nand U23194 (N_23194,N_16593,N_16150);
or U23195 (N_23195,N_19166,N_17128);
and U23196 (N_23196,N_18904,N_16160);
xor U23197 (N_23197,N_16900,N_18758);
and U23198 (N_23198,N_18682,N_19202);
nor U23199 (N_23199,N_15888,N_19327);
or U23200 (N_23200,N_17044,N_17407);
nor U23201 (N_23201,N_16426,N_18253);
and U23202 (N_23202,N_17480,N_17570);
and U23203 (N_23203,N_17616,N_16673);
nor U23204 (N_23204,N_19579,N_19000);
and U23205 (N_23205,N_17642,N_16321);
or U23206 (N_23206,N_18408,N_15983);
nand U23207 (N_23207,N_16966,N_16905);
or U23208 (N_23208,N_19724,N_19969);
and U23209 (N_23209,N_17451,N_16810);
and U23210 (N_23210,N_17548,N_19940);
xnor U23211 (N_23211,N_19760,N_18673);
nor U23212 (N_23212,N_16341,N_16463);
and U23213 (N_23213,N_19358,N_18000);
nand U23214 (N_23214,N_15354,N_17935);
nand U23215 (N_23215,N_15262,N_17310);
nor U23216 (N_23216,N_18698,N_19847);
and U23217 (N_23217,N_19587,N_16714);
xor U23218 (N_23218,N_15990,N_18626);
xnor U23219 (N_23219,N_19757,N_15089);
and U23220 (N_23220,N_19593,N_15524);
nor U23221 (N_23221,N_19924,N_19469);
nand U23222 (N_23222,N_15850,N_15631);
nor U23223 (N_23223,N_18813,N_17934);
or U23224 (N_23224,N_16624,N_18672);
nor U23225 (N_23225,N_19082,N_15028);
nor U23226 (N_23226,N_18385,N_18011);
xor U23227 (N_23227,N_16358,N_18951);
nand U23228 (N_23228,N_17995,N_18050);
xor U23229 (N_23229,N_16279,N_16387);
xor U23230 (N_23230,N_18626,N_19324);
nor U23231 (N_23231,N_15993,N_17733);
nor U23232 (N_23232,N_16062,N_16554);
or U23233 (N_23233,N_18147,N_19918);
xnor U23234 (N_23234,N_18907,N_19786);
xnor U23235 (N_23235,N_16273,N_17535);
xnor U23236 (N_23236,N_15432,N_17645);
and U23237 (N_23237,N_16825,N_17887);
or U23238 (N_23238,N_16488,N_19825);
or U23239 (N_23239,N_16353,N_19059);
nor U23240 (N_23240,N_15247,N_17304);
and U23241 (N_23241,N_16856,N_15568);
xor U23242 (N_23242,N_15037,N_15553);
nand U23243 (N_23243,N_19944,N_18746);
and U23244 (N_23244,N_18991,N_18356);
nand U23245 (N_23245,N_17283,N_19508);
nor U23246 (N_23246,N_15990,N_15791);
nor U23247 (N_23247,N_18822,N_18928);
nor U23248 (N_23248,N_16685,N_17497);
nor U23249 (N_23249,N_18348,N_18568);
nor U23250 (N_23250,N_15952,N_19364);
xor U23251 (N_23251,N_18757,N_16776);
and U23252 (N_23252,N_15912,N_15900);
and U23253 (N_23253,N_15072,N_19767);
and U23254 (N_23254,N_18649,N_19335);
and U23255 (N_23255,N_18325,N_19288);
xnor U23256 (N_23256,N_19765,N_17235);
nand U23257 (N_23257,N_17916,N_19134);
and U23258 (N_23258,N_15556,N_18260);
nor U23259 (N_23259,N_16725,N_17262);
nor U23260 (N_23260,N_19530,N_16090);
nand U23261 (N_23261,N_18092,N_17640);
nand U23262 (N_23262,N_18182,N_18287);
xor U23263 (N_23263,N_19782,N_16024);
xor U23264 (N_23264,N_19066,N_15718);
nand U23265 (N_23265,N_18843,N_17934);
nor U23266 (N_23266,N_15146,N_19645);
xor U23267 (N_23267,N_17967,N_19402);
and U23268 (N_23268,N_17513,N_19294);
or U23269 (N_23269,N_17557,N_15046);
nor U23270 (N_23270,N_15683,N_19468);
and U23271 (N_23271,N_17725,N_15283);
or U23272 (N_23272,N_17071,N_16158);
or U23273 (N_23273,N_19267,N_19138);
nor U23274 (N_23274,N_19948,N_17921);
nor U23275 (N_23275,N_19653,N_19534);
or U23276 (N_23276,N_18141,N_19005);
and U23277 (N_23277,N_17507,N_17607);
nand U23278 (N_23278,N_15367,N_19538);
and U23279 (N_23279,N_15956,N_18332);
xor U23280 (N_23280,N_18457,N_16117);
or U23281 (N_23281,N_15233,N_15978);
or U23282 (N_23282,N_17800,N_19870);
nor U23283 (N_23283,N_15534,N_17685);
nor U23284 (N_23284,N_16606,N_17610);
or U23285 (N_23285,N_16942,N_17315);
or U23286 (N_23286,N_16637,N_16723);
and U23287 (N_23287,N_19409,N_19103);
or U23288 (N_23288,N_18346,N_17257);
nor U23289 (N_23289,N_17566,N_18527);
xor U23290 (N_23290,N_18134,N_19642);
and U23291 (N_23291,N_18011,N_18349);
nand U23292 (N_23292,N_17088,N_19777);
nor U23293 (N_23293,N_18045,N_15438);
nor U23294 (N_23294,N_15396,N_18644);
nand U23295 (N_23295,N_19245,N_18410);
nand U23296 (N_23296,N_18005,N_15180);
xnor U23297 (N_23297,N_17843,N_15082);
nand U23298 (N_23298,N_18003,N_19149);
or U23299 (N_23299,N_15788,N_18291);
nand U23300 (N_23300,N_16633,N_15929);
nand U23301 (N_23301,N_19543,N_18186);
nand U23302 (N_23302,N_16009,N_19199);
xnor U23303 (N_23303,N_17152,N_17293);
or U23304 (N_23304,N_16307,N_19100);
or U23305 (N_23305,N_17012,N_16420);
or U23306 (N_23306,N_15093,N_15245);
and U23307 (N_23307,N_16961,N_17358);
and U23308 (N_23308,N_16977,N_16307);
or U23309 (N_23309,N_17900,N_16263);
or U23310 (N_23310,N_15468,N_19898);
and U23311 (N_23311,N_16032,N_15345);
and U23312 (N_23312,N_17119,N_18288);
nand U23313 (N_23313,N_19054,N_15188);
xor U23314 (N_23314,N_16404,N_16306);
and U23315 (N_23315,N_18297,N_15030);
or U23316 (N_23316,N_17462,N_17267);
or U23317 (N_23317,N_18169,N_16875);
or U23318 (N_23318,N_15585,N_17720);
xor U23319 (N_23319,N_18926,N_17760);
nand U23320 (N_23320,N_15918,N_16673);
or U23321 (N_23321,N_17628,N_15782);
nor U23322 (N_23322,N_15188,N_19756);
and U23323 (N_23323,N_15918,N_18273);
xnor U23324 (N_23324,N_18399,N_16990);
nand U23325 (N_23325,N_17253,N_16292);
nand U23326 (N_23326,N_15567,N_15048);
nor U23327 (N_23327,N_18601,N_18434);
nand U23328 (N_23328,N_16765,N_15893);
nand U23329 (N_23329,N_19691,N_18679);
or U23330 (N_23330,N_16091,N_16736);
nand U23331 (N_23331,N_18923,N_18881);
and U23332 (N_23332,N_17677,N_19026);
or U23333 (N_23333,N_18061,N_17380);
xor U23334 (N_23334,N_16438,N_19888);
xnor U23335 (N_23335,N_17224,N_17945);
and U23336 (N_23336,N_19251,N_16884);
nor U23337 (N_23337,N_17953,N_15770);
xor U23338 (N_23338,N_18563,N_18245);
nor U23339 (N_23339,N_16321,N_17403);
xor U23340 (N_23340,N_17483,N_18724);
or U23341 (N_23341,N_16647,N_18221);
and U23342 (N_23342,N_16263,N_15920);
xnor U23343 (N_23343,N_19838,N_16405);
xor U23344 (N_23344,N_16892,N_17824);
xnor U23345 (N_23345,N_16698,N_16431);
nand U23346 (N_23346,N_17717,N_17543);
or U23347 (N_23347,N_19382,N_15484);
nand U23348 (N_23348,N_16036,N_18809);
and U23349 (N_23349,N_17161,N_15799);
xnor U23350 (N_23350,N_19590,N_15895);
and U23351 (N_23351,N_16033,N_17721);
xor U23352 (N_23352,N_15503,N_17350);
xnor U23353 (N_23353,N_16511,N_18782);
nor U23354 (N_23354,N_15010,N_19107);
nand U23355 (N_23355,N_19231,N_15843);
xnor U23356 (N_23356,N_19508,N_17528);
xnor U23357 (N_23357,N_15163,N_17515);
nand U23358 (N_23358,N_19202,N_15146);
xor U23359 (N_23359,N_16838,N_18044);
or U23360 (N_23360,N_18279,N_15725);
nand U23361 (N_23361,N_18727,N_15867);
or U23362 (N_23362,N_18266,N_16354);
nand U23363 (N_23363,N_16108,N_17617);
or U23364 (N_23364,N_18158,N_17447);
or U23365 (N_23365,N_18003,N_16242);
xnor U23366 (N_23366,N_17505,N_15122);
and U23367 (N_23367,N_19219,N_19218);
nor U23368 (N_23368,N_16324,N_18608);
nor U23369 (N_23369,N_18327,N_18141);
nor U23370 (N_23370,N_19460,N_16768);
or U23371 (N_23371,N_18772,N_16824);
and U23372 (N_23372,N_19720,N_18000);
and U23373 (N_23373,N_15506,N_16428);
xnor U23374 (N_23374,N_18905,N_19469);
nor U23375 (N_23375,N_18412,N_17535);
nor U23376 (N_23376,N_15153,N_18298);
nor U23377 (N_23377,N_19566,N_19845);
nor U23378 (N_23378,N_17594,N_16661);
nor U23379 (N_23379,N_19617,N_17612);
xnor U23380 (N_23380,N_18472,N_17455);
xor U23381 (N_23381,N_19295,N_16914);
or U23382 (N_23382,N_17291,N_16254);
xor U23383 (N_23383,N_18745,N_18401);
nor U23384 (N_23384,N_19046,N_17879);
xnor U23385 (N_23385,N_15023,N_19432);
and U23386 (N_23386,N_15991,N_15807);
or U23387 (N_23387,N_18171,N_16479);
nand U23388 (N_23388,N_19764,N_17202);
xor U23389 (N_23389,N_16220,N_17850);
nor U23390 (N_23390,N_18343,N_17628);
or U23391 (N_23391,N_16283,N_19729);
and U23392 (N_23392,N_16692,N_17965);
or U23393 (N_23393,N_15148,N_17356);
and U23394 (N_23394,N_18229,N_19022);
nand U23395 (N_23395,N_18150,N_19245);
or U23396 (N_23396,N_18077,N_18338);
nor U23397 (N_23397,N_15976,N_16377);
or U23398 (N_23398,N_18300,N_18070);
xnor U23399 (N_23399,N_18113,N_18741);
or U23400 (N_23400,N_19182,N_17968);
nor U23401 (N_23401,N_16851,N_17890);
nand U23402 (N_23402,N_19724,N_16485);
nor U23403 (N_23403,N_17215,N_18316);
nand U23404 (N_23404,N_15186,N_17944);
xnor U23405 (N_23405,N_16537,N_16725);
nand U23406 (N_23406,N_17872,N_18669);
or U23407 (N_23407,N_18206,N_17652);
or U23408 (N_23408,N_16585,N_16525);
nor U23409 (N_23409,N_18080,N_16305);
xnor U23410 (N_23410,N_19840,N_15810);
and U23411 (N_23411,N_16034,N_16114);
nor U23412 (N_23412,N_18347,N_16516);
or U23413 (N_23413,N_17612,N_18791);
or U23414 (N_23414,N_18748,N_16504);
xnor U23415 (N_23415,N_17924,N_15452);
or U23416 (N_23416,N_15698,N_17252);
and U23417 (N_23417,N_18218,N_17561);
nand U23418 (N_23418,N_17688,N_16919);
nor U23419 (N_23419,N_15158,N_18938);
or U23420 (N_23420,N_19175,N_16131);
nand U23421 (N_23421,N_19592,N_17767);
or U23422 (N_23422,N_16516,N_15461);
nor U23423 (N_23423,N_18529,N_15051);
or U23424 (N_23424,N_19719,N_19675);
xor U23425 (N_23425,N_17456,N_18933);
or U23426 (N_23426,N_17100,N_18800);
or U23427 (N_23427,N_16301,N_19994);
nand U23428 (N_23428,N_17095,N_18946);
or U23429 (N_23429,N_15931,N_16425);
xor U23430 (N_23430,N_16476,N_17418);
nand U23431 (N_23431,N_15218,N_17983);
nor U23432 (N_23432,N_16886,N_18250);
and U23433 (N_23433,N_18284,N_16959);
nand U23434 (N_23434,N_19993,N_19639);
nand U23435 (N_23435,N_17567,N_19740);
and U23436 (N_23436,N_16697,N_15364);
and U23437 (N_23437,N_17617,N_18489);
or U23438 (N_23438,N_19013,N_15881);
nor U23439 (N_23439,N_17445,N_16339);
and U23440 (N_23440,N_16470,N_15116);
xor U23441 (N_23441,N_19545,N_17880);
xor U23442 (N_23442,N_19147,N_16251);
xor U23443 (N_23443,N_18248,N_17658);
or U23444 (N_23444,N_17333,N_17929);
nor U23445 (N_23445,N_17025,N_18693);
nand U23446 (N_23446,N_17142,N_17827);
nor U23447 (N_23447,N_18641,N_15712);
or U23448 (N_23448,N_17100,N_16864);
and U23449 (N_23449,N_15821,N_19696);
and U23450 (N_23450,N_15998,N_17073);
nand U23451 (N_23451,N_15861,N_19197);
and U23452 (N_23452,N_18629,N_16103);
xor U23453 (N_23453,N_19940,N_18713);
xor U23454 (N_23454,N_19321,N_17707);
nor U23455 (N_23455,N_16834,N_19873);
nor U23456 (N_23456,N_16567,N_15764);
nand U23457 (N_23457,N_16385,N_17110);
nand U23458 (N_23458,N_19015,N_17196);
nand U23459 (N_23459,N_16078,N_17942);
and U23460 (N_23460,N_16931,N_17171);
or U23461 (N_23461,N_18886,N_15590);
or U23462 (N_23462,N_15970,N_17105);
or U23463 (N_23463,N_15587,N_18714);
nand U23464 (N_23464,N_15168,N_18201);
and U23465 (N_23465,N_17777,N_19740);
xor U23466 (N_23466,N_15855,N_19907);
xnor U23467 (N_23467,N_19052,N_19573);
or U23468 (N_23468,N_18729,N_17635);
nand U23469 (N_23469,N_15650,N_16350);
xnor U23470 (N_23470,N_18930,N_19853);
or U23471 (N_23471,N_16714,N_16030);
nand U23472 (N_23472,N_15232,N_19761);
nand U23473 (N_23473,N_18213,N_15722);
xnor U23474 (N_23474,N_16103,N_16189);
nor U23475 (N_23475,N_15018,N_15781);
or U23476 (N_23476,N_19908,N_16230);
or U23477 (N_23477,N_16544,N_17821);
and U23478 (N_23478,N_17508,N_16742);
xor U23479 (N_23479,N_17603,N_15311);
nand U23480 (N_23480,N_16975,N_19118);
or U23481 (N_23481,N_18221,N_17105);
and U23482 (N_23482,N_18351,N_18864);
and U23483 (N_23483,N_15059,N_19224);
nor U23484 (N_23484,N_17519,N_16141);
or U23485 (N_23485,N_18257,N_17022);
nand U23486 (N_23486,N_19237,N_16176);
and U23487 (N_23487,N_16486,N_19733);
or U23488 (N_23488,N_15521,N_16506);
nand U23489 (N_23489,N_18836,N_17318);
nor U23490 (N_23490,N_19601,N_19906);
nor U23491 (N_23491,N_15501,N_19449);
and U23492 (N_23492,N_16384,N_19041);
xnor U23493 (N_23493,N_19020,N_16012);
nor U23494 (N_23494,N_15634,N_19841);
xor U23495 (N_23495,N_19541,N_15589);
or U23496 (N_23496,N_15813,N_19048);
xnor U23497 (N_23497,N_19692,N_19486);
nor U23498 (N_23498,N_15813,N_18392);
and U23499 (N_23499,N_19625,N_18372);
xor U23500 (N_23500,N_16436,N_18880);
xnor U23501 (N_23501,N_17517,N_15512);
or U23502 (N_23502,N_19558,N_17718);
nand U23503 (N_23503,N_16636,N_18884);
nor U23504 (N_23504,N_15892,N_17547);
xnor U23505 (N_23505,N_16152,N_16498);
nor U23506 (N_23506,N_16127,N_18409);
or U23507 (N_23507,N_15650,N_16118);
and U23508 (N_23508,N_17641,N_18707);
and U23509 (N_23509,N_19526,N_16016);
nand U23510 (N_23510,N_15471,N_19953);
xnor U23511 (N_23511,N_17195,N_18209);
nand U23512 (N_23512,N_19957,N_19336);
or U23513 (N_23513,N_18552,N_16460);
nand U23514 (N_23514,N_17015,N_16812);
and U23515 (N_23515,N_17640,N_18879);
and U23516 (N_23516,N_19835,N_17242);
nor U23517 (N_23517,N_17975,N_18481);
nand U23518 (N_23518,N_19561,N_17694);
xnor U23519 (N_23519,N_18020,N_16656);
nor U23520 (N_23520,N_19873,N_16960);
or U23521 (N_23521,N_16954,N_19732);
or U23522 (N_23522,N_15588,N_18144);
nand U23523 (N_23523,N_19119,N_15253);
and U23524 (N_23524,N_18643,N_15758);
and U23525 (N_23525,N_18317,N_17664);
or U23526 (N_23526,N_18575,N_16762);
and U23527 (N_23527,N_18847,N_16003);
nor U23528 (N_23528,N_16677,N_19950);
nand U23529 (N_23529,N_16939,N_16145);
or U23530 (N_23530,N_19684,N_18207);
nor U23531 (N_23531,N_19766,N_15595);
nand U23532 (N_23532,N_18983,N_15127);
and U23533 (N_23533,N_16097,N_17010);
or U23534 (N_23534,N_19912,N_15700);
nand U23535 (N_23535,N_18799,N_18104);
nor U23536 (N_23536,N_15200,N_16184);
nand U23537 (N_23537,N_17704,N_17828);
nor U23538 (N_23538,N_16766,N_19173);
nor U23539 (N_23539,N_19568,N_19329);
nand U23540 (N_23540,N_19012,N_16129);
xnor U23541 (N_23541,N_19748,N_15204);
and U23542 (N_23542,N_17592,N_17623);
or U23543 (N_23543,N_15381,N_16863);
or U23544 (N_23544,N_15804,N_17059);
xnor U23545 (N_23545,N_17132,N_17504);
nand U23546 (N_23546,N_18627,N_18544);
nand U23547 (N_23547,N_19194,N_15525);
nor U23548 (N_23548,N_18852,N_19005);
nand U23549 (N_23549,N_19824,N_17595);
nor U23550 (N_23550,N_18123,N_16083);
or U23551 (N_23551,N_16820,N_16664);
and U23552 (N_23552,N_16362,N_15042);
and U23553 (N_23553,N_18376,N_17166);
xor U23554 (N_23554,N_15150,N_17877);
nand U23555 (N_23555,N_16480,N_17512);
and U23556 (N_23556,N_18336,N_15127);
nand U23557 (N_23557,N_17780,N_15017);
nor U23558 (N_23558,N_16520,N_18497);
nor U23559 (N_23559,N_17667,N_16326);
and U23560 (N_23560,N_17409,N_16574);
and U23561 (N_23561,N_19376,N_18358);
xnor U23562 (N_23562,N_15454,N_19581);
or U23563 (N_23563,N_19449,N_18353);
and U23564 (N_23564,N_16975,N_17533);
nand U23565 (N_23565,N_19381,N_17235);
nand U23566 (N_23566,N_16499,N_19576);
or U23567 (N_23567,N_17160,N_15912);
or U23568 (N_23568,N_18745,N_15523);
or U23569 (N_23569,N_15432,N_15333);
xor U23570 (N_23570,N_17633,N_18942);
nand U23571 (N_23571,N_19948,N_19943);
and U23572 (N_23572,N_17964,N_19818);
xnor U23573 (N_23573,N_19153,N_16659);
nand U23574 (N_23574,N_19976,N_18224);
xnor U23575 (N_23575,N_17479,N_15280);
nand U23576 (N_23576,N_16166,N_16302);
xnor U23577 (N_23577,N_18825,N_17285);
nor U23578 (N_23578,N_18224,N_18273);
xnor U23579 (N_23579,N_19601,N_17234);
nand U23580 (N_23580,N_15127,N_15996);
nand U23581 (N_23581,N_19074,N_18304);
and U23582 (N_23582,N_19543,N_18323);
or U23583 (N_23583,N_17755,N_18677);
and U23584 (N_23584,N_19639,N_18363);
or U23585 (N_23585,N_19492,N_17231);
and U23586 (N_23586,N_18269,N_16836);
nor U23587 (N_23587,N_19483,N_19372);
and U23588 (N_23588,N_16101,N_18892);
and U23589 (N_23589,N_18734,N_18427);
xnor U23590 (N_23590,N_19509,N_18980);
nor U23591 (N_23591,N_15536,N_19290);
nor U23592 (N_23592,N_19440,N_17735);
xor U23593 (N_23593,N_17602,N_18462);
or U23594 (N_23594,N_18089,N_17969);
nor U23595 (N_23595,N_18072,N_17270);
xnor U23596 (N_23596,N_16838,N_17211);
nand U23597 (N_23597,N_16295,N_18008);
xor U23598 (N_23598,N_18437,N_16518);
nand U23599 (N_23599,N_18608,N_16231);
nor U23600 (N_23600,N_18931,N_18131);
or U23601 (N_23601,N_18226,N_19848);
and U23602 (N_23602,N_19672,N_15694);
and U23603 (N_23603,N_17024,N_17892);
xnor U23604 (N_23604,N_18973,N_19976);
or U23605 (N_23605,N_15278,N_16207);
xnor U23606 (N_23606,N_15615,N_19495);
nor U23607 (N_23607,N_15059,N_15245);
xnor U23608 (N_23608,N_17456,N_18886);
and U23609 (N_23609,N_16203,N_15930);
xor U23610 (N_23610,N_16945,N_16754);
and U23611 (N_23611,N_15764,N_15276);
nand U23612 (N_23612,N_15763,N_15240);
xor U23613 (N_23613,N_16427,N_16306);
and U23614 (N_23614,N_15745,N_15704);
nand U23615 (N_23615,N_18384,N_16172);
or U23616 (N_23616,N_16254,N_17678);
nor U23617 (N_23617,N_18121,N_18667);
xnor U23618 (N_23618,N_16676,N_15211);
or U23619 (N_23619,N_19837,N_18532);
nand U23620 (N_23620,N_16135,N_18023);
xnor U23621 (N_23621,N_15234,N_18626);
xnor U23622 (N_23622,N_16295,N_15507);
and U23623 (N_23623,N_15625,N_15703);
and U23624 (N_23624,N_17500,N_15396);
nor U23625 (N_23625,N_16663,N_18839);
xnor U23626 (N_23626,N_15321,N_18122);
nand U23627 (N_23627,N_17960,N_18852);
and U23628 (N_23628,N_16107,N_16863);
or U23629 (N_23629,N_15403,N_15019);
xnor U23630 (N_23630,N_19320,N_17217);
nand U23631 (N_23631,N_18750,N_19385);
and U23632 (N_23632,N_19317,N_18673);
or U23633 (N_23633,N_17695,N_17786);
and U23634 (N_23634,N_18491,N_17245);
nand U23635 (N_23635,N_18532,N_19239);
or U23636 (N_23636,N_18200,N_17148);
nor U23637 (N_23637,N_16550,N_16258);
nor U23638 (N_23638,N_17427,N_15683);
nor U23639 (N_23639,N_18821,N_19840);
nor U23640 (N_23640,N_17666,N_15870);
nand U23641 (N_23641,N_15249,N_17548);
and U23642 (N_23642,N_15575,N_18732);
and U23643 (N_23643,N_15562,N_16658);
nor U23644 (N_23644,N_17678,N_17632);
and U23645 (N_23645,N_17591,N_16606);
xor U23646 (N_23646,N_17191,N_19982);
xnor U23647 (N_23647,N_17860,N_19706);
and U23648 (N_23648,N_19362,N_15912);
nor U23649 (N_23649,N_18670,N_18802);
xor U23650 (N_23650,N_16058,N_17980);
nor U23651 (N_23651,N_19848,N_16334);
xor U23652 (N_23652,N_16796,N_18546);
nand U23653 (N_23653,N_19409,N_16777);
nand U23654 (N_23654,N_18954,N_17540);
xnor U23655 (N_23655,N_19904,N_16001);
and U23656 (N_23656,N_16905,N_19690);
nor U23657 (N_23657,N_18093,N_16803);
or U23658 (N_23658,N_18187,N_15471);
nor U23659 (N_23659,N_19459,N_17232);
nor U23660 (N_23660,N_16920,N_15270);
or U23661 (N_23661,N_17818,N_19997);
or U23662 (N_23662,N_19132,N_19323);
nor U23663 (N_23663,N_18751,N_15489);
and U23664 (N_23664,N_16848,N_18533);
nor U23665 (N_23665,N_15591,N_15001);
nand U23666 (N_23666,N_18324,N_19863);
nor U23667 (N_23667,N_17905,N_16103);
nand U23668 (N_23668,N_19361,N_16249);
nor U23669 (N_23669,N_17479,N_16905);
or U23670 (N_23670,N_19764,N_17897);
nor U23671 (N_23671,N_19891,N_17858);
nor U23672 (N_23672,N_18230,N_16487);
and U23673 (N_23673,N_17233,N_17600);
and U23674 (N_23674,N_19263,N_15106);
and U23675 (N_23675,N_19554,N_18590);
nor U23676 (N_23676,N_17038,N_16500);
or U23677 (N_23677,N_19756,N_19283);
and U23678 (N_23678,N_16799,N_15693);
or U23679 (N_23679,N_16927,N_19147);
or U23680 (N_23680,N_17605,N_19937);
nor U23681 (N_23681,N_15222,N_18333);
and U23682 (N_23682,N_19518,N_18980);
nand U23683 (N_23683,N_18245,N_15516);
and U23684 (N_23684,N_16655,N_15265);
nor U23685 (N_23685,N_17245,N_16717);
or U23686 (N_23686,N_17889,N_16945);
or U23687 (N_23687,N_17178,N_16093);
nor U23688 (N_23688,N_16988,N_16333);
or U23689 (N_23689,N_18757,N_19051);
nand U23690 (N_23690,N_15130,N_18637);
nand U23691 (N_23691,N_19882,N_19279);
nor U23692 (N_23692,N_18243,N_15842);
or U23693 (N_23693,N_15286,N_16826);
nor U23694 (N_23694,N_15262,N_15706);
nand U23695 (N_23695,N_17619,N_18287);
nand U23696 (N_23696,N_16650,N_18304);
or U23697 (N_23697,N_15464,N_18376);
nand U23698 (N_23698,N_17902,N_18671);
and U23699 (N_23699,N_15742,N_16170);
nand U23700 (N_23700,N_18666,N_15995);
nor U23701 (N_23701,N_17220,N_16565);
nor U23702 (N_23702,N_16370,N_15436);
xnor U23703 (N_23703,N_18954,N_18915);
nor U23704 (N_23704,N_16302,N_18095);
xor U23705 (N_23705,N_15807,N_15102);
and U23706 (N_23706,N_17856,N_19886);
or U23707 (N_23707,N_18846,N_17529);
or U23708 (N_23708,N_19095,N_15140);
nor U23709 (N_23709,N_18221,N_17091);
or U23710 (N_23710,N_19011,N_17292);
xor U23711 (N_23711,N_18397,N_16062);
or U23712 (N_23712,N_17855,N_15899);
xnor U23713 (N_23713,N_17746,N_17780);
and U23714 (N_23714,N_19276,N_15235);
and U23715 (N_23715,N_19490,N_16100);
xnor U23716 (N_23716,N_18814,N_18004);
and U23717 (N_23717,N_17033,N_16121);
nand U23718 (N_23718,N_17884,N_16194);
nand U23719 (N_23719,N_17409,N_15299);
and U23720 (N_23720,N_19194,N_19136);
and U23721 (N_23721,N_18989,N_16207);
xor U23722 (N_23722,N_18559,N_18948);
nor U23723 (N_23723,N_18035,N_19690);
xor U23724 (N_23724,N_15931,N_15689);
xor U23725 (N_23725,N_19255,N_18589);
nand U23726 (N_23726,N_19001,N_17179);
xnor U23727 (N_23727,N_15551,N_18339);
or U23728 (N_23728,N_18447,N_18669);
nand U23729 (N_23729,N_19991,N_15288);
nor U23730 (N_23730,N_16508,N_19694);
and U23731 (N_23731,N_18582,N_18184);
or U23732 (N_23732,N_19990,N_15856);
or U23733 (N_23733,N_15288,N_16896);
xor U23734 (N_23734,N_16677,N_17837);
or U23735 (N_23735,N_17887,N_16121);
nand U23736 (N_23736,N_16560,N_19885);
xnor U23737 (N_23737,N_19042,N_19843);
or U23738 (N_23738,N_17610,N_17615);
nor U23739 (N_23739,N_16776,N_18159);
and U23740 (N_23740,N_15788,N_19797);
and U23741 (N_23741,N_18027,N_17297);
and U23742 (N_23742,N_17277,N_15588);
xnor U23743 (N_23743,N_18338,N_15334);
nor U23744 (N_23744,N_17669,N_17216);
nand U23745 (N_23745,N_19578,N_16614);
xnor U23746 (N_23746,N_19010,N_17929);
xor U23747 (N_23747,N_17355,N_17930);
or U23748 (N_23748,N_19201,N_18193);
xor U23749 (N_23749,N_16121,N_17962);
or U23750 (N_23750,N_16570,N_17337);
or U23751 (N_23751,N_19863,N_18490);
nand U23752 (N_23752,N_15397,N_17087);
and U23753 (N_23753,N_15939,N_16252);
nand U23754 (N_23754,N_15496,N_16685);
and U23755 (N_23755,N_15300,N_19752);
or U23756 (N_23756,N_18777,N_18452);
xor U23757 (N_23757,N_18446,N_16201);
nor U23758 (N_23758,N_17237,N_19410);
or U23759 (N_23759,N_15939,N_17716);
or U23760 (N_23760,N_16180,N_16375);
xor U23761 (N_23761,N_19832,N_19784);
nand U23762 (N_23762,N_16293,N_18548);
nor U23763 (N_23763,N_19087,N_17798);
nand U23764 (N_23764,N_17887,N_18879);
nand U23765 (N_23765,N_15269,N_15705);
and U23766 (N_23766,N_18018,N_17054);
xor U23767 (N_23767,N_17804,N_17404);
nor U23768 (N_23768,N_16624,N_18245);
xor U23769 (N_23769,N_16160,N_19932);
xor U23770 (N_23770,N_15333,N_15162);
nand U23771 (N_23771,N_18218,N_15031);
and U23772 (N_23772,N_17692,N_17417);
nand U23773 (N_23773,N_18098,N_17292);
and U23774 (N_23774,N_18541,N_16170);
or U23775 (N_23775,N_17368,N_16360);
and U23776 (N_23776,N_18847,N_18457);
nand U23777 (N_23777,N_18530,N_19415);
nor U23778 (N_23778,N_19246,N_15746);
nand U23779 (N_23779,N_16907,N_17986);
nand U23780 (N_23780,N_18868,N_16061);
nand U23781 (N_23781,N_19305,N_19450);
or U23782 (N_23782,N_17253,N_17181);
xor U23783 (N_23783,N_16969,N_17704);
nor U23784 (N_23784,N_16808,N_16717);
or U23785 (N_23785,N_15797,N_19743);
nor U23786 (N_23786,N_15977,N_17805);
or U23787 (N_23787,N_15764,N_18760);
or U23788 (N_23788,N_19122,N_18208);
xnor U23789 (N_23789,N_18197,N_17405);
nand U23790 (N_23790,N_19135,N_15602);
nand U23791 (N_23791,N_16272,N_16520);
nor U23792 (N_23792,N_16000,N_18823);
or U23793 (N_23793,N_18294,N_17235);
or U23794 (N_23794,N_17669,N_17471);
and U23795 (N_23795,N_18201,N_18460);
or U23796 (N_23796,N_19269,N_19403);
and U23797 (N_23797,N_18716,N_15558);
xnor U23798 (N_23798,N_17498,N_17432);
or U23799 (N_23799,N_19290,N_15018);
nand U23800 (N_23800,N_16426,N_18820);
nand U23801 (N_23801,N_15664,N_17237);
nand U23802 (N_23802,N_16424,N_18866);
or U23803 (N_23803,N_19125,N_16591);
and U23804 (N_23804,N_18377,N_15804);
and U23805 (N_23805,N_17730,N_19313);
xor U23806 (N_23806,N_15770,N_16076);
or U23807 (N_23807,N_16465,N_15123);
and U23808 (N_23808,N_15926,N_18348);
xnor U23809 (N_23809,N_18732,N_16556);
nor U23810 (N_23810,N_15847,N_15249);
xnor U23811 (N_23811,N_17664,N_19008);
and U23812 (N_23812,N_16052,N_16747);
and U23813 (N_23813,N_15406,N_19184);
nor U23814 (N_23814,N_18056,N_18566);
and U23815 (N_23815,N_17964,N_16762);
and U23816 (N_23816,N_18409,N_15692);
xor U23817 (N_23817,N_19247,N_19012);
or U23818 (N_23818,N_19841,N_16568);
nor U23819 (N_23819,N_19900,N_15098);
nand U23820 (N_23820,N_19331,N_17734);
nand U23821 (N_23821,N_16742,N_18056);
nor U23822 (N_23822,N_16331,N_17773);
or U23823 (N_23823,N_17446,N_15005);
nand U23824 (N_23824,N_17591,N_17904);
and U23825 (N_23825,N_16040,N_17014);
xnor U23826 (N_23826,N_17427,N_19831);
and U23827 (N_23827,N_19312,N_17218);
nor U23828 (N_23828,N_19948,N_18092);
and U23829 (N_23829,N_19040,N_16686);
nor U23830 (N_23830,N_16849,N_19506);
or U23831 (N_23831,N_15341,N_17766);
nor U23832 (N_23832,N_16348,N_19709);
xor U23833 (N_23833,N_19369,N_17257);
or U23834 (N_23834,N_18747,N_16106);
or U23835 (N_23835,N_17761,N_19322);
and U23836 (N_23836,N_19946,N_15683);
and U23837 (N_23837,N_19160,N_18282);
xnor U23838 (N_23838,N_18755,N_16979);
or U23839 (N_23839,N_16293,N_18365);
xor U23840 (N_23840,N_16896,N_18905);
and U23841 (N_23841,N_17042,N_15350);
nand U23842 (N_23842,N_15988,N_18919);
nand U23843 (N_23843,N_16341,N_19589);
or U23844 (N_23844,N_18715,N_19367);
nand U23845 (N_23845,N_15013,N_19857);
xnor U23846 (N_23846,N_16128,N_18706);
or U23847 (N_23847,N_18728,N_15873);
or U23848 (N_23848,N_17154,N_15830);
nor U23849 (N_23849,N_16172,N_16799);
nor U23850 (N_23850,N_19319,N_16460);
or U23851 (N_23851,N_15793,N_19220);
and U23852 (N_23852,N_16927,N_17805);
or U23853 (N_23853,N_18066,N_17465);
nand U23854 (N_23854,N_15272,N_19443);
nand U23855 (N_23855,N_15667,N_16717);
nand U23856 (N_23856,N_15401,N_15974);
nor U23857 (N_23857,N_17386,N_18980);
nor U23858 (N_23858,N_18205,N_16150);
nand U23859 (N_23859,N_19652,N_15868);
nor U23860 (N_23860,N_19461,N_17963);
and U23861 (N_23861,N_16875,N_19251);
or U23862 (N_23862,N_18920,N_15780);
nor U23863 (N_23863,N_19434,N_19865);
and U23864 (N_23864,N_19682,N_16732);
xnor U23865 (N_23865,N_18671,N_16044);
or U23866 (N_23866,N_18518,N_18906);
xor U23867 (N_23867,N_19833,N_15447);
or U23868 (N_23868,N_15265,N_19585);
nor U23869 (N_23869,N_16812,N_16370);
nor U23870 (N_23870,N_17771,N_16499);
or U23871 (N_23871,N_19451,N_15722);
xnor U23872 (N_23872,N_15878,N_16776);
and U23873 (N_23873,N_16192,N_17434);
xor U23874 (N_23874,N_16726,N_16468);
nor U23875 (N_23875,N_18935,N_15802);
and U23876 (N_23876,N_19179,N_17198);
nand U23877 (N_23877,N_18380,N_19130);
or U23878 (N_23878,N_16714,N_15208);
xor U23879 (N_23879,N_17493,N_18007);
xnor U23880 (N_23880,N_18249,N_17541);
xnor U23881 (N_23881,N_16624,N_18073);
or U23882 (N_23882,N_18240,N_18334);
xor U23883 (N_23883,N_16732,N_17572);
xor U23884 (N_23884,N_15421,N_17571);
nor U23885 (N_23885,N_15836,N_16884);
xor U23886 (N_23886,N_18693,N_18518);
or U23887 (N_23887,N_15886,N_16285);
nand U23888 (N_23888,N_17280,N_19949);
or U23889 (N_23889,N_16883,N_19304);
nor U23890 (N_23890,N_19819,N_17211);
nor U23891 (N_23891,N_15582,N_19103);
or U23892 (N_23892,N_16820,N_17397);
xnor U23893 (N_23893,N_16399,N_19884);
nor U23894 (N_23894,N_15302,N_16124);
or U23895 (N_23895,N_19819,N_17081);
xor U23896 (N_23896,N_15588,N_19194);
or U23897 (N_23897,N_19418,N_18115);
xor U23898 (N_23898,N_18961,N_18422);
nor U23899 (N_23899,N_17488,N_16162);
nor U23900 (N_23900,N_19164,N_15719);
nand U23901 (N_23901,N_17452,N_19876);
or U23902 (N_23902,N_18336,N_16693);
nor U23903 (N_23903,N_16811,N_18787);
or U23904 (N_23904,N_15485,N_15856);
nand U23905 (N_23905,N_15370,N_16356);
nand U23906 (N_23906,N_16006,N_18951);
nor U23907 (N_23907,N_18426,N_18969);
nor U23908 (N_23908,N_16711,N_16318);
xor U23909 (N_23909,N_15136,N_18807);
nor U23910 (N_23910,N_17437,N_15555);
nor U23911 (N_23911,N_17573,N_17243);
xor U23912 (N_23912,N_17500,N_19918);
and U23913 (N_23913,N_15604,N_16711);
nor U23914 (N_23914,N_18720,N_18822);
xnor U23915 (N_23915,N_18638,N_19772);
nor U23916 (N_23916,N_17738,N_19384);
nand U23917 (N_23917,N_18313,N_15749);
and U23918 (N_23918,N_17616,N_16061);
and U23919 (N_23919,N_17686,N_17918);
nor U23920 (N_23920,N_17937,N_15532);
nor U23921 (N_23921,N_17879,N_19821);
or U23922 (N_23922,N_16469,N_17444);
nor U23923 (N_23923,N_18230,N_17472);
nand U23924 (N_23924,N_18112,N_15157);
and U23925 (N_23925,N_19408,N_15648);
xor U23926 (N_23926,N_16492,N_16549);
nor U23927 (N_23927,N_18355,N_18599);
and U23928 (N_23928,N_19460,N_16215);
nand U23929 (N_23929,N_18068,N_18477);
xor U23930 (N_23930,N_18247,N_19770);
xnor U23931 (N_23931,N_18935,N_19405);
and U23932 (N_23932,N_17933,N_17112);
or U23933 (N_23933,N_16199,N_15087);
xnor U23934 (N_23934,N_18451,N_17516);
nand U23935 (N_23935,N_18752,N_15967);
or U23936 (N_23936,N_15008,N_18630);
and U23937 (N_23937,N_15834,N_18379);
or U23938 (N_23938,N_17065,N_19588);
xor U23939 (N_23939,N_16924,N_17419);
or U23940 (N_23940,N_19708,N_19264);
and U23941 (N_23941,N_19836,N_17060);
or U23942 (N_23942,N_18886,N_17383);
nor U23943 (N_23943,N_17212,N_15521);
nor U23944 (N_23944,N_19099,N_18608);
or U23945 (N_23945,N_18430,N_18192);
or U23946 (N_23946,N_19214,N_17875);
xnor U23947 (N_23947,N_16727,N_16062);
nand U23948 (N_23948,N_16276,N_18427);
and U23949 (N_23949,N_15759,N_16126);
nor U23950 (N_23950,N_17718,N_16296);
nand U23951 (N_23951,N_16040,N_19911);
and U23952 (N_23952,N_19621,N_18748);
xnor U23953 (N_23953,N_19421,N_16678);
nor U23954 (N_23954,N_15206,N_15454);
xnor U23955 (N_23955,N_15852,N_16853);
or U23956 (N_23956,N_15290,N_15830);
or U23957 (N_23957,N_19901,N_19713);
xnor U23958 (N_23958,N_15733,N_16419);
nand U23959 (N_23959,N_16155,N_19995);
or U23960 (N_23960,N_16668,N_16847);
or U23961 (N_23961,N_15130,N_17462);
nand U23962 (N_23962,N_17676,N_15416);
nor U23963 (N_23963,N_16669,N_18382);
and U23964 (N_23964,N_15610,N_17460);
and U23965 (N_23965,N_18869,N_15891);
or U23966 (N_23966,N_18873,N_17572);
or U23967 (N_23967,N_17514,N_19946);
or U23968 (N_23968,N_16229,N_18501);
or U23969 (N_23969,N_16947,N_16164);
nand U23970 (N_23970,N_18536,N_19928);
and U23971 (N_23971,N_18512,N_19905);
xor U23972 (N_23972,N_19486,N_15430);
nor U23973 (N_23973,N_16756,N_16071);
xnor U23974 (N_23974,N_18773,N_15485);
nand U23975 (N_23975,N_18704,N_17065);
xnor U23976 (N_23976,N_16562,N_18518);
and U23977 (N_23977,N_16122,N_15358);
and U23978 (N_23978,N_19479,N_18417);
nand U23979 (N_23979,N_17940,N_15267);
nand U23980 (N_23980,N_18828,N_16975);
nor U23981 (N_23981,N_19553,N_17204);
nand U23982 (N_23982,N_17378,N_18480);
or U23983 (N_23983,N_15010,N_17061);
nand U23984 (N_23984,N_18578,N_16856);
nor U23985 (N_23985,N_15373,N_16399);
nor U23986 (N_23986,N_16670,N_19901);
or U23987 (N_23987,N_19686,N_16592);
and U23988 (N_23988,N_16482,N_16150);
and U23989 (N_23989,N_19052,N_18459);
xor U23990 (N_23990,N_17989,N_17638);
and U23991 (N_23991,N_16443,N_15502);
and U23992 (N_23992,N_15314,N_18180);
or U23993 (N_23993,N_19796,N_18697);
nor U23994 (N_23994,N_17697,N_17899);
xnor U23995 (N_23995,N_19588,N_17987);
nor U23996 (N_23996,N_18785,N_18480);
and U23997 (N_23997,N_17897,N_17808);
nor U23998 (N_23998,N_19920,N_17182);
or U23999 (N_23999,N_19121,N_15542);
nand U24000 (N_24000,N_17937,N_19550);
nand U24001 (N_24001,N_18572,N_17944);
xnor U24002 (N_24002,N_15735,N_15955);
nand U24003 (N_24003,N_17508,N_19414);
nor U24004 (N_24004,N_18242,N_16537);
nand U24005 (N_24005,N_18531,N_16260);
nor U24006 (N_24006,N_19285,N_16451);
or U24007 (N_24007,N_16962,N_19136);
or U24008 (N_24008,N_15584,N_16653);
xor U24009 (N_24009,N_17506,N_19773);
or U24010 (N_24010,N_15120,N_15449);
nand U24011 (N_24011,N_18213,N_18494);
and U24012 (N_24012,N_19587,N_18427);
nor U24013 (N_24013,N_19217,N_15033);
nand U24014 (N_24014,N_15094,N_17468);
and U24015 (N_24015,N_15930,N_19842);
and U24016 (N_24016,N_16996,N_17534);
nor U24017 (N_24017,N_18174,N_19824);
or U24018 (N_24018,N_19641,N_15460);
or U24019 (N_24019,N_19806,N_19029);
and U24020 (N_24020,N_15715,N_18360);
nand U24021 (N_24021,N_18307,N_18476);
xor U24022 (N_24022,N_18310,N_16739);
or U24023 (N_24023,N_16444,N_19354);
or U24024 (N_24024,N_17776,N_15853);
nand U24025 (N_24025,N_17658,N_16757);
nor U24026 (N_24026,N_15113,N_19574);
xnor U24027 (N_24027,N_18430,N_15470);
nand U24028 (N_24028,N_16118,N_15461);
nand U24029 (N_24029,N_19276,N_16857);
nand U24030 (N_24030,N_18127,N_18176);
xor U24031 (N_24031,N_17266,N_17373);
nand U24032 (N_24032,N_17323,N_17224);
xnor U24033 (N_24033,N_18997,N_16441);
xnor U24034 (N_24034,N_16081,N_19490);
nand U24035 (N_24035,N_19354,N_19897);
or U24036 (N_24036,N_16682,N_16429);
nand U24037 (N_24037,N_17950,N_17656);
nor U24038 (N_24038,N_15365,N_15028);
nand U24039 (N_24039,N_18215,N_15950);
or U24040 (N_24040,N_15259,N_16491);
and U24041 (N_24041,N_19285,N_16465);
nand U24042 (N_24042,N_17061,N_15670);
or U24043 (N_24043,N_18041,N_16502);
xnor U24044 (N_24044,N_17230,N_16374);
nand U24045 (N_24045,N_19513,N_19181);
nand U24046 (N_24046,N_15828,N_18223);
xnor U24047 (N_24047,N_16429,N_19852);
or U24048 (N_24048,N_19618,N_18751);
or U24049 (N_24049,N_16876,N_15525);
and U24050 (N_24050,N_17262,N_17144);
nor U24051 (N_24051,N_17990,N_19643);
and U24052 (N_24052,N_15775,N_18966);
xor U24053 (N_24053,N_19614,N_17896);
and U24054 (N_24054,N_17527,N_18731);
nand U24055 (N_24055,N_18351,N_18611);
nand U24056 (N_24056,N_16675,N_19588);
or U24057 (N_24057,N_15735,N_18135);
and U24058 (N_24058,N_17550,N_15100);
and U24059 (N_24059,N_18483,N_16730);
or U24060 (N_24060,N_19758,N_19895);
or U24061 (N_24061,N_16562,N_17753);
nand U24062 (N_24062,N_18044,N_15070);
nand U24063 (N_24063,N_17755,N_18928);
or U24064 (N_24064,N_18685,N_19484);
nand U24065 (N_24065,N_16341,N_17150);
and U24066 (N_24066,N_19520,N_18495);
or U24067 (N_24067,N_15841,N_17233);
and U24068 (N_24068,N_18299,N_18764);
or U24069 (N_24069,N_19207,N_18652);
and U24070 (N_24070,N_17844,N_17056);
xor U24071 (N_24071,N_17516,N_18845);
xor U24072 (N_24072,N_17304,N_17716);
nand U24073 (N_24073,N_17059,N_19516);
or U24074 (N_24074,N_19193,N_15432);
xnor U24075 (N_24075,N_16914,N_19826);
nand U24076 (N_24076,N_16186,N_15719);
or U24077 (N_24077,N_18100,N_16183);
xnor U24078 (N_24078,N_18335,N_19989);
xnor U24079 (N_24079,N_16744,N_18323);
xnor U24080 (N_24080,N_16402,N_15042);
xnor U24081 (N_24081,N_19342,N_17850);
nand U24082 (N_24082,N_19139,N_16183);
and U24083 (N_24083,N_19962,N_15257);
and U24084 (N_24084,N_19555,N_16773);
nand U24085 (N_24085,N_19739,N_17894);
xnor U24086 (N_24086,N_19682,N_16877);
nand U24087 (N_24087,N_19253,N_16276);
or U24088 (N_24088,N_16051,N_15130);
nor U24089 (N_24089,N_15124,N_15703);
nor U24090 (N_24090,N_19111,N_16027);
xnor U24091 (N_24091,N_16498,N_19857);
or U24092 (N_24092,N_17370,N_16030);
nand U24093 (N_24093,N_19709,N_15473);
xor U24094 (N_24094,N_19100,N_17738);
or U24095 (N_24095,N_18122,N_15694);
or U24096 (N_24096,N_18557,N_15131);
nand U24097 (N_24097,N_19680,N_15247);
or U24098 (N_24098,N_17708,N_16885);
and U24099 (N_24099,N_17164,N_19109);
nor U24100 (N_24100,N_19226,N_19069);
nand U24101 (N_24101,N_19076,N_18308);
xor U24102 (N_24102,N_15151,N_19407);
nor U24103 (N_24103,N_17051,N_16686);
and U24104 (N_24104,N_19580,N_18501);
xnor U24105 (N_24105,N_16492,N_16708);
or U24106 (N_24106,N_15262,N_15000);
nand U24107 (N_24107,N_17229,N_19285);
or U24108 (N_24108,N_19487,N_15198);
xor U24109 (N_24109,N_17050,N_15067);
and U24110 (N_24110,N_17750,N_19776);
xnor U24111 (N_24111,N_15552,N_15646);
nand U24112 (N_24112,N_19065,N_16755);
nor U24113 (N_24113,N_16547,N_15362);
nand U24114 (N_24114,N_15437,N_16655);
and U24115 (N_24115,N_16229,N_16467);
or U24116 (N_24116,N_19289,N_19690);
xnor U24117 (N_24117,N_17549,N_15544);
or U24118 (N_24118,N_16291,N_17686);
xnor U24119 (N_24119,N_15398,N_19994);
nand U24120 (N_24120,N_17624,N_17704);
nand U24121 (N_24121,N_15007,N_15130);
and U24122 (N_24122,N_18506,N_19384);
and U24123 (N_24123,N_17595,N_19731);
nor U24124 (N_24124,N_15718,N_19010);
xnor U24125 (N_24125,N_17588,N_15315);
xor U24126 (N_24126,N_16583,N_19474);
nand U24127 (N_24127,N_16315,N_15320);
nand U24128 (N_24128,N_18005,N_15326);
nor U24129 (N_24129,N_18852,N_15652);
and U24130 (N_24130,N_18895,N_18940);
nand U24131 (N_24131,N_18496,N_16666);
nand U24132 (N_24132,N_17589,N_19282);
or U24133 (N_24133,N_18848,N_17817);
nor U24134 (N_24134,N_16275,N_16819);
nand U24135 (N_24135,N_19584,N_15047);
and U24136 (N_24136,N_19276,N_18193);
and U24137 (N_24137,N_16183,N_17907);
or U24138 (N_24138,N_17663,N_18106);
nand U24139 (N_24139,N_19627,N_15646);
nor U24140 (N_24140,N_15024,N_16206);
or U24141 (N_24141,N_16217,N_19294);
or U24142 (N_24142,N_15186,N_15422);
nand U24143 (N_24143,N_18162,N_15194);
xor U24144 (N_24144,N_17556,N_19578);
or U24145 (N_24145,N_15766,N_15703);
xnor U24146 (N_24146,N_16081,N_16245);
nand U24147 (N_24147,N_17284,N_19181);
nand U24148 (N_24148,N_17764,N_18767);
or U24149 (N_24149,N_16257,N_16245);
and U24150 (N_24150,N_18585,N_17306);
and U24151 (N_24151,N_15841,N_16100);
or U24152 (N_24152,N_18323,N_16969);
nand U24153 (N_24153,N_18188,N_15674);
and U24154 (N_24154,N_16564,N_19442);
xnor U24155 (N_24155,N_16636,N_16274);
or U24156 (N_24156,N_19863,N_15213);
and U24157 (N_24157,N_18773,N_19701);
and U24158 (N_24158,N_19896,N_15588);
nand U24159 (N_24159,N_19975,N_19933);
or U24160 (N_24160,N_15524,N_19074);
and U24161 (N_24161,N_18355,N_19710);
or U24162 (N_24162,N_17981,N_16958);
nand U24163 (N_24163,N_18648,N_17096);
and U24164 (N_24164,N_16985,N_16434);
or U24165 (N_24165,N_16339,N_16925);
and U24166 (N_24166,N_18810,N_19200);
or U24167 (N_24167,N_17629,N_16202);
nand U24168 (N_24168,N_19840,N_16972);
nor U24169 (N_24169,N_19358,N_16307);
nand U24170 (N_24170,N_16175,N_17112);
or U24171 (N_24171,N_15833,N_18845);
and U24172 (N_24172,N_15934,N_18031);
xor U24173 (N_24173,N_15950,N_17726);
xor U24174 (N_24174,N_16087,N_17938);
and U24175 (N_24175,N_19454,N_16041);
xnor U24176 (N_24176,N_16496,N_19093);
or U24177 (N_24177,N_17107,N_19615);
and U24178 (N_24178,N_16391,N_17073);
nor U24179 (N_24179,N_17229,N_17058);
nand U24180 (N_24180,N_15144,N_17322);
nor U24181 (N_24181,N_15029,N_15465);
or U24182 (N_24182,N_15750,N_18603);
nand U24183 (N_24183,N_17022,N_15161);
nand U24184 (N_24184,N_15363,N_16337);
or U24185 (N_24185,N_18825,N_18851);
and U24186 (N_24186,N_15667,N_19131);
or U24187 (N_24187,N_18546,N_16451);
nor U24188 (N_24188,N_16133,N_18907);
or U24189 (N_24189,N_18618,N_19259);
and U24190 (N_24190,N_17998,N_17816);
and U24191 (N_24191,N_16220,N_16215);
nor U24192 (N_24192,N_18887,N_17174);
and U24193 (N_24193,N_15065,N_19551);
xor U24194 (N_24194,N_18180,N_17751);
and U24195 (N_24195,N_15857,N_17780);
nor U24196 (N_24196,N_19852,N_15501);
nand U24197 (N_24197,N_15410,N_19317);
nor U24198 (N_24198,N_18501,N_18035);
xnor U24199 (N_24199,N_18080,N_16020);
xnor U24200 (N_24200,N_19873,N_16105);
nand U24201 (N_24201,N_19154,N_18095);
nor U24202 (N_24202,N_17107,N_15114);
nor U24203 (N_24203,N_15037,N_15407);
nand U24204 (N_24204,N_16151,N_17421);
nor U24205 (N_24205,N_16673,N_18588);
nand U24206 (N_24206,N_17639,N_19530);
and U24207 (N_24207,N_18816,N_15888);
or U24208 (N_24208,N_15479,N_16404);
nand U24209 (N_24209,N_16521,N_17697);
nor U24210 (N_24210,N_18978,N_18164);
and U24211 (N_24211,N_16642,N_15249);
or U24212 (N_24212,N_16107,N_16295);
xor U24213 (N_24213,N_17120,N_19078);
nor U24214 (N_24214,N_15948,N_15894);
nand U24215 (N_24215,N_16009,N_17582);
nor U24216 (N_24216,N_15593,N_19929);
or U24217 (N_24217,N_18024,N_16887);
and U24218 (N_24218,N_16849,N_18627);
and U24219 (N_24219,N_16359,N_15403);
nand U24220 (N_24220,N_19848,N_16471);
or U24221 (N_24221,N_18760,N_19873);
and U24222 (N_24222,N_17198,N_16992);
nor U24223 (N_24223,N_17002,N_18479);
xor U24224 (N_24224,N_19845,N_17185);
xor U24225 (N_24225,N_16456,N_15978);
or U24226 (N_24226,N_16606,N_17553);
or U24227 (N_24227,N_19796,N_18816);
and U24228 (N_24228,N_19326,N_19627);
or U24229 (N_24229,N_16529,N_18069);
and U24230 (N_24230,N_16116,N_18474);
xnor U24231 (N_24231,N_19740,N_18403);
and U24232 (N_24232,N_16698,N_17448);
nor U24233 (N_24233,N_18606,N_16603);
nand U24234 (N_24234,N_19823,N_15995);
nor U24235 (N_24235,N_18318,N_16661);
xnor U24236 (N_24236,N_17219,N_18839);
nor U24237 (N_24237,N_17425,N_18130);
xnor U24238 (N_24238,N_19340,N_16196);
or U24239 (N_24239,N_19843,N_17081);
xor U24240 (N_24240,N_16203,N_17504);
or U24241 (N_24241,N_18478,N_17688);
or U24242 (N_24242,N_16820,N_19395);
and U24243 (N_24243,N_15928,N_15575);
xor U24244 (N_24244,N_15598,N_17211);
and U24245 (N_24245,N_16533,N_15255);
or U24246 (N_24246,N_17715,N_15815);
or U24247 (N_24247,N_16930,N_16836);
nand U24248 (N_24248,N_18673,N_18699);
nand U24249 (N_24249,N_15788,N_15615);
nand U24250 (N_24250,N_16015,N_19052);
xnor U24251 (N_24251,N_16915,N_18852);
xor U24252 (N_24252,N_15099,N_18262);
or U24253 (N_24253,N_15181,N_16144);
nor U24254 (N_24254,N_19788,N_18276);
and U24255 (N_24255,N_15756,N_19638);
xnor U24256 (N_24256,N_17117,N_18984);
nor U24257 (N_24257,N_16092,N_18874);
and U24258 (N_24258,N_18737,N_15228);
nand U24259 (N_24259,N_19073,N_19856);
xnor U24260 (N_24260,N_15456,N_17999);
nand U24261 (N_24261,N_17739,N_16083);
or U24262 (N_24262,N_15447,N_17686);
xor U24263 (N_24263,N_18621,N_18161);
nor U24264 (N_24264,N_17733,N_18454);
nor U24265 (N_24265,N_15090,N_16021);
nand U24266 (N_24266,N_17569,N_17949);
nand U24267 (N_24267,N_19749,N_18237);
xnor U24268 (N_24268,N_17675,N_19420);
nor U24269 (N_24269,N_19279,N_16483);
or U24270 (N_24270,N_15080,N_17847);
and U24271 (N_24271,N_17845,N_15588);
nand U24272 (N_24272,N_16486,N_19356);
nand U24273 (N_24273,N_18013,N_19945);
nand U24274 (N_24274,N_17511,N_19260);
nand U24275 (N_24275,N_16699,N_17705);
or U24276 (N_24276,N_16261,N_15409);
xnor U24277 (N_24277,N_19639,N_16725);
xnor U24278 (N_24278,N_17435,N_17204);
xor U24279 (N_24279,N_19042,N_17581);
nor U24280 (N_24280,N_17683,N_16574);
or U24281 (N_24281,N_19649,N_18713);
xor U24282 (N_24282,N_18889,N_18460);
nor U24283 (N_24283,N_16003,N_19583);
nand U24284 (N_24284,N_19821,N_19022);
xor U24285 (N_24285,N_15920,N_15120);
nor U24286 (N_24286,N_16508,N_15823);
nor U24287 (N_24287,N_17971,N_19301);
nand U24288 (N_24288,N_18753,N_19829);
and U24289 (N_24289,N_16609,N_16979);
xor U24290 (N_24290,N_18112,N_19194);
xnor U24291 (N_24291,N_16176,N_19931);
xnor U24292 (N_24292,N_16751,N_16688);
and U24293 (N_24293,N_18201,N_15806);
and U24294 (N_24294,N_18800,N_18725);
or U24295 (N_24295,N_19817,N_15506);
xor U24296 (N_24296,N_15542,N_16321);
nor U24297 (N_24297,N_17415,N_19331);
xnor U24298 (N_24298,N_15111,N_17465);
nor U24299 (N_24299,N_19598,N_19182);
and U24300 (N_24300,N_15028,N_15419);
and U24301 (N_24301,N_17453,N_15316);
or U24302 (N_24302,N_15007,N_15433);
nor U24303 (N_24303,N_15311,N_18268);
or U24304 (N_24304,N_19912,N_17936);
or U24305 (N_24305,N_16214,N_17947);
xnor U24306 (N_24306,N_18688,N_16977);
and U24307 (N_24307,N_18133,N_19958);
nor U24308 (N_24308,N_16460,N_18193);
xnor U24309 (N_24309,N_19077,N_16708);
nor U24310 (N_24310,N_16757,N_19340);
or U24311 (N_24311,N_16806,N_18644);
or U24312 (N_24312,N_18343,N_16876);
nand U24313 (N_24313,N_16178,N_15475);
nand U24314 (N_24314,N_15837,N_17819);
nor U24315 (N_24315,N_16198,N_17231);
nor U24316 (N_24316,N_17269,N_19759);
or U24317 (N_24317,N_19858,N_15437);
nor U24318 (N_24318,N_19872,N_19643);
nand U24319 (N_24319,N_15872,N_19924);
xor U24320 (N_24320,N_17398,N_19577);
nor U24321 (N_24321,N_16413,N_17999);
nand U24322 (N_24322,N_19052,N_15110);
nand U24323 (N_24323,N_16846,N_18325);
and U24324 (N_24324,N_15803,N_18473);
and U24325 (N_24325,N_18396,N_18289);
xor U24326 (N_24326,N_19049,N_15553);
and U24327 (N_24327,N_15972,N_18757);
xor U24328 (N_24328,N_19649,N_17435);
nor U24329 (N_24329,N_18917,N_18804);
xor U24330 (N_24330,N_17574,N_15587);
or U24331 (N_24331,N_16262,N_17365);
nor U24332 (N_24332,N_18824,N_17360);
or U24333 (N_24333,N_15094,N_15712);
nor U24334 (N_24334,N_15916,N_16854);
nand U24335 (N_24335,N_15707,N_17754);
and U24336 (N_24336,N_15886,N_15246);
and U24337 (N_24337,N_16427,N_18792);
xor U24338 (N_24338,N_16810,N_18300);
nor U24339 (N_24339,N_16155,N_16557);
xor U24340 (N_24340,N_19942,N_16809);
and U24341 (N_24341,N_15981,N_18498);
nand U24342 (N_24342,N_17911,N_16581);
nor U24343 (N_24343,N_17138,N_16293);
nor U24344 (N_24344,N_18618,N_15443);
or U24345 (N_24345,N_18011,N_15447);
and U24346 (N_24346,N_18847,N_17240);
xor U24347 (N_24347,N_17556,N_19183);
and U24348 (N_24348,N_16121,N_19515);
nor U24349 (N_24349,N_15934,N_18862);
xor U24350 (N_24350,N_18158,N_18935);
nor U24351 (N_24351,N_18086,N_17480);
and U24352 (N_24352,N_16676,N_19467);
or U24353 (N_24353,N_18368,N_18204);
and U24354 (N_24354,N_19052,N_16256);
xor U24355 (N_24355,N_17413,N_15404);
xor U24356 (N_24356,N_19909,N_16081);
nand U24357 (N_24357,N_17172,N_18697);
nand U24358 (N_24358,N_15660,N_19597);
and U24359 (N_24359,N_15559,N_15081);
and U24360 (N_24360,N_15776,N_17475);
and U24361 (N_24361,N_18490,N_19964);
and U24362 (N_24362,N_15320,N_17925);
xor U24363 (N_24363,N_15464,N_19462);
nand U24364 (N_24364,N_15673,N_18803);
nand U24365 (N_24365,N_15976,N_18485);
and U24366 (N_24366,N_16640,N_19427);
or U24367 (N_24367,N_15826,N_19519);
xnor U24368 (N_24368,N_16968,N_18845);
nor U24369 (N_24369,N_16328,N_16206);
nand U24370 (N_24370,N_15930,N_19276);
nor U24371 (N_24371,N_19565,N_17210);
nand U24372 (N_24372,N_18638,N_18857);
nor U24373 (N_24373,N_19551,N_19950);
xnor U24374 (N_24374,N_17687,N_15019);
xor U24375 (N_24375,N_15648,N_17890);
nand U24376 (N_24376,N_15589,N_17773);
xor U24377 (N_24377,N_19013,N_15065);
or U24378 (N_24378,N_18314,N_18847);
and U24379 (N_24379,N_19829,N_18749);
and U24380 (N_24380,N_16952,N_15371);
and U24381 (N_24381,N_18950,N_16882);
and U24382 (N_24382,N_15266,N_18323);
nor U24383 (N_24383,N_15233,N_15971);
nand U24384 (N_24384,N_16513,N_18834);
xnor U24385 (N_24385,N_16750,N_15372);
or U24386 (N_24386,N_17939,N_17040);
and U24387 (N_24387,N_16056,N_17876);
nand U24388 (N_24388,N_15899,N_16246);
nand U24389 (N_24389,N_17239,N_17539);
xor U24390 (N_24390,N_19930,N_15091);
nand U24391 (N_24391,N_16076,N_15987);
xnor U24392 (N_24392,N_19253,N_17130);
xor U24393 (N_24393,N_19185,N_15431);
nor U24394 (N_24394,N_18811,N_15024);
nor U24395 (N_24395,N_17622,N_17673);
xnor U24396 (N_24396,N_18797,N_18628);
and U24397 (N_24397,N_17562,N_18708);
xor U24398 (N_24398,N_18681,N_16240);
and U24399 (N_24399,N_19671,N_16128);
xnor U24400 (N_24400,N_19710,N_18524);
xor U24401 (N_24401,N_17015,N_18124);
or U24402 (N_24402,N_16790,N_15715);
nand U24403 (N_24403,N_18134,N_17395);
nor U24404 (N_24404,N_19281,N_19701);
xor U24405 (N_24405,N_17725,N_15886);
or U24406 (N_24406,N_19232,N_15965);
and U24407 (N_24407,N_15192,N_18028);
xnor U24408 (N_24408,N_15526,N_15629);
nand U24409 (N_24409,N_16130,N_18448);
nor U24410 (N_24410,N_17083,N_18998);
or U24411 (N_24411,N_18151,N_16896);
or U24412 (N_24412,N_19812,N_19491);
nor U24413 (N_24413,N_16656,N_17424);
and U24414 (N_24414,N_19829,N_19646);
nand U24415 (N_24415,N_17420,N_17455);
xor U24416 (N_24416,N_17792,N_19192);
nand U24417 (N_24417,N_17323,N_17808);
or U24418 (N_24418,N_15997,N_18901);
nand U24419 (N_24419,N_16663,N_17159);
nor U24420 (N_24420,N_17644,N_19729);
xor U24421 (N_24421,N_15963,N_17570);
or U24422 (N_24422,N_19240,N_17967);
nand U24423 (N_24423,N_16122,N_16282);
or U24424 (N_24424,N_19319,N_17682);
nand U24425 (N_24425,N_19392,N_16351);
nor U24426 (N_24426,N_19270,N_17936);
nor U24427 (N_24427,N_16990,N_19205);
or U24428 (N_24428,N_16461,N_18551);
and U24429 (N_24429,N_16641,N_18254);
nor U24430 (N_24430,N_18616,N_18111);
and U24431 (N_24431,N_17041,N_16169);
nor U24432 (N_24432,N_16408,N_15872);
and U24433 (N_24433,N_18697,N_16285);
xnor U24434 (N_24434,N_16553,N_19490);
and U24435 (N_24435,N_16763,N_18757);
xnor U24436 (N_24436,N_18386,N_16719);
and U24437 (N_24437,N_19459,N_18953);
nor U24438 (N_24438,N_17072,N_19100);
and U24439 (N_24439,N_15603,N_16088);
nor U24440 (N_24440,N_19941,N_16871);
nor U24441 (N_24441,N_17806,N_17196);
and U24442 (N_24442,N_18095,N_17442);
and U24443 (N_24443,N_16641,N_18822);
xnor U24444 (N_24444,N_16706,N_16899);
nand U24445 (N_24445,N_17131,N_18990);
and U24446 (N_24446,N_15749,N_18107);
and U24447 (N_24447,N_15333,N_16152);
and U24448 (N_24448,N_15274,N_17029);
nor U24449 (N_24449,N_18992,N_15518);
xnor U24450 (N_24450,N_15587,N_17914);
nand U24451 (N_24451,N_16329,N_17872);
nor U24452 (N_24452,N_19425,N_19533);
and U24453 (N_24453,N_16951,N_19770);
and U24454 (N_24454,N_17090,N_18246);
or U24455 (N_24455,N_19747,N_18097);
nor U24456 (N_24456,N_18791,N_15515);
or U24457 (N_24457,N_17320,N_17057);
or U24458 (N_24458,N_18510,N_17017);
nand U24459 (N_24459,N_19126,N_15145);
xnor U24460 (N_24460,N_16788,N_19119);
nand U24461 (N_24461,N_17505,N_17145);
nand U24462 (N_24462,N_19160,N_16317);
xnor U24463 (N_24463,N_19096,N_19682);
and U24464 (N_24464,N_19084,N_15339);
nor U24465 (N_24465,N_16925,N_18964);
xor U24466 (N_24466,N_18675,N_17987);
xnor U24467 (N_24467,N_17265,N_19420);
or U24468 (N_24468,N_17419,N_18806);
xor U24469 (N_24469,N_18942,N_15512);
xnor U24470 (N_24470,N_15817,N_15244);
nor U24471 (N_24471,N_16326,N_18257);
nand U24472 (N_24472,N_17075,N_16794);
and U24473 (N_24473,N_17223,N_16934);
or U24474 (N_24474,N_15975,N_17591);
nor U24475 (N_24475,N_19141,N_15901);
or U24476 (N_24476,N_17743,N_18956);
nor U24477 (N_24477,N_18097,N_15737);
xnor U24478 (N_24478,N_16880,N_16118);
and U24479 (N_24479,N_16350,N_17350);
or U24480 (N_24480,N_18160,N_17183);
nor U24481 (N_24481,N_16130,N_18624);
xor U24482 (N_24482,N_19578,N_16479);
nor U24483 (N_24483,N_16311,N_19087);
or U24484 (N_24484,N_18363,N_16662);
nand U24485 (N_24485,N_15032,N_19431);
nand U24486 (N_24486,N_17776,N_19807);
and U24487 (N_24487,N_15869,N_15154);
nand U24488 (N_24488,N_15929,N_15349);
and U24489 (N_24489,N_16365,N_17174);
nor U24490 (N_24490,N_19817,N_16179);
and U24491 (N_24491,N_17200,N_19687);
or U24492 (N_24492,N_19756,N_17197);
or U24493 (N_24493,N_19897,N_16229);
nand U24494 (N_24494,N_19673,N_17402);
xnor U24495 (N_24495,N_15730,N_16720);
and U24496 (N_24496,N_19665,N_15834);
nor U24497 (N_24497,N_19183,N_18593);
and U24498 (N_24498,N_19088,N_16183);
nand U24499 (N_24499,N_16714,N_19172);
nand U24500 (N_24500,N_16193,N_17196);
xnor U24501 (N_24501,N_18400,N_15194);
nand U24502 (N_24502,N_15170,N_15687);
nand U24503 (N_24503,N_19609,N_18646);
or U24504 (N_24504,N_17425,N_18485);
xnor U24505 (N_24505,N_18106,N_16985);
and U24506 (N_24506,N_15470,N_15505);
and U24507 (N_24507,N_16187,N_19177);
nand U24508 (N_24508,N_17556,N_15738);
xnor U24509 (N_24509,N_15108,N_16727);
xor U24510 (N_24510,N_16581,N_19610);
nor U24511 (N_24511,N_18291,N_16306);
and U24512 (N_24512,N_15054,N_16630);
and U24513 (N_24513,N_18641,N_18434);
xnor U24514 (N_24514,N_17897,N_17374);
or U24515 (N_24515,N_18621,N_19445);
and U24516 (N_24516,N_18299,N_17885);
and U24517 (N_24517,N_15088,N_18809);
or U24518 (N_24518,N_19402,N_15076);
or U24519 (N_24519,N_17023,N_19735);
nand U24520 (N_24520,N_19133,N_16214);
or U24521 (N_24521,N_18154,N_17497);
xor U24522 (N_24522,N_18836,N_16473);
and U24523 (N_24523,N_18601,N_18909);
or U24524 (N_24524,N_19436,N_18548);
or U24525 (N_24525,N_16584,N_15923);
and U24526 (N_24526,N_19614,N_15000);
nor U24527 (N_24527,N_16279,N_19714);
nand U24528 (N_24528,N_16643,N_19144);
or U24529 (N_24529,N_18903,N_15735);
or U24530 (N_24530,N_15775,N_15060);
nand U24531 (N_24531,N_18631,N_17187);
and U24532 (N_24532,N_18432,N_16673);
and U24533 (N_24533,N_17050,N_17795);
and U24534 (N_24534,N_15055,N_16237);
or U24535 (N_24535,N_17425,N_16564);
or U24536 (N_24536,N_19808,N_19850);
or U24537 (N_24537,N_16585,N_16741);
nand U24538 (N_24538,N_19380,N_16106);
xnor U24539 (N_24539,N_19955,N_16571);
nor U24540 (N_24540,N_18521,N_16665);
and U24541 (N_24541,N_16977,N_19243);
nor U24542 (N_24542,N_18697,N_15084);
xor U24543 (N_24543,N_15224,N_17291);
xnor U24544 (N_24544,N_17004,N_15442);
nor U24545 (N_24545,N_19161,N_15642);
and U24546 (N_24546,N_19148,N_18494);
and U24547 (N_24547,N_16166,N_19172);
xor U24548 (N_24548,N_16709,N_19089);
and U24549 (N_24549,N_18061,N_16473);
nor U24550 (N_24550,N_15885,N_19520);
xor U24551 (N_24551,N_16842,N_16827);
nor U24552 (N_24552,N_19342,N_15221);
and U24553 (N_24553,N_16921,N_16978);
nand U24554 (N_24554,N_16132,N_15400);
nand U24555 (N_24555,N_15547,N_15417);
nand U24556 (N_24556,N_17637,N_15172);
or U24557 (N_24557,N_18494,N_18055);
xor U24558 (N_24558,N_18280,N_15076);
xor U24559 (N_24559,N_18432,N_16405);
nor U24560 (N_24560,N_18829,N_16550);
or U24561 (N_24561,N_19426,N_18986);
nand U24562 (N_24562,N_16597,N_19293);
nor U24563 (N_24563,N_18818,N_18237);
xor U24564 (N_24564,N_18454,N_18866);
nand U24565 (N_24565,N_18989,N_19959);
and U24566 (N_24566,N_17316,N_16363);
nor U24567 (N_24567,N_15280,N_16262);
nor U24568 (N_24568,N_18027,N_15019);
or U24569 (N_24569,N_19028,N_19587);
xnor U24570 (N_24570,N_19803,N_19725);
xor U24571 (N_24571,N_18151,N_16854);
or U24572 (N_24572,N_17315,N_15967);
or U24573 (N_24573,N_16047,N_19289);
and U24574 (N_24574,N_15388,N_17568);
or U24575 (N_24575,N_16780,N_18114);
xor U24576 (N_24576,N_15494,N_16880);
nor U24577 (N_24577,N_15781,N_15544);
or U24578 (N_24578,N_16722,N_18922);
xor U24579 (N_24579,N_19271,N_16115);
nand U24580 (N_24580,N_18454,N_17928);
or U24581 (N_24581,N_19018,N_15075);
nor U24582 (N_24582,N_15503,N_19018);
and U24583 (N_24583,N_15322,N_15732);
nand U24584 (N_24584,N_16313,N_18107);
and U24585 (N_24585,N_17587,N_15840);
or U24586 (N_24586,N_15462,N_19217);
nor U24587 (N_24587,N_15158,N_17032);
xnor U24588 (N_24588,N_17825,N_18578);
and U24589 (N_24589,N_18185,N_19873);
nor U24590 (N_24590,N_16009,N_19935);
nand U24591 (N_24591,N_19888,N_18828);
nor U24592 (N_24592,N_15441,N_15305);
xnor U24593 (N_24593,N_18093,N_18644);
and U24594 (N_24594,N_19296,N_17243);
nor U24595 (N_24595,N_15829,N_18690);
xnor U24596 (N_24596,N_18953,N_17055);
and U24597 (N_24597,N_15686,N_18860);
nand U24598 (N_24598,N_18708,N_15986);
nor U24599 (N_24599,N_15732,N_18815);
nand U24600 (N_24600,N_18231,N_17976);
nand U24601 (N_24601,N_17734,N_15649);
nand U24602 (N_24602,N_19829,N_15271);
or U24603 (N_24603,N_18025,N_19666);
nand U24604 (N_24604,N_18419,N_15859);
nor U24605 (N_24605,N_15465,N_15907);
nand U24606 (N_24606,N_18394,N_16967);
nor U24607 (N_24607,N_18904,N_18933);
and U24608 (N_24608,N_17225,N_15465);
and U24609 (N_24609,N_18088,N_19745);
xnor U24610 (N_24610,N_15384,N_18196);
or U24611 (N_24611,N_18679,N_15586);
xor U24612 (N_24612,N_16987,N_17048);
nor U24613 (N_24613,N_16689,N_18961);
xnor U24614 (N_24614,N_19787,N_19729);
nor U24615 (N_24615,N_17424,N_15695);
nor U24616 (N_24616,N_18766,N_19166);
xnor U24617 (N_24617,N_17956,N_16371);
nor U24618 (N_24618,N_15967,N_17077);
nand U24619 (N_24619,N_17082,N_18012);
or U24620 (N_24620,N_19111,N_18953);
or U24621 (N_24621,N_17923,N_19119);
and U24622 (N_24622,N_15349,N_19479);
or U24623 (N_24623,N_15003,N_15304);
and U24624 (N_24624,N_15767,N_15532);
or U24625 (N_24625,N_17652,N_16913);
xor U24626 (N_24626,N_19552,N_17767);
nand U24627 (N_24627,N_15142,N_16869);
xnor U24628 (N_24628,N_16646,N_19602);
and U24629 (N_24629,N_16325,N_17624);
and U24630 (N_24630,N_16085,N_17240);
and U24631 (N_24631,N_19609,N_15987);
nor U24632 (N_24632,N_17074,N_15419);
xor U24633 (N_24633,N_15603,N_16351);
nor U24634 (N_24634,N_15803,N_19328);
nand U24635 (N_24635,N_15271,N_16668);
or U24636 (N_24636,N_18872,N_15810);
or U24637 (N_24637,N_16452,N_19289);
and U24638 (N_24638,N_16547,N_15233);
nor U24639 (N_24639,N_17178,N_16058);
nand U24640 (N_24640,N_19174,N_17810);
and U24641 (N_24641,N_15936,N_19449);
xnor U24642 (N_24642,N_16054,N_17464);
nand U24643 (N_24643,N_16470,N_17337);
nand U24644 (N_24644,N_16062,N_15189);
nor U24645 (N_24645,N_17358,N_17260);
or U24646 (N_24646,N_19744,N_16322);
xor U24647 (N_24647,N_19752,N_16476);
xnor U24648 (N_24648,N_15829,N_17409);
nor U24649 (N_24649,N_17875,N_18209);
or U24650 (N_24650,N_16804,N_19056);
xnor U24651 (N_24651,N_19713,N_17073);
or U24652 (N_24652,N_17001,N_19907);
nand U24653 (N_24653,N_15483,N_19897);
nor U24654 (N_24654,N_16252,N_16071);
nand U24655 (N_24655,N_18289,N_17956);
nand U24656 (N_24656,N_16732,N_18954);
or U24657 (N_24657,N_15594,N_16825);
nor U24658 (N_24658,N_19930,N_17187);
or U24659 (N_24659,N_18794,N_18258);
nand U24660 (N_24660,N_19351,N_19236);
or U24661 (N_24661,N_16100,N_19643);
and U24662 (N_24662,N_19209,N_16994);
nor U24663 (N_24663,N_15596,N_18247);
nor U24664 (N_24664,N_18687,N_17967);
nand U24665 (N_24665,N_18636,N_18289);
or U24666 (N_24666,N_16931,N_19208);
or U24667 (N_24667,N_16626,N_16319);
nor U24668 (N_24668,N_17122,N_19763);
and U24669 (N_24669,N_19907,N_19910);
xnor U24670 (N_24670,N_15589,N_19018);
nand U24671 (N_24671,N_19997,N_17557);
xor U24672 (N_24672,N_17198,N_19591);
or U24673 (N_24673,N_16567,N_18038);
nor U24674 (N_24674,N_16255,N_16525);
nand U24675 (N_24675,N_16574,N_15789);
or U24676 (N_24676,N_18036,N_15484);
xor U24677 (N_24677,N_18662,N_18019);
xnor U24678 (N_24678,N_17036,N_18166);
nand U24679 (N_24679,N_16370,N_17160);
nand U24680 (N_24680,N_18433,N_18843);
or U24681 (N_24681,N_15626,N_19529);
xor U24682 (N_24682,N_19575,N_17757);
nor U24683 (N_24683,N_15971,N_16844);
xnor U24684 (N_24684,N_18834,N_16684);
nand U24685 (N_24685,N_18566,N_16021);
or U24686 (N_24686,N_17226,N_16236);
nor U24687 (N_24687,N_18249,N_19271);
or U24688 (N_24688,N_18712,N_15745);
or U24689 (N_24689,N_17060,N_19113);
and U24690 (N_24690,N_19175,N_18257);
nand U24691 (N_24691,N_18361,N_18941);
nor U24692 (N_24692,N_15639,N_15880);
xor U24693 (N_24693,N_17425,N_16998);
or U24694 (N_24694,N_17578,N_18153);
or U24695 (N_24695,N_19576,N_18558);
nor U24696 (N_24696,N_18985,N_18453);
or U24697 (N_24697,N_15496,N_16194);
or U24698 (N_24698,N_16145,N_15325);
xnor U24699 (N_24699,N_18327,N_17323);
nor U24700 (N_24700,N_19904,N_19103);
xnor U24701 (N_24701,N_16775,N_19041);
nand U24702 (N_24702,N_18241,N_16572);
or U24703 (N_24703,N_17811,N_17441);
nor U24704 (N_24704,N_17609,N_17395);
xor U24705 (N_24705,N_16364,N_19929);
or U24706 (N_24706,N_15560,N_15515);
and U24707 (N_24707,N_19694,N_15413);
nand U24708 (N_24708,N_16855,N_18247);
and U24709 (N_24709,N_18182,N_16984);
xor U24710 (N_24710,N_17425,N_17302);
or U24711 (N_24711,N_18698,N_15949);
nand U24712 (N_24712,N_19326,N_17165);
xor U24713 (N_24713,N_15271,N_17819);
or U24714 (N_24714,N_18449,N_16205);
nor U24715 (N_24715,N_19479,N_15544);
xor U24716 (N_24716,N_17207,N_19144);
nor U24717 (N_24717,N_15758,N_18746);
and U24718 (N_24718,N_19930,N_17914);
nand U24719 (N_24719,N_18016,N_18630);
or U24720 (N_24720,N_19865,N_17798);
nor U24721 (N_24721,N_19552,N_16778);
nor U24722 (N_24722,N_17528,N_16308);
or U24723 (N_24723,N_17430,N_15105);
and U24724 (N_24724,N_17856,N_16014);
or U24725 (N_24725,N_15664,N_18017);
nand U24726 (N_24726,N_16714,N_18651);
nor U24727 (N_24727,N_18914,N_16157);
and U24728 (N_24728,N_18843,N_19660);
or U24729 (N_24729,N_16815,N_19049);
xnor U24730 (N_24730,N_16395,N_19584);
xor U24731 (N_24731,N_19837,N_18415);
nand U24732 (N_24732,N_15377,N_15334);
or U24733 (N_24733,N_16053,N_19003);
nand U24734 (N_24734,N_18128,N_17980);
xnor U24735 (N_24735,N_17862,N_15381);
or U24736 (N_24736,N_15874,N_19745);
nor U24737 (N_24737,N_15573,N_15471);
or U24738 (N_24738,N_19657,N_15713);
or U24739 (N_24739,N_16378,N_17212);
xnor U24740 (N_24740,N_18303,N_19310);
nand U24741 (N_24741,N_19961,N_18187);
xor U24742 (N_24742,N_17536,N_19011);
nand U24743 (N_24743,N_19646,N_17752);
xor U24744 (N_24744,N_15965,N_18309);
xnor U24745 (N_24745,N_15232,N_19559);
or U24746 (N_24746,N_18334,N_17090);
nand U24747 (N_24747,N_16776,N_17058);
and U24748 (N_24748,N_18427,N_19339);
or U24749 (N_24749,N_15869,N_18697);
and U24750 (N_24750,N_15931,N_15545);
xnor U24751 (N_24751,N_17044,N_19692);
or U24752 (N_24752,N_17954,N_17347);
xor U24753 (N_24753,N_19028,N_15213);
xor U24754 (N_24754,N_18790,N_16929);
or U24755 (N_24755,N_17923,N_17766);
or U24756 (N_24756,N_18915,N_15875);
xor U24757 (N_24757,N_19842,N_17904);
or U24758 (N_24758,N_18408,N_15379);
and U24759 (N_24759,N_15132,N_16464);
nor U24760 (N_24760,N_18445,N_17710);
nand U24761 (N_24761,N_17916,N_17762);
xnor U24762 (N_24762,N_19444,N_18273);
nor U24763 (N_24763,N_17651,N_15367);
nor U24764 (N_24764,N_19200,N_19652);
and U24765 (N_24765,N_17904,N_15684);
xor U24766 (N_24766,N_19426,N_16376);
xor U24767 (N_24767,N_15056,N_18496);
and U24768 (N_24768,N_15393,N_15482);
nand U24769 (N_24769,N_16502,N_18907);
nor U24770 (N_24770,N_17458,N_17196);
nand U24771 (N_24771,N_18011,N_15086);
or U24772 (N_24772,N_17677,N_18046);
or U24773 (N_24773,N_17876,N_17161);
and U24774 (N_24774,N_15670,N_19085);
xnor U24775 (N_24775,N_16013,N_19899);
and U24776 (N_24776,N_19342,N_19220);
xnor U24777 (N_24777,N_19854,N_19920);
nand U24778 (N_24778,N_19947,N_17139);
nor U24779 (N_24779,N_18097,N_19162);
or U24780 (N_24780,N_16908,N_18523);
xor U24781 (N_24781,N_16818,N_15074);
or U24782 (N_24782,N_19187,N_18975);
xor U24783 (N_24783,N_15086,N_17537);
nor U24784 (N_24784,N_17705,N_19016);
xnor U24785 (N_24785,N_15288,N_19153);
xor U24786 (N_24786,N_18599,N_15996);
and U24787 (N_24787,N_19662,N_18104);
xor U24788 (N_24788,N_17822,N_18559);
nor U24789 (N_24789,N_15035,N_19256);
xnor U24790 (N_24790,N_17352,N_16468);
nand U24791 (N_24791,N_15166,N_15633);
nor U24792 (N_24792,N_16734,N_15439);
nor U24793 (N_24793,N_19445,N_15630);
and U24794 (N_24794,N_18657,N_19670);
nand U24795 (N_24795,N_15628,N_15546);
nor U24796 (N_24796,N_18922,N_15129);
nor U24797 (N_24797,N_15732,N_16307);
or U24798 (N_24798,N_19071,N_17015);
nor U24799 (N_24799,N_17738,N_15911);
nand U24800 (N_24800,N_17468,N_16903);
nand U24801 (N_24801,N_19537,N_16594);
and U24802 (N_24802,N_17649,N_18633);
and U24803 (N_24803,N_18957,N_16429);
or U24804 (N_24804,N_15583,N_19326);
nand U24805 (N_24805,N_18476,N_15224);
nand U24806 (N_24806,N_18800,N_15546);
nand U24807 (N_24807,N_19697,N_19924);
nor U24808 (N_24808,N_16151,N_17215);
nand U24809 (N_24809,N_16013,N_15214);
xnor U24810 (N_24810,N_18963,N_17852);
xnor U24811 (N_24811,N_18931,N_19613);
and U24812 (N_24812,N_16416,N_19101);
and U24813 (N_24813,N_18078,N_17697);
nor U24814 (N_24814,N_17907,N_15367);
xnor U24815 (N_24815,N_17806,N_18519);
nor U24816 (N_24816,N_18642,N_16987);
xnor U24817 (N_24817,N_19295,N_18353);
and U24818 (N_24818,N_17764,N_16101);
nand U24819 (N_24819,N_16473,N_15867);
and U24820 (N_24820,N_17054,N_18474);
xor U24821 (N_24821,N_17923,N_19325);
nand U24822 (N_24822,N_18027,N_18584);
or U24823 (N_24823,N_17748,N_19208);
xnor U24824 (N_24824,N_18551,N_15073);
nor U24825 (N_24825,N_15591,N_15097);
nand U24826 (N_24826,N_16668,N_16335);
or U24827 (N_24827,N_19538,N_15063);
and U24828 (N_24828,N_18901,N_15053);
nor U24829 (N_24829,N_18459,N_15158);
and U24830 (N_24830,N_15101,N_18133);
or U24831 (N_24831,N_17887,N_16204);
and U24832 (N_24832,N_17954,N_19203);
xor U24833 (N_24833,N_19758,N_18752);
or U24834 (N_24834,N_18881,N_16613);
or U24835 (N_24835,N_18128,N_17844);
nor U24836 (N_24836,N_15083,N_15400);
nor U24837 (N_24837,N_19837,N_17319);
xnor U24838 (N_24838,N_16935,N_19044);
or U24839 (N_24839,N_16854,N_17084);
xnor U24840 (N_24840,N_18552,N_16523);
and U24841 (N_24841,N_18504,N_15608);
or U24842 (N_24842,N_17273,N_18101);
nand U24843 (N_24843,N_16008,N_17826);
or U24844 (N_24844,N_17685,N_17723);
nor U24845 (N_24845,N_19669,N_19555);
nor U24846 (N_24846,N_15412,N_15025);
xor U24847 (N_24847,N_19016,N_16461);
nand U24848 (N_24848,N_16731,N_19453);
or U24849 (N_24849,N_18579,N_15967);
and U24850 (N_24850,N_19456,N_19091);
and U24851 (N_24851,N_15274,N_18779);
xor U24852 (N_24852,N_16547,N_19092);
xnor U24853 (N_24853,N_15770,N_18865);
xnor U24854 (N_24854,N_17027,N_19821);
nand U24855 (N_24855,N_16897,N_19065);
or U24856 (N_24856,N_17242,N_18394);
nand U24857 (N_24857,N_19094,N_18220);
xnor U24858 (N_24858,N_19091,N_18937);
or U24859 (N_24859,N_17065,N_16927);
nand U24860 (N_24860,N_17154,N_16922);
nor U24861 (N_24861,N_15655,N_18859);
nand U24862 (N_24862,N_19876,N_16066);
or U24863 (N_24863,N_17796,N_15113);
and U24864 (N_24864,N_15030,N_17728);
or U24865 (N_24865,N_19427,N_15387);
and U24866 (N_24866,N_17284,N_16341);
and U24867 (N_24867,N_18670,N_15920);
xor U24868 (N_24868,N_16733,N_16381);
or U24869 (N_24869,N_15220,N_17518);
or U24870 (N_24870,N_18656,N_17672);
and U24871 (N_24871,N_16899,N_15147);
nor U24872 (N_24872,N_19309,N_17887);
nand U24873 (N_24873,N_15848,N_15570);
or U24874 (N_24874,N_15676,N_15076);
or U24875 (N_24875,N_19218,N_18761);
and U24876 (N_24876,N_18630,N_16989);
nor U24877 (N_24877,N_18352,N_18755);
xor U24878 (N_24878,N_17455,N_18409);
and U24879 (N_24879,N_15313,N_15855);
nor U24880 (N_24880,N_17788,N_19938);
nor U24881 (N_24881,N_19666,N_16017);
xnor U24882 (N_24882,N_18502,N_19354);
xor U24883 (N_24883,N_19059,N_19366);
nand U24884 (N_24884,N_15459,N_17104);
and U24885 (N_24885,N_17036,N_15393);
nand U24886 (N_24886,N_16025,N_17835);
nor U24887 (N_24887,N_15530,N_18263);
nand U24888 (N_24888,N_16238,N_18227);
or U24889 (N_24889,N_15435,N_16670);
xnor U24890 (N_24890,N_15802,N_18124);
nand U24891 (N_24891,N_15569,N_16430);
or U24892 (N_24892,N_19779,N_15773);
and U24893 (N_24893,N_19572,N_17294);
xnor U24894 (N_24894,N_19677,N_16389);
or U24895 (N_24895,N_18697,N_19383);
xnor U24896 (N_24896,N_18999,N_15141);
nand U24897 (N_24897,N_19299,N_17836);
and U24898 (N_24898,N_16751,N_17170);
and U24899 (N_24899,N_18253,N_15671);
nand U24900 (N_24900,N_16398,N_16235);
or U24901 (N_24901,N_17570,N_19157);
nand U24902 (N_24902,N_17398,N_19856);
xnor U24903 (N_24903,N_16693,N_16863);
and U24904 (N_24904,N_16393,N_19578);
nor U24905 (N_24905,N_16941,N_16599);
or U24906 (N_24906,N_17105,N_19524);
nand U24907 (N_24907,N_19803,N_18272);
nor U24908 (N_24908,N_18702,N_19349);
nand U24909 (N_24909,N_17188,N_18705);
nand U24910 (N_24910,N_19435,N_19134);
or U24911 (N_24911,N_18955,N_15551);
xor U24912 (N_24912,N_16555,N_18361);
xnor U24913 (N_24913,N_19754,N_16104);
or U24914 (N_24914,N_16739,N_18463);
or U24915 (N_24915,N_18246,N_17560);
nor U24916 (N_24916,N_16658,N_15389);
and U24917 (N_24917,N_16988,N_17743);
or U24918 (N_24918,N_17050,N_16328);
nor U24919 (N_24919,N_15070,N_18671);
and U24920 (N_24920,N_17915,N_17805);
and U24921 (N_24921,N_19383,N_19483);
xnor U24922 (N_24922,N_16750,N_16824);
and U24923 (N_24923,N_17017,N_15026);
nor U24924 (N_24924,N_16674,N_16996);
xnor U24925 (N_24925,N_18749,N_16442);
xor U24926 (N_24926,N_19997,N_17094);
and U24927 (N_24927,N_17335,N_19766);
nor U24928 (N_24928,N_18487,N_17411);
nand U24929 (N_24929,N_16608,N_18698);
nor U24930 (N_24930,N_19878,N_16534);
or U24931 (N_24931,N_15190,N_18443);
xnor U24932 (N_24932,N_19285,N_19098);
xor U24933 (N_24933,N_17464,N_18351);
xnor U24934 (N_24934,N_16988,N_19829);
nand U24935 (N_24935,N_17718,N_17339);
or U24936 (N_24936,N_18932,N_15698);
xor U24937 (N_24937,N_16299,N_17863);
or U24938 (N_24938,N_19272,N_18338);
or U24939 (N_24939,N_15767,N_18656);
xnor U24940 (N_24940,N_15343,N_19869);
and U24941 (N_24941,N_17424,N_18131);
nand U24942 (N_24942,N_19722,N_19334);
and U24943 (N_24943,N_19490,N_19380);
or U24944 (N_24944,N_15593,N_16292);
nand U24945 (N_24945,N_19436,N_18795);
or U24946 (N_24946,N_18618,N_16732);
nand U24947 (N_24947,N_18922,N_18251);
or U24948 (N_24948,N_17568,N_17082);
xnor U24949 (N_24949,N_19409,N_17812);
or U24950 (N_24950,N_19947,N_15444);
nor U24951 (N_24951,N_19735,N_15021);
or U24952 (N_24952,N_15795,N_19021);
xor U24953 (N_24953,N_16478,N_16423);
nor U24954 (N_24954,N_19638,N_15232);
or U24955 (N_24955,N_16762,N_16777);
and U24956 (N_24956,N_18175,N_18390);
xnor U24957 (N_24957,N_17231,N_18008);
and U24958 (N_24958,N_17574,N_19725);
nor U24959 (N_24959,N_15513,N_17264);
nor U24960 (N_24960,N_18841,N_19172);
nand U24961 (N_24961,N_19779,N_17291);
and U24962 (N_24962,N_15323,N_17895);
or U24963 (N_24963,N_17909,N_18766);
nor U24964 (N_24964,N_15660,N_17453);
nand U24965 (N_24965,N_19412,N_18102);
or U24966 (N_24966,N_19701,N_19413);
xnor U24967 (N_24967,N_18693,N_15159);
and U24968 (N_24968,N_15886,N_17549);
or U24969 (N_24969,N_16578,N_17507);
or U24970 (N_24970,N_19256,N_16119);
xor U24971 (N_24971,N_18798,N_16904);
nand U24972 (N_24972,N_18329,N_16831);
nand U24973 (N_24973,N_15798,N_16257);
xor U24974 (N_24974,N_17872,N_15211);
or U24975 (N_24975,N_17812,N_18737);
nand U24976 (N_24976,N_17922,N_19906);
nor U24977 (N_24977,N_17736,N_15127);
or U24978 (N_24978,N_16601,N_15412);
or U24979 (N_24979,N_17570,N_16616);
nor U24980 (N_24980,N_18224,N_15364);
nor U24981 (N_24981,N_17880,N_16047);
nor U24982 (N_24982,N_16901,N_17280);
and U24983 (N_24983,N_16066,N_19907);
and U24984 (N_24984,N_19733,N_17865);
or U24985 (N_24985,N_16799,N_19953);
and U24986 (N_24986,N_19066,N_18349);
or U24987 (N_24987,N_17563,N_15212);
and U24988 (N_24988,N_16631,N_17242);
and U24989 (N_24989,N_18202,N_17229);
or U24990 (N_24990,N_19669,N_18265);
nand U24991 (N_24991,N_16448,N_17860);
nor U24992 (N_24992,N_19350,N_16167);
nor U24993 (N_24993,N_17183,N_19955);
or U24994 (N_24994,N_16146,N_19719);
xnor U24995 (N_24995,N_19578,N_17031);
and U24996 (N_24996,N_17328,N_17802);
or U24997 (N_24997,N_17122,N_15028);
and U24998 (N_24998,N_16897,N_19724);
and U24999 (N_24999,N_18361,N_15431);
or U25000 (N_25000,N_24393,N_22702);
and U25001 (N_25001,N_23101,N_20351);
and U25002 (N_25002,N_24715,N_23469);
or U25003 (N_25003,N_21771,N_23372);
nor U25004 (N_25004,N_22569,N_24823);
nor U25005 (N_25005,N_22220,N_20867);
nor U25006 (N_25006,N_20022,N_21011);
xnor U25007 (N_25007,N_21733,N_24280);
or U25008 (N_25008,N_22011,N_24883);
xnor U25009 (N_25009,N_21339,N_24077);
and U25010 (N_25010,N_20647,N_22143);
and U25011 (N_25011,N_24194,N_21263);
and U25012 (N_25012,N_22822,N_22033);
nand U25013 (N_25013,N_22082,N_21217);
and U25014 (N_25014,N_22016,N_24915);
and U25015 (N_25015,N_21211,N_20207);
nor U25016 (N_25016,N_20635,N_20159);
and U25017 (N_25017,N_21187,N_22365);
nor U25018 (N_25018,N_21083,N_21895);
xnor U25019 (N_25019,N_20711,N_23261);
xnor U25020 (N_25020,N_21893,N_21849);
nor U25021 (N_25021,N_22744,N_24047);
nand U25022 (N_25022,N_22669,N_21617);
nand U25023 (N_25023,N_24130,N_21111);
nand U25024 (N_25024,N_20276,N_20309);
nor U25025 (N_25025,N_20496,N_22936);
nor U25026 (N_25026,N_22765,N_22230);
xor U25027 (N_25027,N_21941,N_22182);
xnor U25028 (N_25028,N_22328,N_21380);
xor U25029 (N_25029,N_20190,N_20410);
nand U25030 (N_25030,N_21913,N_21678);
and U25031 (N_25031,N_21527,N_23939);
nor U25032 (N_25032,N_20825,N_20521);
nor U25033 (N_25033,N_20893,N_24162);
xnor U25034 (N_25034,N_21786,N_23843);
nand U25035 (N_25035,N_23321,N_22334);
nand U25036 (N_25036,N_23876,N_22157);
xnor U25037 (N_25037,N_20203,N_22199);
nor U25038 (N_25038,N_22565,N_20609);
nand U25039 (N_25039,N_22452,N_23176);
nand U25040 (N_25040,N_23557,N_20117);
xnor U25041 (N_25041,N_20691,N_20097);
nand U25042 (N_25042,N_20044,N_21706);
xor U25043 (N_25043,N_20934,N_23930);
nand U25044 (N_25044,N_22192,N_23524);
nor U25045 (N_25045,N_21062,N_22960);
and U25046 (N_25046,N_22293,N_21983);
nand U25047 (N_25047,N_21647,N_20056);
xnor U25048 (N_25048,N_20155,N_20313);
nor U25049 (N_25049,N_24145,N_22791);
or U25050 (N_25050,N_22392,N_23960);
xnor U25051 (N_25051,N_20085,N_22172);
xor U25052 (N_25052,N_22857,N_23977);
or U25053 (N_25053,N_24377,N_20167);
nand U25054 (N_25054,N_24778,N_23394);
nor U25055 (N_25055,N_21725,N_20606);
and U25056 (N_25056,N_20094,N_23779);
nand U25057 (N_25057,N_21794,N_20418);
and U25058 (N_25058,N_22507,N_20806);
xnor U25059 (N_25059,N_21775,N_20474);
nor U25060 (N_25060,N_21743,N_20305);
xor U25061 (N_25061,N_20288,N_24269);
xnor U25062 (N_25062,N_21136,N_21076);
nand U25063 (N_25063,N_20198,N_24131);
nor U25064 (N_25064,N_24200,N_24770);
nand U25065 (N_25065,N_21521,N_24273);
nor U25066 (N_25066,N_24467,N_21180);
xor U25067 (N_25067,N_22484,N_21319);
and U25068 (N_25068,N_22440,N_21084);
nand U25069 (N_25069,N_23377,N_23645);
and U25070 (N_25070,N_20476,N_20661);
xnor U25071 (N_25071,N_20592,N_24650);
nand U25072 (N_25072,N_20212,N_22542);
nor U25073 (N_25073,N_20375,N_24511);
and U25074 (N_25074,N_21590,N_22938);
and U25075 (N_25075,N_24870,N_21618);
xnor U25076 (N_25076,N_22879,N_20561);
nand U25077 (N_25077,N_20982,N_20581);
and U25078 (N_25078,N_23154,N_20277);
xor U25079 (N_25079,N_24251,N_20736);
and U25080 (N_25080,N_24873,N_21230);
nand U25081 (N_25081,N_22799,N_23126);
nand U25082 (N_25082,N_20243,N_23034);
nor U25083 (N_25083,N_22428,N_22013);
or U25084 (N_25084,N_24239,N_22890);
xor U25085 (N_25085,N_21249,N_21114);
or U25086 (N_25086,N_23453,N_22470);
and U25087 (N_25087,N_22572,N_20009);
nor U25088 (N_25088,N_22737,N_21562);
nand U25089 (N_25089,N_20692,N_21443);
nand U25090 (N_25090,N_20978,N_23595);
nand U25091 (N_25091,N_20485,N_23364);
and U25092 (N_25092,N_24332,N_21639);
or U25093 (N_25093,N_23800,N_23974);
xnor U25094 (N_25094,N_20785,N_20761);
nand U25095 (N_25095,N_24104,N_22102);
nor U25096 (N_25096,N_21251,N_24308);
nand U25097 (N_25097,N_21985,N_20384);
nand U25098 (N_25098,N_23159,N_20489);
nor U25099 (N_25099,N_22894,N_24385);
or U25100 (N_25100,N_24493,N_24381);
and U25101 (N_25101,N_21392,N_24938);
or U25102 (N_25102,N_20929,N_20076);
nor U25103 (N_25103,N_20311,N_22841);
or U25104 (N_25104,N_20787,N_21505);
nand U25105 (N_25105,N_20471,N_21470);
or U25106 (N_25106,N_23702,N_23692);
nor U25107 (N_25107,N_22296,N_23167);
xnor U25108 (N_25108,N_22308,N_21550);
nor U25109 (N_25109,N_21624,N_23265);
nand U25110 (N_25110,N_22026,N_23521);
or U25111 (N_25111,N_21595,N_22282);
or U25112 (N_25112,N_23467,N_20163);
xor U25113 (N_25113,N_22653,N_20538);
nand U25114 (N_25114,N_23984,N_21195);
or U25115 (N_25115,N_24451,N_20646);
or U25116 (N_25116,N_20179,N_23349);
nor U25117 (N_25117,N_21432,N_23809);
or U25118 (N_25118,N_22492,N_22885);
xor U25119 (N_25119,N_24372,N_23587);
xor U25120 (N_25120,N_22895,N_22110);
nor U25121 (N_25121,N_21353,N_24815);
nor U25122 (N_25122,N_24238,N_24888);
nor U25123 (N_25123,N_20693,N_24617);
and U25124 (N_25124,N_23037,N_20219);
xnor U25125 (N_25125,N_24098,N_22394);
xor U25126 (N_25126,N_20140,N_23153);
and U25127 (N_25127,N_20405,N_24429);
or U25128 (N_25128,N_23156,N_21078);
or U25129 (N_25129,N_22886,N_24327);
or U25130 (N_25130,N_23796,N_24922);
or U25131 (N_25131,N_24808,N_24401);
and U25132 (N_25132,N_24809,N_24171);
and U25133 (N_25133,N_24025,N_20686);
xnor U25134 (N_25134,N_22391,N_24363);
nand U25135 (N_25135,N_23805,N_21253);
nor U25136 (N_25136,N_21435,N_21368);
nand U25137 (N_25137,N_21707,N_21371);
nand U25138 (N_25138,N_21765,N_22548);
nand U25139 (N_25139,N_20863,N_22657);
nor U25140 (N_25140,N_24271,N_21218);
nor U25141 (N_25141,N_20017,N_24101);
nor U25142 (N_25142,N_22378,N_23452);
nor U25143 (N_25143,N_20100,N_22380);
or U25144 (N_25144,N_23554,N_23963);
and U25145 (N_25145,N_24865,N_24080);
xnor U25146 (N_25146,N_23282,N_21287);
xor U25147 (N_25147,N_24060,N_21580);
xor U25148 (N_25148,N_20506,N_24800);
and U25149 (N_25149,N_20573,N_20965);
nor U25150 (N_25150,N_23711,N_22904);
xor U25151 (N_25151,N_24563,N_21953);
or U25152 (N_25152,N_23513,N_20949);
and U25153 (N_25153,N_24330,N_21623);
and U25154 (N_25154,N_21110,N_24927);
and U25155 (N_25155,N_24796,N_24916);
nand U25156 (N_25156,N_24484,N_21594);
xor U25157 (N_25157,N_24675,N_24586);
nand U25158 (N_25158,N_24083,N_20399);
xnor U25159 (N_25159,N_22459,N_20388);
nand U25160 (N_25160,N_23373,N_22336);
nor U25161 (N_25161,N_24782,N_20067);
nor U25162 (N_25162,N_24395,N_23136);
or U25163 (N_25163,N_21256,N_24154);
and U25164 (N_25164,N_20481,N_23205);
and U25165 (N_25165,N_23708,N_24213);
nand U25166 (N_25166,N_24307,N_21300);
nor U25167 (N_25167,N_24984,N_20618);
or U25168 (N_25168,N_24411,N_23689);
xnor U25169 (N_25169,N_22774,N_20781);
and U25170 (N_25170,N_23317,N_21607);
and U25171 (N_25171,N_20411,N_21665);
nand U25172 (N_25172,N_23088,N_21567);
nand U25173 (N_25173,N_24515,N_22224);
nand U25174 (N_25174,N_20404,N_23532);
nor U25175 (N_25175,N_21871,N_23393);
nand U25176 (N_25176,N_20488,N_21266);
nor U25177 (N_25177,N_24476,N_22750);
and U25178 (N_25178,N_22728,N_24718);
xor U25179 (N_25179,N_24084,N_20387);
nand U25180 (N_25180,N_21762,N_20712);
nor U25181 (N_25181,N_23725,N_20259);
nor U25182 (N_25182,N_24082,N_22173);
xnor U25183 (N_25183,N_21800,N_20298);
or U25184 (N_25184,N_23878,N_23854);
and U25185 (N_25185,N_22783,N_23647);
and U25186 (N_25186,N_24024,N_21431);
xor U25187 (N_25187,N_24420,N_22880);
nand U25188 (N_25188,N_21804,N_21902);
and U25189 (N_25189,N_21449,N_23583);
xnor U25190 (N_25190,N_22957,N_22631);
and U25191 (N_25191,N_23161,N_23838);
or U25192 (N_25192,N_23486,N_24753);
and U25193 (N_25193,N_23560,N_23283);
xnor U25194 (N_25194,N_23918,N_23801);
nand U25195 (N_25195,N_20397,N_21887);
or U25196 (N_25196,N_22818,N_22761);
nand U25197 (N_25197,N_20162,N_24015);
or U25198 (N_25198,N_23183,N_21519);
or U25199 (N_25199,N_24551,N_20241);
nor U25200 (N_25200,N_23526,N_21198);
or U25201 (N_25201,N_20558,N_22313);
xnor U25202 (N_25202,N_20373,N_22395);
nor U25203 (N_25203,N_22151,N_23889);
nor U25204 (N_25204,N_22367,N_21296);
or U25205 (N_25205,N_24817,N_22208);
xor U25206 (N_25206,N_20763,N_22701);
and U25207 (N_25207,N_24703,N_22798);
nor U25208 (N_25208,N_24295,N_21019);
and U25209 (N_25209,N_22696,N_24137);
and U25210 (N_25210,N_23097,N_22118);
and U25211 (N_25211,N_21112,N_22248);
or U25212 (N_25212,N_20619,N_22431);
and U25213 (N_25213,N_22086,N_21508);
xnor U25214 (N_25214,N_22320,N_22920);
nand U25215 (N_25215,N_23813,N_22268);
nor U25216 (N_25216,N_22022,N_21089);
and U25217 (N_25217,N_23203,N_21032);
xnor U25218 (N_25218,N_23451,N_20026);
nor U25219 (N_25219,N_22836,N_24813);
or U25220 (N_25220,N_20180,N_24366);
xnor U25221 (N_25221,N_21829,N_22263);
or U25222 (N_25222,N_22083,N_20264);
nor U25223 (N_25223,N_21143,N_24686);
nand U25224 (N_25224,N_22374,N_21675);
nor U25225 (N_25225,N_23440,N_21097);
nor U25226 (N_25226,N_23051,N_22029);
and U25227 (N_25227,N_21051,N_22150);
xor U25228 (N_25228,N_22437,N_23833);
nand U25229 (N_25229,N_24757,N_20598);
or U25230 (N_25230,N_23934,N_22038);
nand U25231 (N_25231,N_24764,N_24720);
and U25232 (N_25232,N_24323,N_20060);
nand U25233 (N_25233,N_21163,N_24204);
nand U25234 (N_25234,N_21117,N_22454);
nor U25235 (N_25235,N_22021,N_21899);
or U25236 (N_25236,N_22863,N_21377);
nor U25237 (N_25237,N_23650,N_21701);
nand U25238 (N_25238,N_23040,N_22800);
and U25239 (N_25239,N_23551,N_20877);
or U25240 (N_25240,N_23999,N_23470);
nor U25241 (N_25241,N_20096,N_21576);
nand U25242 (N_25242,N_23355,N_22581);
or U25243 (N_25243,N_20317,N_22113);
and U25244 (N_25244,N_23318,N_20034);
nor U25245 (N_25245,N_21667,N_20192);
xor U25246 (N_25246,N_20665,N_21252);
and U25247 (N_25247,N_22429,N_21669);
and U25248 (N_25248,N_23535,N_22796);
and U25249 (N_25249,N_20401,N_21149);
and U25250 (N_25250,N_23382,N_22499);
and U25251 (N_25251,N_22658,N_23910);
xnor U25252 (N_25252,N_20783,N_23973);
and U25253 (N_25253,N_21698,N_21175);
nor U25254 (N_25254,N_24948,N_22784);
nand U25255 (N_25255,N_22971,N_22698);
nor U25256 (N_25256,N_23134,N_24472);
and U25257 (N_25257,N_23057,N_21789);
nor U25258 (N_25258,N_21404,N_21462);
nand U25259 (N_25259,N_21104,N_21079);
xor U25260 (N_25260,N_24187,N_21495);
or U25261 (N_25261,N_20986,N_20260);
or U25262 (N_25262,N_22115,N_20346);
nand U25263 (N_25263,N_24211,N_23292);
xnor U25264 (N_25264,N_21416,N_22103);
xnor U25265 (N_25265,N_20879,N_24731);
and U25266 (N_25266,N_22238,N_20347);
nand U25267 (N_25267,N_22606,N_23543);
or U25268 (N_25268,N_21972,N_22571);
xor U25269 (N_25269,N_23464,N_22725);
nand U25270 (N_25270,N_24603,N_20383);
or U25271 (N_25271,N_20750,N_20331);
or U25272 (N_25272,N_21182,N_21629);
xnor U25273 (N_25273,N_22262,N_24422);
and U25274 (N_25274,N_24655,N_22662);
or U25275 (N_25275,N_24249,N_20283);
xnor U25276 (N_25276,N_21073,N_21127);
xnor U25277 (N_25277,N_23785,N_22844);
or U25278 (N_25278,N_24337,N_22469);
or U25279 (N_25279,N_20895,N_21812);
nor U25280 (N_25280,N_24351,N_24890);
and U25281 (N_25281,N_21239,N_21369);
and U25282 (N_25282,N_23108,N_22372);
xor U25283 (N_25283,N_21275,N_20596);
nand U25284 (N_25284,N_21709,N_22384);
nor U25285 (N_25285,N_23494,N_22495);
nand U25286 (N_25286,N_20544,N_20040);
xor U25287 (N_25287,N_21003,N_23314);
and U25288 (N_25288,N_23958,N_24496);
xnor U25289 (N_25289,N_22279,N_23380);
or U25290 (N_25290,N_20003,N_20977);
nand U25291 (N_25291,N_22382,N_22540);
nor U25292 (N_25292,N_21419,N_21407);
nor U25293 (N_25293,N_23155,N_24860);
and U25294 (N_25294,N_23832,N_24446);
nand U25295 (N_25295,N_21254,N_23143);
nor U25296 (N_25296,N_24886,N_21870);
and U25297 (N_25297,N_24898,N_21139);
nor U25298 (N_25298,N_21183,N_23677);
and U25299 (N_25299,N_23240,N_20339);
xnor U25300 (N_25300,N_24042,N_20823);
or U25301 (N_25301,N_23403,N_22060);
and U25302 (N_25302,N_21710,N_24168);
or U25303 (N_25303,N_24125,N_20894);
nor U25304 (N_25304,N_24447,N_21045);
xnor U25305 (N_25305,N_24975,N_20111);
and U25306 (N_25306,N_20591,N_21986);
xor U25307 (N_25307,N_24169,N_21224);
or U25308 (N_25308,N_22842,N_22030);
xor U25309 (N_25309,N_24135,N_22341);
nor U25310 (N_25310,N_23411,N_24998);
and U25311 (N_25311,N_21900,N_24606);
xnor U25312 (N_25312,N_21481,N_23309);
nor U25313 (N_25313,N_23625,N_21781);
and U25314 (N_25314,N_23684,N_24408);
nand U25315 (N_25315,N_23267,N_22421);
and U25316 (N_25316,N_20108,N_23922);
nor U25317 (N_25317,N_21641,N_21642);
or U25318 (N_25318,N_21277,N_23271);
or U25319 (N_25319,N_22543,N_23447);
xnor U25320 (N_25320,N_21290,N_22075);
and U25321 (N_25321,N_23158,N_20683);
nor U25322 (N_25322,N_20286,N_20116);
nand U25323 (N_25323,N_23496,N_22637);
nand U25324 (N_25324,N_22810,N_22611);
and U25325 (N_25325,N_20466,N_21199);
nor U25326 (N_25326,N_22024,N_23190);
nand U25327 (N_25327,N_20278,N_24839);
or U25328 (N_25328,N_22181,N_24387);
nor U25329 (N_25329,N_22237,N_24854);
xnor U25330 (N_25330,N_20795,N_22404);
nand U25331 (N_25331,N_20898,N_22628);
and U25332 (N_25332,N_21044,N_22813);
nor U25333 (N_25333,N_20627,N_20991);
and U25334 (N_25334,N_21480,N_24626);
nand U25335 (N_25335,N_22360,N_20491);
nor U25336 (N_25336,N_22937,N_24265);
or U25337 (N_25337,N_20704,N_21945);
and U25338 (N_25338,N_24569,N_20943);
and U25339 (N_25339,N_22315,N_23198);
xor U25340 (N_25340,N_20587,N_22125);
xnor U25341 (N_25341,N_20394,N_24999);
xnor U25342 (N_25342,N_24222,N_23252);
nand U25343 (N_25343,N_23301,N_24763);
xor U25344 (N_25344,N_21050,N_21714);
or U25345 (N_25345,N_24061,N_20759);
xnor U25346 (N_25346,N_24348,N_22035);
or U25347 (N_25347,N_20451,N_23682);
or U25348 (N_25348,N_22148,N_21763);
nand U25349 (N_25349,N_24797,N_24837);
and U25350 (N_25350,N_20454,N_21342);
and U25351 (N_25351,N_22646,N_23588);
xor U25352 (N_25352,N_23771,N_23049);
nand U25353 (N_25353,N_22792,N_21693);
and U25354 (N_25354,N_21184,N_22947);
xnor U25355 (N_25355,N_23676,N_22537);
xnor U25356 (N_25356,N_22223,N_24805);
and U25357 (N_25357,N_24439,N_23219);
and U25358 (N_25358,N_20739,N_21129);
and U25359 (N_25359,N_21194,N_20684);
xnor U25360 (N_25360,N_22165,N_23256);
or U25361 (N_25361,N_23287,N_22759);
and U25362 (N_25362,N_23581,N_20634);
xnor U25363 (N_25363,N_20031,N_23481);
nand U25364 (N_25364,N_20023,N_22708);
or U25365 (N_25365,N_24935,N_20620);
and U25366 (N_25366,N_23839,N_20837);
nand U25367 (N_25367,N_20204,N_23840);
xor U25368 (N_25368,N_23611,N_20751);
xor U25369 (N_25369,N_21950,N_21023);
nor U25370 (N_25370,N_22625,N_23196);
nand U25371 (N_25371,N_20602,N_21272);
nand U25372 (N_25372,N_24554,N_24519);
and U25373 (N_25373,N_23569,N_23722);
nand U25374 (N_25374,N_24696,N_23214);
and U25375 (N_25375,N_22134,N_20379);
or U25376 (N_25376,N_23264,N_23549);
or U25377 (N_25377,N_20719,N_24120);
nor U25378 (N_25378,N_23199,N_21695);
or U25379 (N_25379,N_20328,N_23458);
and U25380 (N_25380,N_22557,N_24150);
and U25381 (N_25381,N_21265,N_21080);
nor U25382 (N_25382,N_20175,N_23728);
nor U25383 (N_25383,N_21186,N_20320);
or U25384 (N_25384,N_24583,N_21359);
and U25385 (N_25385,N_24740,N_24955);
or U25386 (N_25386,N_20642,N_22071);
and U25387 (N_25387,N_24725,N_20295);
xor U25388 (N_25388,N_23504,N_21027);
or U25389 (N_25389,N_21185,N_23825);
and U25390 (N_25390,N_20639,N_22566);
and U25391 (N_25391,N_23150,N_24611);
xnor U25392 (N_25392,N_23241,N_24121);
or U25393 (N_25393,N_20370,N_20492);
and U25394 (N_25394,N_20523,N_24897);
nor U25395 (N_25395,N_24994,N_23208);
nand U25396 (N_25396,N_20516,N_20176);
and U25397 (N_25397,N_23552,N_20791);
nor U25398 (N_25398,N_20348,N_23117);
nand U25399 (N_25399,N_21960,N_21538);
and U25400 (N_25400,N_23618,N_23491);
or U25401 (N_25401,N_22449,N_21212);
and U25402 (N_25402,N_23706,N_24011);
nand U25403 (N_25403,N_22644,N_22913);
nand U25404 (N_25404,N_22532,N_23865);
or U25405 (N_25405,N_21168,N_20367);
and U25406 (N_25406,N_24012,N_20463);
and U25407 (N_25407,N_24349,N_21862);
nor U25408 (N_25408,N_24853,N_24336);
xor U25409 (N_25409,N_22734,N_22821);
nand U25410 (N_25410,N_21378,N_24906);
nand U25411 (N_25411,N_20960,N_20595);
and U25412 (N_25412,N_20435,N_20480);
nand U25413 (N_25413,N_21421,N_24956);
and U25414 (N_25414,N_22955,N_24596);
nand U25415 (N_25415,N_20363,N_23837);
nor U25416 (N_25416,N_22997,N_22408);
nor U25417 (N_25417,N_22139,N_23626);
and U25418 (N_25418,N_22098,N_24728);
xor U25419 (N_25419,N_21038,N_23048);
and U25420 (N_25420,N_21244,N_23443);
nand U25421 (N_25421,N_24094,N_23479);
nor U25422 (N_25422,N_22032,N_23904);
nand U25423 (N_25423,N_24954,N_23738);
or U25424 (N_25424,N_20105,N_20856);
xnor U25425 (N_25425,N_20776,N_21908);
nand U25426 (N_25426,N_24000,N_23766);
and U25427 (N_25427,N_23182,N_24480);
or U25428 (N_25428,N_20838,N_22155);
xor U25429 (N_25429,N_23793,N_20185);
nor U25430 (N_25430,N_21356,N_23402);
nand U25431 (N_25431,N_20654,N_22770);
xnor U25432 (N_25432,N_22697,N_22418);
nand U25433 (N_25433,N_20568,N_24328);
nor U25434 (N_25434,N_21264,N_24007);
nor U25435 (N_25435,N_22138,N_20037);
nand U25436 (N_25436,N_22674,N_22874);
or U25437 (N_25437,N_23811,N_21464);
nor U25438 (N_25438,N_22145,N_21477);
nand U25439 (N_25439,N_22221,N_22815);
or U25440 (N_25440,N_23078,N_21959);
nor U25441 (N_25441,N_24090,N_24777);
xor U25442 (N_25442,N_20730,N_21929);
xor U25443 (N_25443,N_23181,N_20345);
nor U25444 (N_25444,N_23957,N_20782);
and U25445 (N_25445,N_24952,N_21069);
nor U25446 (N_25446,N_22434,N_23721);
nand U25447 (N_25447,N_20225,N_24930);
and U25448 (N_25448,N_20640,N_24582);
and U25449 (N_25449,N_22174,N_24791);
or U25450 (N_25450,N_23400,N_22056);
and U25451 (N_25451,N_22554,N_24445);
nand U25452 (N_25452,N_24185,N_24139);
xor U25453 (N_25453,N_20901,N_24052);
or U25454 (N_25454,N_22838,N_24391);
nor U25455 (N_25455,N_22965,N_22161);
nor U25456 (N_25456,N_22877,N_21592);
or U25457 (N_25457,N_23791,N_23751);
nor U25458 (N_25458,N_24621,N_20417);
or U25459 (N_25459,N_21861,N_20643);
and U25460 (N_25460,N_23937,N_21674);
xor U25461 (N_25461,N_23232,N_24833);
nor U25462 (N_25462,N_22166,N_23542);
nand U25463 (N_25463,N_20557,N_23852);
nor U25464 (N_25464,N_24301,N_22261);
nand U25465 (N_25465,N_21722,N_23556);
nor U25466 (N_25466,N_21311,N_24039);
nor U25467 (N_25467,N_20508,N_22239);
or U25468 (N_25468,N_21004,N_20007);
and U25469 (N_25469,N_23105,N_22501);
or U25470 (N_25470,N_22930,N_22990);
nand U25471 (N_25471,N_23192,N_21029);
and U25472 (N_25472,N_23324,N_20150);
or U25473 (N_25473,N_24876,N_21541);
nand U25474 (N_25474,N_22167,N_21234);
nand U25475 (N_25475,N_23148,N_20932);
nand U25476 (N_25476,N_23065,N_22462);
or U25477 (N_25477,N_22159,N_20672);
or U25478 (N_25478,N_22676,N_22825);
nor U25479 (N_25479,N_24230,N_20115);
nor U25480 (N_25480,N_20762,N_23899);
or U25481 (N_25481,N_22443,N_24164);
and U25482 (N_25482,N_23386,N_21460);
or U25483 (N_25483,N_20584,N_21513);
and U25484 (N_25484,N_22731,N_23311);
or U25485 (N_25485,N_22547,N_22047);
nand U25486 (N_25486,N_22848,N_20069);
or U25487 (N_25487,N_23053,N_22923);
nand U25488 (N_25488,N_24253,N_24322);
nor U25489 (N_25489,N_20141,N_24477);
and U25490 (N_25490,N_22716,N_20866);
nor U25491 (N_25491,N_20586,N_20656);
and U25492 (N_25492,N_22576,N_20679);
and U25493 (N_25493,N_23525,N_21880);
and U25494 (N_25494,N_22819,N_20575);
nand U25495 (N_25495,N_20012,N_20548);
nand U25496 (N_25496,N_24632,N_24013);
xnor U25497 (N_25497,N_23750,N_24262);
or U25498 (N_25498,N_24631,N_22487);
or U25499 (N_25499,N_23804,N_21077);
nand U25500 (N_25500,N_22603,N_20552);
and U25501 (N_25501,N_23142,N_22667);
nor U25502 (N_25502,N_20453,N_23586);
and U25503 (N_25503,N_21821,N_24641);
and U25504 (N_25504,N_21229,N_23485);
or U25505 (N_25505,N_20438,N_22685);
and U25506 (N_25506,N_24623,N_21293);
nand U25507 (N_25507,N_23754,N_24064);
nand U25508 (N_25508,N_22347,N_21235);
nor U25509 (N_25509,N_21341,N_20613);
and U25510 (N_25510,N_22733,N_24318);
nor U25511 (N_25511,N_21984,N_21534);
xor U25512 (N_25512,N_21119,N_20008);
and U25513 (N_25513,N_24561,N_23223);
or U25514 (N_25514,N_22478,N_23913);
xor U25515 (N_25515,N_21987,N_21779);
or U25516 (N_25516,N_24510,N_22080);
nor U25517 (N_25517,N_21213,N_24637);
nand U25518 (N_25518,N_21780,N_24263);
and U25519 (N_25519,N_22414,N_21625);
xnor U25520 (N_25520,N_21058,N_20995);
and U25521 (N_25521,N_23724,N_23893);
and U25522 (N_25522,N_24995,N_20315);
and U25523 (N_25523,N_21888,N_20834);
xnor U25524 (N_25524,N_21917,N_21837);
nand U25525 (N_25525,N_20876,N_24724);
nand U25526 (N_25526,N_22875,N_21150);
and U25527 (N_25527,N_22768,N_20130);
or U25528 (N_25528,N_21686,N_21587);
xnor U25529 (N_25529,N_24929,N_24063);
nor U25530 (N_25530,N_24373,N_22710);
and U25531 (N_25531,N_22991,N_23709);
nand U25532 (N_25532,N_20374,N_24933);
xnor U25533 (N_25533,N_23652,N_20261);
nor U25534 (N_25534,N_22531,N_23130);
nand U25535 (N_25535,N_20341,N_20072);
xor U25536 (N_25536,N_24748,N_21367);
and U25537 (N_25537,N_21022,N_24503);
nand U25538 (N_25538,N_23010,N_23822);
and U25539 (N_25539,N_20999,N_21305);
or U25540 (N_25540,N_23894,N_23576);
and U25541 (N_25541,N_24872,N_22079);
and U25542 (N_25542,N_24457,N_22285);
nor U25543 (N_25543,N_21321,N_22057);
nand U25544 (N_25544,N_20849,N_22077);
nor U25545 (N_25545,N_21593,N_21444);
or U25546 (N_25546,N_22684,N_20519);
and U25547 (N_25547,N_24844,N_20038);
nand U25548 (N_25548,N_21009,N_24688);
nor U25549 (N_25549,N_22041,N_24355);
and U25550 (N_25550,N_24671,N_20870);
and U25551 (N_25551,N_21751,N_21761);
or U25552 (N_25552,N_20030,N_22290);
nor U25553 (N_25553,N_22827,N_23029);
nand U25554 (N_25554,N_24590,N_23092);
or U25555 (N_25555,N_20336,N_21939);
nand U25556 (N_25556,N_24616,N_22114);
nand U25557 (N_25557,N_24434,N_22448);
nor U25558 (N_25558,N_23397,N_22457);
nor U25559 (N_25559,N_23000,N_20985);
or U25560 (N_25560,N_24982,N_23342);
nor U25561 (N_25561,N_22381,N_24378);
xor U25562 (N_25562,N_21206,N_21784);
xnor U25563 (N_25563,N_20902,N_24123);
xor U25564 (N_25564,N_24615,N_22983);
and U25565 (N_25565,N_20820,N_20906);
nor U25566 (N_25566,N_23112,N_22104);
nand U25567 (N_25567,N_20833,N_23480);
and U25568 (N_25568,N_20166,N_22356);
nor U25569 (N_25569,N_23483,N_21756);
or U25570 (N_25570,N_22574,N_20612);
and U25571 (N_25571,N_20565,N_23395);
and U25572 (N_25572,N_20799,N_20836);
nor U25573 (N_25573,N_23033,N_23829);
nor U25574 (N_25574,N_22169,N_22471);
or U25575 (N_25575,N_22642,N_21585);
nand U25576 (N_25576,N_22225,N_23772);
nand U25577 (N_25577,N_20498,N_23905);
xor U25578 (N_25578,N_23590,N_24229);
and U25579 (N_25579,N_22973,N_24970);
xor U25580 (N_25580,N_23060,N_21914);
xnor U25581 (N_25581,N_23871,N_23943);
nand U25582 (N_25582,N_22592,N_20696);
or U25583 (N_25583,N_22982,N_21606);
xor U25584 (N_25584,N_21130,N_22435);
xnor U25585 (N_25585,N_21467,N_21313);
xor U25586 (N_25586,N_22704,N_21994);
xnor U25587 (N_25587,N_23281,N_20662);
nand U25588 (N_25588,N_23877,N_24951);
nor U25589 (N_25589,N_21364,N_20449);
nand U25590 (N_25590,N_23189,N_24241);
nand U25591 (N_25591,N_23369,N_24423);
xnor U25592 (N_25592,N_20892,N_24612);
and U25593 (N_25593,N_22550,N_24959);
or U25594 (N_25594,N_23164,N_22189);
nand U25595 (N_25595,N_22652,N_21512);
nand U25596 (N_25596,N_20222,N_24717);
nand U25597 (N_25597,N_21232,N_22502);
and U25598 (N_25598,N_21554,N_23757);
nand U25599 (N_25599,N_20440,N_22762);
nand U25600 (N_25600,N_24831,N_22197);
nand U25601 (N_25601,N_23606,N_23471);
and U25602 (N_25602,N_24205,N_24140);
xnor U25603 (N_25603,N_24086,N_20483);
xnor U25604 (N_25604,N_24404,N_22465);
and U25605 (N_25605,N_20073,N_21088);
or U25606 (N_25606,N_22267,N_24691);
and U25607 (N_25607,N_21291,N_21052);
or U25608 (N_25608,N_21754,N_23249);
or U25609 (N_25609,N_20061,N_20996);
or U25610 (N_25610,N_23140,N_20577);
nand U25611 (N_25611,N_20503,N_23050);
xnor U25612 (N_25612,N_23008,N_21930);
and U25613 (N_25613,N_22757,N_21724);
and U25614 (N_25614,N_21091,N_21471);
nor U25615 (N_25615,N_23303,N_23310);
nor U25616 (N_25616,N_21901,N_22939);
nand U25617 (N_25617,N_22096,N_21132);
nand U25618 (N_25618,N_23533,N_21651);
nor U25619 (N_25619,N_21708,N_23404);
nand U25620 (N_25620,N_21980,N_23396);
or U25621 (N_25621,N_20318,N_21308);
nand U25622 (N_25622,N_24027,N_20004);
nand U25623 (N_25623,N_20460,N_24051);
nor U25624 (N_25624,N_21996,N_23933);
xor U25625 (N_25625,N_24736,N_23305);
nor U25626 (N_25626,N_20145,N_21497);
xnor U25627 (N_25627,N_24282,N_23648);
xnor U25628 (N_25628,N_20447,N_20290);
or U25629 (N_25629,N_22772,N_21563);
and U25630 (N_25630,N_21816,N_21772);
nand U25631 (N_25631,N_24079,N_21963);
nor U25632 (N_25632,N_21909,N_22726);
and U25633 (N_25633,N_24259,N_21739);
nand U25634 (N_25634,N_21666,N_24679);
xnor U25635 (N_25635,N_20459,N_23884);
and U25636 (N_25636,N_22707,N_22403);
and U25637 (N_25637,N_20525,N_22953);
and U25638 (N_25638,N_20349,N_20221);
xor U25639 (N_25639,N_20967,N_24198);
xor U25640 (N_25640,N_23221,N_23614);
and U25641 (N_25641,N_20478,N_23908);
xor U25642 (N_25642,N_24531,N_24739);
or U25643 (N_25643,N_24682,N_22445);
and U25644 (N_25644,N_20000,N_21528);
xor U25645 (N_25645,N_22088,N_22633);
and U25646 (N_25646,N_24776,N_23284);
or U25647 (N_25647,N_20202,N_22037);
or U25648 (N_25648,N_22820,N_22467);
nor U25649 (N_25649,N_21903,N_24097);
nor U25650 (N_25650,N_22561,N_24115);
or U25651 (N_25651,N_20265,N_24437);
nand U25652 (N_25652,N_22000,N_23815);
nor U25653 (N_25653,N_21634,N_20758);
xnor U25654 (N_25654,N_22563,N_23263);
nand U25655 (N_25655,N_24544,N_20800);
xnor U25656 (N_25656,N_20993,N_24838);
or U25657 (N_25657,N_21720,N_22753);
xor U25658 (N_25658,N_20941,N_23995);
or U25659 (N_25659,N_24525,N_22312);
or U25660 (N_25660,N_22607,N_22120);
nor U25661 (N_25661,N_22583,N_24002);
nor U25662 (N_25662,N_23465,N_23500);
xor U25663 (N_25663,N_20542,N_24672);
or U25664 (N_25664,N_22438,N_20626);
nor U25665 (N_25665,N_22175,N_20864);
nor U25666 (N_25666,N_21360,N_22775);
xnor U25667 (N_25667,N_23202,N_24474);
and U25668 (N_25668,N_23780,N_20081);
or U25669 (N_25669,N_20916,N_21936);
nor U25670 (N_25670,N_24789,N_23497);
nand U25671 (N_25671,N_24977,N_23630);
nand U25672 (N_25672,N_23945,N_24347);
and U25673 (N_25673,N_22579,N_24861);
nor U25674 (N_25674,N_20452,N_23414);
xnor U25675 (N_25675,N_23797,N_24415);
nand U25676 (N_25676,N_20238,N_20631);
nor U25677 (N_25677,N_21210,N_20041);
nand U25678 (N_25678,N_21559,N_20183);
xor U25679 (N_25679,N_21866,N_23792);
or U25680 (N_25680,N_21840,N_23662);
nor U25681 (N_25681,N_22809,N_24708);
nor U25682 (N_25682,N_21652,N_21894);
xnor U25683 (N_25683,N_24223,N_23329);
xnor U25684 (N_25684,N_22689,N_21351);
xor U25685 (N_25685,N_20323,N_21690);
nand U25686 (N_25686,N_21726,N_24288);
nor U25687 (N_25687,N_21581,N_22709);
xor U25688 (N_25688,N_21961,N_23306);
nand U25689 (N_25689,N_20107,N_24571);
and U25690 (N_25690,N_24233,N_24598);
or U25691 (N_25691,N_23858,N_23895);
nor U25692 (N_25692,N_23873,N_22692);
nor U25693 (N_25693,N_20583,N_21398);
and U25694 (N_25694,N_21024,N_23548);
or U25695 (N_25695,N_22626,N_24639);
xor U25696 (N_25696,N_24668,N_21394);
nand U25697 (N_25697,N_21352,N_21545);
xnor U25698 (N_25698,N_22837,N_23613);
and U25699 (N_25699,N_22317,N_21520);
xnor U25700 (N_25700,N_20829,N_23968);
or U25701 (N_25701,N_24343,N_23367);
nand U25702 (N_25702,N_20300,N_24181);
nor U25703 (N_25703,N_21228,N_22956);
xor U25704 (N_25704,N_21925,N_20644);
xnor U25705 (N_25705,N_24279,N_21907);
or U25706 (N_25706,N_23950,N_24785);
and U25707 (N_25707,N_22556,N_24483);
xnor U25708 (N_25708,N_23445,N_20104);
xnor U25709 (N_25709,N_22427,N_20690);
nand U25710 (N_25710,N_24543,N_21502);
nor U25711 (N_25711,N_24031,N_22785);
nand U25712 (N_25712,N_20729,N_20990);
nand U25713 (N_25713,N_20247,N_23109);
or U25714 (N_25714,N_22912,N_23007);
and U25715 (N_25715,N_20790,N_20842);
xnor U25716 (N_25716,N_22413,N_21049);
nor U25717 (N_25717,N_20887,N_21619);
nand U25718 (N_25718,N_24836,N_21096);
nand U25719 (N_25719,N_21848,N_22823);
and U25720 (N_25720,N_23519,N_23949);
nor U25721 (N_25721,N_20102,N_22952);
and U25722 (N_25722,N_21276,N_22859);
nor U25723 (N_25723,N_22524,N_22007);
nor U25724 (N_25724,N_22379,N_22406);
or U25725 (N_25725,N_20925,N_21452);
xor U25726 (N_25726,N_21219,N_20827);
xnor U25727 (N_25727,N_23068,N_20727);
and U25728 (N_25728,N_20668,N_22348);
nand U25729 (N_25729,N_20968,N_21299);
or U25730 (N_25730,N_21696,N_20118);
xnor U25731 (N_25731,N_24005,N_22276);
nand U25732 (N_25732,N_22089,N_23157);
nor U25733 (N_25733,N_20873,N_23175);
and U25734 (N_25734,N_24798,N_24431);
nor U25735 (N_25735,N_20294,N_21525);
xnor U25736 (N_25736,N_21588,N_20354);
nor U25737 (N_25737,N_21773,N_22108);
and U25738 (N_25738,N_23786,N_22255);
or U25739 (N_25739,N_23687,N_22234);
nand U25740 (N_25740,N_21396,N_20182);
and U25741 (N_25741,N_23777,N_24712);
xor U25742 (N_25742,N_24680,N_23169);
or U25743 (N_25743,N_23017,N_20844);
nand U25744 (N_25744,N_23629,N_23201);
nand U25745 (N_25745,N_20784,N_20585);
xnor U25746 (N_25746,N_24878,N_23222);
and U25747 (N_25747,N_22729,N_24647);
and U25748 (N_25748,N_21328,N_23063);
xor U25749 (N_25749,N_23238,N_23730);
nor U25750 (N_25750,N_24662,N_20019);
nor U25751 (N_25751,N_24206,N_24119);
and U25752 (N_25752,N_24350,N_20549);
and U25753 (N_25753,N_24329,N_22295);
and U25754 (N_25754,N_23089,N_23589);
or U25755 (N_25755,N_20063,N_24673);
nand U25756 (N_25756,N_21638,N_23312);
or U25757 (N_25757,N_23919,N_22451);
or U25758 (N_25758,N_20214,N_21067);
nor U25759 (N_25759,N_23315,N_23354);
and U25760 (N_25760,N_24742,N_21685);
or U25761 (N_25761,N_22473,N_22570);
nor U25762 (N_25762,N_22474,N_24314);
or U25763 (N_25763,N_22962,N_20251);
nor U25764 (N_25764,N_23512,N_23041);
nor U25765 (N_25765,N_24407,N_20456);
nor U25766 (N_25766,N_23992,N_23900);
or U25767 (N_25767,N_21297,N_20032);
nand U25768 (N_25768,N_22647,N_20423);
nand U25769 (N_25769,N_22195,N_24594);
xnor U25770 (N_25770,N_23932,N_23690);
and U25771 (N_25771,N_20882,N_23947);
or U25772 (N_25772,N_24790,N_24961);
and U25773 (N_25773,N_20649,N_22141);
nand U25774 (N_25774,N_23719,N_24441);
and U25775 (N_25775,N_22078,N_20988);
or U25776 (N_25776,N_21331,N_22858);
nand U25777 (N_25777,N_22853,N_24089);
or U25778 (N_25778,N_21262,N_21557);
xnor U25779 (N_25779,N_22536,N_21068);
nand U25780 (N_25780,N_21493,N_24697);
nor U25781 (N_25781,N_21140,N_22357);
xor U25782 (N_25782,N_23013,N_22472);
xnor U25783 (N_25783,N_21036,N_23082);
nand U25784 (N_25784,N_21145,N_20448);
or U25785 (N_25785,N_20236,N_24360);
xor U25786 (N_25786,N_23683,N_20119);
or U25787 (N_25787,N_23444,N_22968);
and U25788 (N_25788,N_24444,N_23901);
and U25789 (N_25789,N_20289,N_22420);
and U25790 (N_25790,N_21522,N_21982);
nor U25791 (N_25791,N_24516,N_24532);
nand U25792 (N_25792,N_20871,N_23638);
xor U25793 (N_25793,N_21834,N_21115);
nor U25794 (N_25794,N_24417,N_24996);
nor U25795 (N_25795,N_22363,N_23866);
or U25796 (N_25796,N_20770,N_22130);
and U25797 (N_25797,N_21161,N_23149);
xnor U25798 (N_25798,N_20457,N_20616);
or U25799 (N_25799,N_22680,N_23986);
and U25800 (N_25800,N_20223,N_20702);
and U25801 (N_25801,N_23376,N_20989);
xor U25802 (N_25802,N_24071,N_24689);
or U25803 (N_25803,N_21492,N_23331);
and U25804 (N_25804,N_22959,N_22538);
nor U25805 (N_25805,N_20918,N_21260);
nor U25806 (N_25806,N_20997,N_21047);
nand U25807 (N_25807,N_24772,N_20614);
nand U25808 (N_25808,N_21702,N_20006);
or U25809 (N_25809,N_21723,N_22807);
or U25810 (N_25810,N_20926,N_24627);
nand U25811 (N_25811,N_21334,N_24699);
and U25812 (N_25812,N_23285,N_24473);
and U25813 (N_25813,N_21007,N_21531);
and U25814 (N_25814,N_23015,N_22458);
and U25815 (N_25815,N_24442,N_24193);
and U25816 (N_25816,N_22422,N_24852);
or U25817 (N_25817,N_20897,N_23416);
or U25818 (N_25818,N_24156,N_24158);
nand U25819 (N_25819,N_23511,N_24315);
nor U25820 (N_25820,N_23036,N_23610);
nor U25821 (N_25821,N_23350,N_22398);
xor U25822 (N_25822,N_24055,N_20256);
nor U25823 (N_25823,N_24950,N_23023);
or U25824 (N_25824,N_22934,N_24869);
nor U25825 (N_25825,N_20629,N_23966);
or U25826 (N_25826,N_23253,N_22084);
and U25827 (N_25827,N_24324,N_24868);
nor U25828 (N_25828,N_21179,N_20658);
xnor U25829 (N_25829,N_20050,N_20740);
nor U25830 (N_25830,N_24232,N_24920);
nor U25831 (N_25831,N_20930,N_20957);
nand U25832 (N_25832,N_23093,N_21819);
xor U25833 (N_25833,N_21361,N_22567);
or U25834 (N_25834,N_23213,N_24147);
nor U25835 (N_25835,N_22596,N_24487);
nor U25836 (N_25836,N_24840,N_21268);
and U25837 (N_25837,N_24536,N_24726);
or U25838 (N_25838,N_20197,N_21556);
or U25839 (N_25839,N_24409,N_23897);
or U25840 (N_25840,N_24362,N_21700);
xnor U25841 (N_25841,N_23924,N_23915);
nor U25842 (N_25842,N_23427,N_20412);
xnor U25843 (N_25843,N_23670,N_23432);
nand U25844 (N_25844,N_20433,N_22814);
or U25845 (N_25845,N_20302,N_22711);
nor U25846 (N_25846,N_21876,N_24286);
nand U25847 (N_25847,N_22872,N_20853);
or U25848 (N_25848,N_20392,N_21620);
or U25849 (N_25849,N_23753,N_23747);
nand U25850 (N_25850,N_24481,N_22584);
xnor U25851 (N_25851,N_22012,N_24023);
nand U25852 (N_25852,N_24514,N_20172);
or U25853 (N_25853,N_20589,N_22146);
nand U25854 (N_25854,N_24069,N_20766);
xnor U25855 (N_25855,N_23259,N_21659);
nand U25856 (N_25856,N_21434,N_23289);
or U25857 (N_25857,N_21082,N_21614);
xor U25858 (N_25858,N_20490,N_24709);
nand U25859 (N_25859,N_23679,N_23431);
nand U25860 (N_25860,N_20905,N_24368);
nand U25861 (N_25861,N_20811,N_21459);
nor U25862 (N_25862,N_21515,N_22849);
and U25863 (N_25863,N_23236,N_20134);
xor U25864 (N_25864,N_20036,N_24614);
xor U25865 (N_25865,N_22941,N_24352);
or U25866 (N_25866,N_22643,N_24281);
xnor U25867 (N_25867,N_21247,N_24522);
xor U25868 (N_25868,N_24706,N_24215);
nor U25869 (N_25869,N_20725,N_22812);
nor U25870 (N_25870,N_24166,N_23756);
nand U25871 (N_25871,N_21711,N_21318);
or U25872 (N_25872,N_23011,N_23846);
nor U25873 (N_25873,N_21169,N_20406);
nor U25874 (N_25874,N_21170,N_24862);
xnor U25875 (N_25875,N_20588,N_23269);
xnor U25876 (N_25876,N_21787,N_21918);
nor U25877 (N_25877,N_24105,N_20254);
nand U25878 (N_25878,N_21879,N_22627);
and U25879 (N_25879,N_20694,N_21615);
xor U25880 (N_25880,N_22549,N_21575);
and U25881 (N_25881,N_23333,N_22789);
or U25882 (N_25882,N_21817,N_20518);
or U25883 (N_25883,N_24928,N_21978);
xor U25884 (N_25884,N_22826,N_20522);
or U25885 (N_25885,N_23424,N_22998);
or U25886 (N_25886,N_22183,N_23642);
nand U25887 (N_25887,N_21040,N_22046);
nor U25888 (N_25888,N_21037,N_24979);
nor U25889 (N_25889,N_21301,N_23812);
xor U25890 (N_25890,N_24413,N_23336);
xor U25891 (N_25891,N_24176,N_24850);
nand U25892 (N_25892,N_22740,N_22464);
xor U25893 (N_25893,N_23861,N_20801);
xor U25894 (N_25894,N_20628,N_20270);
nor U25895 (N_25895,N_22824,N_21688);
and U25896 (N_25896,N_22091,N_23659);
and U25897 (N_25897,N_24932,N_21968);
and U25898 (N_25898,N_22216,N_22829);
or U25899 (N_25899,N_24983,N_22954);
xor U25900 (N_25900,N_24660,N_22342);
nor U25901 (N_25901,N_22140,N_23917);
and U25902 (N_25902,N_23523,N_22958);
xor U25903 (N_25903,N_23052,N_21383);
or U25904 (N_25904,N_24884,N_20755);
or U25905 (N_25905,N_22992,N_24524);
and U25906 (N_25906,N_21086,N_24997);
nor U25907 (N_25907,N_23823,N_20299);
and U25908 (N_25908,N_20580,N_24219);
nor U25909 (N_25909,N_20715,N_24702);
and U25910 (N_25910,N_21752,N_20599);
nand U25911 (N_25911,N_24658,N_20975);
nand U25912 (N_25912,N_21973,N_20560);
xnor U25913 (N_25913,N_22214,N_20721);
nor U25914 (N_25914,N_21967,N_20622);
and U25915 (N_25915,N_23300,N_21373);
and U25916 (N_25916,N_24867,N_22610);
and U25917 (N_25917,N_21261,N_21859);
nand U25918 (N_25918,N_20413,N_23807);
or U25919 (N_25919,N_24520,N_20535);
nor U25920 (N_25920,N_21354,N_20826);
and U25921 (N_25921,N_20603,N_21571);
xnor U25922 (N_25922,N_22278,N_21586);
or U25923 (N_25923,N_24609,N_20409);
nor U25924 (N_25924,N_23674,N_24856);
xnor U25925 (N_25925,N_23844,N_24388);
nor U25926 (N_25926,N_20623,N_24779);
xnor U25927 (N_25927,N_21060,N_21072);
or U25928 (N_25928,N_22778,N_22703);
xnor U25929 (N_25929,N_24313,N_21750);
or U25930 (N_25930,N_20958,N_20437);
and U25931 (N_25931,N_20952,N_23026);
nor U25932 (N_25932,N_23802,N_21409);
and U25933 (N_25933,N_22335,N_20329);
or U25934 (N_25934,N_22326,N_23270);
and U25935 (N_25935,N_20342,N_20537);
nand U25936 (N_25936,N_21796,N_21671);
and U25937 (N_25937,N_22925,N_20899);
nor U25938 (N_25938,N_20732,N_24317);
xor U25939 (N_25939,N_21094,N_24085);
and U25940 (N_25940,N_20778,N_20499);
or U25941 (N_25941,N_22005,N_22700);
nand U25942 (N_25942,N_24062,N_21898);
and U25943 (N_25943,N_24877,N_23848);
nand U25944 (N_25944,N_22743,N_23868);
nor U25945 (N_25945,N_21957,N_20529);
or U25946 (N_25946,N_22156,N_24894);
or U25947 (N_25947,N_20312,N_24136);
xnor U25948 (N_25948,N_24547,N_22226);
and U25949 (N_25949,N_20567,N_24070);
xnor U25950 (N_25950,N_24828,N_21484);
nand U25951 (N_25951,N_24550,N_23454);
nand U25952 (N_25952,N_23360,N_21504);
xnor U25953 (N_25953,N_20292,N_24184);
or U25954 (N_25954,N_22333,N_20291);
nand U25955 (N_25955,N_23579,N_22050);
xor U25956 (N_25956,N_21633,N_23566);
nor U25957 (N_25957,N_23686,N_23983);
and U25958 (N_25958,N_22417,N_21947);
or U25959 (N_25959,N_20604,N_22589);
or U25960 (N_25960,N_21738,N_22660);
xor U25961 (N_25961,N_20579,N_21197);
nor U25962 (N_25962,N_24226,N_20600);
xor U25963 (N_25963,N_22620,N_24542);
xor U25964 (N_25964,N_21034,N_24704);
and U25965 (N_25965,N_22788,N_20666);
nor U25966 (N_25966,N_20128,N_21637);
nor U25967 (N_25967,N_22201,N_22803);
nor U25968 (N_25968,N_24624,N_23898);
and U25969 (N_25969,N_22860,N_21043);
nor U25970 (N_25970,N_20886,N_20652);
and U25971 (N_25971,N_21441,N_24591);
xnor U25972 (N_25972,N_23209,N_20804);
xnor U25973 (N_25973,N_20507,N_23472);
and U25974 (N_25974,N_21551,N_20158);
and U25975 (N_25975,N_20099,N_22097);
or U25976 (N_25976,N_23737,N_24234);
or U25977 (N_25977,N_21209,N_20706);
nand U25978 (N_25978,N_21236,N_21306);
nor U25979 (N_25979,N_23831,N_23032);
nor U25980 (N_25980,N_21860,N_21863);
and U25981 (N_25981,N_24399,N_21568);
nor U25982 (N_25982,N_22769,N_24306);
nand U25983 (N_25983,N_21355,N_21137);
nor U25984 (N_25984,N_21374,N_23215);
and U25985 (N_25985,N_23964,N_23712);
nand U25986 (N_25986,N_22222,N_22188);
or U25987 (N_25987,N_22305,N_22987);
and U25988 (N_25988,N_23628,N_22903);
or U25989 (N_25989,N_21160,N_23517);
nand U25990 (N_25990,N_20120,N_21455);
and U25991 (N_25991,N_22739,N_20900);
or U25992 (N_25992,N_21475,N_20186);
and U25993 (N_25993,N_20720,N_23651);
nor U25994 (N_25994,N_22695,N_22758);
and U25995 (N_25995,N_20874,N_24964);
xor U25996 (N_25996,N_23851,N_24258);
and U25997 (N_25997,N_20981,N_24009);
or U25998 (N_25998,N_22025,N_20881);
nor U25999 (N_25999,N_20124,N_23699);
or U26000 (N_26000,N_20688,N_21802);
nor U26001 (N_26001,N_20364,N_24196);
nor U26002 (N_26002,N_23225,N_21430);
nor U26003 (N_26003,N_23325,N_21524);
or U26004 (N_26004,N_21174,N_24613);
nor U26005 (N_26005,N_20551,N_24112);
nand U26006 (N_26006,N_20297,N_24386);
and U26007 (N_26007,N_22419,N_24568);
xnor U26008 (N_26008,N_20053,N_21343);
xnor U26009 (N_26009,N_23773,N_21010);
nand U26010 (N_26010,N_20213,N_21897);
or U26011 (N_26011,N_24521,N_24567);
nor U26012 (N_26012,N_22539,N_24812);
xnor U26013 (N_26013,N_22588,N_23695);
nor U26014 (N_26014,N_21923,N_23768);
and U26015 (N_26015,N_24138,N_21118);
nand U26016 (N_26016,N_21348,N_23132);
nor U26017 (N_26017,N_24298,N_24905);
nor U26018 (N_26018,N_24529,N_22855);
nand U26019 (N_26019,N_21993,N_24114);
nor U26020 (N_26020,N_20942,N_22442);
nor U26021 (N_26021,N_24499,N_20333);
nand U26022 (N_26022,N_24958,N_22309);
nor U26023 (N_26023,N_21687,N_22523);
xor U26024 (N_26024,N_22250,N_21875);
nor U26025 (N_26025,N_21835,N_21400);
or U26026 (N_26026,N_20722,N_23280);
nand U26027 (N_26027,N_21494,N_24491);
or U26028 (N_26028,N_20563,N_20816);
and U26029 (N_26029,N_24578,N_24498);
nand U26030 (N_26030,N_22617,N_22517);
and U26031 (N_26031,N_23463,N_24186);
xnor U26032 (N_26032,N_24128,N_21405);
nand U26033 (N_26033,N_22070,N_22715);
and U26034 (N_26034,N_20168,N_21790);
nor U26035 (N_26035,N_22892,N_23363);
nor U26036 (N_26036,N_22127,N_23969);
xor U26037 (N_26037,N_21869,N_20268);
or U26038 (N_26038,N_20780,N_24141);
nand U26039 (N_26039,N_22624,N_20296);
or U26040 (N_26040,N_21946,N_24541);
nor U26041 (N_26041,N_22582,N_20093);
and U26042 (N_26042,N_22439,N_21439);
nor U26043 (N_26043,N_22777,N_20086);
or U26044 (N_26044,N_21281,N_24546);
xnor U26045 (N_26045,N_21246,N_23294);
nor U26046 (N_26046,N_20819,N_21727);
nor U26047 (N_26047,N_21795,N_21844);
nor U26048 (N_26048,N_24968,N_22996);
nor U26049 (N_26049,N_22042,N_21839);
nand U26050 (N_26050,N_22608,N_21144);
or U26051 (N_26051,N_21622,N_21440);
or U26052 (N_26052,N_20909,N_21192);
nand U26053 (N_26053,N_24901,N_24559);
and U26054 (N_26054,N_20464,N_24354);
xor U26055 (N_26055,N_23061,N_20486);
or U26056 (N_26056,N_23931,N_24045);
and U26057 (N_26057,N_21558,N_23307);
xnor U26058 (N_26058,N_23279,N_24244);
or U26059 (N_26059,N_23952,N_20689);
or U26060 (N_26060,N_22901,N_24584);
nand U26061 (N_26061,N_24365,N_22651);
or U26062 (N_26062,N_20550,N_21326);
or U26063 (N_26063,N_22665,N_24191);
or U26064 (N_26064,N_23334,N_21158);
xor U26065 (N_26065,N_21797,N_24267);
xnor U26066 (N_26066,N_23459,N_21616);
xnor U26067 (N_26067,N_22274,N_20590);
and U26068 (N_26068,N_24425,N_20880);
nor U26069 (N_26069,N_23520,N_24163);
or U26070 (N_26070,N_23887,N_24610);
or U26071 (N_26071,N_23038,N_21288);
nor U26072 (N_26072,N_20042,N_23954);
and U26073 (N_26073,N_23492,N_20350);
nand U26074 (N_26074,N_20232,N_23857);
nand U26075 (N_26075,N_24394,N_24339);
nand U26076 (N_26076,N_24227,N_20461);
and U26077 (N_26077,N_24657,N_21926);
or U26078 (N_26078,N_22252,N_23981);
or U26079 (N_26079,N_23004,N_23530);
nand U26080 (N_26080,N_23600,N_22794);
nand U26081 (N_26081,N_22202,N_21506);
nor U26082 (N_26082,N_22318,N_23428);
xnor U26083 (N_26083,N_21691,N_20258);
nand U26084 (N_26084,N_20301,N_24973);
nand U26085 (N_26085,N_20998,N_21496);
nor U26086 (N_26086,N_24303,N_22602);
nand U26087 (N_26087,N_22254,N_21827);
nand U26088 (N_26088,N_22286,N_21454);
xnor U26089 (N_26089,N_22373,N_21657);
or U26090 (N_26090,N_20582,N_23173);
nor U26091 (N_26091,N_22525,N_22215);
or U26092 (N_26092,N_21487,N_23455);
nor U26093 (N_26093,N_21874,N_24644);
or U26094 (N_26094,N_20777,N_23081);
nand U26095 (N_26095,N_20101,N_20255);
and U26096 (N_26096,N_21649,N_21740);
and U26097 (N_26097,N_23216,N_24342);
nand U26098 (N_26098,N_21388,N_24490);
nand U26099 (N_26099,N_24693,N_23608);
or U26100 (N_26100,N_22797,N_20959);
and U26101 (N_26101,N_23392,N_20429);
xnor U26102 (N_26102,N_21333,N_20330);
nor U26103 (N_26103,N_24122,N_20504);
nand U26104 (N_26104,N_24034,N_20127);
or U26105 (N_26105,N_21384,N_20153);
and U26106 (N_26106,N_23170,N_24835);
or U26107 (N_26107,N_23298,N_22974);
xor U26108 (N_26108,N_24767,N_21491);
or U26109 (N_26109,N_20847,N_20966);
nor U26110 (N_26110,N_24981,N_21741);
or U26111 (N_26111,N_23299,N_23572);
xor U26112 (N_26112,N_22897,N_20143);
xor U26113 (N_26113,N_23425,N_21231);
nand U26114 (N_26114,N_24826,N_22970);
and U26115 (N_26115,N_22362,N_21856);
and U26116 (N_26116,N_24971,N_20467);
xnor U26117 (N_26117,N_21857,N_23075);
xor U26118 (N_26118,N_23658,N_22376);
nor U26119 (N_26119,N_24752,N_20933);
nand U26120 (N_26120,N_20123,N_22663);
nand U26121 (N_26121,N_23923,N_24871);
and U26122 (N_26122,N_20025,N_23104);
nand U26123 (N_26123,N_22801,N_24945);
nor U26124 (N_26124,N_20638,N_23599);
xnor U26125 (N_26125,N_20520,N_24762);
nand U26126 (N_26126,N_24296,N_20114);
or U26127 (N_26127,N_21056,N_21777);
nor U26128 (N_26128,N_23365,N_24161);
or U26129 (N_26129,N_20677,N_20814);
or U26130 (N_26130,N_20088,N_20377);
or U26131 (N_26131,N_21878,N_20632);
nand U26132 (N_26132,N_23046,N_23850);
xor U26133 (N_26133,N_24099,N_21366);
and U26134 (N_26134,N_21259,N_24769);
nor U26135 (N_26135,N_23559,N_21309);
nor U26136 (N_26136,N_24414,N_20678);
nor U26137 (N_26137,N_23340,N_21851);
nand U26138 (N_26138,N_24539,N_21805);
and U26139 (N_26139,N_21566,N_23174);
or U26140 (N_26140,N_22518,N_24486);
nand U26141 (N_26141,N_20226,N_20227);
or U26142 (N_26142,N_23817,N_23563);
and U26143 (N_26143,N_21650,N_22945);
and U26144 (N_26144,N_22905,N_21589);
xnor U26145 (N_26145,N_21503,N_22771);
and U26146 (N_26146,N_22980,N_21548);
nor U26147 (N_26147,N_23226,N_24050);
and U26148 (N_26148,N_22375,N_24889);
nor U26149 (N_26149,N_20284,N_22401);
or U26150 (N_26150,N_23024,N_24987);
xor U26151 (N_26151,N_22720,N_22677);
nor U26152 (N_26152,N_20240,N_23680);
xnor U26153 (N_26153,N_22755,N_23135);
and U26154 (N_26154,N_23107,N_20726);
nand U26155 (N_26155,N_24482,N_20458);
and U26156 (N_26156,N_24435,N_23358);
nor U26157 (N_26157,N_23477,N_21415);
nand U26158 (N_26158,N_24814,N_24842);
or U26159 (N_26159,N_21516,N_23818);
and U26160 (N_26160,N_22928,N_24361);
nor U26161 (N_26161,N_24786,N_20380);
nor U26162 (N_26162,N_21386,N_21041);
or U26163 (N_26163,N_23534,N_23094);
xor U26164 (N_26164,N_23636,N_22943);
nor U26165 (N_26165,N_24299,N_23609);
xnor U26166 (N_26166,N_20391,N_24272);
xor U26167 (N_26167,N_24325,N_24302);
nor U26168 (N_26168,N_22149,N_21099);
nor U26169 (N_26169,N_24750,N_21087);
or U26170 (N_26170,N_24618,N_21853);
or U26171 (N_26171,N_21542,N_23025);
nand U26172 (N_26172,N_21178,N_24919);
and U26173 (N_26173,N_20868,N_23129);
and U26174 (N_26174,N_22259,N_22245);
and U26175 (N_26175,N_20015,N_21269);
and U26176 (N_26176,N_24081,N_24537);
nor U26177 (N_26177,N_24666,N_24066);
nor U26178 (N_26178,N_22323,N_22111);
and U26179 (N_26179,N_21793,N_23806);
nor U26180 (N_26180,N_24321,N_24564);
nand U26181 (N_26181,N_22179,N_21215);
or U26182 (N_26182,N_20136,N_21017);
nand U26183 (N_26183,N_24291,N_24058);
nor U26184 (N_26184,N_21138,N_22485);
and U26185 (N_26185,N_24903,N_20536);
nand U26186 (N_26186,N_22763,N_21838);
and U26187 (N_26187,N_22178,N_21141);
nand U26188 (N_26188,N_21882,N_23193);
and U26189 (N_26189,N_24479,N_21891);
or U26190 (N_26190,N_24730,N_21372);
nand U26191 (N_26191,N_23555,N_21177);
nor U26192 (N_26192,N_21465,N_23540);
xnor U26193 (N_26193,N_24562,N_21561);
and U26194 (N_26194,N_24635,N_21843);
and U26195 (N_26195,N_23383,N_23714);
nor U26196 (N_26196,N_20442,N_23946);
xnor U26197 (N_26197,N_21403,N_21937);
nor U26198 (N_26198,N_21715,N_20734);
xor U26199 (N_26199,N_22241,N_24412);
or U26200 (N_26200,N_20737,N_24029);
xnor U26201 (N_26201,N_21482,N_23975);
nand U26202 (N_26202,N_22116,N_22388);
nor U26203 (N_26203,N_23286,N_22450);
xor U26204 (N_26204,N_23058,N_21573);
nor U26205 (N_26205,N_22854,N_22719);
nand U26206 (N_26206,N_20547,N_20500);
nor U26207 (N_26207,N_22655,N_24100);
and U26208 (N_26208,N_21433,N_23824);
nand U26209 (N_26209,N_23230,N_21608);
nor U26210 (N_26210,N_22756,N_22993);
or U26211 (N_26211,N_21021,N_20337);
xnor U26212 (N_26212,N_20748,N_23028);
nand U26213 (N_26213,N_23778,N_21329);
or U26214 (N_26214,N_23816,N_23921);
xnor U26215 (N_26215,N_24751,N_21042);
or U26216 (N_26216,N_24940,N_20205);
and U26217 (N_26217,N_20151,N_22490);
or U26218 (N_26218,N_23095,N_23180);
and U26219 (N_26219,N_23009,N_22340);
and U26220 (N_26220,N_21488,N_23362);
and U26221 (N_26221,N_21684,N_22851);
nor U26222 (N_26222,N_24209,N_24581);
nor U26223 (N_26223,N_21799,N_20964);
nand U26224 (N_26224,N_20497,N_23388);
xnor U26225 (N_26225,N_22106,N_24863);
nor U26226 (N_26226,N_21498,N_23347);
xnor U26227 (N_26227,N_22425,N_20133);
and U26228 (N_26228,N_23565,N_24383);
nor U26229 (N_26229,N_20855,N_24924);
nor U26230 (N_26230,N_23688,N_20428);
nor U26231 (N_26231,N_24038,N_24896);
and U26232 (N_26232,N_22830,N_23604);
xnor U26233 (N_26233,N_24684,N_20249);
or U26234 (N_26234,N_22891,N_22981);
nor U26235 (N_26235,N_21451,N_24893);
or U26236 (N_26236,N_23407,N_22867);
nor U26237 (N_26237,N_24133,N_22343);
or U26238 (N_26238,N_22039,N_23819);
or U26239 (N_26239,N_22541,N_20951);
and U26240 (N_26240,N_22527,N_23484);
xnor U26241 (N_26241,N_23538,N_22888);
and U26242 (N_26242,N_21292,N_23607);
nand U26243 (N_26243,N_23255,N_20533);
or U26244 (N_26244,N_22618,N_22534);
xor U26245 (N_26245,N_21867,N_21537);
or U26246 (N_26246,N_22847,N_20961);
nor U26247 (N_26247,N_24649,N_23390);
nor U26248 (N_26248,N_21402,N_23508);
nand U26249 (N_26249,N_23744,N_24707);
and U26250 (N_26250,N_20470,N_23627);
and U26251 (N_26251,N_22142,N_21964);
nand U26252 (N_26252,N_20956,N_23641);
and U26253 (N_26253,N_22590,N_23152);
and U26254 (N_26254,N_23195,N_21273);
nand U26255 (N_26255,N_20576,N_23242);
nor U26256 (N_26256,N_21549,N_21518);
nor U26257 (N_26257,N_21147,N_20340);
nand U26258 (N_26258,N_23617,N_22940);
xor U26259 (N_26259,N_22074,N_24257);
or U26260 (N_26260,N_20002,N_23457);
or U26261 (N_26261,N_20872,N_24057);
and U26262 (N_26262,N_22275,N_21054);
and U26263 (N_26263,N_24986,N_23277);
and U26264 (N_26264,N_20733,N_22645);
nor U26265 (N_26265,N_21417,N_20891);
nor U26266 (N_26266,N_20048,N_23217);
xor U26267 (N_26267,N_24001,N_20910);
or U26268 (N_26268,N_23495,N_23955);
or U26269 (N_26269,N_23302,N_23022);
nor U26270 (N_26270,N_24892,N_22718);
and U26271 (N_26271,N_24026,N_20382);
xnor U26272 (N_26272,N_22736,N_23474);
nor U26273 (N_26273,N_21610,N_24822);
nand U26274 (N_26274,N_23870,N_20029);
nand U26275 (N_26275,N_20083,N_23501);
nor U26276 (N_26276,N_22144,N_21414);
xnor U26277 (N_26277,N_22122,N_22247);
nor U26278 (N_26278,N_21966,N_20344);
or U26279 (N_26279,N_23119,N_24687);
and U26280 (N_26280,N_20234,N_20669);
and U26281 (N_26281,N_21716,N_21788);
nor U26282 (N_26282,N_20039,N_21681);
or U26283 (N_26283,N_20695,N_24738);
nand U26284 (N_26284,N_23678,N_24021);
nand U26285 (N_26285,N_22902,N_22741);
or U26286 (N_26286,N_20915,N_22100);
or U26287 (N_26287,N_23187,N_20005);
or U26288 (N_26288,N_21828,N_21154);
or U26289 (N_26289,N_21428,N_24749);
nor U26290 (N_26290,N_20065,N_23080);
xnor U26291 (N_26291,N_20796,N_22533);
and U26292 (N_26292,N_24465,N_21981);
or U26293 (N_26293,N_21108,N_23133);
and U26294 (N_26294,N_21307,N_23620);
nand U26295 (N_26295,N_21105,N_24848);
nor U26296 (N_26296,N_23585,N_23351);
xnor U26297 (N_26297,N_20731,N_22002);
and U26298 (N_26298,N_21523,N_24032);
xor U26299 (N_26299,N_20954,N_23435);
and U26300 (N_26300,N_22018,N_23257);
nor U26301 (N_26301,N_24700,N_23228);
xor U26302 (N_26302,N_22754,N_24787);
or U26303 (N_26303,N_22893,N_22512);
xor U26304 (N_26304,N_20420,N_23660);
and U26305 (N_26305,N_22508,N_23421);
nand U26306 (N_26306,N_21020,N_21507);
or U26307 (N_26307,N_21815,N_24670);
xor U26308 (N_26308,N_20938,N_23781);
or U26309 (N_26309,N_21999,N_21189);
xnor U26310 (N_26310,N_21379,N_21782);
or U26311 (N_26311,N_21103,N_24622);
xor U26312 (N_26312,N_20830,N_21221);
nand U26313 (N_26313,N_23783,N_22995);
or U26314 (N_26314,N_22246,N_23755);
or U26315 (N_26315,N_20194,N_20152);
or U26316 (N_26316,N_21030,N_20098);
nor U26317 (N_26317,N_24841,N_23059);
nand U26318 (N_26318,N_21632,N_21832);
or U26319 (N_26319,N_21489,N_24173);
xnor U26320 (N_26320,N_22929,N_22961);
xnor U26321 (N_26321,N_21071,N_20431);
or U26322 (N_26322,N_20395,N_22722);
and U26323 (N_26323,N_22889,N_21658);
xnor U26324 (N_26324,N_20177,N_22976);
and U26325 (N_26325,N_21227,N_24759);
or U26326 (N_26326,N_21511,N_24497);
nand U26327 (N_26327,N_23920,N_24418);
or U26328 (N_26328,N_20272,N_22306);
or U26329 (N_26329,N_23948,N_22244);
and U26330 (N_26330,N_23681,N_23545);
or U26331 (N_26331,N_23558,N_20858);
nand U26332 (N_26332,N_22714,N_23740);
or U26333 (N_26333,N_20472,N_22233);
and U26334 (N_26334,N_22273,N_22526);
xnor U26335 (N_26335,N_24557,N_24646);
nand U26336 (N_26336,N_20064,N_21237);
nand U26337 (N_26337,N_20419,N_22509);
nor U26338 (N_26338,N_21046,N_21370);
or U26339 (N_26339,N_20744,N_23584);
xor U26340 (N_26340,N_24743,N_23056);
and U26341 (N_26341,N_21801,N_24620);
or U26342 (N_26342,N_20233,N_20416);
xnor U26343 (N_26343,N_22869,N_20980);
nor U26344 (N_26344,N_20969,N_20135);
and U26345 (N_26345,N_22460,N_21535);
or U26346 (N_26346,N_22558,N_21544);
xor U26347 (N_26347,N_23976,N_20852);
and U26348 (N_26348,N_22137,N_24921);
and U26349 (N_26349,N_20517,N_21220);
and U26350 (N_26350,N_22463,N_22316);
or U26351 (N_26351,N_20554,N_23212);
or U26352 (N_26352,N_24643,N_20524);
nor U26353 (N_26353,N_20747,N_21438);
and U26354 (N_26354,N_24713,N_24102);
nand U26355 (N_26355,N_23064,N_22067);
nor U26356 (N_26356,N_23021,N_20314);
xor U26357 (N_26357,N_23030,N_22498);
nand U26358 (N_26358,N_24607,N_21717);
nor U26359 (N_26359,N_24846,N_22969);
nand U26360 (N_26360,N_23944,N_22191);
or U26361 (N_26361,N_20070,N_22632);
nand U26362 (N_26362,N_23759,N_20400);
nor U26363 (N_26363,N_23956,N_21526);
or U26364 (N_26364,N_21683,N_24502);
xnor U26365 (N_26365,N_20199,N_21005);
and U26366 (N_26366,N_23482,N_21601);
and U26367 (N_26367,N_23574,N_22031);
or U26368 (N_26368,N_21338,N_20450);
or U26369 (N_26369,N_20436,N_20122);
nand U26370 (N_26370,N_24811,N_20355);
nor U26371 (N_26371,N_22587,N_23827);
nand U26372 (N_26372,N_24819,N_24276);
or U26373 (N_26373,N_20572,N_21676);
nand U26374 (N_26374,N_22535,N_20555);
nand U26375 (N_26375,N_24463,N_22004);
nor U26376 (N_26376,N_23178,N_22519);
nand U26377 (N_26377,N_24980,N_22668);
xor U26378 (N_26378,N_23928,N_22264);
nor U26379 (N_26379,N_20228,N_21461);
nor U26380 (N_26380,N_21131,N_21113);
or U26381 (N_26381,N_21948,N_24092);
or U26382 (N_26382,N_22271,N_22481);
and U26383 (N_26383,N_21436,N_21483);
or U26384 (N_26384,N_24247,N_23732);
nand U26385 (N_26385,N_22843,N_22069);
nand U26386 (N_26386,N_20724,N_22896);
or U26387 (N_26387,N_22866,N_24628);
or U26388 (N_26388,N_21845,N_20465);
nor U26389 (N_26389,N_24044,N_24741);
nor U26390 (N_26390,N_22387,N_24183);
nand U26391 (N_26391,N_23575,N_21553);
xnor U26392 (N_26392,N_22006,N_20282);
or U26393 (N_26393,N_20422,N_22738);
or U26394 (N_26394,N_22015,N_24638);
or U26395 (N_26395,N_24488,N_24157);
xor U26396 (N_26396,N_21798,N_21699);
nand U26397 (N_26397,N_22713,N_24608);
xnor U26398 (N_26398,N_20106,N_24297);
nor U26399 (N_26399,N_22724,N_23316);
xor U26400 (N_26400,N_22808,N_21842);
and U26401 (N_26401,N_23997,N_21362);
or U26402 (N_26402,N_24719,N_23834);
nand U26403 (N_26403,N_24018,N_21582);
or U26404 (N_26404,N_22614,N_23499);
nor U26405 (N_26405,N_22986,N_23409);
or U26406 (N_26406,N_21753,N_22402);
nand U26407 (N_26407,N_22121,N_20513);
nand U26408 (N_26408,N_23361,N_21223);
or U26409 (N_26409,N_21612,N_24960);
nor U26410 (N_26410,N_20667,N_23206);
nand U26411 (N_26411,N_21453,N_23020);
or U26412 (N_26412,N_24416,N_23961);
nand U26413 (N_26413,N_22833,N_23278);
nor U26414 (N_26414,N_24268,N_22339);
or U26415 (N_26415,N_21825,N_22034);
xnor U26416 (N_26416,N_20462,N_20764);
and U26417 (N_26417,N_23774,N_24284);
and U26418 (N_26418,N_24788,N_22862);
nand U26419 (N_26419,N_24041,N_22870);
nand U26420 (N_26420,N_21282,N_22061);
xor U26421 (N_26421,N_23596,N_22212);
nor U26422 (N_26422,N_20477,N_22599);
nand U26423 (N_26423,N_24469,N_21905);
or U26424 (N_26424,N_21646,N_20562);
xnor U26425 (N_26425,N_20723,N_20403);
nand U26426 (N_26426,N_23836,N_23054);
and U26427 (N_26427,N_21324,N_21931);
or U26428 (N_26428,N_20502,N_23890);
and U26429 (N_26429,N_23741,N_23940);
nor U26430 (N_26430,N_22926,N_20209);
and U26431 (N_26431,N_22107,N_23539);
nand U26432 (N_26432,N_22314,N_22281);
or U26433 (N_26433,N_24640,N_22455);
nor U26434 (N_26434,N_23510,N_21075);
nor U26435 (N_26435,N_24904,N_22307);
and U26436 (N_26436,N_20904,N_21424);
and U26437 (N_26437,N_20845,N_24874);
nand U26438 (N_26438,N_20773,N_24619);
nand U26439 (N_26439,N_23327,N_20660);
nor U26440 (N_26440,N_21133,N_20035);
and U26441 (N_26441,N_22390,N_21442);
nor U26442 (N_26442,N_22480,N_24766);
xnor U26443 (N_26443,N_21764,N_20125);
and U26444 (N_26444,N_20421,N_20633);
xor U26445 (N_26445,N_20285,N_24866);
and U26446 (N_26446,N_22023,N_24116);
xnor U26447 (N_26447,N_21423,N_21193);
or U26448 (N_26448,N_23084,N_24556);
xor U26449 (N_26449,N_20269,N_21977);
nand U26450 (N_26450,N_20907,N_23433);
xor U26451 (N_26451,N_23006,N_22613);
xor U26452 (N_26452,N_20425,N_23856);
xnor U26453 (N_26453,N_22575,N_20371);
nor U26454 (N_26454,N_20824,N_24941);
nor U26455 (N_26455,N_21284,N_24264);
nand U26456 (N_26456,N_24891,N_21943);
and U26457 (N_26457,N_23664,N_20512);
or U26458 (N_26458,N_22678,N_24661);
or U26459 (N_26459,N_22162,N_23503);
nor U26460 (N_26460,N_23166,N_21196);
nor U26461 (N_26461,N_21603,N_21572);
or U26462 (N_26462,N_20788,N_21074);
or U26463 (N_26463,N_21809,N_20113);
or U26464 (N_26464,N_20839,N_22839);
or U26465 (N_26465,N_23248,N_24756);
nor U26466 (N_26466,N_20338,N_23106);
and U26467 (N_26467,N_20280,N_23332);
nor U26468 (N_26468,N_23546,N_20859);
xnor U26469 (N_26469,N_24374,N_20257);
nor U26470 (N_26470,N_23379,N_24701);
nand U26471 (N_26471,N_23436,N_24587);
nand U26472 (N_26472,N_24807,N_22003);
or U26473 (N_26473,N_21949,N_23391);
nor U26474 (N_26474,N_24358,N_23859);
and U26475 (N_26475,N_21758,N_24019);
and U26476 (N_26476,N_24780,N_24126);
xor U26477 (N_26477,N_21357,N_21998);
xnor U26478 (N_26478,N_23655,N_24734);
nand U26479 (N_26479,N_21735,N_22489);
nor U26480 (N_26480,N_24651,N_24535);
nor U26481 (N_26481,N_24438,N_23116);
nand U26482 (N_26482,N_24634,N_24555);
xor U26483 (N_26483,N_21271,N_22355);
nand U26484 (N_26484,N_24585,N_22520);
nor U26485 (N_26485,N_21769,N_23603);
nand U26486 (N_26486,N_21152,N_20043);
nand U26487 (N_26487,N_24925,N_23375);
nor U26488 (N_26488,N_21703,N_20815);
or U26489 (N_26489,N_23353,N_22407);
nand U26490 (N_26490,N_24832,N_23810);
and U26491 (N_26491,N_20112,N_20919);
or U26492 (N_26492,N_24326,N_23147);
nor U26493 (N_26493,N_22568,N_23874);
nor U26494 (N_26494,N_23234,N_22482);
xnor U26495 (N_26495,N_24907,N_22371);
nand U26496 (N_26496,N_20701,N_22028);
xor U26497 (N_26497,N_20319,N_23764);
xnor U26498 (N_26498,N_21768,N_24452);
nand U26499 (N_26499,N_20408,N_23319);
xor U26500 (N_26500,N_20287,N_24669);
and U26501 (N_26501,N_21349,N_21656);
and U26502 (N_26502,N_24129,N_22058);
nor U26503 (N_26503,N_24017,N_22400);
xnor U26504 (N_26504,N_21836,N_20432);
nand U26505 (N_26505,N_20326,N_23505);
xor U26506 (N_26506,N_24604,N_22491);
nor U26507 (N_26507,N_20054,N_20316);
xnor U26508 (N_26508,N_24430,N_21469);
and U26509 (N_26509,N_24217,N_22898);
xor U26510 (N_26510,N_22236,N_20090);
nor U26511 (N_26511,N_24579,N_20156);
or U26512 (N_26512,N_20252,N_24722);
nand U26513 (N_26513,N_24875,N_20671);
nor U26514 (N_26514,N_23448,N_22207);
xor U26515 (N_26515,N_23987,N_22564);
and U26516 (N_26516,N_22598,N_23529);
nor U26517 (N_26517,N_22393,N_21473);
or U26518 (N_26518,N_22299,N_24400);
or U26519 (N_26519,N_21742,N_20971);
or U26520 (N_26520,N_22359,N_23262);
and U26521 (N_26521,N_22019,N_22092);
xnor U26522 (N_26522,N_23567,N_20430);
xnor U26523 (N_26523,N_22064,N_24428);
xnor U26524 (N_26524,N_20841,N_23909);
nor U26525 (N_26525,N_20267,N_22914);
nand U26526 (N_26526,N_20047,N_22605);
nor U26527 (N_26527,N_21065,N_21390);
or U26528 (N_26528,N_24988,N_20057);
nand U26529 (N_26529,N_22063,N_20396);
or U26530 (N_26530,N_21093,N_22746);
nor U26531 (N_26531,N_20774,N_20970);
or U26532 (N_26532,N_24830,N_23401);
nand U26533 (N_26533,N_21574,N_21655);
nand U26534 (N_26534,N_21810,N_22972);
nand U26535 (N_26535,N_23912,N_23959);
or U26536 (N_26536,N_23713,N_21200);
or U26537 (N_26537,N_21746,N_24188);
nand U26538 (N_26538,N_21736,N_20752);
or U26539 (N_26539,N_23478,N_22416);
xnor U26540 (N_26540,N_20889,N_20685);
and U26541 (N_26541,N_22483,N_20860);
nand U26542 (N_26542,N_21095,N_22933);
nand U26543 (N_26543,N_21940,N_21303);
nor U26544 (N_26544,N_23016,N_20651);
nand U26545 (N_26545,N_23413,N_23765);
nor U26546 (N_26546,N_20621,N_21928);
nand U26547 (N_26547,N_23438,N_24910);
nor U26548 (N_26548,N_20129,N_24527);
or U26549 (N_26549,N_22353,N_23622);
nor U26550 (N_26550,N_22546,N_23027);
xnor U26551 (N_26551,N_23531,N_22679);
or U26552 (N_26552,N_21164,N_23518);
nor U26553 (N_26553,N_21911,N_24533);
nor U26554 (N_26554,N_20366,N_24818);
nand U26555 (N_26555,N_21989,N_24334);
and U26556 (N_26556,N_24588,N_22650);
or U26557 (N_26557,N_24509,N_20922);
nor U26558 (N_26558,N_21935,N_24654);
xor U26559 (N_26559,N_21092,N_24152);
and U26560 (N_26560,N_22864,N_23516);
or U26561 (N_26561,N_21546,N_21910);
nor U26562 (N_26562,N_20875,N_21270);
xor U26563 (N_26563,N_23892,N_20878);
xnor U26564 (N_26564,N_22468,N_23761);
or U26565 (N_26565,N_24127,N_23710);
nor U26566 (N_26566,N_24795,N_20973);
nor U26567 (N_26567,N_20574,N_22975);
nor U26568 (N_26568,N_24335,N_23514);
and U26569 (N_26569,N_22670,N_22604);
and U26570 (N_26570,N_24216,N_22500);
and U26571 (N_26571,N_24124,N_23862);
nand U26572 (N_26572,N_21201,N_24806);
nor U26573 (N_26573,N_23564,N_21734);
nand U26574 (N_26574,N_23337,N_22338);
xnor U26575 (N_26575,N_23661,N_23207);
nor U26576 (N_26576,N_21892,N_23430);
xnor U26577 (N_26577,N_21745,N_21956);
nand U26578 (N_26578,N_23210,N_24246);
nor U26579 (N_26579,N_24175,N_24008);
nor U26580 (N_26580,N_20850,N_20274);
nand U26581 (N_26581,N_22257,N_22369);
nor U26582 (N_26582,N_20630,N_23014);
xnor U26583 (N_26583,N_24605,N_21732);
xnor U26584 (N_26584,N_24443,N_23634);
nor U26585 (N_26585,N_20149,N_24177);
nor U26586 (N_26586,N_23735,N_23442);
or U26587 (N_26587,N_20645,N_23784);
or U26588 (N_26588,N_24937,N_22153);
nand U26589 (N_26589,N_22505,N_24242);
nand U26590 (N_26590,N_20757,N_20947);
or U26591 (N_26591,N_24248,N_23293);
or U26592 (N_26592,N_22456,N_20570);
or U26593 (N_26593,N_22717,N_20709);
or U26594 (N_26594,N_22171,N_22595);
xnor U26595 (N_26595,N_23297,N_22073);
nand U26596 (N_26596,N_20673,N_20173);
nor U26597 (N_26597,N_20253,N_24851);
nand U26598 (N_26598,N_21626,N_24471);
or U26599 (N_26599,N_20362,N_20714);
and U26600 (N_26600,N_23012,N_22446);
nor U26601 (N_26601,N_24648,N_21418);
and U26602 (N_26602,N_21053,N_21974);
nand U26603 (N_26603,N_23864,N_24450);
xor U26604 (N_26604,N_24802,N_24059);
nor U26605 (N_26605,N_21807,N_21830);
nor U26606 (N_26606,N_21162,N_23437);
and U26607 (N_26607,N_23100,N_21654);
nand U26608 (N_26608,N_20077,N_24338);
or U26609 (N_26609,N_20325,N_20169);
or U26610 (N_26610,N_20215,N_21886);
and U26611 (N_26611,N_23951,N_22573);
nand U26612 (N_26612,N_24310,N_20132);
or U26613 (N_26613,N_22270,N_22209);
nor U26614 (N_26614,N_21942,N_24111);
or U26615 (N_26615,N_21012,N_20443);
xor U26616 (N_26616,N_20808,N_23113);
nor U26617 (N_26617,N_23729,N_21001);
xnor U26618 (N_26618,N_23124,N_23926);
or U26619 (N_26619,N_22242,N_23775);
nor U26620 (N_26620,N_21205,N_21014);
nor U26621 (N_26621,N_20848,N_20170);
xnor U26622 (N_26622,N_20831,N_24056);
nor U26623 (N_26623,N_20515,N_23694);
xnor U26624 (N_26624,N_22931,N_23748);
nand U26625 (N_26625,N_21167,N_20680);
xnor U26626 (N_26626,N_20553,N_21952);
xor U26627 (N_26627,N_20505,N_23602);
or U26628 (N_26628,N_21791,N_22664);
or U26629 (N_26629,N_22256,N_20636);
and U26630 (N_26630,N_23637,N_20948);
and U26631 (N_26631,N_22522,N_21668);
nor U26632 (N_26632,N_23123,N_22129);
xnor U26633 (N_26633,N_24270,N_20767);
xnor U26634 (N_26634,N_22368,N_20578);
nor U26635 (N_26635,N_22612,N_24470);
nor U26636 (N_26636,N_23875,N_24274);
or U26637 (N_26637,N_22052,N_21776);
nand U26638 (N_26638,N_22793,N_22919);
nand U26639 (N_26639,N_20912,N_24825);
xor U26640 (N_26640,N_23527,N_23705);
or U26641 (N_26641,N_23980,N_23916);
nand U26642 (N_26642,N_20045,N_22630);
xnor U26643 (N_26643,N_21921,N_21295);
nor U26644 (N_26644,N_20924,N_20191);
or U26645 (N_26645,N_21694,N_20262);
xnor U26646 (N_26646,N_21596,N_20195);
nand U26647 (N_26647,N_22303,N_23667);
xor U26648 (N_26648,N_24091,N_21100);
nor U26649 (N_26649,N_23731,N_24345);
or U26650 (N_26650,N_22946,N_23619);
nor U26651 (N_26651,N_24464,N_24953);
nor U26652 (N_26652,N_24885,N_23745);
and U26653 (N_26653,N_20703,N_20705);
and U26654 (N_26654,N_23879,N_24652);
nand U26655 (N_26655,N_23144,N_21662);
and U26656 (N_26656,N_20230,N_23162);
xor U26657 (N_26657,N_23460,N_22193);
nor U26658 (N_26658,N_22001,N_24683);
or U26659 (N_26659,N_20310,N_21035);
nand U26660 (N_26660,N_22486,N_23218);
nor U26661 (N_26661,N_20352,N_24492);
or U26662 (N_26662,N_21992,N_20540);
xor U26663 (N_26663,N_20812,N_20089);
nand U26664 (N_26664,N_21824,N_22324);
xnor U26665 (N_26665,N_21336,N_23399);
or U26666 (N_26666,N_22922,N_21474);
nand U26667 (N_26667,N_21889,N_23896);
nand U26668 (N_26668,N_23099,N_23808);
or U26669 (N_26669,N_24746,N_21486);
and U26670 (N_26670,N_22721,N_20360);
nand U26671 (N_26671,N_22742,N_22062);
and U26672 (N_26672,N_23406,N_24580);
xnor U26673 (N_26673,N_21411,N_24574);
nand U26674 (N_26674,N_20308,N_22132);
nor U26675 (N_26675,N_22918,N_20920);
or U26676 (N_26676,N_23697,N_22693);
nor U26677 (N_26677,N_21570,N_22619);
xor U26678 (N_26678,N_24192,N_20509);
and U26679 (N_26679,N_23734,N_21479);
xor U26680 (N_26680,N_22672,N_23863);
nor U26681 (N_26681,N_23326,N_22910);
xnor U26682 (N_26682,N_24716,N_24642);
nand U26683 (N_26683,N_23665,N_22727);
or U26684 (N_26684,N_22515,N_23942);
nor U26685 (N_26685,N_20657,N_20137);
nand U26686 (N_26686,N_20923,N_20148);
xor U26687 (N_26687,N_21151,N_20681);
nand U26688 (N_26688,N_24771,N_21597);
xnor U26689 (N_26689,N_22979,N_22232);
and U26690 (N_26690,N_20511,N_24167);
nand U26691 (N_26691,N_20381,N_24760);
nand U26692 (N_26692,N_23578,N_21279);
or U26693 (N_26693,N_20390,N_22900);
and U26694 (N_26694,N_22426,N_22351);
nor U26695 (N_26695,N_21997,N_21855);
nor U26696 (N_26696,N_24534,N_23487);
xnor U26697 (N_26697,N_23716,N_20792);
nor U26698 (N_26698,N_21689,N_21958);
nand U26699 (N_26699,N_23313,N_24207);
or U26700 (N_26700,N_21712,N_21532);
xor U26701 (N_26701,N_23700,N_24732);
nor U26702 (N_26702,N_22545,N_20494);
nor U26703 (N_26703,N_23121,N_24500);
xor U26704 (N_26704,N_23821,N_20913);
xor U26705 (N_26705,N_23419,N_22811);
nand U26706 (N_26706,N_21833,N_21222);
xnor U26707 (N_26707,N_22383,N_21081);
nor U26708 (N_26708,N_23743,N_24595);
xor U26709 (N_26709,N_23989,N_21636);
and U26710 (N_26710,N_21285,N_22330);
nand U26711 (N_26711,N_21344,N_22066);
nor U26712 (N_26712,N_23185,N_23907);
and U26713 (N_26713,N_22453,N_22051);
or U26714 (N_26714,N_24485,N_22585);
and U26715 (N_26715,N_22272,N_20564);
and U26716 (N_26716,N_21705,N_21640);
nor U26717 (N_26717,N_20157,N_24513);
and U26718 (N_26718,N_22988,N_20962);
xnor U26719 (N_26719,N_22845,N_20832);
or U26720 (N_26720,N_24565,N_20530);
nor U26721 (N_26721,N_22036,N_20160);
or U26722 (N_26722,N_21427,N_23727);
nand U26723 (N_26723,N_23547,N_21450);
nor U26724 (N_26724,N_22366,N_20444);
nor U26725 (N_26725,N_23842,N_23536);
xnor U26726 (N_26726,N_21510,N_20700);
or U26727 (N_26727,N_20532,N_23883);
or U26728 (N_26728,N_23826,N_22349);
or U26729 (N_26729,N_23979,N_21823);
nand U26730 (N_26730,N_21335,N_24858);
and U26731 (N_26731,N_20246,N_20945);
or U26732 (N_26732,N_24203,N_21298);
and U26733 (N_26733,N_20955,N_20765);
nor U26734 (N_26734,N_20546,N_24371);
and U26735 (N_26735,N_21172,N_24212);
and U26736 (N_26736,N_24043,N_20332);
or U26737 (N_26737,N_24035,N_22396);
nor U26738 (N_26738,N_21002,N_23019);
nand U26739 (N_26739,N_23322,N_20810);
and U26740 (N_26740,N_23243,N_20650);
nand U26741 (N_26741,N_23541,N_22010);
xnor U26742 (N_26742,N_20479,N_23601);
or U26743 (N_26743,N_24552,N_22055);
nand U26744 (N_26744,N_24653,N_23929);
and U26745 (N_26745,N_20514,N_24939);
nor U26746 (N_26746,N_21033,N_21547);
nand U26747 (N_26747,N_21425,N_22180);
and U26748 (N_26748,N_22397,N_21447);
xnor U26749 (N_26749,N_21747,N_21245);
xnor U26750 (N_26750,N_23128,N_23356);
and U26751 (N_26751,N_23449,N_22878);
nand U26752 (N_26752,N_22345,N_22213);
and U26753 (N_26753,N_21116,N_24455);
and U26754 (N_26754,N_23623,N_24406);
and U26755 (N_26755,N_21059,N_22609);
nor U26756 (N_26756,N_22154,N_21951);
xor U26757 (N_26757,N_20178,N_23001);
nand U26758 (N_26758,N_23790,N_23412);
nor U26759 (N_26759,N_20675,N_20426);
nor U26760 (N_26760,N_22177,N_24659);
or U26761 (N_26761,N_20789,N_21248);
nor U26762 (N_26762,N_23643,N_22090);
or U26763 (N_26763,N_24190,N_20266);
nor U26764 (N_26764,N_20569,N_22834);
and U26765 (N_26765,N_21385,N_23074);
xor U26766 (N_26766,N_22732,N_21729);
and U26767 (N_26767,N_22640,N_21013);
nand U26768 (N_26768,N_21286,N_20271);
nand U26769 (N_26769,N_21238,N_23882);
xor U26770 (N_26770,N_22514,N_24316);
or U26771 (N_26771,N_21730,N_22683);
or U26772 (N_26772,N_23098,N_22691);
nand U26773 (N_26773,N_24711,N_20953);
or U26774 (N_26774,N_24727,N_23869);
nand U26775 (N_26775,N_23577,N_23605);
xor U26776 (N_26776,N_22020,N_23646);
nor U26777 (N_26777,N_21188,N_24911);
nor U26778 (N_26778,N_22999,N_23633);
nor U26779 (N_26779,N_22861,N_22240);
or U26780 (N_26780,N_23231,N_23461);
or U26781 (N_26781,N_22072,N_24677);
xor U26782 (N_26782,N_24453,N_21971);
nand U26783 (N_26783,N_23591,N_24172);
nor U26784 (N_26784,N_22099,N_23296);
nand U26785 (N_26785,N_23509,N_24754);
and U26786 (N_26786,N_23220,N_21602);
or U26787 (N_26787,N_20687,N_23378);
nand U26788 (N_26788,N_20768,N_24436);
xor U26789 (N_26789,N_23936,N_24245);
or U26790 (N_26790,N_22944,N_24340);
and U26791 (N_26791,N_20559,N_24159);
or U26792 (N_26792,N_24506,N_21121);
and U26793 (N_26793,N_21456,N_24370);
nor U26794 (N_26794,N_23860,N_21680);
nor U26795 (N_26795,N_21025,N_20171);
xor U26796 (N_26796,N_21583,N_24424);
nor U26797 (N_26797,N_22319,N_21304);
xor U26798 (N_26798,N_20641,N_20164);
xnor U26799 (N_26799,N_23339,N_23090);
xnor U26800 (N_26800,N_22280,N_20368);
or U26801 (N_26801,N_24046,N_24305);
nor U26802 (N_26802,N_20674,N_20193);
and U26803 (N_26803,N_24426,N_21630);
nand U26804 (N_26804,N_23649,N_21858);
nand U26805 (N_26805,N_22730,N_21604);
xnor U26806 (N_26806,N_21591,N_24573);
nand U26807 (N_26807,N_20427,N_22951);
nor U26808 (N_26808,N_21697,N_22087);
xnor U26809 (N_26809,N_21672,N_23830);
and U26810 (N_26810,N_21757,N_20802);
nand U26811 (N_26811,N_23598,N_22217);
xnor U26812 (N_26812,N_24182,N_22593);
xnor U26813 (N_26813,N_24461,N_24076);
nand U26814 (N_26814,N_20369,N_21055);
or U26815 (N_26815,N_20775,N_22044);
or U26816 (N_26816,N_22735,N_24110);
and U26817 (N_26817,N_20021,N_24320);
nor U26818 (N_26818,N_23417,N_23227);
nor U26819 (N_26819,N_20196,N_21128);
nor U26820 (N_26820,N_22723,N_20244);
nor U26821 (N_26821,N_24990,N_20543);
nand U26822 (N_26822,N_23717,N_21258);
nor U26823 (N_26823,N_22105,N_22409);
and U26824 (N_26824,N_23739,N_20931);
nor U26825 (N_26825,N_20103,N_23127);
nand U26826 (N_26826,N_20220,N_24692);
nor U26827 (N_26827,N_24575,N_21257);
nand U26828 (N_26828,N_21171,N_21243);
nor U26829 (N_26829,N_22218,N_22168);
xor U26830 (N_26830,N_20605,N_23456);
or U26831 (N_26831,N_20235,N_23072);
nor U26832 (N_26832,N_23597,N_23462);
nor U26833 (N_26833,N_22186,N_23703);
nor U26834 (N_26834,N_20911,N_22528);
and U26835 (N_26835,N_21552,N_24468);
nor U26836 (N_26836,N_23125,N_22673);
nand U26837 (N_26837,N_20869,N_22551);
xor U26838 (N_26838,N_21852,N_21920);
or U26839 (N_26839,N_21207,N_21778);
nor U26840 (N_26840,N_23204,N_22580);
or U26841 (N_26841,N_20245,N_23814);
and U26842 (N_26842,N_24344,N_21478);
xnor U26843 (N_26843,N_22690,N_23069);
or U26844 (N_26844,N_21584,N_24597);
or U26845 (N_26845,N_22249,N_22634);
and U26846 (N_26846,N_23237,N_24236);
and U26847 (N_26847,N_24398,N_23782);
nor U26848 (N_26848,N_22040,N_22586);
nand U26849 (N_26849,N_24816,N_20357);
or U26850 (N_26850,N_23693,N_24601);
or U26851 (N_26851,N_22964,N_23003);
xor U26852 (N_26852,N_22136,N_24151);
and U26853 (N_26853,N_23005,N_24523);
xor U26854 (N_26854,N_22331,N_20917);
nand U26855 (N_26855,N_21536,N_22776);
xor U26856 (N_26856,N_22048,N_24144);
nand U26857 (N_26857,N_21135,N_22950);
nand U26858 (N_26858,N_21555,N_23631);
nor U26859 (N_26859,N_21472,N_23880);
xor U26860 (N_26860,N_20455,N_20888);
xnor U26861 (N_26861,N_24240,N_21106);
or U26862 (N_26862,N_22053,N_22511);
xor U26863 (N_26863,N_23122,N_24095);
nor U26864 (N_26864,N_20527,N_20534);
xor U26865 (N_26865,N_20545,N_22310);
and U26866 (N_26866,N_24917,N_20950);
xnor U26867 (N_26867,N_23644,N_21315);
nand U26868 (N_26868,N_22552,N_24847);
or U26869 (N_26869,N_22269,N_20769);
or U26870 (N_26870,N_23675,N_23911);
and U26871 (N_26871,N_20756,N_20386);
nand U26872 (N_26872,N_21190,N_24962);
or U26873 (N_26873,N_21422,N_22049);
or U26874 (N_26874,N_23953,N_22405);
nor U26875 (N_26875,N_21569,N_23544);
nor U26876 (N_26876,N_23275,N_22656);
or U26877 (N_26877,N_20742,N_23762);
and U26878 (N_26878,N_20217,N_22831);
nor U26879 (N_26879,N_22160,N_24972);
and U26880 (N_26880,N_24645,N_23962);
and U26881 (N_26881,N_24224,N_22344);
xnor U26882 (N_26882,N_24501,N_23568);
nand U26883 (N_26883,N_21242,N_21458);
nor U26884 (N_26884,N_23160,N_22095);
or U26885 (N_26885,N_23763,N_23967);
and U26886 (N_26886,N_23723,N_22300);
nand U26887 (N_26887,N_23357,N_22641);
nand U26888 (N_26888,N_24747,N_20469);
nor U26889 (N_26889,N_21774,N_24505);
nor U26890 (N_26890,N_24440,N_24075);
nand U26891 (N_26891,N_20126,N_20468);
nor U26892 (N_26892,N_20921,N_21346);
or U26893 (N_26893,N_22477,N_24201);
and U26894 (N_26894,N_22884,N_23276);
or U26895 (N_26895,N_23191,N_24881);
or U26896 (N_26896,N_20181,N_23522);
nand U26897 (N_26897,N_21274,N_21468);
nand U26898 (N_26898,N_22745,N_20139);
or U26899 (N_26899,N_23151,N_24676);
nand U26900 (N_26900,N_23076,N_24195);
or U26901 (N_26901,N_22187,N_22760);
or U26902 (N_26902,N_21490,N_24278);
or U26903 (N_26903,N_24855,N_22828);
or U26904 (N_26904,N_20944,N_20708);
xnor U26905 (N_26905,N_20343,N_20144);
nand U26906 (N_26906,N_21704,N_24287);
nor U26907 (N_26907,N_22530,N_24006);
xor U26908 (N_26908,N_20018,N_22510);
nand U26909 (N_26909,N_20786,N_24625);
nand U26910 (N_26910,N_23177,N_24410);
or U26911 (N_26911,N_23704,N_22158);
xnor U26912 (N_26912,N_23338,N_23669);
nor U26913 (N_26913,N_22433,N_21533);
or U26914 (N_26914,N_22909,N_24113);
nor U26915 (N_26915,N_24495,N_20187);
or U26916 (N_26916,N_23798,N_23701);
nor U26917 (N_26917,N_21877,N_23561);
nand U26918 (N_26918,N_20110,N_22915);
nand U26919 (N_26919,N_21347,N_24218);
nor U26920 (N_26920,N_24359,N_22621);
nor U26921 (N_26921,N_22850,N_24784);
nor U26922 (N_26922,N_20092,N_22008);
and U26923 (N_26923,N_23616,N_22206);
or U26924 (N_26924,N_22852,N_20013);
nor U26925 (N_26925,N_23570,N_23408);
xnor U26926 (N_26926,N_20927,N_23398);
nor U26927 (N_26927,N_22832,N_24134);
nand U26928 (N_26928,N_23426,N_23200);
or U26929 (N_26929,N_24228,N_21102);
or U26930 (N_26930,N_24285,N_24985);
and U26931 (N_26931,N_22287,N_23434);
and U26932 (N_26932,N_22479,N_24403);
nor U26933 (N_26933,N_24108,N_21962);
xnor U26934 (N_26934,N_22635,N_20389);
or U26935 (N_26935,N_23079,N_22311);
and U26936 (N_26936,N_20231,N_20963);
and U26937 (N_26937,N_22076,N_21397);
and U26938 (N_26938,N_20011,N_22430);
and U26939 (N_26939,N_23685,N_23668);
or U26940 (N_26940,N_21517,N_22322);
xnor U26941 (N_26941,N_24966,N_23274);
or U26942 (N_26942,N_21323,N_24942);
xor U26943 (N_26943,N_20078,N_20809);
nand U26944 (N_26944,N_24729,N_21677);
nor U26945 (N_26945,N_23787,N_24243);
and U26946 (N_26946,N_21783,N_21429);
nor U26947 (N_26947,N_23389,N_23239);
and U26948 (N_26948,N_21294,N_24947);
nand U26949 (N_26949,N_23330,N_20327);
nand U26950 (N_26950,N_23553,N_24781);
nand U26951 (N_26951,N_24593,N_24592);
nand U26952 (N_26952,N_22493,N_20843);
or U26953 (N_26953,N_20441,N_20303);
or U26954 (N_26954,N_23828,N_22235);
xor U26955 (N_26955,N_24016,N_21955);
and U26956 (N_26956,N_22194,N_21148);
nand U26957 (N_26957,N_24829,N_24664);
or U26958 (N_26958,N_21320,N_21760);
nor U26959 (N_26959,N_24252,N_22294);
xor U26960 (N_26960,N_24548,N_22112);
xnor U26961 (N_26961,N_23841,N_22688);
nor U26962 (N_26962,N_24834,N_24526);
or U26963 (N_26963,N_20147,N_20805);
nor U26964 (N_26964,N_20321,N_24974);
nor U26965 (N_26965,N_22258,N_21988);
xnor U26966 (N_26966,N_20335,N_22009);
nand U26967 (N_26967,N_23502,N_20016);
nor U26968 (N_26968,N_24794,N_24577);
nand U26969 (N_26969,N_23925,N_21854);
and U26970 (N_26970,N_23146,N_24967);
nor U26971 (N_26971,N_20760,N_23385);
or U26972 (N_26972,N_22577,N_21066);
nand U26973 (N_26973,N_22399,N_24518);
and U26974 (N_26974,N_24448,N_22924);
and U26975 (N_26975,N_24078,N_22370);
or U26976 (N_26976,N_21381,N_24231);
nor U26977 (N_26977,N_20001,N_21173);
nor U26978 (N_26978,N_21820,N_24765);
nand U26979 (N_26979,N_21806,N_20446);
nand U26980 (N_26980,N_21008,N_22027);
nor U26981 (N_26981,N_22638,N_20239);
nand U26982 (N_26982,N_24965,N_21208);
nand U26983 (N_26983,N_24913,N_22883);
nand U26984 (N_26984,N_24433,N_20728);
xnor U26985 (N_26985,N_24504,N_20735);
or U26986 (N_26986,N_24824,N_23673);
and U26987 (N_26987,N_20840,N_22560);
or U26988 (N_26988,N_20746,N_21302);
nand U26989 (N_26989,N_21159,N_23266);
and U26990 (N_26990,N_22868,N_24180);
and U26991 (N_26991,N_21332,N_21560);
and U26992 (N_26992,N_24202,N_22304);
and U26993 (N_26993,N_23171,N_21463);
and U26994 (N_26994,N_23268,N_22476);
or U26995 (N_26995,N_20608,N_24820);
and U26996 (N_26996,N_23849,N_23418);
nand U26997 (N_26997,N_23137,N_24949);
xnor U26998 (N_26998,N_21831,N_22699);
nand U26999 (N_26999,N_24036,N_22846);
xor U27000 (N_27000,N_20398,N_22661);
xnor U27001 (N_27001,N_23855,N_22795);
and U27002 (N_27002,N_21598,N_21410);
xnor U27003 (N_27003,N_21125,N_24220);
and U27004 (N_27004,N_20772,N_23988);
or U27005 (N_27005,N_24600,N_23489);
nand U27006 (N_27006,N_21682,N_23592);
or U27007 (N_27007,N_24466,N_23971);
or U27008 (N_27008,N_22917,N_20242);
nand U27009 (N_27009,N_22623,N_20992);
nand U27010 (N_27010,N_20084,N_22461);
xor U27011 (N_27011,N_24155,N_24723);
nor U27012 (N_27012,N_23420,N_20865);
nand U27013 (N_27013,N_20208,N_20716);
nor U27014 (N_27014,N_24589,N_24449);
nor U27015 (N_27015,N_24508,N_22364);
nor U27016 (N_27016,N_23612,N_23423);
and U27017 (N_27017,N_22350,N_21543);
or U27018 (N_27018,N_22117,N_23422);
nor U27019 (N_27019,N_20484,N_21181);
or U27020 (N_27020,N_22410,N_23184);
or U27021 (N_27021,N_24289,N_24918);
and U27022 (N_27022,N_24199,N_24803);
and U27023 (N_27023,N_22927,N_21822);
nor U27024 (N_27024,N_20049,N_20020);
and U27025 (N_27025,N_20051,N_24028);
or U27026 (N_27026,N_20648,N_22597);
or U27027 (N_27027,N_22412,N_22694);
nor U27028 (N_27028,N_21635,N_24963);
nor U27029 (N_27029,N_20071,N_21509);
nand U27030 (N_27030,N_24773,N_21728);
and U27031 (N_27031,N_20079,N_24294);
xnor U27032 (N_27032,N_20676,N_24599);
and U27033 (N_27033,N_23387,N_24768);
or U27034 (N_27034,N_22984,N_21445);
xnor U27035 (N_27035,N_22773,N_23663);
nor U27036 (N_27036,N_23323,N_21499);
nand U27037 (N_27037,N_21605,N_22014);
nand U27038 (N_27038,N_20028,N_22686);
xor U27039 (N_27039,N_23229,N_24943);
nand U27040 (N_27040,N_20304,N_20862);
nor U27041 (N_27041,N_22764,N_21107);
xnor U27042 (N_27042,N_21737,N_21767);
and U27043 (N_27043,N_23736,N_23043);
nand U27044 (N_27044,N_24880,N_21965);
nand U27045 (N_27045,N_21395,N_22126);
or U27046 (N_27046,N_24117,N_23039);
nor U27047 (N_27047,N_22681,N_24462);
nor U27048 (N_27048,N_20402,N_22985);
nand U27049 (N_27049,N_24560,N_21564);
xnor U27050 (N_27050,N_22671,N_20293);
xnor U27051 (N_27051,N_22358,N_21376);
and U27052 (N_27052,N_22639,N_23872);
xor U27053 (N_27053,N_22441,N_20407);
xnor U27054 (N_27054,N_22135,N_24636);
xor U27055 (N_27055,N_23582,N_23273);
nand U27056 (N_27056,N_24040,N_24053);
nand U27057 (N_27057,N_22906,N_24405);
nand U27058 (N_27058,N_24106,N_22277);
nor U27059 (N_27059,N_20939,N_20617);
nor U27060 (N_27060,N_20087,N_20854);
xnor U27061 (N_27061,N_24096,N_23348);
or U27062 (N_27062,N_21310,N_24512);
and U27063 (N_27063,N_24392,N_21933);
nand U27064 (N_27064,N_21191,N_22147);
nor U27065 (N_27065,N_20741,N_23488);
or U27066 (N_27066,N_20052,N_21393);
or U27067 (N_27067,N_24197,N_20597);
or U27068 (N_27068,N_24721,N_23803);
nor U27069 (N_27069,N_21808,N_22266);
or U27070 (N_27070,N_24899,N_20903);
nand U27071 (N_27071,N_20594,N_20984);
or U27072 (N_27072,N_22283,N_24923);
nor U27073 (N_27073,N_21915,N_23233);
nor U27074 (N_27074,N_21864,N_24143);
nand U27075 (N_27075,N_20699,N_20121);
or U27076 (N_27076,N_21064,N_21401);
nand U27077 (N_27077,N_21719,N_23493);
and U27078 (N_27078,N_21382,N_21124);
nand U27079 (N_27079,N_23343,N_22210);
nand U27080 (N_27080,N_21609,N_20861);
and U27081 (N_27081,N_20174,N_23903);
nor U27082 (N_27082,N_22555,N_21437);
nand U27083 (N_27083,N_20161,N_22682);
and U27084 (N_27084,N_23114,N_20210);
nor U27085 (N_27085,N_20154,N_23163);
xor U27086 (N_27086,N_23141,N_24421);
and U27087 (N_27087,N_24275,N_24957);
nor U27088 (N_27088,N_23194,N_24048);
and U27089 (N_27089,N_20415,N_22687);
nand U27090 (N_27090,N_22389,N_21283);
xor U27091 (N_27091,N_21904,N_21312);
xor U27092 (N_27092,N_23749,N_24010);
nor U27093 (N_27093,N_20928,N_23165);
or U27094 (N_27094,N_22329,N_20414);
xor U27095 (N_27095,N_22907,N_24250);
nor U27096 (N_27096,N_24065,N_20109);
nand U27097 (N_27097,N_22288,N_24926);
nand U27098 (N_27098,N_20987,N_24293);
xnor U27099 (N_27099,N_23439,N_24946);
or U27100 (N_27100,N_21916,N_20754);
and U27101 (N_27101,N_22017,N_22747);
nor U27102 (N_27102,N_23888,N_22128);
and U27103 (N_27103,N_22806,N_22601);
nor U27104 (N_27104,N_20475,N_21766);
xnor U27105 (N_27105,N_24072,N_21731);
and U27106 (N_27106,N_20356,N_24189);
or U27107 (N_27107,N_24745,N_23304);
and U27108 (N_27108,N_24235,N_24319);
and U27109 (N_27109,N_23476,N_21906);
or U27110 (N_27110,N_21944,N_23580);
or U27111 (N_27111,N_23746,N_21814);
nor U27112 (N_27112,N_23067,N_22133);
nand U27113 (N_27113,N_21885,N_23758);
or U27114 (N_27114,N_23062,N_22887);
or U27115 (N_27115,N_24074,N_24944);
and U27116 (N_27116,N_22544,N_23341);
nor U27117 (N_27117,N_23891,N_21176);
nand U27118 (N_27118,N_23498,N_24733);
nor U27119 (N_27119,N_22200,N_24277);
nand U27120 (N_27120,N_24478,N_23632);
nand U27121 (N_27121,N_23254,N_22513);
or U27122 (N_27122,N_20095,N_20743);
or U27123 (N_27123,N_24304,N_24902);
xnor U27124 (N_27124,N_20883,N_20983);
nor U27125 (N_27125,N_24629,N_22594);
nand U27126 (N_27126,N_24801,N_23776);
or U27127 (N_27127,N_24367,N_21718);
or U27128 (N_27128,N_21600,N_22325);
xor U27129 (N_27129,N_21000,N_21216);
and U27130 (N_27130,N_22298,N_22488);
or U27131 (N_27131,N_21938,N_22219);
nor U27132 (N_27132,N_24237,N_21912);
xor U27133 (N_27133,N_21627,N_21061);
or U27134 (N_27134,N_23715,N_23197);
or U27135 (N_27135,N_24030,N_21165);
xor U27136 (N_27136,N_22496,N_21579);
and U27137 (N_27137,N_24993,N_21358);
xnor U27138 (N_27138,N_20615,N_23770);
and U27139 (N_27139,N_23742,N_22094);
or U27140 (N_27140,N_20828,N_24456);
or U27141 (N_27141,N_21233,N_23131);
nor U27142 (N_27142,N_20908,N_24528);
and U27143 (N_27143,N_24549,N_20797);
xor U27144 (N_27144,N_23847,N_20424);
nand U27145 (N_27145,N_24737,N_24879);
and U27146 (N_27146,N_23639,N_23002);
nor U27147 (N_27147,N_22916,N_20793);
xnor U27148 (N_27148,N_24283,N_24356);
and U27149 (N_27149,N_24107,N_23047);
and U27150 (N_27150,N_22600,N_22751);
xor U27151 (N_27151,N_24857,N_22871);
nand U27152 (N_27152,N_24068,N_22045);
xor U27153 (N_27153,N_21350,N_21847);
nor U27154 (N_27154,N_20324,N_22321);
or U27155 (N_27155,N_21098,N_22243);
or U27156 (N_27156,N_22559,N_22948);
nor U27157 (N_27157,N_20359,N_20066);
and U27158 (N_27158,N_20445,N_24774);
xnor U27159 (N_27159,N_20473,N_20493);
and U27160 (N_27160,N_22205,N_24266);
xor U27161 (N_27161,N_23537,N_24256);
nand U27162 (N_27162,N_22840,N_20138);
xor U27163 (N_27163,N_21500,N_23235);
nand U27164 (N_27164,N_23820,N_22251);
or U27165 (N_27165,N_23726,N_24909);
or U27166 (N_27166,N_24292,N_23799);
nor U27167 (N_27167,N_21166,N_21826);
xnor U27168 (N_27168,N_23086,N_22068);
xnor U27169 (N_27169,N_22466,N_21970);
and U27170 (N_27170,N_24936,N_23594);
nor U27171 (N_27171,N_21322,N_20372);
xnor U27172 (N_27172,N_20358,N_22856);
nor U27173 (N_27173,N_21214,N_21868);
nor U27174 (N_27174,N_22562,N_23902);
and U27175 (N_27175,N_24912,N_23982);
or U27176 (N_27176,N_21426,N_21811);
xor U27177 (N_27177,N_21679,N_22123);
or U27178 (N_27178,N_24333,N_21969);
or U27179 (N_27179,N_21990,N_22301);
nor U27180 (N_27180,N_21628,N_24827);
and U27181 (N_27181,N_23991,N_21363);
xor U27182 (N_27182,N_21934,N_21466);
nor U27183 (N_27183,N_22170,N_23345);
nand U27184 (N_27184,N_24775,N_22881);
or U27185 (N_27185,N_23138,N_20201);
nand U27186 (N_27186,N_23927,N_23970);
nand U27187 (N_27187,N_22423,N_22164);
nor U27188 (N_27188,N_20976,N_20142);
xnor U27189 (N_27189,N_24384,N_23468);
xnor U27190 (N_27190,N_23077,N_23384);
xor U27191 (N_27191,N_23291,N_20749);
nand U27192 (N_27192,N_23941,N_23168);
xnor U27193 (N_27193,N_20091,N_21389);
and U27194 (N_27194,N_24900,N_23490);
nor U27195 (N_27195,N_23359,N_21932);
nand U27196 (N_27196,N_21240,N_20501);
and U27197 (N_27197,N_20818,N_22377);
or U27198 (N_27198,N_23272,N_20082);
nand U27199 (N_27199,N_24538,N_22119);
nor U27200 (N_27200,N_23720,N_22835);
nand U27201 (N_27201,N_22327,N_23346);
xnor U27202 (N_27202,N_23752,N_21613);
and U27203 (N_27203,N_24755,N_24698);
nand U27204 (N_27204,N_21785,N_21413);
and U27205 (N_27205,N_24887,N_20322);
nor U27206 (N_27206,N_22415,N_22054);
nor U27207 (N_27207,N_21226,N_24346);
and U27208 (N_27208,N_22385,N_20817);
and U27209 (N_27209,N_23672,N_23441);
nand U27210 (N_27210,N_22804,N_23370);
and U27211 (N_27211,N_24174,N_20281);
nor U27212 (N_27212,N_21530,N_24376);
nand U27213 (N_27213,N_20273,N_24103);
nand U27214 (N_27214,N_20365,N_21644);
nand U27215 (N_27215,N_21203,N_23188);
or U27216 (N_27216,N_21090,N_24254);
xnor U27217 (N_27217,N_21539,N_22332);
nand U27218 (N_27218,N_24633,N_24976);
xnor U27219 (N_27219,N_21039,N_24037);
nor U27220 (N_27220,N_24369,N_20994);
xnor U27221 (N_27221,N_23656,N_22043);
nand U27222 (N_27222,N_20237,N_21653);
or U27223 (N_27223,N_21412,N_24165);
or U27224 (N_27224,N_23085,N_23290);
xnor U27225 (N_27225,N_21578,N_20062);
xor U27226 (N_27226,N_23562,N_21420);
nor U27227 (N_27227,N_20771,N_24694);
xor U27228 (N_27228,N_20055,N_22185);
and U27229 (N_27229,N_21156,N_22093);
xnor U27230 (N_27230,N_22899,N_24402);
or U27231 (N_27231,N_22654,N_24255);
and U27232 (N_27232,N_20439,N_20625);
xor U27233 (N_27233,N_20637,N_24225);
nand U27234 (N_27234,N_20376,N_21621);
nor U27235 (N_27235,N_21337,N_23996);
nand U27236 (N_27236,N_21976,N_23045);
or U27237 (N_27237,N_22497,N_20896);
or U27238 (N_27238,N_23073,N_24067);
xor U27239 (N_27239,N_23671,N_24300);
and U27240 (N_27240,N_22284,N_21954);
nor U27241 (N_27241,N_20885,N_20248);
or U27242 (N_27242,N_20080,N_22616);
nor U27243 (N_27243,N_23224,N_24142);
nor U27244 (N_27244,N_22648,N_22882);
xnor U27245 (N_27245,N_22712,N_20663);
and U27246 (N_27246,N_24992,N_24459);
nand U27247 (N_27247,N_23446,N_20541);
or U27248 (N_27248,N_21884,N_21142);
nand U27249 (N_27249,N_23845,N_21476);
xnor U27250 (N_27250,N_23044,N_23698);
or U27251 (N_27251,N_20659,N_21063);
nand U27252 (N_27252,N_20697,N_24382);
nand U27253 (N_27253,N_21070,N_24357);
xnor U27254 (N_27254,N_20713,N_23055);
nand U27255 (N_27255,N_21922,N_22706);
and U27256 (N_27256,N_20385,N_20601);
xor U27257 (N_27257,N_21599,N_21330);
xor U27258 (N_27258,N_23111,N_21241);
nand U27259 (N_27259,N_24118,N_21850);
or U27260 (N_27260,N_20707,N_23139);
xor U27261 (N_27261,N_23691,N_24311);
nor U27262 (N_27262,N_22963,N_22190);
nor U27263 (N_27263,N_21663,N_23640);
or U27264 (N_27264,N_24364,N_20165);
nand U27265 (N_27265,N_20526,N_24845);
nand U27266 (N_27266,N_23507,N_20014);
or U27267 (N_27267,N_21408,N_20531);
nand U27268 (N_27268,N_21155,N_23914);
nor U27269 (N_27269,N_24148,N_20846);
nand U27270 (N_27270,N_22292,N_22989);
and U27271 (N_27271,N_23145,N_24553);
and U27272 (N_27272,N_24049,N_23978);
nand U27273 (N_27273,N_22749,N_24390);
nor U27274 (N_27274,N_22591,N_22911);
nand U27275 (N_27275,N_20607,N_22649);
or U27276 (N_27276,N_21015,N_21565);
nor U27277 (N_27277,N_21485,N_24991);
nor U27278 (N_27278,N_20024,N_21317);
nor U27279 (N_27279,N_22354,N_21841);
or U27280 (N_27280,N_20250,N_23042);
nand U27281 (N_27281,N_23083,N_21813);
xor U27282 (N_27282,N_22748,N_22436);
or U27283 (N_27283,N_22196,N_23473);
and U27284 (N_27284,N_21345,N_22816);
xnor U27285 (N_27285,N_20393,N_21123);
and U27286 (N_27286,N_20353,N_23718);
or U27287 (N_27287,N_22817,N_21109);
and U27288 (N_27288,N_24290,N_24793);
xnor U27289 (N_27289,N_20593,N_24475);
or U27290 (N_27290,N_20884,N_21890);
xor U27291 (N_27291,N_20482,N_23410);
or U27292 (N_27292,N_24630,N_24379);
nand U27293 (N_27293,N_21101,N_23405);
xor U27294 (N_27294,N_22411,N_24895);
nand U27295 (N_27295,N_23070,N_23881);
nor U27296 (N_27296,N_24665,N_24908);
nor U27297 (N_27297,N_24714,N_23250);
nand U27298 (N_27298,N_22198,N_23260);
xnor U27299 (N_27299,N_22908,N_21387);
xor U27300 (N_27300,N_20940,N_22444);
or U27301 (N_27301,N_20835,N_22506);
nor U27302 (N_27302,N_24087,N_22786);
xor U27303 (N_27303,N_20753,N_20611);
nor U27304 (N_27304,N_24458,N_21670);
or U27305 (N_27305,N_24178,N_22529);
or U27306 (N_27306,N_23071,N_21611);
or U27307 (N_27307,N_22447,N_24761);
and U27308 (N_27308,N_20556,N_20655);
xnor U27309 (N_27309,N_20803,N_21792);
nor U27310 (N_27310,N_24969,N_22622);
or U27311 (N_27311,N_21975,N_24572);
and U27312 (N_27312,N_20798,N_20610);
nor U27313 (N_27313,N_20074,N_21018);
nor U27314 (N_27314,N_24353,N_22781);
nand U27315 (N_27315,N_21755,N_23087);
and U27316 (N_27316,N_21126,N_24210);
xnor U27317 (N_27317,N_22059,N_24389);
or U27318 (N_27318,N_20745,N_23031);
and U27319 (N_27319,N_24602,N_22805);
nor U27320 (N_27320,N_24758,N_22124);
or U27321 (N_27321,N_21406,N_21399);
nand U27322 (N_27322,N_23789,N_21031);
nand U27323 (N_27323,N_20510,N_21202);
nand U27324 (N_27324,N_21529,N_23295);
nor U27325 (N_27325,N_20010,N_23994);
xor U27326 (N_27326,N_21316,N_24397);
or U27327 (N_27327,N_23571,N_24093);
nor U27328 (N_27328,N_23621,N_21692);
xnor U27329 (N_27329,N_23506,N_20974);
xor U27330 (N_27330,N_23938,N_22932);
xnor U27331 (N_27331,N_21631,N_24710);
and U27332 (N_27332,N_24432,N_22229);
nand U27333 (N_27333,N_23657,N_21375);
nor U27334 (N_27334,N_24735,N_24656);
nor U27335 (N_27335,N_20624,N_23993);
or U27336 (N_27336,N_24132,N_23935);
nand U27337 (N_27337,N_23172,N_23246);
nor U27338 (N_27338,N_21744,N_23288);
or U27339 (N_27339,N_20937,N_24073);
and U27340 (N_27340,N_21365,N_20528);
and U27341 (N_27341,N_22361,N_24799);
or U27342 (N_27342,N_20670,N_23429);
and U27343 (N_27343,N_22966,N_22184);
and U27344 (N_27344,N_22666,N_24160);
and U27345 (N_27345,N_23066,N_23118);
nand U27346 (N_27346,N_22790,N_24570);
or U27347 (N_27347,N_21391,N_24695);
or U27348 (N_27348,N_20229,N_24821);
or U27349 (N_27349,N_22705,N_23103);
and U27350 (N_27350,N_23179,N_22978);
nor U27351 (N_27351,N_23352,N_24375);
nand U27352 (N_27352,N_20216,N_20027);
xnor U27353 (N_27353,N_23115,N_21577);
nor U27354 (N_27354,N_24859,N_22994);
nor U27355 (N_27355,N_24849,N_23760);
nand U27356 (N_27356,N_24576,N_24014);
and U27357 (N_27357,N_20131,N_20361);
or U27358 (N_27358,N_24566,N_21664);
nand U27359 (N_27359,N_21225,N_24545);
and U27360 (N_27360,N_24530,N_21048);
nand U27361 (N_27361,N_20698,N_23247);
nor U27362 (N_27362,N_21749,N_23475);
nand U27363 (N_27363,N_20224,N_24341);
nand U27364 (N_27364,N_23415,N_20033);
or U27365 (N_27365,N_20857,N_21006);
nor U27366 (N_27366,N_20495,N_24674);
and U27367 (N_27367,N_24681,N_24020);
xor U27368 (N_27368,N_23211,N_24744);
and U27369 (N_27369,N_20434,N_24221);
or U27370 (N_27370,N_21873,N_21289);
and U27371 (N_27371,N_23366,N_22949);
xnor U27372 (N_27372,N_23245,N_21514);
nor U27373 (N_27373,N_23450,N_23102);
or U27374 (N_27374,N_23853,N_23573);
xor U27375 (N_27375,N_22352,N_23344);
nand U27376 (N_27376,N_24088,N_23794);
xor U27377 (N_27377,N_20682,N_21540);
or U27378 (N_27378,N_21721,N_22675);
xnor U27379 (N_27379,N_20378,N_20058);
nand U27380 (N_27380,N_24380,N_22228);
nor U27381 (N_27381,N_23035,N_22101);
nand U27382 (N_27382,N_23320,N_22346);
nand U27383 (N_27383,N_22386,N_22767);
or U27384 (N_27384,N_23244,N_22521);
nand U27385 (N_27385,N_21204,N_20188);
nand U27386 (N_27386,N_23018,N_21120);
nand U27387 (N_27387,N_24054,N_24494);
or U27388 (N_27388,N_24914,N_22504);
xnor U27389 (N_27389,N_22615,N_22659);
or U27390 (N_27390,N_23867,N_21250);
and U27391 (N_27391,N_21146,N_20972);
nor U27392 (N_27392,N_21016,N_23328);
nor U27393 (N_27393,N_21846,N_20822);
nand U27394 (N_27394,N_21991,N_23788);
and U27395 (N_27395,N_20718,N_20068);
or U27396 (N_27396,N_23335,N_22253);
and U27397 (N_27397,N_20306,N_23528);
or U27398 (N_27398,N_22065,N_22636);
or U27399 (N_27399,N_22494,N_21927);
and U27400 (N_27400,N_21872,N_24690);
or U27401 (N_27401,N_23371,N_20184);
and U27402 (N_27402,N_21340,N_22503);
and U27403 (N_27403,N_24783,N_21919);
xnor U27404 (N_27404,N_20200,N_22578);
or U27405 (N_27405,N_22163,N_23985);
and U27406 (N_27406,N_21881,N_24934);
nand U27407 (N_27407,N_22752,N_21134);
and U27408 (N_27408,N_20813,N_21896);
nor U27409 (N_27409,N_23707,N_21648);
or U27410 (N_27410,N_20935,N_23258);
xnor U27411 (N_27411,N_24864,N_23615);
nor U27412 (N_27412,N_24261,N_23990);
nand U27413 (N_27413,N_24705,N_20189);
or U27414 (N_27414,N_20146,N_24489);
or U27415 (N_27415,N_23998,N_22782);
nor U27416 (N_27416,N_23120,N_21770);
nand U27417 (N_27417,N_22081,N_24260);
and U27418 (N_27418,N_22152,N_22876);
and U27419 (N_27419,N_24153,N_24882);
nand U27420 (N_27420,N_24003,N_22203);
xor U27421 (N_27421,N_24685,N_20046);
and U27422 (N_27422,N_23308,N_24214);
or U27423 (N_27423,N_24931,N_22553);
and U27424 (N_27424,N_22977,N_24146);
and U27425 (N_27425,N_20807,N_21645);
or U27426 (N_27426,N_22231,N_24667);
nor U27427 (N_27427,N_24663,N_23666);
nor U27428 (N_27428,N_23381,N_22873);
xor U27429 (N_27429,N_23733,N_22779);
nor U27430 (N_27430,N_21501,N_21673);
nand U27431 (N_27431,N_20851,N_21803);
nand U27432 (N_27432,N_21883,N_23515);
nor U27433 (N_27433,N_21267,N_24792);
and U27434 (N_27434,N_20717,N_21643);
or U27435 (N_27435,N_20059,N_21327);
or U27436 (N_27436,N_23906,N_23885);
nor U27437 (N_27437,N_23110,N_21153);
nand U27438 (N_27438,N_22921,N_21979);
nand U27439 (N_27439,N_20279,N_24978);
nand U27440 (N_27440,N_24454,N_23550);
or U27441 (N_27441,N_21661,N_24843);
or U27442 (N_27442,N_20571,N_21028);
xor U27443 (N_27443,N_23374,N_22176);
nand U27444 (N_27444,N_22227,N_22297);
or U27445 (N_27445,N_23091,N_22935);
nor U27446 (N_27446,N_22265,N_21057);
xnor U27447 (N_27447,N_22085,N_23368);
and U27448 (N_27448,N_23624,N_20263);
nand U27449 (N_27449,N_21446,N_23635);
nand U27450 (N_27450,N_23972,N_22204);
or U27451 (N_27451,N_20539,N_20936);
nand U27452 (N_27452,N_21995,N_20307);
nand U27453 (N_27453,N_24396,N_21713);
or U27454 (N_27454,N_22780,N_22424);
and U27455 (N_27455,N_22475,N_24540);
or U27456 (N_27456,N_22766,N_24179);
nor U27457 (N_27457,N_23795,N_20821);
nor U27458 (N_27458,N_22291,N_22131);
xnor U27459 (N_27459,N_23096,N_20738);
or U27460 (N_27460,N_22865,N_24460);
xnor U27461 (N_27461,N_23186,N_24427);
nor U27462 (N_27462,N_21325,N_24517);
xnor U27463 (N_27463,N_21660,N_23696);
and U27464 (N_27464,N_24331,N_23653);
and U27465 (N_27465,N_24309,N_21457);
nand U27466 (N_27466,N_23654,N_20946);
and U27467 (N_27467,N_22787,N_20206);
and U27468 (N_27468,N_21759,N_23886);
and U27469 (N_27469,N_24558,N_21314);
xor U27470 (N_27470,N_24419,N_20890);
nor U27471 (N_27471,N_22516,N_22289);
and U27472 (N_27472,N_20794,N_20566);
and U27473 (N_27473,N_20218,N_21085);
or U27474 (N_27474,N_20275,N_21278);
xnor U27475 (N_27475,N_21818,N_24208);
nand U27476 (N_27476,N_24004,N_22302);
nor U27477 (N_27477,N_22629,N_22260);
nor U27478 (N_27478,N_20914,N_20334);
or U27479 (N_27479,N_21122,N_20779);
and U27480 (N_27480,N_24033,N_21865);
nor U27481 (N_27481,N_24312,N_24804);
xor U27482 (N_27482,N_20075,N_21157);
xnor U27483 (N_27483,N_21924,N_20979);
nand U27484 (N_27484,N_23251,N_21280);
and U27485 (N_27485,N_21448,N_24810);
or U27486 (N_27486,N_21255,N_23767);
nor U27487 (N_27487,N_21748,N_24507);
nor U27488 (N_27488,N_24149,N_21026);
nor U27489 (N_27489,N_24678,N_20487);
or U27490 (N_27490,N_22109,N_24022);
or U27491 (N_27491,N_23769,N_22432);
and U27492 (N_27492,N_22942,N_24989);
nor U27493 (N_27493,N_23835,N_22967);
nand U27494 (N_27494,N_20653,N_23466);
and U27495 (N_27495,N_22337,N_20211);
and U27496 (N_27496,N_22802,N_24170);
nor U27497 (N_27497,N_20710,N_22211);
nor U27498 (N_27498,N_20664,N_23593);
nand U27499 (N_27499,N_23965,N_24109);
or U27500 (N_27500,N_22941,N_21320);
nor U27501 (N_27501,N_23581,N_21495);
and U27502 (N_27502,N_21085,N_23046);
nor U27503 (N_27503,N_22983,N_23747);
or U27504 (N_27504,N_20377,N_21961);
xnor U27505 (N_27505,N_22071,N_22375);
or U27506 (N_27506,N_22948,N_23293);
nand U27507 (N_27507,N_20465,N_20169);
nand U27508 (N_27508,N_20074,N_23786);
nor U27509 (N_27509,N_22512,N_21801);
or U27510 (N_27510,N_21519,N_21335);
and U27511 (N_27511,N_20045,N_21524);
and U27512 (N_27512,N_21990,N_23257);
nand U27513 (N_27513,N_22461,N_20572);
nand U27514 (N_27514,N_23990,N_24524);
and U27515 (N_27515,N_24348,N_22426);
xnor U27516 (N_27516,N_22777,N_20705);
nor U27517 (N_27517,N_20094,N_23447);
or U27518 (N_27518,N_24326,N_21902);
nor U27519 (N_27519,N_22339,N_21827);
nand U27520 (N_27520,N_21514,N_22819);
nor U27521 (N_27521,N_23430,N_23044);
nand U27522 (N_27522,N_21438,N_24154);
nand U27523 (N_27523,N_22498,N_21486);
and U27524 (N_27524,N_20437,N_20204);
nand U27525 (N_27525,N_24340,N_22300);
and U27526 (N_27526,N_24938,N_23371);
nand U27527 (N_27527,N_21625,N_20460);
nand U27528 (N_27528,N_21604,N_22442);
or U27529 (N_27529,N_24302,N_23104);
nand U27530 (N_27530,N_20572,N_20662);
or U27531 (N_27531,N_20146,N_24495);
xor U27532 (N_27532,N_24088,N_20854);
or U27533 (N_27533,N_22857,N_23187);
nor U27534 (N_27534,N_22272,N_20495);
nor U27535 (N_27535,N_21049,N_24504);
or U27536 (N_27536,N_23494,N_21749);
nand U27537 (N_27537,N_22328,N_21937);
nor U27538 (N_27538,N_21720,N_20667);
and U27539 (N_27539,N_22230,N_22667);
and U27540 (N_27540,N_24390,N_21259);
or U27541 (N_27541,N_23006,N_20664);
or U27542 (N_27542,N_23509,N_24619);
xnor U27543 (N_27543,N_21907,N_23932);
nor U27544 (N_27544,N_24260,N_21405);
nand U27545 (N_27545,N_22425,N_21342);
nor U27546 (N_27546,N_23354,N_24435);
xor U27547 (N_27547,N_23755,N_24105);
nor U27548 (N_27548,N_24532,N_20560);
xor U27549 (N_27549,N_20002,N_22213);
xnor U27550 (N_27550,N_22662,N_20616);
or U27551 (N_27551,N_21343,N_20706);
or U27552 (N_27552,N_21862,N_23879);
and U27553 (N_27553,N_23440,N_24989);
and U27554 (N_27554,N_24774,N_20684);
xor U27555 (N_27555,N_24511,N_23493);
and U27556 (N_27556,N_21039,N_20503);
nor U27557 (N_27557,N_24043,N_24939);
or U27558 (N_27558,N_22479,N_23487);
nor U27559 (N_27559,N_20132,N_22315);
and U27560 (N_27560,N_20137,N_21481);
and U27561 (N_27561,N_23921,N_23868);
and U27562 (N_27562,N_23081,N_23996);
nand U27563 (N_27563,N_23752,N_20089);
and U27564 (N_27564,N_22098,N_24567);
nor U27565 (N_27565,N_20812,N_23502);
and U27566 (N_27566,N_20011,N_24199);
or U27567 (N_27567,N_21947,N_23855);
nand U27568 (N_27568,N_21289,N_21643);
xor U27569 (N_27569,N_21178,N_23083);
xnor U27570 (N_27570,N_21084,N_23954);
nor U27571 (N_27571,N_24653,N_23416);
or U27572 (N_27572,N_21480,N_20818);
or U27573 (N_27573,N_22495,N_21498);
nand U27574 (N_27574,N_23881,N_22463);
or U27575 (N_27575,N_22086,N_22561);
or U27576 (N_27576,N_22980,N_22981);
or U27577 (N_27577,N_21148,N_20517);
nor U27578 (N_27578,N_24826,N_24244);
xnor U27579 (N_27579,N_24502,N_23213);
nand U27580 (N_27580,N_21723,N_21317);
and U27581 (N_27581,N_22577,N_22491);
nand U27582 (N_27582,N_22632,N_21571);
or U27583 (N_27583,N_20868,N_24747);
and U27584 (N_27584,N_22374,N_24494);
nand U27585 (N_27585,N_22694,N_21065);
or U27586 (N_27586,N_23280,N_24198);
or U27587 (N_27587,N_21113,N_23435);
and U27588 (N_27588,N_23849,N_23653);
or U27589 (N_27589,N_21515,N_20536);
and U27590 (N_27590,N_20819,N_22358);
xnor U27591 (N_27591,N_23825,N_24851);
nand U27592 (N_27592,N_20137,N_23677);
nand U27593 (N_27593,N_20757,N_20611);
and U27594 (N_27594,N_20082,N_20264);
or U27595 (N_27595,N_22318,N_22434);
nor U27596 (N_27596,N_22246,N_20542);
or U27597 (N_27597,N_22602,N_22860);
and U27598 (N_27598,N_22741,N_23559);
nor U27599 (N_27599,N_20106,N_23170);
and U27600 (N_27600,N_20443,N_22029);
or U27601 (N_27601,N_22995,N_22996);
nand U27602 (N_27602,N_24690,N_20354);
nor U27603 (N_27603,N_24709,N_20783);
and U27604 (N_27604,N_20578,N_23516);
and U27605 (N_27605,N_24428,N_21223);
or U27606 (N_27606,N_24789,N_24346);
nand U27607 (N_27607,N_24404,N_22655);
and U27608 (N_27608,N_23688,N_23374);
xor U27609 (N_27609,N_20584,N_23887);
and U27610 (N_27610,N_23520,N_21319);
nand U27611 (N_27611,N_21954,N_21491);
nor U27612 (N_27612,N_20849,N_20586);
nor U27613 (N_27613,N_23074,N_20960);
nand U27614 (N_27614,N_23767,N_24438);
nand U27615 (N_27615,N_23289,N_23927);
nor U27616 (N_27616,N_20862,N_20452);
nor U27617 (N_27617,N_22819,N_20757);
nor U27618 (N_27618,N_20285,N_23145);
and U27619 (N_27619,N_22134,N_24804);
nand U27620 (N_27620,N_21968,N_24469);
nand U27621 (N_27621,N_22503,N_21068);
nor U27622 (N_27622,N_23958,N_23452);
nor U27623 (N_27623,N_21140,N_22408);
nand U27624 (N_27624,N_24262,N_24043);
nand U27625 (N_27625,N_23110,N_24517);
or U27626 (N_27626,N_23580,N_21992);
nand U27627 (N_27627,N_22411,N_21488);
nor U27628 (N_27628,N_21117,N_23719);
nor U27629 (N_27629,N_22569,N_21446);
and U27630 (N_27630,N_24716,N_20396);
nor U27631 (N_27631,N_22758,N_23949);
and U27632 (N_27632,N_22930,N_22041);
or U27633 (N_27633,N_22588,N_24792);
xor U27634 (N_27634,N_21044,N_24435);
xor U27635 (N_27635,N_22741,N_23161);
and U27636 (N_27636,N_20291,N_22646);
or U27637 (N_27637,N_23582,N_20098);
nor U27638 (N_27638,N_20334,N_24545);
or U27639 (N_27639,N_21941,N_23105);
nor U27640 (N_27640,N_24547,N_23406);
nor U27641 (N_27641,N_22883,N_21056);
and U27642 (N_27642,N_21037,N_22586);
xor U27643 (N_27643,N_24453,N_22498);
xnor U27644 (N_27644,N_21529,N_21575);
and U27645 (N_27645,N_23362,N_23019);
nor U27646 (N_27646,N_22826,N_21862);
nor U27647 (N_27647,N_20293,N_21922);
xnor U27648 (N_27648,N_21283,N_23070);
and U27649 (N_27649,N_23956,N_23061);
and U27650 (N_27650,N_21755,N_24961);
and U27651 (N_27651,N_20487,N_20813);
xor U27652 (N_27652,N_22132,N_21525);
nor U27653 (N_27653,N_23983,N_22510);
nor U27654 (N_27654,N_23725,N_20238);
nand U27655 (N_27655,N_22839,N_23854);
nand U27656 (N_27656,N_22407,N_24540);
and U27657 (N_27657,N_24504,N_24574);
and U27658 (N_27658,N_20979,N_21768);
xnor U27659 (N_27659,N_23539,N_21072);
nor U27660 (N_27660,N_22462,N_21617);
or U27661 (N_27661,N_23943,N_21516);
or U27662 (N_27662,N_24350,N_23399);
xnor U27663 (N_27663,N_23867,N_22575);
xor U27664 (N_27664,N_20315,N_23439);
nand U27665 (N_27665,N_20833,N_21645);
xnor U27666 (N_27666,N_22753,N_21701);
or U27667 (N_27667,N_22915,N_21583);
and U27668 (N_27668,N_22284,N_23332);
nand U27669 (N_27669,N_24670,N_21684);
or U27670 (N_27670,N_21124,N_21225);
or U27671 (N_27671,N_24865,N_24405);
nor U27672 (N_27672,N_20194,N_22126);
and U27673 (N_27673,N_21575,N_24290);
or U27674 (N_27674,N_22175,N_24059);
and U27675 (N_27675,N_24257,N_23562);
and U27676 (N_27676,N_23366,N_20135);
and U27677 (N_27677,N_21240,N_24888);
or U27678 (N_27678,N_20924,N_23682);
or U27679 (N_27679,N_22549,N_21954);
nand U27680 (N_27680,N_24697,N_20400);
xor U27681 (N_27681,N_22437,N_20003);
nand U27682 (N_27682,N_24233,N_23347);
nand U27683 (N_27683,N_24747,N_24217);
xnor U27684 (N_27684,N_24835,N_22426);
xnor U27685 (N_27685,N_23339,N_20878);
or U27686 (N_27686,N_21637,N_22293);
nor U27687 (N_27687,N_21316,N_21514);
or U27688 (N_27688,N_20108,N_21842);
nor U27689 (N_27689,N_24470,N_21398);
nor U27690 (N_27690,N_23056,N_21059);
xnor U27691 (N_27691,N_21841,N_22646);
or U27692 (N_27692,N_21947,N_21928);
nand U27693 (N_27693,N_20250,N_23127);
nand U27694 (N_27694,N_20057,N_20401);
nor U27695 (N_27695,N_20382,N_21168);
and U27696 (N_27696,N_23246,N_24418);
nand U27697 (N_27697,N_24833,N_22863);
and U27698 (N_27698,N_20265,N_23625);
nand U27699 (N_27699,N_22752,N_20020);
or U27700 (N_27700,N_21315,N_24960);
or U27701 (N_27701,N_24819,N_22813);
and U27702 (N_27702,N_20528,N_24486);
nand U27703 (N_27703,N_21079,N_24743);
nor U27704 (N_27704,N_21914,N_20952);
nand U27705 (N_27705,N_22557,N_20936);
and U27706 (N_27706,N_23700,N_22499);
xor U27707 (N_27707,N_21919,N_20379);
xnor U27708 (N_27708,N_20687,N_20828);
and U27709 (N_27709,N_22206,N_21506);
or U27710 (N_27710,N_24844,N_21751);
nand U27711 (N_27711,N_21376,N_24445);
nand U27712 (N_27712,N_21645,N_23449);
nor U27713 (N_27713,N_21036,N_24502);
nor U27714 (N_27714,N_20002,N_23818);
nor U27715 (N_27715,N_23881,N_23326);
nor U27716 (N_27716,N_20453,N_21258);
nand U27717 (N_27717,N_21979,N_23836);
xor U27718 (N_27718,N_24916,N_22430);
nand U27719 (N_27719,N_21801,N_24616);
nand U27720 (N_27720,N_24295,N_22846);
xor U27721 (N_27721,N_21654,N_20495);
or U27722 (N_27722,N_24079,N_23772);
and U27723 (N_27723,N_24599,N_21742);
nor U27724 (N_27724,N_23372,N_24583);
xor U27725 (N_27725,N_20811,N_21734);
nor U27726 (N_27726,N_22081,N_22055);
or U27727 (N_27727,N_23074,N_22542);
nor U27728 (N_27728,N_24272,N_22547);
and U27729 (N_27729,N_24618,N_23877);
xnor U27730 (N_27730,N_23106,N_20314);
nor U27731 (N_27731,N_24369,N_22382);
nor U27732 (N_27732,N_20940,N_24019);
xor U27733 (N_27733,N_23264,N_24097);
nor U27734 (N_27734,N_22865,N_24924);
or U27735 (N_27735,N_24137,N_22237);
nand U27736 (N_27736,N_23797,N_22317);
xor U27737 (N_27737,N_24174,N_23361);
xor U27738 (N_27738,N_24710,N_21321);
and U27739 (N_27739,N_20946,N_23258);
or U27740 (N_27740,N_23574,N_20853);
or U27741 (N_27741,N_20514,N_24631);
nor U27742 (N_27742,N_23337,N_24790);
and U27743 (N_27743,N_21711,N_24159);
and U27744 (N_27744,N_23180,N_21862);
xnor U27745 (N_27745,N_22681,N_20703);
or U27746 (N_27746,N_22804,N_23902);
xor U27747 (N_27747,N_23688,N_23821);
nand U27748 (N_27748,N_21323,N_21162);
xnor U27749 (N_27749,N_23377,N_21658);
nand U27750 (N_27750,N_21188,N_23684);
nor U27751 (N_27751,N_21338,N_21326);
or U27752 (N_27752,N_22520,N_24172);
nor U27753 (N_27753,N_20696,N_21279);
nand U27754 (N_27754,N_21577,N_24356);
or U27755 (N_27755,N_23661,N_21340);
xnor U27756 (N_27756,N_20779,N_22501);
nor U27757 (N_27757,N_23591,N_24840);
or U27758 (N_27758,N_20310,N_21844);
or U27759 (N_27759,N_22521,N_21532);
nor U27760 (N_27760,N_24465,N_22633);
nand U27761 (N_27761,N_24738,N_20772);
and U27762 (N_27762,N_24078,N_21451);
nand U27763 (N_27763,N_20959,N_20532);
and U27764 (N_27764,N_22363,N_24195);
and U27765 (N_27765,N_24853,N_22413);
nand U27766 (N_27766,N_22462,N_21559);
nand U27767 (N_27767,N_21223,N_21111);
xor U27768 (N_27768,N_21463,N_24728);
and U27769 (N_27769,N_20603,N_24711);
nand U27770 (N_27770,N_24563,N_22850);
or U27771 (N_27771,N_23303,N_21446);
and U27772 (N_27772,N_24299,N_23817);
xor U27773 (N_27773,N_20089,N_23022);
or U27774 (N_27774,N_24275,N_21090);
nor U27775 (N_27775,N_21666,N_23631);
or U27776 (N_27776,N_21755,N_22926);
nor U27777 (N_27777,N_22819,N_24626);
xor U27778 (N_27778,N_22974,N_22798);
nor U27779 (N_27779,N_24211,N_20370);
xor U27780 (N_27780,N_21288,N_23860);
or U27781 (N_27781,N_20380,N_21456);
nand U27782 (N_27782,N_22257,N_22513);
or U27783 (N_27783,N_23299,N_23179);
xor U27784 (N_27784,N_24100,N_22491);
and U27785 (N_27785,N_22813,N_21894);
nor U27786 (N_27786,N_20654,N_24842);
nand U27787 (N_27787,N_20159,N_22951);
nor U27788 (N_27788,N_21572,N_23035);
and U27789 (N_27789,N_22198,N_21194);
nor U27790 (N_27790,N_24473,N_22442);
xnor U27791 (N_27791,N_24265,N_22846);
and U27792 (N_27792,N_20071,N_20003);
nor U27793 (N_27793,N_20016,N_22305);
xnor U27794 (N_27794,N_23416,N_23397);
and U27795 (N_27795,N_22385,N_24460);
and U27796 (N_27796,N_20174,N_23062);
nand U27797 (N_27797,N_23636,N_21605);
or U27798 (N_27798,N_24297,N_22191);
nor U27799 (N_27799,N_23915,N_23232);
nor U27800 (N_27800,N_22453,N_21486);
xor U27801 (N_27801,N_22273,N_20242);
and U27802 (N_27802,N_20064,N_21395);
and U27803 (N_27803,N_20173,N_23388);
nand U27804 (N_27804,N_21674,N_23807);
and U27805 (N_27805,N_23728,N_20500);
or U27806 (N_27806,N_20062,N_20501);
and U27807 (N_27807,N_24367,N_20230);
nor U27808 (N_27808,N_21147,N_20143);
and U27809 (N_27809,N_20995,N_24288);
or U27810 (N_27810,N_21197,N_23201);
nand U27811 (N_27811,N_24298,N_21646);
and U27812 (N_27812,N_20397,N_21078);
nor U27813 (N_27813,N_21018,N_22539);
xnor U27814 (N_27814,N_23417,N_22678);
nor U27815 (N_27815,N_23541,N_22303);
and U27816 (N_27816,N_24713,N_21056);
nor U27817 (N_27817,N_20234,N_22801);
and U27818 (N_27818,N_20024,N_23799);
nand U27819 (N_27819,N_23771,N_24633);
and U27820 (N_27820,N_21867,N_21296);
nor U27821 (N_27821,N_23685,N_23651);
xnor U27822 (N_27822,N_24005,N_23718);
xnor U27823 (N_27823,N_22754,N_22128);
nand U27824 (N_27824,N_21279,N_20797);
and U27825 (N_27825,N_20352,N_20885);
nor U27826 (N_27826,N_21818,N_23371);
nor U27827 (N_27827,N_22528,N_20503);
nand U27828 (N_27828,N_21762,N_20303);
and U27829 (N_27829,N_22146,N_22321);
nor U27830 (N_27830,N_23565,N_21311);
xor U27831 (N_27831,N_21734,N_21356);
nand U27832 (N_27832,N_24672,N_21648);
nand U27833 (N_27833,N_22371,N_22100);
nand U27834 (N_27834,N_24520,N_23961);
xor U27835 (N_27835,N_21969,N_21199);
nand U27836 (N_27836,N_21498,N_24596);
nor U27837 (N_27837,N_21534,N_24199);
nand U27838 (N_27838,N_21342,N_24076);
or U27839 (N_27839,N_21440,N_23750);
and U27840 (N_27840,N_24380,N_20348);
nand U27841 (N_27841,N_24229,N_24591);
xnor U27842 (N_27842,N_20752,N_22005);
or U27843 (N_27843,N_20308,N_21155);
nor U27844 (N_27844,N_22472,N_20866);
nor U27845 (N_27845,N_23935,N_23219);
or U27846 (N_27846,N_23022,N_20753);
nor U27847 (N_27847,N_21405,N_21907);
xnor U27848 (N_27848,N_24722,N_23440);
nand U27849 (N_27849,N_22498,N_20008);
and U27850 (N_27850,N_23045,N_22167);
xnor U27851 (N_27851,N_24104,N_22133);
or U27852 (N_27852,N_21712,N_20993);
xnor U27853 (N_27853,N_22181,N_20554);
and U27854 (N_27854,N_22436,N_24737);
nor U27855 (N_27855,N_24331,N_20616);
nor U27856 (N_27856,N_24230,N_23564);
or U27857 (N_27857,N_22001,N_21524);
nand U27858 (N_27858,N_20385,N_21778);
nor U27859 (N_27859,N_22847,N_20525);
nand U27860 (N_27860,N_20549,N_21658);
nor U27861 (N_27861,N_22456,N_22339);
nand U27862 (N_27862,N_24911,N_20948);
nand U27863 (N_27863,N_21822,N_22980);
nor U27864 (N_27864,N_21236,N_23149);
and U27865 (N_27865,N_23172,N_24927);
nor U27866 (N_27866,N_24843,N_20453);
nor U27867 (N_27867,N_24403,N_23671);
nor U27868 (N_27868,N_21816,N_21850);
xor U27869 (N_27869,N_24439,N_24137);
or U27870 (N_27870,N_21032,N_20744);
or U27871 (N_27871,N_24899,N_23193);
and U27872 (N_27872,N_20318,N_24578);
nor U27873 (N_27873,N_22386,N_20448);
or U27874 (N_27874,N_22788,N_20314);
and U27875 (N_27875,N_24069,N_23451);
xor U27876 (N_27876,N_24088,N_20244);
nor U27877 (N_27877,N_21384,N_21176);
nand U27878 (N_27878,N_21533,N_22177);
and U27879 (N_27879,N_24213,N_21857);
or U27880 (N_27880,N_23557,N_24862);
nor U27881 (N_27881,N_20638,N_22516);
nand U27882 (N_27882,N_20820,N_22879);
and U27883 (N_27883,N_20916,N_21927);
nor U27884 (N_27884,N_20989,N_23364);
nor U27885 (N_27885,N_22851,N_20547);
xnor U27886 (N_27886,N_24693,N_23724);
nand U27887 (N_27887,N_21562,N_22129);
xnor U27888 (N_27888,N_21028,N_23642);
nand U27889 (N_27889,N_23171,N_21420);
nor U27890 (N_27890,N_22206,N_21471);
nand U27891 (N_27891,N_24673,N_22093);
xor U27892 (N_27892,N_20893,N_24741);
nor U27893 (N_27893,N_22964,N_21534);
nor U27894 (N_27894,N_21592,N_22011);
or U27895 (N_27895,N_20931,N_22525);
nor U27896 (N_27896,N_22898,N_20659);
xnor U27897 (N_27897,N_20935,N_21841);
or U27898 (N_27898,N_23043,N_22656);
xor U27899 (N_27899,N_24058,N_22466);
nor U27900 (N_27900,N_21715,N_20901);
or U27901 (N_27901,N_24276,N_22294);
or U27902 (N_27902,N_21459,N_24486);
xor U27903 (N_27903,N_22128,N_20639);
and U27904 (N_27904,N_20517,N_23754);
or U27905 (N_27905,N_20687,N_23438);
nand U27906 (N_27906,N_23083,N_22622);
xnor U27907 (N_27907,N_23928,N_23742);
or U27908 (N_27908,N_23218,N_22650);
nand U27909 (N_27909,N_21792,N_20047);
xnor U27910 (N_27910,N_21703,N_22370);
nor U27911 (N_27911,N_22823,N_21113);
nand U27912 (N_27912,N_20914,N_21202);
or U27913 (N_27913,N_24362,N_24531);
nand U27914 (N_27914,N_20942,N_21819);
and U27915 (N_27915,N_23416,N_24593);
nor U27916 (N_27916,N_21258,N_23317);
xor U27917 (N_27917,N_21564,N_23259);
nor U27918 (N_27918,N_20664,N_24436);
nor U27919 (N_27919,N_20840,N_22227);
xor U27920 (N_27920,N_24909,N_24684);
and U27921 (N_27921,N_22643,N_22545);
and U27922 (N_27922,N_20884,N_21796);
and U27923 (N_27923,N_24440,N_22109);
or U27924 (N_27924,N_21816,N_24189);
xor U27925 (N_27925,N_21196,N_21851);
and U27926 (N_27926,N_22997,N_23950);
and U27927 (N_27927,N_24121,N_21718);
nor U27928 (N_27928,N_23506,N_21346);
nand U27929 (N_27929,N_20100,N_24809);
or U27930 (N_27930,N_22045,N_23278);
xor U27931 (N_27931,N_24621,N_20265);
nand U27932 (N_27932,N_23008,N_24775);
nor U27933 (N_27933,N_24508,N_24517);
xor U27934 (N_27934,N_20059,N_21116);
nor U27935 (N_27935,N_20352,N_24261);
xnor U27936 (N_27936,N_23512,N_22189);
nand U27937 (N_27937,N_21494,N_22253);
nor U27938 (N_27938,N_21635,N_20020);
xnor U27939 (N_27939,N_23309,N_24019);
xor U27940 (N_27940,N_21917,N_23965);
or U27941 (N_27941,N_23365,N_21512);
nand U27942 (N_27942,N_22385,N_22829);
or U27943 (N_27943,N_21465,N_20455);
or U27944 (N_27944,N_21954,N_24893);
nand U27945 (N_27945,N_20594,N_24639);
or U27946 (N_27946,N_22437,N_21344);
and U27947 (N_27947,N_22524,N_22883);
nor U27948 (N_27948,N_23993,N_24306);
or U27949 (N_27949,N_23217,N_21631);
and U27950 (N_27950,N_20290,N_21262);
xnor U27951 (N_27951,N_21141,N_22679);
and U27952 (N_27952,N_23499,N_20095);
nand U27953 (N_27953,N_20377,N_20525);
or U27954 (N_27954,N_24034,N_21415);
xor U27955 (N_27955,N_22223,N_20270);
or U27956 (N_27956,N_24741,N_20799);
or U27957 (N_27957,N_24548,N_24642);
nor U27958 (N_27958,N_20435,N_20295);
nor U27959 (N_27959,N_22145,N_20872);
and U27960 (N_27960,N_23093,N_23997);
xor U27961 (N_27961,N_22098,N_24012);
and U27962 (N_27962,N_21754,N_23115);
xnor U27963 (N_27963,N_20945,N_24223);
nand U27964 (N_27964,N_22866,N_24962);
nand U27965 (N_27965,N_21978,N_22426);
nand U27966 (N_27966,N_20930,N_24943);
xor U27967 (N_27967,N_21994,N_20617);
and U27968 (N_27968,N_24800,N_20837);
xor U27969 (N_27969,N_22126,N_21674);
or U27970 (N_27970,N_23951,N_23877);
and U27971 (N_27971,N_20348,N_20461);
xnor U27972 (N_27972,N_21066,N_20332);
or U27973 (N_27973,N_21545,N_23269);
xor U27974 (N_27974,N_24381,N_21787);
xor U27975 (N_27975,N_20876,N_22908);
nor U27976 (N_27976,N_23979,N_24705);
xor U27977 (N_27977,N_24741,N_20651);
nand U27978 (N_27978,N_20983,N_23014);
and U27979 (N_27979,N_24595,N_20315);
or U27980 (N_27980,N_24436,N_24158);
and U27981 (N_27981,N_21419,N_21563);
nor U27982 (N_27982,N_20775,N_24010);
nand U27983 (N_27983,N_22174,N_24330);
and U27984 (N_27984,N_23278,N_24148);
nand U27985 (N_27985,N_21564,N_24396);
nor U27986 (N_27986,N_21097,N_24032);
and U27987 (N_27987,N_23084,N_21318);
nand U27988 (N_27988,N_22215,N_24725);
xor U27989 (N_27989,N_23708,N_20740);
nor U27990 (N_27990,N_23388,N_22164);
xnor U27991 (N_27991,N_21078,N_22994);
and U27992 (N_27992,N_21709,N_20175);
and U27993 (N_27993,N_22239,N_20947);
nand U27994 (N_27994,N_20587,N_21410);
nand U27995 (N_27995,N_23194,N_22079);
xor U27996 (N_27996,N_24767,N_22395);
or U27997 (N_27997,N_24618,N_20132);
nor U27998 (N_27998,N_20277,N_20212);
xor U27999 (N_27999,N_21974,N_22423);
xor U28000 (N_28000,N_24638,N_20702);
and U28001 (N_28001,N_22503,N_21157);
xnor U28002 (N_28002,N_21041,N_21605);
xnor U28003 (N_28003,N_21646,N_23678);
xor U28004 (N_28004,N_24797,N_23668);
nor U28005 (N_28005,N_23479,N_21188);
or U28006 (N_28006,N_23444,N_24894);
xnor U28007 (N_28007,N_21592,N_23476);
nand U28008 (N_28008,N_23607,N_23319);
or U28009 (N_28009,N_21961,N_20010);
and U28010 (N_28010,N_21474,N_22604);
or U28011 (N_28011,N_23898,N_20122);
xor U28012 (N_28012,N_22627,N_22450);
and U28013 (N_28013,N_21296,N_23527);
nand U28014 (N_28014,N_21297,N_24854);
nor U28015 (N_28015,N_21326,N_22063);
or U28016 (N_28016,N_21572,N_20199);
and U28017 (N_28017,N_21656,N_23294);
and U28018 (N_28018,N_23930,N_22290);
or U28019 (N_28019,N_20280,N_24145);
or U28020 (N_28020,N_23262,N_24206);
and U28021 (N_28021,N_20606,N_22781);
or U28022 (N_28022,N_22346,N_21794);
nor U28023 (N_28023,N_23996,N_20355);
nor U28024 (N_28024,N_23548,N_24154);
or U28025 (N_28025,N_24875,N_21156);
nor U28026 (N_28026,N_21399,N_21186);
nor U28027 (N_28027,N_24760,N_22317);
and U28028 (N_28028,N_20749,N_22511);
and U28029 (N_28029,N_24684,N_22833);
nand U28030 (N_28030,N_24699,N_24009);
or U28031 (N_28031,N_20901,N_20523);
and U28032 (N_28032,N_20158,N_24179);
and U28033 (N_28033,N_21103,N_23801);
or U28034 (N_28034,N_20158,N_22610);
or U28035 (N_28035,N_22476,N_20417);
and U28036 (N_28036,N_20271,N_20731);
or U28037 (N_28037,N_23539,N_21698);
nand U28038 (N_28038,N_23803,N_24844);
nor U28039 (N_28039,N_21922,N_24370);
xor U28040 (N_28040,N_21418,N_24334);
or U28041 (N_28041,N_20552,N_24731);
and U28042 (N_28042,N_24246,N_23494);
nand U28043 (N_28043,N_20984,N_23587);
nand U28044 (N_28044,N_21679,N_22503);
nand U28045 (N_28045,N_24227,N_23556);
or U28046 (N_28046,N_21774,N_21024);
and U28047 (N_28047,N_20474,N_24964);
or U28048 (N_28048,N_24212,N_24606);
nand U28049 (N_28049,N_23231,N_24493);
nor U28050 (N_28050,N_23903,N_21854);
nand U28051 (N_28051,N_22666,N_24655);
or U28052 (N_28052,N_23143,N_23021);
and U28053 (N_28053,N_23319,N_24157);
and U28054 (N_28054,N_24840,N_23044);
nor U28055 (N_28055,N_24974,N_21315);
or U28056 (N_28056,N_24587,N_22451);
xor U28057 (N_28057,N_24522,N_20053);
nor U28058 (N_28058,N_23866,N_24347);
nor U28059 (N_28059,N_22710,N_21421);
or U28060 (N_28060,N_21928,N_23392);
or U28061 (N_28061,N_24740,N_24858);
nor U28062 (N_28062,N_23449,N_23202);
nand U28063 (N_28063,N_21203,N_21679);
nor U28064 (N_28064,N_22329,N_21061);
xnor U28065 (N_28065,N_21709,N_20957);
nor U28066 (N_28066,N_22564,N_21355);
nor U28067 (N_28067,N_21751,N_20420);
nor U28068 (N_28068,N_24850,N_22241);
or U28069 (N_28069,N_23616,N_23949);
nand U28070 (N_28070,N_23835,N_20981);
and U28071 (N_28071,N_21966,N_21363);
nor U28072 (N_28072,N_23844,N_23808);
nor U28073 (N_28073,N_22179,N_20269);
or U28074 (N_28074,N_23641,N_21400);
and U28075 (N_28075,N_20211,N_21519);
nand U28076 (N_28076,N_23026,N_23268);
or U28077 (N_28077,N_24725,N_20143);
and U28078 (N_28078,N_23438,N_22248);
xnor U28079 (N_28079,N_20878,N_22401);
and U28080 (N_28080,N_22415,N_23565);
nor U28081 (N_28081,N_20811,N_24479);
and U28082 (N_28082,N_21985,N_23489);
and U28083 (N_28083,N_20348,N_20676);
or U28084 (N_28084,N_23705,N_23090);
and U28085 (N_28085,N_23200,N_20463);
xor U28086 (N_28086,N_21538,N_21566);
and U28087 (N_28087,N_20106,N_22023);
and U28088 (N_28088,N_22371,N_24845);
and U28089 (N_28089,N_24074,N_20337);
or U28090 (N_28090,N_24412,N_23857);
or U28091 (N_28091,N_23662,N_20188);
or U28092 (N_28092,N_23432,N_20551);
nand U28093 (N_28093,N_22482,N_22274);
and U28094 (N_28094,N_22712,N_23055);
xor U28095 (N_28095,N_23141,N_23223);
nor U28096 (N_28096,N_23834,N_21434);
nor U28097 (N_28097,N_23345,N_22352);
nand U28098 (N_28098,N_20658,N_21708);
nand U28099 (N_28099,N_23847,N_21128);
nand U28100 (N_28100,N_24863,N_22814);
and U28101 (N_28101,N_23822,N_23619);
or U28102 (N_28102,N_21183,N_24732);
or U28103 (N_28103,N_23835,N_21912);
or U28104 (N_28104,N_24421,N_24752);
xor U28105 (N_28105,N_24332,N_20333);
xor U28106 (N_28106,N_24477,N_23133);
xnor U28107 (N_28107,N_20233,N_24391);
nand U28108 (N_28108,N_24695,N_21309);
xnor U28109 (N_28109,N_23255,N_21470);
xnor U28110 (N_28110,N_21758,N_23648);
and U28111 (N_28111,N_24473,N_24381);
nor U28112 (N_28112,N_24108,N_22794);
xnor U28113 (N_28113,N_23167,N_20863);
and U28114 (N_28114,N_22046,N_21881);
nand U28115 (N_28115,N_20099,N_23913);
or U28116 (N_28116,N_23058,N_24201);
nor U28117 (N_28117,N_21629,N_22991);
nor U28118 (N_28118,N_21634,N_20902);
nand U28119 (N_28119,N_24437,N_21370);
nor U28120 (N_28120,N_20718,N_22053);
nor U28121 (N_28121,N_22366,N_24899);
or U28122 (N_28122,N_22276,N_24027);
or U28123 (N_28123,N_20594,N_21824);
xnor U28124 (N_28124,N_23497,N_20914);
xor U28125 (N_28125,N_24852,N_23916);
xor U28126 (N_28126,N_22530,N_22121);
xor U28127 (N_28127,N_23243,N_24425);
or U28128 (N_28128,N_20812,N_23039);
and U28129 (N_28129,N_20860,N_24473);
and U28130 (N_28130,N_22815,N_23827);
nor U28131 (N_28131,N_24717,N_21435);
or U28132 (N_28132,N_23620,N_20178);
or U28133 (N_28133,N_20758,N_23881);
xor U28134 (N_28134,N_21490,N_21602);
xnor U28135 (N_28135,N_20063,N_20983);
xor U28136 (N_28136,N_22353,N_23871);
or U28137 (N_28137,N_20398,N_24586);
nand U28138 (N_28138,N_23680,N_22231);
nor U28139 (N_28139,N_22391,N_24601);
xor U28140 (N_28140,N_20351,N_24743);
and U28141 (N_28141,N_21524,N_24615);
and U28142 (N_28142,N_21901,N_24329);
or U28143 (N_28143,N_24530,N_21788);
xor U28144 (N_28144,N_24942,N_21953);
or U28145 (N_28145,N_23116,N_24226);
and U28146 (N_28146,N_23648,N_22342);
nor U28147 (N_28147,N_23066,N_21869);
nand U28148 (N_28148,N_24147,N_20232);
nor U28149 (N_28149,N_20362,N_23967);
nand U28150 (N_28150,N_23081,N_22961);
nor U28151 (N_28151,N_21327,N_23247);
or U28152 (N_28152,N_20958,N_20184);
nand U28153 (N_28153,N_20663,N_23496);
and U28154 (N_28154,N_24214,N_20835);
nor U28155 (N_28155,N_23936,N_20689);
nand U28156 (N_28156,N_20276,N_24249);
or U28157 (N_28157,N_23481,N_23403);
nor U28158 (N_28158,N_22715,N_24516);
or U28159 (N_28159,N_20141,N_22044);
nor U28160 (N_28160,N_20892,N_22561);
and U28161 (N_28161,N_24258,N_21200);
nor U28162 (N_28162,N_23303,N_23165);
or U28163 (N_28163,N_24302,N_22526);
xnor U28164 (N_28164,N_20741,N_20916);
nor U28165 (N_28165,N_24252,N_22650);
and U28166 (N_28166,N_21736,N_20153);
xor U28167 (N_28167,N_23846,N_23673);
or U28168 (N_28168,N_22811,N_24632);
xor U28169 (N_28169,N_20728,N_24765);
or U28170 (N_28170,N_21828,N_22419);
nor U28171 (N_28171,N_24676,N_20546);
and U28172 (N_28172,N_20824,N_21201);
or U28173 (N_28173,N_23476,N_23389);
nand U28174 (N_28174,N_20630,N_22818);
and U28175 (N_28175,N_24134,N_23847);
and U28176 (N_28176,N_21175,N_23650);
or U28177 (N_28177,N_20019,N_21564);
nand U28178 (N_28178,N_23205,N_20109);
and U28179 (N_28179,N_22321,N_20818);
nand U28180 (N_28180,N_22247,N_22876);
xor U28181 (N_28181,N_20182,N_21535);
or U28182 (N_28182,N_20549,N_20849);
nand U28183 (N_28183,N_20363,N_22964);
or U28184 (N_28184,N_21301,N_21557);
nand U28185 (N_28185,N_21308,N_22606);
nor U28186 (N_28186,N_21398,N_22610);
or U28187 (N_28187,N_24478,N_23578);
nand U28188 (N_28188,N_21986,N_24803);
nand U28189 (N_28189,N_21935,N_22579);
and U28190 (N_28190,N_20129,N_24028);
nor U28191 (N_28191,N_20203,N_24818);
or U28192 (N_28192,N_22468,N_22259);
or U28193 (N_28193,N_20084,N_23996);
xor U28194 (N_28194,N_23451,N_20182);
nand U28195 (N_28195,N_21742,N_23272);
nand U28196 (N_28196,N_22496,N_21135);
nand U28197 (N_28197,N_20071,N_22452);
and U28198 (N_28198,N_21255,N_23135);
or U28199 (N_28199,N_20904,N_20354);
nor U28200 (N_28200,N_22278,N_20666);
nand U28201 (N_28201,N_23089,N_24049);
xnor U28202 (N_28202,N_24999,N_24376);
nand U28203 (N_28203,N_20159,N_20271);
nor U28204 (N_28204,N_24978,N_20106);
xor U28205 (N_28205,N_22459,N_23445);
nand U28206 (N_28206,N_23193,N_23469);
nand U28207 (N_28207,N_20301,N_22059);
or U28208 (N_28208,N_21578,N_24470);
xnor U28209 (N_28209,N_21206,N_22279);
or U28210 (N_28210,N_24093,N_20634);
nand U28211 (N_28211,N_20402,N_20525);
nor U28212 (N_28212,N_21137,N_20748);
nand U28213 (N_28213,N_22884,N_22089);
xor U28214 (N_28214,N_22942,N_22779);
and U28215 (N_28215,N_24154,N_23041);
xor U28216 (N_28216,N_22181,N_22894);
xor U28217 (N_28217,N_20133,N_22103);
xnor U28218 (N_28218,N_21307,N_20146);
xnor U28219 (N_28219,N_20864,N_21089);
nand U28220 (N_28220,N_24630,N_20474);
xor U28221 (N_28221,N_22463,N_24227);
xnor U28222 (N_28222,N_24532,N_23928);
xor U28223 (N_28223,N_21941,N_23195);
and U28224 (N_28224,N_22865,N_23313);
nand U28225 (N_28225,N_23712,N_23462);
nor U28226 (N_28226,N_21970,N_22185);
nand U28227 (N_28227,N_22938,N_21836);
or U28228 (N_28228,N_21970,N_23773);
and U28229 (N_28229,N_23164,N_20819);
nand U28230 (N_28230,N_24162,N_24096);
nand U28231 (N_28231,N_20086,N_21074);
and U28232 (N_28232,N_23100,N_22001);
and U28233 (N_28233,N_22643,N_24939);
and U28234 (N_28234,N_23992,N_20224);
nor U28235 (N_28235,N_22525,N_21463);
nand U28236 (N_28236,N_24131,N_22117);
xor U28237 (N_28237,N_20714,N_21422);
or U28238 (N_28238,N_20809,N_23794);
nor U28239 (N_28239,N_21753,N_21999);
nand U28240 (N_28240,N_20086,N_22455);
xor U28241 (N_28241,N_22753,N_20702);
or U28242 (N_28242,N_24188,N_22837);
and U28243 (N_28243,N_22886,N_21919);
or U28244 (N_28244,N_22906,N_23643);
or U28245 (N_28245,N_24555,N_24244);
nor U28246 (N_28246,N_23690,N_20646);
and U28247 (N_28247,N_20215,N_23823);
nor U28248 (N_28248,N_20121,N_20020);
nor U28249 (N_28249,N_21597,N_24227);
nor U28250 (N_28250,N_24420,N_20648);
xor U28251 (N_28251,N_22896,N_24668);
xor U28252 (N_28252,N_23622,N_23357);
xnor U28253 (N_28253,N_22477,N_21563);
nor U28254 (N_28254,N_24577,N_23111);
nand U28255 (N_28255,N_22377,N_24487);
and U28256 (N_28256,N_20781,N_23674);
nand U28257 (N_28257,N_22418,N_24898);
xnor U28258 (N_28258,N_21937,N_21546);
or U28259 (N_28259,N_21881,N_20796);
nand U28260 (N_28260,N_21322,N_24667);
or U28261 (N_28261,N_21983,N_20469);
or U28262 (N_28262,N_21738,N_21908);
and U28263 (N_28263,N_24811,N_24594);
nor U28264 (N_28264,N_21450,N_21242);
or U28265 (N_28265,N_24030,N_24012);
and U28266 (N_28266,N_23069,N_22081);
and U28267 (N_28267,N_21137,N_20600);
xnor U28268 (N_28268,N_23898,N_21289);
or U28269 (N_28269,N_22267,N_24633);
and U28270 (N_28270,N_22944,N_23133);
nor U28271 (N_28271,N_24564,N_24200);
or U28272 (N_28272,N_21306,N_22917);
nand U28273 (N_28273,N_22299,N_22035);
xor U28274 (N_28274,N_24273,N_22355);
and U28275 (N_28275,N_24749,N_22778);
and U28276 (N_28276,N_24722,N_24933);
and U28277 (N_28277,N_24152,N_21346);
nor U28278 (N_28278,N_24159,N_21926);
nor U28279 (N_28279,N_20005,N_24596);
xnor U28280 (N_28280,N_23759,N_21045);
nand U28281 (N_28281,N_21055,N_21992);
nor U28282 (N_28282,N_21292,N_22258);
xnor U28283 (N_28283,N_20707,N_24766);
and U28284 (N_28284,N_20689,N_23517);
nor U28285 (N_28285,N_22966,N_23005);
xor U28286 (N_28286,N_24220,N_23427);
and U28287 (N_28287,N_24229,N_20987);
nand U28288 (N_28288,N_22472,N_20514);
nand U28289 (N_28289,N_20729,N_21174);
nand U28290 (N_28290,N_23611,N_20181);
or U28291 (N_28291,N_23593,N_24787);
xnor U28292 (N_28292,N_22464,N_20825);
nand U28293 (N_28293,N_20741,N_20063);
nor U28294 (N_28294,N_20302,N_22530);
xor U28295 (N_28295,N_20982,N_21967);
and U28296 (N_28296,N_20106,N_20476);
and U28297 (N_28297,N_23498,N_24176);
or U28298 (N_28298,N_22889,N_23229);
or U28299 (N_28299,N_22498,N_23144);
nand U28300 (N_28300,N_24297,N_20862);
and U28301 (N_28301,N_23031,N_22480);
and U28302 (N_28302,N_21201,N_21437);
and U28303 (N_28303,N_24391,N_21087);
or U28304 (N_28304,N_22282,N_22525);
nand U28305 (N_28305,N_20953,N_22617);
xor U28306 (N_28306,N_21744,N_21488);
nand U28307 (N_28307,N_23153,N_20046);
or U28308 (N_28308,N_23879,N_24671);
xnor U28309 (N_28309,N_24464,N_24964);
or U28310 (N_28310,N_22421,N_24838);
nand U28311 (N_28311,N_20866,N_20805);
xnor U28312 (N_28312,N_22117,N_21072);
and U28313 (N_28313,N_22127,N_23857);
xnor U28314 (N_28314,N_23026,N_23244);
xnor U28315 (N_28315,N_24300,N_23379);
or U28316 (N_28316,N_23926,N_22484);
or U28317 (N_28317,N_24421,N_23480);
or U28318 (N_28318,N_21234,N_20448);
and U28319 (N_28319,N_20085,N_23296);
or U28320 (N_28320,N_22428,N_20873);
and U28321 (N_28321,N_20213,N_22915);
nand U28322 (N_28322,N_20112,N_20707);
or U28323 (N_28323,N_23256,N_20691);
nor U28324 (N_28324,N_22590,N_24525);
nor U28325 (N_28325,N_24984,N_21220);
or U28326 (N_28326,N_21439,N_23285);
nor U28327 (N_28327,N_20050,N_20260);
nand U28328 (N_28328,N_23720,N_20089);
nand U28329 (N_28329,N_24981,N_20929);
nand U28330 (N_28330,N_23100,N_22994);
nand U28331 (N_28331,N_21122,N_20162);
nor U28332 (N_28332,N_23026,N_21796);
nor U28333 (N_28333,N_21006,N_23981);
xor U28334 (N_28334,N_20387,N_22516);
nor U28335 (N_28335,N_23826,N_20147);
nor U28336 (N_28336,N_24807,N_20353);
nor U28337 (N_28337,N_23098,N_24208);
xor U28338 (N_28338,N_23124,N_21950);
and U28339 (N_28339,N_21504,N_23303);
nor U28340 (N_28340,N_22877,N_21187);
nand U28341 (N_28341,N_20138,N_23155);
nor U28342 (N_28342,N_24804,N_20215);
or U28343 (N_28343,N_20566,N_21927);
xor U28344 (N_28344,N_23313,N_23884);
or U28345 (N_28345,N_20669,N_21278);
nand U28346 (N_28346,N_23318,N_24865);
or U28347 (N_28347,N_23776,N_24454);
nand U28348 (N_28348,N_20094,N_21998);
nor U28349 (N_28349,N_23454,N_24465);
and U28350 (N_28350,N_21309,N_21534);
nor U28351 (N_28351,N_24424,N_21844);
nor U28352 (N_28352,N_20415,N_24932);
and U28353 (N_28353,N_20278,N_20622);
or U28354 (N_28354,N_23298,N_23020);
xnor U28355 (N_28355,N_24478,N_20842);
xor U28356 (N_28356,N_23925,N_22556);
or U28357 (N_28357,N_24152,N_21609);
nand U28358 (N_28358,N_24177,N_24416);
xnor U28359 (N_28359,N_24920,N_22450);
xnor U28360 (N_28360,N_20931,N_23188);
or U28361 (N_28361,N_20711,N_21683);
or U28362 (N_28362,N_21724,N_20133);
xor U28363 (N_28363,N_20246,N_24465);
or U28364 (N_28364,N_24697,N_22337);
nor U28365 (N_28365,N_21996,N_24523);
nor U28366 (N_28366,N_20128,N_23994);
nor U28367 (N_28367,N_20468,N_20528);
or U28368 (N_28368,N_24404,N_22973);
xnor U28369 (N_28369,N_22126,N_23123);
xnor U28370 (N_28370,N_23268,N_20838);
xnor U28371 (N_28371,N_21333,N_21334);
xnor U28372 (N_28372,N_23547,N_24320);
nor U28373 (N_28373,N_24620,N_21616);
or U28374 (N_28374,N_22550,N_21566);
xor U28375 (N_28375,N_20263,N_22126);
or U28376 (N_28376,N_20844,N_22253);
and U28377 (N_28377,N_23207,N_22667);
xnor U28378 (N_28378,N_22568,N_22271);
xor U28379 (N_28379,N_24004,N_24519);
xnor U28380 (N_28380,N_23771,N_22916);
or U28381 (N_28381,N_20311,N_22568);
and U28382 (N_28382,N_20455,N_20207);
nor U28383 (N_28383,N_21838,N_24196);
nand U28384 (N_28384,N_22693,N_22912);
xor U28385 (N_28385,N_22196,N_22344);
nor U28386 (N_28386,N_22354,N_20446);
and U28387 (N_28387,N_22047,N_24834);
and U28388 (N_28388,N_20833,N_22013);
xnor U28389 (N_28389,N_22516,N_22166);
xnor U28390 (N_28390,N_21635,N_24954);
and U28391 (N_28391,N_22119,N_20400);
or U28392 (N_28392,N_20078,N_22107);
nor U28393 (N_28393,N_21320,N_22940);
or U28394 (N_28394,N_24666,N_20538);
xor U28395 (N_28395,N_23215,N_22175);
xnor U28396 (N_28396,N_21644,N_24034);
or U28397 (N_28397,N_22920,N_22113);
and U28398 (N_28398,N_20510,N_21554);
xnor U28399 (N_28399,N_24354,N_23195);
xor U28400 (N_28400,N_24013,N_20889);
nor U28401 (N_28401,N_24362,N_23896);
or U28402 (N_28402,N_24741,N_23739);
or U28403 (N_28403,N_23148,N_24220);
or U28404 (N_28404,N_22282,N_24800);
xnor U28405 (N_28405,N_21138,N_20256);
and U28406 (N_28406,N_21120,N_21249);
nand U28407 (N_28407,N_20917,N_21725);
and U28408 (N_28408,N_22835,N_24067);
and U28409 (N_28409,N_20598,N_22464);
or U28410 (N_28410,N_24341,N_21256);
or U28411 (N_28411,N_21597,N_22846);
nor U28412 (N_28412,N_23539,N_21130);
nor U28413 (N_28413,N_22119,N_20217);
or U28414 (N_28414,N_20417,N_23481);
and U28415 (N_28415,N_24215,N_22887);
nor U28416 (N_28416,N_23771,N_22868);
and U28417 (N_28417,N_20728,N_20158);
nor U28418 (N_28418,N_24447,N_22642);
nor U28419 (N_28419,N_23222,N_20318);
or U28420 (N_28420,N_23550,N_22866);
or U28421 (N_28421,N_20386,N_22798);
nand U28422 (N_28422,N_24230,N_23830);
nor U28423 (N_28423,N_24812,N_24723);
nor U28424 (N_28424,N_22661,N_22359);
or U28425 (N_28425,N_23795,N_22450);
or U28426 (N_28426,N_22846,N_20857);
nand U28427 (N_28427,N_23384,N_21040);
and U28428 (N_28428,N_20518,N_20894);
nor U28429 (N_28429,N_21349,N_22134);
nor U28430 (N_28430,N_23190,N_22272);
xor U28431 (N_28431,N_20261,N_20387);
nand U28432 (N_28432,N_23750,N_22977);
and U28433 (N_28433,N_24322,N_23485);
nor U28434 (N_28434,N_20752,N_24238);
xnor U28435 (N_28435,N_23886,N_20601);
nor U28436 (N_28436,N_21110,N_23257);
and U28437 (N_28437,N_21631,N_20442);
xnor U28438 (N_28438,N_23892,N_24721);
and U28439 (N_28439,N_21608,N_23037);
and U28440 (N_28440,N_20015,N_20637);
or U28441 (N_28441,N_24952,N_21778);
nand U28442 (N_28442,N_22097,N_24195);
and U28443 (N_28443,N_20301,N_22474);
nor U28444 (N_28444,N_23713,N_24105);
and U28445 (N_28445,N_24561,N_22956);
nand U28446 (N_28446,N_20230,N_23339);
nand U28447 (N_28447,N_22717,N_24160);
nand U28448 (N_28448,N_21123,N_23223);
nand U28449 (N_28449,N_23663,N_24559);
and U28450 (N_28450,N_24717,N_20792);
and U28451 (N_28451,N_21200,N_20269);
or U28452 (N_28452,N_21523,N_20463);
xor U28453 (N_28453,N_20873,N_24909);
and U28454 (N_28454,N_20689,N_23157);
xor U28455 (N_28455,N_22147,N_23520);
and U28456 (N_28456,N_22774,N_24413);
and U28457 (N_28457,N_20415,N_21395);
xor U28458 (N_28458,N_23697,N_24508);
nor U28459 (N_28459,N_20142,N_20830);
and U28460 (N_28460,N_24639,N_21884);
or U28461 (N_28461,N_23859,N_20006);
nor U28462 (N_28462,N_20892,N_21701);
or U28463 (N_28463,N_21478,N_23854);
or U28464 (N_28464,N_24894,N_23726);
nand U28465 (N_28465,N_22022,N_24257);
xnor U28466 (N_28466,N_22472,N_24436);
or U28467 (N_28467,N_20419,N_24550);
xor U28468 (N_28468,N_22358,N_24208);
xor U28469 (N_28469,N_23328,N_20890);
or U28470 (N_28470,N_23641,N_23704);
nor U28471 (N_28471,N_21821,N_22429);
or U28472 (N_28472,N_23439,N_20251);
or U28473 (N_28473,N_20050,N_23778);
or U28474 (N_28474,N_24577,N_24285);
and U28475 (N_28475,N_20596,N_21003);
or U28476 (N_28476,N_21763,N_23745);
xnor U28477 (N_28477,N_24204,N_22109);
xnor U28478 (N_28478,N_21627,N_22798);
xor U28479 (N_28479,N_20749,N_21177);
xnor U28480 (N_28480,N_21580,N_24594);
nand U28481 (N_28481,N_23352,N_23221);
or U28482 (N_28482,N_23978,N_24266);
nor U28483 (N_28483,N_20333,N_21132);
or U28484 (N_28484,N_24304,N_21044);
nor U28485 (N_28485,N_21476,N_22833);
nor U28486 (N_28486,N_20676,N_20444);
xor U28487 (N_28487,N_20204,N_22528);
or U28488 (N_28488,N_22537,N_22199);
xor U28489 (N_28489,N_22647,N_20486);
nor U28490 (N_28490,N_20544,N_21823);
and U28491 (N_28491,N_23181,N_22787);
or U28492 (N_28492,N_23322,N_20941);
or U28493 (N_28493,N_23346,N_21252);
nand U28494 (N_28494,N_23790,N_24944);
xor U28495 (N_28495,N_20137,N_20845);
nor U28496 (N_28496,N_20410,N_23190);
nor U28497 (N_28497,N_23826,N_22100);
nand U28498 (N_28498,N_24801,N_20772);
or U28499 (N_28499,N_21432,N_21784);
and U28500 (N_28500,N_21812,N_20264);
or U28501 (N_28501,N_20442,N_23958);
and U28502 (N_28502,N_22732,N_24053);
or U28503 (N_28503,N_24156,N_24099);
nand U28504 (N_28504,N_21559,N_20385);
nor U28505 (N_28505,N_20575,N_20668);
or U28506 (N_28506,N_20689,N_24561);
nor U28507 (N_28507,N_24457,N_23324);
nor U28508 (N_28508,N_23773,N_23761);
xor U28509 (N_28509,N_20081,N_23896);
and U28510 (N_28510,N_22710,N_23652);
or U28511 (N_28511,N_21934,N_23804);
nor U28512 (N_28512,N_23166,N_21471);
and U28513 (N_28513,N_21541,N_20690);
xnor U28514 (N_28514,N_23907,N_20255);
xor U28515 (N_28515,N_23864,N_22313);
and U28516 (N_28516,N_23920,N_22517);
nand U28517 (N_28517,N_24742,N_21168);
nor U28518 (N_28518,N_20503,N_23701);
or U28519 (N_28519,N_23724,N_24830);
nand U28520 (N_28520,N_23018,N_23876);
nand U28521 (N_28521,N_22498,N_24394);
nor U28522 (N_28522,N_22702,N_20290);
nand U28523 (N_28523,N_22286,N_24212);
and U28524 (N_28524,N_23693,N_21943);
or U28525 (N_28525,N_23643,N_20695);
xor U28526 (N_28526,N_22819,N_24314);
and U28527 (N_28527,N_24549,N_20058);
or U28528 (N_28528,N_21960,N_22456);
xor U28529 (N_28529,N_24950,N_23573);
or U28530 (N_28530,N_22976,N_24974);
xor U28531 (N_28531,N_22055,N_24947);
nor U28532 (N_28532,N_21542,N_24500);
and U28533 (N_28533,N_21252,N_24622);
and U28534 (N_28534,N_21231,N_20704);
nand U28535 (N_28535,N_24974,N_23471);
and U28536 (N_28536,N_24743,N_21243);
or U28537 (N_28537,N_24232,N_22086);
xnor U28538 (N_28538,N_24739,N_24352);
nor U28539 (N_28539,N_22733,N_22627);
nor U28540 (N_28540,N_22984,N_23772);
nor U28541 (N_28541,N_23047,N_24602);
and U28542 (N_28542,N_20377,N_23425);
nand U28543 (N_28543,N_22874,N_22442);
nor U28544 (N_28544,N_23274,N_21687);
and U28545 (N_28545,N_20127,N_20839);
nand U28546 (N_28546,N_22864,N_22520);
nor U28547 (N_28547,N_22469,N_23317);
xnor U28548 (N_28548,N_21206,N_21566);
nand U28549 (N_28549,N_24146,N_22323);
nor U28550 (N_28550,N_22362,N_24298);
nor U28551 (N_28551,N_24166,N_24232);
nor U28552 (N_28552,N_21506,N_20956);
and U28553 (N_28553,N_20010,N_21318);
xnor U28554 (N_28554,N_22283,N_24224);
and U28555 (N_28555,N_23643,N_22175);
nor U28556 (N_28556,N_23456,N_21440);
and U28557 (N_28557,N_24418,N_22651);
or U28558 (N_28558,N_23349,N_20790);
nor U28559 (N_28559,N_20327,N_21761);
xnor U28560 (N_28560,N_20243,N_23052);
xnor U28561 (N_28561,N_22665,N_21193);
or U28562 (N_28562,N_20331,N_20872);
or U28563 (N_28563,N_21764,N_21275);
nor U28564 (N_28564,N_22606,N_24435);
nand U28565 (N_28565,N_22443,N_24919);
nor U28566 (N_28566,N_22919,N_21213);
xor U28567 (N_28567,N_20838,N_20481);
or U28568 (N_28568,N_24329,N_22750);
nor U28569 (N_28569,N_21116,N_21756);
nand U28570 (N_28570,N_22159,N_23677);
nand U28571 (N_28571,N_23151,N_22622);
nor U28572 (N_28572,N_20018,N_22217);
or U28573 (N_28573,N_20033,N_22295);
nor U28574 (N_28574,N_23482,N_21914);
xnor U28575 (N_28575,N_24089,N_24898);
nand U28576 (N_28576,N_20872,N_24659);
nand U28577 (N_28577,N_24797,N_21113);
and U28578 (N_28578,N_24715,N_21975);
nand U28579 (N_28579,N_21452,N_22790);
and U28580 (N_28580,N_21424,N_23455);
and U28581 (N_28581,N_23334,N_21046);
or U28582 (N_28582,N_21993,N_22629);
or U28583 (N_28583,N_20657,N_22715);
and U28584 (N_28584,N_21932,N_20976);
and U28585 (N_28585,N_24906,N_21765);
nand U28586 (N_28586,N_20482,N_22174);
xor U28587 (N_28587,N_22292,N_24593);
xor U28588 (N_28588,N_22811,N_24391);
nor U28589 (N_28589,N_23650,N_21647);
xnor U28590 (N_28590,N_21904,N_22012);
or U28591 (N_28591,N_24357,N_21826);
and U28592 (N_28592,N_24250,N_21189);
nand U28593 (N_28593,N_24220,N_20412);
and U28594 (N_28594,N_21086,N_23809);
and U28595 (N_28595,N_22914,N_24164);
nor U28596 (N_28596,N_23690,N_24035);
xnor U28597 (N_28597,N_24028,N_22061);
nor U28598 (N_28598,N_23363,N_23695);
and U28599 (N_28599,N_24957,N_21908);
xor U28600 (N_28600,N_24512,N_21947);
nand U28601 (N_28601,N_22504,N_23295);
xnor U28602 (N_28602,N_23544,N_20033);
xnor U28603 (N_28603,N_21730,N_22588);
nor U28604 (N_28604,N_24735,N_21361);
nor U28605 (N_28605,N_22637,N_22083);
xnor U28606 (N_28606,N_24856,N_24699);
nor U28607 (N_28607,N_22314,N_24458);
xnor U28608 (N_28608,N_20294,N_20441);
nor U28609 (N_28609,N_20852,N_21697);
nand U28610 (N_28610,N_22220,N_21651);
nand U28611 (N_28611,N_21396,N_20089);
and U28612 (N_28612,N_21418,N_22091);
nand U28613 (N_28613,N_22100,N_21293);
nand U28614 (N_28614,N_24946,N_24741);
nand U28615 (N_28615,N_21984,N_22632);
xor U28616 (N_28616,N_21898,N_24215);
nand U28617 (N_28617,N_24133,N_24202);
and U28618 (N_28618,N_23238,N_24822);
nor U28619 (N_28619,N_20301,N_24292);
nand U28620 (N_28620,N_23506,N_23548);
xnor U28621 (N_28621,N_21566,N_23518);
nor U28622 (N_28622,N_23673,N_21250);
or U28623 (N_28623,N_22519,N_23527);
nor U28624 (N_28624,N_22159,N_20171);
nand U28625 (N_28625,N_22708,N_24556);
or U28626 (N_28626,N_20389,N_20982);
nor U28627 (N_28627,N_20142,N_24062);
nor U28628 (N_28628,N_22683,N_22317);
nand U28629 (N_28629,N_20826,N_24728);
or U28630 (N_28630,N_24835,N_20266);
and U28631 (N_28631,N_21347,N_22838);
and U28632 (N_28632,N_22530,N_22162);
and U28633 (N_28633,N_24808,N_22242);
nand U28634 (N_28634,N_22021,N_20443);
nand U28635 (N_28635,N_21745,N_23294);
xor U28636 (N_28636,N_20039,N_23673);
xnor U28637 (N_28637,N_24472,N_21980);
nand U28638 (N_28638,N_24641,N_22686);
or U28639 (N_28639,N_22456,N_24075);
nor U28640 (N_28640,N_22867,N_24932);
nor U28641 (N_28641,N_24197,N_20527);
xor U28642 (N_28642,N_24593,N_23795);
nor U28643 (N_28643,N_21334,N_24836);
nor U28644 (N_28644,N_22983,N_22559);
nor U28645 (N_28645,N_24569,N_23624);
nand U28646 (N_28646,N_22163,N_20039);
nor U28647 (N_28647,N_23960,N_22422);
nand U28648 (N_28648,N_22754,N_22667);
nor U28649 (N_28649,N_22229,N_23311);
xnor U28650 (N_28650,N_22600,N_20787);
and U28651 (N_28651,N_22525,N_24832);
xor U28652 (N_28652,N_22631,N_24955);
nor U28653 (N_28653,N_21079,N_22495);
nand U28654 (N_28654,N_23080,N_23251);
xor U28655 (N_28655,N_22755,N_24688);
nand U28656 (N_28656,N_23628,N_21025);
and U28657 (N_28657,N_23263,N_22258);
or U28658 (N_28658,N_20239,N_20037);
and U28659 (N_28659,N_22587,N_21663);
xor U28660 (N_28660,N_23158,N_21882);
or U28661 (N_28661,N_23641,N_22425);
or U28662 (N_28662,N_22129,N_23100);
nor U28663 (N_28663,N_24260,N_23804);
xor U28664 (N_28664,N_23448,N_20476);
xnor U28665 (N_28665,N_20391,N_23995);
or U28666 (N_28666,N_24909,N_24661);
nand U28667 (N_28667,N_21710,N_20499);
nor U28668 (N_28668,N_23701,N_20591);
nand U28669 (N_28669,N_23613,N_22172);
or U28670 (N_28670,N_20858,N_21001);
xor U28671 (N_28671,N_24743,N_22858);
nor U28672 (N_28672,N_23613,N_23658);
nand U28673 (N_28673,N_24564,N_23039);
or U28674 (N_28674,N_20239,N_24185);
and U28675 (N_28675,N_24181,N_22077);
and U28676 (N_28676,N_22907,N_23088);
xor U28677 (N_28677,N_23255,N_21879);
nand U28678 (N_28678,N_23442,N_21944);
xnor U28679 (N_28679,N_22358,N_20420);
nand U28680 (N_28680,N_21710,N_21769);
xnor U28681 (N_28681,N_23623,N_22464);
nand U28682 (N_28682,N_22397,N_24789);
and U28683 (N_28683,N_20869,N_23097);
and U28684 (N_28684,N_22196,N_21195);
nor U28685 (N_28685,N_23269,N_23793);
or U28686 (N_28686,N_23409,N_24343);
xnor U28687 (N_28687,N_23926,N_24964);
nor U28688 (N_28688,N_22151,N_24563);
xnor U28689 (N_28689,N_24386,N_21953);
nand U28690 (N_28690,N_23663,N_21283);
nand U28691 (N_28691,N_21927,N_22072);
and U28692 (N_28692,N_24057,N_24431);
nor U28693 (N_28693,N_24388,N_22745);
nor U28694 (N_28694,N_20454,N_22009);
nand U28695 (N_28695,N_24221,N_23996);
or U28696 (N_28696,N_23195,N_21113);
or U28697 (N_28697,N_23082,N_21645);
and U28698 (N_28698,N_22487,N_22948);
nor U28699 (N_28699,N_21943,N_22485);
xnor U28700 (N_28700,N_20498,N_23926);
nor U28701 (N_28701,N_21480,N_23615);
nand U28702 (N_28702,N_20304,N_24172);
nor U28703 (N_28703,N_24140,N_20599);
nand U28704 (N_28704,N_23669,N_20125);
nor U28705 (N_28705,N_20239,N_23091);
nor U28706 (N_28706,N_21037,N_21635);
nor U28707 (N_28707,N_22826,N_20794);
or U28708 (N_28708,N_21062,N_24757);
xor U28709 (N_28709,N_22563,N_23305);
nor U28710 (N_28710,N_23177,N_22484);
xnor U28711 (N_28711,N_21238,N_21839);
xor U28712 (N_28712,N_24780,N_23087);
nor U28713 (N_28713,N_23246,N_21063);
xor U28714 (N_28714,N_22781,N_23161);
nand U28715 (N_28715,N_23170,N_24724);
nand U28716 (N_28716,N_20352,N_24489);
xnor U28717 (N_28717,N_22391,N_22038);
or U28718 (N_28718,N_24831,N_23299);
or U28719 (N_28719,N_24037,N_24351);
or U28720 (N_28720,N_23401,N_20705);
nor U28721 (N_28721,N_24108,N_22636);
and U28722 (N_28722,N_22817,N_24536);
nand U28723 (N_28723,N_23521,N_24110);
and U28724 (N_28724,N_23899,N_20205);
xnor U28725 (N_28725,N_21858,N_21637);
nand U28726 (N_28726,N_23047,N_23635);
and U28727 (N_28727,N_22301,N_22006);
or U28728 (N_28728,N_22944,N_23551);
and U28729 (N_28729,N_20826,N_24514);
nor U28730 (N_28730,N_24090,N_23819);
and U28731 (N_28731,N_20816,N_21759);
and U28732 (N_28732,N_24083,N_24823);
nand U28733 (N_28733,N_22269,N_20844);
nand U28734 (N_28734,N_22719,N_22521);
nor U28735 (N_28735,N_22383,N_23939);
or U28736 (N_28736,N_23728,N_22099);
nor U28737 (N_28737,N_21706,N_24114);
nand U28738 (N_28738,N_22699,N_21219);
or U28739 (N_28739,N_21490,N_20547);
or U28740 (N_28740,N_22675,N_20807);
xor U28741 (N_28741,N_23916,N_21813);
xor U28742 (N_28742,N_21009,N_22060);
nand U28743 (N_28743,N_21447,N_20614);
nand U28744 (N_28744,N_22623,N_23907);
nor U28745 (N_28745,N_21116,N_21150);
or U28746 (N_28746,N_22442,N_23430);
or U28747 (N_28747,N_22786,N_23204);
or U28748 (N_28748,N_20712,N_24877);
nor U28749 (N_28749,N_23074,N_23140);
xnor U28750 (N_28750,N_22018,N_23143);
xor U28751 (N_28751,N_23683,N_20579);
nor U28752 (N_28752,N_20759,N_23307);
nor U28753 (N_28753,N_20438,N_23149);
nand U28754 (N_28754,N_23470,N_21626);
nor U28755 (N_28755,N_22914,N_20170);
or U28756 (N_28756,N_22971,N_21287);
and U28757 (N_28757,N_22311,N_20208);
and U28758 (N_28758,N_21797,N_24097);
xnor U28759 (N_28759,N_21205,N_21000);
nor U28760 (N_28760,N_23154,N_24581);
nand U28761 (N_28761,N_22108,N_23860);
nand U28762 (N_28762,N_20168,N_23344);
nand U28763 (N_28763,N_24883,N_21832);
nand U28764 (N_28764,N_22128,N_24982);
nand U28765 (N_28765,N_20818,N_20873);
nor U28766 (N_28766,N_24469,N_23538);
nand U28767 (N_28767,N_24581,N_21292);
or U28768 (N_28768,N_22622,N_23087);
nand U28769 (N_28769,N_21920,N_20285);
or U28770 (N_28770,N_20614,N_22031);
nand U28771 (N_28771,N_21055,N_20575);
nand U28772 (N_28772,N_24280,N_21044);
and U28773 (N_28773,N_24831,N_24274);
and U28774 (N_28774,N_20039,N_21066);
xnor U28775 (N_28775,N_22347,N_24005);
or U28776 (N_28776,N_24411,N_24246);
nand U28777 (N_28777,N_22942,N_23119);
nand U28778 (N_28778,N_23460,N_23913);
xnor U28779 (N_28779,N_21791,N_23860);
nand U28780 (N_28780,N_24988,N_24361);
and U28781 (N_28781,N_23736,N_22978);
nand U28782 (N_28782,N_23722,N_23384);
and U28783 (N_28783,N_21652,N_20026);
or U28784 (N_28784,N_21169,N_21208);
nand U28785 (N_28785,N_21059,N_22745);
or U28786 (N_28786,N_22909,N_24610);
and U28787 (N_28787,N_22769,N_24127);
or U28788 (N_28788,N_24033,N_22816);
xor U28789 (N_28789,N_20489,N_24490);
or U28790 (N_28790,N_23020,N_24766);
nand U28791 (N_28791,N_21174,N_20544);
and U28792 (N_28792,N_23396,N_23793);
nand U28793 (N_28793,N_22075,N_21076);
xnor U28794 (N_28794,N_24741,N_23814);
or U28795 (N_28795,N_23866,N_24527);
or U28796 (N_28796,N_24679,N_24105);
and U28797 (N_28797,N_20998,N_24945);
nand U28798 (N_28798,N_24935,N_20799);
and U28799 (N_28799,N_21497,N_21953);
or U28800 (N_28800,N_20066,N_24004);
or U28801 (N_28801,N_21221,N_21937);
or U28802 (N_28802,N_23606,N_20307);
or U28803 (N_28803,N_24790,N_20350);
nand U28804 (N_28804,N_23026,N_22370);
and U28805 (N_28805,N_22043,N_23734);
xnor U28806 (N_28806,N_20566,N_24795);
nand U28807 (N_28807,N_24236,N_24419);
or U28808 (N_28808,N_24932,N_24976);
nor U28809 (N_28809,N_21024,N_24399);
xor U28810 (N_28810,N_23411,N_24130);
and U28811 (N_28811,N_23000,N_21747);
or U28812 (N_28812,N_20567,N_20672);
or U28813 (N_28813,N_21297,N_20161);
xnor U28814 (N_28814,N_22265,N_20818);
xor U28815 (N_28815,N_23075,N_20369);
or U28816 (N_28816,N_20934,N_20097);
xor U28817 (N_28817,N_21994,N_23762);
or U28818 (N_28818,N_22853,N_23007);
and U28819 (N_28819,N_23036,N_23926);
and U28820 (N_28820,N_20078,N_20460);
nor U28821 (N_28821,N_20488,N_21397);
xnor U28822 (N_28822,N_20218,N_20889);
or U28823 (N_28823,N_24989,N_22336);
xnor U28824 (N_28824,N_20802,N_22285);
nand U28825 (N_28825,N_20333,N_20859);
xnor U28826 (N_28826,N_21825,N_24336);
nand U28827 (N_28827,N_22634,N_24080);
xor U28828 (N_28828,N_20385,N_24494);
nor U28829 (N_28829,N_24573,N_23962);
nand U28830 (N_28830,N_22187,N_21409);
or U28831 (N_28831,N_23020,N_23562);
or U28832 (N_28832,N_21638,N_21269);
nor U28833 (N_28833,N_24559,N_22719);
nand U28834 (N_28834,N_24366,N_22748);
xor U28835 (N_28835,N_22289,N_23658);
xor U28836 (N_28836,N_24180,N_23788);
xnor U28837 (N_28837,N_24384,N_21793);
xor U28838 (N_28838,N_22562,N_24512);
nor U28839 (N_28839,N_24619,N_24102);
xor U28840 (N_28840,N_21604,N_24349);
and U28841 (N_28841,N_23437,N_22607);
nand U28842 (N_28842,N_24378,N_23808);
nand U28843 (N_28843,N_22580,N_22779);
and U28844 (N_28844,N_21413,N_20501);
nand U28845 (N_28845,N_20094,N_21328);
nand U28846 (N_28846,N_23058,N_22099);
nor U28847 (N_28847,N_20867,N_22640);
nand U28848 (N_28848,N_23946,N_23534);
or U28849 (N_28849,N_23895,N_24643);
xnor U28850 (N_28850,N_22274,N_20600);
nor U28851 (N_28851,N_20369,N_23029);
nor U28852 (N_28852,N_24297,N_24475);
and U28853 (N_28853,N_21750,N_20012);
xor U28854 (N_28854,N_23947,N_20170);
and U28855 (N_28855,N_22124,N_23036);
or U28856 (N_28856,N_23589,N_23731);
or U28857 (N_28857,N_24140,N_24176);
xor U28858 (N_28858,N_24716,N_21963);
xnor U28859 (N_28859,N_20900,N_23841);
nor U28860 (N_28860,N_23692,N_21443);
or U28861 (N_28861,N_24940,N_21231);
nor U28862 (N_28862,N_21641,N_20767);
and U28863 (N_28863,N_22911,N_23588);
xor U28864 (N_28864,N_24674,N_21323);
nand U28865 (N_28865,N_23680,N_22001);
and U28866 (N_28866,N_20017,N_22720);
nand U28867 (N_28867,N_24787,N_23835);
nand U28868 (N_28868,N_22940,N_23250);
or U28869 (N_28869,N_22491,N_23295);
nand U28870 (N_28870,N_22293,N_22735);
or U28871 (N_28871,N_20617,N_21531);
xnor U28872 (N_28872,N_20632,N_24192);
or U28873 (N_28873,N_23152,N_24329);
and U28874 (N_28874,N_24646,N_21803);
or U28875 (N_28875,N_23152,N_22508);
nand U28876 (N_28876,N_24025,N_22258);
and U28877 (N_28877,N_22609,N_21572);
nand U28878 (N_28878,N_20135,N_22500);
nand U28879 (N_28879,N_22530,N_22206);
nand U28880 (N_28880,N_21904,N_24365);
and U28881 (N_28881,N_22500,N_24432);
or U28882 (N_28882,N_22214,N_23253);
nor U28883 (N_28883,N_20078,N_24445);
xnor U28884 (N_28884,N_23475,N_22837);
or U28885 (N_28885,N_23086,N_23385);
and U28886 (N_28886,N_24832,N_21608);
or U28887 (N_28887,N_22848,N_21959);
or U28888 (N_28888,N_21702,N_22099);
nor U28889 (N_28889,N_23076,N_24293);
nor U28890 (N_28890,N_22498,N_22630);
nor U28891 (N_28891,N_24167,N_24569);
and U28892 (N_28892,N_23785,N_21158);
nand U28893 (N_28893,N_23283,N_20010);
xor U28894 (N_28894,N_23165,N_24601);
or U28895 (N_28895,N_21367,N_24338);
and U28896 (N_28896,N_23760,N_22626);
nand U28897 (N_28897,N_22048,N_21958);
and U28898 (N_28898,N_22167,N_24524);
and U28899 (N_28899,N_23278,N_24112);
nor U28900 (N_28900,N_22851,N_22123);
and U28901 (N_28901,N_23812,N_20238);
and U28902 (N_28902,N_21129,N_20488);
xnor U28903 (N_28903,N_21302,N_24531);
nand U28904 (N_28904,N_21590,N_20243);
and U28905 (N_28905,N_21804,N_23109);
and U28906 (N_28906,N_23398,N_23723);
nor U28907 (N_28907,N_20279,N_23812);
xnor U28908 (N_28908,N_20237,N_20006);
nor U28909 (N_28909,N_24564,N_24818);
nand U28910 (N_28910,N_21950,N_21368);
nand U28911 (N_28911,N_21140,N_21398);
or U28912 (N_28912,N_20791,N_24048);
or U28913 (N_28913,N_21368,N_22836);
nor U28914 (N_28914,N_21187,N_20651);
nor U28915 (N_28915,N_22819,N_20628);
xnor U28916 (N_28916,N_24262,N_23831);
and U28917 (N_28917,N_20088,N_20831);
nand U28918 (N_28918,N_20281,N_24021);
nand U28919 (N_28919,N_21816,N_23423);
xor U28920 (N_28920,N_21556,N_22974);
and U28921 (N_28921,N_21337,N_23617);
xor U28922 (N_28922,N_21558,N_22795);
nor U28923 (N_28923,N_21212,N_22542);
xor U28924 (N_28924,N_21104,N_20581);
xor U28925 (N_28925,N_24483,N_21391);
nor U28926 (N_28926,N_21317,N_20246);
nor U28927 (N_28927,N_23258,N_23414);
or U28928 (N_28928,N_22919,N_21200);
xnor U28929 (N_28929,N_24080,N_23672);
xnor U28930 (N_28930,N_22549,N_21187);
or U28931 (N_28931,N_22704,N_24392);
and U28932 (N_28932,N_23893,N_23105);
or U28933 (N_28933,N_22183,N_22740);
and U28934 (N_28934,N_21674,N_23306);
nand U28935 (N_28935,N_20274,N_21098);
xnor U28936 (N_28936,N_21870,N_22413);
nand U28937 (N_28937,N_22392,N_24960);
nand U28938 (N_28938,N_22947,N_20596);
xor U28939 (N_28939,N_23808,N_21739);
xnor U28940 (N_28940,N_23230,N_23353);
nand U28941 (N_28941,N_24004,N_23151);
or U28942 (N_28942,N_21247,N_22906);
nor U28943 (N_28943,N_23176,N_20304);
or U28944 (N_28944,N_20467,N_20659);
nand U28945 (N_28945,N_24275,N_20531);
xnor U28946 (N_28946,N_20417,N_21535);
and U28947 (N_28947,N_20470,N_20969);
and U28948 (N_28948,N_21412,N_23526);
and U28949 (N_28949,N_23038,N_20992);
nor U28950 (N_28950,N_21802,N_20540);
or U28951 (N_28951,N_23255,N_22990);
and U28952 (N_28952,N_22326,N_24041);
and U28953 (N_28953,N_23420,N_21533);
or U28954 (N_28954,N_20996,N_22987);
and U28955 (N_28955,N_21519,N_20473);
nand U28956 (N_28956,N_21703,N_21523);
nand U28957 (N_28957,N_24470,N_20911);
and U28958 (N_28958,N_20492,N_21405);
and U28959 (N_28959,N_20539,N_23235);
nor U28960 (N_28960,N_23700,N_22221);
xor U28961 (N_28961,N_23686,N_21009);
and U28962 (N_28962,N_22920,N_21482);
nor U28963 (N_28963,N_24781,N_24873);
nor U28964 (N_28964,N_20917,N_20043);
and U28965 (N_28965,N_23117,N_21315);
or U28966 (N_28966,N_22004,N_24630);
xnor U28967 (N_28967,N_22215,N_20814);
nand U28968 (N_28968,N_22362,N_24620);
xnor U28969 (N_28969,N_24871,N_22734);
nor U28970 (N_28970,N_24511,N_20404);
nor U28971 (N_28971,N_20458,N_22276);
xnor U28972 (N_28972,N_21114,N_20476);
and U28973 (N_28973,N_20599,N_21955);
nor U28974 (N_28974,N_24004,N_24432);
xnor U28975 (N_28975,N_22054,N_20225);
or U28976 (N_28976,N_20074,N_24406);
xnor U28977 (N_28977,N_21133,N_21681);
xor U28978 (N_28978,N_24959,N_21362);
xnor U28979 (N_28979,N_21119,N_21403);
xor U28980 (N_28980,N_23111,N_24795);
nor U28981 (N_28981,N_21654,N_24147);
nand U28982 (N_28982,N_22028,N_20791);
and U28983 (N_28983,N_23700,N_24852);
nand U28984 (N_28984,N_22601,N_23476);
nor U28985 (N_28985,N_23082,N_24537);
and U28986 (N_28986,N_23326,N_24519);
nand U28987 (N_28987,N_22155,N_22676);
nor U28988 (N_28988,N_20061,N_22260);
and U28989 (N_28989,N_23438,N_21407);
and U28990 (N_28990,N_23527,N_23763);
nor U28991 (N_28991,N_24746,N_21605);
xor U28992 (N_28992,N_24705,N_24593);
and U28993 (N_28993,N_23671,N_22306);
and U28994 (N_28994,N_23763,N_20021);
or U28995 (N_28995,N_20579,N_23836);
nor U28996 (N_28996,N_24480,N_20622);
nand U28997 (N_28997,N_21304,N_23502);
xor U28998 (N_28998,N_22677,N_23672);
xnor U28999 (N_28999,N_24073,N_22221);
and U29000 (N_29000,N_20781,N_20280);
nor U29001 (N_29001,N_20580,N_22843);
or U29002 (N_29002,N_24948,N_24087);
and U29003 (N_29003,N_20545,N_24045);
xor U29004 (N_29004,N_24024,N_21118);
xor U29005 (N_29005,N_23749,N_23229);
xnor U29006 (N_29006,N_22115,N_24279);
nand U29007 (N_29007,N_22790,N_20618);
nand U29008 (N_29008,N_20465,N_21670);
nand U29009 (N_29009,N_24986,N_21236);
nand U29010 (N_29010,N_21822,N_24613);
xnor U29011 (N_29011,N_22781,N_22598);
nor U29012 (N_29012,N_20713,N_23163);
and U29013 (N_29013,N_22554,N_24516);
or U29014 (N_29014,N_20947,N_20283);
nor U29015 (N_29015,N_20366,N_23881);
xnor U29016 (N_29016,N_21213,N_22647);
and U29017 (N_29017,N_23888,N_20473);
and U29018 (N_29018,N_24889,N_21598);
nor U29019 (N_29019,N_20092,N_22504);
or U29020 (N_29020,N_21857,N_24016);
xnor U29021 (N_29021,N_21414,N_23154);
xnor U29022 (N_29022,N_24709,N_22390);
xnor U29023 (N_29023,N_20067,N_20608);
xor U29024 (N_29024,N_22296,N_23445);
xor U29025 (N_29025,N_23616,N_20739);
and U29026 (N_29026,N_24754,N_23787);
and U29027 (N_29027,N_24923,N_24241);
nor U29028 (N_29028,N_23762,N_22408);
or U29029 (N_29029,N_20099,N_21945);
nor U29030 (N_29030,N_21009,N_23479);
or U29031 (N_29031,N_24479,N_24461);
nor U29032 (N_29032,N_20723,N_24538);
nand U29033 (N_29033,N_20518,N_20207);
and U29034 (N_29034,N_20247,N_20179);
or U29035 (N_29035,N_20558,N_22380);
xor U29036 (N_29036,N_22932,N_22419);
and U29037 (N_29037,N_20952,N_23785);
xor U29038 (N_29038,N_20393,N_23115);
nand U29039 (N_29039,N_20237,N_24566);
nand U29040 (N_29040,N_22387,N_21141);
xnor U29041 (N_29041,N_22178,N_21271);
nor U29042 (N_29042,N_21940,N_24835);
xnor U29043 (N_29043,N_22623,N_23798);
and U29044 (N_29044,N_24798,N_24689);
nand U29045 (N_29045,N_22722,N_22116);
xnor U29046 (N_29046,N_24586,N_24784);
xor U29047 (N_29047,N_20977,N_23850);
and U29048 (N_29048,N_23932,N_24595);
nor U29049 (N_29049,N_24598,N_21223);
xor U29050 (N_29050,N_24253,N_23064);
nand U29051 (N_29051,N_22636,N_22303);
or U29052 (N_29052,N_22043,N_21043);
or U29053 (N_29053,N_20969,N_24616);
and U29054 (N_29054,N_21301,N_23163);
nor U29055 (N_29055,N_21150,N_20012);
nand U29056 (N_29056,N_21611,N_20742);
nor U29057 (N_29057,N_22538,N_23418);
and U29058 (N_29058,N_23544,N_23159);
and U29059 (N_29059,N_21276,N_21943);
and U29060 (N_29060,N_24038,N_21783);
nor U29061 (N_29061,N_20958,N_24960);
and U29062 (N_29062,N_23480,N_21348);
and U29063 (N_29063,N_22542,N_20301);
and U29064 (N_29064,N_20873,N_20415);
xor U29065 (N_29065,N_23055,N_22970);
nand U29066 (N_29066,N_21194,N_20717);
or U29067 (N_29067,N_20755,N_21904);
nand U29068 (N_29068,N_23429,N_20727);
nand U29069 (N_29069,N_24228,N_20808);
xor U29070 (N_29070,N_22179,N_22564);
and U29071 (N_29071,N_22668,N_20169);
nor U29072 (N_29072,N_24724,N_21940);
and U29073 (N_29073,N_22756,N_23469);
or U29074 (N_29074,N_20184,N_21944);
nand U29075 (N_29075,N_22621,N_21886);
or U29076 (N_29076,N_23710,N_24059);
nor U29077 (N_29077,N_20272,N_21477);
xor U29078 (N_29078,N_24008,N_20766);
nand U29079 (N_29079,N_21959,N_21078);
and U29080 (N_29080,N_21864,N_22509);
or U29081 (N_29081,N_23436,N_23176);
and U29082 (N_29082,N_20333,N_20354);
and U29083 (N_29083,N_22445,N_24215);
or U29084 (N_29084,N_24306,N_22792);
nor U29085 (N_29085,N_20235,N_22508);
and U29086 (N_29086,N_21328,N_24622);
nand U29087 (N_29087,N_23304,N_21348);
xnor U29088 (N_29088,N_21352,N_24938);
xor U29089 (N_29089,N_23490,N_23782);
xnor U29090 (N_29090,N_21107,N_21531);
or U29091 (N_29091,N_21099,N_22600);
nand U29092 (N_29092,N_22534,N_20512);
xnor U29093 (N_29093,N_21514,N_23767);
nor U29094 (N_29094,N_23602,N_20314);
or U29095 (N_29095,N_22435,N_22510);
nor U29096 (N_29096,N_22980,N_22235);
nor U29097 (N_29097,N_23952,N_23693);
nor U29098 (N_29098,N_21724,N_21059);
nand U29099 (N_29099,N_23194,N_20339);
xor U29100 (N_29100,N_24138,N_23852);
nand U29101 (N_29101,N_22576,N_23872);
or U29102 (N_29102,N_22094,N_22025);
nand U29103 (N_29103,N_23849,N_22179);
nand U29104 (N_29104,N_20165,N_21286);
xnor U29105 (N_29105,N_22467,N_22737);
nand U29106 (N_29106,N_23475,N_21922);
and U29107 (N_29107,N_22748,N_20106);
xor U29108 (N_29108,N_20042,N_20726);
xnor U29109 (N_29109,N_22188,N_21295);
nand U29110 (N_29110,N_24628,N_23198);
and U29111 (N_29111,N_23099,N_20846);
or U29112 (N_29112,N_23406,N_23253);
or U29113 (N_29113,N_24747,N_23654);
xnor U29114 (N_29114,N_21742,N_22419);
nor U29115 (N_29115,N_22066,N_24402);
or U29116 (N_29116,N_22340,N_21464);
and U29117 (N_29117,N_24507,N_20462);
nor U29118 (N_29118,N_21629,N_24104);
xnor U29119 (N_29119,N_23915,N_22552);
or U29120 (N_29120,N_20187,N_22451);
xor U29121 (N_29121,N_21791,N_24443);
or U29122 (N_29122,N_23067,N_22087);
and U29123 (N_29123,N_20111,N_20814);
or U29124 (N_29124,N_23204,N_23492);
nor U29125 (N_29125,N_20546,N_23305);
nor U29126 (N_29126,N_21848,N_21782);
xnor U29127 (N_29127,N_23571,N_20712);
and U29128 (N_29128,N_20551,N_20421);
and U29129 (N_29129,N_20338,N_22948);
xnor U29130 (N_29130,N_23378,N_24971);
nand U29131 (N_29131,N_24988,N_21483);
nand U29132 (N_29132,N_24118,N_21428);
or U29133 (N_29133,N_22901,N_21457);
or U29134 (N_29134,N_22128,N_20928);
nand U29135 (N_29135,N_20651,N_23667);
and U29136 (N_29136,N_20710,N_24663);
xor U29137 (N_29137,N_22179,N_20854);
and U29138 (N_29138,N_20945,N_24077);
and U29139 (N_29139,N_23834,N_24285);
and U29140 (N_29140,N_24078,N_22437);
nor U29141 (N_29141,N_23123,N_21395);
or U29142 (N_29142,N_20020,N_22151);
nor U29143 (N_29143,N_23774,N_24452);
nand U29144 (N_29144,N_24923,N_20457);
or U29145 (N_29145,N_24022,N_23063);
and U29146 (N_29146,N_22506,N_20459);
nor U29147 (N_29147,N_20080,N_21877);
nand U29148 (N_29148,N_22717,N_22407);
nand U29149 (N_29149,N_24708,N_23301);
xnor U29150 (N_29150,N_20796,N_20998);
nor U29151 (N_29151,N_23089,N_21740);
nor U29152 (N_29152,N_23008,N_24259);
and U29153 (N_29153,N_22478,N_24919);
or U29154 (N_29154,N_21711,N_20065);
or U29155 (N_29155,N_20547,N_20710);
nor U29156 (N_29156,N_22604,N_23323);
nand U29157 (N_29157,N_22763,N_22665);
nor U29158 (N_29158,N_21191,N_24206);
nor U29159 (N_29159,N_21104,N_24414);
nor U29160 (N_29160,N_21192,N_24129);
and U29161 (N_29161,N_24101,N_23492);
xnor U29162 (N_29162,N_23628,N_22767);
or U29163 (N_29163,N_20739,N_22604);
xor U29164 (N_29164,N_23627,N_20245);
nand U29165 (N_29165,N_22014,N_23079);
nand U29166 (N_29166,N_20901,N_24980);
or U29167 (N_29167,N_21221,N_20677);
or U29168 (N_29168,N_22641,N_21967);
or U29169 (N_29169,N_20936,N_24306);
nand U29170 (N_29170,N_22270,N_21151);
xor U29171 (N_29171,N_21521,N_21784);
and U29172 (N_29172,N_23743,N_22539);
or U29173 (N_29173,N_21047,N_22538);
nand U29174 (N_29174,N_22208,N_23349);
or U29175 (N_29175,N_24130,N_24749);
nor U29176 (N_29176,N_22945,N_24891);
nor U29177 (N_29177,N_23310,N_21218);
nand U29178 (N_29178,N_21074,N_21705);
nor U29179 (N_29179,N_23262,N_24653);
xnor U29180 (N_29180,N_21073,N_22966);
or U29181 (N_29181,N_24042,N_24479);
xor U29182 (N_29182,N_21453,N_24274);
or U29183 (N_29183,N_24523,N_20198);
nand U29184 (N_29184,N_24026,N_24886);
and U29185 (N_29185,N_21567,N_20276);
and U29186 (N_29186,N_21193,N_21586);
or U29187 (N_29187,N_20278,N_22349);
xor U29188 (N_29188,N_22059,N_20658);
or U29189 (N_29189,N_24314,N_21124);
or U29190 (N_29190,N_22911,N_24466);
xnor U29191 (N_29191,N_23843,N_22695);
xor U29192 (N_29192,N_23487,N_20155);
xnor U29193 (N_29193,N_22758,N_23323);
nand U29194 (N_29194,N_23505,N_22334);
nand U29195 (N_29195,N_20062,N_22055);
and U29196 (N_29196,N_23673,N_21725);
nand U29197 (N_29197,N_22512,N_23017);
or U29198 (N_29198,N_24084,N_20880);
nand U29199 (N_29199,N_24340,N_24084);
xor U29200 (N_29200,N_21471,N_22539);
nor U29201 (N_29201,N_20986,N_23934);
or U29202 (N_29202,N_21907,N_22838);
nor U29203 (N_29203,N_24723,N_20991);
nand U29204 (N_29204,N_20046,N_21510);
and U29205 (N_29205,N_24293,N_21287);
or U29206 (N_29206,N_21822,N_22294);
and U29207 (N_29207,N_21343,N_23447);
nand U29208 (N_29208,N_22481,N_21778);
or U29209 (N_29209,N_24292,N_24405);
and U29210 (N_29210,N_21532,N_21453);
or U29211 (N_29211,N_21072,N_20087);
nand U29212 (N_29212,N_20398,N_21640);
and U29213 (N_29213,N_21882,N_24172);
or U29214 (N_29214,N_24116,N_21920);
nand U29215 (N_29215,N_24196,N_20434);
and U29216 (N_29216,N_21700,N_22943);
and U29217 (N_29217,N_24630,N_20455);
and U29218 (N_29218,N_22510,N_21209);
nor U29219 (N_29219,N_23223,N_20562);
nand U29220 (N_29220,N_24340,N_22486);
xor U29221 (N_29221,N_24779,N_24239);
and U29222 (N_29222,N_24652,N_21675);
and U29223 (N_29223,N_20271,N_22132);
nand U29224 (N_29224,N_21561,N_22350);
xnor U29225 (N_29225,N_23509,N_24101);
nand U29226 (N_29226,N_24383,N_21768);
or U29227 (N_29227,N_21566,N_20211);
and U29228 (N_29228,N_23352,N_24445);
nand U29229 (N_29229,N_21443,N_24915);
nor U29230 (N_29230,N_24003,N_24069);
or U29231 (N_29231,N_21562,N_23005);
nand U29232 (N_29232,N_24665,N_20482);
or U29233 (N_29233,N_21690,N_22876);
or U29234 (N_29234,N_24725,N_22669);
and U29235 (N_29235,N_22954,N_24012);
nor U29236 (N_29236,N_24479,N_21976);
and U29237 (N_29237,N_23810,N_21469);
and U29238 (N_29238,N_23062,N_21952);
nand U29239 (N_29239,N_20909,N_24378);
nor U29240 (N_29240,N_22506,N_20372);
or U29241 (N_29241,N_21623,N_22403);
nand U29242 (N_29242,N_24096,N_21310);
nor U29243 (N_29243,N_22782,N_24933);
nand U29244 (N_29244,N_20766,N_23755);
xor U29245 (N_29245,N_20209,N_20471);
nor U29246 (N_29246,N_22160,N_24312);
xor U29247 (N_29247,N_22032,N_21193);
nand U29248 (N_29248,N_21880,N_23336);
or U29249 (N_29249,N_24136,N_21253);
nor U29250 (N_29250,N_22361,N_23302);
nand U29251 (N_29251,N_24326,N_22178);
nor U29252 (N_29252,N_20636,N_23301);
nor U29253 (N_29253,N_22388,N_22321);
or U29254 (N_29254,N_20323,N_20888);
and U29255 (N_29255,N_20756,N_21830);
or U29256 (N_29256,N_20209,N_23206);
nand U29257 (N_29257,N_21986,N_24194);
nor U29258 (N_29258,N_20642,N_24405);
xor U29259 (N_29259,N_21706,N_21666);
nor U29260 (N_29260,N_24244,N_22107);
xnor U29261 (N_29261,N_21129,N_21746);
nand U29262 (N_29262,N_22374,N_23114);
or U29263 (N_29263,N_24283,N_24281);
and U29264 (N_29264,N_24753,N_22024);
nor U29265 (N_29265,N_22547,N_20826);
nand U29266 (N_29266,N_20147,N_24624);
and U29267 (N_29267,N_22920,N_23775);
nor U29268 (N_29268,N_22039,N_23183);
xor U29269 (N_29269,N_20460,N_20724);
xor U29270 (N_29270,N_22503,N_23868);
or U29271 (N_29271,N_23074,N_24409);
nor U29272 (N_29272,N_21499,N_24387);
xnor U29273 (N_29273,N_22090,N_21694);
nand U29274 (N_29274,N_24749,N_23150);
or U29275 (N_29275,N_23814,N_20621);
or U29276 (N_29276,N_23989,N_22359);
or U29277 (N_29277,N_24531,N_24785);
nand U29278 (N_29278,N_21856,N_22405);
nor U29279 (N_29279,N_24351,N_20398);
nor U29280 (N_29280,N_21244,N_23331);
and U29281 (N_29281,N_24334,N_22796);
nand U29282 (N_29282,N_22402,N_22391);
or U29283 (N_29283,N_22795,N_22591);
nor U29284 (N_29284,N_21948,N_20714);
nor U29285 (N_29285,N_21996,N_23155);
nand U29286 (N_29286,N_24248,N_22190);
nand U29287 (N_29287,N_23330,N_21401);
xor U29288 (N_29288,N_20843,N_21692);
and U29289 (N_29289,N_21622,N_24074);
nor U29290 (N_29290,N_22653,N_24359);
nor U29291 (N_29291,N_20887,N_22784);
and U29292 (N_29292,N_20374,N_20269);
nand U29293 (N_29293,N_21797,N_23575);
nor U29294 (N_29294,N_20728,N_20922);
nand U29295 (N_29295,N_22428,N_22769);
nand U29296 (N_29296,N_20921,N_24595);
nor U29297 (N_29297,N_24977,N_20758);
xnor U29298 (N_29298,N_23174,N_22433);
nor U29299 (N_29299,N_21463,N_21457);
or U29300 (N_29300,N_20656,N_21955);
or U29301 (N_29301,N_23606,N_21322);
and U29302 (N_29302,N_20148,N_23474);
nand U29303 (N_29303,N_21089,N_24668);
xnor U29304 (N_29304,N_24356,N_23163);
nand U29305 (N_29305,N_23400,N_24261);
nor U29306 (N_29306,N_20948,N_23272);
or U29307 (N_29307,N_20596,N_24542);
xor U29308 (N_29308,N_20240,N_24166);
and U29309 (N_29309,N_22376,N_20659);
and U29310 (N_29310,N_21104,N_22118);
nand U29311 (N_29311,N_24211,N_21770);
nor U29312 (N_29312,N_22569,N_21333);
and U29313 (N_29313,N_20764,N_24622);
or U29314 (N_29314,N_20986,N_24165);
or U29315 (N_29315,N_23408,N_22669);
nor U29316 (N_29316,N_20999,N_24414);
and U29317 (N_29317,N_23616,N_23138);
nor U29318 (N_29318,N_24214,N_24195);
and U29319 (N_29319,N_22522,N_23893);
nand U29320 (N_29320,N_20939,N_23386);
nand U29321 (N_29321,N_24930,N_20530);
and U29322 (N_29322,N_22439,N_21398);
xor U29323 (N_29323,N_22119,N_21903);
and U29324 (N_29324,N_24342,N_22007);
or U29325 (N_29325,N_22712,N_20951);
nor U29326 (N_29326,N_20983,N_22632);
nor U29327 (N_29327,N_24873,N_24172);
nor U29328 (N_29328,N_22982,N_20077);
nor U29329 (N_29329,N_24202,N_22143);
nand U29330 (N_29330,N_21068,N_24940);
and U29331 (N_29331,N_20484,N_23920);
nor U29332 (N_29332,N_20548,N_22100);
and U29333 (N_29333,N_23584,N_21104);
xnor U29334 (N_29334,N_20999,N_20746);
or U29335 (N_29335,N_24402,N_20789);
nand U29336 (N_29336,N_24561,N_23474);
nand U29337 (N_29337,N_24795,N_24711);
nand U29338 (N_29338,N_24918,N_24285);
nand U29339 (N_29339,N_24061,N_22914);
xor U29340 (N_29340,N_22159,N_23330);
nor U29341 (N_29341,N_23929,N_20047);
xor U29342 (N_29342,N_23626,N_23939);
or U29343 (N_29343,N_24886,N_22783);
nand U29344 (N_29344,N_24084,N_21077);
nor U29345 (N_29345,N_21777,N_23469);
nor U29346 (N_29346,N_24207,N_21658);
xnor U29347 (N_29347,N_23987,N_23227);
and U29348 (N_29348,N_21272,N_22415);
xor U29349 (N_29349,N_22004,N_21863);
and U29350 (N_29350,N_22246,N_21092);
and U29351 (N_29351,N_22148,N_22864);
xor U29352 (N_29352,N_20100,N_22100);
or U29353 (N_29353,N_22050,N_24214);
and U29354 (N_29354,N_21391,N_23956);
xor U29355 (N_29355,N_20593,N_23893);
and U29356 (N_29356,N_21223,N_20972);
nand U29357 (N_29357,N_20678,N_23930);
or U29358 (N_29358,N_20589,N_24875);
nor U29359 (N_29359,N_24941,N_21550);
xor U29360 (N_29360,N_20234,N_20605);
nor U29361 (N_29361,N_22968,N_23447);
nand U29362 (N_29362,N_23748,N_20536);
or U29363 (N_29363,N_24241,N_24480);
or U29364 (N_29364,N_22468,N_24829);
or U29365 (N_29365,N_20747,N_21775);
and U29366 (N_29366,N_20044,N_21200);
nand U29367 (N_29367,N_24717,N_21736);
or U29368 (N_29368,N_24081,N_20305);
xor U29369 (N_29369,N_20021,N_24748);
nand U29370 (N_29370,N_21629,N_21901);
nand U29371 (N_29371,N_24100,N_20194);
or U29372 (N_29372,N_23743,N_21110);
or U29373 (N_29373,N_21682,N_23836);
and U29374 (N_29374,N_22984,N_21125);
xor U29375 (N_29375,N_22214,N_23128);
nor U29376 (N_29376,N_24077,N_24971);
or U29377 (N_29377,N_24672,N_21660);
nand U29378 (N_29378,N_22272,N_21893);
nor U29379 (N_29379,N_24437,N_24476);
or U29380 (N_29380,N_20575,N_22118);
and U29381 (N_29381,N_23743,N_23009);
nand U29382 (N_29382,N_23615,N_24580);
and U29383 (N_29383,N_22473,N_20137);
xnor U29384 (N_29384,N_23278,N_20060);
xor U29385 (N_29385,N_24533,N_22543);
or U29386 (N_29386,N_20638,N_23593);
xnor U29387 (N_29387,N_21082,N_24732);
nor U29388 (N_29388,N_22479,N_20459);
xnor U29389 (N_29389,N_20339,N_21632);
nand U29390 (N_29390,N_20556,N_22546);
xor U29391 (N_29391,N_24649,N_21226);
or U29392 (N_29392,N_24031,N_22115);
xnor U29393 (N_29393,N_22688,N_24974);
xnor U29394 (N_29394,N_21966,N_22487);
or U29395 (N_29395,N_23226,N_22437);
nand U29396 (N_29396,N_20548,N_23583);
nand U29397 (N_29397,N_21453,N_20691);
or U29398 (N_29398,N_22498,N_23201);
nand U29399 (N_29399,N_24483,N_22953);
nand U29400 (N_29400,N_21601,N_23884);
and U29401 (N_29401,N_21403,N_20628);
xnor U29402 (N_29402,N_24180,N_22545);
nand U29403 (N_29403,N_20198,N_24948);
xnor U29404 (N_29404,N_22492,N_21910);
and U29405 (N_29405,N_22089,N_22099);
nor U29406 (N_29406,N_20100,N_22763);
nor U29407 (N_29407,N_22751,N_22636);
or U29408 (N_29408,N_21785,N_21432);
nand U29409 (N_29409,N_23785,N_20872);
and U29410 (N_29410,N_22194,N_24954);
nand U29411 (N_29411,N_23863,N_23470);
and U29412 (N_29412,N_23790,N_21760);
and U29413 (N_29413,N_22566,N_20818);
or U29414 (N_29414,N_22694,N_20949);
nor U29415 (N_29415,N_20322,N_23798);
and U29416 (N_29416,N_23474,N_20678);
or U29417 (N_29417,N_24457,N_23390);
and U29418 (N_29418,N_21139,N_23860);
nand U29419 (N_29419,N_20790,N_21981);
nor U29420 (N_29420,N_20574,N_23011);
nand U29421 (N_29421,N_24672,N_20263);
nand U29422 (N_29422,N_22217,N_21337);
and U29423 (N_29423,N_24391,N_23998);
nand U29424 (N_29424,N_24619,N_23086);
nand U29425 (N_29425,N_21975,N_23412);
nor U29426 (N_29426,N_21688,N_23906);
nor U29427 (N_29427,N_20388,N_20615);
xor U29428 (N_29428,N_22755,N_24456);
nor U29429 (N_29429,N_20068,N_23625);
nand U29430 (N_29430,N_20994,N_21879);
or U29431 (N_29431,N_22296,N_21562);
xor U29432 (N_29432,N_22082,N_24225);
and U29433 (N_29433,N_24274,N_21949);
nand U29434 (N_29434,N_22122,N_24480);
xor U29435 (N_29435,N_21842,N_21978);
nor U29436 (N_29436,N_20122,N_23258);
xnor U29437 (N_29437,N_21440,N_21328);
and U29438 (N_29438,N_24165,N_23868);
nor U29439 (N_29439,N_21161,N_24052);
nor U29440 (N_29440,N_21949,N_21334);
nand U29441 (N_29441,N_20055,N_22778);
or U29442 (N_29442,N_20723,N_20421);
or U29443 (N_29443,N_21244,N_24393);
nand U29444 (N_29444,N_24279,N_20778);
xnor U29445 (N_29445,N_22542,N_20358);
and U29446 (N_29446,N_24931,N_20793);
xor U29447 (N_29447,N_20868,N_23628);
and U29448 (N_29448,N_21035,N_23549);
nand U29449 (N_29449,N_23385,N_21169);
nand U29450 (N_29450,N_23440,N_22222);
or U29451 (N_29451,N_22395,N_20792);
xnor U29452 (N_29452,N_21365,N_24337);
nor U29453 (N_29453,N_23106,N_21298);
nand U29454 (N_29454,N_22903,N_20153);
and U29455 (N_29455,N_20168,N_21957);
nand U29456 (N_29456,N_21129,N_23259);
nor U29457 (N_29457,N_23901,N_23841);
or U29458 (N_29458,N_20706,N_20007);
or U29459 (N_29459,N_20529,N_20771);
nand U29460 (N_29460,N_21448,N_21973);
and U29461 (N_29461,N_22105,N_20631);
nand U29462 (N_29462,N_24812,N_21367);
nor U29463 (N_29463,N_23561,N_24427);
nand U29464 (N_29464,N_20512,N_22914);
or U29465 (N_29465,N_24683,N_20189);
xnor U29466 (N_29466,N_21414,N_20162);
and U29467 (N_29467,N_20351,N_22265);
nor U29468 (N_29468,N_22604,N_24947);
nor U29469 (N_29469,N_23292,N_21736);
or U29470 (N_29470,N_20241,N_20859);
and U29471 (N_29471,N_22444,N_21854);
and U29472 (N_29472,N_23630,N_22688);
or U29473 (N_29473,N_20372,N_22705);
nand U29474 (N_29474,N_20507,N_20311);
nand U29475 (N_29475,N_23686,N_21119);
and U29476 (N_29476,N_23295,N_20962);
nand U29477 (N_29477,N_24335,N_21904);
nor U29478 (N_29478,N_23228,N_20918);
nor U29479 (N_29479,N_21709,N_22089);
nand U29480 (N_29480,N_21029,N_21411);
nand U29481 (N_29481,N_20901,N_20250);
and U29482 (N_29482,N_24398,N_20845);
or U29483 (N_29483,N_24983,N_20577);
xor U29484 (N_29484,N_23842,N_20617);
xnor U29485 (N_29485,N_23821,N_24583);
xnor U29486 (N_29486,N_22297,N_21136);
xnor U29487 (N_29487,N_23485,N_21777);
nand U29488 (N_29488,N_21063,N_21568);
nand U29489 (N_29489,N_20028,N_20400);
nand U29490 (N_29490,N_20392,N_21719);
or U29491 (N_29491,N_23909,N_22496);
nand U29492 (N_29492,N_21297,N_20308);
and U29493 (N_29493,N_24975,N_24446);
nand U29494 (N_29494,N_21341,N_23056);
or U29495 (N_29495,N_23087,N_24567);
nor U29496 (N_29496,N_21473,N_21644);
or U29497 (N_29497,N_21510,N_24903);
or U29498 (N_29498,N_21078,N_22026);
xor U29499 (N_29499,N_23604,N_23591);
or U29500 (N_29500,N_24859,N_20748);
nand U29501 (N_29501,N_21006,N_22200);
or U29502 (N_29502,N_22447,N_23305);
nand U29503 (N_29503,N_22567,N_22740);
and U29504 (N_29504,N_21302,N_20337);
nand U29505 (N_29505,N_21582,N_20388);
xnor U29506 (N_29506,N_21202,N_23790);
and U29507 (N_29507,N_24088,N_22907);
or U29508 (N_29508,N_23262,N_21484);
nor U29509 (N_29509,N_21708,N_20425);
nor U29510 (N_29510,N_23708,N_22008);
nor U29511 (N_29511,N_23505,N_24688);
xor U29512 (N_29512,N_24206,N_20945);
or U29513 (N_29513,N_21261,N_22179);
or U29514 (N_29514,N_21835,N_24632);
nand U29515 (N_29515,N_23974,N_23407);
and U29516 (N_29516,N_24290,N_24278);
nor U29517 (N_29517,N_23014,N_22802);
xnor U29518 (N_29518,N_22734,N_24233);
nor U29519 (N_29519,N_22241,N_20001);
or U29520 (N_29520,N_24216,N_22620);
nand U29521 (N_29521,N_21854,N_20058);
nor U29522 (N_29522,N_24462,N_23704);
nand U29523 (N_29523,N_22117,N_23956);
or U29524 (N_29524,N_23973,N_23512);
xor U29525 (N_29525,N_24180,N_21527);
and U29526 (N_29526,N_24061,N_21563);
or U29527 (N_29527,N_20293,N_21313);
and U29528 (N_29528,N_22238,N_23362);
xor U29529 (N_29529,N_24471,N_23122);
nand U29530 (N_29530,N_21808,N_23688);
or U29531 (N_29531,N_22360,N_21258);
xnor U29532 (N_29532,N_21373,N_21085);
nor U29533 (N_29533,N_21081,N_23959);
or U29534 (N_29534,N_23392,N_20686);
xnor U29535 (N_29535,N_23712,N_20940);
and U29536 (N_29536,N_21810,N_22849);
nand U29537 (N_29537,N_24240,N_21303);
xnor U29538 (N_29538,N_22626,N_20272);
and U29539 (N_29539,N_23469,N_23685);
nand U29540 (N_29540,N_21112,N_20218);
and U29541 (N_29541,N_23232,N_22672);
or U29542 (N_29542,N_22335,N_20915);
or U29543 (N_29543,N_21723,N_21581);
nand U29544 (N_29544,N_21891,N_22671);
or U29545 (N_29545,N_20290,N_24635);
nor U29546 (N_29546,N_21522,N_23833);
nor U29547 (N_29547,N_20676,N_24491);
nor U29548 (N_29548,N_22351,N_20563);
or U29549 (N_29549,N_23978,N_22288);
nor U29550 (N_29550,N_24410,N_23798);
xor U29551 (N_29551,N_20678,N_20526);
and U29552 (N_29552,N_20043,N_20897);
nor U29553 (N_29553,N_22355,N_20649);
nand U29554 (N_29554,N_23774,N_24418);
nor U29555 (N_29555,N_20470,N_20239);
nor U29556 (N_29556,N_20375,N_23130);
xnor U29557 (N_29557,N_24433,N_22749);
nor U29558 (N_29558,N_23374,N_20930);
and U29559 (N_29559,N_20019,N_22104);
nor U29560 (N_29560,N_24569,N_21185);
xnor U29561 (N_29561,N_20411,N_23898);
nor U29562 (N_29562,N_24555,N_21040);
and U29563 (N_29563,N_24637,N_21858);
or U29564 (N_29564,N_21513,N_21200);
or U29565 (N_29565,N_22063,N_22077);
nand U29566 (N_29566,N_23492,N_23627);
or U29567 (N_29567,N_22173,N_21432);
and U29568 (N_29568,N_24153,N_23425);
or U29569 (N_29569,N_24874,N_23825);
xor U29570 (N_29570,N_21949,N_23439);
or U29571 (N_29571,N_22493,N_20827);
or U29572 (N_29572,N_23381,N_22966);
and U29573 (N_29573,N_20982,N_21146);
nor U29574 (N_29574,N_20029,N_20190);
nor U29575 (N_29575,N_23856,N_21790);
nand U29576 (N_29576,N_24254,N_22330);
nor U29577 (N_29577,N_23968,N_22609);
and U29578 (N_29578,N_22329,N_24804);
or U29579 (N_29579,N_22299,N_24291);
and U29580 (N_29580,N_21008,N_24276);
nor U29581 (N_29581,N_20103,N_22596);
or U29582 (N_29582,N_24483,N_24469);
nand U29583 (N_29583,N_20090,N_21050);
nand U29584 (N_29584,N_23689,N_24589);
nand U29585 (N_29585,N_24648,N_20079);
nor U29586 (N_29586,N_21747,N_21767);
xnor U29587 (N_29587,N_24484,N_23572);
nor U29588 (N_29588,N_20249,N_21482);
nand U29589 (N_29589,N_22433,N_24206);
nand U29590 (N_29590,N_21453,N_20926);
nor U29591 (N_29591,N_23240,N_21480);
and U29592 (N_29592,N_21166,N_20073);
nor U29593 (N_29593,N_23882,N_21915);
nand U29594 (N_29594,N_21655,N_23985);
or U29595 (N_29595,N_23528,N_24516);
or U29596 (N_29596,N_24632,N_20078);
and U29597 (N_29597,N_24821,N_23105);
nor U29598 (N_29598,N_24760,N_22134);
nand U29599 (N_29599,N_22891,N_21222);
and U29600 (N_29600,N_21633,N_24815);
xnor U29601 (N_29601,N_20372,N_24176);
xnor U29602 (N_29602,N_23419,N_21931);
nand U29603 (N_29603,N_20274,N_22843);
or U29604 (N_29604,N_23713,N_21728);
nand U29605 (N_29605,N_23328,N_20142);
xnor U29606 (N_29606,N_24538,N_22983);
nand U29607 (N_29607,N_24284,N_24405);
xnor U29608 (N_29608,N_22347,N_21154);
nor U29609 (N_29609,N_23827,N_22991);
xor U29610 (N_29610,N_22443,N_21272);
nor U29611 (N_29611,N_22256,N_20524);
and U29612 (N_29612,N_20421,N_23556);
nor U29613 (N_29613,N_21658,N_24114);
nor U29614 (N_29614,N_20264,N_22791);
or U29615 (N_29615,N_20685,N_23197);
xnor U29616 (N_29616,N_20820,N_20241);
xnor U29617 (N_29617,N_20656,N_24134);
or U29618 (N_29618,N_24248,N_22913);
nand U29619 (N_29619,N_21795,N_20193);
or U29620 (N_29620,N_20193,N_20998);
or U29621 (N_29621,N_22098,N_22414);
or U29622 (N_29622,N_24936,N_20461);
and U29623 (N_29623,N_24366,N_23767);
xor U29624 (N_29624,N_24418,N_24265);
nor U29625 (N_29625,N_23596,N_24621);
xnor U29626 (N_29626,N_24318,N_20976);
nand U29627 (N_29627,N_20888,N_23667);
or U29628 (N_29628,N_23539,N_21226);
and U29629 (N_29629,N_21243,N_23663);
xor U29630 (N_29630,N_20874,N_21166);
nor U29631 (N_29631,N_20679,N_20774);
nand U29632 (N_29632,N_23037,N_22223);
or U29633 (N_29633,N_24422,N_20075);
and U29634 (N_29634,N_23073,N_21378);
xnor U29635 (N_29635,N_24012,N_23685);
xnor U29636 (N_29636,N_22480,N_23023);
nand U29637 (N_29637,N_24659,N_21559);
nor U29638 (N_29638,N_23933,N_24391);
nor U29639 (N_29639,N_22578,N_23901);
or U29640 (N_29640,N_22851,N_24077);
xnor U29641 (N_29641,N_21654,N_24882);
or U29642 (N_29642,N_20083,N_23376);
xnor U29643 (N_29643,N_22103,N_23392);
xnor U29644 (N_29644,N_20538,N_22981);
or U29645 (N_29645,N_24257,N_21117);
xnor U29646 (N_29646,N_20452,N_20541);
and U29647 (N_29647,N_24920,N_23677);
nand U29648 (N_29648,N_20858,N_24534);
and U29649 (N_29649,N_20133,N_23542);
nand U29650 (N_29650,N_21105,N_22987);
xor U29651 (N_29651,N_24110,N_20160);
or U29652 (N_29652,N_23957,N_20742);
nor U29653 (N_29653,N_22777,N_23812);
or U29654 (N_29654,N_21488,N_20377);
xor U29655 (N_29655,N_22088,N_24134);
xor U29656 (N_29656,N_23239,N_20403);
xor U29657 (N_29657,N_21224,N_21002);
nor U29658 (N_29658,N_20828,N_21871);
nor U29659 (N_29659,N_21281,N_20330);
or U29660 (N_29660,N_20966,N_22435);
or U29661 (N_29661,N_22429,N_24209);
and U29662 (N_29662,N_20161,N_23655);
nor U29663 (N_29663,N_23121,N_24394);
and U29664 (N_29664,N_22767,N_23346);
or U29665 (N_29665,N_22883,N_23541);
or U29666 (N_29666,N_24059,N_20283);
xnor U29667 (N_29667,N_22472,N_21864);
and U29668 (N_29668,N_24085,N_21868);
nor U29669 (N_29669,N_24427,N_23413);
nor U29670 (N_29670,N_23747,N_23110);
nor U29671 (N_29671,N_20446,N_21763);
or U29672 (N_29672,N_24538,N_23324);
xnor U29673 (N_29673,N_20701,N_22835);
or U29674 (N_29674,N_24034,N_23546);
xnor U29675 (N_29675,N_24385,N_20853);
or U29676 (N_29676,N_23280,N_22728);
nand U29677 (N_29677,N_20158,N_23788);
nand U29678 (N_29678,N_20050,N_21085);
xor U29679 (N_29679,N_23904,N_23192);
nor U29680 (N_29680,N_20861,N_24866);
xnor U29681 (N_29681,N_23578,N_20692);
nor U29682 (N_29682,N_21238,N_22683);
nor U29683 (N_29683,N_24823,N_24935);
and U29684 (N_29684,N_24737,N_21977);
nor U29685 (N_29685,N_22637,N_21904);
nand U29686 (N_29686,N_22565,N_23015);
nand U29687 (N_29687,N_24137,N_23484);
xor U29688 (N_29688,N_22189,N_23245);
nor U29689 (N_29689,N_20698,N_21109);
xnor U29690 (N_29690,N_23597,N_22630);
nand U29691 (N_29691,N_20366,N_22261);
or U29692 (N_29692,N_24339,N_23547);
or U29693 (N_29693,N_22578,N_20445);
nand U29694 (N_29694,N_23349,N_22167);
xnor U29695 (N_29695,N_24302,N_23206);
nand U29696 (N_29696,N_22929,N_22395);
nor U29697 (N_29697,N_24156,N_22908);
nor U29698 (N_29698,N_24226,N_20019);
or U29699 (N_29699,N_21664,N_20877);
or U29700 (N_29700,N_23165,N_23204);
and U29701 (N_29701,N_20877,N_20823);
or U29702 (N_29702,N_23118,N_21908);
nand U29703 (N_29703,N_23566,N_22560);
xor U29704 (N_29704,N_21218,N_21857);
xor U29705 (N_29705,N_20150,N_22289);
nand U29706 (N_29706,N_22695,N_20896);
or U29707 (N_29707,N_23716,N_21510);
or U29708 (N_29708,N_24235,N_20165);
and U29709 (N_29709,N_24226,N_23960);
nor U29710 (N_29710,N_22725,N_24075);
xor U29711 (N_29711,N_20441,N_21748);
nand U29712 (N_29712,N_22933,N_21538);
nor U29713 (N_29713,N_23444,N_23786);
xnor U29714 (N_29714,N_22092,N_20439);
xor U29715 (N_29715,N_21646,N_20610);
nand U29716 (N_29716,N_23536,N_23334);
nor U29717 (N_29717,N_22035,N_24622);
or U29718 (N_29718,N_20409,N_20431);
nor U29719 (N_29719,N_20226,N_24889);
nand U29720 (N_29720,N_20021,N_23330);
nand U29721 (N_29721,N_23907,N_24340);
nor U29722 (N_29722,N_21720,N_22156);
or U29723 (N_29723,N_23297,N_24046);
and U29724 (N_29724,N_21193,N_21067);
or U29725 (N_29725,N_20987,N_21686);
nor U29726 (N_29726,N_21944,N_20290);
or U29727 (N_29727,N_20393,N_22977);
nor U29728 (N_29728,N_22775,N_23070);
nor U29729 (N_29729,N_21933,N_20532);
or U29730 (N_29730,N_20010,N_22386);
and U29731 (N_29731,N_20497,N_23573);
xor U29732 (N_29732,N_21772,N_22669);
nor U29733 (N_29733,N_22973,N_22436);
or U29734 (N_29734,N_20834,N_23551);
nor U29735 (N_29735,N_21816,N_20533);
nand U29736 (N_29736,N_24879,N_23178);
xor U29737 (N_29737,N_23590,N_24322);
or U29738 (N_29738,N_21923,N_20222);
xnor U29739 (N_29739,N_24016,N_23172);
nor U29740 (N_29740,N_24979,N_20844);
or U29741 (N_29741,N_23799,N_23658);
xor U29742 (N_29742,N_21510,N_20470);
nor U29743 (N_29743,N_21327,N_21810);
nand U29744 (N_29744,N_21742,N_22094);
and U29745 (N_29745,N_22381,N_22484);
nand U29746 (N_29746,N_24225,N_23217);
and U29747 (N_29747,N_21933,N_24549);
and U29748 (N_29748,N_20277,N_20792);
or U29749 (N_29749,N_23409,N_24561);
and U29750 (N_29750,N_21795,N_22632);
nor U29751 (N_29751,N_21680,N_20686);
xor U29752 (N_29752,N_22151,N_23410);
xnor U29753 (N_29753,N_23983,N_22321);
nor U29754 (N_29754,N_21698,N_24304);
nand U29755 (N_29755,N_20707,N_24225);
nor U29756 (N_29756,N_22348,N_24845);
xor U29757 (N_29757,N_20339,N_23107);
and U29758 (N_29758,N_21793,N_23777);
or U29759 (N_29759,N_23173,N_20001);
or U29760 (N_29760,N_22541,N_21120);
xnor U29761 (N_29761,N_22465,N_24769);
nor U29762 (N_29762,N_24992,N_21709);
nor U29763 (N_29763,N_24116,N_21902);
xor U29764 (N_29764,N_22809,N_23392);
and U29765 (N_29765,N_24793,N_21606);
nor U29766 (N_29766,N_20659,N_23130);
nand U29767 (N_29767,N_21892,N_24890);
nor U29768 (N_29768,N_21503,N_22903);
xnor U29769 (N_29769,N_24901,N_21958);
nand U29770 (N_29770,N_22307,N_21091);
xnor U29771 (N_29771,N_23090,N_24915);
nor U29772 (N_29772,N_21477,N_21363);
nor U29773 (N_29773,N_24762,N_20605);
and U29774 (N_29774,N_21062,N_21124);
nor U29775 (N_29775,N_23292,N_22164);
or U29776 (N_29776,N_21371,N_21746);
or U29777 (N_29777,N_22054,N_20907);
xnor U29778 (N_29778,N_22907,N_20497);
or U29779 (N_29779,N_21764,N_22859);
nor U29780 (N_29780,N_21077,N_23758);
and U29781 (N_29781,N_22406,N_20556);
nor U29782 (N_29782,N_22767,N_20880);
or U29783 (N_29783,N_20155,N_22029);
and U29784 (N_29784,N_20110,N_23204);
xnor U29785 (N_29785,N_22310,N_24534);
nand U29786 (N_29786,N_21842,N_24111);
xnor U29787 (N_29787,N_24640,N_23443);
xnor U29788 (N_29788,N_22508,N_23480);
and U29789 (N_29789,N_21749,N_21944);
nand U29790 (N_29790,N_23143,N_20392);
nor U29791 (N_29791,N_23912,N_21109);
or U29792 (N_29792,N_20108,N_23636);
and U29793 (N_29793,N_20444,N_22493);
nand U29794 (N_29794,N_24852,N_21999);
or U29795 (N_29795,N_21553,N_20746);
nor U29796 (N_29796,N_23172,N_23542);
nand U29797 (N_29797,N_21428,N_24775);
or U29798 (N_29798,N_23815,N_20773);
nor U29799 (N_29799,N_23061,N_20947);
nor U29800 (N_29800,N_23517,N_20623);
and U29801 (N_29801,N_21754,N_21110);
nand U29802 (N_29802,N_20238,N_23195);
and U29803 (N_29803,N_21606,N_21035);
xor U29804 (N_29804,N_20327,N_20855);
nor U29805 (N_29805,N_21838,N_22534);
nor U29806 (N_29806,N_20212,N_23046);
or U29807 (N_29807,N_23652,N_24747);
nand U29808 (N_29808,N_24999,N_24796);
nor U29809 (N_29809,N_22570,N_20445);
xnor U29810 (N_29810,N_20260,N_22206);
xor U29811 (N_29811,N_23554,N_20194);
nand U29812 (N_29812,N_22197,N_22697);
and U29813 (N_29813,N_23208,N_23961);
and U29814 (N_29814,N_24746,N_20447);
or U29815 (N_29815,N_24804,N_20946);
and U29816 (N_29816,N_22020,N_20943);
xnor U29817 (N_29817,N_24971,N_21410);
and U29818 (N_29818,N_21563,N_24474);
nand U29819 (N_29819,N_21891,N_23634);
xor U29820 (N_29820,N_23205,N_24028);
and U29821 (N_29821,N_23577,N_23148);
xor U29822 (N_29822,N_21121,N_21407);
nor U29823 (N_29823,N_24478,N_23718);
nor U29824 (N_29824,N_23069,N_21601);
nand U29825 (N_29825,N_22388,N_21369);
nand U29826 (N_29826,N_23993,N_20590);
nand U29827 (N_29827,N_21349,N_22538);
nand U29828 (N_29828,N_22594,N_24717);
and U29829 (N_29829,N_21804,N_24346);
nor U29830 (N_29830,N_21087,N_24462);
xnor U29831 (N_29831,N_21853,N_21979);
and U29832 (N_29832,N_22847,N_20776);
or U29833 (N_29833,N_23259,N_23701);
nor U29834 (N_29834,N_22541,N_24583);
xor U29835 (N_29835,N_22568,N_20367);
or U29836 (N_29836,N_23290,N_22846);
nor U29837 (N_29837,N_23196,N_21341);
nand U29838 (N_29838,N_24761,N_20591);
and U29839 (N_29839,N_24411,N_23995);
or U29840 (N_29840,N_20072,N_22412);
nand U29841 (N_29841,N_22751,N_23154);
nor U29842 (N_29842,N_24005,N_24263);
nand U29843 (N_29843,N_23855,N_20602);
or U29844 (N_29844,N_21523,N_22979);
nand U29845 (N_29845,N_22710,N_23357);
or U29846 (N_29846,N_20474,N_22973);
nor U29847 (N_29847,N_23326,N_22298);
nor U29848 (N_29848,N_24588,N_23419);
nor U29849 (N_29849,N_23578,N_20680);
nor U29850 (N_29850,N_21039,N_24591);
xnor U29851 (N_29851,N_20691,N_24787);
or U29852 (N_29852,N_24326,N_23668);
nor U29853 (N_29853,N_21769,N_21752);
nand U29854 (N_29854,N_24106,N_20425);
or U29855 (N_29855,N_23167,N_22151);
or U29856 (N_29856,N_22475,N_22589);
or U29857 (N_29857,N_21506,N_23734);
or U29858 (N_29858,N_24778,N_22950);
or U29859 (N_29859,N_20529,N_24873);
or U29860 (N_29860,N_20157,N_21872);
nand U29861 (N_29861,N_24399,N_20041);
xnor U29862 (N_29862,N_22272,N_22688);
xor U29863 (N_29863,N_22144,N_24418);
nand U29864 (N_29864,N_21816,N_21805);
nor U29865 (N_29865,N_24588,N_22218);
and U29866 (N_29866,N_20215,N_24792);
xnor U29867 (N_29867,N_22895,N_21583);
or U29868 (N_29868,N_22427,N_23346);
xor U29869 (N_29869,N_24460,N_21705);
and U29870 (N_29870,N_22281,N_23902);
nand U29871 (N_29871,N_22801,N_23886);
and U29872 (N_29872,N_22988,N_23992);
and U29873 (N_29873,N_22041,N_24492);
and U29874 (N_29874,N_24314,N_22655);
xor U29875 (N_29875,N_21588,N_23840);
xor U29876 (N_29876,N_24569,N_23200);
or U29877 (N_29877,N_20943,N_23234);
nor U29878 (N_29878,N_24728,N_23846);
or U29879 (N_29879,N_24477,N_22464);
or U29880 (N_29880,N_20871,N_22058);
xnor U29881 (N_29881,N_20544,N_21380);
nand U29882 (N_29882,N_20092,N_24329);
nand U29883 (N_29883,N_24840,N_20926);
and U29884 (N_29884,N_22508,N_20748);
and U29885 (N_29885,N_20432,N_22986);
nand U29886 (N_29886,N_20034,N_23386);
xnor U29887 (N_29887,N_23582,N_21449);
or U29888 (N_29888,N_22802,N_24673);
nand U29889 (N_29889,N_23079,N_24441);
nor U29890 (N_29890,N_23048,N_23609);
nand U29891 (N_29891,N_24695,N_22087);
or U29892 (N_29892,N_21638,N_22408);
nand U29893 (N_29893,N_20268,N_23420);
nor U29894 (N_29894,N_23244,N_23021);
xor U29895 (N_29895,N_23994,N_21637);
and U29896 (N_29896,N_20414,N_21762);
or U29897 (N_29897,N_23152,N_23514);
nand U29898 (N_29898,N_22124,N_24693);
xnor U29899 (N_29899,N_23114,N_20738);
nor U29900 (N_29900,N_24537,N_21605);
nand U29901 (N_29901,N_23471,N_21542);
and U29902 (N_29902,N_22543,N_24871);
and U29903 (N_29903,N_22716,N_24923);
nor U29904 (N_29904,N_24815,N_24254);
nand U29905 (N_29905,N_21322,N_24473);
nor U29906 (N_29906,N_23921,N_23321);
and U29907 (N_29907,N_23972,N_24885);
or U29908 (N_29908,N_23254,N_21039);
nand U29909 (N_29909,N_20350,N_20085);
or U29910 (N_29910,N_20027,N_24488);
nand U29911 (N_29911,N_24085,N_22588);
nand U29912 (N_29912,N_21272,N_20561);
and U29913 (N_29913,N_20659,N_20929);
or U29914 (N_29914,N_22590,N_22658);
nand U29915 (N_29915,N_24260,N_20767);
nand U29916 (N_29916,N_20392,N_21490);
and U29917 (N_29917,N_21336,N_21706);
nand U29918 (N_29918,N_22961,N_22447);
and U29919 (N_29919,N_22141,N_24947);
nor U29920 (N_29920,N_24986,N_23027);
nor U29921 (N_29921,N_20386,N_20109);
nand U29922 (N_29922,N_23471,N_22060);
nand U29923 (N_29923,N_22758,N_24084);
xnor U29924 (N_29924,N_20937,N_23229);
nor U29925 (N_29925,N_24355,N_24290);
and U29926 (N_29926,N_20034,N_21566);
xnor U29927 (N_29927,N_24206,N_20283);
xnor U29928 (N_29928,N_20433,N_22070);
xor U29929 (N_29929,N_23037,N_23668);
or U29930 (N_29930,N_22928,N_23042);
nand U29931 (N_29931,N_22658,N_24323);
or U29932 (N_29932,N_24274,N_21025);
and U29933 (N_29933,N_22393,N_23814);
nor U29934 (N_29934,N_22963,N_24495);
nand U29935 (N_29935,N_23955,N_24163);
and U29936 (N_29936,N_24694,N_22323);
and U29937 (N_29937,N_20220,N_22652);
and U29938 (N_29938,N_24749,N_20935);
nor U29939 (N_29939,N_23041,N_24728);
xnor U29940 (N_29940,N_24729,N_23487);
or U29941 (N_29941,N_22878,N_23480);
or U29942 (N_29942,N_20198,N_22527);
or U29943 (N_29943,N_22959,N_22152);
and U29944 (N_29944,N_22062,N_20063);
nand U29945 (N_29945,N_24036,N_22001);
nor U29946 (N_29946,N_20327,N_20969);
nand U29947 (N_29947,N_20140,N_22901);
or U29948 (N_29948,N_21393,N_24351);
nor U29949 (N_29949,N_24096,N_20337);
or U29950 (N_29950,N_24823,N_24124);
nor U29951 (N_29951,N_20211,N_23774);
xnor U29952 (N_29952,N_20598,N_24011);
or U29953 (N_29953,N_22127,N_22178);
or U29954 (N_29954,N_22165,N_20695);
and U29955 (N_29955,N_22840,N_21340);
nor U29956 (N_29956,N_21443,N_21321);
nand U29957 (N_29957,N_24600,N_22223);
and U29958 (N_29958,N_22836,N_23700);
and U29959 (N_29959,N_21699,N_23720);
nor U29960 (N_29960,N_23503,N_21937);
nor U29961 (N_29961,N_24670,N_21274);
xor U29962 (N_29962,N_21369,N_23728);
nor U29963 (N_29963,N_21330,N_20476);
and U29964 (N_29964,N_23781,N_23329);
nor U29965 (N_29965,N_23644,N_24053);
nor U29966 (N_29966,N_21161,N_21552);
nand U29967 (N_29967,N_21255,N_22731);
xor U29968 (N_29968,N_20189,N_20452);
nor U29969 (N_29969,N_21037,N_23791);
xnor U29970 (N_29970,N_21332,N_22340);
or U29971 (N_29971,N_20053,N_24696);
and U29972 (N_29972,N_24649,N_23368);
nand U29973 (N_29973,N_23853,N_22170);
or U29974 (N_29974,N_21583,N_20941);
and U29975 (N_29975,N_24235,N_20957);
xor U29976 (N_29976,N_20842,N_20098);
xnor U29977 (N_29977,N_23338,N_22360);
xnor U29978 (N_29978,N_22337,N_20437);
and U29979 (N_29979,N_20951,N_22638);
nand U29980 (N_29980,N_23582,N_24693);
and U29981 (N_29981,N_24918,N_21475);
xnor U29982 (N_29982,N_20846,N_24495);
and U29983 (N_29983,N_21058,N_22010);
nand U29984 (N_29984,N_22518,N_24908);
xor U29985 (N_29985,N_24816,N_23091);
or U29986 (N_29986,N_20919,N_22571);
and U29987 (N_29987,N_24159,N_23107);
or U29988 (N_29988,N_20246,N_21227);
or U29989 (N_29989,N_22288,N_24843);
and U29990 (N_29990,N_24075,N_24250);
nor U29991 (N_29991,N_21568,N_24308);
nand U29992 (N_29992,N_23239,N_20881);
and U29993 (N_29993,N_23532,N_22925);
nor U29994 (N_29994,N_21298,N_23503);
nor U29995 (N_29995,N_23254,N_21907);
xor U29996 (N_29996,N_24251,N_23851);
or U29997 (N_29997,N_21985,N_24617);
nand U29998 (N_29998,N_23047,N_23855);
and U29999 (N_29999,N_22649,N_20565);
xnor UO_0 (O_0,N_28238,N_25696);
nand UO_1 (O_1,N_28953,N_27218);
nor UO_2 (O_2,N_29845,N_27528);
and UO_3 (O_3,N_28555,N_27914);
nand UO_4 (O_4,N_26541,N_28370);
nand UO_5 (O_5,N_26677,N_27205);
xor UO_6 (O_6,N_29691,N_26087);
nor UO_7 (O_7,N_26288,N_29987);
and UO_8 (O_8,N_29697,N_27074);
xnor UO_9 (O_9,N_29455,N_27171);
nand UO_10 (O_10,N_25121,N_29238);
nor UO_11 (O_11,N_28703,N_25953);
nand UO_12 (O_12,N_29144,N_27012);
xnor UO_13 (O_13,N_25449,N_27891);
and UO_14 (O_14,N_28835,N_27249);
or UO_15 (O_15,N_26638,N_29486);
and UO_16 (O_16,N_26049,N_27427);
and UO_17 (O_17,N_25137,N_29459);
nand UO_18 (O_18,N_25555,N_29430);
or UO_19 (O_19,N_25367,N_26194);
and UO_20 (O_20,N_26322,N_29873);
and UO_21 (O_21,N_26934,N_26601);
or UO_22 (O_22,N_25721,N_29300);
or UO_23 (O_23,N_25909,N_29299);
or UO_24 (O_24,N_29327,N_26690);
or UO_25 (O_25,N_29470,N_25044);
nor UO_26 (O_26,N_27037,N_29035);
xor UO_27 (O_27,N_27731,N_27335);
xor UO_28 (O_28,N_28795,N_29946);
or UO_29 (O_29,N_26961,N_25285);
and UO_30 (O_30,N_28520,N_29022);
xnor UO_31 (O_31,N_25215,N_27926);
nor UO_32 (O_32,N_29335,N_29159);
and UO_33 (O_33,N_28163,N_26596);
or UO_34 (O_34,N_26767,N_29775);
nor UO_35 (O_35,N_26533,N_29563);
nor UO_36 (O_36,N_27820,N_27388);
nor UO_37 (O_37,N_26667,N_29718);
nor UO_38 (O_38,N_26821,N_27202);
nor UO_39 (O_39,N_27059,N_28450);
xnor UO_40 (O_40,N_27472,N_25875);
xnor UO_41 (O_41,N_28205,N_25673);
nor UO_42 (O_42,N_29654,N_29853);
nand UO_43 (O_43,N_28718,N_28600);
nor UO_44 (O_44,N_29239,N_26800);
nand UO_45 (O_45,N_26815,N_26469);
or UO_46 (O_46,N_28379,N_26010);
xnor UO_47 (O_47,N_29389,N_29284);
and UO_48 (O_48,N_26666,N_25090);
nor UO_49 (O_49,N_27295,N_29085);
xor UO_50 (O_50,N_28235,N_27157);
or UO_51 (O_51,N_28566,N_26905);
nor UO_52 (O_52,N_28498,N_28049);
nor UO_53 (O_53,N_29446,N_26932);
nand UO_54 (O_54,N_26197,N_28920);
nand UO_55 (O_55,N_26594,N_25489);
nand UO_56 (O_56,N_27281,N_25782);
nand UO_57 (O_57,N_26652,N_27756);
or UO_58 (O_58,N_29900,N_25657);
or UO_59 (O_59,N_25799,N_27901);
nor UO_60 (O_60,N_25227,N_29168);
nand UO_61 (O_61,N_27258,N_25779);
or UO_62 (O_62,N_26367,N_29994);
and UO_63 (O_63,N_26226,N_29259);
xor UO_64 (O_64,N_26552,N_27095);
or UO_65 (O_65,N_26656,N_26101);
or UO_66 (O_66,N_29029,N_29972);
nand UO_67 (O_67,N_29793,N_27562);
xor UO_68 (O_68,N_28115,N_28131);
nand UO_69 (O_69,N_26037,N_27390);
nand UO_70 (O_70,N_27821,N_28224);
nand UO_71 (O_71,N_28458,N_25101);
nor UO_72 (O_72,N_25115,N_27878);
or UO_73 (O_73,N_28322,N_29315);
nor UO_74 (O_74,N_29426,N_27723);
or UO_75 (O_75,N_28804,N_25297);
nor UO_76 (O_76,N_27898,N_26181);
nand UO_77 (O_77,N_28505,N_26917);
and UO_78 (O_78,N_27452,N_29700);
and UO_79 (O_79,N_26429,N_26270);
and UO_80 (O_80,N_28992,N_28032);
and UO_81 (O_81,N_27918,N_25607);
or UO_82 (O_82,N_28808,N_25582);
xnor UO_83 (O_83,N_26224,N_25569);
nor UO_84 (O_84,N_26501,N_29161);
or UO_85 (O_85,N_27827,N_25588);
and UO_86 (O_86,N_26833,N_25364);
nor UO_87 (O_87,N_25440,N_26295);
xnor UO_88 (O_88,N_28975,N_26355);
and UO_89 (O_89,N_25506,N_29863);
or UO_90 (O_90,N_25811,N_27481);
or UO_91 (O_91,N_25100,N_28468);
xnor UO_92 (O_92,N_29655,N_26870);
and UO_93 (O_93,N_26175,N_27711);
nor UO_94 (O_94,N_29776,N_26737);
and UO_95 (O_95,N_27771,N_26869);
xor UO_96 (O_96,N_29608,N_25086);
or UO_97 (O_97,N_26949,N_25881);
nor UO_98 (O_98,N_27178,N_25651);
and UO_99 (O_99,N_25703,N_29686);
nor UO_100 (O_100,N_26370,N_27759);
and UO_101 (O_101,N_26188,N_28510);
nor UO_102 (O_102,N_29626,N_26456);
and UO_103 (O_103,N_29541,N_28028);
nor UO_104 (O_104,N_25772,N_29857);
nor UO_105 (O_105,N_25357,N_29616);
or UO_106 (O_106,N_27434,N_25258);
xnor UO_107 (O_107,N_25608,N_25293);
or UO_108 (O_108,N_28276,N_28685);
or UO_109 (O_109,N_25382,N_27988);
nand UO_110 (O_110,N_29865,N_28757);
nor UO_111 (O_111,N_27102,N_28381);
nor UO_112 (O_112,N_25464,N_28169);
xor UO_113 (O_113,N_29796,N_25046);
nor UO_114 (O_114,N_26202,N_27526);
or UO_115 (O_115,N_26482,N_27641);
nand UO_116 (O_116,N_26867,N_26589);
or UO_117 (O_117,N_29534,N_26225);
nor UO_118 (O_118,N_27397,N_26184);
and UO_119 (O_119,N_27986,N_28026);
nand UO_120 (O_120,N_25733,N_25063);
nor UO_121 (O_121,N_28576,N_26222);
or UO_122 (O_122,N_26110,N_29941);
nand UO_123 (O_123,N_26450,N_29832);
nand UO_124 (O_124,N_25337,N_25028);
xnor UO_125 (O_125,N_27063,N_25848);
or UO_126 (O_126,N_27385,N_26699);
nor UO_127 (O_127,N_28193,N_26228);
and UO_128 (O_128,N_26962,N_25004);
nand UO_129 (O_129,N_25565,N_26956);
xor UO_130 (O_130,N_26873,N_28960);
xnor UO_131 (O_131,N_29309,N_27927);
xnor UO_132 (O_132,N_29329,N_29944);
or UO_133 (O_133,N_26984,N_29550);
or UO_134 (O_134,N_25697,N_28110);
xor UO_135 (O_135,N_26365,N_27071);
nand UO_136 (O_136,N_27439,N_27426);
or UO_137 (O_137,N_29514,N_29343);
nand UO_138 (O_138,N_26190,N_26169);
nor UO_139 (O_139,N_29305,N_27964);
nand UO_140 (O_140,N_28832,N_29247);
or UO_141 (O_141,N_29760,N_28504);
and UO_142 (O_142,N_28400,N_26626);
nor UO_143 (O_143,N_28681,N_26102);
or UO_144 (O_144,N_25062,N_26597);
and UO_145 (O_145,N_29033,N_29293);
nor UO_146 (O_146,N_28708,N_25053);
xnor UO_147 (O_147,N_28326,N_27129);
nor UO_148 (O_148,N_29172,N_29543);
xor UO_149 (O_149,N_27230,N_28796);
nand UO_150 (O_150,N_27677,N_29158);
or UO_151 (O_151,N_27140,N_26458);
nor UO_152 (O_152,N_29968,N_28419);
and UO_153 (O_153,N_27318,N_25050);
nor UO_154 (O_154,N_25678,N_29133);
xor UO_155 (O_155,N_25214,N_26358);
xnor UO_156 (O_156,N_28740,N_29767);
nor UO_157 (O_157,N_28754,N_26282);
nor UO_158 (O_158,N_25034,N_26515);
nand UO_159 (O_159,N_28892,N_25975);
and UO_160 (O_160,N_28569,N_28812);
or UO_161 (O_161,N_25150,N_26974);
and UO_162 (O_162,N_29585,N_25778);
or UO_163 (O_163,N_29047,N_28562);
nor UO_164 (O_164,N_26001,N_28060);
nand UO_165 (O_165,N_28319,N_27131);
xor UO_166 (O_166,N_27995,N_25160);
or UO_167 (O_167,N_25240,N_28003);
and UO_168 (O_168,N_25813,N_26980);
nand UO_169 (O_169,N_27703,N_25687);
or UO_170 (O_170,N_26341,N_25809);
xnor UO_171 (O_171,N_25271,N_27273);
and UO_172 (O_172,N_27297,N_29586);
and UO_173 (O_173,N_26850,N_26234);
xnor UO_174 (O_174,N_25596,N_25768);
and UO_175 (O_175,N_25662,N_26292);
or UO_176 (O_176,N_29082,N_25106);
xnor UO_177 (O_177,N_25076,N_28958);
xnor UO_178 (O_178,N_25295,N_28854);
nor UO_179 (O_179,N_28923,N_28233);
nor UO_180 (O_180,N_26535,N_29165);
nand UO_181 (O_181,N_28696,N_25385);
nand UO_182 (O_182,N_25840,N_29289);
nand UO_183 (O_183,N_26381,N_26751);
nor UO_184 (O_184,N_26303,N_27806);
or UO_185 (O_185,N_26035,N_25108);
nand UO_186 (O_186,N_25350,N_28385);
or UO_187 (O_187,N_28340,N_26498);
xnor UO_188 (O_188,N_28102,N_29848);
or UO_189 (O_189,N_25553,N_27045);
nand UO_190 (O_190,N_26513,N_27590);
nor UO_191 (O_191,N_25660,N_25991);
xor UO_192 (O_192,N_25111,N_28291);
nand UO_193 (O_193,N_27116,N_28980);
nand UO_194 (O_194,N_29193,N_28646);
xnor UO_195 (O_195,N_26912,N_27994);
or UO_196 (O_196,N_29531,N_26418);
nand UO_197 (O_197,N_27358,N_26307);
xnor UO_198 (O_198,N_26852,N_26025);
xnor UO_199 (O_199,N_28420,N_25908);
nor UO_200 (O_200,N_29021,N_27517);
nor UO_201 (O_201,N_28219,N_26030);
and UO_202 (O_202,N_29434,N_25427);
xnor UO_203 (O_203,N_25451,N_28616);
or UO_204 (O_204,N_25445,N_25276);
nor UO_205 (O_205,N_25623,N_29366);
and UO_206 (O_206,N_25459,N_25835);
nand UO_207 (O_207,N_26167,N_25784);
and UO_208 (O_208,N_25170,N_26473);
or UO_209 (O_209,N_28273,N_25310);
nor UO_210 (O_210,N_26454,N_29162);
or UO_211 (O_211,N_29003,N_25737);
nor UO_212 (O_212,N_25174,N_28924);
or UO_213 (O_213,N_27279,N_29581);
or UO_214 (O_214,N_26174,N_27149);
nand UO_215 (O_215,N_29245,N_25461);
xnor UO_216 (O_216,N_27316,N_27495);
nand UO_217 (O_217,N_29286,N_29780);
or UO_218 (O_218,N_29904,N_26144);
or UO_219 (O_219,N_29125,N_29668);
or UO_220 (O_220,N_28671,N_26260);
or UO_221 (O_221,N_26470,N_26346);
nor UO_222 (O_222,N_25886,N_27599);
or UO_223 (O_223,N_25021,N_27530);
xnor UO_224 (O_224,N_27367,N_25689);
nor UO_225 (O_225,N_25491,N_26123);
xnor UO_226 (O_226,N_26521,N_27086);
nor UO_227 (O_227,N_29087,N_25573);
nand UO_228 (O_228,N_26308,N_27817);
nand UO_229 (O_229,N_25575,N_27728);
nand UO_230 (O_230,N_29818,N_26388);
xor UO_231 (O_231,N_26318,N_26770);
xor UO_232 (O_232,N_28410,N_29248);
nor UO_233 (O_233,N_27029,N_29516);
nor UO_234 (O_234,N_29601,N_25524);
or UO_235 (O_235,N_26743,N_25612);
nor UO_236 (O_236,N_29886,N_27604);
nor UO_237 (O_237,N_29128,N_29020);
or UO_238 (O_238,N_25722,N_28515);
nor UO_239 (O_239,N_27299,N_25441);
or UO_240 (O_240,N_26608,N_26653);
nor UO_241 (O_241,N_29105,N_28399);
or UO_242 (O_242,N_28056,N_28132);
xor UO_243 (O_243,N_25003,N_29549);
and UO_244 (O_244,N_28974,N_28277);
xor UO_245 (O_245,N_28001,N_29219);
nor UO_246 (O_246,N_25734,N_28814);
nand UO_247 (O_247,N_28043,N_26304);
nor UO_248 (O_248,N_28727,N_29448);
and UO_249 (O_249,N_27490,N_25710);
nand UO_250 (O_250,N_29062,N_29090);
or UO_251 (O_251,N_27863,N_27609);
nand UO_252 (O_252,N_28143,N_27939);
nor UO_253 (O_253,N_25705,N_27253);
nand UO_254 (O_254,N_27169,N_29837);
xnor UO_255 (O_255,N_27608,N_28313);
or UO_256 (O_256,N_28246,N_25676);
or UO_257 (O_257,N_26890,N_29160);
xor UO_258 (O_258,N_26054,N_25430);
and UO_259 (O_259,N_29342,N_29474);
nand UO_260 (O_260,N_27035,N_29226);
and UO_261 (O_261,N_27324,N_25685);
nand UO_262 (O_262,N_27675,N_29617);
nor UO_263 (O_263,N_28155,N_29562);
nand UO_264 (O_264,N_25900,N_27987);
nand UO_265 (O_265,N_29175,N_26200);
nand UO_266 (O_266,N_25262,N_26402);
nand UO_267 (O_267,N_28365,N_28767);
and UO_268 (O_268,N_25526,N_28013);
nor UO_269 (O_269,N_28643,N_26196);
xnor UO_270 (O_270,N_26128,N_28452);
nor UO_271 (O_271,N_27264,N_28464);
nand UO_272 (O_272,N_25644,N_28630);
nand UO_273 (O_273,N_25584,N_27466);
or UO_274 (O_274,N_26803,N_25712);
or UO_275 (O_275,N_28011,N_27651);
nor UO_276 (O_276,N_28429,N_29892);
or UO_277 (O_277,N_26384,N_25518);
or UO_278 (O_278,N_27755,N_28781);
and UO_279 (O_279,N_26543,N_28388);
nor UO_280 (O_280,N_27596,N_26544);
xor UO_281 (O_281,N_29801,N_26462);
and UO_282 (O_282,N_29319,N_28288);
and UO_283 (O_283,N_29618,N_26272);
nand UO_284 (O_284,N_27443,N_25955);
or UO_285 (O_285,N_28380,N_26802);
or UO_286 (O_286,N_28888,N_27550);
and UO_287 (O_287,N_27935,N_27315);
xnor UO_288 (O_288,N_27851,N_25861);
nor UO_289 (O_289,N_25387,N_29424);
xnor UO_290 (O_290,N_29728,N_25147);
or UO_291 (O_291,N_27673,N_29217);
xnor UO_292 (O_292,N_27183,N_25736);
nand UO_293 (O_293,N_26373,N_26909);
or UO_294 (O_294,N_28284,N_25514);
xor UO_295 (O_295,N_28517,N_26701);
nand UO_296 (O_296,N_26259,N_27478);
or UO_297 (O_297,N_26117,N_27201);
nor UO_298 (O_298,N_27573,N_27139);
nand UO_299 (O_299,N_26564,N_28104);
xnor UO_300 (O_300,N_26334,N_25235);
and UO_301 (O_301,N_26960,N_26438);
nand UO_302 (O_302,N_25009,N_26306);
or UO_303 (O_303,N_25473,N_26721);
and UO_304 (O_304,N_29577,N_28112);
or UO_305 (O_305,N_25493,N_26391);
or UO_306 (O_306,N_27189,N_26248);
nor UO_307 (O_307,N_28665,N_26107);
nor UO_308 (O_308,N_26579,N_26636);
or UO_309 (O_309,N_25726,N_28040);
nand UO_310 (O_310,N_26132,N_26165);
xnor UO_311 (O_311,N_28443,N_27482);
or UO_312 (O_312,N_28275,N_27135);
or UO_313 (O_313,N_25587,N_29467);
or UO_314 (O_314,N_28782,N_26790);
nand UO_315 (O_315,N_26941,N_29421);
and UO_316 (O_316,N_29896,N_27525);
nor UO_317 (O_317,N_26674,N_29603);
or UO_318 (O_318,N_28462,N_25424);
nand UO_319 (O_319,N_25475,N_29263);
and UO_320 (O_320,N_28945,N_29742);
or UO_321 (O_321,N_29701,N_28896);
nand UO_322 (O_322,N_29485,N_25810);
or UO_323 (O_323,N_25426,N_26603);
xnor UO_324 (O_324,N_25118,N_28943);
nand UO_325 (O_325,N_27893,N_29212);
or UO_326 (O_326,N_29472,N_29901);
or UO_327 (O_327,N_28034,N_26383);
or UO_328 (O_328,N_28442,N_25503);
and UO_329 (O_329,N_25414,N_27293);
nor UO_330 (O_330,N_28783,N_26265);
xnor UO_331 (O_331,N_26137,N_28647);
or UO_332 (O_332,N_28819,N_25682);
xor UO_333 (O_333,N_26857,N_26403);
or UO_334 (O_334,N_26465,N_27807);
nor UO_335 (O_335,N_25672,N_25610);
nand UO_336 (O_336,N_27666,N_29210);
nand UO_337 (O_337,N_26882,N_26809);
or UO_338 (O_338,N_28145,N_26192);
nand UO_339 (O_339,N_26828,N_29076);
or UO_340 (O_340,N_29827,N_27580);
xor UO_341 (O_341,N_26539,N_27501);
or UO_342 (O_342,N_29526,N_28862);
nor UO_343 (O_343,N_29334,N_29926);
or UO_344 (O_344,N_29321,N_25457);
and UO_345 (O_345,N_28000,N_28651);
nor UO_346 (O_346,N_26162,N_29919);
xnor UO_347 (O_347,N_27799,N_25237);
nand UO_348 (O_348,N_28598,N_29053);
nand UO_349 (O_349,N_28282,N_27812);
nand UO_350 (O_350,N_25648,N_29377);
nand UO_351 (O_351,N_26022,N_28707);
and UO_352 (O_352,N_27797,N_29380);
or UO_353 (O_353,N_27973,N_29754);
nand UO_354 (O_354,N_26179,N_29273);
or UO_355 (O_355,N_26424,N_29184);
nor UO_356 (O_356,N_29348,N_27196);
xnor UO_357 (O_357,N_26204,N_26178);
nor UO_358 (O_358,N_26240,N_27742);
nor UO_359 (O_359,N_26460,N_25042);
nor UO_360 (O_360,N_27393,N_29116);
or UO_361 (O_361,N_29709,N_26777);
xnor UO_362 (O_362,N_29648,N_25333);
xor UO_363 (O_363,N_25329,N_28689);
nor UO_364 (O_364,N_26886,N_27244);
or UO_365 (O_365,N_28371,N_26063);
nor UO_366 (O_366,N_28871,N_25795);
xnor UO_367 (O_367,N_27304,N_28788);
nand UO_368 (O_368,N_26964,N_28077);
and UO_369 (O_369,N_28912,N_29819);
xor UO_370 (O_370,N_27475,N_27614);
or UO_371 (O_371,N_27676,N_26553);
nor UO_372 (O_372,N_26231,N_28969);
xnor UO_373 (O_373,N_29791,N_25636);
nand UO_374 (O_374,N_26710,N_25929);
nor UO_375 (O_375,N_28964,N_25129);
and UO_376 (O_376,N_28876,N_25225);
xnor UO_377 (O_377,N_25674,N_29403);
or UO_378 (O_378,N_26512,N_29822);
or UO_379 (O_379,N_26029,N_27301);
nor UO_380 (O_380,N_27681,N_25856);
and UO_381 (O_381,N_27944,N_25116);
nor UO_382 (O_382,N_25266,N_27360);
xor UO_383 (O_383,N_28702,N_26868);
or UO_384 (O_384,N_27162,N_25085);
and UO_385 (O_385,N_25937,N_29536);
nor UO_386 (O_386,N_27831,N_27702);
nand UO_387 (O_387,N_27032,N_26439);
nand UO_388 (O_388,N_28928,N_29639);
or UO_389 (O_389,N_29318,N_28485);
xnor UO_390 (O_390,N_28167,N_29500);
and UO_391 (O_391,N_28154,N_29503);
nor UO_392 (O_392,N_27379,N_29001);
nand UO_393 (O_393,N_29741,N_25966);
and UO_394 (O_394,N_27764,N_26496);
nand UO_395 (O_395,N_28966,N_29610);
or UO_396 (O_396,N_25932,N_28502);
nand UO_397 (O_397,N_26746,N_25331);
or UO_398 (O_398,N_26431,N_29713);
nand UO_399 (O_399,N_29887,N_27587);
and UO_400 (O_400,N_29340,N_25589);
and UO_401 (O_401,N_27598,N_29042);
xor UO_402 (O_402,N_25056,N_26177);
nor UO_403 (O_403,N_27521,N_27752);
xor UO_404 (O_404,N_27068,N_26935);
nand UO_405 (O_405,N_25438,N_25663);
nand UO_406 (O_406,N_28775,N_25072);
and UO_407 (O_407,N_29658,N_26368);
or UO_408 (O_408,N_29030,N_26831);
nand UO_409 (O_409,N_28318,N_27322);
or UO_410 (O_410,N_29496,N_27122);
and UO_411 (O_411,N_25131,N_28158);
nand UO_412 (O_412,N_25097,N_27127);
nor UO_413 (O_413,N_29561,N_29894);
and UO_414 (O_414,N_28030,N_27084);
xor UO_415 (O_415,N_26269,N_29824);
nor UO_416 (O_416,N_25957,N_28579);
and UO_417 (O_417,N_29740,N_25781);
or UO_418 (O_418,N_28506,N_28108);
xnor UO_419 (O_419,N_29140,N_27663);
xnor UO_420 (O_420,N_26289,N_27809);
nand UO_421 (O_421,N_27730,N_26262);
and UO_422 (O_422,N_28355,N_28401);
xor UO_423 (O_423,N_26399,N_27996);
xnor UO_424 (O_424,N_26058,N_29759);
or UO_425 (O_425,N_28567,N_25926);
nand UO_426 (O_426,N_27446,N_29379);
nand UO_427 (O_427,N_28471,N_25643);
or UO_428 (O_428,N_29049,N_27593);
nor UO_429 (O_429,N_26628,N_27910);
and UO_430 (O_430,N_29778,N_26085);
or UO_431 (O_431,N_28677,N_25155);
and UO_432 (O_432,N_28025,N_28432);
and UO_433 (O_433,N_29489,N_25185);
or UO_434 (O_434,N_29557,N_29565);
xor UO_435 (O_435,N_27700,N_29669);
and UO_436 (O_436,N_25997,N_28500);
or UO_437 (O_437,N_28185,N_25562);
or UO_438 (O_438,N_25910,N_29625);
or UO_439 (O_439,N_27509,N_29027);
xnor UO_440 (O_440,N_29440,N_25967);
xnor UO_441 (O_441,N_25241,N_26452);
or UO_442 (O_442,N_26939,N_26753);
or UO_443 (O_443,N_28454,N_25015);
xor UO_444 (O_444,N_28961,N_27979);
xnor UO_445 (O_445,N_29057,N_26898);
and UO_446 (O_446,N_26419,N_26310);
nor UO_447 (O_447,N_25545,N_29437);
xnor UO_448 (O_448,N_28096,N_28800);
nor UO_449 (O_449,N_27125,N_28343);
nand UO_450 (O_450,N_27533,N_29382);
xnor UO_451 (O_451,N_26766,N_26120);
nor UO_452 (O_452,N_29338,N_25369);
and UO_453 (O_453,N_25352,N_25762);
or UO_454 (O_454,N_26786,N_27349);
or UO_455 (O_455,N_29523,N_27882);
nand UO_456 (O_456,N_27136,N_27929);
nand UO_457 (O_457,N_27552,N_25007);
and UO_458 (O_458,N_27254,N_28846);
nand UO_459 (O_459,N_25231,N_25994);
xnor UO_460 (O_460,N_28861,N_29269);
nor UO_461 (O_461,N_26537,N_29738);
xor UO_462 (O_462,N_26779,N_25070);
nor UO_463 (O_463,N_28247,N_27761);
nor UO_464 (O_464,N_29748,N_26689);
nor UO_465 (O_465,N_26919,N_28303);
or UO_466 (O_466,N_25186,N_29692);
xor UO_467 (O_467,N_25405,N_27652);
and UO_468 (O_468,N_29737,N_27257);
xnor UO_469 (O_469,N_25701,N_29215);
and UO_470 (O_470,N_25775,N_26526);
or UO_471 (O_471,N_28877,N_27107);
or UO_472 (O_472,N_26261,N_26559);
or UO_473 (O_473,N_28117,N_27856);
nand UO_474 (O_474,N_25209,N_26755);
nor UO_475 (O_475,N_25260,N_29736);
xor UO_476 (O_476,N_28111,N_26854);
or UO_477 (O_477,N_27558,N_27883);
nor UO_478 (O_478,N_28254,N_29673);
nand UO_479 (O_479,N_29992,N_26353);
nand UO_480 (O_480,N_26125,N_29990);
nor UO_481 (O_481,N_26442,N_29034);
xnor UO_482 (O_482,N_25264,N_27389);
or UO_483 (O_483,N_25005,N_25330);
nand UO_484 (O_484,N_27020,N_28007);
xor UO_485 (O_485,N_26284,N_28310);
nand UO_486 (O_486,N_27559,N_25363);
or UO_487 (O_487,N_26203,N_27422);
xnor UO_488 (O_488,N_27660,N_28421);
or UO_489 (O_489,N_25247,N_26435);
xnor UO_490 (O_490,N_26880,N_27826);
xnor UO_491 (O_491,N_27765,N_27143);
and UO_492 (O_492,N_27622,N_28490);
nand UO_493 (O_493,N_26256,N_25704);
or UO_494 (O_494,N_25622,N_28907);
nand UO_495 (O_495,N_26915,N_28161);
or UO_496 (O_496,N_28890,N_25802);
or UO_497 (O_497,N_28885,N_27329);
and UO_498 (O_498,N_27298,N_28843);
nand UO_499 (O_499,N_26019,N_25537);
nor UO_500 (O_500,N_26795,N_26807);
or UO_501 (O_501,N_27674,N_29466);
nor UO_502 (O_502,N_27160,N_26508);
and UO_503 (O_503,N_29260,N_28884);
and UO_504 (O_504,N_29689,N_29519);
nor UO_505 (O_505,N_25082,N_26302);
and UO_506 (O_506,N_26255,N_28237);
nor UO_507 (O_507,N_26842,N_27537);
nor UO_508 (O_508,N_27500,N_27184);
nor UO_509 (O_509,N_27965,N_25924);
xor UO_510 (O_510,N_29429,N_29522);
xnor UO_511 (O_511,N_29189,N_28572);
and UO_512 (O_512,N_27081,N_26816);
nor UO_513 (O_513,N_25113,N_28496);
or UO_514 (O_514,N_28157,N_25743);
xor UO_515 (O_515,N_29782,N_27860);
nor UO_516 (O_516,N_28734,N_29469);
xor UO_517 (O_517,N_27924,N_25995);
nand UO_518 (O_518,N_29264,N_25495);
xnor UO_519 (O_519,N_29789,N_27459);
or UO_520 (O_520,N_25444,N_26237);
xnor UO_521 (O_521,N_29011,N_26104);
nor UO_522 (O_522,N_25362,N_25968);
nand UO_523 (O_523,N_27770,N_28712);
xnor UO_524 (O_524,N_27378,N_28827);
nand UO_525 (O_525,N_29449,N_26719);
and UO_526 (O_526,N_25741,N_28830);
nor UO_527 (O_527,N_29488,N_27252);
and UO_528 (O_528,N_27117,N_28501);
or UO_529 (O_529,N_27607,N_26952);
nand UO_530 (O_530,N_26449,N_28552);
nand UO_531 (O_531,N_25962,N_26372);
or UO_532 (O_532,N_25725,N_26422);
nand UO_533 (O_533,N_27085,N_29383);
and UO_534 (O_534,N_28372,N_26468);
nand UO_535 (O_535,N_26033,N_29898);
nand UO_536 (O_536,N_25785,N_27999);
nand UO_537 (O_537,N_26414,N_28204);
nand UO_538 (O_538,N_25755,N_26342);
nor UO_539 (O_539,N_28268,N_25360);
nor UO_540 (O_540,N_27553,N_28127);
nor UO_541 (O_541,N_25328,N_27516);
nand UO_542 (O_542,N_28292,N_27738);
xor UO_543 (O_543,N_26745,N_28751);
nor UO_544 (O_544,N_27621,N_29445);
nand UO_545 (O_545,N_29115,N_28699);
or UO_546 (O_546,N_28839,N_29113);
nand UO_547 (O_547,N_25057,N_28051);
nor UO_548 (O_548,N_29490,N_25500);
nor UO_549 (O_549,N_29411,N_27691);
nand UO_550 (O_550,N_27578,N_25691);
xnor UO_551 (O_551,N_28129,N_27998);
and UO_552 (O_552,N_26976,N_29502);
or UO_553 (O_553,N_29934,N_25838);
or UO_554 (O_554,N_26871,N_27100);
nand UO_555 (O_555,N_29266,N_28359);
nor UO_556 (O_556,N_28455,N_29220);
and UO_557 (O_557,N_26523,N_28722);
xor UO_558 (O_558,N_26154,N_29556);
nand UO_559 (O_559,N_29831,N_27386);
nor UO_560 (O_560,N_25572,N_27172);
and UO_561 (O_561,N_26569,N_26293);
nand UO_562 (O_562,N_29276,N_26718);
nand UO_563 (O_563,N_26472,N_25508);
or UO_564 (O_564,N_29173,N_28672);
and UO_565 (O_565,N_28947,N_29204);
nand UO_566 (O_566,N_28956,N_28136);
xnor UO_567 (O_567,N_25885,N_26349);
nor UO_568 (O_568,N_26834,N_28587);
nor UO_569 (O_569,N_25951,N_26096);
or UO_570 (O_570,N_25378,N_25318);
nand UO_571 (O_571,N_29091,N_25177);
or UO_572 (O_572,N_26671,N_29707);
and UO_573 (O_573,N_26863,N_25980);
xnor UO_574 (O_574,N_28036,N_29346);
nand UO_575 (O_575,N_28239,N_28213);
and UO_576 (O_576,N_28210,N_28467);
nand UO_577 (O_577,N_25550,N_25467);
and UO_578 (O_578,N_29055,N_26811);
and UO_579 (O_579,N_26524,N_26706);
or UO_580 (O_580,N_29180,N_25706);
nor UO_581 (O_581,N_25758,N_29629);
or UO_582 (O_582,N_27502,N_25554);
xnor UO_583 (O_583,N_27680,N_26499);
nor UO_584 (O_584,N_26404,N_25591);
or UO_585 (O_585,N_29254,N_28621);
nor UO_586 (O_586,N_29296,N_25770);
or UO_587 (O_587,N_26208,N_29364);
and UO_588 (O_588,N_28695,N_27232);
or UO_589 (O_589,N_29513,N_27123);
xor UO_590 (O_590,N_29907,N_26650);
nand UO_591 (O_591,N_26778,N_25808);
nor UO_592 (O_592,N_28825,N_29839);
nor UO_593 (O_593,N_25409,N_28666);
or UO_594 (O_594,N_27876,N_26206);
nor UO_595 (O_595,N_25190,N_29535);
or UO_596 (O_596,N_27698,N_26928);
xor UO_597 (O_597,N_29080,N_27520);
or UO_598 (O_598,N_29590,N_25857);
xnor UO_599 (O_599,N_26958,N_25080);
xor UO_600 (O_600,N_26480,N_25091);
nand UO_601 (O_601,N_27028,N_28258);
and UO_602 (O_602,N_26055,N_29255);
nand UO_603 (O_603,N_28889,N_25477);
xnor UO_604 (O_604,N_27888,N_26220);
or UO_605 (O_605,N_28852,N_29607);
nor UO_606 (O_606,N_25233,N_29982);
or UO_607 (O_607,N_27331,N_29404);
nor UO_608 (O_608,N_28618,N_28847);
or UO_609 (O_609,N_28064,N_25187);
and UO_610 (O_610,N_28017,N_25166);
xnor UO_611 (O_611,N_28955,N_26697);
and UO_612 (O_612,N_28391,N_26799);
or UO_613 (O_613,N_26648,N_29725);
and UO_614 (O_614,N_26091,N_25059);
or UO_615 (O_615,N_29921,N_29632);
or UO_616 (O_616,N_29277,N_27276);
nor UO_617 (O_617,N_29287,N_27611);
nor UO_618 (O_618,N_28350,N_29595);
nand UO_619 (O_619,N_28358,N_29142);
or UO_620 (O_620,N_25964,N_28570);
or UO_621 (O_621,N_29785,N_29533);
and UO_622 (O_622,N_29064,N_28690);
nand UO_623 (O_623,N_27941,N_29362);
and UO_624 (O_624,N_28818,N_26233);
or UO_625 (O_625,N_29758,N_28608);
nand UO_626 (O_626,N_27793,N_28218);
and UO_627 (O_627,N_27777,N_28709);
or UO_628 (O_628,N_26378,N_25040);
nor UO_629 (O_629,N_28543,N_25393);
or UO_630 (O_630,N_28267,N_28897);
nand UO_631 (O_631,N_25944,N_28873);
nand UO_632 (O_632,N_26474,N_27338);
xor UO_633 (O_633,N_25316,N_25096);
nor UO_634 (O_634,N_27519,N_25157);
or UO_635 (O_635,N_27348,N_25641);
or UO_636 (O_636,N_28134,N_28586);
xor UO_637 (O_637,N_25306,N_26122);
and UO_638 (O_638,N_26660,N_26632);
or UO_639 (O_639,N_25940,N_28918);
nor UO_640 (O_640,N_27073,N_26395);
or UO_641 (O_641,N_29636,N_28250);
xnor UO_642 (O_642,N_29576,N_29480);
xnor UO_643 (O_643,N_28774,N_28470);
and UO_644 (O_644,N_25273,N_29794);
and UO_645 (O_645,N_25659,N_27591);
or UO_646 (O_646,N_29333,N_25000);
and UO_647 (O_647,N_27671,N_26116);
xor UO_648 (O_648,N_27656,N_25763);
nor UO_649 (O_649,N_29132,N_28440);
or UO_650 (O_650,N_25898,N_25110);
nand UO_651 (O_651,N_25067,N_29570);
and UO_652 (O_652,N_25533,N_26772);
or UO_653 (O_653,N_26313,N_26810);
or UO_654 (O_654,N_28589,N_26605);
or UO_655 (O_655,N_28279,N_26607);
nand UO_656 (O_656,N_26971,N_27000);
nor UO_657 (O_657,N_28212,N_26115);
nor UO_658 (O_658,N_26028,N_28753);
xor UO_659 (O_659,N_29152,N_25023);
or UO_660 (O_660,N_25877,N_27488);
nand UO_661 (O_661,N_27869,N_29391);
nand UO_662 (O_662,N_26506,N_27704);
and UO_663 (O_663,N_25019,N_26897);
xnor UO_664 (O_664,N_26386,N_28609);
xor UO_665 (O_665,N_26351,N_27819);
nor UO_666 (O_666,N_27772,N_26332);
nor UO_667 (O_667,N_27450,N_25436);
or UO_668 (O_668,N_25071,N_26981);
and UO_669 (O_669,N_27133,N_29007);
or UO_670 (O_670,N_29871,N_27374);
and UO_671 (O_671,N_29866,N_28556);
or UO_672 (O_672,N_26039,N_26965);
and UO_673 (O_673,N_25728,N_27104);
or UO_674 (O_674,N_27395,N_27413);
nand UO_675 (O_675,N_27239,N_27250);
xor UO_676 (O_676,N_25780,N_29574);
xnor UO_677 (O_677,N_28551,N_26545);
nand UO_678 (O_678,N_27707,N_25277);
nor UO_679 (O_679,N_27346,N_28613);
nand UO_680 (O_680,N_25801,N_27341);
xor UO_681 (O_681,N_27997,N_29119);
or UO_682 (O_682,N_27906,N_29963);
xnor UO_683 (O_683,N_29288,N_28475);
or UO_684 (O_684,N_28195,N_29928);
nand UO_685 (O_685,N_25774,N_26056);
xor UO_686 (O_686,N_26051,N_27256);
nor UO_687 (O_687,N_28536,N_27286);
nand UO_688 (O_688,N_28124,N_25248);
or UO_689 (O_689,N_25078,N_27498);
xor UO_690 (O_690,N_25354,N_28487);
nand UO_691 (O_691,N_28721,N_26788);
nand UO_692 (O_692,N_26077,N_26083);
and UO_693 (O_693,N_29752,N_27938);
nor UO_694 (O_694,N_25434,N_29812);
nand UO_695 (O_695,N_26159,N_25880);
nor UO_696 (O_696,N_29704,N_26970);
nor UO_697 (O_697,N_28393,N_27152);
xor UO_698 (O_698,N_29317,N_26407);
xnor UO_699 (O_699,N_28465,N_27945);
and UO_700 (O_700,N_26189,N_29641);
xnor UO_701 (O_701,N_25549,N_27231);
and UO_702 (O_702,N_28300,N_27420);
nand UO_703 (O_703,N_25020,N_28747);
and UO_704 (O_704,N_27602,N_29527);
nand UO_705 (O_705,N_26139,N_25411);
nand UO_706 (O_706,N_25894,N_26567);
and UO_707 (O_707,N_26210,N_27483);
nor UO_708 (O_708,N_27515,N_27017);
nand UO_709 (O_709,N_28236,N_27991);
xor UO_710 (O_710,N_27804,N_29249);
and UO_711 (O_711,N_27234,N_29661);
and UO_712 (O_712,N_27757,N_29414);
xnor UO_713 (O_713,N_26557,N_28121);
or UO_714 (O_714,N_27853,N_27949);
nor UO_715 (O_715,N_29110,N_28577);
nand UO_716 (O_716,N_25421,N_25595);
and UO_717 (O_717,N_29451,N_26073);
or UO_718 (O_718,N_26574,N_27108);
nand UO_719 (O_719,N_27586,N_29815);
or UO_720 (O_720,N_28405,N_26611);
nor UO_721 (O_721,N_26698,N_28002);
and UO_722 (O_722,N_26443,N_26774);
nand UO_723 (O_723,N_28750,N_27636);
or UO_724 (O_724,N_27147,N_28164);
and UO_725 (O_725,N_29409,N_25542);
and UO_726 (O_726,N_29745,N_27810);
and UO_727 (O_727,N_28460,N_26445);
or UO_728 (O_728,N_28211,N_27209);
and UO_729 (O_729,N_27203,N_29773);
nor UO_730 (O_730,N_29991,N_29202);
nor UO_731 (O_731,N_27565,N_25730);
and UO_732 (O_732,N_29267,N_25342);
or UO_733 (O_733,N_28459,N_27428);
xor UO_734 (O_734,N_29274,N_28597);
nor UO_735 (O_735,N_26781,N_25124);
xnor UO_736 (O_736,N_27740,N_28408);
nor UO_737 (O_737,N_26630,N_25917);
nor UO_738 (O_738,N_28050,N_25637);
nor UO_739 (O_739,N_25844,N_25876);
and UO_740 (O_740,N_26455,N_28412);
xnor UO_741 (O_741,N_28741,N_26166);
xnor UO_742 (O_742,N_25482,N_28585);
and UO_743 (O_743,N_26088,N_26312);
or UO_744 (O_744,N_28222,N_28637);
or UO_745 (O_745,N_27679,N_25825);
xnor UO_746 (O_746,N_26625,N_25510);
nor UO_747 (O_747,N_28674,N_25729);
or UO_748 (O_748,N_29197,N_29962);
nor UO_749 (O_749,N_29123,N_27263);
and UO_750 (O_750,N_28771,N_26356);
or UO_751 (O_751,N_26441,N_28149);
nor UO_752 (O_752,N_25903,N_25504);
xor UO_753 (O_753,N_26783,N_27845);
or UO_754 (O_754,N_28801,N_29587);
xnor UO_755 (O_755,N_25642,N_26722);
nor UO_756 (O_756,N_27334,N_26299);
nand UO_757 (O_757,N_25098,N_28635);
xnor UO_758 (O_758,N_28075,N_25650);
xnor UO_759 (O_759,N_25356,N_27146);
or UO_760 (O_760,N_27534,N_27556);
or UO_761 (O_761,N_25632,N_25171);
and UO_762 (O_762,N_28856,N_28976);
nand UO_763 (O_763,N_25012,N_26972);
and UO_764 (O_764,N_26094,N_29947);
nand UO_765 (O_765,N_26572,N_25192);
nand UO_766 (O_766,N_26230,N_25724);
and UO_767 (O_767,N_27892,N_25165);
nor UO_768 (O_768,N_25915,N_29730);
or UO_769 (O_769,N_28021,N_27958);
and UO_770 (O_770,N_29860,N_26263);
or UO_771 (O_771,N_29073,N_26340);
and UO_772 (O_772,N_26043,N_28434);
xnor UO_773 (O_773,N_29957,N_25038);
and UO_774 (O_774,N_25646,N_26420);
xnor UO_775 (O_775,N_27199,N_27846);
nand UO_776 (O_776,N_25244,N_28398);
nor UO_777 (O_777,N_28148,N_28287);
nand UO_778 (O_778,N_29710,N_28761);
xnor UO_779 (O_779,N_26813,N_28525);
or UO_780 (O_780,N_28999,N_26542);
or UO_781 (O_781,N_27392,N_28626);
nand UO_782 (O_782,N_28508,N_27091);
nor UO_783 (O_783,N_29065,N_25407);
or UO_784 (O_784,N_28760,N_26151);
and UO_785 (O_785,N_28346,N_29914);
xor UO_786 (O_786,N_28954,N_27855);
nor UO_787 (O_787,N_27916,N_28448);
nor UO_788 (O_788,N_25617,N_25727);
or UO_789 (O_789,N_29281,N_29088);
nand UO_790 (O_790,N_28676,N_25788);
nand UO_791 (O_791,N_29181,N_28269);
or UO_792 (O_792,N_26610,N_26736);
or UO_793 (O_793,N_26959,N_28479);
xor UO_794 (O_794,N_28617,N_28101);
nor UO_795 (O_795,N_29929,N_25911);
nor UO_796 (O_796,N_28069,N_28374);
and UO_797 (O_797,N_28334,N_28528);
and UO_798 (O_798,N_29178,N_28008);
xnor UO_799 (O_799,N_27285,N_29179);
nor UO_800 (O_800,N_26074,N_27406);
nor UO_801 (O_801,N_28762,N_27153);
nor UO_802 (O_802,N_29835,N_28144);
nand UO_803 (O_803,N_26437,N_25487);
nand UO_804 (O_804,N_28090,N_27654);
and UO_805 (O_805,N_29913,N_28870);
xor UO_806 (O_806,N_26111,N_27760);
nand UO_807 (O_807,N_29083,N_28230);
and UO_808 (O_808,N_29802,N_29771);
nand UO_809 (O_809,N_27119,N_28926);
and UO_810 (O_810,N_29599,N_27105);
and UO_811 (O_811,N_26245,N_28328);
and UO_812 (O_812,N_27235,N_26103);
or UO_813 (O_813,N_27842,N_28872);
nor UO_814 (O_814,N_29937,N_29664);
nand UO_815 (O_815,N_29156,N_28395);
and UO_816 (O_816,N_28497,N_25359);
nor UO_817 (O_817,N_28191,N_26294);
nor UO_818 (O_818,N_28542,N_29194);
and UO_819 (O_819,N_29952,N_28680);
xor UO_820 (O_820,N_26851,N_28335);
or UO_821 (O_821,N_28638,N_27384);
nand UO_822 (O_822,N_26347,N_25977);
or UO_823 (O_823,N_26902,N_25052);
xnor UO_824 (O_824,N_28995,N_26683);
xor UO_825 (O_825,N_28176,N_27937);
and UO_826 (O_826,N_29498,N_26007);
nor UO_827 (O_827,N_25420,N_29787);
and UO_828 (O_828,N_27527,N_29207);
or UO_829 (O_829,N_29878,N_29439);
nor UO_830 (O_830,N_28733,N_25583);
xnor UO_831 (O_831,N_27259,N_26002);
nand UO_832 (O_832,N_26005,N_25008);
xnor UO_833 (O_833,N_29660,N_28331);
nor UO_834 (O_834,N_25684,N_26013);
or UO_835 (O_835,N_28826,N_29208);
or UO_836 (O_836,N_25745,N_26339);
nor UO_837 (O_837,N_27693,N_29242);
nand UO_838 (O_838,N_29094,N_29099);
nand UO_839 (O_839,N_29885,N_26872);
nor UO_840 (O_840,N_28667,N_26938);
nor UO_841 (O_841,N_27726,N_27921);
and UO_842 (O_842,N_26629,N_25439);
and UO_843 (O_843,N_26273,N_29923);
or UO_844 (O_844,N_26408,N_28661);
nor UO_845 (O_845,N_28012,N_27371);
xnor UO_846 (O_846,N_27188,N_29882);
nor UO_847 (O_847,N_28731,N_28207);
nand UO_848 (O_848,N_27626,N_29138);
nand UO_849 (O_849,N_28725,N_27717);
and UO_850 (O_850,N_29997,N_26804);
or UO_851 (O_851,N_29983,N_26138);
and UO_852 (O_852,N_25647,N_28984);
or UO_853 (O_853,N_29931,N_27634);
xnor UO_854 (O_854,N_29890,N_26829);
nor UO_855 (O_855,N_29508,N_27690);
or UO_856 (O_856,N_25718,N_29463);
or UO_857 (O_857,N_29188,N_27083);
xnor UO_858 (O_858,N_25272,N_27966);
nand UO_859 (O_859,N_28917,N_28234);
nand UO_860 (O_860,N_26943,N_26348);
or UO_861 (O_861,N_28192,N_28438);
or UO_862 (O_862,N_26791,N_28338);
nand UO_863 (O_863,N_25323,N_25390);
or UO_864 (O_864,N_28841,N_28092);
xor UO_865 (O_865,N_28732,N_26018);
or UO_866 (O_866,N_27486,N_27214);
nand UO_867 (O_867,N_26859,N_25523);
nor UO_868 (O_868,N_27266,N_29653);
nor UO_869 (O_869,N_26691,N_28794);
and UO_870 (O_870,N_25576,N_28086);
nand UO_871 (O_871,N_26801,N_29515);
nor UO_872 (O_872,N_29528,N_28855);
or UO_873 (O_873,N_26153,N_27992);
xor UO_874 (O_874,N_28559,N_28998);
nor UO_875 (O_875,N_28251,N_27404);
nand UO_876 (O_876,N_25292,N_28325);
nor UO_877 (O_877,N_27271,N_29390);
and UO_878 (O_878,N_27735,N_26510);
nor UO_879 (O_879,N_25918,N_28991);
and UO_880 (O_880,N_25852,N_25351);
nand UO_881 (O_881,N_27441,N_25027);
or UO_882 (O_882,N_26711,N_27811);
nor UO_883 (O_883,N_28182,N_29387);
nor UO_884 (O_884,N_27243,N_25036);
nor UO_885 (O_885,N_26891,N_28035);
xnor UO_886 (O_886,N_27889,N_25895);
or UO_887 (O_887,N_25792,N_26631);
xor UO_888 (O_888,N_26241,N_29044);
and UO_889 (O_889,N_29524,N_29392);
xnor UO_890 (O_890,N_27303,N_28905);
nor UO_891 (O_891,N_25184,N_26050);
nor UO_892 (O_892,N_28772,N_28324);
or UO_893 (O_893,N_27454,N_29015);
xnor UO_894 (O_894,N_28748,N_25453);
xnor UO_895 (O_895,N_25982,N_28682);
nor UO_896 (O_896,N_28407,N_26908);
xor UO_897 (O_897,N_25930,N_28738);
nand UO_898 (O_898,N_28053,N_28809);
nand UO_899 (O_899,N_29419,N_25018);
nand UO_900 (O_900,N_25089,N_27103);
and UO_901 (O_901,N_28684,N_25289);
and UO_902 (O_902,N_27192,N_28105);
nand UO_903 (O_903,N_25904,N_28316);
or UO_904 (O_904,N_26780,N_27638);
nand UO_905 (O_905,N_25827,N_28070);
xor UO_906 (O_906,N_29059,N_25948);
nand UO_907 (O_907,N_29621,N_29698);
or UO_908 (O_908,N_29545,N_27978);
and UO_909 (O_909,N_29955,N_27368);
and UO_910 (O_910,N_28240,N_25821);
xor UO_911 (O_911,N_29679,N_29344);
nand UO_912 (O_912,N_29988,N_25942);
or UO_913 (O_913,N_25959,N_26848);
or UO_914 (O_914,N_25887,N_29897);
nand UO_915 (O_915,N_29600,N_25334);
xnor UO_916 (O_916,N_29271,N_26808);
xnor UO_917 (O_917,N_29285,N_25638);
nor UO_918 (O_918,N_29218,N_26173);
or UO_919 (O_919,N_29627,N_26830);
nor UO_920 (O_920,N_26847,N_28138);
or UO_921 (O_921,N_25671,N_28038);
xnor UO_922 (O_922,N_26993,N_29695);
xor UO_923 (O_923,N_29766,N_27983);
xor UO_924 (O_924,N_27850,N_26979);
nor UO_925 (O_925,N_27568,N_26195);
or UO_926 (O_926,N_29539,N_28529);
nor UO_927 (O_927,N_29114,N_26827);
and UO_928 (O_928,N_25343,N_28527);
nor UO_929 (O_929,N_29762,N_29229);
nand UO_930 (O_930,N_25102,N_27433);
xor UO_931 (O_931,N_28894,N_28027);
or UO_932 (O_932,N_27411,N_28323);
nand UO_933 (O_933,N_27226,N_25347);
nor UO_934 (O_934,N_28076,N_25479);
and UO_935 (O_935,N_28387,N_29117);
nand UO_936 (O_936,N_26991,N_27212);
nor UO_937 (O_937,N_28491,N_29611);
nor UO_938 (O_938,N_29985,N_28209);
nand UO_939 (O_939,N_28764,N_26146);
and UO_940 (O_940,N_27313,N_26734);
nor UO_941 (O_941,N_27321,N_29507);
xnor UO_942 (O_942,N_28298,N_26466);
or UO_943 (O_943,N_29927,N_28296);
nor UO_944 (O_944,N_29650,N_26158);
and UO_945 (O_945,N_26969,N_29699);
and UO_946 (O_946,N_27034,N_29996);
or UO_947 (O_947,N_28368,N_26733);
nor UO_948 (O_948,N_26663,N_28549);
nand UO_949 (O_949,N_27824,N_25965);
nand UO_950 (O_950,N_25606,N_28231);
and UO_951 (O_951,N_29657,N_29491);
nor UO_952 (O_952,N_29604,N_28486);
nand UO_953 (O_953,N_26841,N_26876);
nor UO_954 (O_954,N_28194,N_26182);
or UO_955 (O_955,N_26118,N_28792);
nand UO_956 (O_956,N_25077,N_28831);
and UO_957 (O_957,N_25372,N_25014);
nand UO_958 (O_958,N_29394,N_25144);
and UO_959 (O_959,N_29244,N_28189);
or UO_960 (O_960,N_27540,N_25084);
nand UO_961 (O_961,N_25164,N_27942);
nand UO_962 (O_962,N_28320,N_25891);
nand UO_963 (O_963,N_25851,N_25103);
and UO_964 (O_964,N_25458,N_29004);
nand UO_965 (O_965,N_26092,N_27026);
xor UO_966 (O_966,N_28180,N_28437);
xnor UO_967 (O_967,N_29232,N_25973);
nor UO_968 (O_968,N_27078,N_25598);
xnor UO_969 (O_969,N_29719,N_25958);
xnor UO_970 (O_970,N_25379,N_25590);
or UO_971 (O_971,N_25654,N_26525);
or UO_972 (O_972,N_25158,N_25655);
xnor UO_973 (O_973,N_28773,N_27507);
xnor UO_974 (O_974,N_28057,N_29569);
nand UO_975 (O_975,N_27200,N_25145);
or UO_976 (O_976,N_25138,N_27217);
and UO_977 (O_977,N_27403,N_29331);
nor UO_978 (O_978,N_25092,N_26627);
xnor UO_979 (O_979,N_27167,N_25901);
or UO_980 (O_980,N_27727,N_26421);
nand UO_981 (O_981,N_25068,N_26727);
and UO_982 (O_982,N_28135,N_27323);
or UO_983 (O_983,N_27610,N_27213);
and UO_984 (O_984,N_26738,N_29041);
nand UO_985 (O_985,N_25899,N_26027);
or UO_986 (O_986,N_26840,N_28241);
nor UO_987 (O_987,N_25026,N_26413);
and UO_988 (O_988,N_28880,N_27142);
and UO_989 (O_989,N_29372,N_28940);
or UO_990 (O_990,N_28866,N_26004);
nor UO_991 (O_991,N_27957,N_28908);
nor UO_992 (O_992,N_27002,N_27174);
and UO_993 (O_993,N_26749,N_28593);
or UO_994 (O_994,N_29540,N_28197);
nor UO_995 (O_995,N_29084,N_28899);
and UO_996 (O_996,N_26659,N_29790);
or UO_997 (O_997,N_26536,N_28749);
and UO_998 (O_998,N_27376,N_28752);
or UO_999 (O_999,N_26489,N_28147);
nor UO_1000 (O_1000,N_26921,N_28710);
xnor UO_1001 (O_1001,N_26686,N_29016);
and UO_1002 (O_1002,N_25159,N_27745);
and UO_1003 (O_1003,N_25313,N_26032);
nand UO_1004 (O_1004,N_28547,N_25925);
nor UO_1005 (O_1005,N_25579,N_25578);
nor UO_1006 (O_1006,N_28172,N_25670);
and UO_1007 (O_1007,N_27242,N_27685);
or UO_1008 (O_1008,N_26947,N_29056);
and UO_1009 (O_1009,N_29240,N_26853);
xor UO_1010 (O_1010,N_28623,N_26114);
or UO_1011 (O_1011,N_29257,N_26075);
nor UO_1012 (O_1012,N_25298,N_26726);
and UO_1013 (O_1013,N_29492,N_29642);
nor UO_1014 (O_1014,N_26999,N_29487);
xnor UO_1015 (O_1015,N_28916,N_25874);
nor UO_1016 (O_1016,N_26773,N_27040);
nand UO_1017 (O_1017,N_26183,N_25709);
nor UO_1018 (O_1018,N_29844,N_26978);
or UO_1019 (O_1019,N_29756,N_25253);
and UO_1020 (O_1020,N_27504,N_28347);
or UO_1021 (O_1021,N_27126,N_29385);
nor UO_1022 (O_1022,N_28376,N_25580);
nor UO_1023 (O_1023,N_26119,N_25934);
nor UO_1024 (O_1024,N_26664,N_27222);
or UO_1025 (O_1025,N_25597,N_28962);
nand UO_1026 (O_1026,N_27976,N_27198);
xnor UO_1027 (O_1027,N_28988,N_27060);
or UO_1028 (O_1028,N_26942,N_28700);
xor UO_1029 (O_1029,N_26742,N_29241);
xor UO_1030 (O_1030,N_25558,N_29118);
nand UO_1031 (O_1031,N_25478,N_28978);
or UO_1032 (O_1032,N_26385,N_29578);
nor UO_1033 (O_1033,N_29292,N_26588);
xor UO_1034 (O_1034,N_29295,N_29093);
xor UO_1035 (O_1035,N_27541,N_28242);
and UO_1036 (O_1036,N_25817,N_28302);
or UO_1037 (O_1037,N_27524,N_27603);
nor UO_1038 (O_1038,N_28972,N_26319);
xnor UO_1039 (O_1039,N_25093,N_25945);
and UO_1040 (O_1040,N_27005,N_27776);
nand UO_1041 (O_1041,N_25816,N_29283);
xnor UO_1042 (O_1042,N_26301,N_25791);
nor UO_1043 (O_1043,N_27047,N_26590);
xnor UO_1044 (O_1044,N_25547,N_28228);
nor UO_1045 (O_1045,N_26130,N_28171);
nor UO_1046 (O_1046,N_25540,N_27963);
nand UO_1047 (O_1047,N_27721,N_28390);
nand UO_1048 (O_1048,N_27087,N_28297);
or UO_1049 (O_1049,N_26992,N_25757);
nand UO_1050 (O_1050,N_29750,N_29930);
xor UO_1051 (O_1051,N_28023,N_27545);
or UO_1052 (O_1052,N_25618,N_28997);
nand UO_1053 (O_1053,N_26883,N_27150);
nor UO_1054 (O_1054,N_25088,N_26006);
nor UO_1055 (O_1055,N_25502,N_29765);
nor UO_1056 (O_1056,N_28047,N_26712);
and UO_1057 (O_1057,N_27134,N_27601);
and UO_1058 (O_1058,N_25624,N_25872);
and UO_1059 (O_1059,N_29149,N_29129);
xnor UO_1060 (O_1060,N_29659,N_25707);
nor UO_1061 (O_1061,N_29628,N_27859);
nand UO_1062 (O_1062,N_28829,N_29917);
nor UO_1063 (O_1063,N_26702,N_26352);
nand UO_1064 (O_1064,N_28369,N_27251);
nor UO_1065 (O_1065,N_25287,N_28083);
or UO_1066 (O_1066,N_27090,N_29442);
and UO_1067 (O_1067,N_25574,N_25832);
nor UO_1068 (O_1068,N_27260,N_26731);
and UO_1069 (O_1069,N_29684,N_26835);
and UO_1070 (O_1070,N_26546,N_28533);
and UO_1071 (O_1071,N_28140,N_25567);
nor UO_1072 (O_1072,N_27186,N_25265);
or UO_1073 (O_1073,N_25047,N_27689);
nand UO_1074 (O_1074,N_29150,N_27984);
nor UO_1075 (O_1075,N_26447,N_26502);
or UO_1076 (O_1076,N_27332,N_29324);
or UO_1077 (O_1077,N_27391,N_29211);
xor UO_1078 (O_1078,N_29779,N_27781);
nor UO_1079 (O_1079,N_25831,N_27861);
nor UO_1080 (O_1080,N_28848,N_26641);
xnor UO_1081 (O_1081,N_25213,N_27968);
or UO_1082 (O_1082,N_28348,N_28952);
and UO_1083 (O_1083,N_28833,N_29956);
or UO_1084 (O_1084,N_27544,N_28820);
or UO_1085 (O_1085,N_28986,N_26236);
nand UO_1086 (O_1086,N_29870,N_29497);
or UO_1087 (O_1087,N_25754,N_26657);
nor UO_1088 (O_1088,N_28706,N_25677);
nand UO_1089 (O_1089,N_25279,N_26155);
and UO_1090 (O_1090,N_27158,N_28604);
or UO_1091 (O_1091,N_28822,N_27132);
or UO_1092 (O_1092,N_25470,N_25206);
nor UO_1093 (O_1093,N_25060,N_25974);
xnor UO_1094 (O_1094,N_26658,N_29544);
or UO_1095 (O_1095,N_28564,N_29357);
or UO_1096 (O_1096,N_26359,N_26587);
nor UO_1097 (O_1097,N_28285,N_28605);
nand UO_1098 (O_1098,N_28378,N_26267);
and UO_1099 (O_1099,N_25255,N_26031);
or UO_1100 (O_1100,N_27030,N_27695);
and UO_1101 (O_1101,N_28615,N_26250);
xnor UO_1102 (O_1102,N_29397,N_26614);
nand UO_1103 (O_1103,N_28174,N_27072);
or UO_1104 (O_1104,N_27872,N_28919);
nor UO_1105 (O_1105,N_25751,N_28392);
and UO_1106 (O_1106,N_26760,N_25529);
nor UO_1107 (O_1107,N_29732,N_27911);
xnor UO_1108 (O_1108,N_26345,N_26152);
xor UO_1109 (O_1109,N_29332,N_29237);
nor UO_1110 (O_1110,N_27484,N_25471);
nor UO_1111 (O_1111,N_26276,N_29918);
or UO_1112 (O_1112,N_25256,N_29107);
and UO_1113 (O_1113,N_26794,N_29712);
or UO_1114 (O_1114,N_27325,N_25916);
and UO_1115 (O_1115,N_25245,N_27007);
nand UO_1116 (O_1116,N_26497,N_26843);
nand UO_1117 (O_1117,N_29989,N_27623);
nand UO_1118 (O_1118,N_25920,N_25806);
and UO_1119 (O_1119,N_26362,N_28196);
nand UO_1120 (O_1120,N_25229,N_26575);
nand UO_1121 (O_1121,N_26433,N_29975);
nor UO_1122 (O_1122,N_26291,N_29402);
nor UO_1123 (O_1123,N_29935,N_28015);
and UO_1124 (O_1124,N_28107,N_27027);
nand UO_1125 (O_1125,N_28875,N_29879);
xnor UO_1126 (O_1126,N_28509,N_27175);
nand UO_1127 (O_1127,N_29518,N_29396);
and UO_1128 (O_1128,N_26983,N_27631);
nand UO_1129 (O_1129,N_28963,N_27019);
nor UO_1130 (O_1130,N_28935,N_27067);
and UO_1131 (O_1131,N_29398,N_26592);
nor UO_1132 (O_1132,N_26082,N_26892);
xnor UO_1133 (O_1133,N_25167,N_28416);
nor UO_1134 (O_1134,N_27787,N_28599);
nand UO_1135 (O_1135,N_26495,N_27880);
or UO_1136 (O_1136,N_28628,N_29501);
or UO_1137 (O_1137,N_28321,N_29783);
nor UO_1138 (O_1138,N_28759,N_29417);
or UO_1139 (O_1139,N_28444,N_27410);
nor UO_1140 (O_1140,N_27549,N_27647);
or UO_1141 (O_1141,N_26814,N_29031);
or UO_1142 (O_1142,N_26042,N_29602);
and UO_1143 (O_1143,N_26099,N_26215);
or UO_1144 (O_1144,N_26487,N_26948);
and UO_1145 (O_1145,N_25134,N_26558);
nand UO_1146 (O_1146,N_25132,N_28068);
and UO_1147 (O_1147,N_25442,N_26500);
or UO_1148 (O_1148,N_29071,N_25604);
nor UO_1149 (O_1149,N_26223,N_27884);
nand UO_1150 (O_1150,N_29724,N_26822);
and UO_1151 (O_1151,N_26321,N_25544);
or UO_1152 (O_1152,N_25228,N_26668);
nor UO_1153 (O_1153,N_28691,N_26164);
nor UO_1154 (O_1154,N_26817,N_29388);
or UO_1155 (O_1155,N_27461,N_29013);
nor UO_1156 (O_1156,N_25850,N_29095);
nor UO_1157 (O_1157,N_25226,N_28511);
nand UO_1158 (O_1158,N_27288,N_26268);
nand UO_1159 (O_1159,N_25969,N_27669);
nand UO_1160 (O_1160,N_29948,N_28625);
or UO_1161 (O_1161,N_25715,N_26717);
nor UO_1162 (O_1162,N_28717,N_27262);
and UO_1163 (O_1163,N_29222,N_28850);
and UO_1164 (O_1164,N_26540,N_29788);
nor UO_1165 (O_1165,N_29644,N_27261);
xor UO_1166 (O_1166,N_25447,N_29272);
nand UO_1167 (O_1167,N_29572,N_28198);
nor UO_1168 (O_1168,N_27282,N_25868);
xnor UO_1169 (O_1169,N_26205,N_25818);
xor UO_1170 (O_1170,N_27692,N_25312);
xor UO_1171 (O_1171,N_28133,N_29376);
nor UO_1172 (O_1172,N_28375,N_27487);
nand UO_1173 (O_1173,N_25854,N_25747);
nand UO_1174 (O_1174,N_26448,N_26577);
nor UO_1175 (O_1175,N_27361,N_25865);
and UO_1176 (O_1176,N_25683,N_25773);
and UO_1177 (O_1177,N_26081,N_29354);
and UO_1178 (O_1178,N_28603,N_26693);
xor UO_1179 (O_1179,N_26729,N_25708);
and UO_1180 (O_1180,N_29743,N_26534);
and UO_1181 (O_1181,N_26899,N_25667);
and UO_1182 (O_1182,N_27605,N_26316);
nand UO_1183 (O_1183,N_26624,N_25928);
or UO_1184 (O_1184,N_29720,N_26730);
and UO_1185 (O_1185,N_29460,N_28307);
nand UO_1186 (O_1186,N_25560,N_29703);
or UO_1187 (O_1187,N_28886,N_27946);
or UO_1188 (O_1188,N_27786,N_29475);
xor UO_1189 (O_1189,N_29032,N_27930);
or UO_1190 (O_1190,N_25614,N_28697);
and UO_1191 (O_1191,N_26071,N_25481);
nand UO_1192 (O_1192,N_25760,N_25049);
nor UO_1193 (O_1193,N_28927,N_27342);
nor UO_1194 (O_1194,N_27187,N_28816);
xor UO_1195 (O_1195,N_25275,N_25396);
or UO_1196 (O_1196,N_27832,N_29018);
xor UO_1197 (O_1197,N_27789,N_28736);
nor UO_1198 (O_1198,N_28878,N_26673);
nor UO_1199 (O_1199,N_26966,N_27670);
or UO_1200 (O_1200,N_26595,N_26326);
nor UO_1201 (O_1201,N_25217,N_25123);
nand UO_1202 (O_1202,N_25702,N_27920);
nor UO_1203 (O_1203,N_27344,N_29619);
nand UO_1204 (O_1204,N_28922,N_28704);
or UO_1205 (O_1205,N_26131,N_26765);
nor UO_1206 (O_1206,N_25448,N_29872);
or UO_1207 (O_1207,N_26286,N_29816);
nand UO_1208 (O_1208,N_25224,N_29201);
xnor UO_1209 (O_1209,N_26147,N_26271);
and UO_1210 (O_1210,N_25864,N_25301);
or UO_1211 (O_1211,N_29715,N_26343);
xor UO_1212 (O_1212,N_28039,N_25349);
nor UO_1213 (O_1213,N_25548,N_27112);
xor UO_1214 (O_1214,N_25949,N_25163);
nand UO_1215 (O_1215,N_27124,N_25480);
xnor UO_1216 (O_1216,N_29120,N_27802);
nand UO_1217 (O_1217,N_25862,N_28996);
nor UO_1218 (O_1218,N_29147,N_26411);
and UO_1219 (O_1219,N_25290,N_25740);
and UO_1220 (O_1220,N_29614,N_25566);
nand UO_1221 (O_1221,N_26750,N_27470);
or UO_1222 (O_1222,N_27907,N_29798);
or UO_1223 (O_1223,N_28179,N_29717);
xnor UO_1224 (O_1224,N_29412,N_26060);
or UO_1225 (O_1225,N_26425,N_26931);
xnor UO_1226 (O_1226,N_25551,N_29268);
and UO_1227 (O_1227,N_28836,N_28278);
nand UO_1228 (O_1228,N_29203,N_29227);
and UO_1229 (O_1229,N_25790,N_25001);
or UO_1230 (O_1230,N_26207,N_26640);
and UO_1231 (O_1231,N_28633,N_27275);
and UO_1232 (O_1232,N_26937,N_28948);
nand UO_1233 (O_1233,N_26887,N_25355);
nor UO_1234 (O_1234,N_28645,N_25561);
and UO_1235 (O_1235,N_28851,N_29579);
and UO_1236 (O_1236,N_27857,N_25404);
or UO_1237 (O_1237,N_26547,N_29182);
nor UO_1238 (O_1238,N_29096,N_27401);
xnor UO_1239 (O_1239,N_28578,N_25054);
nor UO_1240 (O_1240,N_28170,N_27210);
xnor UO_1241 (O_1241,N_26275,N_27955);
nand UO_1242 (O_1242,N_28644,N_27033);
nor UO_1243 (O_1243,N_25183,N_26725);
nor UO_1244 (O_1244,N_27359,N_28423);
xor UO_1245 (O_1245,N_27570,N_28177);
nand UO_1246 (O_1246,N_25570,N_25979);
and UO_1247 (O_1247,N_26995,N_28020);
or UO_1248 (O_1248,N_26366,N_26926);
nor UO_1249 (O_1249,N_26661,N_28305);
xor UO_1250 (O_1250,N_25153,N_26703);
nor UO_1251 (O_1251,N_28669,N_27456);
xor UO_1252 (O_1252,N_28655,N_28639);
xor UO_1253 (O_1253,N_25935,N_26838);
nor UO_1254 (O_1254,N_27364,N_29596);
xor UO_1255 (O_1255,N_27661,N_29510);
nand UO_1256 (O_1256,N_25201,N_27606);
and UO_1257 (O_1257,N_25653,N_27712);
or UO_1258 (O_1258,N_26161,N_25345);
xnor UO_1259 (O_1259,N_25594,N_25029);
nand UO_1260 (O_1260,N_29308,N_28150);
or UO_1261 (O_1261,N_27457,N_29185);
xnor UO_1262 (O_1262,N_25543,N_26337);
and UO_1263 (O_1263,N_26585,N_27159);
and UO_1264 (O_1264,N_29473,N_29864);
and UO_1265 (O_1265,N_25242,N_27041);
xor UO_1266 (O_1266,N_26405,N_25520);
xor UO_1267 (O_1267,N_26100,N_26708);
nor UO_1268 (O_1268,N_28165,N_25173);
nor UO_1269 (O_1269,N_28356,N_25317);
nand UO_1270 (O_1270,N_29856,N_28445);
and UO_1271 (O_1271,N_29949,N_25938);
xnor UO_1272 (O_1272,N_26655,N_29834);
and UO_1273 (O_1273,N_27294,N_28815);
nand UO_1274 (O_1274,N_25066,N_29384);
and UO_1275 (O_1275,N_26281,N_28424);
nor UO_1276 (O_1276,N_28849,N_27718);
and UO_1277 (O_1277,N_26826,N_25120);
nor UO_1278 (O_1278,N_29481,N_25521);
nand UO_1279 (O_1279,N_27477,N_29582);
or UO_1280 (O_1280,N_27722,N_25065);
nand UO_1281 (O_1281,N_29721,N_26369);
nand UO_1282 (O_1282,N_29768,N_28009);
nor UO_1283 (O_1283,N_26121,N_27415);
or UO_1284 (O_1284,N_29810,N_25699);
xor UO_1285 (O_1285,N_29529,N_29061);
nand UO_1286 (O_1286,N_25361,N_28526);
nor UO_1287 (O_1287,N_29876,N_28201);
xor UO_1288 (O_1288,N_25499,N_29063);
or UO_1289 (O_1289,N_27051,N_29341);
nand UO_1290 (O_1290,N_26212,N_29792);
nand UO_1291 (O_1291,N_28675,N_29542);
nand UO_1292 (O_1292,N_27069,N_26688);
or UO_1293 (O_1293,N_28620,N_27833);
xor UO_1294 (O_1294,N_26895,N_25767);
nor UO_1295 (O_1295,N_29705,N_26020);
xor UO_1296 (O_1296,N_29854,N_27099);
or UO_1297 (O_1297,N_29969,N_28022);
xnor UO_1298 (O_1298,N_27438,N_26444);
or UO_1299 (O_1299,N_25883,N_25429);
or UO_1300 (O_1300,N_26300,N_27302);
and UO_1301 (O_1301,N_26901,N_26896);
nor UO_1302 (O_1302,N_29592,N_25819);
xor UO_1303 (O_1303,N_27061,N_25095);
nand UO_1304 (O_1304,N_28245,N_29646);
xnor UO_1305 (O_1305,N_26079,N_26048);
nor UO_1306 (O_1306,N_26023,N_29405);
xnor UO_1307 (O_1307,N_29068,N_26866);
nand UO_1308 (O_1308,N_28363,N_25454);
nor UO_1309 (O_1309,N_26675,N_28742);
and UO_1310 (O_1310,N_28687,N_26335);
nand UO_1311 (O_1311,N_26432,N_26113);
nor UO_1312 (O_1312,N_29905,N_27098);
xnor UO_1313 (O_1313,N_28584,N_28087);
or UO_1314 (O_1314,N_27161,N_29855);
or UO_1315 (O_1315,N_27985,N_25532);
or UO_1316 (O_1316,N_26044,N_25223);
xor UO_1317 (O_1317,N_25284,N_26112);
or UO_1318 (O_1318,N_27814,N_26150);
xnor UO_1319 (O_1319,N_28489,N_28223);
or UO_1320 (O_1320,N_27923,N_29108);
xnor UO_1321 (O_1321,N_27491,N_29637);
xor UO_1322 (O_1322,N_26457,N_27775);
and UO_1323 (O_1323,N_28660,N_26467);
nand UO_1324 (O_1324,N_25314,N_29640);
and UO_1325 (O_1325,N_26768,N_27649);
and UO_1326 (O_1326,N_26538,N_25621);
xor UO_1327 (O_1327,N_28834,N_26759);
xor UO_1328 (O_1328,N_28869,N_26602);
xor UO_1329 (O_1329,N_26186,N_28100);
or UO_1330 (O_1330,N_29048,N_29407);
xnor UO_1331 (O_1331,N_26637,N_25139);
and UO_1332 (O_1332,N_27511,N_25987);
nand UO_1333 (O_1333,N_29176,N_26639);
xnor UO_1334 (O_1334,N_28394,N_28364);
xor UO_1335 (O_1335,N_28404,N_25593);
nor UO_1336 (O_1336,N_25383,N_29051);
nor UO_1337 (O_1337,N_28859,N_25829);
and UO_1338 (O_1338,N_27168,N_25238);
and UO_1339 (O_1339,N_27766,N_28967);
or UO_1340 (O_1340,N_27628,N_27220);
nor UO_1341 (O_1341,N_28981,N_29711);
nor UO_1342 (O_1342,N_26529,N_26062);
nor UO_1343 (O_1343,N_29575,N_27278);
nor UO_1344 (O_1344,N_25536,N_27453);
or UO_1345 (O_1345,N_25978,N_27445);
nor UO_1346 (O_1346,N_27118,N_29371);
or UO_1347 (O_1347,N_27245,N_26518);
nor UO_1348 (O_1348,N_27873,N_28913);
xor UO_1349 (O_1349,N_25180,N_28844);
nand UO_1350 (O_1350,N_27227,N_27319);
or UO_1351 (O_1351,N_25205,N_28006);
nor UO_1352 (O_1352,N_27070,N_29505);
nor UO_1353 (O_1353,N_25376,N_25336);
and UO_1354 (O_1354,N_28141,N_27497);
xnor UO_1355 (O_1355,N_29213,N_28484);
nor UO_1356 (O_1356,N_25749,N_29631);
xor UO_1357 (O_1357,N_29965,N_25402);
nor UO_1358 (O_1358,N_26878,N_26486);
nor UO_1359 (O_1359,N_27508,N_26604);
and UO_1360 (O_1360,N_27557,N_29747);
nand UO_1361 (O_1361,N_29320,N_29546);
and UO_1362 (O_1362,N_27803,N_28929);
and UO_1363 (O_1363,N_28989,N_26277);
nor UO_1364 (O_1364,N_27138,N_26551);
xnor UO_1365 (O_1365,N_25679,N_29888);
or UO_1366 (O_1366,N_26503,N_25753);
nor UO_1367 (O_1367,N_27705,N_27128);
or UO_1368 (O_1368,N_25195,N_26409);
nor UO_1369 (O_1369,N_29422,N_28342);
or UO_1370 (O_1370,N_26519,N_25933);
nor UO_1371 (O_1371,N_25353,N_27890);
nor UO_1372 (O_1372,N_29137,N_25528);
nand UO_1373 (O_1373,N_26246,N_25824);
xor UO_1374 (O_1374,N_28314,N_28730);
xnor UO_1375 (O_1375,N_29676,N_25472);
nand UO_1376 (O_1376,N_29356,N_27182);
or UO_1377 (O_1377,N_28565,N_26925);
and UO_1378 (O_1378,N_28903,N_29312);
nor UO_1379 (O_1379,N_26330,N_26600);
nor UO_1380 (O_1380,N_27451,N_28539);
xor UO_1381 (O_1381,N_25652,N_27270);
nor UO_1382 (O_1382,N_25395,N_25130);
nor UO_1383 (O_1383,N_27082,N_25981);
and UO_1384 (O_1384,N_25649,N_29199);
or UO_1385 (O_1385,N_28162,N_26744);
or UO_1386 (O_1386,N_28139,N_29131);
nand UO_1387 (O_1387,N_26397,N_28642);
xnor UO_1388 (O_1388,N_28874,N_25114);
nand UO_1389 (O_1389,N_27079,N_25871);
and UO_1390 (O_1390,N_27769,N_28495);
xor UO_1391 (O_1391,N_27006,N_26016);
or UO_1392 (O_1392,N_25794,N_26819);
and UO_1393 (O_1393,N_29960,N_25972);
nand UO_1394 (O_1394,N_25803,N_25603);
nand UO_1395 (O_1395,N_28611,N_28864);
nand UO_1396 (O_1396,N_27970,N_26761);
or UO_1397 (O_1397,N_25896,N_28766);
and UO_1398 (O_1398,N_25303,N_29799);
nand UO_1399 (O_1399,N_29932,N_25249);
xnor UO_1400 (O_1400,N_25083,N_29262);
or UO_1401 (O_1401,N_26287,N_26193);
and UO_1402 (O_1402,N_27440,N_25308);
nor UO_1403 (O_1403,N_25146,N_26148);
and UO_1404 (O_1404,N_28336,N_29304);
or UO_1405 (O_1405,N_26704,N_26561);
and UO_1406 (O_1406,N_27485,N_25546);
and UO_1407 (O_1407,N_29261,N_28590);
nand UO_1408 (O_1408,N_28895,N_25805);
and UO_1409 (O_1409,N_29593,N_28386);
xor UO_1410 (O_1410,N_25797,N_27982);
or UO_1411 (O_1411,N_28248,N_27377);
and UO_1412 (O_1412,N_29134,N_25432);
nor UO_1413 (O_1413,N_27835,N_27064);
xnor UO_1414 (O_1414,N_29290,N_28867);
xnor UO_1415 (O_1415,N_28031,N_29221);
xnor UO_1416 (O_1416,N_27709,N_25443);
and UO_1417 (O_1417,N_29558,N_27398);
or UO_1418 (O_1418,N_25633,N_26257);
and UO_1419 (O_1419,N_27881,N_25571);
nor UO_1420 (O_1420,N_28304,N_25882);
xnor UO_1421 (O_1421,N_25216,N_26459);
nand UO_1422 (O_1422,N_26549,N_25634);
and UO_1423 (O_1423,N_29933,N_29911);
or UO_1424 (O_1424,N_28058,N_25283);
or UO_1425 (O_1425,N_28779,N_25830);
or UO_1426 (O_1426,N_29591,N_28281);
and UO_1427 (O_1427,N_29167,N_26216);
or UO_1428 (O_1428,N_25585,N_27629);
or UO_1429 (O_1429,N_28936,N_29685);
or UO_1430 (O_1430,N_25497,N_27009);
or UO_1431 (O_1431,N_29735,N_25413);
or UO_1432 (O_1432,N_26957,N_29190);
nand UO_1433 (O_1433,N_29781,N_27363);
or UO_1434 (O_1434,N_25126,N_25199);
and UO_1435 (O_1435,N_27683,N_25280);
nor UO_1436 (O_1436,N_27494,N_28557);
xnor UO_1437 (O_1437,N_26918,N_25338);
nor UO_1438 (O_1438,N_25168,N_29899);
and UO_1439 (O_1439,N_26927,N_25403);
nand UO_1440 (O_1440,N_27837,N_28054);
or UO_1441 (O_1441,N_29253,N_29124);
and UO_1442 (O_1442,N_26855,N_28519);
or UO_1443 (O_1443,N_28535,N_25148);
xnor UO_1444 (O_1444,N_25022,N_27630);
nor UO_1445 (O_1445,N_26492,N_25064);
xor UO_1446 (O_1446,N_26528,N_25221);
or UO_1447 (O_1447,N_28473,N_26285);
nor UO_1448 (O_1448,N_29339,N_28705);
or UO_1449 (O_1449,N_27576,N_25455);
and UO_1450 (O_1450,N_26619,N_29025);
nor UO_1451 (O_1451,N_26428,N_27808);
nor UO_1452 (O_1452,N_29532,N_26198);
nand UO_1453 (O_1453,N_28592,N_25732);
nor UO_1454 (O_1454,N_26160,N_25136);
xor UO_1455 (O_1455,N_29674,N_29454);
and UO_1456 (O_1456,N_27013,N_27736);
nor UO_1457 (O_1457,N_28130,N_27518);
nor UO_1458 (O_1458,N_28931,N_27546);
nor UO_1459 (O_1459,N_29830,N_25474);
and UO_1460 (O_1460,N_27539,N_25370);
or UO_1461 (O_1461,N_27579,N_25268);
or UO_1462 (O_1462,N_27655,N_29279);
xnor UO_1463 (O_1463,N_29216,N_27154);
and UO_1464 (O_1464,N_28845,N_28037);
xor UO_1465 (O_1465,N_28446,N_29186);
and UO_1466 (O_1466,N_28042,N_27431);
and UO_1467 (O_1467,N_29163,N_25422);
nand UO_1468 (O_1468,N_25996,N_29326);
or UO_1469 (O_1469,N_27408,N_27375);
nor UO_1470 (O_1470,N_25156,N_28199);
and UO_1471 (O_1471,N_27414,N_26798);
xnor UO_1472 (O_1472,N_29101,N_27337);
xnor UO_1473 (O_1473,N_27801,N_27699);
nand UO_1474 (O_1474,N_27345,N_29205);
and UO_1475 (O_1475,N_25182,N_28447);
nand UO_1476 (O_1476,N_26283,N_25870);
nor UO_1477 (O_1477,N_28349,N_25983);
nand UO_1478 (O_1478,N_27989,N_26954);
or UO_1479 (O_1479,N_28119,N_26328);
and UO_1480 (O_1480,N_25863,N_26163);
nand UO_1481 (O_1481,N_29008,N_29683);
or UO_1482 (O_1482,N_26806,N_25815);
or UO_1483 (O_1483,N_25380,N_27642);
nand UO_1484 (O_1484,N_28838,N_25866);
and UO_1485 (O_1485,N_28857,N_25849);
or UO_1486 (O_1486,N_29813,N_27754);
nor UO_1487 (O_1487,N_25535,N_27645);
nand UO_1488 (O_1488,N_26784,N_29630);
xnor UO_1489 (O_1489,N_28280,N_26471);
and UO_1490 (O_1490,N_29656,N_25823);
or UO_1491 (O_1491,N_27751,N_25202);
or UO_1492 (O_1492,N_27862,N_28415);
or UO_1493 (O_1493,N_29881,N_29148);
or UO_1494 (O_1494,N_29980,N_26338);
nor UO_1495 (O_1495,N_26922,N_25074);
nand UO_1496 (O_1496,N_29072,N_25346);
nand UO_1497 (O_1497,N_25204,N_29764);
xor UO_1498 (O_1498,N_25412,N_27176);
nand UO_1499 (O_1499,N_27542,N_25519);
nand UO_1500 (O_1500,N_26622,N_27571);
and UO_1501 (O_1501,N_29425,N_26488);
nor UO_1502 (O_1502,N_29645,N_28457);
and UO_1503 (O_1503,N_25586,N_28573);
or UO_1504 (O_1504,N_25625,N_25386);
nor UO_1505 (O_1505,N_26436,N_26705);
nand UO_1506 (O_1506,N_26775,N_25640);
and UO_1507 (O_1507,N_29458,N_29014);
nor UO_1508 (O_1508,N_27902,N_28694);
or UO_1509 (O_1509,N_29954,N_27828);
nor UO_1510 (O_1510,N_28944,N_25239);
xor UO_1511 (O_1511,N_26209,N_25620);
or UO_1512 (O_1512,N_28881,N_26647);
xnor UO_1513 (O_1513,N_29479,N_29995);
or UO_1514 (O_1514,N_28807,N_27437);
nor UO_1515 (O_1515,N_27145,N_29859);
nand UO_1516 (O_1516,N_29433,N_29075);
nor UO_1517 (O_1517,N_29432,N_29568);
and UO_1518 (O_1518,N_26440,N_29077);
xor UO_1519 (O_1519,N_25194,N_25694);
or UO_1520 (O_1520,N_27236,N_26410);
nand UO_1521 (O_1521,N_27233,N_27714);
nor UO_1522 (O_1522,N_25992,N_28417);
nand UO_1523 (O_1523,N_29846,N_29912);
or UO_1524 (O_1524,N_27056,N_25616);
nand UO_1525 (O_1525,N_27416,N_26124);
nand UO_1526 (O_1526,N_27419,N_26633);
xor UO_1527 (O_1527,N_27269,N_26278);
nor UO_1528 (O_1528,N_25486,N_25626);
nor UO_1529 (O_1529,N_25534,N_26752);
and UO_1530 (O_1530,N_25208,N_25176);
xor UO_1531 (O_1531,N_26565,N_29006);
or UO_1532 (O_1532,N_29233,N_26920);
or UO_1533 (O_1533,N_25203,N_28299);
nor UO_1534 (O_1534,N_27177,N_26645);
or UO_1535 (O_1535,N_29311,N_28403);
and UO_1536 (O_1536,N_28122,N_27493);
nand UO_1537 (O_1537,N_26740,N_28711);
and UO_1538 (O_1538,N_29374,N_27782);
nand UO_1539 (O_1539,N_26180,N_25761);
nor UO_1540 (O_1540,N_27659,N_25912);
nand UO_1541 (O_1541,N_29939,N_29693);
or UO_1542 (O_1542,N_28345,N_25483);
or UO_1543 (O_1543,N_27615,N_27165);
xor UO_1544 (O_1544,N_26011,N_25752);
nand UO_1545 (O_1545,N_28357,N_25243);
or UO_1546 (O_1546,N_27448,N_26888);
nor UO_1547 (O_1547,N_25236,N_29971);
xnor UO_1548 (O_1548,N_29097,N_29726);
nand UO_1549 (O_1549,N_28901,N_29889);
or UO_1550 (O_1550,N_25669,N_27290);
nor UO_1551 (O_1551,N_27585,N_25399);
and UO_1552 (O_1552,N_27635,N_26982);
nor UO_1553 (O_1553,N_29951,N_26903);
nand UO_1554 (O_1554,N_29554,N_29200);
or UO_1555 (O_1555,N_27109,N_25140);
and UO_1556 (O_1556,N_29643,N_28190);
nand UO_1557 (O_1557,N_27931,N_28072);
nor UO_1558 (O_1558,N_29447,N_25954);
nand UO_1559 (O_1559,N_26679,N_26694);
or UO_1560 (O_1560,N_28634,N_29821);
xnor UO_1561 (O_1561,N_28453,N_25720);
xor UO_1562 (O_1562,N_26862,N_28581);
xor UO_1563 (O_1563,N_26696,N_26229);
and UO_1564 (O_1564,N_27194,N_25117);
nand UO_1565 (O_1565,N_25043,N_28377);
nor UO_1566 (O_1566,N_25456,N_25563);
and UO_1567 (O_1567,N_27387,N_26963);
or UO_1568 (O_1568,N_26423,N_29058);
nand UO_1569 (O_1569,N_27024,N_29100);
and UO_1570 (O_1570,N_27823,N_28828);
and UO_1571 (O_1571,N_25196,N_29106);
or UO_1572 (O_1572,N_29347,N_26724);
nor UO_1573 (O_1573,N_27043,N_25494);
nor UO_1574 (O_1574,N_26008,N_28494);
or UO_1575 (O_1575,N_29838,N_26911);
nor UO_1576 (O_1576,N_26105,N_25406);
xnor UO_1577 (O_1577,N_29325,N_26676);
nor UO_1578 (O_1578,N_29651,N_26218);
nor UO_1579 (O_1579,N_29191,N_25515);
or UO_1580 (O_1580,N_29482,N_28005);
or UO_1581 (O_1581,N_27421,N_29236);
nand UO_1582 (O_1582,N_25922,N_28950);
nand UO_1583 (O_1583,N_29511,N_26593);
and UO_1584 (O_1584,N_27697,N_27932);
and UO_1585 (O_1585,N_25921,N_25024);
or UO_1586 (O_1586,N_27904,N_29537);
xnor UO_1587 (O_1587,N_27382,N_29594);
or UO_1588 (O_1588,N_27088,N_27746);
or UO_1589 (O_1589,N_27114,N_26581);
and UO_1590 (O_1590,N_29580,N_26599);
xor UO_1591 (O_1591,N_27773,N_27228);
and UO_1592 (O_1592,N_29753,N_26621);
nand UO_1593 (O_1593,N_28949,N_26350);
nand UO_1594 (O_1594,N_27458,N_28093);
and UO_1595 (O_1595,N_29520,N_26061);
or UO_1596 (O_1596,N_26849,N_25611);
xnor UO_1597 (O_1597,N_26623,N_27582);
or UO_1598 (O_1598,N_26548,N_29102);
nand UO_1599 (O_1599,N_28142,N_29512);
nor UO_1600 (O_1600,N_29583,N_29386);
xor UO_1601 (O_1601,N_25320,N_25858);
xor UO_1602 (O_1602,N_27156,N_27003);
and UO_1603 (O_1603,N_25250,N_26907);
and UO_1604 (O_1604,N_27330,N_27326);
and UO_1605 (O_1605,N_25032,N_29171);
and UO_1606 (O_1606,N_26463,N_26357);
nand UO_1607 (O_1607,N_28389,N_28959);
nand UO_1608 (O_1608,N_25581,N_27317);
xnor UO_1609 (O_1609,N_29566,N_27981);
nand UO_1610 (O_1610,N_27022,N_26389);
nand UO_1611 (O_1611,N_27225,N_28737);
nand UO_1612 (O_1612,N_28206,N_26695);
nand UO_1613 (O_1613,N_27619,N_28765);
or UO_1614 (O_1614,N_27204,N_26331);
nor UO_1615 (O_1615,N_29401,N_26836);
or UO_1616 (O_1616,N_26065,N_26135);
xor UO_1617 (O_1617,N_27743,N_26108);
xnor UO_1618 (O_1618,N_28469,N_29423);
xnor UO_1619 (O_1619,N_29234,N_29688);
nor UO_1620 (O_1620,N_29360,N_29925);
and UO_1621 (O_1621,N_26127,N_26881);
nand UO_1622 (O_1622,N_27505,N_29483);
nand UO_1623 (O_1623,N_28574,N_25388);
and UO_1624 (O_1624,N_25750,N_27058);
xnor UO_1625 (O_1625,N_26371,N_25309);
and UO_1626 (O_1626,N_25274,N_27977);
nand UO_1627 (O_1627,N_27463,N_27871);
nor UO_1628 (O_1628,N_29224,N_28756);
xor UO_1629 (O_1629,N_27791,N_28120);
nand UO_1630 (O_1630,N_26003,N_26274);
and UO_1631 (O_1631,N_25511,N_29453);
or UO_1632 (O_1632,N_29795,N_28538);
nor UO_1633 (O_1633,N_29243,N_28272);
nand UO_1634 (O_1634,N_28518,N_27075);
or UO_1635 (O_1635,N_26889,N_27166);
or UO_1636 (O_1636,N_25220,N_27181);
and UO_1637 (O_1637,N_26955,N_26475);
nor UO_1638 (O_1638,N_26662,N_27356);
xnor UO_1639 (O_1639,N_28921,N_26427);
xnor UO_1640 (O_1640,N_28341,N_25789);
nor UO_1641 (O_1641,N_27287,N_29192);
xor UO_1642 (O_1642,N_27583,N_29974);
nand UO_1643 (O_1643,N_29609,N_27447);
nor UO_1644 (O_1644,N_29069,N_28560);
or UO_1645 (O_1645,N_27307,N_28575);
nand UO_1646 (O_1646,N_28123,N_28344);
or UO_1647 (O_1647,N_25484,N_29842);
and UO_1648 (O_1648,N_29195,N_27848);
xor UO_1649 (O_1649,N_28776,N_28214);
xnor UO_1650 (O_1650,N_28353,N_25505);
or UO_1651 (O_1651,N_29155,N_26217);
and UO_1652 (O_1652,N_28312,N_29265);
and UO_1653 (O_1653,N_29850,N_25476);
nand UO_1654 (O_1654,N_29410,N_25288);
and UO_1655 (O_1655,N_28580,N_25807);
and UO_1656 (O_1656,N_26191,N_28089);
xnor UO_1657 (O_1657,N_25259,N_25218);
or UO_1658 (O_1658,N_26839,N_29230);
xnor UO_1659 (O_1659,N_27912,N_27778);
nor UO_1660 (O_1660,N_28588,N_26136);
xor UO_1661 (O_1661,N_25919,N_25435);
and UO_1662 (O_1662,N_26171,N_29495);
xnor UO_1663 (O_1663,N_25989,N_29769);
nand UO_1664 (O_1664,N_28985,N_25756);
nand UO_1665 (O_1665,N_25742,N_25315);
or UO_1666 (O_1666,N_29943,N_28910);
nand UO_1667 (O_1667,N_26000,N_27618);
nand UO_1668 (O_1668,N_28595,N_28582);
and UO_1669 (O_1669,N_28583,N_26479);
nand UO_1670 (O_1670,N_27284,N_25031);
or UO_1671 (O_1671,N_25629,N_27947);
xor UO_1672 (O_1672,N_28499,N_28360);
xor UO_1673 (O_1673,N_25366,N_25041);
nor UO_1674 (O_1674,N_25468,N_28571);
or UO_1675 (O_1675,N_29151,N_27974);
or UO_1676 (O_1676,N_28906,N_27952);
and UO_1677 (O_1677,N_28081,N_26059);
xnor UO_1678 (O_1678,N_25814,N_28932);
nor UO_1679 (O_1679,N_28640,N_25906);
or UO_1680 (O_1680,N_29345,N_25197);
xor UO_1681 (O_1681,N_25193,N_26680);
xnor UO_1682 (O_1682,N_26877,N_28656);
xnor UO_1683 (O_1683,N_29739,N_25010);
nand UO_1684 (O_1684,N_29400,N_29761);
or UO_1685 (O_1685,N_27206,N_28636);
nor UO_1686 (O_1686,N_28439,N_28270);
or UO_1687 (O_1687,N_28946,N_28662);
nand UO_1688 (O_1688,N_27362,N_28425);
nor UO_1689 (O_1689,N_27687,N_28253);
xnor UO_1690 (O_1690,N_25246,N_29903);
nor UO_1691 (O_1691,N_25270,N_28293);
nor UO_1692 (O_1692,N_28065,N_25943);
or UO_1693 (O_1693,N_29687,N_29938);
nand UO_1694 (O_1694,N_28729,N_26258);
nor UO_1695 (O_1695,N_28979,N_25415);
nor UO_1696 (O_1696,N_26913,N_29297);
and UO_1697 (O_1697,N_27328,N_29298);
xor UO_1698 (O_1698,N_27148,N_26530);
and UO_1699 (O_1699,N_29039,N_27900);
nor UO_1700 (O_1700,N_28882,N_25094);
nand UO_1701 (O_1701,N_27829,N_29045);
and UO_1702 (O_1702,N_28688,N_29744);
nor UO_1703 (O_1703,N_27879,N_27788);
nor UO_1704 (O_1704,N_28522,N_27370);
or UO_1705 (O_1705,N_29862,N_25219);
nand UO_1706 (O_1706,N_29973,N_27841);
or UO_1707 (O_1707,N_26747,N_28482);
and UO_1708 (O_1708,N_29420,N_27779);
or UO_1709 (O_1709,N_28939,N_25999);
nand UO_1710 (O_1710,N_29079,N_26700);
or UO_1711 (O_1711,N_25731,N_26580);
xnor UO_1712 (O_1712,N_29589,N_26390);
and UO_1713 (O_1713,N_26238,N_29567);
nand UO_1714 (O_1714,N_28085,N_25488);
nand UO_1715 (O_1715,N_28373,N_28911);
and UO_1716 (O_1716,N_28965,N_25914);
nor UO_1717 (O_1717,N_25107,N_26232);
or UO_1718 (O_1718,N_27971,N_29349);
or UO_1719 (O_1719,N_27719,N_29986);
and UO_1720 (O_1720,N_25963,N_29672);
xor UO_1721 (O_1721,N_25717,N_25281);
nand UO_1722 (O_1722,N_26670,N_27369);
or UO_1723 (O_1723,N_29573,N_25700);
or UO_1724 (O_1724,N_27798,N_26015);
xnor UO_1725 (O_1725,N_28441,N_28244);
or UO_1726 (O_1726,N_26531,N_29922);
nor UO_1727 (O_1727,N_29098,N_28337);
nand UO_1728 (O_1728,N_29352,N_26320);
nand UO_1729 (O_1729,N_25485,N_26996);
nand UO_1730 (O_1730,N_25656,N_29457);
nand UO_1731 (O_1731,N_26570,N_28607);
nor UO_1732 (O_1732,N_29959,N_28354);
xor UO_1733 (O_1733,N_27653,N_26247);
nand UO_1734 (O_1734,N_29465,N_27224);
xnor UO_1735 (O_1735,N_29126,N_29122);
or UO_1736 (O_1736,N_29869,N_28033);
nor UO_1737 (O_1737,N_27455,N_29258);
or UO_1738 (O_1738,N_26789,N_28397);
or UO_1739 (O_1739,N_27739,N_28046);
nand UO_1740 (O_1740,N_27333,N_28187);
nor UO_1741 (O_1741,N_27057,N_25105);
nand UO_1742 (O_1742,N_25516,N_29836);
xor UO_1743 (O_1743,N_25766,N_26451);
and UO_1744 (O_1744,N_27492,N_28714);
xnor UO_1745 (O_1745,N_29828,N_26017);
nand UO_1746 (O_1746,N_29858,N_26586);
and UO_1747 (O_1747,N_26832,N_29353);
nor UO_1748 (O_1748,N_27554,N_28071);
and UO_1749 (O_1749,N_27678,N_27336);
xor UO_1750 (O_1750,N_29749,N_28183);
xor UO_1751 (O_1751,N_28266,N_27733);
xnor UO_1752 (O_1752,N_28891,N_25263);
nand UO_1753 (O_1753,N_28786,N_28693);
xor UO_1754 (O_1754,N_29849,N_28799);
and UO_1755 (O_1755,N_26556,N_28306);
nor UO_1756 (O_1756,N_25956,N_29633);
nor UO_1757 (O_1757,N_25398,N_27016);
and UO_1758 (O_1758,N_27758,N_29906);
and UO_1759 (O_1759,N_27616,N_28014);
and UO_1760 (O_1760,N_26884,N_27080);
and UO_1761 (O_1761,N_29584,N_28548);
nor UO_1762 (O_1762,N_25278,N_26994);
and UO_1763 (O_1763,N_26975,N_28673);
nor UO_1764 (O_1764,N_25033,N_25419);
and UO_1765 (O_1765,N_28221,N_28061);
xor UO_1766 (O_1766,N_25452,N_28942);
and UO_1767 (O_1767,N_25602,N_27396);
nor UO_1768 (O_1768,N_25860,N_25300);
nand UO_1769 (O_1769,N_29024,N_25371);
and UO_1770 (O_1770,N_28553,N_27240);
or UO_1771 (O_1771,N_29678,N_25391);
xor UO_1772 (O_1772,N_27380,N_25776);
xnor UO_1773 (O_1773,N_27877,N_29250);
nor UO_1774 (O_1774,N_28853,N_27767);
xnor UO_1775 (O_1775,N_28811,N_25261);
or UO_1776 (O_1776,N_28817,N_27852);
and UO_1777 (O_1777,N_29435,N_28078);
and UO_1778 (O_1778,N_25680,N_25099);
and UO_1779 (O_1779,N_29843,N_28329);
nor UO_1780 (O_1780,N_28203,N_28803);
nand UO_1781 (O_1781,N_26392,N_27617);
and UO_1782 (O_1782,N_25971,N_29714);
xor UO_1783 (O_1783,N_27658,N_28274);
xnor UO_1784 (O_1784,N_25011,N_26170);
and UO_1785 (O_1785,N_29187,N_29037);
xor UO_1786 (O_1786,N_27155,N_27990);
nand UO_1787 (O_1787,N_26649,N_26672);
nand UO_1788 (O_1788,N_27665,N_25796);
nor UO_1789 (O_1789,N_29373,N_27014);
or UO_1790 (O_1790,N_29111,N_25665);
xnor UO_1791 (O_1791,N_29136,N_29322);
nand UO_1792 (O_1792,N_26514,N_25836);
and UO_1793 (O_1793,N_27748,N_26823);
nor UO_1794 (O_1794,N_29729,N_29146);
xnor UO_1795 (O_1795,N_29504,N_27637);
nor UO_1796 (O_1796,N_28106,N_25693);
nor UO_1797 (O_1797,N_25327,N_29089);
xor UO_1798 (O_1798,N_27049,N_27474);
or UO_1799 (O_1799,N_25675,N_26089);
or UO_1800 (O_1800,N_27589,N_28654);
nor UO_1801 (O_1801,N_28900,N_26616);
nor UO_1802 (O_1802,N_29231,N_26634);
xor UO_1803 (O_1803,N_26651,N_25613);
nand UO_1804 (O_1804,N_28428,N_29464);
and UO_1805 (O_1805,N_29924,N_25492);
xnor UO_1806 (O_1806,N_27896,N_28067);
nand UO_1807 (O_1807,N_27750,N_28925);
xor UO_1808 (O_1808,N_29967,N_25061);
xnor UO_1809 (O_1809,N_29884,N_25127);
nor UO_1810 (O_1810,N_25230,N_28629);
xor UO_1811 (O_1811,N_27221,N_27940);
nand UO_1812 (O_1812,N_27308,N_28987);
nor UO_1813 (O_1813,N_25961,N_26713);
nand UO_1814 (O_1814,N_25048,N_27265);
xor UO_1815 (O_1815,N_27897,N_29978);
and UO_1816 (O_1816,N_28409,N_29092);
and UO_1817 (O_1817,N_28181,N_27110);
xnor UO_1818 (O_1818,N_29727,N_28823);
or UO_1819 (O_1819,N_28118,N_27928);
nor UO_1820 (O_1820,N_29734,N_28103);
or UO_1821 (O_1821,N_25319,N_26945);
and UO_1822 (O_1822,N_29154,N_25189);
xor UO_1823 (O_1823,N_28080,N_26507);
and UO_1824 (O_1824,N_27885,N_27339);
or UO_1825 (O_1825,N_28545,N_29494);
and UO_1826 (O_1826,N_27915,N_25539);
xnor UO_1827 (O_1827,N_29624,N_27381);
xor UO_1828 (O_1828,N_28200,N_25841);
nand UO_1829 (O_1829,N_29395,N_27716);
nor UO_1830 (O_1830,N_28084,N_29450);
and UO_1831 (O_1831,N_25307,N_28516);
or UO_1832 (O_1832,N_28554,N_26522);
xnor UO_1833 (O_1833,N_29046,N_29909);
nand UO_1834 (O_1834,N_28720,N_28798);
xnor UO_1835 (O_1835,N_27048,N_28983);
and UO_1836 (O_1836,N_28982,N_27469);
or UO_1837 (O_1837,N_28622,N_28243);
xnor UO_1838 (O_1838,N_29443,N_29477);
nor UO_1839 (O_1839,N_26967,N_27094);
nor UO_1840 (O_1840,N_28128,N_25960);
nor UO_1841 (O_1841,N_29365,N_27274);
nor UO_1842 (O_1842,N_25941,N_26620);
and UO_1843 (O_1843,N_29139,N_27151);
nand UO_1844 (O_1844,N_27969,N_26785);
nand UO_1845 (O_1845,N_27624,N_29337);
nand UO_1846 (O_1846,N_25142,N_29647);
or UO_1847 (O_1847,N_28724,N_28466);
or UO_1848 (O_1848,N_27600,N_28422);
nand UO_1849 (O_1849,N_26707,N_26856);
nand UO_1850 (O_1850,N_25296,N_29086);
or UO_1851 (O_1851,N_26560,N_28653);
nand UO_1852 (O_1852,N_27792,N_27046);
or UO_1853 (O_1853,N_26253,N_27936);
nor UO_1854 (O_1854,N_28216,N_26379);
nand UO_1855 (O_1855,N_25986,N_28787);
xnor UO_1856 (O_1856,N_27836,N_26364);
and UO_1857 (O_1857,N_25985,N_26953);
and UO_1858 (O_1858,N_26064,N_25890);
xor UO_1859 (O_1859,N_25222,N_27708);
or UO_1860 (O_1860,N_26324,N_25559);
nor UO_1861 (O_1861,N_26097,N_25198);
nor UO_1862 (O_1862,N_29950,N_27818);
or UO_1863 (O_1863,N_27741,N_29302);
xnor UO_1864 (O_1864,N_27197,N_28286);
or UO_1865 (O_1865,N_28789,N_25299);
nand UO_1866 (O_1866,N_29428,N_28726);
or UO_1867 (O_1867,N_27424,N_28650);
and UO_1868 (O_1868,N_25269,N_27170);
nand UO_1869 (O_1869,N_27706,N_27734);
or UO_1870 (O_1870,N_27834,N_26327);
or UO_1871 (O_1871,N_27870,N_28074);
or UO_1872 (O_1872,N_26311,N_25377);
xor UO_1873 (O_1873,N_28166,N_26026);
and UO_1874 (O_1874,N_25304,N_25787);
or UO_1875 (O_1875,N_25635,N_27038);
or UO_1876 (O_1876,N_28860,N_26793);
xor UO_1877 (O_1877,N_26516,N_26681);
nand UO_1878 (O_1878,N_25417,N_29009);
and UO_1879 (O_1879,N_27473,N_28159);
nand UO_1880 (O_1880,N_26394,N_28426);
or UO_1881 (O_1881,N_25746,N_28641);
nor UO_1882 (O_1882,N_26532,N_25384);
nor UO_1883 (O_1883,N_28879,N_29235);
or UO_1884 (O_1884,N_28383,N_26797);
nor UO_1885 (O_1885,N_27657,N_26987);
xor UO_1886 (O_1886,N_29351,N_28480);
nand UO_1887 (O_1887,N_25557,N_29945);
nand UO_1888 (O_1888,N_27312,N_26251);
nor UO_1889 (O_1889,N_28793,N_25512);
nor UO_1890 (O_1890,N_28366,N_28483);
nand UO_1891 (O_1891,N_26490,N_28156);
nor UO_1892 (O_1892,N_29809,N_26998);
and UO_1893 (O_1893,N_26199,N_27668);
nor UO_1894 (O_1894,N_25619,N_28362);
nand UO_1895 (O_1895,N_26446,N_29803);
nand UO_1896 (O_1896,N_26052,N_25690);
and UO_1897 (O_1897,N_28778,N_29066);
nand UO_1898 (O_1898,N_28806,N_28746);
nor UO_1899 (O_1899,N_28202,N_28805);
xor UO_1900 (O_1900,N_28664,N_25175);
and UO_1901 (O_1901,N_25905,N_28887);
nor UO_1902 (O_1902,N_27866,N_28594);
or UO_1903 (O_1903,N_25257,N_27551);
or UO_1904 (O_1904,N_28898,N_29662);
nor UO_1905 (O_1905,N_29010,N_26758);
nand UO_1906 (O_1906,N_29530,N_26417);
nor UO_1907 (O_1907,N_28016,N_28840);
or UO_1908 (O_1908,N_27311,N_28744);
or UO_1909 (O_1909,N_28097,N_26036);
or UO_1910 (O_1910,N_29206,N_29806);
and UO_1911 (O_1911,N_25210,N_26875);
and UO_1912 (O_1912,N_28029,N_28938);
nor UO_1913 (O_1913,N_27868,N_27815);
or UO_1914 (O_1914,N_29820,N_29251);
or UO_1915 (O_1915,N_27215,N_26554);
nand UO_1916 (O_1916,N_28648,N_28478);
and UO_1917 (O_1917,N_27121,N_26824);
nand UO_1918 (O_1918,N_28435,N_28868);
nand UO_1919 (O_1919,N_26505,N_26511);
nand UO_1920 (O_1920,N_29868,N_29183);
or UO_1921 (O_1921,N_25976,N_27223);
or UO_1922 (O_1922,N_29043,N_26156);
xnor UO_1923 (O_1923,N_29993,N_28257);
nand UO_1924 (O_1924,N_26796,N_28631);
nand UO_1925 (O_1925,N_25902,N_25234);
nor UO_1926 (O_1926,N_28758,N_28537);
and UO_1927 (O_1927,N_27682,N_25878);
or UO_1928 (O_1928,N_27503,N_27612);
nor UO_1929 (O_1929,N_26715,N_26709);
xnor UO_1930 (O_1930,N_28544,N_27467);
and UO_1931 (O_1931,N_28802,N_25711);
xor UO_1932 (O_1932,N_28521,N_25859);
and UO_1933 (O_1933,N_25897,N_27768);
nand UO_1934 (O_1934,N_26046,N_26988);
and UO_1935 (O_1935,N_25469,N_25658);
xnor UO_1936 (O_1936,N_27725,N_29670);
nor UO_1937 (O_1937,N_29355,N_25907);
or UO_1938 (O_1938,N_25735,N_28339);
xor UO_1939 (O_1939,N_28973,N_28225);
nand UO_1940 (O_1940,N_29336,N_25045);
or UO_1941 (O_1941,N_26582,N_26252);
or UO_1942 (O_1942,N_29559,N_28260);
xor UO_1943 (O_1943,N_29961,N_25143);
and UO_1944 (O_1944,N_28062,N_28791);
nor UO_1945 (O_1945,N_27468,N_28723);
nand UO_1946 (O_1946,N_26374,N_28116);
xnor UO_1947 (O_1947,N_27464,N_29548);
xnor UO_1948 (O_1948,N_25428,N_26145);
xor UO_1949 (O_1949,N_25869,N_27255);
and UO_1950 (O_1950,N_27327,N_26618);
xor UO_1951 (O_1951,N_27442,N_29301);
nand UO_1952 (O_1952,N_26254,N_29307);
or UO_1953 (O_1953,N_28951,N_28596);
and UO_1954 (O_1954,N_27510,N_28481);
nand UO_1955 (O_1955,N_26985,N_27886);
xnor UO_1956 (O_1956,N_29456,N_26084);
or UO_1957 (O_1957,N_27962,N_29228);
or UO_1958 (O_1958,N_26453,N_26720);
and UO_1959 (O_1959,N_29209,N_29127);
or UO_1960 (O_1960,N_25759,N_26916);
nand UO_1961 (O_1961,N_26825,N_28503);
and UO_1962 (O_1962,N_25748,N_26900);
nor UO_1963 (O_1963,N_25847,N_26176);
nand UO_1964 (O_1964,N_25668,N_29826);
or UO_1965 (O_1965,N_29915,N_26249);
or UO_1966 (O_1966,N_26149,N_29805);
xor UO_1967 (O_1967,N_25936,N_28406);
xnor UO_1968 (O_1968,N_28659,N_27350);
xor UO_1969 (O_1969,N_26893,N_27664);
or UO_1970 (O_1970,N_26776,N_26606);
nand UO_1971 (O_1971,N_25339,N_25692);
and UO_1972 (O_1972,N_25112,N_26635);
xnor UO_1973 (O_1973,N_26764,N_25025);
and UO_1974 (O_1974,N_26739,N_25325);
nand UO_1975 (O_1975,N_27737,N_29153);
xor UO_1976 (O_1976,N_27096,N_28670);
nor UO_1977 (O_1977,N_27306,N_28755);
nand UO_1978 (O_1978,N_28658,N_27975);
nor UO_1979 (O_1979,N_28476,N_27062);
nor UO_1980 (O_1980,N_25418,N_28137);
xnor UO_1981 (O_1981,N_25017,N_29038);
or UO_1982 (O_1982,N_27762,N_27449);
nand UO_1983 (O_1983,N_27825,N_29358);
and UO_1984 (O_1984,N_29811,N_27352);
nor UO_1985 (O_1985,N_27732,N_25713);
nand UO_1986 (O_1986,N_27588,N_25804);
and UO_1987 (O_1987,N_25666,N_25311);
or UO_1988 (O_1988,N_29145,N_27948);
or UO_1989 (O_1989,N_28858,N_27830);
nor UO_1990 (O_1990,N_25207,N_25568);
nor UO_1991 (O_1991,N_28125,N_27753);
or UO_1992 (O_1992,N_25771,N_27594);
or UO_1993 (O_1993,N_29104,N_27805);
or UO_1994 (O_1994,N_28114,N_28259);
xor UO_1995 (O_1995,N_25397,N_25990);
and UO_1996 (O_1996,N_28052,N_25931);
nor UO_1997 (O_1997,N_25820,N_27444);
xor UO_1998 (O_1998,N_25282,N_27514);
or UO_1999 (O_1999,N_25564,N_28941);
and UO_2000 (O_2000,N_27018,N_28739);
and UO_2001 (O_2001,N_28735,N_26997);
or UO_2002 (O_2002,N_29436,N_27101);
xnor UO_2003 (O_2003,N_29246,N_28716);
nand UO_2004 (O_2004,N_27355,N_27052);
nor UO_2005 (O_2005,N_28295,N_27120);
xor UO_2006 (O_2006,N_28797,N_25055);
or UO_2007 (O_2007,N_28333,N_28957);
and UO_2008 (O_2008,N_27919,N_28262);
nand UO_2009 (O_2009,N_25552,N_28126);
xnor UO_2010 (O_2010,N_27366,N_28220);
and UO_2011 (O_2011,N_28619,N_25035);
and UO_2012 (O_2012,N_26728,N_28837);
nor UO_2013 (O_2013,N_29861,N_29958);
nor UO_2014 (O_2014,N_29666,N_29521);
nor UO_2015 (O_2015,N_26009,N_27115);
nor UO_2016 (O_2016,N_27584,N_27208);
and UO_2017 (O_2017,N_27407,N_28431);
and UO_2018 (O_2018,N_27111,N_27347);
or UO_2019 (O_2019,N_27887,N_28657);
and UO_2020 (O_2020,N_29406,N_27838);
nand UO_2021 (O_2021,N_25688,N_26643);
nor UO_2022 (O_2022,N_26944,N_27039);
or UO_2023 (O_2023,N_25149,N_28019);
and UO_2024 (O_2024,N_29314,N_25509);
or UO_2025 (O_2025,N_29755,N_28472);
nand UO_2026 (O_2026,N_25125,N_28018);
and UO_2027 (O_2027,N_25843,N_28265);
xor UO_2028 (O_2028,N_26280,N_27011);
nand UO_2029 (O_2029,N_27272,N_27476);
and UO_2030 (O_2030,N_28692,N_29040);
nor UO_2031 (O_2031,N_27092,N_27246);
or UO_2032 (O_2032,N_26047,N_25793);
or UO_2033 (O_2033,N_26684,N_27430);
xnor UO_2034 (O_2034,N_26415,N_28541);
or UO_2035 (O_2035,N_26864,N_25592);
nor UO_2036 (O_2036,N_27036,N_28082);
nand UO_2037 (O_2037,N_25525,N_25846);
nand UO_2038 (O_2038,N_29370,N_26483);
nor UO_2039 (O_2039,N_29399,N_28863);
or UO_2040 (O_2040,N_28309,N_25358);
nand UO_2041 (O_2041,N_25952,N_25425);
nand UO_2042 (O_2042,N_28561,N_27280);
or UO_2043 (O_2043,N_29823,N_25211);
or UO_2044 (O_2044,N_25341,N_29525);
and UO_2045 (O_2045,N_27597,N_27499);
nand UO_2046 (O_2046,N_26219,N_28994);
xnor UO_2047 (O_2047,N_29060,N_26363);
and UO_2048 (O_2048,N_27646,N_28249);
xnor UO_2049 (O_2049,N_29649,N_25577);
nand UO_2050 (O_2050,N_26732,N_27908);
nor UO_2051 (O_2051,N_28044,N_27353);
and UO_2052 (O_2052,N_26024,N_27211);
nor UO_2053 (O_2053,N_28532,N_26951);
and UO_2054 (O_2054,N_29635,N_28713);
nand UO_2055 (O_2055,N_29804,N_27800);
nand UO_2056 (O_2056,N_27639,N_25075);
or UO_2057 (O_2057,N_27567,N_25723);
nand UO_2058 (O_2058,N_25037,N_25783);
xor UO_2059 (O_2059,N_28294,N_28610);
nor UO_2060 (O_2060,N_29552,N_27961);
and UO_2061 (O_2061,N_29350,N_25884);
nor UO_2062 (O_2062,N_27813,N_27875);
or UO_2063 (O_2063,N_27044,N_25104);
or UO_2064 (O_2064,N_27193,N_26568);
xnor UO_2065 (O_2065,N_26290,N_26904);
or UO_2066 (O_2066,N_25888,N_27531);
nor UO_2067 (O_2067,N_29112,N_28683);
nor UO_2068 (O_2068,N_29623,N_29028);
xnor UO_2069 (O_2069,N_25769,N_27247);
and UO_2070 (O_2070,N_25152,N_29000);
nor UO_2071 (O_2071,N_27854,N_27015);
or UO_2072 (O_2072,N_29597,N_28263);
nand UO_2073 (O_2073,N_29634,N_27686);
and UO_2074 (O_2074,N_29143,N_27053);
nand UO_2075 (O_2075,N_27423,N_28099);
or UO_2076 (O_2076,N_29164,N_28601);
and UO_2077 (O_2077,N_28686,N_25002);
or UO_2078 (O_2078,N_26879,N_25433);
nand UO_2079 (O_2079,N_28461,N_26933);
nand UO_2080 (O_2080,N_28785,N_26771);
xor UO_2081 (O_2081,N_29829,N_27314);
or UO_2082 (O_2082,N_29036,N_29613);
nor UO_2083 (O_2083,N_28990,N_27010);
or UO_2084 (O_2084,N_26820,N_27429);
or UO_2085 (O_2085,N_27684,N_29833);
nand UO_2086 (O_2086,N_28079,N_26239);
nor UO_2087 (O_2087,N_29940,N_25294);
xor UO_2088 (O_2088,N_28048,N_27839);
xor UO_2089 (O_2089,N_29681,N_25081);
xor UO_2090 (O_2090,N_25400,N_28010);
xnor UO_2091 (O_2091,N_27959,N_25695);
xnor UO_2092 (O_2092,N_29772,N_27180);
nand UO_2093 (O_2093,N_27089,N_26950);
and UO_2094 (O_2094,N_27694,N_27418);
xor UO_2095 (O_2095,N_25188,N_25267);
xor UO_2096 (O_2096,N_26382,N_28524);
nand UO_2097 (O_2097,N_25450,N_27840);
xor UO_2098 (O_2098,N_27268,N_28563);
or UO_2099 (O_2099,N_26309,N_27566);
xor UO_2100 (O_2100,N_27462,N_26106);
nor UO_2101 (O_2101,N_27563,N_29694);
nand UO_2102 (O_2102,N_28632,N_26142);
xnor UO_2103 (O_2103,N_29622,N_26126);
and UO_2104 (O_2104,N_29444,N_27523);
xnor UO_2105 (O_2105,N_25490,N_29067);
nand UO_2106 (O_2106,N_25305,N_28315);
nand UO_2107 (O_2107,N_28088,N_29612);
and UO_2108 (O_2108,N_26214,N_29680);
nand UO_2109 (O_2109,N_28531,N_28790);
and UO_2110 (O_2110,N_27425,N_28367);
or UO_2111 (O_2111,N_25605,N_28971);
and UO_2112 (O_2112,N_26687,N_27267);
nor UO_2113 (O_2113,N_28507,N_27320);
nand UO_2114 (O_2114,N_25162,N_28055);
nand UO_2115 (O_2115,N_27513,N_29310);
or UO_2116 (O_2116,N_29078,N_26973);
xnor UO_2117 (O_2117,N_28152,N_25993);
nand UO_2118 (O_2118,N_27394,N_29368);
nor UO_2119 (O_2119,N_25365,N_28719);
nor UO_2120 (O_2120,N_29367,N_28512);
nand UO_2121 (O_2121,N_27402,N_25744);
nand UO_2122 (O_2122,N_28668,N_25892);
nand UO_2123 (O_2123,N_25254,N_27633);
and UO_2124 (O_2124,N_27238,N_27592);
xnor UO_2125 (O_2125,N_29476,N_25291);
and UO_2126 (O_2126,N_28433,N_28215);
xor UO_2127 (O_2127,N_26325,N_26380);
xnor UO_2128 (O_2128,N_29002,N_28558);
and UO_2129 (O_2129,N_25374,N_26227);
or UO_2130 (O_2130,N_28045,N_29891);
nand UO_2131 (O_2131,N_25058,N_25939);
and UO_2132 (O_2132,N_27522,N_28934);
xor UO_2133 (O_2133,N_29770,N_28550);
or UO_2134 (O_2134,N_28865,N_29605);
xnor UO_2135 (O_2135,N_26143,N_25609);
and UO_2136 (O_2136,N_25200,N_26093);
xnor UO_2137 (O_2137,N_29198,N_26562);
xor UO_2138 (O_2138,N_27190,N_29883);
and UO_2139 (O_2139,N_27763,N_26329);
or UO_2140 (O_2140,N_28743,N_26654);
nor UO_2141 (O_2141,N_28612,N_25051);
nor UO_2142 (O_2142,N_26478,N_27816);
and UO_2143 (O_2143,N_29225,N_29984);
xnor UO_2144 (O_2144,N_28290,N_27093);
nand UO_2145 (O_2145,N_28777,N_25719);
xnor UO_2146 (O_2146,N_25839,N_29121);
and UO_2147 (O_2147,N_27943,N_25822);
nand UO_2148 (O_2148,N_27688,N_27951);
nor UO_2149 (O_2149,N_28449,N_27672);
nand UO_2150 (O_2150,N_28813,N_29252);
and UO_2151 (O_2151,N_27383,N_25714);
or UO_2152 (O_2152,N_29598,N_27191);
or UO_2153 (O_2153,N_25879,N_27173);
nand UO_2154 (O_2154,N_27950,N_26133);
or UO_2155 (O_2155,N_29052,N_25834);
or UO_2156 (O_2156,N_29223,N_29282);
xnor UO_2157 (O_2157,N_26067,N_27543);
and UO_2158 (O_2158,N_27667,N_29509);
xnor UO_2159 (O_2159,N_26874,N_26014);
xnor UO_2160 (O_2160,N_26080,N_29517);
or UO_2161 (O_2161,N_26989,N_26504);
xor UO_2162 (O_2162,N_25889,N_29588);
or UO_2163 (O_2163,N_28113,N_27065);
or UO_2164 (O_2164,N_28311,N_28591);
nor UO_2165 (O_2165,N_29979,N_27575);
nand UO_2166 (O_2166,N_29359,N_26885);
xnor UO_2167 (O_2167,N_28523,N_28414);
or UO_2168 (O_2168,N_27972,N_27343);
nand UO_2169 (O_2169,N_28477,N_25530);
nand UO_2170 (O_2170,N_26929,N_25800);
or UO_2171 (O_2171,N_25030,N_27277);
xnor UO_2172 (O_2172,N_28627,N_27529);
nand UO_2173 (O_2173,N_27536,N_26109);
and UO_2174 (O_2174,N_29682,N_27357);
or UO_2175 (O_2175,N_28351,N_25286);
or UO_2176 (O_2176,N_28883,N_29270);
or UO_2177 (O_2177,N_27796,N_26914);
and UO_2178 (O_2178,N_25777,N_28893);
nor UO_2179 (O_2179,N_25340,N_26527);
nand UO_2180 (O_2180,N_27296,N_26615);
and UO_2181 (O_2181,N_28066,N_26090);
nor UO_2182 (O_2182,N_27713,N_28063);
xnor UO_2183 (O_2183,N_27163,N_29665);
nand UO_2184 (O_2184,N_26858,N_29330);
xor UO_2185 (O_2185,N_26936,N_29468);
nand UO_2186 (O_2186,N_27564,N_27535);
or UO_2187 (O_2187,N_26072,N_26168);
xnor UO_2188 (O_2188,N_28255,N_29716);
nand UO_2189 (O_2189,N_25739,N_28678);
nor UO_2190 (O_2190,N_27701,N_29303);
nor UO_2191 (O_2191,N_28094,N_25812);
nor UO_2192 (O_2192,N_26787,N_25686);
and UO_2193 (O_2193,N_27632,N_26393);
xor UO_2194 (O_2194,N_28530,N_29023);
xnor UO_2195 (O_2195,N_26484,N_28810);
nor UO_2196 (O_2196,N_26053,N_29571);
xnor UO_2197 (O_2197,N_27909,N_27847);
or UO_2198 (O_2198,N_26201,N_26323);
nor UO_2199 (O_2199,N_28418,N_27309);
or UO_2200 (O_2200,N_29538,N_27822);
or UO_2201 (O_2201,N_27548,N_27780);
nor UO_2202 (O_2202,N_26792,N_26566);
or UO_2203 (O_2203,N_25119,N_25335);
or UO_2204 (O_2204,N_27436,N_27409);
and UO_2205 (O_2205,N_26612,N_27008);
nor UO_2206 (O_2206,N_28352,N_25006);
xnor UO_2207 (O_2207,N_26837,N_28624);
xnor UO_2208 (O_2208,N_29702,N_29757);
and UO_2209 (O_2209,N_28073,N_26314);
nand UO_2210 (O_2210,N_29800,N_25381);
xnor UO_2211 (O_2211,N_28513,N_27195);
nand UO_2212 (O_2212,N_25716,N_25466);
xnor UO_2213 (O_2213,N_25541,N_26266);
xnor UO_2214 (O_2214,N_29438,N_27744);
nor UO_2215 (O_2215,N_25513,N_29328);
xnor UO_2216 (O_2216,N_25855,N_28024);
nand UO_2217 (O_2217,N_28780,N_28256);
nand UO_2218 (O_2218,N_29413,N_25556);
and UO_2219 (O_2219,N_26041,N_26805);
nor UO_2220 (O_2220,N_25232,N_26021);
nor UO_2221 (O_2221,N_25039,N_28488);
or UO_2222 (O_2222,N_25324,N_29169);
xnor UO_2223 (O_2223,N_27412,N_28261);
or UO_2224 (O_2224,N_28728,N_28915);
and UO_2225 (O_2225,N_28382,N_29942);
or UO_2226 (O_2226,N_27785,N_26434);
and UO_2227 (O_2227,N_28175,N_27720);
or UO_2228 (O_2228,N_29976,N_26844);
or UO_2229 (O_2229,N_26279,N_27054);
or UO_2230 (O_2230,N_26716,N_26493);
nor UO_2231 (O_2231,N_28474,N_26264);
xnor UO_2232 (O_2232,N_25321,N_29910);
and UO_2233 (O_2233,N_27843,N_27248);
and UO_2234 (O_2234,N_29547,N_29416);
xor UO_2235 (O_2235,N_29777,N_27292);
nor UO_2236 (O_2236,N_25798,N_27917);
nand UO_2237 (O_2237,N_29157,N_26769);
nand UO_2238 (O_2238,N_28095,N_28402);
and UO_2239 (O_2239,N_26398,N_28264);
or UO_2240 (O_2240,N_28698,N_26069);
nand UO_2241 (O_2241,N_25946,N_25079);
and UO_2242 (O_2242,N_29363,N_29054);
nor UO_2243 (O_2243,N_27023,N_29431);
and UO_2244 (O_2244,N_27724,N_28968);
or UO_2245 (O_2245,N_26665,N_27077);
or UO_2246 (O_2246,N_25122,N_28178);
xor UO_2247 (O_2247,N_29418,N_28933);
nor UO_2248 (O_2248,N_29019,N_28546);
nand UO_2249 (O_2249,N_29408,N_29381);
or UO_2250 (O_2250,N_28663,N_29427);
nor UO_2251 (O_2251,N_25073,N_28606);
or UO_2252 (O_2252,N_26757,N_25837);
xnor UO_2253 (O_2253,N_25375,N_28271);
and UO_2254 (O_2254,N_27858,N_26573);
xor UO_2255 (O_2255,N_25416,N_26714);
nor UO_2256 (O_2256,N_25501,N_29135);
or UO_2257 (O_2257,N_28902,N_27310);
nor UO_2258 (O_2258,N_29103,N_27512);
and UO_2259 (O_2259,N_26141,N_26517);
xor UO_2260 (O_2260,N_29471,N_25446);
nand UO_2261 (O_2261,N_29615,N_28091);
nor UO_2262 (O_2262,N_26609,N_26845);
or UO_2263 (O_2263,N_27613,N_27648);
and UO_2264 (O_2264,N_26578,N_28188);
and UO_2265 (O_2265,N_29786,N_27351);
nand UO_2266 (O_2266,N_27577,N_29551);
nand UO_2267 (O_2267,N_26735,N_29323);
nand UO_2268 (O_2268,N_26243,N_25016);
nor UO_2269 (O_2269,N_26040,N_27899);
xnor UO_2270 (O_2270,N_27538,N_29278);
or UO_2271 (O_2271,N_26140,N_25527);
xnor UO_2272 (O_2272,N_26550,N_25368);
xor UO_2273 (O_2273,N_26187,N_29663);
nand UO_2274 (O_2274,N_25615,N_29441);
nor UO_2275 (O_2275,N_25302,N_28151);
nand UO_2276 (O_2276,N_25599,N_25087);
nor UO_2277 (O_2277,N_26333,N_27581);
xor UO_2278 (O_2278,N_26211,N_28384);
or UO_2279 (O_2279,N_29880,N_25465);
or UO_2280 (O_2280,N_29874,N_29751);
xor UO_2281 (O_2281,N_28153,N_27874);
or UO_2282 (O_2282,N_29696,N_29867);
xnor UO_2283 (O_2283,N_26235,N_26317);
nor UO_2284 (O_2284,N_29275,N_29808);
and UO_2285 (O_2285,N_25181,N_26782);
xor UO_2286 (O_2286,N_29214,N_29070);
xor UO_2287 (O_2287,N_27953,N_29499);
or UO_2288 (O_2288,N_28283,N_26129);
and UO_2289 (O_2289,N_27460,N_29763);
and UO_2290 (O_2290,N_25141,N_25462);
and UO_2291 (O_2291,N_29671,N_25842);
nor UO_2292 (O_2292,N_25873,N_26583);
and UO_2293 (O_2293,N_29908,N_27066);
nor UO_2294 (O_2294,N_26305,N_25069);
and UO_2295 (O_2295,N_26430,N_29895);
or UO_2296 (O_2296,N_27137,N_25927);
or UO_2297 (O_2297,N_26426,N_28146);
nand UO_2298 (O_2298,N_28232,N_25913);
nand UO_2299 (O_2299,N_25013,N_26818);
nand UO_2300 (O_2300,N_27644,N_26076);
xnor UO_2301 (O_2301,N_29807,N_29652);
nand UO_2302 (O_2302,N_26669,N_28914);
xor UO_2303 (O_2303,N_26086,N_28463);
and UO_2304 (O_2304,N_27913,N_25845);
xnor UO_2305 (O_2305,N_25833,N_27229);
nor UO_2306 (O_2306,N_27795,N_28614);
xnor UO_2307 (O_2307,N_25601,N_28109);
xor UO_2308 (O_2308,N_27749,N_27216);
or UO_2309 (O_2309,N_26336,N_29369);
nor UO_2310 (O_2310,N_26376,N_27783);
or UO_2311 (O_2311,N_27465,N_28652);
xnor UO_2312 (O_2312,N_26485,N_28411);
xnor UO_2313 (O_2313,N_25631,N_27237);
or UO_2314 (O_2314,N_27956,N_25698);
or UO_2315 (O_2315,N_27300,N_25496);
nor UO_2316 (O_2316,N_27354,N_29731);
xor UO_2317 (O_2317,N_27489,N_25984);
xor UO_2318 (O_2318,N_27219,N_25154);
or UO_2319 (O_2319,N_28227,N_26946);
or UO_2320 (O_2320,N_26412,N_27185);
nand UO_2321 (O_2321,N_26070,N_29361);
nand UO_2322 (O_2322,N_25988,N_29784);
nor UO_2323 (O_2323,N_26906,N_26968);
nor UO_2324 (O_2324,N_27640,N_27696);
or UO_2325 (O_2325,N_28173,N_26400);
or UO_2326 (O_2326,N_29012,N_28308);
nor UO_2327 (O_2327,N_25517,N_29774);
or UO_2328 (O_2328,N_29840,N_25661);
xnor UO_2329 (O_2329,N_26923,N_28715);
nand UO_2330 (O_2330,N_27643,N_29916);
nor UO_2331 (O_2331,N_27560,N_28217);
nor UO_2332 (O_2332,N_26591,N_27865);
nand UO_2333 (O_2333,N_29415,N_25212);
nand UO_2334 (O_2334,N_26012,N_27790);
nand UO_2335 (O_2335,N_26298,N_29081);
nand UO_2336 (O_2336,N_27373,N_27747);
nand UO_2337 (O_2337,N_29797,N_29378);
and UO_2338 (O_2338,N_27715,N_25765);
nor UO_2339 (O_2339,N_26613,N_28904);
nor UO_2340 (O_2340,N_29291,N_27435);
or UO_2341 (O_2341,N_28436,N_28649);
nor UO_2342 (O_2342,N_26723,N_25600);
nand UO_2343 (O_2343,N_27106,N_27595);
nand UO_2344 (O_2344,N_29553,N_25498);
xnor UO_2345 (O_2345,N_27532,N_27903);
and UO_2346 (O_2346,N_25786,N_26464);
nand UO_2347 (O_2347,N_27922,N_29493);
or UO_2348 (O_2348,N_27934,N_25251);
nand UO_2349 (O_2349,N_25394,N_26646);
or UO_2350 (O_2350,N_25332,N_27496);
or UO_2351 (O_2351,N_28184,N_29966);
nand UO_2352 (O_2352,N_26509,N_29723);
xor UO_2353 (O_2353,N_26494,N_27774);
xnor UO_2354 (O_2354,N_29170,N_27283);
nand UO_2355 (O_2355,N_26754,N_26762);
nand UO_2356 (O_2356,N_25389,N_27113);
or UO_2357 (O_2357,N_26157,N_28413);
and UO_2358 (O_2358,N_29564,N_25179);
or UO_2359 (O_2359,N_28679,N_26763);
nor UO_2360 (O_2360,N_27980,N_29814);
and UO_2361 (O_2361,N_28768,N_28824);
nand UO_2362 (O_2362,N_28602,N_28252);
xor UO_2363 (O_2363,N_27561,N_28514);
xor UO_2364 (O_2364,N_26354,N_25437);
and UO_2365 (O_2365,N_29877,N_27993);
xnor UO_2366 (O_2366,N_28229,N_26865);
nor UO_2367 (O_2367,N_27627,N_27055);
xnor UO_2368 (O_2368,N_29902,N_26563);
xnor UO_2369 (O_2369,N_28098,N_27849);
xor UO_2370 (O_2370,N_29964,N_28361);
nand UO_2371 (O_2371,N_26068,N_27954);
or UO_2372 (O_2372,N_29722,N_29484);
and UO_2373 (O_2373,N_25463,N_25738);
nand UO_2374 (O_2374,N_29050,N_29920);
and UO_2375 (O_2375,N_27399,N_27400);
and UO_2376 (O_2376,N_26756,N_27471);
or UO_2377 (O_2377,N_28492,N_27164);
and UO_2378 (O_2378,N_29825,N_28289);
or UO_2379 (O_2379,N_27207,N_29017);
xnor UO_2380 (O_2380,N_25950,N_27555);
xnor UO_2381 (O_2381,N_28842,N_28930);
xnor UO_2382 (O_2382,N_28332,N_25423);
nand UO_2383 (O_2383,N_26461,N_28770);
and UO_2384 (O_2384,N_27547,N_27130);
nand UO_2385 (O_2385,N_26172,N_27662);
nand UO_2386 (O_2386,N_28745,N_29998);
nand UO_2387 (O_2387,N_26584,N_29690);
or UO_2388 (O_2388,N_29166,N_29620);
and UO_2389 (O_2389,N_26375,N_26185);
nand UO_2390 (O_2390,N_27241,N_26678);
nor UO_2391 (O_2391,N_26057,N_29953);
nand UO_2392 (O_2392,N_29174,N_29638);
and UO_2393 (O_2393,N_26555,N_26406);
and UO_2394 (O_2394,N_26066,N_25322);
or UO_2395 (O_2395,N_26344,N_28821);
xnor UO_2396 (O_2396,N_26571,N_27289);
and UO_2397 (O_2397,N_28160,N_26598);
nor UO_2398 (O_2398,N_25161,N_26377);
nand UO_2399 (O_2399,N_29970,N_28301);
nand UO_2400 (O_2400,N_27960,N_27305);
xnor UO_2401 (O_2401,N_25826,N_27895);
or UO_2402 (O_2402,N_28970,N_25531);
nand UO_2403 (O_2403,N_26034,N_27844);
nand UO_2404 (O_2404,N_25410,N_29478);
and UO_2405 (O_2405,N_29256,N_28937);
xor UO_2406 (O_2406,N_29294,N_25522);
xnor UO_2407 (O_2407,N_28493,N_26401);
nor UO_2408 (O_2408,N_26861,N_27097);
nor UO_2409 (O_2409,N_29606,N_28059);
nand UO_2410 (O_2410,N_25151,N_29555);
or UO_2411 (O_2411,N_29109,N_26812);
xnor UO_2412 (O_2412,N_26977,N_29875);
nor UO_2413 (O_2413,N_27141,N_29506);
nor UO_2414 (O_2414,N_27042,N_25460);
or UO_2415 (O_2415,N_27569,N_26685);
and UO_2416 (O_2416,N_25645,N_27179);
nand UO_2417 (O_2417,N_25392,N_26213);
and UO_2418 (O_2418,N_27864,N_25828);
or UO_2419 (O_2419,N_25664,N_28769);
nand UO_2420 (O_2420,N_26476,N_27967);
or UO_2421 (O_2421,N_28427,N_25172);
xnor UO_2422 (O_2422,N_26221,N_26682);
and UO_2423 (O_2423,N_26297,N_29893);
nand UO_2424 (O_2424,N_29936,N_26491);
or UO_2425 (O_2425,N_29733,N_27894);
and UO_2426 (O_2426,N_28977,N_26692);
xnor UO_2427 (O_2427,N_29851,N_27432);
or UO_2428 (O_2428,N_28208,N_25133);
or UO_2429 (O_2429,N_25627,N_29130);
nand UO_2430 (O_2430,N_25853,N_26387);
nand UO_2431 (O_2431,N_29074,N_26045);
xnor UO_2432 (O_2432,N_27004,N_27480);
nor UO_2433 (O_2433,N_26098,N_29852);
nor UO_2434 (O_2434,N_27001,N_29005);
or UO_2435 (O_2435,N_26242,N_25681);
and UO_2436 (O_2436,N_25348,N_27025);
nand UO_2437 (O_2437,N_28186,N_25639);
nand UO_2438 (O_2438,N_26894,N_28168);
nand UO_2439 (O_2439,N_27405,N_28430);
xnor UO_2440 (O_2440,N_26930,N_26134);
nor UO_2441 (O_2441,N_25507,N_26990);
xnor UO_2442 (O_2442,N_29847,N_28701);
and UO_2443 (O_2443,N_26396,N_26360);
nor UO_2444 (O_2444,N_26986,N_26296);
nand UO_2445 (O_2445,N_26910,N_26477);
and UO_2446 (O_2446,N_25893,N_27365);
nor UO_2447 (O_2447,N_25401,N_28327);
nand UO_2448 (O_2448,N_27650,N_25191);
xnor UO_2449 (O_2449,N_28396,N_26846);
nand UO_2450 (O_2450,N_28317,N_25135);
xor UO_2451 (O_2451,N_28993,N_26244);
and UO_2452 (O_2452,N_25128,N_26741);
nor UO_2453 (O_2453,N_29026,N_25970);
and UO_2454 (O_2454,N_28456,N_28226);
nor UO_2455 (O_2455,N_28004,N_28330);
or UO_2456 (O_2456,N_27794,N_29316);
xor UO_2457 (O_2457,N_29280,N_26644);
nand UO_2458 (O_2458,N_29313,N_25169);
or UO_2459 (O_2459,N_27729,N_25628);
nand UO_2460 (O_2460,N_25344,N_26416);
nor UO_2461 (O_2461,N_25109,N_28451);
nand UO_2462 (O_2462,N_25630,N_28568);
and UO_2463 (O_2463,N_26860,N_27905);
or UO_2464 (O_2464,N_28784,N_28534);
or UO_2465 (O_2465,N_29177,N_27076);
and UO_2466 (O_2466,N_27417,N_29999);
nor UO_2467 (O_2467,N_25538,N_29306);
or UO_2468 (O_2468,N_29708,N_28540);
nor UO_2469 (O_2469,N_29841,N_27021);
xor UO_2470 (O_2470,N_26481,N_27710);
nand UO_2471 (O_2471,N_26940,N_29817);
and UO_2472 (O_2472,N_25764,N_29675);
nand UO_2473 (O_2473,N_25947,N_26924);
nor UO_2474 (O_2474,N_27620,N_29746);
and UO_2475 (O_2475,N_28041,N_29461);
xnor UO_2476 (O_2476,N_27574,N_25408);
or UO_2477 (O_2477,N_27050,N_26748);
nor UO_2478 (O_2478,N_29981,N_26078);
and UO_2479 (O_2479,N_27784,N_28763);
xor UO_2480 (O_2480,N_27933,N_27340);
or UO_2481 (O_2481,N_25326,N_25923);
nand UO_2482 (O_2482,N_25178,N_26361);
xor UO_2483 (O_2483,N_26038,N_29706);
and UO_2484 (O_2484,N_27506,N_27144);
or UO_2485 (O_2485,N_26520,N_27625);
and UO_2486 (O_2486,N_25998,N_25431);
xnor UO_2487 (O_2487,N_26315,N_27291);
nand UO_2488 (O_2488,N_26095,N_27925);
nor UO_2489 (O_2489,N_28909,N_25867);
xor UO_2490 (O_2490,N_29560,N_26642);
nand UO_2491 (O_2491,N_26576,N_27572);
nand UO_2492 (O_2492,N_29452,N_26617);
nand UO_2493 (O_2493,N_27867,N_29667);
and UO_2494 (O_2494,N_27031,N_29141);
xor UO_2495 (O_2495,N_29677,N_29977);
or UO_2496 (O_2496,N_29462,N_27372);
or UO_2497 (O_2497,N_29393,N_25373);
and UO_2498 (O_2498,N_29375,N_25252);
and UO_2499 (O_2499,N_29196,N_27479);
nand UO_2500 (O_2500,N_27448,N_26294);
nand UO_2501 (O_2501,N_27909,N_28440);
nand UO_2502 (O_2502,N_25893,N_25381);
xor UO_2503 (O_2503,N_26995,N_25952);
nor UO_2504 (O_2504,N_25710,N_25660);
or UO_2505 (O_2505,N_26006,N_26683);
nand UO_2506 (O_2506,N_27217,N_29559);
nor UO_2507 (O_2507,N_27879,N_28184);
and UO_2508 (O_2508,N_26710,N_29715);
xnor UO_2509 (O_2509,N_29872,N_28755);
and UO_2510 (O_2510,N_29451,N_28954);
and UO_2511 (O_2511,N_27909,N_25683);
nor UO_2512 (O_2512,N_26830,N_25868);
xor UO_2513 (O_2513,N_25080,N_25915);
xnor UO_2514 (O_2514,N_28268,N_28681);
nand UO_2515 (O_2515,N_29031,N_26630);
or UO_2516 (O_2516,N_26989,N_26268);
nor UO_2517 (O_2517,N_29246,N_25941);
nor UO_2518 (O_2518,N_26231,N_26822);
nor UO_2519 (O_2519,N_28828,N_27877);
or UO_2520 (O_2520,N_26266,N_29740);
or UO_2521 (O_2521,N_25896,N_26528);
or UO_2522 (O_2522,N_26744,N_26877);
or UO_2523 (O_2523,N_29338,N_29725);
or UO_2524 (O_2524,N_27516,N_26279);
and UO_2525 (O_2525,N_26466,N_28563);
nor UO_2526 (O_2526,N_25613,N_29481);
xnor UO_2527 (O_2527,N_29982,N_27817);
nand UO_2528 (O_2528,N_27048,N_25605);
nand UO_2529 (O_2529,N_25947,N_25213);
nand UO_2530 (O_2530,N_28797,N_26905);
xnor UO_2531 (O_2531,N_29901,N_28662);
nand UO_2532 (O_2532,N_29327,N_27083);
nand UO_2533 (O_2533,N_29304,N_28271);
nor UO_2534 (O_2534,N_27759,N_29910);
xor UO_2535 (O_2535,N_29632,N_28170);
or UO_2536 (O_2536,N_25631,N_29781);
nand UO_2537 (O_2537,N_25574,N_29948);
or UO_2538 (O_2538,N_25011,N_26997);
nand UO_2539 (O_2539,N_27574,N_28191);
xor UO_2540 (O_2540,N_27011,N_26304);
nor UO_2541 (O_2541,N_28107,N_25420);
or UO_2542 (O_2542,N_29545,N_25658);
nor UO_2543 (O_2543,N_29575,N_25851);
nor UO_2544 (O_2544,N_28445,N_29498);
nand UO_2545 (O_2545,N_27914,N_26019);
and UO_2546 (O_2546,N_26290,N_25259);
xor UO_2547 (O_2547,N_28383,N_27352);
nand UO_2548 (O_2548,N_27409,N_29287);
nor UO_2549 (O_2549,N_27671,N_27227);
nor UO_2550 (O_2550,N_25388,N_26259);
or UO_2551 (O_2551,N_27897,N_29439);
and UO_2552 (O_2552,N_27116,N_26571);
xnor UO_2553 (O_2553,N_25758,N_25937);
xnor UO_2554 (O_2554,N_28059,N_28218);
nor UO_2555 (O_2555,N_28610,N_28516);
nor UO_2556 (O_2556,N_28265,N_29738);
xor UO_2557 (O_2557,N_26563,N_26772);
nor UO_2558 (O_2558,N_26438,N_28695);
and UO_2559 (O_2559,N_27086,N_29205);
nand UO_2560 (O_2560,N_29984,N_29748);
nand UO_2561 (O_2561,N_26022,N_26822);
xnor UO_2562 (O_2562,N_27185,N_29798);
nand UO_2563 (O_2563,N_26619,N_25353);
nor UO_2564 (O_2564,N_27138,N_29270);
or UO_2565 (O_2565,N_27585,N_28947);
and UO_2566 (O_2566,N_25122,N_28751);
nor UO_2567 (O_2567,N_29541,N_26322);
or UO_2568 (O_2568,N_29222,N_28402);
nand UO_2569 (O_2569,N_26831,N_29158);
or UO_2570 (O_2570,N_28288,N_27994);
nor UO_2571 (O_2571,N_28794,N_26065);
nand UO_2572 (O_2572,N_27037,N_27803);
nand UO_2573 (O_2573,N_28284,N_25987);
xnor UO_2574 (O_2574,N_25603,N_26197);
nand UO_2575 (O_2575,N_27182,N_27228);
nand UO_2576 (O_2576,N_27794,N_26015);
and UO_2577 (O_2577,N_26298,N_27520);
or UO_2578 (O_2578,N_25769,N_26912);
nor UO_2579 (O_2579,N_26880,N_29003);
nor UO_2580 (O_2580,N_28822,N_28792);
xor UO_2581 (O_2581,N_27690,N_25977);
nor UO_2582 (O_2582,N_25797,N_28354);
xor UO_2583 (O_2583,N_26216,N_25795);
nand UO_2584 (O_2584,N_25811,N_27776);
and UO_2585 (O_2585,N_27262,N_26462);
and UO_2586 (O_2586,N_28083,N_28482);
xnor UO_2587 (O_2587,N_28936,N_27754);
xnor UO_2588 (O_2588,N_27735,N_28710);
xnor UO_2589 (O_2589,N_26102,N_25164);
nand UO_2590 (O_2590,N_29797,N_28049);
and UO_2591 (O_2591,N_29387,N_26879);
nor UO_2592 (O_2592,N_28556,N_26773);
nand UO_2593 (O_2593,N_29387,N_27867);
and UO_2594 (O_2594,N_29655,N_28317);
nand UO_2595 (O_2595,N_26858,N_28744);
or UO_2596 (O_2596,N_28404,N_28524);
and UO_2597 (O_2597,N_25794,N_29570);
nand UO_2598 (O_2598,N_26050,N_25460);
xnor UO_2599 (O_2599,N_28812,N_26655);
nand UO_2600 (O_2600,N_25764,N_29850);
and UO_2601 (O_2601,N_26198,N_26605);
nand UO_2602 (O_2602,N_28957,N_27555);
xnor UO_2603 (O_2603,N_28744,N_25386);
and UO_2604 (O_2604,N_26013,N_29553);
xnor UO_2605 (O_2605,N_25987,N_29923);
nor UO_2606 (O_2606,N_28835,N_26869);
and UO_2607 (O_2607,N_26188,N_26318);
nand UO_2608 (O_2608,N_28130,N_26947);
nand UO_2609 (O_2609,N_26116,N_27873);
nor UO_2610 (O_2610,N_29765,N_26366);
or UO_2611 (O_2611,N_27987,N_26979);
xnor UO_2612 (O_2612,N_27374,N_28055);
nand UO_2613 (O_2613,N_25845,N_27352);
nor UO_2614 (O_2614,N_29881,N_28896);
xor UO_2615 (O_2615,N_28035,N_25807);
nand UO_2616 (O_2616,N_25555,N_25353);
nor UO_2617 (O_2617,N_29387,N_27804);
and UO_2618 (O_2618,N_26853,N_26346);
or UO_2619 (O_2619,N_29842,N_29795);
or UO_2620 (O_2620,N_26190,N_25088);
nor UO_2621 (O_2621,N_26980,N_29007);
and UO_2622 (O_2622,N_27498,N_28042);
nor UO_2623 (O_2623,N_25128,N_29159);
or UO_2624 (O_2624,N_25820,N_26697);
nand UO_2625 (O_2625,N_27273,N_28091);
and UO_2626 (O_2626,N_25499,N_29117);
and UO_2627 (O_2627,N_29213,N_29021);
or UO_2628 (O_2628,N_27366,N_28916);
xor UO_2629 (O_2629,N_27038,N_29892);
xnor UO_2630 (O_2630,N_27076,N_26582);
and UO_2631 (O_2631,N_26218,N_27785);
xor UO_2632 (O_2632,N_29608,N_25497);
or UO_2633 (O_2633,N_26153,N_25763);
xor UO_2634 (O_2634,N_26374,N_26077);
nor UO_2635 (O_2635,N_28500,N_27173);
nand UO_2636 (O_2636,N_26115,N_28842);
or UO_2637 (O_2637,N_29830,N_28129);
xnor UO_2638 (O_2638,N_27446,N_29736);
xnor UO_2639 (O_2639,N_29576,N_29993);
xor UO_2640 (O_2640,N_25875,N_27303);
xor UO_2641 (O_2641,N_25998,N_27629);
and UO_2642 (O_2642,N_29868,N_29796);
nand UO_2643 (O_2643,N_25808,N_28131);
xor UO_2644 (O_2644,N_25191,N_26122);
or UO_2645 (O_2645,N_29562,N_25512);
or UO_2646 (O_2646,N_25349,N_28391);
or UO_2647 (O_2647,N_26091,N_25483);
nand UO_2648 (O_2648,N_27571,N_29013);
and UO_2649 (O_2649,N_28621,N_27514);
or UO_2650 (O_2650,N_25555,N_27693);
or UO_2651 (O_2651,N_26276,N_28313);
nor UO_2652 (O_2652,N_29265,N_28120);
nand UO_2653 (O_2653,N_25368,N_29016);
and UO_2654 (O_2654,N_28472,N_27024);
xor UO_2655 (O_2655,N_29082,N_26666);
nor UO_2656 (O_2656,N_25757,N_26121);
and UO_2657 (O_2657,N_28305,N_29086);
nand UO_2658 (O_2658,N_28202,N_26151);
nand UO_2659 (O_2659,N_29294,N_27070);
xnor UO_2660 (O_2660,N_25460,N_26573);
nand UO_2661 (O_2661,N_29383,N_28085);
nor UO_2662 (O_2662,N_28455,N_25037);
nand UO_2663 (O_2663,N_26437,N_28260);
nand UO_2664 (O_2664,N_25130,N_25618);
and UO_2665 (O_2665,N_28108,N_25995);
xnor UO_2666 (O_2666,N_27081,N_28254);
nor UO_2667 (O_2667,N_26498,N_25795);
and UO_2668 (O_2668,N_25706,N_29877);
xnor UO_2669 (O_2669,N_25225,N_27075);
xor UO_2670 (O_2670,N_26385,N_28346);
or UO_2671 (O_2671,N_26439,N_26694);
nor UO_2672 (O_2672,N_26098,N_28622);
xor UO_2673 (O_2673,N_27928,N_25415);
nand UO_2674 (O_2674,N_25952,N_26289);
and UO_2675 (O_2675,N_26686,N_28621);
and UO_2676 (O_2676,N_25189,N_27630);
nor UO_2677 (O_2677,N_25310,N_27395);
xnor UO_2678 (O_2678,N_25282,N_26925);
xor UO_2679 (O_2679,N_28789,N_29040);
nand UO_2680 (O_2680,N_28565,N_25934);
nor UO_2681 (O_2681,N_26598,N_28290);
xor UO_2682 (O_2682,N_28438,N_25625);
and UO_2683 (O_2683,N_28074,N_29775);
or UO_2684 (O_2684,N_26663,N_28462);
or UO_2685 (O_2685,N_25936,N_28246);
xnor UO_2686 (O_2686,N_28065,N_28496);
and UO_2687 (O_2687,N_25015,N_26858);
nand UO_2688 (O_2688,N_26215,N_29369);
nor UO_2689 (O_2689,N_27633,N_27963);
and UO_2690 (O_2690,N_25454,N_29456);
nor UO_2691 (O_2691,N_29313,N_25348);
nand UO_2692 (O_2692,N_26422,N_26933);
nor UO_2693 (O_2693,N_28413,N_25448);
or UO_2694 (O_2694,N_29664,N_29461);
nor UO_2695 (O_2695,N_27771,N_29914);
xor UO_2696 (O_2696,N_29663,N_27032);
nor UO_2697 (O_2697,N_29345,N_27378);
nand UO_2698 (O_2698,N_25275,N_26286);
and UO_2699 (O_2699,N_29929,N_26588);
and UO_2700 (O_2700,N_29903,N_29137);
and UO_2701 (O_2701,N_26760,N_26860);
nor UO_2702 (O_2702,N_25964,N_27765);
nand UO_2703 (O_2703,N_26367,N_29423);
xor UO_2704 (O_2704,N_29018,N_28067);
and UO_2705 (O_2705,N_25468,N_25598);
xor UO_2706 (O_2706,N_25006,N_28529);
and UO_2707 (O_2707,N_27197,N_27242);
nor UO_2708 (O_2708,N_28981,N_25242);
nor UO_2709 (O_2709,N_29858,N_29221);
or UO_2710 (O_2710,N_27469,N_26249);
or UO_2711 (O_2711,N_28769,N_25835);
nor UO_2712 (O_2712,N_25317,N_29422);
or UO_2713 (O_2713,N_25568,N_25273);
nand UO_2714 (O_2714,N_26024,N_26664);
xnor UO_2715 (O_2715,N_27924,N_26321);
nor UO_2716 (O_2716,N_25388,N_27222);
nor UO_2717 (O_2717,N_25452,N_27291);
or UO_2718 (O_2718,N_28351,N_29489);
nor UO_2719 (O_2719,N_26076,N_25447);
and UO_2720 (O_2720,N_28978,N_29972);
xor UO_2721 (O_2721,N_26563,N_28448);
xor UO_2722 (O_2722,N_27796,N_27461);
xnor UO_2723 (O_2723,N_25912,N_29735);
nand UO_2724 (O_2724,N_26789,N_28187);
nand UO_2725 (O_2725,N_27158,N_29404);
nor UO_2726 (O_2726,N_29399,N_27758);
or UO_2727 (O_2727,N_29605,N_26198);
nand UO_2728 (O_2728,N_26343,N_27948);
or UO_2729 (O_2729,N_27078,N_25562);
or UO_2730 (O_2730,N_29008,N_26811);
xor UO_2731 (O_2731,N_28377,N_29380);
xor UO_2732 (O_2732,N_28457,N_29766);
and UO_2733 (O_2733,N_25965,N_25868);
or UO_2734 (O_2734,N_29992,N_25612);
xor UO_2735 (O_2735,N_28885,N_28805);
or UO_2736 (O_2736,N_28647,N_27795);
xor UO_2737 (O_2737,N_29963,N_29288);
nand UO_2738 (O_2738,N_26580,N_25699);
xnor UO_2739 (O_2739,N_28384,N_29882);
xnor UO_2740 (O_2740,N_28034,N_25207);
xnor UO_2741 (O_2741,N_25142,N_25674);
or UO_2742 (O_2742,N_29787,N_28622);
nor UO_2743 (O_2743,N_27797,N_28908);
xor UO_2744 (O_2744,N_28804,N_29811);
and UO_2745 (O_2745,N_26887,N_27313);
nand UO_2746 (O_2746,N_29313,N_26687);
nand UO_2747 (O_2747,N_27679,N_25660);
and UO_2748 (O_2748,N_27052,N_28490);
nand UO_2749 (O_2749,N_26648,N_28918);
or UO_2750 (O_2750,N_27434,N_25330);
or UO_2751 (O_2751,N_27644,N_27426);
xor UO_2752 (O_2752,N_29619,N_28184);
or UO_2753 (O_2753,N_28407,N_28607);
nand UO_2754 (O_2754,N_25781,N_27826);
or UO_2755 (O_2755,N_25418,N_26400);
and UO_2756 (O_2756,N_25837,N_25825);
nor UO_2757 (O_2757,N_26689,N_29932);
or UO_2758 (O_2758,N_27684,N_29624);
or UO_2759 (O_2759,N_28858,N_28616);
nor UO_2760 (O_2760,N_25526,N_29139);
nand UO_2761 (O_2761,N_26852,N_27007);
and UO_2762 (O_2762,N_29016,N_28531);
or UO_2763 (O_2763,N_25584,N_27080);
or UO_2764 (O_2764,N_25026,N_27280);
or UO_2765 (O_2765,N_25307,N_29537);
xor UO_2766 (O_2766,N_27773,N_29346);
xor UO_2767 (O_2767,N_27600,N_26592);
and UO_2768 (O_2768,N_28410,N_26515);
and UO_2769 (O_2769,N_25862,N_25846);
and UO_2770 (O_2770,N_27818,N_25165);
or UO_2771 (O_2771,N_28188,N_25718);
nor UO_2772 (O_2772,N_26187,N_27806);
and UO_2773 (O_2773,N_25993,N_25602);
and UO_2774 (O_2774,N_28171,N_29837);
xor UO_2775 (O_2775,N_26187,N_26403);
or UO_2776 (O_2776,N_29743,N_29128);
or UO_2777 (O_2777,N_27785,N_25752);
nor UO_2778 (O_2778,N_25943,N_25939);
and UO_2779 (O_2779,N_27769,N_25170);
nor UO_2780 (O_2780,N_27350,N_25515);
and UO_2781 (O_2781,N_27249,N_29020);
nand UO_2782 (O_2782,N_28166,N_27708);
xor UO_2783 (O_2783,N_25470,N_29349);
nor UO_2784 (O_2784,N_25706,N_28901);
and UO_2785 (O_2785,N_28916,N_29499);
nand UO_2786 (O_2786,N_27671,N_28984);
or UO_2787 (O_2787,N_26880,N_26838);
or UO_2788 (O_2788,N_26602,N_25809);
nor UO_2789 (O_2789,N_27307,N_29422);
or UO_2790 (O_2790,N_29697,N_25024);
xor UO_2791 (O_2791,N_26690,N_27809);
or UO_2792 (O_2792,N_27174,N_29000);
nor UO_2793 (O_2793,N_27743,N_29144);
or UO_2794 (O_2794,N_29260,N_27585);
or UO_2795 (O_2795,N_26879,N_27768);
xor UO_2796 (O_2796,N_28843,N_26923);
nand UO_2797 (O_2797,N_26012,N_25611);
xnor UO_2798 (O_2798,N_25559,N_27695);
nand UO_2799 (O_2799,N_29538,N_28905);
nand UO_2800 (O_2800,N_26483,N_25787);
nor UO_2801 (O_2801,N_29027,N_25679);
and UO_2802 (O_2802,N_25170,N_25735);
nor UO_2803 (O_2803,N_29832,N_27432);
xor UO_2804 (O_2804,N_25359,N_25075);
or UO_2805 (O_2805,N_27458,N_26527);
or UO_2806 (O_2806,N_26988,N_27593);
or UO_2807 (O_2807,N_27052,N_26421);
xnor UO_2808 (O_2808,N_28934,N_28408);
nor UO_2809 (O_2809,N_28252,N_29976);
and UO_2810 (O_2810,N_28561,N_28347);
nor UO_2811 (O_2811,N_28133,N_29656);
xor UO_2812 (O_2812,N_25042,N_29598);
and UO_2813 (O_2813,N_28690,N_27523);
or UO_2814 (O_2814,N_27456,N_27439);
and UO_2815 (O_2815,N_27664,N_27540);
or UO_2816 (O_2816,N_26858,N_25424);
and UO_2817 (O_2817,N_25824,N_26535);
nand UO_2818 (O_2818,N_28441,N_25416);
xnor UO_2819 (O_2819,N_27790,N_27306);
or UO_2820 (O_2820,N_26886,N_26853);
nand UO_2821 (O_2821,N_27697,N_25400);
nand UO_2822 (O_2822,N_25369,N_28721);
nor UO_2823 (O_2823,N_26812,N_29811);
or UO_2824 (O_2824,N_27345,N_29679);
xor UO_2825 (O_2825,N_25792,N_29025);
xnor UO_2826 (O_2826,N_27736,N_29748);
and UO_2827 (O_2827,N_27398,N_26780);
or UO_2828 (O_2828,N_27597,N_26696);
nor UO_2829 (O_2829,N_27141,N_27414);
and UO_2830 (O_2830,N_28806,N_27651);
xor UO_2831 (O_2831,N_27873,N_27975);
nor UO_2832 (O_2832,N_29296,N_27101);
or UO_2833 (O_2833,N_28655,N_27540);
and UO_2834 (O_2834,N_28266,N_26034);
or UO_2835 (O_2835,N_26564,N_29187);
or UO_2836 (O_2836,N_28263,N_28736);
nand UO_2837 (O_2837,N_27723,N_28372);
and UO_2838 (O_2838,N_26948,N_27192);
xnor UO_2839 (O_2839,N_28297,N_25005);
xor UO_2840 (O_2840,N_25066,N_28012);
or UO_2841 (O_2841,N_25494,N_25296);
nor UO_2842 (O_2842,N_25816,N_27900);
and UO_2843 (O_2843,N_28021,N_25128);
and UO_2844 (O_2844,N_28153,N_28370);
or UO_2845 (O_2845,N_29273,N_29206);
or UO_2846 (O_2846,N_29546,N_26569);
and UO_2847 (O_2847,N_26293,N_29663);
nor UO_2848 (O_2848,N_27980,N_28382);
xor UO_2849 (O_2849,N_25434,N_29859);
nor UO_2850 (O_2850,N_26518,N_25947);
and UO_2851 (O_2851,N_25353,N_26549);
and UO_2852 (O_2852,N_29556,N_27921);
xnor UO_2853 (O_2853,N_29047,N_25262);
xnor UO_2854 (O_2854,N_27139,N_28894);
nand UO_2855 (O_2855,N_29747,N_26570);
xnor UO_2856 (O_2856,N_26153,N_28200);
xor UO_2857 (O_2857,N_28374,N_25558);
nor UO_2858 (O_2858,N_28317,N_25070);
and UO_2859 (O_2859,N_27670,N_26082);
and UO_2860 (O_2860,N_28536,N_25367);
or UO_2861 (O_2861,N_27417,N_26565);
and UO_2862 (O_2862,N_25567,N_26173);
or UO_2863 (O_2863,N_25784,N_27781);
or UO_2864 (O_2864,N_25850,N_27945);
or UO_2865 (O_2865,N_27156,N_29692);
xnor UO_2866 (O_2866,N_29370,N_25017);
nand UO_2867 (O_2867,N_29664,N_27425);
or UO_2868 (O_2868,N_28668,N_27153);
xnor UO_2869 (O_2869,N_28757,N_29344);
and UO_2870 (O_2870,N_27380,N_25054);
nor UO_2871 (O_2871,N_25347,N_29776);
xor UO_2872 (O_2872,N_25355,N_26111);
nor UO_2873 (O_2873,N_28744,N_25616);
xnor UO_2874 (O_2874,N_27132,N_26473);
xor UO_2875 (O_2875,N_27453,N_25502);
nor UO_2876 (O_2876,N_27611,N_29969);
and UO_2877 (O_2877,N_26747,N_28951);
nand UO_2878 (O_2878,N_28043,N_26659);
nand UO_2879 (O_2879,N_25684,N_26733);
or UO_2880 (O_2880,N_25192,N_29048);
nor UO_2881 (O_2881,N_26185,N_25606);
or UO_2882 (O_2882,N_27464,N_27383);
xor UO_2883 (O_2883,N_27663,N_25608);
nand UO_2884 (O_2884,N_29260,N_27536);
or UO_2885 (O_2885,N_28992,N_25048);
nand UO_2886 (O_2886,N_26285,N_28394);
and UO_2887 (O_2887,N_28384,N_25506);
xnor UO_2888 (O_2888,N_28683,N_25132);
xnor UO_2889 (O_2889,N_27747,N_26488);
and UO_2890 (O_2890,N_28143,N_27895);
or UO_2891 (O_2891,N_28108,N_25205);
and UO_2892 (O_2892,N_29735,N_26426);
and UO_2893 (O_2893,N_25563,N_29703);
nand UO_2894 (O_2894,N_28601,N_25233);
and UO_2895 (O_2895,N_27701,N_29580);
and UO_2896 (O_2896,N_29520,N_29398);
and UO_2897 (O_2897,N_28776,N_29910);
and UO_2898 (O_2898,N_26397,N_28350);
nor UO_2899 (O_2899,N_27050,N_28193);
and UO_2900 (O_2900,N_25144,N_28873);
nor UO_2901 (O_2901,N_26433,N_26114);
and UO_2902 (O_2902,N_27904,N_29544);
xor UO_2903 (O_2903,N_26939,N_25496);
and UO_2904 (O_2904,N_27508,N_25416);
nor UO_2905 (O_2905,N_29710,N_28835);
nor UO_2906 (O_2906,N_26314,N_26739);
or UO_2907 (O_2907,N_25155,N_28147);
xor UO_2908 (O_2908,N_25019,N_29041);
and UO_2909 (O_2909,N_26327,N_28121);
and UO_2910 (O_2910,N_28740,N_26335);
nor UO_2911 (O_2911,N_28732,N_26552);
xor UO_2912 (O_2912,N_29681,N_29138);
or UO_2913 (O_2913,N_29533,N_27424);
nor UO_2914 (O_2914,N_25162,N_29800);
and UO_2915 (O_2915,N_27163,N_29636);
and UO_2916 (O_2916,N_25522,N_27883);
or UO_2917 (O_2917,N_28997,N_29277);
nand UO_2918 (O_2918,N_28691,N_27161);
xnor UO_2919 (O_2919,N_28287,N_26974);
nor UO_2920 (O_2920,N_29219,N_27778);
xnor UO_2921 (O_2921,N_28244,N_25316);
and UO_2922 (O_2922,N_25022,N_29566);
and UO_2923 (O_2923,N_28478,N_29013);
xnor UO_2924 (O_2924,N_26530,N_27795);
nand UO_2925 (O_2925,N_25935,N_28269);
xor UO_2926 (O_2926,N_26256,N_27669);
and UO_2927 (O_2927,N_28187,N_28579);
xnor UO_2928 (O_2928,N_27328,N_25618);
or UO_2929 (O_2929,N_29011,N_25159);
and UO_2930 (O_2930,N_25715,N_29929);
and UO_2931 (O_2931,N_29241,N_29181);
and UO_2932 (O_2932,N_29083,N_28127);
nor UO_2933 (O_2933,N_25877,N_28842);
or UO_2934 (O_2934,N_27468,N_29855);
nor UO_2935 (O_2935,N_27543,N_25403);
nor UO_2936 (O_2936,N_26536,N_28210);
and UO_2937 (O_2937,N_25077,N_26946);
nand UO_2938 (O_2938,N_26689,N_27413);
nand UO_2939 (O_2939,N_26961,N_29697);
and UO_2940 (O_2940,N_29895,N_29225);
xnor UO_2941 (O_2941,N_28129,N_25718);
xnor UO_2942 (O_2942,N_29747,N_29476);
nand UO_2943 (O_2943,N_26284,N_28587);
nor UO_2944 (O_2944,N_25162,N_26038);
xnor UO_2945 (O_2945,N_29731,N_26459);
xor UO_2946 (O_2946,N_28338,N_28890);
or UO_2947 (O_2947,N_27473,N_26805);
xor UO_2948 (O_2948,N_27052,N_28186);
and UO_2949 (O_2949,N_25884,N_26122);
or UO_2950 (O_2950,N_28083,N_28640);
or UO_2951 (O_2951,N_27947,N_25845);
or UO_2952 (O_2952,N_26389,N_26851);
or UO_2953 (O_2953,N_28960,N_26395);
xnor UO_2954 (O_2954,N_25423,N_29987);
nand UO_2955 (O_2955,N_25402,N_25508);
nand UO_2956 (O_2956,N_26551,N_27787);
nand UO_2957 (O_2957,N_28085,N_27675);
and UO_2958 (O_2958,N_29373,N_25063);
nor UO_2959 (O_2959,N_29499,N_29395);
and UO_2960 (O_2960,N_29614,N_25016);
and UO_2961 (O_2961,N_25532,N_25638);
nand UO_2962 (O_2962,N_28005,N_27177);
or UO_2963 (O_2963,N_27434,N_25798);
nand UO_2964 (O_2964,N_27571,N_29212);
nor UO_2965 (O_2965,N_26614,N_29831);
xnor UO_2966 (O_2966,N_29496,N_28903);
nand UO_2967 (O_2967,N_28306,N_27377);
and UO_2968 (O_2968,N_28491,N_25295);
or UO_2969 (O_2969,N_25766,N_28572);
or UO_2970 (O_2970,N_29534,N_29649);
nand UO_2971 (O_2971,N_28400,N_28768);
nand UO_2972 (O_2972,N_28938,N_27338);
and UO_2973 (O_2973,N_25488,N_28736);
xnor UO_2974 (O_2974,N_26584,N_27324);
nand UO_2975 (O_2975,N_26158,N_29138);
or UO_2976 (O_2976,N_27771,N_29175);
and UO_2977 (O_2977,N_28368,N_25207);
and UO_2978 (O_2978,N_29011,N_29695);
nor UO_2979 (O_2979,N_29489,N_25176);
and UO_2980 (O_2980,N_26268,N_27733);
and UO_2981 (O_2981,N_28725,N_28483);
nor UO_2982 (O_2982,N_28468,N_25283);
xor UO_2983 (O_2983,N_25734,N_26654);
or UO_2984 (O_2984,N_28494,N_29966);
and UO_2985 (O_2985,N_27313,N_29912);
xor UO_2986 (O_2986,N_27182,N_25315);
or UO_2987 (O_2987,N_26368,N_27508);
and UO_2988 (O_2988,N_28105,N_29677);
and UO_2989 (O_2989,N_25139,N_29055);
or UO_2990 (O_2990,N_28849,N_27683);
nor UO_2991 (O_2991,N_28534,N_26188);
nor UO_2992 (O_2992,N_29298,N_26937);
and UO_2993 (O_2993,N_25202,N_29994);
xor UO_2994 (O_2994,N_25747,N_29247);
nand UO_2995 (O_2995,N_29690,N_26483);
xor UO_2996 (O_2996,N_27934,N_27312);
nor UO_2997 (O_2997,N_25524,N_25828);
nor UO_2998 (O_2998,N_29566,N_27709);
and UO_2999 (O_2999,N_28235,N_26526);
nand UO_3000 (O_3000,N_27206,N_27427);
xnor UO_3001 (O_3001,N_25286,N_27761);
nor UO_3002 (O_3002,N_27029,N_25493);
nor UO_3003 (O_3003,N_27521,N_29103);
xor UO_3004 (O_3004,N_29072,N_29025);
or UO_3005 (O_3005,N_29242,N_29880);
nand UO_3006 (O_3006,N_25948,N_27889);
xor UO_3007 (O_3007,N_28355,N_25666);
nor UO_3008 (O_3008,N_25095,N_29988);
nor UO_3009 (O_3009,N_29379,N_26334);
or UO_3010 (O_3010,N_28584,N_29761);
and UO_3011 (O_3011,N_26987,N_26891);
nand UO_3012 (O_3012,N_27095,N_26280);
or UO_3013 (O_3013,N_29145,N_28254);
nor UO_3014 (O_3014,N_28066,N_26722);
or UO_3015 (O_3015,N_29597,N_25046);
or UO_3016 (O_3016,N_25417,N_26675);
xnor UO_3017 (O_3017,N_28567,N_25714);
nor UO_3018 (O_3018,N_25499,N_29874);
nand UO_3019 (O_3019,N_26188,N_25476);
and UO_3020 (O_3020,N_27627,N_28302);
and UO_3021 (O_3021,N_27426,N_25759);
nand UO_3022 (O_3022,N_27308,N_27708);
nor UO_3023 (O_3023,N_27040,N_29760);
or UO_3024 (O_3024,N_27566,N_27848);
nand UO_3025 (O_3025,N_29590,N_28207);
nand UO_3026 (O_3026,N_25447,N_25512);
or UO_3027 (O_3027,N_25859,N_29493);
or UO_3028 (O_3028,N_25372,N_25898);
xor UO_3029 (O_3029,N_29483,N_26301);
and UO_3030 (O_3030,N_27239,N_27759);
or UO_3031 (O_3031,N_27729,N_29765);
nor UO_3032 (O_3032,N_25878,N_27877);
nor UO_3033 (O_3033,N_27155,N_25095);
xor UO_3034 (O_3034,N_28831,N_25971);
nor UO_3035 (O_3035,N_28566,N_29137);
or UO_3036 (O_3036,N_28352,N_29682);
nand UO_3037 (O_3037,N_25679,N_25434);
or UO_3038 (O_3038,N_27254,N_26763);
and UO_3039 (O_3039,N_25732,N_27011);
nand UO_3040 (O_3040,N_28871,N_26777);
or UO_3041 (O_3041,N_26854,N_27029);
xnor UO_3042 (O_3042,N_27091,N_26454);
nor UO_3043 (O_3043,N_27786,N_26106);
and UO_3044 (O_3044,N_25032,N_29383);
xnor UO_3045 (O_3045,N_29833,N_26645);
nor UO_3046 (O_3046,N_28951,N_26626);
nor UO_3047 (O_3047,N_27713,N_29045);
xnor UO_3048 (O_3048,N_25212,N_27395);
nand UO_3049 (O_3049,N_28911,N_28737);
nand UO_3050 (O_3050,N_26614,N_27309);
nor UO_3051 (O_3051,N_27194,N_25883);
xnor UO_3052 (O_3052,N_27790,N_25678);
or UO_3053 (O_3053,N_28261,N_26719);
nor UO_3054 (O_3054,N_25600,N_27451);
nand UO_3055 (O_3055,N_27250,N_25246);
or UO_3056 (O_3056,N_28609,N_26762);
nand UO_3057 (O_3057,N_26359,N_28311);
nand UO_3058 (O_3058,N_27880,N_29724);
or UO_3059 (O_3059,N_29431,N_27328);
xnor UO_3060 (O_3060,N_27479,N_29272);
nor UO_3061 (O_3061,N_26345,N_28991);
nor UO_3062 (O_3062,N_28653,N_25364);
and UO_3063 (O_3063,N_28918,N_25630);
and UO_3064 (O_3064,N_25558,N_27325);
nor UO_3065 (O_3065,N_28686,N_26507);
and UO_3066 (O_3066,N_25150,N_26220);
or UO_3067 (O_3067,N_26262,N_27807);
nand UO_3068 (O_3068,N_28382,N_27253);
and UO_3069 (O_3069,N_26011,N_29195);
and UO_3070 (O_3070,N_26133,N_26358);
and UO_3071 (O_3071,N_29700,N_28608);
nor UO_3072 (O_3072,N_29204,N_29627);
xnor UO_3073 (O_3073,N_25424,N_28061);
and UO_3074 (O_3074,N_29116,N_27340);
and UO_3075 (O_3075,N_27993,N_29509);
nand UO_3076 (O_3076,N_27438,N_27412);
nand UO_3077 (O_3077,N_27255,N_29717);
xnor UO_3078 (O_3078,N_26404,N_28182);
xnor UO_3079 (O_3079,N_26951,N_27755);
nand UO_3080 (O_3080,N_26815,N_25263);
and UO_3081 (O_3081,N_29512,N_28163);
or UO_3082 (O_3082,N_26732,N_28855);
or UO_3083 (O_3083,N_26705,N_26014);
nor UO_3084 (O_3084,N_27735,N_27461);
or UO_3085 (O_3085,N_28579,N_28765);
or UO_3086 (O_3086,N_29578,N_29533);
xnor UO_3087 (O_3087,N_26478,N_26221);
nand UO_3088 (O_3088,N_26105,N_25641);
xnor UO_3089 (O_3089,N_26610,N_28029);
and UO_3090 (O_3090,N_29721,N_27656);
nand UO_3091 (O_3091,N_29299,N_25544);
nor UO_3092 (O_3092,N_28644,N_27485);
nand UO_3093 (O_3093,N_28751,N_28441);
nor UO_3094 (O_3094,N_28695,N_26423);
nor UO_3095 (O_3095,N_28384,N_29553);
nor UO_3096 (O_3096,N_26307,N_26700);
xnor UO_3097 (O_3097,N_28791,N_27422);
and UO_3098 (O_3098,N_26706,N_25407);
or UO_3099 (O_3099,N_27699,N_26416);
nor UO_3100 (O_3100,N_25048,N_25569);
and UO_3101 (O_3101,N_25184,N_29411);
xor UO_3102 (O_3102,N_26028,N_25244);
or UO_3103 (O_3103,N_25392,N_26989);
or UO_3104 (O_3104,N_29127,N_25569);
and UO_3105 (O_3105,N_28941,N_25324);
xnor UO_3106 (O_3106,N_26262,N_28748);
nand UO_3107 (O_3107,N_26101,N_27340);
nand UO_3108 (O_3108,N_25470,N_25112);
xnor UO_3109 (O_3109,N_27855,N_28236);
xor UO_3110 (O_3110,N_27559,N_28070);
and UO_3111 (O_3111,N_28772,N_28372);
or UO_3112 (O_3112,N_25152,N_27603);
xor UO_3113 (O_3113,N_28897,N_25085);
xor UO_3114 (O_3114,N_26641,N_25177);
and UO_3115 (O_3115,N_28276,N_27441);
or UO_3116 (O_3116,N_26947,N_28310);
nor UO_3117 (O_3117,N_29810,N_26443);
or UO_3118 (O_3118,N_25716,N_26582);
nand UO_3119 (O_3119,N_25302,N_25468);
or UO_3120 (O_3120,N_27748,N_26715);
nand UO_3121 (O_3121,N_25244,N_26033);
or UO_3122 (O_3122,N_25482,N_25020);
xor UO_3123 (O_3123,N_27369,N_25915);
and UO_3124 (O_3124,N_28626,N_28137);
xnor UO_3125 (O_3125,N_25799,N_25660);
nand UO_3126 (O_3126,N_29116,N_26514);
nand UO_3127 (O_3127,N_26794,N_26540);
xnor UO_3128 (O_3128,N_25368,N_25182);
or UO_3129 (O_3129,N_29924,N_27467);
and UO_3130 (O_3130,N_29310,N_29795);
xnor UO_3131 (O_3131,N_27404,N_29661);
xnor UO_3132 (O_3132,N_25216,N_29449);
or UO_3133 (O_3133,N_29128,N_26946);
or UO_3134 (O_3134,N_29518,N_27531);
nand UO_3135 (O_3135,N_27599,N_25746);
and UO_3136 (O_3136,N_26026,N_27671);
xor UO_3137 (O_3137,N_27752,N_26242);
nor UO_3138 (O_3138,N_25565,N_25766);
or UO_3139 (O_3139,N_25663,N_29498);
or UO_3140 (O_3140,N_25480,N_25087);
and UO_3141 (O_3141,N_26398,N_29387);
xnor UO_3142 (O_3142,N_25199,N_27053);
nor UO_3143 (O_3143,N_29659,N_25568);
nand UO_3144 (O_3144,N_25440,N_29490);
or UO_3145 (O_3145,N_26599,N_25091);
nand UO_3146 (O_3146,N_28846,N_26875);
nand UO_3147 (O_3147,N_26198,N_25058);
nor UO_3148 (O_3148,N_26476,N_27466);
nand UO_3149 (O_3149,N_29845,N_29658);
xor UO_3150 (O_3150,N_25008,N_25574);
xor UO_3151 (O_3151,N_28034,N_25195);
and UO_3152 (O_3152,N_25290,N_25110);
nand UO_3153 (O_3153,N_26500,N_27947);
and UO_3154 (O_3154,N_25015,N_29859);
or UO_3155 (O_3155,N_26047,N_27671);
nor UO_3156 (O_3156,N_28348,N_27550);
or UO_3157 (O_3157,N_26322,N_26800);
xnor UO_3158 (O_3158,N_25633,N_28712);
xnor UO_3159 (O_3159,N_26980,N_28576);
or UO_3160 (O_3160,N_28360,N_29217);
nand UO_3161 (O_3161,N_28444,N_26082);
nand UO_3162 (O_3162,N_27462,N_25593);
and UO_3163 (O_3163,N_27076,N_29568);
nor UO_3164 (O_3164,N_28984,N_25994);
or UO_3165 (O_3165,N_27556,N_27240);
or UO_3166 (O_3166,N_28768,N_27279);
nand UO_3167 (O_3167,N_26571,N_25995);
and UO_3168 (O_3168,N_28749,N_27177);
and UO_3169 (O_3169,N_28602,N_27487);
and UO_3170 (O_3170,N_26161,N_25912);
nor UO_3171 (O_3171,N_27707,N_25098);
nand UO_3172 (O_3172,N_26985,N_25321);
nor UO_3173 (O_3173,N_29297,N_28175);
and UO_3174 (O_3174,N_25103,N_27889);
or UO_3175 (O_3175,N_26072,N_26018);
or UO_3176 (O_3176,N_28600,N_27827);
nor UO_3177 (O_3177,N_25198,N_28627);
or UO_3178 (O_3178,N_26391,N_28720);
nand UO_3179 (O_3179,N_26433,N_25851);
xor UO_3180 (O_3180,N_26599,N_29761);
nand UO_3181 (O_3181,N_27635,N_26112);
nand UO_3182 (O_3182,N_25107,N_29201);
or UO_3183 (O_3183,N_29372,N_25193);
nor UO_3184 (O_3184,N_29619,N_28298);
nor UO_3185 (O_3185,N_25464,N_27434);
nand UO_3186 (O_3186,N_29034,N_25182);
xnor UO_3187 (O_3187,N_26259,N_27358);
xor UO_3188 (O_3188,N_26838,N_27121);
xnor UO_3189 (O_3189,N_26402,N_25467);
nor UO_3190 (O_3190,N_28148,N_27893);
and UO_3191 (O_3191,N_27745,N_28063);
nand UO_3192 (O_3192,N_29588,N_26292);
and UO_3193 (O_3193,N_29731,N_25898);
xnor UO_3194 (O_3194,N_29194,N_28857);
or UO_3195 (O_3195,N_26140,N_29980);
nor UO_3196 (O_3196,N_28122,N_27735);
nand UO_3197 (O_3197,N_25287,N_25361);
or UO_3198 (O_3198,N_27806,N_28957);
xor UO_3199 (O_3199,N_25604,N_29019);
nor UO_3200 (O_3200,N_25927,N_29408);
nor UO_3201 (O_3201,N_25643,N_28841);
nand UO_3202 (O_3202,N_29023,N_29386);
xor UO_3203 (O_3203,N_29155,N_29685);
nand UO_3204 (O_3204,N_27444,N_27023);
xnor UO_3205 (O_3205,N_27316,N_26126);
and UO_3206 (O_3206,N_26448,N_28050);
or UO_3207 (O_3207,N_27725,N_29888);
xnor UO_3208 (O_3208,N_28253,N_26448);
nand UO_3209 (O_3209,N_27293,N_25251);
and UO_3210 (O_3210,N_27956,N_29936);
nor UO_3211 (O_3211,N_25073,N_25288);
or UO_3212 (O_3212,N_27051,N_28380);
nor UO_3213 (O_3213,N_28109,N_25443);
or UO_3214 (O_3214,N_26275,N_28303);
xor UO_3215 (O_3215,N_26608,N_28321);
xnor UO_3216 (O_3216,N_27939,N_29377);
nand UO_3217 (O_3217,N_28667,N_26836);
nand UO_3218 (O_3218,N_27808,N_26381);
xnor UO_3219 (O_3219,N_25114,N_25311);
xor UO_3220 (O_3220,N_25310,N_27405);
nor UO_3221 (O_3221,N_28229,N_25606);
nor UO_3222 (O_3222,N_29583,N_28980);
or UO_3223 (O_3223,N_27545,N_25264);
nand UO_3224 (O_3224,N_25761,N_28737);
xor UO_3225 (O_3225,N_25096,N_28645);
xor UO_3226 (O_3226,N_28023,N_29639);
xor UO_3227 (O_3227,N_25648,N_26904);
or UO_3228 (O_3228,N_28050,N_25248);
or UO_3229 (O_3229,N_28190,N_27150);
and UO_3230 (O_3230,N_25421,N_29096);
or UO_3231 (O_3231,N_27251,N_27985);
nor UO_3232 (O_3232,N_29485,N_26380);
xor UO_3233 (O_3233,N_25476,N_29431);
xor UO_3234 (O_3234,N_27540,N_28530);
nor UO_3235 (O_3235,N_26355,N_27571);
xor UO_3236 (O_3236,N_27978,N_27939);
xor UO_3237 (O_3237,N_29809,N_25877);
or UO_3238 (O_3238,N_28177,N_29697);
and UO_3239 (O_3239,N_28363,N_25131);
or UO_3240 (O_3240,N_28773,N_29660);
nor UO_3241 (O_3241,N_26755,N_26685);
or UO_3242 (O_3242,N_28337,N_26927);
or UO_3243 (O_3243,N_28841,N_27029);
nand UO_3244 (O_3244,N_28079,N_28906);
or UO_3245 (O_3245,N_25018,N_28630);
or UO_3246 (O_3246,N_27530,N_25404);
xnor UO_3247 (O_3247,N_25916,N_27272);
and UO_3248 (O_3248,N_26033,N_29582);
nand UO_3249 (O_3249,N_26070,N_27379);
nor UO_3250 (O_3250,N_29383,N_27777);
xnor UO_3251 (O_3251,N_29447,N_26860);
xor UO_3252 (O_3252,N_27270,N_25228);
and UO_3253 (O_3253,N_27826,N_27865);
nor UO_3254 (O_3254,N_25419,N_27049);
nand UO_3255 (O_3255,N_27198,N_29628);
nor UO_3256 (O_3256,N_26906,N_25171);
nand UO_3257 (O_3257,N_28985,N_28631);
and UO_3258 (O_3258,N_27770,N_26912);
or UO_3259 (O_3259,N_26356,N_26649);
nand UO_3260 (O_3260,N_26718,N_29400);
or UO_3261 (O_3261,N_26195,N_29975);
and UO_3262 (O_3262,N_27093,N_25962);
xor UO_3263 (O_3263,N_28316,N_29129);
xor UO_3264 (O_3264,N_25530,N_29044);
or UO_3265 (O_3265,N_26444,N_27242);
nand UO_3266 (O_3266,N_29324,N_27987);
and UO_3267 (O_3267,N_28974,N_26065);
xor UO_3268 (O_3268,N_27241,N_28638);
and UO_3269 (O_3269,N_28187,N_26307);
or UO_3270 (O_3270,N_26093,N_29162);
and UO_3271 (O_3271,N_26011,N_25898);
and UO_3272 (O_3272,N_28924,N_26177);
and UO_3273 (O_3273,N_26955,N_25172);
or UO_3274 (O_3274,N_29709,N_29025);
nor UO_3275 (O_3275,N_28446,N_25837);
xnor UO_3276 (O_3276,N_27368,N_25705);
nor UO_3277 (O_3277,N_29690,N_27094);
or UO_3278 (O_3278,N_28232,N_28337);
xor UO_3279 (O_3279,N_25894,N_28996);
nand UO_3280 (O_3280,N_27584,N_29707);
xnor UO_3281 (O_3281,N_27583,N_27183);
xor UO_3282 (O_3282,N_26560,N_25146);
or UO_3283 (O_3283,N_25683,N_27947);
nand UO_3284 (O_3284,N_28035,N_25248);
nor UO_3285 (O_3285,N_27768,N_25895);
nand UO_3286 (O_3286,N_25647,N_29945);
xnor UO_3287 (O_3287,N_28801,N_28128);
nor UO_3288 (O_3288,N_29726,N_28691);
and UO_3289 (O_3289,N_26702,N_27954);
or UO_3290 (O_3290,N_28945,N_28791);
nand UO_3291 (O_3291,N_29950,N_29144);
nand UO_3292 (O_3292,N_25867,N_29800);
and UO_3293 (O_3293,N_25495,N_25984);
nand UO_3294 (O_3294,N_27187,N_25902);
and UO_3295 (O_3295,N_27162,N_28075);
and UO_3296 (O_3296,N_28490,N_27790);
and UO_3297 (O_3297,N_28223,N_25250);
nor UO_3298 (O_3298,N_29998,N_25420);
nand UO_3299 (O_3299,N_29566,N_29917);
or UO_3300 (O_3300,N_25458,N_28909);
xor UO_3301 (O_3301,N_29987,N_28206);
and UO_3302 (O_3302,N_27425,N_27279);
nor UO_3303 (O_3303,N_26688,N_26991);
and UO_3304 (O_3304,N_29200,N_25378);
and UO_3305 (O_3305,N_26969,N_29732);
nor UO_3306 (O_3306,N_25502,N_25518);
nand UO_3307 (O_3307,N_27397,N_26555);
nor UO_3308 (O_3308,N_25461,N_27662);
nor UO_3309 (O_3309,N_29296,N_25677);
nor UO_3310 (O_3310,N_25805,N_29500);
nand UO_3311 (O_3311,N_29804,N_28284);
and UO_3312 (O_3312,N_28368,N_25076);
and UO_3313 (O_3313,N_25224,N_28810);
nor UO_3314 (O_3314,N_29110,N_26484);
nand UO_3315 (O_3315,N_25857,N_26569);
or UO_3316 (O_3316,N_28926,N_28714);
and UO_3317 (O_3317,N_27339,N_28952);
nor UO_3318 (O_3318,N_29168,N_25016);
nor UO_3319 (O_3319,N_29951,N_27883);
nand UO_3320 (O_3320,N_28503,N_29452);
or UO_3321 (O_3321,N_28620,N_25757);
xnor UO_3322 (O_3322,N_29111,N_26538);
nor UO_3323 (O_3323,N_27080,N_29737);
and UO_3324 (O_3324,N_27578,N_27202);
nor UO_3325 (O_3325,N_29584,N_26252);
and UO_3326 (O_3326,N_27083,N_29536);
or UO_3327 (O_3327,N_27255,N_26269);
nand UO_3328 (O_3328,N_27540,N_27517);
or UO_3329 (O_3329,N_29622,N_27240);
xor UO_3330 (O_3330,N_25770,N_26747);
and UO_3331 (O_3331,N_26578,N_29985);
or UO_3332 (O_3332,N_26827,N_25356);
or UO_3333 (O_3333,N_25396,N_25767);
nand UO_3334 (O_3334,N_26085,N_29588);
nor UO_3335 (O_3335,N_25061,N_28076);
nor UO_3336 (O_3336,N_28573,N_29160);
nand UO_3337 (O_3337,N_27202,N_29543);
nand UO_3338 (O_3338,N_27655,N_28415);
nand UO_3339 (O_3339,N_25063,N_29454);
or UO_3340 (O_3340,N_26594,N_28995);
and UO_3341 (O_3341,N_27709,N_28146);
and UO_3342 (O_3342,N_27813,N_29334);
nor UO_3343 (O_3343,N_28193,N_25659);
and UO_3344 (O_3344,N_26141,N_26061);
and UO_3345 (O_3345,N_28744,N_29560);
and UO_3346 (O_3346,N_26510,N_28737);
xnor UO_3347 (O_3347,N_27078,N_27124);
nand UO_3348 (O_3348,N_28092,N_26091);
xnor UO_3349 (O_3349,N_27009,N_25569);
or UO_3350 (O_3350,N_29880,N_28213);
and UO_3351 (O_3351,N_27005,N_29953);
and UO_3352 (O_3352,N_29286,N_27301);
or UO_3353 (O_3353,N_26137,N_28304);
nand UO_3354 (O_3354,N_27254,N_26551);
nor UO_3355 (O_3355,N_26344,N_25654);
and UO_3356 (O_3356,N_29269,N_26395);
and UO_3357 (O_3357,N_25986,N_25552);
xor UO_3358 (O_3358,N_25600,N_28568);
xnor UO_3359 (O_3359,N_26125,N_28153);
xor UO_3360 (O_3360,N_26418,N_27329);
and UO_3361 (O_3361,N_27536,N_29247);
nand UO_3362 (O_3362,N_27918,N_27446);
nand UO_3363 (O_3363,N_28662,N_27990);
nor UO_3364 (O_3364,N_26339,N_28383);
or UO_3365 (O_3365,N_27435,N_27654);
and UO_3366 (O_3366,N_26486,N_29739);
nor UO_3367 (O_3367,N_25441,N_27855);
and UO_3368 (O_3368,N_29297,N_25472);
nand UO_3369 (O_3369,N_26514,N_25257);
nor UO_3370 (O_3370,N_26721,N_25375);
or UO_3371 (O_3371,N_28464,N_29267);
nand UO_3372 (O_3372,N_29637,N_25171);
and UO_3373 (O_3373,N_27572,N_28274);
nor UO_3374 (O_3374,N_27356,N_25982);
or UO_3375 (O_3375,N_29157,N_26321);
or UO_3376 (O_3376,N_27528,N_25815);
or UO_3377 (O_3377,N_28912,N_25124);
nor UO_3378 (O_3378,N_29296,N_25059);
nor UO_3379 (O_3379,N_28396,N_26988);
nand UO_3380 (O_3380,N_28543,N_28551);
nor UO_3381 (O_3381,N_27518,N_28411);
nor UO_3382 (O_3382,N_25783,N_28351);
nor UO_3383 (O_3383,N_28838,N_27904);
or UO_3384 (O_3384,N_26617,N_28784);
nand UO_3385 (O_3385,N_29967,N_26616);
xor UO_3386 (O_3386,N_26075,N_28552);
nor UO_3387 (O_3387,N_27076,N_25399);
nor UO_3388 (O_3388,N_25104,N_29756);
and UO_3389 (O_3389,N_25850,N_29132);
and UO_3390 (O_3390,N_25181,N_27020);
nand UO_3391 (O_3391,N_29671,N_29200);
and UO_3392 (O_3392,N_28250,N_27504);
xor UO_3393 (O_3393,N_29820,N_28931);
xor UO_3394 (O_3394,N_27910,N_28847);
xor UO_3395 (O_3395,N_29758,N_28953);
xor UO_3396 (O_3396,N_25433,N_26145);
or UO_3397 (O_3397,N_25233,N_28678);
nor UO_3398 (O_3398,N_25780,N_27860);
nor UO_3399 (O_3399,N_26003,N_26240);
nor UO_3400 (O_3400,N_29167,N_27436);
nor UO_3401 (O_3401,N_26359,N_28770);
nor UO_3402 (O_3402,N_28696,N_27607);
nand UO_3403 (O_3403,N_27620,N_26977);
or UO_3404 (O_3404,N_26211,N_29514);
and UO_3405 (O_3405,N_28840,N_25557);
xor UO_3406 (O_3406,N_28356,N_25449);
xor UO_3407 (O_3407,N_29642,N_25913);
nand UO_3408 (O_3408,N_25952,N_27829);
xnor UO_3409 (O_3409,N_25387,N_27277);
nor UO_3410 (O_3410,N_28998,N_25669);
or UO_3411 (O_3411,N_28455,N_25998);
nor UO_3412 (O_3412,N_29923,N_28035);
nor UO_3413 (O_3413,N_25907,N_26338);
and UO_3414 (O_3414,N_29061,N_26265);
or UO_3415 (O_3415,N_25623,N_28970);
nor UO_3416 (O_3416,N_27636,N_26628);
nand UO_3417 (O_3417,N_29287,N_29685);
nand UO_3418 (O_3418,N_27292,N_25439);
xnor UO_3419 (O_3419,N_29401,N_25728);
nand UO_3420 (O_3420,N_25775,N_26646);
xor UO_3421 (O_3421,N_29632,N_25683);
and UO_3422 (O_3422,N_25038,N_29325);
and UO_3423 (O_3423,N_26622,N_26694);
xnor UO_3424 (O_3424,N_26942,N_29145);
nor UO_3425 (O_3425,N_29491,N_26082);
or UO_3426 (O_3426,N_29726,N_25286);
xor UO_3427 (O_3427,N_27237,N_27515);
nand UO_3428 (O_3428,N_25806,N_28730);
or UO_3429 (O_3429,N_25813,N_29679);
or UO_3430 (O_3430,N_28463,N_26269);
xor UO_3431 (O_3431,N_28092,N_27016);
xnor UO_3432 (O_3432,N_29229,N_29022);
or UO_3433 (O_3433,N_27937,N_28169);
or UO_3434 (O_3434,N_25138,N_27226);
or UO_3435 (O_3435,N_25488,N_27572);
and UO_3436 (O_3436,N_29976,N_26086);
nor UO_3437 (O_3437,N_29701,N_27455);
nor UO_3438 (O_3438,N_25711,N_26546);
and UO_3439 (O_3439,N_28571,N_26168);
or UO_3440 (O_3440,N_28740,N_28562);
xnor UO_3441 (O_3441,N_29903,N_25578);
nor UO_3442 (O_3442,N_25773,N_26336);
and UO_3443 (O_3443,N_27037,N_26951);
xor UO_3444 (O_3444,N_25368,N_27432);
xnor UO_3445 (O_3445,N_25967,N_27588);
nor UO_3446 (O_3446,N_28957,N_27194);
xnor UO_3447 (O_3447,N_29794,N_28105);
nand UO_3448 (O_3448,N_27515,N_27959);
nor UO_3449 (O_3449,N_25043,N_28066);
nor UO_3450 (O_3450,N_26633,N_29488);
xor UO_3451 (O_3451,N_28100,N_26681);
xor UO_3452 (O_3452,N_29561,N_27244);
nand UO_3453 (O_3453,N_26367,N_27581);
nand UO_3454 (O_3454,N_27574,N_25050);
nor UO_3455 (O_3455,N_26568,N_26761);
nand UO_3456 (O_3456,N_27719,N_29030);
or UO_3457 (O_3457,N_28427,N_29810);
nand UO_3458 (O_3458,N_27672,N_29900);
and UO_3459 (O_3459,N_26437,N_25088);
and UO_3460 (O_3460,N_27318,N_27904);
or UO_3461 (O_3461,N_26914,N_28165);
and UO_3462 (O_3462,N_25232,N_25351);
or UO_3463 (O_3463,N_27747,N_28354);
nor UO_3464 (O_3464,N_26791,N_27629);
or UO_3465 (O_3465,N_28809,N_29289);
nor UO_3466 (O_3466,N_29936,N_26155);
and UO_3467 (O_3467,N_29992,N_28477);
or UO_3468 (O_3468,N_27922,N_28698);
or UO_3469 (O_3469,N_29080,N_28116);
nand UO_3470 (O_3470,N_26294,N_29144);
nor UO_3471 (O_3471,N_26510,N_26129);
xor UO_3472 (O_3472,N_26296,N_29462);
xor UO_3473 (O_3473,N_29688,N_26841);
nand UO_3474 (O_3474,N_25284,N_28253);
nor UO_3475 (O_3475,N_25053,N_25514);
xor UO_3476 (O_3476,N_25841,N_25269);
and UO_3477 (O_3477,N_29609,N_27795);
nor UO_3478 (O_3478,N_26641,N_26586);
nand UO_3479 (O_3479,N_27914,N_25875);
xnor UO_3480 (O_3480,N_25677,N_29095);
nor UO_3481 (O_3481,N_27728,N_27365);
and UO_3482 (O_3482,N_26126,N_27480);
nor UO_3483 (O_3483,N_27054,N_25038);
nand UO_3484 (O_3484,N_25500,N_27822);
nor UO_3485 (O_3485,N_25113,N_26630);
nand UO_3486 (O_3486,N_27267,N_28993);
xor UO_3487 (O_3487,N_28195,N_25789);
nor UO_3488 (O_3488,N_25139,N_25126);
nor UO_3489 (O_3489,N_29442,N_29873);
nor UO_3490 (O_3490,N_29614,N_27564);
nor UO_3491 (O_3491,N_27188,N_29545);
nand UO_3492 (O_3492,N_28425,N_25985);
or UO_3493 (O_3493,N_27592,N_29891);
and UO_3494 (O_3494,N_28996,N_29062);
and UO_3495 (O_3495,N_29290,N_25357);
nor UO_3496 (O_3496,N_25510,N_26313);
or UO_3497 (O_3497,N_25142,N_27347);
or UO_3498 (O_3498,N_29800,N_27656);
nand UO_3499 (O_3499,N_28784,N_29531);
endmodule