module basic_500_3000_500_5_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_3,In_211);
and U1 (N_1,In_282,In_415);
nand U2 (N_2,In_223,In_274);
nor U3 (N_3,In_479,In_158);
nand U4 (N_4,In_459,In_498);
xnor U5 (N_5,In_252,In_388);
or U6 (N_6,In_412,In_447);
nand U7 (N_7,In_35,In_324);
xnor U8 (N_8,In_221,In_393);
and U9 (N_9,In_308,In_234);
xor U10 (N_10,In_164,In_244);
xor U11 (N_11,In_454,In_178);
or U12 (N_12,In_475,In_362);
or U13 (N_13,In_105,In_203);
nand U14 (N_14,In_314,In_61);
xor U15 (N_15,In_92,In_167);
nand U16 (N_16,In_48,In_251);
and U17 (N_17,In_477,In_346);
nand U18 (N_18,In_494,In_46);
nor U19 (N_19,In_224,In_204);
nand U20 (N_20,In_127,In_411);
nand U21 (N_21,In_33,In_267);
nand U22 (N_22,In_481,In_330);
xnor U23 (N_23,In_396,In_209);
and U24 (N_24,In_117,In_166);
nand U25 (N_25,In_446,In_76);
nand U26 (N_26,In_163,In_339);
nor U27 (N_27,In_94,In_275);
nand U28 (N_28,In_417,In_305);
nor U29 (N_29,In_291,In_56);
nand U30 (N_30,In_325,In_80);
and U31 (N_31,In_302,In_90);
nor U32 (N_32,In_287,In_156);
xor U33 (N_33,In_6,In_122);
nand U34 (N_34,In_180,In_23);
or U35 (N_35,In_217,In_67);
or U36 (N_36,In_320,In_458);
xnor U37 (N_37,In_216,In_248);
and U38 (N_38,In_378,In_496);
nand U39 (N_39,In_148,In_371);
nand U40 (N_40,In_181,In_311);
nor U41 (N_41,In_108,In_34);
nand U42 (N_42,In_38,In_7);
nor U43 (N_43,In_174,In_335);
nor U44 (N_44,In_161,In_289);
xnor U45 (N_45,In_124,In_199);
nand U46 (N_46,In_97,In_243);
nand U47 (N_47,In_52,In_309);
nor U48 (N_48,In_408,In_256);
nand U49 (N_49,In_183,In_318);
and U50 (N_50,In_194,In_231);
and U51 (N_51,In_352,In_421);
nand U52 (N_52,In_64,In_344);
nand U53 (N_53,In_192,In_294);
or U54 (N_54,In_208,In_160);
xnor U55 (N_55,In_402,In_228);
nor U56 (N_56,In_196,In_136);
or U57 (N_57,In_22,In_72);
or U58 (N_58,In_100,In_345);
nand U59 (N_59,In_395,In_301);
nor U60 (N_60,In_106,In_467);
or U61 (N_61,In_60,In_2);
or U62 (N_62,In_188,In_202);
and U63 (N_63,In_1,In_348);
xnor U64 (N_64,In_20,In_226);
nand U65 (N_65,In_31,In_112);
nor U66 (N_66,In_426,In_230);
xor U67 (N_67,In_384,In_409);
xnor U68 (N_68,In_43,In_261);
or U69 (N_69,In_336,In_0);
or U70 (N_70,In_403,In_142);
xor U71 (N_71,In_75,In_65);
or U72 (N_72,In_141,In_214);
nand U73 (N_73,In_441,In_103);
nand U74 (N_74,In_281,In_394);
nand U75 (N_75,In_438,In_413);
nand U76 (N_76,In_427,In_176);
nand U77 (N_77,In_16,In_307);
or U78 (N_78,In_120,In_169);
xnor U79 (N_79,In_277,In_316);
nor U80 (N_80,In_349,In_292);
nor U81 (N_81,In_375,In_385);
and U82 (N_82,In_470,In_74);
or U83 (N_83,In_66,In_58);
nor U84 (N_84,In_215,In_300);
nor U85 (N_85,In_165,In_280);
xor U86 (N_86,In_63,In_337);
and U87 (N_87,In_342,In_357);
nor U88 (N_88,In_478,In_14);
nor U89 (N_89,In_153,In_206);
and U90 (N_90,In_240,In_400);
nor U91 (N_91,In_455,In_207);
nor U92 (N_92,In_284,In_430);
and U93 (N_93,In_259,In_482);
xor U94 (N_94,In_488,In_113);
nand U95 (N_95,In_460,In_489);
nand U96 (N_96,In_5,In_55);
nand U97 (N_97,In_205,In_419);
nand U98 (N_98,In_270,In_98);
nand U99 (N_99,In_383,In_431);
or U100 (N_100,In_404,In_326);
xor U101 (N_101,In_29,In_463);
nand U102 (N_102,In_130,In_382);
and U103 (N_103,In_238,In_129);
xor U104 (N_104,In_125,In_295);
and U105 (N_105,In_49,In_179);
or U106 (N_106,In_30,In_442);
nor U107 (N_107,In_422,In_297);
nor U108 (N_108,In_88,In_424);
nor U109 (N_109,In_343,In_476);
or U110 (N_110,In_116,In_239);
nor U111 (N_111,In_182,In_247);
nand U112 (N_112,In_77,In_36);
nand U113 (N_113,In_323,In_304);
nand U114 (N_114,In_134,In_45);
nand U115 (N_115,In_145,In_131);
or U116 (N_116,In_351,In_109);
and U117 (N_117,In_364,In_186);
xor U118 (N_118,In_229,In_397);
nand U119 (N_119,In_47,In_59);
nor U120 (N_120,In_128,In_12);
nand U121 (N_121,In_474,In_296);
nand U122 (N_122,In_51,In_95);
or U123 (N_123,In_185,In_99);
xnor U124 (N_124,In_456,In_450);
xnor U125 (N_125,In_200,In_245);
xnor U126 (N_126,In_269,In_487);
or U127 (N_127,In_233,In_448);
or U128 (N_128,In_386,In_170);
nor U129 (N_129,In_84,In_439);
nor U130 (N_130,In_437,In_468);
xor U131 (N_131,In_480,In_387);
nor U132 (N_132,In_187,In_283);
nand U133 (N_133,In_15,In_273);
nor U134 (N_134,In_132,In_25);
nand U135 (N_135,In_338,In_418);
xnor U136 (N_136,In_11,In_490);
or U137 (N_137,In_327,In_368);
or U138 (N_138,In_451,In_78);
or U139 (N_139,In_360,In_86);
xnor U140 (N_140,In_333,In_288);
nor U141 (N_141,In_341,In_389);
nand U142 (N_142,In_365,In_62);
nor U143 (N_143,In_328,In_361);
or U144 (N_144,In_443,In_126);
nand U145 (N_145,In_253,In_401);
xor U146 (N_146,In_276,In_81);
or U147 (N_147,In_114,In_249);
nand U148 (N_148,In_453,In_57);
and U149 (N_149,In_260,In_173);
nor U150 (N_150,In_315,In_286);
nor U151 (N_151,In_266,In_429);
nand U152 (N_152,In_306,In_71);
and U153 (N_153,In_50,In_104);
nand U154 (N_154,In_213,In_440);
nor U155 (N_155,In_299,In_171);
nor U156 (N_156,In_332,In_313);
nor U157 (N_157,In_189,In_17);
xor U158 (N_158,In_150,In_497);
and U159 (N_159,In_172,In_82);
nand U160 (N_160,In_310,In_359);
xor U161 (N_161,In_8,In_26);
nor U162 (N_162,In_374,In_492);
nand U163 (N_163,In_380,In_491);
xor U164 (N_164,In_9,In_19);
xor U165 (N_165,In_197,In_40);
xor U166 (N_166,In_373,In_83);
or U167 (N_167,In_369,In_139);
nand U168 (N_168,In_322,In_366);
nor U169 (N_169,In_390,In_18);
and U170 (N_170,In_191,In_235);
nor U171 (N_171,In_119,In_246);
nand U172 (N_172,In_363,In_133);
nor U173 (N_173,In_184,In_219);
nor U174 (N_174,In_499,In_398);
xor U175 (N_175,In_87,In_268);
and U176 (N_176,In_358,In_70);
and U177 (N_177,In_111,In_272);
xnor U178 (N_178,In_483,In_312);
and U179 (N_179,In_271,In_159);
nand U180 (N_180,In_212,In_484);
or U181 (N_181,In_262,In_89);
and U182 (N_182,In_118,In_255);
nor U183 (N_183,In_279,In_392);
nand U184 (N_184,In_465,In_329);
and U185 (N_185,In_405,In_28);
and U186 (N_186,In_190,In_293);
or U187 (N_187,In_140,In_298);
and U188 (N_188,In_68,In_376);
nand U189 (N_189,In_347,In_218);
or U190 (N_190,In_420,In_263);
nor U191 (N_191,In_466,In_321);
and U192 (N_192,In_39,In_101);
nor U193 (N_193,In_250,In_462);
nor U194 (N_194,In_472,In_121);
or U195 (N_195,In_391,In_242);
nor U196 (N_196,In_152,In_73);
nand U197 (N_197,In_435,In_254);
and U198 (N_198,In_222,In_69);
xnor U199 (N_199,In_41,In_154);
or U200 (N_200,In_53,In_37);
nand U201 (N_201,In_227,In_85);
and U202 (N_202,In_428,In_96);
or U203 (N_203,In_157,In_471);
or U204 (N_204,In_210,In_461);
nor U205 (N_205,In_265,In_13);
or U206 (N_206,In_79,In_457);
and U207 (N_207,In_464,In_93);
nand U208 (N_208,In_155,In_372);
or U209 (N_209,In_473,In_290);
or U210 (N_210,In_317,In_399);
nor U211 (N_211,In_423,In_162);
and U212 (N_212,In_367,In_485);
xor U213 (N_213,In_54,In_264);
and U214 (N_214,In_198,In_407);
nand U215 (N_215,In_377,In_445);
nor U216 (N_216,In_355,In_370);
nand U217 (N_217,In_433,In_319);
nand U218 (N_218,In_278,In_143);
or U219 (N_219,In_138,In_110);
or U220 (N_220,In_432,In_237);
xor U221 (N_221,In_285,In_353);
nand U222 (N_222,In_469,In_425);
and U223 (N_223,In_144,In_436);
or U224 (N_224,In_452,In_303);
nor U225 (N_225,In_241,In_24);
and U226 (N_226,In_168,In_175);
nor U227 (N_227,In_414,In_10);
and U228 (N_228,In_444,In_379);
nand U229 (N_229,In_449,In_410);
nand U230 (N_230,In_123,In_334);
and U231 (N_231,In_4,In_193);
nor U232 (N_232,In_258,In_149);
and U233 (N_233,In_495,In_220);
nand U234 (N_234,In_416,In_381);
or U235 (N_235,In_42,In_493);
nand U236 (N_236,In_225,In_236);
or U237 (N_237,In_356,In_406);
xor U238 (N_238,In_107,In_151);
nor U239 (N_239,In_257,In_21);
and U240 (N_240,In_486,In_102);
nor U241 (N_241,In_32,In_331);
nor U242 (N_242,In_340,In_177);
nor U243 (N_243,In_146,In_147);
nand U244 (N_244,In_354,In_27);
xnor U245 (N_245,In_44,In_115);
nor U246 (N_246,In_135,In_201);
nand U247 (N_247,In_232,In_195);
or U248 (N_248,In_350,In_137);
nor U249 (N_249,In_91,In_434);
xnor U250 (N_250,In_28,In_118);
and U251 (N_251,In_40,In_143);
and U252 (N_252,In_302,In_262);
and U253 (N_253,In_361,In_484);
nand U254 (N_254,In_176,In_301);
nor U255 (N_255,In_481,In_439);
xor U256 (N_256,In_325,In_142);
and U257 (N_257,In_438,In_279);
nor U258 (N_258,In_378,In_241);
nor U259 (N_259,In_344,In_309);
nor U260 (N_260,In_167,In_300);
or U261 (N_261,In_382,In_161);
or U262 (N_262,In_404,In_1);
xnor U263 (N_263,In_144,In_37);
and U264 (N_264,In_201,In_160);
and U265 (N_265,In_27,In_316);
nand U266 (N_266,In_331,In_110);
nor U267 (N_267,In_418,In_64);
and U268 (N_268,In_45,In_319);
or U269 (N_269,In_93,In_394);
xnor U270 (N_270,In_100,In_55);
xnor U271 (N_271,In_401,In_422);
nand U272 (N_272,In_462,In_179);
and U273 (N_273,In_450,In_245);
nor U274 (N_274,In_169,In_411);
or U275 (N_275,In_495,In_31);
nor U276 (N_276,In_258,In_423);
and U277 (N_277,In_17,In_377);
nand U278 (N_278,In_63,In_364);
and U279 (N_279,In_452,In_104);
nand U280 (N_280,In_314,In_92);
xnor U281 (N_281,In_307,In_174);
or U282 (N_282,In_251,In_183);
and U283 (N_283,In_69,In_401);
xnor U284 (N_284,In_77,In_283);
and U285 (N_285,In_359,In_319);
xor U286 (N_286,In_3,In_449);
nand U287 (N_287,In_187,In_104);
nand U288 (N_288,In_244,In_119);
and U289 (N_289,In_105,In_411);
nand U290 (N_290,In_374,In_262);
and U291 (N_291,In_321,In_48);
and U292 (N_292,In_440,In_241);
nor U293 (N_293,In_219,In_297);
xnor U294 (N_294,In_439,In_187);
and U295 (N_295,In_249,In_482);
nor U296 (N_296,In_246,In_443);
nor U297 (N_297,In_135,In_409);
nand U298 (N_298,In_207,In_389);
xor U299 (N_299,In_316,In_14);
or U300 (N_300,In_168,In_71);
xor U301 (N_301,In_483,In_100);
and U302 (N_302,In_313,In_427);
nor U303 (N_303,In_368,In_293);
nand U304 (N_304,In_258,In_473);
nor U305 (N_305,In_301,In_177);
nor U306 (N_306,In_174,In_224);
or U307 (N_307,In_83,In_190);
or U308 (N_308,In_190,In_194);
nand U309 (N_309,In_495,In_482);
or U310 (N_310,In_169,In_109);
nor U311 (N_311,In_22,In_297);
xor U312 (N_312,In_352,In_417);
nor U313 (N_313,In_485,In_396);
and U314 (N_314,In_492,In_144);
or U315 (N_315,In_447,In_442);
or U316 (N_316,In_44,In_186);
nor U317 (N_317,In_169,In_66);
or U318 (N_318,In_310,In_284);
nand U319 (N_319,In_488,In_438);
nand U320 (N_320,In_15,In_12);
xnor U321 (N_321,In_400,In_217);
and U322 (N_322,In_85,In_258);
nor U323 (N_323,In_292,In_120);
or U324 (N_324,In_237,In_114);
and U325 (N_325,In_46,In_170);
and U326 (N_326,In_356,In_269);
or U327 (N_327,In_214,In_393);
nand U328 (N_328,In_189,In_396);
xnor U329 (N_329,In_96,In_304);
or U330 (N_330,In_478,In_217);
or U331 (N_331,In_304,In_106);
nand U332 (N_332,In_145,In_340);
nand U333 (N_333,In_406,In_265);
xor U334 (N_334,In_447,In_300);
nor U335 (N_335,In_368,In_349);
xnor U336 (N_336,In_483,In_272);
or U337 (N_337,In_192,In_30);
nor U338 (N_338,In_410,In_349);
and U339 (N_339,In_283,In_345);
xor U340 (N_340,In_88,In_63);
nand U341 (N_341,In_472,In_119);
nand U342 (N_342,In_460,In_343);
or U343 (N_343,In_231,In_361);
or U344 (N_344,In_218,In_288);
nand U345 (N_345,In_488,In_128);
xor U346 (N_346,In_316,In_190);
xnor U347 (N_347,In_32,In_466);
or U348 (N_348,In_185,In_434);
and U349 (N_349,In_289,In_125);
or U350 (N_350,In_332,In_495);
nor U351 (N_351,In_476,In_380);
nand U352 (N_352,In_163,In_409);
and U353 (N_353,In_306,In_301);
or U354 (N_354,In_63,In_248);
or U355 (N_355,In_488,In_440);
xor U356 (N_356,In_342,In_300);
nor U357 (N_357,In_368,In_344);
nand U358 (N_358,In_341,In_106);
nor U359 (N_359,In_137,In_24);
or U360 (N_360,In_23,In_252);
and U361 (N_361,In_218,In_31);
xor U362 (N_362,In_217,In_63);
and U363 (N_363,In_356,In_54);
and U364 (N_364,In_146,In_474);
nand U365 (N_365,In_237,In_297);
xnor U366 (N_366,In_407,In_13);
nand U367 (N_367,In_81,In_105);
nor U368 (N_368,In_160,In_430);
xnor U369 (N_369,In_143,In_32);
nor U370 (N_370,In_102,In_148);
xnor U371 (N_371,In_208,In_57);
or U372 (N_372,In_220,In_371);
xnor U373 (N_373,In_108,In_271);
xor U374 (N_374,In_134,In_343);
xnor U375 (N_375,In_145,In_256);
nor U376 (N_376,In_136,In_63);
xnor U377 (N_377,In_63,In_321);
and U378 (N_378,In_404,In_388);
or U379 (N_379,In_336,In_366);
nand U380 (N_380,In_469,In_125);
and U381 (N_381,In_136,In_19);
or U382 (N_382,In_202,In_232);
nor U383 (N_383,In_465,In_275);
nand U384 (N_384,In_421,In_167);
and U385 (N_385,In_247,In_238);
and U386 (N_386,In_235,In_395);
xnor U387 (N_387,In_276,In_426);
and U388 (N_388,In_286,In_73);
nand U389 (N_389,In_105,In_60);
xnor U390 (N_390,In_339,In_449);
and U391 (N_391,In_425,In_314);
xnor U392 (N_392,In_260,In_292);
nor U393 (N_393,In_49,In_135);
or U394 (N_394,In_154,In_187);
nor U395 (N_395,In_15,In_279);
nor U396 (N_396,In_417,In_326);
nor U397 (N_397,In_28,In_44);
or U398 (N_398,In_347,In_55);
nor U399 (N_399,In_373,In_104);
or U400 (N_400,In_55,In_461);
or U401 (N_401,In_323,In_242);
or U402 (N_402,In_475,In_244);
nand U403 (N_403,In_335,In_1);
xor U404 (N_404,In_497,In_185);
nor U405 (N_405,In_318,In_457);
nor U406 (N_406,In_186,In_258);
nand U407 (N_407,In_343,In_213);
or U408 (N_408,In_275,In_123);
and U409 (N_409,In_473,In_53);
xor U410 (N_410,In_236,In_214);
and U411 (N_411,In_362,In_27);
xnor U412 (N_412,In_373,In_432);
nor U413 (N_413,In_470,In_168);
nand U414 (N_414,In_313,In_341);
and U415 (N_415,In_262,In_125);
or U416 (N_416,In_262,In_203);
or U417 (N_417,In_401,In_443);
and U418 (N_418,In_84,In_327);
and U419 (N_419,In_471,In_393);
or U420 (N_420,In_310,In_0);
or U421 (N_421,In_130,In_420);
nand U422 (N_422,In_250,In_325);
xor U423 (N_423,In_121,In_338);
nand U424 (N_424,In_469,In_384);
xnor U425 (N_425,In_76,In_262);
and U426 (N_426,In_351,In_390);
nand U427 (N_427,In_130,In_191);
and U428 (N_428,In_153,In_410);
and U429 (N_429,In_480,In_435);
nor U430 (N_430,In_220,In_496);
nor U431 (N_431,In_488,In_60);
nand U432 (N_432,In_266,In_411);
or U433 (N_433,In_408,In_479);
nor U434 (N_434,In_442,In_332);
xor U435 (N_435,In_163,In_482);
nor U436 (N_436,In_210,In_272);
nor U437 (N_437,In_205,In_338);
xor U438 (N_438,In_54,In_496);
or U439 (N_439,In_260,In_25);
nand U440 (N_440,In_29,In_293);
and U441 (N_441,In_7,In_423);
nor U442 (N_442,In_251,In_115);
or U443 (N_443,In_420,In_68);
or U444 (N_444,In_327,In_259);
nand U445 (N_445,In_160,In_240);
and U446 (N_446,In_492,In_319);
nor U447 (N_447,In_353,In_151);
and U448 (N_448,In_122,In_34);
nand U449 (N_449,In_342,In_388);
nand U450 (N_450,In_489,In_292);
or U451 (N_451,In_66,In_30);
or U452 (N_452,In_167,In_133);
nor U453 (N_453,In_216,In_116);
or U454 (N_454,In_325,In_95);
or U455 (N_455,In_383,In_427);
xnor U456 (N_456,In_243,In_254);
nor U457 (N_457,In_73,In_266);
and U458 (N_458,In_34,In_179);
nor U459 (N_459,In_484,In_290);
xor U460 (N_460,In_253,In_470);
nor U461 (N_461,In_124,In_205);
and U462 (N_462,In_492,In_242);
nand U463 (N_463,In_50,In_108);
nand U464 (N_464,In_195,In_351);
or U465 (N_465,In_13,In_226);
xor U466 (N_466,In_237,In_350);
nand U467 (N_467,In_81,In_20);
and U468 (N_468,In_270,In_7);
nand U469 (N_469,In_322,In_214);
nor U470 (N_470,In_252,In_155);
nor U471 (N_471,In_163,In_207);
xor U472 (N_472,In_366,In_5);
or U473 (N_473,In_31,In_392);
nand U474 (N_474,In_200,In_145);
nor U475 (N_475,In_253,In_187);
nor U476 (N_476,In_84,In_421);
or U477 (N_477,In_182,In_123);
and U478 (N_478,In_151,In_204);
and U479 (N_479,In_327,In_161);
xnor U480 (N_480,In_120,In_382);
or U481 (N_481,In_247,In_324);
nand U482 (N_482,In_208,In_92);
and U483 (N_483,In_35,In_122);
and U484 (N_484,In_149,In_371);
nor U485 (N_485,In_124,In_413);
nor U486 (N_486,In_116,In_40);
nor U487 (N_487,In_134,In_196);
and U488 (N_488,In_463,In_155);
nand U489 (N_489,In_141,In_455);
nor U490 (N_490,In_345,In_148);
and U491 (N_491,In_14,In_277);
and U492 (N_492,In_303,In_436);
xor U493 (N_493,In_365,In_103);
nand U494 (N_494,In_104,In_73);
or U495 (N_495,In_409,In_96);
and U496 (N_496,In_173,In_14);
nand U497 (N_497,In_324,In_356);
or U498 (N_498,In_167,In_86);
nand U499 (N_499,In_66,In_451);
or U500 (N_500,In_480,In_332);
xor U501 (N_501,In_222,In_419);
nand U502 (N_502,In_261,In_83);
and U503 (N_503,In_383,In_432);
xnor U504 (N_504,In_98,In_164);
nand U505 (N_505,In_197,In_223);
nor U506 (N_506,In_391,In_145);
nand U507 (N_507,In_438,In_464);
nor U508 (N_508,In_80,In_157);
or U509 (N_509,In_253,In_4);
nor U510 (N_510,In_460,In_203);
xnor U511 (N_511,In_423,In_47);
xnor U512 (N_512,In_101,In_475);
and U513 (N_513,In_287,In_419);
nand U514 (N_514,In_233,In_20);
xnor U515 (N_515,In_309,In_253);
or U516 (N_516,In_65,In_277);
nand U517 (N_517,In_392,In_52);
or U518 (N_518,In_229,In_251);
nand U519 (N_519,In_178,In_194);
nand U520 (N_520,In_96,In_206);
nor U521 (N_521,In_55,In_400);
and U522 (N_522,In_13,In_203);
nand U523 (N_523,In_204,In_394);
or U524 (N_524,In_465,In_78);
and U525 (N_525,In_143,In_185);
nand U526 (N_526,In_63,In_353);
and U527 (N_527,In_422,In_229);
or U528 (N_528,In_332,In_404);
nor U529 (N_529,In_427,In_460);
and U530 (N_530,In_410,In_159);
nor U531 (N_531,In_474,In_291);
and U532 (N_532,In_96,In_242);
nor U533 (N_533,In_46,In_204);
nand U534 (N_534,In_276,In_225);
xnor U535 (N_535,In_298,In_485);
xnor U536 (N_536,In_375,In_320);
nand U537 (N_537,In_65,In_16);
nand U538 (N_538,In_469,In_120);
and U539 (N_539,In_490,In_379);
nand U540 (N_540,In_29,In_441);
or U541 (N_541,In_130,In_367);
nor U542 (N_542,In_240,In_388);
or U543 (N_543,In_255,In_220);
nor U544 (N_544,In_477,In_196);
nor U545 (N_545,In_205,In_188);
or U546 (N_546,In_112,In_117);
and U547 (N_547,In_248,In_60);
nand U548 (N_548,In_486,In_180);
nand U549 (N_549,In_26,In_252);
xnor U550 (N_550,In_150,In_377);
and U551 (N_551,In_356,In_464);
xor U552 (N_552,In_355,In_53);
nor U553 (N_553,In_399,In_377);
xnor U554 (N_554,In_467,In_322);
and U555 (N_555,In_96,In_478);
and U556 (N_556,In_470,In_98);
or U557 (N_557,In_192,In_416);
and U558 (N_558,In_13,In_482);
and U559 (N_559,In_302,In_363);
and U560 (N_560,In_269,In_33);
xor U561 (N_561,In_231,In_322);
nor U562 (N_562,In_189,In_348);
or U563 (N_563,In_319,In_282);
xor U564 (N_564,In_93,In_158);
or U565 (N_565,In_154,In_226);
xnor U566 (N_566,In_183,In_289);
nor U567 (N_567,In_418,In_354);
nand U568 (N_568,In_380,In_490);
nand U569 (N_569,In_444,In_335);
nor U570 (N_570,In_350,In_467);
xnor U571 (N_571,In_96,In_197);
or U572 (N_572,In_404,In_284);
or U573 (N_573,In_293,In_463);
and U574 (N_574,In_420,In_368);
xnor U575 (N_575,In_283,In_420);
nand U576 (N_576,In_236,In_448);
or U577 (N_577,In_14,In_139);
or U578 (N_578,In_62,In_236);
nand U579 (N_579,In_284,In_55);
nand U580 (N_580,In_178,In_160);
and U581 (N_581,In_19,In_118);
and U582 (N_582,In_147,In_160);
nand U583 (N_583,In_248,In_416);
and U584 (N_584,In_144,In_272);
nand U585 (N_585,In_145,In_63);
and U586 (N_586,In_322,In_396);
or U587 (N_587,In_207,In_321);
or U588 (N_588,In_301,In_404);
nor U589 (N_589,In_104,In_86);
nor U590 (N_590,In_48,In_237);
xor U591 (N_591,In_128,In_106);
and U592 (N_592,In_22,In_312);
xnor U593 (N_593,In_382,In_165);
nand U594 (N_594,In_245,In_269);
and U595 (N_595,In_84,In_262);
or U596 (N_596,In_379,In_2);
or U597 (N_597,In_267,In_498);
or U598 (N_598,In_261,In_434);
and U599 (N_599,In_135,In_188);
nor U600 (N_600,N_568,N_262);
and U601 (N_601,N_193,N_274);
xnor U602 (N_602,N_153,N_225);
nand U603 (N_603,N_339,N_552);
or U604 (N_604,N_53,N_369);
and U605 (N_605,N_11,N_215);
and U606 (N_606,N_363,N_290);
and U607 (N_607,N_594,N_165);
nand U608 (N_608,N_146,N_522);
nand U609 (N_609,N_521,N_370);
nand U610 (N_610,N_387,N_134);
and U611 (N_611,N_212,N_122);
nor U612 (N_612,N_286,N_504);
nor U613 (N_613,N_404,N_580);
nor U614 (N_614,N_156,N_564);
and U615 (N_615,N_467,N_419);
nand U616 (N_616,N_551,N_358);
and U617 (N_617,N_338,N_344);
nand U618 (N_618,N_257,N_380);
nor U619 (N_619,N_571,N_410);
or U620 (N_620,N_538,N_301);
or U621 (N_621,N_559,N_195);
nor U622 (N_622,N_180,N_245);
nand U623 (N_623,N_174,N_459);
nor U624 (N_624,N_411,N_528);
or U625 (N_625,N_557,N_132);
nor U626 (N_626,N_461,N_261);
and U627 (N_627,N_545,N_445);
or U628 (N_628,N_343,N_373);
and U629 (N_629,N_575,N_412);
or U630 (N_630,N_359,N_396);
nand U631 (N_631,N_295,N_456);
nand U632 (N_632,N_263,N_120);
or U633 (N_633,N_392,N_105);
and U634 (N_634,N_171,N_535);
or U635 (N_635,N_511,N_474);
and U636 (N_636,N_138,N_320);
xor U637 (N_637,N_310,N_409);
nand U638 (N_638,N_251,N_349);
or U639 (N_639,N_469,N_94);
nor U640 (N_640,N_311,N_523);
or U641 (N_641,N_207,N_450);
xnor U642 (N_642,N_536,N_36);
xnor U643 (N_643,N_140,N_247);
xnor U644 (N_644,N_484,N_583);
nor U645 (N_645,N_141,N_435);
xor U646 (N_646,N_326,N_51);
nand U647 (N_647,N_509,N_208);
nor U648 (N_648,N_307,N_487);
nand U649 (N_649,N_576,N_391);
nor U650 (N_650,N_114,N_309);
xnor U651 (N_651,N_577,N_345);
and U652 (N_652,N_476,N_315);
and U653 (N_653,N_164,N_176);
nor U654 (N_654,N_33,N_240);
or U655 (N_655,N_151,N_73);
xnor U656 (N_656,N_490,N_25);
or U657 (N_657,N_477,N_492);
and U658 (N_658,N_252,N_88);
and U659 (N_659,N_3,N_330);
nor U660 (N_660,N_386,N_289);
xor U661 (N_661,N_353,N_434);
nand U662 (N_662,N_50,N_161);
or U663 (N_663,N_139,N_43);
xor U664 (N_664,N_590,N_187);
and U665 (N_665,N_26,N_52);
nor U666 (N_666,N_76,N_133);
and U667 (N_667,N_107,N_77);
nor U668 (N_668,N_220,N_287);
xor U669 (N_669,N_554,N_483);
nand U670 (N_670,N_291,N_230);
nand U671 (N_671,N_273,N_28);
nor U672 (N_672,N_70,N_425);
xor U673 (N_673,N_92,N_281);
nor U674 (N_674,N_599,N_259);
and U675 (N_675,N_123,N_341);
nand U676 (N_676,N_278,N_317);
nor U677 (N_677,N_78,N_238);
xnor U678 (N_678,N_178,N_405);
or U679 (N_679,N_335,N_495);
or U680 (N_680,N_464,N_532);
or U681 (N_681,N_424,N_206);
and U682 (N_682,N_546,N_596);
or U683 (N_683,N_398,N_471);
or U684 (N_684,N_480,N_444);
nand U685 (N_685,N_381,N_155);
nor U686 (N_686,N_525,N_201);
xnor U687 (N_687,N_457,N_473);
xnor U688 (N_688,N_248,N_427);
nor U689 (N_689,N_529,N_272);
and U690 (N_690,N_555,N_589);
xor U691 (N_691,N_573,N_403);
nor U692 (N_692,N_58,N_54);
or U693 (N_693,N_169,N_19);
nor U694 (N_694,N_585,N_159);
nor U695 (N_695,N_100,N_510);
xor U696 (N_696,N_16,N_109);
nor U697 (N_697,N_285,N_86);
nor U698 (N_698,N_519,N_270);
xnor U699 (N_699,N_482,N_130);
xnor U700 (N_700,N_18,N_539);
xor U701 (N_701,N_277,N_305);
xnor U702 (N_702,N_125,N_237);
and U703 (N_703,N_64,N_524);
nor U704 (N_704,N_574,N_17);
and U705 (N_705,N_232,N_362);
and U706 (N_706,N_60,N_160);
or U707 (N_707,N_421,N_79);
or U708 (N_708,N_269,N_390);
xnor U709 (N_709,N_560,N_31);
nand U710 (N_710,N_219,N_593);
nor U711 (N_711,N_111,N_550);
nand U712 (N_712,N_361,N_508);
and U713 (N_713,N_266,N_297);
nand U714 (N_714,N_163,N_246);
nand U715 (N_715,N_365,N_197);
nand U716 (N_716,N_177,N_222);
xor U717 (N_717,N_352,N_470);
nand U718 (N_718,N_556,N_260);
and U719 (N_719,N_158,N_84);
xnor U720 (N_720,N_194,N_55);
nand U721 (N_721,N_417,N_181);
xor U722 (N_722,N_85,N_385);
nand U723 (N_723,N_401,N_20);
xor U724 (N_724,N_384,N_302);
and U725 (N_725,N_436,N_292);
or U726 (N_726,N_318,N_265);
or U727 (N_727,N_209,N_357);
nor U728 (N_728,N_527,N_418);
nor U729 (N_729,N_399,N_451);
xnor U730 (N_730,N_96,N_414);
or U731 (N_731,N_14,N_595);
nand U732 (N_732,N_127,N_95);
nor U733 (N_733,N_440,N_598);
nor U734 (N_734,N_4,N_423);
or U735 (N_735,N_2,N_465);
nand U736 (N_736,N_558,N_377);
or U737 (N_737,N_347,N_67);
nor U738 (N_738,N_332,N_516);
nor U739 (N_739,N_323,N_101);
nand U740 (N_740,N_98,N_388);
nand U741 (N_741,N_400,N_253);
nand U742 (N_742,N_6,N_162);
nor U743 (N_743,N_561,N_42);
and U744 (N_744,N_513,N_533);
nor U745 (N_745,N_507,N_249);
nor U746 (N_746,N_23,N_542);
nor U747 (N_747,N_514,N_202);
nor U748 (N_748,N_588,N_62);
and U749 (N_749,N_38,N_144);
xnor U750 (N_750,N_422,N_548);
nor U751 (N_751,N_453,N_75);
nand U752 (N_752,N_89,N_441);
xnor U753 (N_753,N_40,N_366);
xor U754 (N_754,N_540,N_63);
and U755 (N_755,N_7,N_21);
and U756 (N_756,N_211,N_406);
xnor U757 (N_757,N_314,N_280);
nand U758 (N_758,N_231,N_526);
nand U759 (N_759,N_108,N_382);
xor U760 (N_760,N_41,N_397);
or U761 (N_761,N_129,N_44);
nor U762 (N_762,N_426,N_47);
and U763 (N_763,N_56,N_69);
and U764 (N_764,N_367,N_498);
xor U765 (N_765,N_446,N_110);
nand U766 (N_766,N_543,N_192);
and U767 (N_767,N_429,N_586);
or U768 (N_768,N_488,N_346);
nand U769 (N_769,N_515,N_175);
nor U770 (N_770,N_582,N_49);
xor U771 (N_771,N_503,N_226);
nand U772 (N_772,N_87,N_15);
xnor U773 (N_773,N_452,N_393);
and U774 (N_774,N_82,N_499);
nand U775 (N_775,N_472,N_170);
nor U776 (N_776,N_117,N_566);
nand U777 (N_777,N_184,N_152);
xnor U778 (N_778,N_126,N_199);
nand U779 (N_779,N_416,N_572);
and U780 (N_780,N_13,N_213);
and U781 (N_781,N_420,N_221);
and U782 (N_782,N_481,N_27);
nor U783 (N_783,N_534,N_433);
nand U784 (N_784,N_135,N_282);
xnor U785 (N_785,N_321,N_379);
xnor U786 (N_786,N_579,N_35);
xnor U787 (N_787,N_137,N_271);
xor U788 (N_788,N_506,N_549);
nor U789 (N_789,N_131,N_188);
xnor U790 (N_790,N_413,N_218);
and U791 (N_791,N_375,N_447);
nor U792 (N_792,N_570,N_167);
nor U793 (N_793,N_61,N_210);
nor U794 (N_794,N_355,N_83);
xnor U795 (N_795,N_22,N_115);
nand U796 (N_796,N_368,N_243);
nor U797 (N_797,N_402,N_242);
nand U798 (N_798,N_442,N_500);
nand U799 (N_799,N_319,N_5);
xor U800 (N_800,N_371,N_223);
and U801 (N_801,N_298,N_166);
or U802 (N_802,N_531,N_428);
nor U803 (N_803,N_342,N_333);
or U804 (N_804,N_196,N_97);
nand U805 (N_805,N_591,N_541);
or U806 (N_806,N_205,N_112);
xnor U807 (N_807,N_71,N_217);
nand U808 (N_808,N_157,N_430);
xnor U809 (N_809,N_374,N_66);
and U810 (N_810,N_408,N_173);
nand U811 (N_811,N_443,N_168);
nand U812 (N_812,N_48,N_306);
and U813 (N_813,N_239,N_597);
and U814 (N_814,N_494,N_113);
xnor U815 (N_815,N_454,N_284);
xor U816 (N_816,N_74,N_254);
or U817 (N_817,N_186,N_395);
xnor U818 (N_818,N_150,N_241);
and U819 (N_819,N_283,N_581);
or U820 (N_820,N_485,N_91);
xnor U821 (N_821,N_308,N_530);
or U822 (N_822,N_10,N_104);
or U823 (N_823,N_90,N_296);
nor U824 (N_824,N_93,N_275);
and U825 (N_825,N_475,N_147);
or U826 (N_826,N_32,N_148);
or U827 (N_827,N_154,N_518);
and U828 (N_828,N_293,N_479);
nor U829 (N_829,N_316,N_415);
and U830 (N_830,N_303,N_299);
nor U831 (N_831,N_118,N_276);
or U832 (N_832,N_149,N_1);
nand U833 (N_833,N_493,N_204);
or U834 (N_834,N_455,N_121);
nand U835 (N_835,N_200,N_565);
xor U836 (N_836,N_466,N_562);
nand U837 (N_837,N_29,N_360);
nand U838 (N_838,N_304,N_438);
and U839 (N_839,N_145,N_578);
nand U840 (N_840,N_517,N_431);
or U841 (N_841,N_128,N_136);
or U842 (N_842,N_119,N_57);
or U843 (N_843,N_224,N_45);
nand U844 (N_844,N_547,N_313);
nor U845 (N_845,N_234,N_235);
nor U846 (N_846,N_372,N_142);
or U847 (N_847,N_244,N_300);
nor U848 (N_848,N_389,N_68);
and U849 (N_849,N_106,N_183);
nand U850 (N_850,N_227,N_65);
nor U851 (N_851,N_331,N_185);
or U852 (N_852,N_279,N_103);
and U853 (N_853,N_288,N_460);
and U854 (N_854,N_364,N_255);
xor U855 (N_855,N_99,N_383);
or U856 (N_856,N_312,N_264);
or U857 (N_857,N_437,N_407);
and U858 (N_858,N_334,N_351);
nand U859 (N_859,N_350,N_563);
and U860 (N_860,N_143,N_256);
nand U861 (N_861,N_329,N_228);
or U862 (N_862,N_37,N_80);
xnor U863 (N_863,N_72,N_394);
nand U864 (N_864,N_432,N_322);
or U865 (N_865,N_268,N_267);
nor U866 (N_866,N_486,N_449);
or U867 (N_867,N_102,N_340);
nor U868 (N_868,N_489,N_81);
nand U869 (N_869,N_124,N_182);
nand U870 (N_870,N_376,N_501);
and U871 (N_871,N_229,N_236);
nand U872 (N_872,N_378,N_458);
nand U873 (N_873,N_584,N_328);
nand U874 (N_874,N_294,N_198);
nor U875 (N_875,N_569,N_325);
nor U876 (N_876,N_348,N_258);
nor U877 (N_877,N_491,N_172);
and U878 (N_878,N_191,N_9);
and U879 (N_879,N_30,N_354);
xor U880 (N_880,N_439,N_214);
or U881 (N_881,N_24,N_537);
or U882 (N_882,N_587,N_463);
xnor U883 (N_883,N_12,N_502);
and U884 (N_884,N_496,N_337);
or U885 (N_885,N_233,N_520);
xor U886 (N_886,N_512,N_189);
or U887 (N_887,N_203,N_59);
nand U888 (N_888,N_553,N_462);
nor U889 (N_889,N_336,N_216);
nand U890 (N_890,N_327,N_8);
nand U891 (N_891,N_0,N_497);
nor U892 (N_892,N_324,N_567);
and U893 (N_893,N_190,N_544);
or U894 (N_894,N_468,N_356);
nand U895 (N_895,N_116,N_39);
and U896 (N_896,N_34,N_250);
and U897 (N_897,N_448,N_478);
nand U898 (N_898,N_592,N_505);
and U899 (N_899,N_179,N_46);
nor U900 (N_900,N_56,N_14);
nor U901 (N_901,N_501,N_67);
nor U902 (N_902,N_446,N_290);
xor U903 (N_903,N_67,N_343);
nor U904 (N_904,N_372,N_508);
nand U905 (N_905,N_375,N_294);
xnor U906 (N_906,N_218,N_558);
nand U907 (N_907,N_88,N_471);
xor U908 (N_908,N_272,N_260);
nor U909 (N_909,N_348,N_127);
nand U910 (N_910,N_415,N_572);
nand U911 (N_911,N_582,N_34);
or U912 (N_912,N_61,N_244);
nor U913 (N_913,N_318,N_279);
or U914 (N_914,N_296,N_352);
nor U915 (N_915,N_98,N_333);
and U916 (N_916,N_54,N_177);
and U917 (N_917,N_26,N_54);
and U918 (N_918,N_344,N_496);
nand U919 (N_919,N_1,N_436);
xnor U920 (N_920,N_29,N_489);
nand U921 (N_921,N_499,N_361);
nand U922 (N_922,N_275,N_301);
xnor U923 (N_923,N_272,N_162);
xor U924 (N_924,N_311,N_213);
or U925 (N_925,N_287,N_90);
xnor U926 (N_926,N_534,N_372);
nor U927 (N_927,N_509,N_245);
or U928 (N_928,N_303,N_396);
xnor U929 (N_929,N_241,N_288);
or U930 (N_930,N_385,N_80);
or U931 (N_931,N_518,N_142);
and U932 (N_932,N_479,N_311);
or U933 (N_933,N_517,N_450);
xnor U934 (N_934,N_353,N_229);
nand U935 (N_935,N_325,N_468);
and U936 (N_936,N_524,N_313);
or U937 (N_937,N_61,N_323);
or U938 (N_938,N_436,N_576);
xnor U939 (N_939,N_217,N_38);
nor U940 (N_940,N_125,N_207);
xor U941 (N_941,N_594,N_303);
or U942 (N_942,N_535,N_0);
xnor U943 (N_943,N_212,N_175);
xor U944 (N_944,N_339,N_46);
or U945 (N_945,N_417,N_62);
nand U946 (N_946,N_29,N_140);
nand U947 (N_947,N_96,N_259);
nand U948 (N_948,N_437,N_479);
or U949 (N_949,N_571,N_110);
xnor U950 (N_950,N_293,N_462);
and U951 (N_951,N_17,N_154);
and U952 (N_952,N_530,N_426);
xor U953 (N_953,N_285,N_575);
xor U954 (N_954,N_573,N_331);
or U955 (N_955,N_203,N_79);
xnor U956 (N_956,N_420,N_10);
and U957 (N_957,N_96,N_399);
or U958 (N_958,N_28,N_190);
xnor U959 (N_959,N_521,N_322);
or U960 (N_960,N_54,N_66);
nor U961 (N_961,N_62,N_549);
xor U962 (N_962,N_159,N_140);
nand U963 (N_963,N_300,N_137);
xor U964 (N_964,N_286,N_333);
nor U965 (N_965,N_113,N_259);
nor U966 (N_966,N_146,N_277);
or U967 (N_967,N_227,N_121);
or U968 (N_968,N_562,N_271);
and U969 (N_969,N_423,N_267);
and U970 (N_970,N_392,N_324);
xor U971 (N_971,N_187,N_390);
nor U972 (N_972,N_213,N_573);
nand U973 (N_973,N_380,N_60);
xnor U974 (N_974,N_208,N_288);
nand U975 (N_975,N_549,N_56);
nand U976 (N_976,N_318,N_463);
nor U977 (N_977,N_259,N_440);
or U978 (N_978,N_163,N_390);
or U979 (N_979,N_173,N_192);
nor U980 (N_980,N_146,N_54);
nor U981 (N_981,N_478,N_217);
nand U982 (N_982,N_234,N_360);
nor U983 (N_983,N_266,N_111);
xor U984 (N_984,N_352,N_192);
xnor U985 (N_985,N_457,N_5);
xor U986 (N_986,N_327,N_232);
nor U987 (N_987,N_253,N_102);
or U988 (N_988,N_457,N_241);
and U989 (N_989,N_235,N_145);
or U990 (N_990,N_32,N_463);
nor U991 (N_991,N_455,N_340);
xor U992 (N_992,N_584,N_432);
xor U993 (N_993,N_228,N_218);
nor U994 (N_994,N_417,N_189);
nor U995 (N_995,N_17,N_29);
nor U996 (N_996,N_321,N_111);
or U997 (N_997,N_100,N_280);
xnor U998 (N_998,N_587,N_419);
xor U999 (N_999,N_76,N_445);
nand U1000 (N_1000,N_98,N_345);
nand U1001 (N_1001,N_443,N_394);
or U1002 (N_1002,N_28,N_120);
nor U1003 (N_1003,N_146,N_599);
nor U1004 (N_1004,N_308,N_265);
nand U1005 (N_1005,N_386,N_117);
and U1006 (N_1006,N_109,N_592);
nand U1007 (N_1007,N_265,N_33);
nand U1008 (N_1008,N_232,N_383);
and U1009 (N_1009,N_384,N_473);
and U1010 (N_1010,N_491,N_145);
or U1011 (N_1011,N_453,N_413);
nand U1012 (N_1012,N_564,N_195);
nand U1013 (N_1013,N_99,N_64);
xnor U1014 (N_1014,N_542,N_496);
or U1015 (N_1015,N_23,N_28);
or U1016 (N_1016,N_144,N_472);
or U1017 (N_1017,N_355,N_222);
nor U1018 (N_1018,N_98,N_463);
or U1019 (N_1019,N_224,N_46);
nand U1020 (N_1020,N_510,N_243);
or U1021 (N_1021,N_87,N_411);
xor U1022 (N_1022,N_287,N_588);
and U1023 (N_1023,N_593,N_206);
xor U1024 (N_1024,N_65,N_330);
and U1025 (N_1025,N_517,N_289);
and U1026 (N_1026,N_45,N_79);
and U1027 (N_1027,N_316,N_335);
or U1028 (N_1028,N_423,N_244);
or U1029 (N_1029,N_430,N_57);
and U1030 (N_1030,N_117,N_16);
nor U1031 (N_1031,N_132,N_471);
or U1032 (N_1032,N_187,N_338);
xnor U1033 (N_1033,N_453,N_467);
nand U1034 (N_1034,N_574,N_598);
nand U1035 (N_1035,N_335,N_191);
nor U1036 (N_1036,N_484,N_464);
nand U1037 (N_1037,N_369,N_47);
nor U1038 (N_1038,N_231,N_3);
or U1039 (N_1039,N_230,N_34);
or U1040 (N_1040,N_167,N_471);
and U1041 (N_1041,N_333,N_78);
xnor U1042 (N_1042,N_17,N_354);
or U1043 (N_1043,N_380,N_195);
nand U1044 (N_1044,N_3,N_186);
or U1045 (N_1045,N_49,N_261);
and U1046 (N_1046,N_131,N_392);
and U1047 (N_1047,N_244,N_331);
nor U1048 (N_1048,N_267,N_191);
xnor U1049 (N_1049,N_58,N_325);
and U1050 (N_1050,N_561,N_120);
nand U1051 (N_1051,N_412,N_385);
nand U1052 (N_1052,N_235,N_458);
or U1053 (N_1053,N_312,N_562);
or U1054 (N_1054,N_165,N_29);
or U1055 (N_1055,N_404,N_267);
nand U1056 (N_1056,N_515,N_427);
and U1057 (N_1057,N_135,N_240);
nand U1058 (N_1058,N_401,N_154);
and U1059 (N_1059,N_572,N_241);
or U1060 (N_1060,N_248,N_261);
xor U1061 (N_1061,N_163,N_560);
xor U1062 (N_1062,N_182,N_28);
and U1063 (N_1063,N_580,N_480);
nor U1064 (N_1064,N_434,N_337);
and U1065 (N_1065,N_442,N_81);
or U1066 (N_1066,N_527,N_332);
xnor U1067 (N_1067,N_151,N_410);
and U1068 (N_1068,N_222,N_375);
nor U1069 (N_1069,N_324,N_37);
xnor U1070 (N_1070,N_347,N_424);
nor U1071 (N_1071,N_391,N_194);
nor U1072 (N_1072,N_475,N_198);
and U1073 (N_1073,N_386,N_236);
and U1074 (N_1074,N_536,N_336);
xor U1075 (N_1075,N_2,N_119);
nand U1076 (N_1076,N_43,N_579);
or U1077 (N_1077,N_189,N_539);
xor U1078 (N_1078,N_572,N_284);
and U1079 (N_1079,N_436,N_369);
nand U1080 (N_1080,N_588,N_332);
nand U1081 (N_1081,N_425,N_355);
or U1082 (N_1082,N_196,N_150);
nand U1083 (N_1083,N_404,N_205);
or U1084 (N_1084,N_487,N_492);
nand U1085 (N_1085,N_491,N_365);
and U1086 (N_1086,N_342,N_319);
nand U1087 (N_1087,N_442,N_429);
nor U1088 (N_1088,N_106,N_78);
or U1089 (N_1089,N_109,N_192);
nor U1090 (N_1090,N_276,N_423);
nor U1091 (N_1091,N_378,N_531);
nand U1092 (N_1092,N_476,N_398);
xnor U1093 (N_1093,N_383,N_517);
xnor U1094 (N_1094,N_519,N_458);
nand U1095 (N_1095,N_503,N_260);
nand U1096 (N_1096,N_246,N_269);
nand U1097 (N_1097,N_106,N_566);
or U1098 (N_1098,N_226,N_214);
or U1099 (N_1099,N_97,N_87);
or U1100 (N_1100,N_515,N_591);
nand U1101 (N_1101,N_533,N_17);
or U1102 (N_1102,N_346,N_589);
and U1103 (N_1103,N_237,N_422);
and U1104 (N_1104,N_525,N_490);
nor U1105 (N_1105,N_592,N_421);
nor U1106 (N_1106,N_315,N_267);
or U1107 (N_1107,N_293,N_102);
nand U1108 (N_1108,N_114,N_40);
or U1109 (N_1109,N_169,N_305);
or U1110 (N_1110,N_54,N_451);
or U1111 (N_1111,N_273,N_90);
nand U1112 (N_1112,N_174,N_92);
nand U1113 (N_1113,N_513,N_483);
nand U1114 (N_1114,N_305,N_190);
xor U1115 (N_1115,N_298,N_384);
and U1116 (N_1116,N_269,N_548);
xor U1117 (N_1117,N_47,N_145);
xnor U1118 (N_1118,N_392,N_241);
xor U1119 (N_1119,N_270,N_246);
nor U1120 (N_1120,N_420,N_38);
nor U1121 (N_1121,N_305,N_350);
and U1122 (N_1122,N_332,N_385);
or U1123 (N_1123,N_103,N_548);
and U1124 (N_1124,N_377,N_497);
xor U1125 (N_1125,N_480,N_515);
nand U1126 (N_1126,N_338,N_26);
and U1127 (N_1127,N_215,N_533);
and U1128 (N_1128,N_412,N_211);
and U1129 (N_1129,N_316,N_468);
nor U1130 (N_1130,N_484,N_3);
nand U1131 (N_1131,N_168,N_315);
nand U1132 (N_1132,N_92,N_496);
nand U1133 (N_1133,N_315,N_592);
and U1134 (N_1134,N_463,N_20);
and U1135 (N_1135,N_364,N_573);
nand U1136 (N_1136,N_276,N_264);
and U1137 (N_1137,N_258,N_290);
nor U1138 (N_1138,N_53,N_415);
xnor U1139 (N_1139,N_449,N_573);
and U1140 (N_1140,N_539,N_263);
nor U1141 (N_1141,N_429,N_180);
and U1142 (N_1142,N_283,N_431);
xor U1143 (N_1143,N_290,N_373);
nand U1144 (N_1144,N_230,N_281);
nor U1145 (N_1145,N_133,N_50);
nand U1146 (N_1146,N_297,N_130);
nand U1147 (N_1147,N_135,N_221);
nor U1148 (N_1148,N_31,N_523);
or U1149 (N_1149,N_139,N_390);
nor U1150 (N_1150,N_18,N_103);
nand U1151 (N_1151,N_303,N_360);
nand U1152 (N_1152,N_486,N_230);
nor U1153 (N_1153,N_478,N_233);
nand U1154 (N_1154,N_565,N_194);
and U1155 (N_1155,N_270,N_128);
and U1156 (N_1156,N_430,N_125);
and U1157 (N_1157,N_233,N_98);
nor U1158 (N_1158,N_323,N_547);
xor U1159 (N_1159,N_186,N_430);
xnor U1160 (N_1160,N_376,N_340);
nand U1161 (N_1161,N_361,N_337);
nor U1162 (N_1162,N_532,N_428);
or U1163 (N_1163,N_499,N_516);
xnor U1164 (N_1164,N_141,N_399);
or U1165 (N_1165,N_242,N_321);
xnor U1166 (N_1166,N_209,N_453);
nand U1167 (N_1167,N_342,N_71);
nor U1168 (N_1168,N_313,N_181);
nand U1169 (N_1169,N_21,N_590);
nor U1170 (N_1170,N_32,N_78);
and U1171 (N_1171,N_57,N_297);
nor U1172 (N_1172,N_324,N_235);
or U1173 (N_1173,N_453,N_563);
or U1174 (N_1174,N_534,N_31);
and U1175 (N_1175,N_7,N_281);
or U1176 (N_1176,N_310,N_394);
and U1177 (N_1177,N_20,N_49);
xnor U1178 (N_1178,N_55,N_37);
and U1179 (N_1179,N_54,N_372);
xnor U1180 (N_1180,N_342,N_427);
nor U1181 (N_1181,N_136,N_198);
nor U1182 (N_1182,N_90,N_101);
nand U1183 (N_1183,N_344,N_475);
xnor U1184 (N_1184,N_372,N_326);
xnor U1185 (N_1185,N_329,N_91);
or U1186 (N_1186,N_355,N_323);
xor U1187 (N_1187,N_162,N_349);
nor U1188 (N_1188,N_294,N_108);
xor U1189 (N_1189,N_481,N_511);
nand U1190 (N_1190,N_2,N_523);
and U1191 (N_1191,N_395,N_376);
nand U1192 (N_1192,N_433,N_476);
xor U1193 (N_1193,N_204,N_302);
nor U1194 (N_1194,N_63,N_52);
or U1195 (N_1195,N_303,N_496);
nor U1196 (N_1196,N_373,N_91);
nor U1197 (N_1197,N_124,N_364);
and U1198 (N_1198,N_374,N_98);
or U1199 (N_1199,N_195,N_327);
nand U1200 (N_1200,N_845,N_945);
nor U1201 (N_1201,N_654,N_915);
or U1202 (N_1202,N_1153,N_601);
and U1203 (N_1203,N_780,N_1136);
or U1204 (N_1204,N_1115,N_640);
nand U1205 (N_1205,N_1196,N_981);
xor U1206 (N_1206,N_1046,N_665);
nand U1207 (N_1207,N_899,N_810);
nand U1208 (N_1208,N_628,N_600);
or U1209 (N_1209,N_1175,N_1064);
nor U1210 (N_1210,N_1089,N_952);
xnor U1211 (N_1211,N_902,N_713);
nor U1212 (N_1212,N_834,N_839);
xor U1213 (N_1213,N_1066,N_919);
and U1214 (N_1214,N_956,N_924);
xnor U1215 (N_1215,N_605,N_710);
xor U1216 (N_1216,N_758,N_846);
or U1217 (N_1217,N_662,N_609);
nor U1218 (N_1218,N_630,N_1096);
nor U1219 (N_1219,N_664,N_1053);
xnor U1220 (N_1220,N_1116,N_741);
or U1221 (N_1221,N_1137,N_769);
nand U1222 (N_1222,N_675,N_682);
nand U1223 (N_1223,N_909,N_660);
nand U1224 (N_1224,N_696,N_680);
nor U1225 (N_1225,N_983,N_926);
and U1226 (N_1226,N_1018,N_724);
nor U1227 (N_1227,N_1067,N_782);
nor U1228 (N_1228,N_1155,N_714);
nand U1229 (N_1229,N_905,N_1114);
nand U1230 (N_1230,N_908,N_1073);
nor U1231 (N_1231,N_932,N_975);
or U1232 (N_1232,N_770,N_999);
xor U1233 (N_1233,N_1080,N_1022);
nand U1234 (N_1234,N_1060,N_923);
nor U1235 (N_1235,N_745,N_816);
nor U1236 (N_1236,N_737,N_783);
and U1237 (N_1237,N_1152,N_937);
nand U1238 (N_1238,N_762,N_973);
nor U1239 (N_1239,N_726,N_644);
nor U1240 (N_1240,N_1000,N_732);
and U1241 (N_1241,N_1168,N_1005);
or U1242 (N_1242,N_1058,N_1130);
and U1243 (N_1243,N_832,N_750);
xnor U1244 (N_1244,N_976,N_1122);
nor U1245 (N_1245,N_962,N_1113);
nand U1246 (N_1246,N_969,N_950);
nor U1247 (N_1247,N_970,N_1144);
and U1248 (N_1248,N_616,N_704);
and U1249 (N_1249,N_638,N_916);
nor U1250 (N_1250,N_1062,N_815);
xor U1251 (N_1251,N_844,N_864);
or U1252 (N_1252,N_798,N_1140);
xor U1253 (N_1253,N_865,N_1104);
nor U1254 (N_1254,N_851,N_1019);
nand U1255 (N_1255,N_636,N_869);
or U1256 (N_1256,N_1121,N_1183);
xnor U1257 (N_1257,N_876,N_727);
nand U1258 (N_1258,N_1108,N_820);
nor U1259 (N_1259,N_688,N_1128);
and U1260 (N_1260,N_951,N_868);
xor U1261 (N_1261,N_1097,N_875);
nor U1262 (N_1262,N_928,N_943);
nor U1263 (N_1263,N_610,N_803);
nor U1264 (N_1264,N_1186,N_870);
or U1265 (N_1265,N_944,N_1041);
nor U1266 (N_1266,N_1030,N_786);
and U1267 (N_1267,N_645,N_717);
xnor U1268 (N_1268,N_1143,N_883);
and U1269 (N_1269,N_1059,N_775);
xnor U1270 (N_1270,N_754,N_894);
nor U1271 (N_1271,N_625,N_957);
xnor U1272 (N_1272,N_812,N_1055);
xor U1273 (N_1273,N_1156,N_854);
xnor U1274 (N_1274,N_1195,N_994);
nor U1275 (N_1275,N_1159,N_1161);
xor U1276 (N_1276,N_1012,N_639);
and U1277 (N_1277,N_871,N_1024);
and U1278 (N_1278,N_1095,N_1149);
nand U1279 (N_1279,N_1084,N_1038);
nor U1280 (N_1280,N_708,N_931);
nor U1281 (N_1281,N_980,N_1169);
xnor U1282 (N_1282,N_760,N_930);
xnor U1283 (N_1283,N_720,N_692);
xor U1284 (N_1284,N_697,N_860);
nand U1285 (N_1285,N_825,N_764);
nand U1286 (N_1286,N_964,N_992);
nor U1287 (N_1287,N_1166,N_723);
nand U1288 (N_1288,N_650,N_721);
xnor U1289 (N_1289,N_1052,N_706);
or U1290 (N_1290,N_824,N_1174);
nand U1291 (N_1291,N_814,N_1070);
xnor U1292 (N_1292,N_800,N_1001);
and U1293 (N_1293,N_1151,N_672);
and U1294 (N_1294,N_1162,N_757);
nand U1295 (N_1295,N_913,N_1016);
xnor U1296 (N_1296,N_1043,N_1150);
nand U1297 (N_1297,N_779,N_888);
nor U1298 (N_1298,N_698,N_797);
and U1299 (N_1299,N_748,N_1184);
xor U1300 (N_1300,N_1085,N_668);
nor U1301 (N_1301,N_968,N_895);
and U1302 (N_1302,N_1083,N_1033);
xnor U1303 (N_1303,N_1106,N_848);
nand U1304 (N_1304,N_1111,N_847);
nor U1305 (N_1305,N_1123,N_744);
xnor U1306 (N_1306,N_1103,N_614);
nand U1307 (N_1307,N_882,N_922);
nand U1308 (N_1308,N_947,N_1126);
or U1309 (N_1309,N_648,N_903);
nor U1310 (N_1310,N_821,N_763);
or U1311 (N_1311,N_687,N_1146);
and U1312 (N_1312,N_773,N_877);
nand U1313 (N_1313,N_948,N_655);
xnor U1314 (N_1314,N_778,N_828);
and U1315 (N_1315,N_889,N_850);
or U1316 (N_1316,N_604,N_606);
nor U1317 (N_1317,N_707,N_852);
or U1318 (N_1318,N_646,N_700);
or U1319 (N_1319,N_901,N_1118);
and U1320 (N_1320,N_771,N_986);
xor U1321 (N_1321,N_751,N_796);
nand U1322 (N_1322,N_1142,N_965);
and U1323 (N_1323,N_1119,N_642);
and U1324 (N_1324,N_772,N_730);
nor U1325 (N_1325,N_794,N_629);
and U1326 (N_1326,N_1002,N_792);
and U1327 (N_1327,N_1050,N_920);
nand U1328 (N_1328,N_728,N_934);
or U1329 (N_1329,N_898,N_925);
and U1330 (N_1330,N_653,N_1177);
xnor U1331 (N_1331,N_1091,N_607);
xnor U1332 (N_1332,N_1117,N_966);
nor U1333 (N_1333,N_826,N_971);
and U1334 (N_1334,N_613,N_1078);
xor U1335 (N_1335,N_656,N_693);
and U1336 (N_1336,N_939,N_768);
or U1337 (N_1337,N_749,N_1093);
nor U1338 (N_1338,N_1160,N_702);
nand U1339 (N_1339,N_1132,N_1071);
xor U1340 (N_1340,N_1061,N_695);
nor U1341 (N_1341,N_1129,N_1029);
and U1342 (N_1342,N_1098,N_1020);
nor U1343 (N_1343,N_1063,N_1148);
or U1344 (N_1344,N_1110,N_1023);
xnor U1345 (N_1345,N_880,N_892);
nor U1346 (N_1346,N_1185,N_1191);
nor U1347 (N_1347,N_960,N_1188);
nor U1348 (N_1348,N_1090,N_685);
xnor U1349 (N_1349,N_997,N_1009);
nor U1350 (N_1350,N_718,N_837);
xnor U1351 (N_1351,N_761,N_603);
nor U1352 (N_1352,N_719,N_840);
nand U1353 (N_1353,N_1057,N_705);
nor U1354 (N_1354,N_701,N_1049);
nor U1355 (N_1355,N_990,N_1036);
nor U1356 (N_1356,N_855,N_953);
and U1357 (N_1357,N_1109,N_878);
xor U1358 (N_1358,N_801,N_678);
nand U1359 (N_1359,N_791,N_716);
nand U1360 (N_1360,N_862,N_1154);
nor U1361 (N_1361,N_918,N_1021);
and U1362 (N_1362,N_681,N_793);
and U1363 (N_1363,N_1105,N_831);
nand U1364 (N_1364,N_808,N_784);
nor U1365 (N_1365,N_979,N_776);
nand U1366 (N_1366,N_729,N_740);
nand U1367 (N_1367,N_1079,N_881);
nor U1368 (N_1368,N_673,N_711);
or U1369 (N_1369,N_1141,N_900);
nor U1370 (N_1370,N_1145,N_627);
nand U1371 (N_1371,N_1170,N_1164);
nand U1372 (N_1372,N_1147,N_1176);
and U1373 (N_1373,N_958,N_838);
or U1374 (N_1374,N_818,N_1194);
nand U1375 (N_1375,N_799,N_617);
or U1376 (N_1376,N_746,N_1139);
xor U1377 (N_1377,N_1100,N_735);
or U1378 (N_1378,N_941,N_977);
xnor U1379 (N_1379,N_927,N_914);
and U1380 (N_1380,N_835,N_1013);
nor U1381 (N_1381,N_805,N_954);
nor U1382 (N_1382,N_911,N_658);
nand U1383 (N_1383,N_1075,N_813);
xor U1384 (N_1384,N_946,N_1127);
nor U1385 (N_1385,N_804,N_703);
xor U1386 (N_1386,N_1192,N_1158);
nor U1387 (N_1387,N_1172,N_993);
xnor U1388 (N_1388,N_829,N_912);
nor U1389 (N_1389,N_766,N_972);
and U1390 (N_1390,N_1068,N_679);
xor U1391 (N_1391,N_1008,N_929);
nand U1392 (N_1392,N_1081,N_666);
or U1393 (N_1393,N_822,N_1134);
or U1394 (N_1394,N_1056,N_663);
nor U1395 (N_1395,N_989,N_857);
or U1396 (N_1396,N_1037,N_674);
and U1397 (N_1397,N_949,N_873);
xor U1398 (N_1398,N_1015,N_1042);
or U1399 (N_1399,N_615,N_942);
nand U1400 (N_1400,N_1133,N_643);
or U1401 (N_1401,N_1167,N_1007);
and U1402 (N_1402,N_1125,N_1044);
or U1403 (N_1403,N_1112,N_1047);
or U1404 (N_1404,N_885,N_1035);
nand U1405 (N_1405,N_955,N_620);
or U1406 (N_1406,N_1011,N_1025);
and U1407 (N_1407,N_752,N_910);
xor U1408 (N_1408,N_623,N_802);
nor U1409 (N_1409,N_747,N_670);
nor U1410 (N_1410,N_1102,N_1039);
and U1411 (N_1411,N_836,N_1124);
xnor U1412 (N_1412,N_1028,N_686);
xor U1413 (N_1413,N_709,N_933);
nor U1414 (N_1414,N_1006,N_1077);
nand U1415 (N_1415,N_677,N_611);
and U1416 (N_1416,N_842,N_982);
or U1417 (N_1417,N_1069,N_1187);
or U1418 (N_1418,N_1086,N_1198);
nand U1419 (N_1419,N_866,N_1180);
or U1420 (N_1420,N_1082,N_887);
xor U1421 (N_1421,N_785,N_959);
or U1422 (N_1422,N_936,N_907);
or U1423 (N_1423,N_988,N_987);
xor U1424 (N_1424,N_753,N_1048);
xnor U1425 (N_1425,N_635,N_890);
xor U1426 (N_1426,N_830,N_938);
nor U1427 (N_1427,N_1027,N_1190);
nor U1428 (N_1428,N_742,N_739);
nand U1429 (N_1429,N_632,N_684);
and U1430 (N_1430,N_691,N_647);
or U1431 (N_1431,N_633,N_1120);
or U1432 (N_1432,N_1054,N_1010);
nand U1433 (N_1433,N_995,N_722);
xnor U1434 (N_1434,N_634,N_1131);
xor U1435 (N_1435,N_1157,N_734);
and U1436 (N_1436,N_891,N_811);
and U1437 (N_1437,N_1199,N_884);
and U1438 (N_1438,N_897,N_906);
nand U1439 (N_1439,N_861,N_712);
xor U1440 (N_1440,N_817,N_940);
or U1441 (N_1441,N_823,N_1088);
nand U1442 (N_1442,N_602,N_659);
and U1443 (N_1443,N_649,N_756);
or U1444 (N_1444,N_859,N_1173);
and U1445 (N_1445,N_781,N_765);
xor U1446 (N_1446,N_879,N_789);
or U1447 (N_1447,N_841,N_1003);
xnor U1448 (N_1448,N_671,N_843);
nand U1449 (N_1449,N_774,N_984);
or U1450 (N_1450,N_809,N_874);
and U1451 (N_1451,N_657,N_985);
xor U1452 (N_1452,N_624,N_967);
and U1453 (N_1453,N_1076,N_612);
or U1454 (N_1454,N_991,N_618);
and U1455 (N_1455,N_996,N_690);
or U1456 (N_1456,N_699,N_715);
or U1457 (N_1457,N_1101,N_858);
or U1458 (N_1458,N_736,N_651);
and U1459 (N_1459,N_725,N_790);
nand U1460 (N_1460,N_819,N_652);
xnor U1461 (N_1461,N_1179,N_1197);
nand U1462 (N_1462,N_893,N_637);
and U1463 (N_1463,N_863,N_1163);
and U1464 (N_1464,N_1034,N_689);
or U1465 (N_1465,N_1017,N_1040);
xor U1466 (N_1466,N_683,N_1031);
or U1467 (N_1467,N_853,N_694);
xnor U1468 (N_1468,N_849,N_974);
xor U1469 (N_1469,N_1182,N_669);
and U1470 (N_1470,N_641,N_896);
or U1471 (N_1471,N_1045,N_1032);
and U1472 (N_1472,N_743,N_1087);
or U1473 (N_1473,N_807,N_1171);
and U1474 (N_1474,N_755,N_759);
and U1475 (N_1475,N_733,N_978);
and U1476 (N_1476,N_856,N_622);
or U1477 (N_1477,N_787,N_1189);
nand U1478 (N_1478,N_961,N_1193);
nor U1479 (N_1479,N_767,N_1138);
nand U1480 (N_1480,N_795,N_872);
xor U1481 (N_1481,N_833,N_608);
and U1482 (N_1482,N_676,N_963);
or U1483 (N_1483,N_1092,N_1099);
and U1484 (N_1484,N_867,N_886);
nand U1485 (N_1485,N_806,N_1072);
and U1486 (N_1486,N_661,N_626);
nor U1487 (N_1487,N_1165,N_1135);
nor U1488 (N_1488,N_935,N_788);
xor U1489 (N_1489,N_1107,N_1026);
nand U1490 (N_1490,N_731,N_1181);
or U1491 (N_1491,N_1178,N_621);
nand U1492 (N_1492,N_917,N_631);
and U1493 (N_1493,N_619,N_904);
and U1494 (N_1494,N_827,N_1051);
xor U1495 (N_1495,N_1014,N_1004);
nand U1496 (N_1496,N_998,N_921);
nand U1497 (N_1497,N_1074,N_738);
or U1498 (N_1498,N_777,N_667);
or U1499 (N_1499,N_1065,N_1094);
and U1500 (N_1500,N_697,N_927);
and U1501 (N_1501,N_710,N_715);
nand U1502 (N_1502,N_1180,N_1118);
xnor U1503 (N_1503,N_1105,N_945);
or U1504 (N_1504,N_1129,N_1087);
nand U1505 (N_1505,N_862,N_940);
or U1506 (N_1506,N_651,N_847);
nand U1507 (N_1507,N_991,N_1166);
nor U1508 (N_1508,N_683,N_640);
and U1509 (N_1509,N_954,N_1076);
xnor U1510 (N_1510,N_1115,N_1118);
or U1511 (N_1511,N_1069,N_994);
xnor U1512 (N_1512,N_641,N_1015);
and U1513 (N_1513,N_928,N_835);
xor U1514 (N_1514,N_629,N_924);
or U1515 (N_1515,N_1019,N_1018);
and U1516 (N_1516,N_895,N_1002);
nor U1517 (N_1517,N_1117,N_920);
nand U1518 (N_1518,N_638,N_883);
nor U1519 (N_1519,N_708,N_1026);
xor U1520 (N_1520,N_678,N_1103);
xnor U1521 (N_1521,N_699,N_719);
or U1522 (N_1522,N_1190,N_620);
nand U1523 (N_1523,N_749,N_1186);
xor U1524 (N_1524,N_1160,N_698);
and U1525 (N_1525,N_792,N_1017);
nand U1526 (N_1526,N_699,N_789);
nor U1527 (N_1527,N_1112,N_933);
xor U1528 (N_1528,N_648,N_626);
and U1529 (N_1529,N_840,N_695);
nand U1530 (N_1530,N_974,N_695);
xnor U1531 (N_1531,N_959,N_762);
xnor U1532 (N_1532,N_1085,N_841);
and U1533 (N_1533,N_1016,N_648);
or U1534 (N_1534,N_1123,N_673);
xor U1535 (N_1535,N_627,N_1126);
nor U1536 (N_1536,N_768,N_798);
xor U1537 (N_1537,N_1165,N_1047);
or U1538 (N_1538,N_850,N_603);
nand U1539 (N_1539,N_1075,N_953);
nand U1540 (N_1540,N_932,N_974);
xnor U1541 (N_1541,N_665,N_1014);
nor U1542 (N_1542,N_1196,N_655);
or U1543 (N_1543,N_790,N_805);
and U1544 (N_1544,N_989,N_600);
nor U1545 (N_1545,N_691,N_704);
and U1546 (N_1546,N_948,N_861);
and U1547 (N_1547,N_693,N_927);
and U1548 (N_1548,N_954,N_702);
and U1549 (N_1549,N_1173,N_744);
nand U1550 (N_1550,N_746,N_846);
xnor U1551 (N_1551,N_628,N_1108);
or U1552 (N_1552,N_921,N_1004);
nand U1553 (N_1553,N_983,N_1164);
and U1554 (N_1554,N_1117,N_1091);
xor U1555 (N_1555,N_897,N_633);
nand U1556 (N_1556,N_1119,N_757);
nand U1557 (N_1557,N_837,N_746);
or U1558 (N_1558,N_799,N_908);
and U1559 (N_1559,N_830,N_715);
or U1560 (N_1560,N_1026,N_764);
nand U1561 (N_1561,N_608,N_1114);
and U1562 (N_1562,N_1195,N_1164);
xnor U1563 (N_1563,N_698,N_977);
xnor U1564 (N_1564,N_947,N_961);
and U1565 (N_1565,N_1163,N_938);
xor U1566 (N_1566,N_679,N_768);
xor U1567 (N_1567,N_982,N_687);
xor U1568 (N_1568,N_1057,N_762);
nor U1569 (N_1569,N_997,N_778);
xor U1570 (N_1570,N_884,N_1060);
nand U1571 (N_1571,N_681,N_1047);
nand U1572 (N_1572,N_1114,N_1139);
xnor U1573 (N_1573,N_1174,N_1163);
or U1574 (N_1574,N_1011,N_759);
xor U1575 (N_1575,N_1032,N_772);
and U1576 (N_1576,N_935,N_809);
xnor U1577 (N_1577,N_693,N_673);
or U1578 (N_1578,N_1143,N_1132);
and U1579 (N_1579,N_1029,N_1137);
xnor U1580 (N_1580,N_1163,N_1177);
and U1581 (N_1581,N_853,N_1111);
and U1582 (N_1582,N_1033,N_1196);
nand U1583 (N_1583,N_865,N_1000);
nand U1584 (N_1584,N_1067,N_967);
or U1585 (N_1585,N_1089,N_780);
and U1586 (N_1586,N_775,N_874);
and U1587 (N_1587,N_881,N_728);
xnor U1588 (N_1588,N_1032,N_804);
nor U1589 (N_1589,N_760,N_1153);
nand U1590 (N_1590,N_1163,N_922);
or U1591 (N_1591,N_1109,N_1039);
xor U1592 (N_1592,N_918,N_766);
or U1593 (N_1593,N_811,N_1081);
xnor U1594 (N_1594,N_875,N_642);
xor U1595 (N_1595,N_621,N_817);
or U1596 (N_1596,N_1104,N_864);
xnor U1597 (N_1597,N_855,N_644);
xnor U1598 (N_1598,N_602,N_647);
xnor U1599 (N_1599,N_1048,N_873);
or U1600 (N_1600,N_1188,N_768);
nor U1601 (N_1601,N_852,N_877);
and U1602 (N_1602,N_709,N_640);
xnor U1603 (N_1603,N_1151,N_961);
and U1604 (N_1604,N_1124,N_816);
nor U1605 (N_1605,N_741,N_948);
nor U1606 (N_1606,N_807,N_769);
or U1607 (N_1607,N_946,N_822);
xnor U1608 (N_1608,N_903,N_874);
nor U1609 (N_1609,N_1052,N_899);
xor U1610 (N_1610,N_939,N_1105);
and U1611 (N_1611,N_842,N_862);
nand U1612 (N_1612,N_713,N_787);
nand U1613 (N_1613,N_1051,N_1006);
or U1614 (N_1614,N_948,N_779);
xnor U1615 (N_1615,N_952,N_788);
xnor U1616 (N_1616,N_1093,N_838);
and U1617 (N_1617,N_998,N_827);
and U1618 (N_1618,N_656,N_715);
nor U1619 (N_1619,N_1010,N_1154);
xor U1620 (N_1620,N_1072,N_1032);
nor U1621 (N_1621,N_850,N_992);
nor U1622 (N_1622,N_1113,N_682);
and U1623 (N_1623,N_926,N_802);
xor U1624 (N_1624,N_997,N_965);
and U1625 (N_1625,N_651,N_1108);
nor U1626 (N_1626,N_1127,N_934);
or U1627 (N_1627,N_875,N_727);
or U1628 (N_1628,N_810,N_877);
nor U1629 (N_1629,N_881,N_795);
nor U1630 (N_1630,N_696,N_962);
nor U1631 (N_1631,N_763,N_818);
xor U1632 (N_1632,N_1096,N_994);
and U1633 (N_1633,N_625,N_853);
and U1634 (N_1634,N_1098,N_1104);
or U1635 (N_1635,N_1097,N_1174);
or U1636 (N_1636,N_897,N_1100);
nor U1637 (N_1637,N_1174,N_1147);
nor U1638 (N_1638,N_959,N_834);
nor U1639 (N_1639,N_695,N_716);
xnor U1640 (N_1640,N_830,N_1111);
nand U1641 (N_1641,N_987,N_752);
nor U1642 (N_1642,N_630,N_1187);
and U1643 (N_1643,N_789,N_656);
nand U1644 (N_1644,N_1122,N_862);
and U1645 (N_1645,N_604,N_845);
nand U1646 (N_1646,N_1002,N_627);
xnor U1647 (N_1647,N_921,N_1066);
and U1648 (N_1648,N_1189,N_1102);
xnor U1649 (N_1649,N_814,N_829);
xnor U1650 (N_1650,N_855,N_856);
or U1651 (N_1651,N_1069,N_919);
or U1652 (N_1652,N_1023,N_1066);
xor U1653 (N_1653,N_744,N_1079);
or U1654 (N_1654,N_741,N_659);
nand U1655 (N_1655,N_855,N_653);
or U1656 (N_1656,N_1083,N_833);
nor U1657 (N_1657,N_1133,N_749);
and U1658 (N_1658,N_1005,N_966);
xnor U1659 (N_1659,N_656,N_808);
or U1660 (N_1660,N_901,N_849);
xor U1661 (N_1661,N_728,N_1056);
and U1662 (N_1662,N_1194,N_609);
xor U1663 (N_1663,N_910,N_720);
nand U1664 (N_1664,N_776,N_985);
xnor U1665 (N_1665,N_1019,N_810);
xnor U1666 (N_1666,N_1064,N_1152);
nor U1667 (N_1667,N_830,N_1008);
and U1668 (N_1668,N_821,N_1025);
or U1669 (N_1669,N_897,N_641);
xnor U1670 (N_1670,N_737,N_1058);
nand U1671 (N_1671,N_1144,N_944);
nand U1672 (N_1672,N_959,N_683);
nor U1673 (N_1673,N_718,N_1167);
nand U1674 (N_1674,N_1155,N_1082);
or U1675 (N_1675,N_628,N_1059);
nor U1676 (N_1676,N_627,N_1123);
xnor U1677 (N_1677,N_970,N_791);
nor U1678 (N_1678,N_860,N_1029);
nand U1679 (N_1679,N_692,N_645);
nor U1680 (N_1680,N_691,N_1165);
or U1681 (N_1681,N_1028,N_1097);
xnor U1682 (N_1682,N_982,N_840);
xnor U1683 (N_1683,N_829,N_1148);
nor U1684 (N_1684,N_1177,N_626);
nand U1685 (N_1685,N_890,N_687);
nand U1686 (N_1686,N_655,N_1042);
nand U1687 (N_1687,N_608,N_1015);
or U1688 (N_1688,N_629,N_846);
and U1689 (N_1689,N_657,N_821);
and U1690 (N_1690,N_1123,N_833);
or U1691 (N_1691,N_903,N_772);
and U1692 (N_1692,N_679,N_783);
nor U1693 (N_1693,N_1029,N_853);
nor U1694 (N_1694,N_921,N_736);
and U1695 (N_1695,N_696,N_1135);
nand U1696 (N_1696,N_1063,N_738);
nor U1697 (N_1697,N_1001,N_1048);
nor U1698 (N_1698,N_1072,N_995);
and U1699 (N_1699,N_1092,N_719);
nor U1700 (N_1700,N_854,N_860);
nand U1701 (N_1701,N_811,N_1102);
and U1702 (N_1702,N_876,N_980);
xnor U1703 (N_1703,N_659,N_983);
xor U1704 (N_1704,N_746,N_641);
or U1705 (N_1705,N_1059,N_972);
nand U1706 (N_1706,N_789,N_873);
nand U1707 (N_1707,N_879,N_781);
xnor U1708 (N_1708,N_848,N_1005);
and U1709 (N_1709,N_640,N_990);
xor U1710 (N_1710,N_1077,N_1083);
and U1711 (N_1711,N_963,N_1109);
xnor U1712 (N_1712,N_1057,N_660);
xor U1713 (N_1713,N_1040,N_1068);
or U1714 (N_1714,N_648,N_674);
or U1715 (N_1715,N_690,N_838);
or U1716 (N_1716,N_868,N_952);
or U1717 (N_1717,N_926,N_1146);
nand U1718 (N_1718,N_601,N_1057);
nand U1719 (N_1719,N_1128,N_604);
nand U1720 (N_1720,N_653,N_1153);
nand U1721 (N_1721,N_1192,N_1130);
nand U1722 (N_1722,N_1177,N_869);
xor U1723 (N_1723,N_848,N_983);
and U1724 (N_1724,N_1062,N_1122);
and U1725 (N_1725,N_790,N_716);
nand U1726 (N_1726,N_704,N_682);
nor U1727 (N_1727,N_1085,N_964);
and U1728 (N_1728,N_1002,N_790);
and U1729 (N_1729,N_1195,N_792);
or U1730 (N_1730,N_912,N_844);
and U1731 (N_1731,N_943,N_876);
xnor U1732 (N_1732,N_1019,N_1029);
nand U1733 (N_1733,N_1081,N_1129);
or U1734 (N_1734,N_1127,N_763);
and U1735 (N_1735,N_814,N_635);
and U1736 (N_1736,N_810,N_612);
and U1737 (N_1737,N_889,N_672);
xnor U1738 (N_1738,N_974,N_669);
or U1739 (N_1739,N_688,N_1193);
or U1740 (N_1740,N_1109,N_982);
nor U1741 (N_1741,N_1180,N_718);
nand U1742 (N_1742,N_753,N_1102);
nor U1743 (N_1743,N_807,N_948);
nand U1744 (N_1744,N_1092,N_695);
nor U1745 (N_1745,N_1006,N_1054);
or U1746 (N_1746,N_900,N_1169);
nand U1747 (N_1747,N_759,N_885);
nor U1748 (N_1748,N_1051,N_1088);
nand U1749 (N_1749,N_1088,N_744);
or U1750 (N_1750,N_702,N_1016);
nor U1751 (N_1751,N_1130,N_671);
and U1752 (N_1752,N_799,N_666);
or U1753 (N_1753,N_1029,N_967);
nor U1754 (N_1754,N_792,N_840);
and U1755 (N_1755,N_889,N_710);
nand U1756 (N_1756,N_1101,N_1021);
nor U1757 (N_1757,N_1171,N_648);
or U1758 (N_1758,N_802,N_870);
xnor U1759 (N_1759,N_1191,N_663);
nand U1760 (N_1760,N_781,N_1092);
and U1761 (N_1761,N_820,N_777);
nand U1762 (N_1762,N_1075,N_920);
and U1763 (N_1763,N_1045,N_1153);
nor U1764 (N_1764,N_613,N_808);
and U1765 (N_1765,N_900,N_706);
nor U1766 (N_1766,N_1175,N_614);
xor U1767 (N_1767,N_1060,N_1158);
nand U1768 (N_1768,N_688,N_847);
or U1769 (N_1769,N_756,N_1162);
nor U1770 (N_1770,N_886,N_997);
or U1771 (N_1771,N_1177,N_888);
nor U1772 (N_1772,N_941,N_696);
xnor U1773 (N_1773,N_652,N_967);
or U1774 (N_1774,N_771,N_845);
or U1775 (N_1775,N_1123,N_845);
or U1776 (N_1776,N_732,N_1016);
nor U1777 (N_1777,N_1156,N_723);
xor U1778 (N_1778,N_879,N_829);
nand U1779 (N_1779,N_1035,N_975);
nor U1780 (N_1780,N_767,N_908);
xnor U1781 (N_1781,N_625,N_1109);
xnor U1782 (N_1782,N_1074,N_973);
or U1783 (N_1783,N_974,N_636);
or U1784 (N_1784,N_1198,N_663);
and U1785 (N_1785,N_953,N_942);
xor U1786 (N_1786,N_651,N_913);
or U1787 (N_1787,N_642,N_600);
xnor U1788 (N_1788,N_895,N_865);
or U1789 (N_1789,N_668,N_873);
nand U1790 (N_1790,N_1172,N_1077);
nand U1791 (N_1791,N_971,N_979);
xor U1792 (N_1792,N_1117,N_628);
nor U1793 (N_1793,N_953,N_834);
and U1794 (N_1794,N_1000,N_996);
xnor U1795 (N_1795,N_661,N_879);
nand U1796 (N_1796,N_1047,N_1163);
and U1797 (N_1797,N_942,N_1191);
nor U1798 (N_1798,N_1001,N_612);
and U1799 (N_1799,N_1011,N_856);
nor U1800 (N_1800,N_1359,N_1427);
nor U1801 (N_1801,N_1662,N_1680);
nand U1802 (N_1802,N_1306,N_1297);
xor U1803 (N_1803,N_1565,N_1489);
and U1804 (N_1804,N_1780,N_1686);
and U1805 (N_1805,N_1731,N_1323);
xor U1806 (N_1806,N_1512,N_1606);
xor U1807 (N_1807,N_1472,N_1574);
or U1808 (N_1808,N_1794,N_1553);
xor U1809 (N_1809,N_1246,N_1313);
xnor U1810 (N_1810,N_1714,N_1629);
nand U1811 (N_1811,N_1201,N_1231);
nor U1812 (N_1812,N_1652,N_1228);
or U1813 (N_1813,N_1307,N_1727);
nand U1814 (N_1814,N_1703,N_1263);
or U1815 (N_1815,N_1719,N_1690);
and U1816 (N_1816,N_1309,N_1315);
nor U1817 (N_1817,N_1508,N_1345);
and U1818 (N_1818,N_1344,N_1599);
nand U1819 (N_1819,N_1774,N_1608);
and U1820 (N_1820,N_1486,N_1239);
or U1821 (N_1821,N_1535,N_1772);
xnor U1822 (N_1822,N_1651,N_1378);
nor U1823 (N_1823,N_1254,N_1337);
or U1824 (N_1824,N_1640,N_1401);
xnor U1825 (N_1825,N_1663,N_1426);
and U1826 (N_1826,N_1412,N_1525);
and U1827 (N_1827,N_1406,N_1795);
or U1828 (N_1828,N_1745,N_1206);
nand U1829 (N_1829,N_1767,N_1236);
nand U1830 (N_1830,N_1351,N_1335);
nand U1831 (N_1831,N_1783,N_1583);
nand U1832 (N_1832,N_1593,N_1630);
nand U1833 (N_1833,N_1688,N_1717);
nand U1834 (N_1834,N_1367,N_1229);
or U1835 (N_1835,N_1682,N_1476);
nand U1836 (N_1836,N_1329,N_1558);
and U1837 (N_1837,N_1726,N_1591);
or U1838 (N_1838,N_1789,N_1528);
nand U1839 (N_1839,N_1289,N_1654);
or U1840 (N_1840,N_1245,N_1338);
and U1841 (N_1841,N_1437,N_1483);
or U1842 (N_1842,N_1220,N_1756);
or U1843 (N_1843,N_1222,N_1432);
or U1844 (N_1844,N_1271,N_1475);
and U1845 (N_1845,N_1588,N_1276);
nand U1846 (N_1846,N_1739,N_1385);
nand U1847 (N_1847,N_1649,N_1537);
xnor U1848 (N_1848,N_1672,N_1562);
and U1849 (N_1849,N_1339,N_1734);
nor U1850 (N_1850,N_1752,N_1658);
xnor U1851 (N_1851,N_1761,N_1624);
or U1852 (N_1852,N_1454,N_1763);
or U1853 (N_1853,N_1350,N_1547);
and U1854 (N_1854,N_1242,N_1718);
nor U1855 (N_1855,N_1365,N_1623);
xor U1856 (N_1856,N_1700,N_1511);
and U1857 (N_1857,N_1790,N_1711);
nor U1858 (N_1858,N_1447,N_1346);
xnor U1859 (N_1859,N_1601,N_1459);
nor U1860 (N_1860,N_1667,N_1358);
and U1861 (N_1861,N_1393,N_1516);
or U1862 (N_1862,N_1692,N_1261);
and U1863 (N_1863,N_1747,N_1764);
nand U1864 (N_1864,N_1320,N_1650);
nand U1865 (N_1865,N_1278,N_1466);
nor U1866 (N_1866,N_1434,N_1460);
xnor U1867 (N_1867,N_1545,N_1636);
or U1868 (N_1868,N_1736,N_1744);
or U1869 (N_1869,N_1281,N_1694);
nand U1870 (N_1870,N_1491,N_1549);
and U1871 (N_1871,N_1380,N_1404);
and U1872 (N_1872,N_1270,N_1304);
or U1873 (N_1873,N_1387,N_1542);
and U1874 (N_1874,N_1587,N_1217);
or U1875 (N_1875,N_1334,N_1439);
and U1876 (N_1876,N_1594,N_1693);
xnor U1877 (N_1877,N_1341,N_1527);
nor U1878 (N_1878,N_1474,N_1219);
or U1879 (N_1879,N_1247,N_1312);
and U1880 (N_1880,N_1259,N_1453);
and U1881 (N_1881,N_1240,N_1251);
nand U1882 (N_1882,N_1584,N_1514);
nand U1883 (N_1883,N_1522,N_1531);
and U1884 (N_1884,N_1668,N_1523);
or U1885 (N_1885,N_1269,N_1684);
xor U1886 (N_1886,N_1610,N_1664);
nand U1887 (N_1887,N_1518,N_1695);
and U1888 (N_1888,N_1445,N_1742);
and U1889 (N_1889,N_1696,N_1235);
and U1890 (N_1890,N_1602,N_1382);
nand U1891 (N_1891,N_1328,N_1567);
nand U1892 (N_1892,N_1478,N_1233);
nand U1893 (N_1893,N_1619,N_1493);
and U1894 (N_1894,N_1291,N_1332);
xor U1895 (N_1895,N_1321,N_1376);
nor U1896 (N_1896,N_1792,N_1796);
nor U1897 (N_1897,N_1502,N_1784);
or U1898 (N_1898,N_1748,N_1670);
nor U1899 (N_1899,N_1722,N_1521);
xnor U1900 (N_1900,N_1749,N_1230);
xor U1901 (N_1901,N_1616,N_1685);
and U1902 (N_1902,N_1347,N_1279);
and U1903 (N_1903,N_1632,N_1373);
or U1904 (N_1904,N_1433,N_1724);
xor U1905 (N_1905,N_1300,N_1721);
xor U1906 (N_1906,N_1555,N_1410);
or U1907 (N_1907,N_1557,N_1755);
xnor U1908 (N_1908,N_1462,N_1637);
or U1909 (N_1909,N_1793,N_1620);
nor U1910 (N_1910,N_1762,N_1471);
nor U1911 (N_1911,N_1260,N_1589);
nor U1912 (N_1912,N_1701,N_1311);
xnor U1913 (N_1913,N_1504,N_1324);
nor U1914 (N_1914,N_1372,N_1213);
nand U1915 (N_1915,N_1325,N_1733);
or U1916 (N_1916,N_1543,N_1364);
nor U1917 (N_1917,N_1292,N_1465);
and U1918 (N_1918,N_1209,N_1458);
xor U1919 (N_1919,N_1787,N_1729);
or U1920 (N_1920,N_1529,N_1609);
nor U1921 (N_1921,N_1411,N_1530);
xor U1922 (N_1922,N_1698,N_1409);
and U1923 (N_1923,N_1282,N_1419);
nand U1924 (N_1924,N_1286,N_1550);
nor U1925 (N_1925,N_1635,N_1687);
xnor U1926 (N_1926,N_1446,N_1255);
or U1927 (N_1927,N_1314,N_1705);
nand U1928 (N_1928,N_1211,N_1730);
nand U1929 (N_1929,N_1503,N_1782);
and U1930 (N_1930,N_1732,N_1571);
or U1931 (N_1931,N_1781,N_1797);
nor U1932 (N_1932,N_1226,N_1786);
and U1933 (N_1933,N_1538,N_1354);
xor U1934 (N_1934,N_1425,N_1488);
and U1935 (N_1935,N_1671,N_1681);
nand U1936 (N_1936,N_1519,N_1451);
nor U1937 (N_1937,N_1738,N_1467);
nand U1938 (N_1938,N_1622,N_1218);
nor U1939 (N_1939,N_1495,N_1268);
nand U1940 (N_1940,N_1487,N_1704);
nor U1941 (N_1941,N_1368,N_1507);
or U1942 (N_1942,N_1417,N_1431);
nand U1943 (N_1943,N_1713,N_1441);
nand U1944 (N_1944,N_1423,N_1390);
or U1945 (N_1945,N_1227,N_1444);
xor U1946 (N_1946,N_1596,N_1643);
nor U1947 (N_1947,N_1646,N_1580);
or U1948 (N_1948,N_1536,N_1352);
and U1949 (N_1949,N_1340,N_1470);
and U1950 (N_1950,N_1208,N_1674);
and U1951 (N_1951,N_1520,N_1293);
nand U1952 (N_1952,N_1277,N_1225);
or U1953 (N_1953,N_1430,N_1689);
or U1954 (N_1954,N_1485,N_1232);
and U1955 (N_1955,N_1707,N_1319);
nor U1956 (N_1956,N_1216,N_1394);
and U1957 (N_1957,N_1655,N_1750);
or U1958 (N_1958,N_1505,N_1777);
or U1959 (N_1959,N_1768,N_1765);
and U1960 (N_1960,N_1515,N_1443);
xnor U1961 (N_1961,N_1403,N_1564);
xnor U1962 (N_1962,N_1613,N_1611);
nand U1963 (N_1963,N_1205,N_1280);
and U1964 (N_1964,N_1723,N_1284);
and U1965 (N_1965,N_1665,N_1395);
nand U1966 (N_1966,N_1362,N_1577);
nor U1967 (N_1967,N_1308,N_1449);
nor U1968 (N_1968,N_1627,N_1375);
nor U1969 (N_1969,N_1464,N_1510);
and U1970 (N_1970,N_1590,N_1773);
nand U1971 (N_1971,N_1473,N_1285);
nand U1972 (N_1972,N_1391,N_1746);
xnor U1973 (N_1973,N_1679,N_1303);
and U1974 (N_1974,N_1371,N_1469);
nor U1975 (N_1975,N_1612,N_1678);
or U1976 (N_1976,N_1477,N_1617);
nand U1977 (N_1977,N_1200,N_1581);
xnor U1978 (N_1978,N_1429,N_1221);
xor U1979 (N_1979,N_1625,N_1356);
xnor U1980 (N_1980,N_1283,N_1657);
nand U1981 (N_1981,N_1592,N_1585);
and U1982 (N_1982,N_1386,N_1603);
or U1983 (N_1983,N_1779,N_1264);
xnor U1984 (N_1984,N_1573,N_1258);
nor U1985 (N_1985,N_1384,N_1570);
or U1986 (N_1986,N_1331,N_1420);
or U1987 (N_1987,N_1490,N_1494);
xor U1988 (N_1988,N_1638,N_1691);
xor U1989 (N_1989,N_1342,N_1397);
xnor U1990 (N_1990,N_1252,N_1699);
nand U1991 (N_1991,N_1374,N_1215);
nand U1992 (N_1992,N_1578,N_1353);
or U1993 (N_1993,N_1526,N_1396);
and U1994 (N_1994,N_1501,N_1524);
or U1995 (N_1995,N_1275,N_1257);
and U1996 (N_1996,N_1753,N_1563);
nand U1997 (N_1997,N_1759,N_1559);
nor U1998 (N_1998,N_1442,N_1568);
nor U1999 (N_1999,N_1541,N_1641);
nand U2000 (N_2000,N_1720,N_1725);
xnor U2001 (N_2001,N_1569,N_1408);
nand U2002 (N_2002,N_1597,N_1496);
nand U2003 (N_2003,N_1653,N_1272);
or U2004 (N_2004,N_1677,N_1572);
nand U2005 (N_2005,N_1204,N_1712);
nand U2006 (N_2006,N_1421,N_1506);
nor U2007 (N_2007,N_1492,N_1295);
nor U2008 (N_2008,N_1539,N_1560);
or U2009 (N_2009,N_1452,N_1288);
xor U2010 (N_2010,N_1702,N_1710);
or U2011 (N_2011,N_1660,N_1399);
or U2012 (N_2012,N_1634,N_1754);
xor U2013 (N_2013,N_1238,N_1301);
xor U2014 (N_2014,N_1428,N_1673);
and U2015 (N_2015,N_1644,N_1366);
xor U2016 (N_2016,N_1256,N_1751);
and U2017 (N_2017,N_1604,N_1413);
nand U2018 (N_2018,N_1659,N_1455);
nor U2019 (N_2019,N_1214,N_1212);
and U2020 (N_2020,N_1669,N_1241);
xor U2021 (N_2021,N_1683,N_1298);
or U2022 (N_2022,N_1639,N_1513);
nand U2023 (N_2023,N_1361,N_1322);
nand U2024 (N_2024,N_1207,N_1737);
xor U2025 (N_2025,N_1438,N_1363);
xor U2026 (N_2026,N_1273,N_1633);
or U2027 (N_2027,N_1243,N_1457);
nor U2028 (N_2028,N_1566,N_1336);
xor U2029 (N_2029,N_1631,N_1480);
xnor U2030 (N_2030,N_1310,N_1798);
nor U2031 (N_2031,N_1575,N_1728);
nor U2032 (N_2032,N_1461,N_1381);
nor U2033 (N_2033,N_1715,N_1333);
xor U2034 (N_2034,N_1648,N_1771);
xor U2035 (N_2035,N_1377,N_1741);
nand U2036 (N_2036,N_1482,N_1370);
nor U2037 (N_2037,N_1586,N_1267);
nand U2038 (N_2038,N_1675,N_1436);
nand U2039 (N_2039,N_1440,N_1330);
xor U2040 (N_2040,N_1349,N_1595);
and U2041 (N_2041,N_1498,N_1621);
nor U2042 (N_2042,N_1661,N_1379);
and U2043 (N_2043,N_1360,N_1642);
or U2044 (N_2044,N_1407,N_1224);
and U2045 (N_2045,N_1766,N_1706);
or U2046 (N_2046,N_1223,N_1418);
xor U2047 (N_2047,N_1355,N_1509);
nor U2048 (N_2048,N_1626,N_1775);
and U2049 (N_2049,N_1249,N_1210);
or U2050 (N_2050,N_1614,N_1785);
nand U2051 (N_2051,N_1383,N_1484);
xor U2052 (N_2052,N_1697,N_1645);
or U2053 (N_2053,N_1369,N_1576);
xnor U2054 (N_2054,N_1348,N_1769);
nand U2055 (N_2055,N_1532,N_1615);
and U2056 (N_2056,N_1400,N_1388);
nor U2057 (N_2057,N_1316,N_1605);
nand U2058 (N_2058,N_1343,N_1237);
xnor U2059 (N_2059,N_1551,N_1234);
xor U2060 (N_2060,N_1422,N_1456);
and U2061 (N_2061,N_1253,N_1357);
nor U2062 (N_2062,N_1758,N_1244);
nand U2063 (N_2063,N_1600,N_1287);
xor U2064 (N_2064,N_1463,N_1540);
or U2065 (N_2065,N_1628,N_1517);
nor U2066 (N_2066,N_1424,N_1556);
nand U2067 (N_2067,N_1450,N_1776);
nand U2068 (N_2068,N_1305,N_1544);
xnor U2069 (N_2069,N_1266,N_1548);
or U2070 (N_2070,N_1416,N_1740);
nor U2071 (N_2071,N_1735,N_1326);
or U2072 (N_2072,N_1248,N_1552);
nor U2073 (N_2073,N_1389,N_1757);
nand U2074 (N_2074,N_1760,N_1647);
and U2075 (N_2075,N_1294,N_1398);
nor U2076 (N_2076,N_1770,N_1799);
xor U2077 (N_2077,N_1579,N_1666);
nand U2078 (N_2078,N_1561,N_1716);
or U2079 (N_2079,N_1250,N_1415);
or U2080 (N_2080,N_1468,N_1709);
or U2081 (N_2081,N_1317,N_1203);
nor U2082 (N_2082,N_1296,N_1607);
nand U2083 (N_2083,N_1479,N_1435);
nand U2084 (N_2084,N_1500,N_1405);
or U2085 (N_2085,N_1290,N_1327);
nor U2086 (N_2086,N_1448,N_1743);
or U2087 (N_2087,N_1791,N_1656);
or U2088 (N_2088,N_1676,N_1554);
nor U2089 (N_2089,N_1274,N_1534);
nand U2090 (N_2090,N_1533,N_1392);
nor U2091 (N_2091,N_1582,N_1481);
and U2092 (N_2092,N_1546,N_1265);
or U2093 (N_2093,N_1318,N_1598);
nand U2094 (N_2094,N_1262,N_1497);
nor U2095 (N_2095,N_1402,N_1414);
and U2096 (N_2096,N_1302,N_1708);
nor U2097 (N_2097,N_1202,N_1299);
and U2098 (N_2098,N_1499,N_1778);
xor U2099 (N_2099,N_1788,N_1618);
nor U2100 (N_2100,N_1474,N_1243);
xnor U2101 (N_2101,N_1465,N_1434);
xnor U2102 (N_2102,N_1278,N_1409);
and U2103 (N_2103,N_1522,N_1277);
and U2104 (N_2104,N_1797,N_1610);
and U2105 (N_2105,N_1263,N_1638);
xor U2106 (N_2106,N_1204,N_1399);
and U2107 (N_2107,N_1393,N_1254);
nand U2108 (N_2108,N_1289,N_1386);
or U2109 (N_2109,N_1359,N_1749);
or U2110 (N_2110,N_1263,N_1556);
nor U2111 (N_2111,N_1285,N_1659);
xor U2112 (N_2112,N_1793,N_1342);
and U2113 (N_2113,N_1415,N_1352);
or U2114 (N_2114,N_1403,N_1766);
nand U2115 (N_2115,N_1744,N_1562);
or U2116 (N_2116,N_1247,N_1385);
nor U2117 (N_2117,N_1474,N_1700);
and U2118 (N_2118,N_1529,N_1590);
xnor U2119 (N_2119,N_1705,N_1345);
and U2120 (N_2120,N_1529,N_1654);
nor U2121 (N_2121,N_1441,N_1236);
xor U2122 (N_2122,N_1216,N_1489);
and U2123 (N_2123,N_1715,N_1615);
xor U2124 (N_2124,N_1358,N_1503);
nand U2125 (N_2125,N_1407,N_1274);
and U2126 (N_2126,N_1297,N_1575);
nand U2127 (N_2127,N_1767,N_1393);
nand U2128 (N_2128,N_1687,N_1622);
or U2129 (N_2129,N_1619,N_1284);
or U2130 (N_2130,N_1724,N_1233);
nor U2131 (N_2131,N_1431,N_1419);
or U2132 (N_2132,N_1436,N_1793);
or U2133 (N_2133,N_1419,N_1788);
nand U2134 (N_2134,N_1576,N_1454);
or U2135 (N_2135,N_1629,N_1207);
or U2136 (N_2136,N_1591,N_1795);
xnor U2137 (N_2137,N_1618,N_1651);
nand U2138 (N_2138,N_1520,N_1503);
or U2139 (N_2139,N_1735,N_1758);
or U2140 (N_2140,N_1630,N_1779);
and U2141 (N_2141,N_1695,N_1372);
nor U2142 (N_2142,N_1688,N_1287);
or U2143 (N_2143,N_1763,N_1713);
or U2144 (N_2144,N_1760,N_1676);
xor U2145 (N_2145,N_1633,N_1593);
or U2146 (N_2146,N_1613,N_1461);
or U2147 (N_2147,N_1797,N_1303);
nand U2148 (N_2148,N_1442,N_1319);
xnor U2149 (N_2149,N_1578,N_1274);
and U2150 (N_2150,N_1660,N_1402);
xnor U2151 (N_2151,N_1652,N_1499);
and U2152 (N_2152,N_1633,N_1613);
and U2153 (N_2153,N_1562,N_1549);
or U2154 (N_2154,N_1573,N_1537);
nor U2155 (N_2155,N_1697,N_1710);
or U2156 (N_2156,N_1799,N_1630);
and U2157 (N_2157,N_1570,N_1408);
nand U2158 (N_2158,N_1230,N_1777);
xnor U2159 (N_2159,N_1328,N_1224);
and U2160 (N_2160,N_1508,N_1538);
xor U2161 (N_2161,N_1300,N_1256);
nand U2162 (N_2162,N_1243,N_1536);
nand U2163 (N_2163,N_1348,N_1482);
xnor U2164 (N_2164,N_1397,N_1408);
or U2165 (N_2165,N_1661,N_1792);
and U2166 (N_2166,N_1544,N_1610);
xnor U2167 (N_2167,N_1219,N_1252);
nor U2168 (N_2168,N_1301,N_1440);
xor U2169 (N_2169,N_1420,N_1656);
or U2170 (N_2170,N_1613,N_1417);
or U2171 (N_2171,N_1641,N_1750);
nand U2172 (N_2172,N_1415,N_1697);
xor U2173 (N_2173,N_1577,N_1392);
nand U2174 (N_2174,N_1286,N_1369);
and U2175 (N_2175,N_1683,N_1360);
and U2176 (N_2176,N_1693,N_1255);
xor U2177 (N_2177,N_1379,N_1526);
xnor U2178 (N_2178,N_1675,N_1247);
nand U2179 (N_2179,N_1387,N_1578);
and U2180 (N_2180,N_1242,N_1224);
nor U2181 (N_2181,N_1719,N_1669);
nor U2182 (N_2182,N_1512,N_1247);
and U2183 (N_2183,N_1456,N_1359);
nor U2184 (N_2184,N_1539,N_1335);
xor U2185 (N_2185,N_1640,N_1712);
xnor U2186 (N_2186,N_1448,N_1570);
nand U2187 (N_2187,N_1282,N_1351);
nand U2188 (N_2188,N_1302,N_1714);
nand U2189 (N_2189,N_1643,N_1495);
or U2190 (N_2190,N_1317,N_1229);
xor U2191 (N_2191,N_1695,N_1525);
nor U2192 (N_2192,N_1598,N_1483);
nor U2193 (N_2193,N_1670,N_1673);
or U2194 (N_2194,N_1797,N_1239);
or U2195 (N_2195,N_1281,N_1234);
xor U2196 (N_2196,N_1774,N_1617);
or U2197 (N_2197,N_1260,N_1255);
nor U2198 (N_2198,N_1433,N_1723);
xor U2199 (N_2199,N_1405,N_1417);
xor U2200 (N_2200,N_1300,N_1613);
nor U2201 (N_2201,N_1513,N_1442);
or U2202 (N_2202,N_1389,N_1500);
and U2203 (N_2203,N_1283,N_1214);
and U2204 (N_2204,N_1489,N_1533);
nor U2205 (N_2205,N_1393,N_1203);
or U2206 (N_2206,N_1388,N_1619);
and U2207 (N_2207,N_1646,N_1497);
nor U2208 (N_2208,N_1276,N_1411);
nand U2209 (N_2209,N_1738,N_1596);
nor U2210 (N_2210,N_1283,N_1410);
and U2211 (N_2211,N_1230,N_1299);
xor U2212 (N_2212,N_1472,N_1390);
or U2213 (N_2213,N_1521,N_1522);
nand U2214 (N_2214,N_1577,N_1201);
or U2215 (N_2215,N_1705,N_1206);
xnor U2216 (N_2216,N_1252,N_1512);
xor U2217 (N_2217,N_1329,N_1644);
and U2218 (N_2218,N_1426,N_1754);
or U2219 (N_2219,N_1553,N_1363);
nand U2220 (N_2220,N_1390,N_1381);
and U2221 (N_2221,N_1760,N_1548);
and U2222 (N_2222,N_1365,N_1284);
nor U2223 (N_2223,N_1221,N_1795);
and U2224 (N_2224,N_1267,N_1718);
nor U2225 (N_2225,N_1458,N_1252);
nor U2226 (N_2226,N_1355,N_1784);
or U2227 (N_2227,N_1778,N_1375);
nor U2228 (N_2228,N_1383,N_1378);
and U2229 (N_2229,N_1278,N_1431);
nor U2230 (N_2230,N_1510,N_1319);
nor U2231 (N_2231,N_1606,N_1332);
xnor U2232 (N_2232,N_1631,N_1237);
nor U2233 (N_2233,N_1676,N_1790);
xnor U2234 (N_2234,N_1372,N_1486);
xor U2235 (N_2235,N_1334,N_1378);
xnor U2236 (N_2236,N_1580,N_1230);
xor U2237 (N_2237,N_1769,N_1291);
and U2238 (N_2238,N_1258,N_1456);
and U2239 (N_2239,N_1274,N_1564);
or U2240 (N_2240,N_1426,N_1690);
xor U2241 (N_2241,N_1769,N_1780);
nor U2242 (N_2242,N_1545,N_1384);
and U2243 (N_2243,N_1341,N_1634);
and U2244 (N_2244,N_1246,N_1300);
nand U2245 (N_2245,N_1347,N_1522);
nand U2246 (N_2246,N_1456,N_1467);
xor U2247 (N_2247,N_1393,N_1538);
nand U2248 (N_2248,N_1331,N_1501);
or U2249 (N_2249,N_1633,N_1563);
or U2250 (N_2250,N_1763,N_1362);
xnor U2251 (N_2251,N_1571,N_1445);
and U2252 (N_2252,N_1654,N_1599);
nand U2253 (N_2253,N_1208,N_1458);
and U2254 (N_2254,N_1715,N_1655);
xor U2255 (N_2255,N_1719,N_1412);
and U2256 (N_2256,N_1242,N_1577);
or U2257 (N_2257,N_1572,N_1489);
nor U2258 (N_2258,N_1709,N_1737);
nor U2259 (N_2259,N_1418,N_1310);
xor U2260 (N_2260,N_1630,N_1485);
nand U2261 (N_2261,N_1380,N_1720);
xnor U2262 (N_2262,N_1371,N_1769);
nand U2263 (N_2263,N_1227,N_1589);
or U2264 (N_2264,N_1792,N_1428);
nand U2265 (N_2265,N_1473,N_1526);
nand U2266 (N_2266,N_1437,N_1632);
nor U2267 (N_2267,N_1234,N_1586);
and U2268 (N_2268,N_1341,N_1481);
or U2269 (N_2269,N_1599,N_1619);
and U2270 (N_2270,N_1255,N_1342);
nand U2271 (N_2271,N_1551,N_1662);
or U2272 (N_2272,N_1650,N_1298);
and U2273 (N_2273,N_1630,N_1266);
xor U2274 (N_2274,N_1463,N_1323);
nand U2275 (N_2275,N_1524,N_1205);
or U2276 (N_2276,N_1556,N_1461);
and U2277 (N_2277,N_1436,N_1294);
xor U2278 (N_2278,N_1658,N_1218);
and U2279 (N_2279,N_1783,N_1317);
nand U2280 (N_2280,N_1361,N_1502);
nand U2281 (N_2281,N_1650,N_1739);
nand U2282 (N_2282,N_1391,N_1333);
nand U2283 (N_2283,N_1598,N_1510);
and U2284 (N_2284,N_1490,N_1226);
nand U2285 (N_2285,N_1362,N_1639);
xor U2286 (N_2286,N_1388,N_1416);
or U2287 (N_2287,N_1528,N_1509);
xor U2288 (N_2288,N_1279,N_1381);
xnor U2289 (N_2289,N_1222,N_1572);
nor U2290 (N_2290,N_1201,N_1425);
xor U2291 (N_2291,N_1291,N_1599);
and U2292 (N_2292,N_1517,N_1243);
and U2293 (N_2293,N_1280,N_1636);
and U2294 (N_2294,N_1526,N_1748);
nand U2295 (N_2295,N_1280,N_1508);
nand U2296 (N_2296,N_1245,N_1406);
nand U2297 (N_2297,N_1207,N_1599);
nand U2298 (N_2298,N_1737,N_1747);
nor U2299 (N_2299,N_1691,N_1258);
and U2300 (N_2300,N_1797,N_1475);
nor U2301 (N_2301,N_1781,N_1351);
xnor U2302 (N_2302,N_1547,N_1730);
and U2303 (N_2303,N_1319,N_1670);
and U2304 (N_2304,N_1235,N_1385);
or U2305 (N_2305,N_1461,N_1318);
nor U2306 (N_2306,N_1471,N_1450);
or U2307 (N_2307,N_1302,N_1416);
xor U2308 (N_2308,N_1766,N_1778);
and U2309 (N_2309,N_1280,N_1710);
nor U2310 (N_2310,N_1338,N_1616);
nand U2311 (N_2311,N_1553,N_1799);
or U2312 (N_2312,N_1565,N_1685);
nand U2313 (N_2313,N_1203,N_1737);
nand U2314 (N_2314,N_1314,N_1656);
xor U2315 (N_2315,N_1501,N_1610);
and U2316 (N_2316,N_1366,N_1298);
or U2317 (N_2317,N_1218,N_1562);
nand U2318 (N_2318,N_1377,N_1388);
nand U2319 (N_2319,N_1485,N_1388);
xor U2320 (N_2320,N_1478,N_1201);
and U2321 (N_2321,N_1799,N_1558);
nor U2322 (N_2322,N_1772,N_1396);
nand U2323 (N_2323,N_1499,N_1530);
and U2324 (N_2324,N_1399,N_1727);
or U2325 (N_2325,N_1524,N_1779);
or U2326 (N_2326,N_1787,N_1587);
and U2327 (N_2327,N_1382,N_1785);
and U2328 (N_2328,N_1589,N_1441);
xnor U2329 (N_2329,N_1737,N_1497);
or U2330 (N_2330,N_1516,N_1327);
or U2331 (N_2331,N_1744,N_1460);
nor U2332 (N_2332,N_1227,N_1588);
xnor U2333 (N_2333,N_1422,N_1655);
or U2334 (N_2334,N_1499,N_1592);
xor U2335 (N_2335,N_1766,N_1313);
xnor U2336 (N_2336,N_1611,N_1449);
xnor U2337 (N_2337,N_1634,N_1667);
nand U2338 (N_2338,N_1655,N_1447);
and U2339 (N_2339,N_1716,N_1398);
or U2340 (N_2340,N_1435,N_1691);
xnor U2341 (N_2341,N_1738,N_1301);
xor U2342 (N_2342,N_1607,N_1527);
xnor U2343 (N_2343,N_1528,N_1289);
or U2344 (N_2344,N_1460,N_1599);
nor U2345 (N_2345,N_1386,N_1498);
xnor U2346 (N_2346,N_1460,N_1536);
or U2347 (N_2347,N_1690,N_1511);
nand U2348 (N_2348,N_1561,N_1599);
nor U2349 (N_2349,N_1636,N_1575);
or U2350 (N_2350,N_1714,N_1255);
nand U2351 (N_2351,N_1357,N_1260);
or U2352 (N_2352,N_1679,N_1595);
or U2353 (N_2353,N_1310,N_1507);
nand U2354 (N_2354,N_1257,N_1681);
or U2355 (N_2355,N_1222,N_1254);
nand U2356 (N_2356,N_1385,N_1492);
and U2357 (N_2357,N_1280,N_1359);
and U2358 (N_2358,N_1736,N_1205);
nor U2359 (N_2359,N_1790,N_1485);
and U2360 (N_2360,N_1341,N_1353);
xnor U2361 (N_2361,N_1258,N_1637);
or U2362 (N_2362,N_1452,N_1387);
and U2363 (N_2363,N_1605,N_1208);
and U2364 (N_2364,N_1335,N_1295);
nor U2365 (N_2365,N_1467,N_1636);
nand U2366 (N_2366,N_1577,N_1304);
and U2367 (N_2367,N_1262,N_1279);
and U2368 (N_2368,N_1422,N_1616);
nand U2369 (N_2369,N_1678,N_1654);
xnor U2370 (N_2370,N_1340,N_1780);
xnor U2371 (N_2371,N_1581,N_1363);
nand U2372 (N_2372,N_1759,N_1554);
nand U2373 (N_2373,N_1736,N_1480);
or U2374 (N_2374,N_1603,N_1456);
or U2375 (N_2375,N_1307,N_1326);
or U2376 (N_2376,N_1633,N_1773);
and U2377 (N_2377,N_1400,N_1510);
and U2378 (N_2378,N_1246,N_1519);
and U2379 (N_2379,N_1432,N_1424);
and U2380 (N_2380,N_1258,N_1771);
nand U2381 (N_2381,N_1623,N_1547);
and U2382 (N_2382,N_1534,N_1284);
nor U2383 (N_2383,N_1462,N_1697);
or U2384 (N_2384,N_1584,N_1368);
and U2385 (N_2385,N_1589,N_1712);
nor U2386 (N_2386,N_1223,N_1444);
xnor U2387 (N_2387,N_1215,N_1613);
nand U2388 (N_2388,N_1472,N_1260);
nand U2389 (N_2389,N_1519,N_1438);
nor U2390 (N_2390,N_1696,N_1296);
and U2391 (N_2391,N_1714,N_1434);
xnor U2392 (N_2392,N_1454,N_1615);
and U2393 (N_2393,N_1280,N_1492);
xor U2394 (N_2394,N_1678,N_1230);
nor U2395 (N_2395,N_1654,N_1629);
nand U2396 (N_2396,N_1286,N_1359);
or U2397 (N_2397,N_1780,N_1348);
and U2398 (N_2398,N_1487,N_1775);
or U2399 (N_2399,N_1757,N_1292);
xor U2400 (N_2400,N_2217,N_2308);
xor U2401 (N_2401,N_2231,N_1991);
nand U2402 (N_2402,N_2198,N_2366);
nand U2403 (N_2403,N_2139,N_2383);
nand U2404 (N_2404,N_1926,N_1811);
xor U2405 (N_2405,N_2253,N_2149);
nand U2406 (N_2406,N_2173,N_1843);
and U2407 (N_2407,N_2057,N_2098);
nand U2408 (N_2408,N_2014,N_1817);
or U2409 (N_2409,N_2386,N_1890);
nor U2410 (N_2410,N_1831,N_2189);
nand U2411 (N_2411,N_1921,N_2232);
nand U2412 (N_2412,N_1813,N_2262);
and U2413 (N_2413,N_1964,N_2355);
and U2414 (N_2414,N_1875,N_2134);
nor U2415 (N_2415,N_1878,N_2390);
and U2416 (N_2416,N_1854,N_1844);
nor U2417 (N_2417,N_2279,N_1877);
nor U2418 (N_2418,N_2342,N_2181);
nor U2419 (N_2419,N_2011,N_1975);
nand U2420 (N_2420,N_2353,N_2347);
and U2421 (N_2421,N_1856,N_1892);
nor U2422 (N_2422,N_2377,N_2058);
or U2423 (N_2423,N_2184,N_2106);
or U2424 (N_2424,N_1942,N_2395);
and U2425 (N_2425,N_2305,N_2091);
and U2426 (N_2426,N_1818,N_2048);
nand U2427 (N_2427,N_2238,N_2041);
nand U2428 (N_2428,N_1901,N_1963);
and U2429 (N_2429,N_2274,N_2102);
xor U2430 (N_2430,N_1951,N_2154);
and U2431 (N_2431,N_2079,N_2157);
nand U2432 (N_2432,N_2069,N_1873);
nand U2433 (N_2433,N_2151,N_2278);
nor U2434 (N_2434,N_2153,N_2172);
nor U2435 (N_2435,N_2197,N_1931);
xnor U2436 (N_2436,N_1803,N_2247);
and U2437 (N_2437,N_2280,N_2376);
or U2438 (N_2438,N_2375,N_2191);
nand U2439 (N_2439,N_2371,N_1801);
or U2440 (N_2440,N_1816,N_2019);
or U2441 (N_2441,N_2257,N_2175);
nor U2442 (N_2442,N_1809,N_1893);
xnor U2443 (N_2443,N_2169,N_2147);
nand U2444 (N_2444,N_2334,N_2290);
xor U2445 (N_2445,N_1895,N_2382);
or U2446 (N_2446,N_2391,N_2089);
nor U2447 (N_2447,N_1968,N_1995);
and U2448 (N_2448,N_1955,N_2165);
xnor U2449 (N_2449,N_2204,N_1940);
nand U2450 (N_2450,N_1967,N_2267);
xor U2451 (N_2451,N_1832,N_2252);
xor U2452 (N_2452,N_2071,N_2365);
nand U2453 (N_2453,N_2150,N_2316);
and U2454 (N_2454,N_1861,N_1999);
nand U2455 (N_2455,N_2162,N_1851);
and U2456 (N_2456,N_2320,N_2061);
nand U2457 (N_2457,N_1922,N_2275);
nand U2458 (N_2458,N_1973,N_1910);
xor U2459 (N_2459,N_2276,N_1907);
nand U2460 (N_2460,N_2369,N_1947);
or U2461 (N_2461,N_2055,N_2009);
xnor U2462 (N_2462,N_2380,N_1938);
nand U2463 (N_2463,N_1885,N_1883);
or U2464 (N_2464,N_1996,N_2078);
nor U2465 (N_2465,N_2260,N_1905);
or U2466 (N_2466,N_2345,N_2220);
nand U2467 (N_2467,N_2392,N_1962);
nand U2468 (N_2468,N_2287,N_2319);
nor U2469 (N_2469,N_1934,N_2285);
nor U2470 (N_2470,N_2143,N_1985);
nand U2471 (N_2471,N_1913,N_1992);
and U2472 (N_2472,N_2388,N_2022);
nand U2473 (N_2473,N_2114,N_2052);
nand U2474 (N_2474,N_2059,N_2393);
or U2475 (N_2475,N_1932,N_1966);
xor U2476 (N_2476,N_1810,N_2020);
nor U2477 (N_2477,N_2062,N_2180);
xnor U2478 (N_2478,N_2145,N_2115);
nor U2479 (N_2479,N_1916,N_2108);
or U2480 (N_2480,N_2167,N_1899);
and U2481 (N_2481,N_1859,N_1886);
or U2482 (N_2482,N_1912,N_1927);
nand U2483 (N_2483,N_1970,N_2178);
and U2484 (N_2484,N_2258,N_2211);
or U2485 (N_2485,N_2187,N_2292);
nand U2486 (N_2486,N_1949,N_2036);
nand U2487 (N_2487,N_2354,N_2083);
or U2488 (N_2488,N_2378,N_1808);
xor U2489 (N_2489,N_1945,N_2124);
and U2490 (N_2490,N_2360,N_2335);
nand U2491 (N_2491,N_1998,N_2337);
and U2492 (N_2492,N_2133,N_1882);
nand U2493 (N_2493,N_1952,N_2295);
xor U2494 (N_2494,N_1868,N_2268);
or U2495 (N_2495,N_2284,N_2381);
and U2496 (N_2496,N_1821,N_1853);
and U2497 (N_2497,N_2321,N_2081);
and U2498 (N_2498,N_2039,N_2343);
nand U2499 (N_2499,N_2200,N_2363);
and U2500 (N_2500,N_1911,N_1888);
and U2501 (N_2501,N_1954,N_2349);
nand U2502 (N_2502,N_2007,N_2113);
or U2503 (N_2503,N_2087,N_1880);
and U2504 (N_2504,N_1943,N_1879);
and U2505 (N_2505,N_1835,N_2293);
nand U2506 (N_2506,N_2140,N_1857);
and U2507 (N_2507,N_2196,N_1867);
xor U2508 (N_2508,N_2100,N_2065);
xor U2509 (N_2509,N_1953,N_2021);
and U2510 (N_2510,N_1976,N_2084);
xor U2511 (N_2511,N_1806,N_1978);
nor U2512 (N_2512,N_2384,N_1933);
nand U2513 (N_2513,N_1974,N_1830);
and U2514 (N_2514,N_2324,N_2156);
nand U2515 (N_2515,N_1815,N_2364);
xor U2516 (N_2516,N_2033,N_2026);
nor U2517 (N_2517,N_2005,N_2146);
nor U2518 (N_2518,N_2070,N_1827);
nand U2519 (N_2519,N_2088,N_2074);
xnor U2520 (N_2520,N_1812,N_2051);
xor U2521 (N_2521,N_1804,N_2199);
xor U2522 (N_2522,N_1900,N_1820);
xor U2523 (N_2523,N_2248,N_2346);
and U2524 (N_2524,N_2073,N_2245);
xor U2525 (N_2525,N_1928,N_2372);
nor U2526 (N_2526,N_2018,N_1863);
and U2527 (N_2527,N_2060,N_1889);
nand U2528 (N_2528,N_2277,N_2221);
nand U2529 (N_2529,N_2129,N_1935);
nor U2530 (N_2530,N_2194,N_2044);
nor U2531 (N_2531,N_2307,N_2313);
and U2532 (N_2532,N_2265,N_2125);
or U2533 (N_2533,N_2144,N_2101);
or U2534 (N_2534,N_2177,N_2155);
or U2535 (N_2535,N_2000,N_2077);
and U2536 (N_2536,N_2179,N_2336);
nor U2537 (N_2537,N_1979,N_2017);
or U2538 (N_2538,N_1860,N_2135);
xnor U2539 (N_2539,N_2362,N_1842);
or U2540 (N_2540,N_2242,N_2348);
and U2541 (N_2541,N_2104,N_2168);
and U2542 (N_2542,N_1884,N_1898);
nand U2543 (N_2543,N_2122,N_2214);
or U2544 (N_2544,N_2158,N_2288);
xor U2545 (N_2545,N_1891,N_2099);
xnor U2546 (N_2546,N_2357,N_2256);
xnor U2547 (N_2547,N_2255,N_2235);
or U2548 (N_2548,N_2182,N_1865);
nor U2549 (N_2549,N_1850,N_1838);
and U2550 (N_2550,N_2185,N_1959);
and U2551 (N_2551,N_1833,N_2207);
and U2552 (N_2552,N_1925,N_2210);
and U2553 (N_2553,N_2001,N_2298);
or U2554 (N_2554,N_2399,N_2086);
nand U2555 (N_2555,N_2269,N_2306);
and U2556 (N_2556,N_1987,N_2170);
nand U2557 (N_2557,N_2008,N_1841);
nand U2558 (N_2558,N_1814,N_1983);
xor U2559 (N_2559,N_2300,N_2118);
or U2560 (N_2560,N_1840,N_2034);
xnor U2561 (N_2561,N_2166,N_2224);
xor U2562 (N_2562,N_2358,N_1941);
or U2563 (N_2563,N_2367,N_1915);
or U2564 (N_2564,N_2037,N_2085);
xnor U2565 (N_2565,N_2107,N_2394);
or U2566 (N_2566,N_1969,N_2246);
nor U2567 (N_2567,N_2128,N_1896);
xnor U2568 (N_2568,N_2183,N_2186);
nand U2569 (N_2569,N_2216,N_2176);
and U2570 (N_2570,N_1872,N_1981);
and U2571 (N_2571,N_1960,N_2195);
and U2572 (N_2572,N_1936,N_2002);
and U2573 (N_2573,N_1870,N_2093);
nor U2574 (N_2574,N_2152,N_2031);
and U2575 (N_2575,N_2028,N_2063);
nand U2576 (N_2576,N_1887,N_2304);
or U2577 (N_2577,N_2236,N_2266);
nand U2578 (N_2578,N_2322,N_2035);
and U2579 (N_2579,N_2163,N_2132);
xor U2580 (N_2580,N_2315,N_2341);
xor U2581 (N_2581,N_2281,N_1972);
xor U2582 (N_2582,N_2301,N_2064);
or U2583 (N_2583,N_1946,N_1903);
nand U2584 (N_2584,N_1956,N_2309);
and U2585 (N_2585,N_1836,N_2229);
xor U2586 (N_2586,N_2126,N_2050);
or U2587 (N_2587,N_2286,N_1825);
and U2588 (N_2588,N_1852,N_2212);
or U2589 (N_2589,N_2303,N_2243);
xnor U2590 (N_2590,N_2328,N_2097);
nor U2591 (N_2591,N_2373,N_2352);
xor U2592 (N_2592,N_1894,N_1881);
nor U2593 (N_2593,N_1918,N_2080);
and U2594 (N_2594,N_2056,N_2318);
and U2595 (N_2595,N_1908,N_2263);
nor U2596 (N_2596,N_2092,N_2249);
or U2597 (N_2597,N_2234,N_2188);
nand U2598 (N_2598,N_2029,N_2379);
nand U2599 (N_2599,N_2270,N_2244);
or U2600 (N_2600,N_1997,N_1989);
and U2601 (N_2601,N_2006,N_2130);
xnor U2602 (N_2602,N_1802,N_2015);
nor U2603 (N_2603,N_1807,N_2117);
and U2604 (N_2604,N_2127,N_2094);
or U2605 (N_2605,N_1923,N_2013);
nand U2606 (N_2606,N_2103,N_2273);
xnor U2607 (N_2607,N_2161,N_2038);
or U2608 (N_2608,N_1937,N_1939);
or U2609 (N_2609,N_2174,N_2067);
and U2610 (N_2610,N_2202,N_2259);
nand U2611 (N_2611,N_1858,N_2047);
or U2612 (N_2612,N_2046,N_1822);
and U2613 (N_2613,N_2193,N_2333);
nand U2614 (N_2614,N_2356,N_2230);
or U2615 (N_2615,N_1862,N_1906);
nor U2616 (N_2616,N_2330,N_1965);
or U2617 (N_2617,N_1948,N_2398);
and U2618 (N_2618,N_1845,N_1839);
xor U2619 (N_2619,N_2283,N_2226);
nand U2620 (N_2620,N_2251,N_1977);
and U2621 (N_2621,N_2164,N_2136);
nand U2622 (N_2622,N_2331,N_1902);
or U2623 (N_2623,N_1826,N_2201);
nand U2624 (N_2624,N_2012,N_2314);
nor U2625 (N_2625,N_2312,N_2040);
xnor U2626 (N_2626,N_2302,N_2141);
nor U2627 (N_2627,N_2241,N_1950);
nor U2628 (N_2628,N_2205,N_1847);
and U2629 (N_2629,N_2049,N_2310);
nor U2630 (N_2630,N_1855,N_2327);
or U2631 (N_2631,N_1848,N_2219);
and U2632 (N_2632,N_1824,N_2192);
xor U2633 (N_2633,N_1930,N_2237);
xnor U2634 (N_2634,N_1904,N_2250);
xor U2635 (N_2635,N_2095,N_2209);
and U2636 (N_2636,N_2137,N_1819);
xor U2637 (N_2637,N_2329,N_2233);
nand U2638 (N_2638,N_1917,N_2032);
nor U2639 (N_2639,N_1961,N_2016);
and U2640 (N_2640,N_2206,N_2159);
nor U2641 (N_2641,N_2042,N_2385);
nand U2642 (N_2642,N_2344,N_1805);
nor U2643 (N_2643,N_1829,N_2054);
nor U2644 (N_2644,N_2361,N_1924);
nand U2645 (N_2645,N_2227,N_2350);
xor U2646 (N_2646,N_1846,N_1874);
nor U2647 (N_2647,N_2066,N_1909);
and U2648 (N_2648,N_2294,N_2389);
and U2649 (N_2649,N_2138,N_2082);
nor U2650 (N_2650,N_2203,N_2208);
and U2651 (N_2651,N_1984,N_2148);
nand U2652 (N_2652,N_2215,N_2326);
xnor U2653 (N_2653,N_2004,N_2374);
xor U2654 (N_2654,N_2296,N_2323);
nand U2655 (N_2655,N_2111,N_2239);
nor U2656 (N_2656,N_2272,N_1958);
xor U2657 (N_2657,N_1849,N_2339);
nor U2658 (N_2658,N_2396,N_1993);
nand U2659 (N_2659,N_1897,N_2223);
and U2660 (N_2660,N_2311,N_2332);
xor U2661 (N_2661,N_2075,N_2025);
nor U2662 (N_2662,N_1834,N_2387);
nand U2663 (N_2663,N_1828,N_2109);
or U2664 (N_2664,N_1919,N_2010);
nor U2665 (N_2665,N_2368,N_2116);
xor U2666 (N_2666,N_2090,N_2043);
xor U2667 (N_2667,N_1990,N_1876);
nand U2668 (N_2668,N_1914,N_2282);
nor U2669 (N_2669,N_2110,N_2160);
nand U2670 (N_2670,N_1980,N_2338);
nand U2671 (N_2671,N_2024,N_1944);
or U2672 (N_2672,N_1994,N_1871);
and U2673 (N_2673,N_1869,N_2351);
and U2674 (N_2674,N_1971,N_2254);
xor U2675 (N_2675,N_2027,N_1864);
nor U2676 (N_2676,N_2112,N_2119);
nand U2677 (N_2677,N_2213,N_2271);
and U2678 (N_2678,N_2023,N_1988);
xor U2679 (N_2679,N_2072,N_2190);
nand U2680 (N_2680,N_2121,N_1837);
or U2681 (N_2681,N_2370,N_2297);
nor U2682 (N_2682,N_2003,N_2045);
nor U2683 (N_2683,N_2359,N_1986);
nor U2684 (N_2684,N_2068,N_1929);
nor U2685 (N_2685,N_2225,N_2096);
or U2686 (N_2686,N_2120,N_2291);
xor U2687 (N_2687,N_2289,N_2131);
or U2688 (N_2688,N_2076,N_1866);
or U2689 (N_2689,N_2218,N_1823);
or U2690 (N_2690,N_2105,N_2261);
xor U2691 (N_2691,N_2030,N_1920);
or U2692 (N_2692,N_1957,N_2123);
or U2693 (N_2693,N_1982,N_2317);
xnor U2694 (N_2694,N_2397,N_2171);
nand U2695 (N_2695,N_2142,N_2222);
or U2696 (N_2696,N_1800,N_2264);
or U2697 (N_2697,N_2228,N_2299);
or U2698 (N_2698,N_2325,N_2240);
nand U2699 (N_2699,N_2340,N_2053);
xor U2700 (N_2700,N_2345,N_2255);
and U2701 (N_2701,N_2348,N_2363);
nand U2702 (N_2702,N_2179,N_2106);
or U2703 (N_2703,N_1984,N_1857);
nor U2704 (N_2704,N_1885,N_2223);
and U2705 (N_2705,N_1914,N_1959);
and U2706 (N_2706,N_2152,N_1909);
nand U2707 (N_2707,N_2280,N_2015);
or U2708 (N_2708,N_2369,N_2252);
nor U2709 (N_2709,N_2102,N_2248);
nor U2710 (N_2710,N_2076,N_2280);
nor U2711 (N_2711,N_2385,N_2073);
nor U2712 (N_2712,N_1837,N_1803);
nor U2713 (N_2713,N_1969,N_1922);
nor U2714 (N_2714,N_1945,N_1901);
nor U2715 (N_2715,N_2387,N_2277);
nor U2716 (N_2716,N_1933,N_2336);
nor U2717 (N_2717,N_2396,N_2102);
xor U2718 (N_2718,N_2298,N_2275);
and U2719 (N_2719,N_1869,N_1871);
nor U2720 (N_2720,N_2169,N_2160);
xnor U2721 (N_2721,N_2286,N_2295);
nand U2722 (N_2722,N_2049,N_2329);
nand U2723 (N_2723,N_2299,N_1891);
nor U2724 (N_2724,N_2214,N_1879);
nor U2725 (N_2725,N_2063,N_2040);
nand U2726 (N_2726,N_2214,N_2393);
or U2727 (N_2727,N_2098,N_1824);
nand U2728 (N_2728,N_2287,N_2220);
or U2729 (N_2729,N_1934,N_2359);
or U2730 (N_2730,N_2303,N_1934);
xnor U2731 (N_2731,N_2393,N_2051);
nor U2732 (N_2732,N_2314,N_2282);
nor U2733 (N_2733,N_1864,N_2076);
or U2734 (N_2734,N_1807,N_2012);
xnor U2735 (N_2735,N_2175,N_1814);
nand U2736 (N_2736,N_2199,N_2184);
xor U2737 (N_2737,N_2286,N_2011);
nand U2738 (N_2738,N_2030,N_2397);
nor U2739 (N_2739,N_1844,N_2005);
or U2740 (N_2740,N_1864,N_2186);
xor U2741 (N_2741,N_2183,N_2057);
nand U2742 (N_2742,N_2082,N_2316);
nand U2743 (N_2743,N_1807,N_2297);
nor U2744 (N_2744,N_2360,N_1952);
nand U2745 (N_2745,N_2071,N_2218);
nand U2746 (N_2746,N_2123,N_1828);
nor U2747 (N_2747,N_2199,N_2136);
nand U2748 (N_2748,N_1887,N_2378);
or U2749 (N_2749,N_2172,N_2268);
and U2750 (N_2750,N_2352,N_2253);
nor U2751 (N_2751,N_2257,N_2158);
xnor U2752 (N_2752,N_2064,N_1881);
and U2753 (N_2753,N_2294,N_1823);
xnor U2754 (N_2754,N_1814,N_1862);
or U2755 (N_2755,N_2398,N_2045);
xnor U2756 (N_2756,N_2178,N_2152);
or U2757 (N_2757,N_2043,N_2376);
xor U2758 (N_2758,N_2364,N_2155);
xor U2759 (N_2759,N_2248,N_1990);
nand U2760 (N_2760,N_2380,N_2394);
and U2761 (N_2761,N_2278,N_2338);
and U2762 (N_2762,N_1817,N_2175);
xor U2763 (N_2763,N_2352,N_2357);
nand U2764 (N_2764,N_2260,N_2174);
and U2765 (N_2765,N_2243,N_1935);
or U2766 (N_2766,N_2031,N_2093);
nand U2767 (N_2767,N_2077,N_2375);
nor U2768 (N_2768,N_1812,N_1905);
xnor U2769 (N_2769,N_2341,N_2079);
nor U2770 (N_2770,N_2374,N_2152);
nor U2771 (N_2771,N_1846,N_1937);
xor U2772 (N_2772,N_2155,N_2304);
xnor U2773 (N_2773,N_2390,N_2079);
and U2774 (N_2774,N_2073,N_2267);
xnor U2775 (N_2775,N_1849,N_2152);
nor U2776 (N_2776,N_1947,N_1861);
nor U2777 (N_2777,N_2084,N_2075);
nand U2778 (N_2778,N_2388,N_2195);
xor U2779 (N_2779,N_1970,N_2099);
nor U2780 (N_2780,N_2175,N_2054);
and U2781 (N_2781,N_1949,N_1852);
nand U2782 (N_2782,N_2387,N_1915);
nand U2783 (N_2783,N_2390,N_2168);
or U2784 (N_2784,N_2391,N_2229);
nand U2785 (N_2785,N_2149,N_2180);
xor U2786 (N_2786,N_2399,N_1965);
xor U2787 (N_2787,N_2048,N_2206);
or U2788 (N_2788,N_1972,N_2142);
nor U2789 (N_2789,N_2064,N_1868);
nor U2790 (N_2790,N_2392,N_1880);
or U2791 (N_2791,N_1998,N_2383);
or U2792 (N_2792,N_2042,N_2252);
or U2793 (N_2793,N_2285,N_1972);
or U2794 (N_2794,N_1820,N_2175);
xnor U2795 (N_2795,N_1834,N_2100);
or U2796 (N_2796,N_2338,N_2334);
and U2797 (N_2797,N_2307,N_2091);
xor U2798 (N_2798,N_2143,N_2044);
xnor U2799 (N_2799,N_2318,N_1890);
nor U2800 (N_2800,N_2135,N_1990);
nand U2801 (N_2801,N_1867,N_1900);
xor U2802 (N_2802,N_1988,N_2040);
or U2803 (N_2803,N_2235,N_2291);
xor U2804 (N_2804,N_2011,N_2038);
nor U2805 (N_2805,N_2398,N_1887);
nor U2806 (N_2806,N_1947,N_2182);
or U2807 (N_2807,N_2347,N_2366);
or U2808 (N_2808,N_1854,N_2218);
nand U2809 (N_2809,N_2377,N_1866);
xnor U2810 (N_2810,N_2044,N_2392);
or U2811 (N_2811,N_1884,N_1984);
or U2812 (N_2812,N_2127,N_1816);
and U2813 (N_2813,N_2064,N_2153);
and U2814 (N_2814,N_2340,N_2037);
xor U2815 (N_2815,N_1930,N_2351);
xor U2816 (N_2816,N_2356,N_2007);
and U2817 (N_2817,N_1908,N_2306);
xnor U2818 (N_2818,N_2064,N_2338);
and U2819 (N_2819,N_1915,N_2347);
xor U2820 (N_2820,N_2026,N_1911);
xor U2821 (N_2821,N_2051,N_2061);
nor U2822 (N_2822,N_2396,N_2160);
nor U2823 (N_2823,N_2227,N_1827);
and U2824 (N_2824,N_2158,N_1938);
and U2825 (N_2825,N_1969,N_1809);
xnor U2826 (N_2826,N_1921,N_1903);
and U2827 (N_2827,N_1819,N_1808);
xnor U2828 (N_2828,N_2067,N_1889);
xor U2829 (N_2829,N_2054,N_1934);
or U2830 (N_2830,N_2383,N_2318);
and U2831 (N_2831,N_2351,N_1982);
and U2832 (N_2832,N_1866,N_2036);
nor U2833 (N_2833,N_1839,N_2005);
xnor U2834 (N_2834,N_2224,N_2265);
or U2835 (N_2835,N_2167,N_2090);
nor U2836 (N_2836,N_2108,N_1941);
or U2837 (N_2837,N_2028,N_2196);
xor U2838 (N_2838,N_2018,N_2094);
xor U2839 (N_2839,N_1919,N_1806);
xnor U2840 (N_2840,N_2064,N_2213);
nand U2841 (N_2841,N_2321,N_2314);
and U2842 (N_2842,N_1839,N_2182);
nand U2843 (N_2843,N_2254,N_1845);
nand U2844 (N_2844,N_2202,N_2354);
and U2845 (N_2845,N_1875,N_2070);
nand U2846 (N_2846,N_1871,N_1947);
nand U2847 (N_2847,N_2371,N_2007);
xor U2848 (N_2848,N_2005,N_1833);
nor U2849 (N_2849,N_2201,N_1897);
nor U2850 (N_2850,N_2353,N_2124);
xor U2851 (N_2851,N_1823,N_1983);
nor U2852 (N_2852,N_1964,N_1948);
nand U2853 (N_2853,N_2321,N_2069);
xor U2854 (N_2854,N_2102,N_1839);
xor U2855 (N_2855,N_2241,N_2265);
nand U2856 (N_2856,N_1976,N_1998);
and U2857 (N_2857,N_1961,N_2142);
or U2858 (N_2858,N_1886,N_1823);
nand U2859 (N_2859,N_2330,N_2256);
nor U2860 (N_2860,N_2033,N_2364);
xor U2861 (N_2861,N_2237,N_2307);
nor U2862 (N_2862,N_2129,N_2316);
nor U2863 (N_2863,N_1847,N_1860);
and U2864 (N_2864,N_1979,N_2333);
and U2865 (N_2865,N_2287,N_2218);
or U2866 (N_2866,N_2048,N_1979);
xor U2867 (N_2867,N_1826,N_2356);
nand U2868 (N_2868,N_2070,N_2163);
nand U2869 (N_2869,N_2187,N_2096);
nand U2870 (N_2870,N_1999,N_1800);
and U2871 (N_2871,N_2021,N_1872);
nand U2872 (N_2872,N_2293,N_2092);
or U2873 (N_2873,N_2271,N_1986);
and U2874 (N_2874,N_2161,N_2104);
nor U2875 (N_2875,N_2275,N_1851);
and U2876 (N_2876,N_1991,N_1856);
and U2877 (N_2877,N_2354,N_2176);
nand U2878 (N_2878,N_1978,N_1850);
and U2879 (N_2879,N_1851,N_2114);
nor U2880 (N_2880,N_1911,N_2152);
xor U2881 (N_2881,N_2049,N_1811);
nor U2882 (N_2882,N_1886,N_1952);
or U2883 (N_2883,N_2293,N_1895);
nor U2884 (N_2884,N_2273,N_2374);
nor U2885 (N_2885,N_2118,N_2195);
or U2886 (N_2886,N_2241,N_2251);
nand U2887 (N_2887,N_1960,N_2144);
nor U2888 (N_2888,N_2004,N_2125);
xor U2889 (N_2889,N_2396,N_2268);
or U2890 (N_2890,N_1936,N_2086);
xor U2891 (N_2891,N_2211,N_2022);
and U2892 (N_2892,N_1810,N_2301);
and U2893 (N_2893,N_2256,N_2142);
nand U2894 (N_2894,N_2192,N_2130);
and U2895 (N_2895,N_2064,N_1802);
nand U2896 (N_2896,N_1952,N_2005);
nand U2897 (N_2897,N_2054,N_2071);
nand U2898 (N_2898,N_1829,N_2399);
nand U2899 (N_2899,N_2329,N_2288);
nand U2900 (N_2900,N_2241,N_2178);
or U2901 (N_2901,N_2134,N_2092);
nand U2902 (N_2902,N_2135,N_1919);
or U2903 (N_2903,N_2074,N_1906);
nand U2904 (N_2904,N_2385,N_1876);
and U2905 (N_2905,N_2127,N_1878);
and U2906 (N_2906,N_2120,N_1873);
xnor U2907 (N_2907,N_1985,N_1991);
nand U2908 (N_2908,N_2167,N_2136);
nand U2909 (N_2909,N_2300,N_2095);
and U2910 (N_2910,N_1850,N_2240);
and U2911 (N_2911,N_1939,N_2285);
and U2912 (N_2912,N_1824,N_2086);
nor U2913 (N_2913,N_2216,N_2088);
or U2914 (N_2914,N_2206,N_2094);
nor U2915 (N_2915,N_1876,N_2142);
nor U2916 (N_2916,N_2115,N_2385);
or U2917 (N_2917,N_1832,N_2028);
nor U2918 (N_2918,N_1990,N_1821);
or U2919 (N_2919,N_1908,N_2334);
and U2920 (N_2920,N_2311,N_2066);
nor U2921 (N_2921,N_2134,N_2232);
and U2922 (N_2922,N_2230,N_2311);
nor U2923 (N_2923,N_2044,N_2252);
xor U2924 (N_2924,N_2173,N_2018);
xnor U2925 (N_2925,N_2117,N_1995);
nor U2926 (N_2926,N_2339,N_2329);
nand U2927 (N_2927,N_1967,N_2182);
nor U2928 (N_2928,N_1926,N_2057);
nor U2929 (N_2929,N_1982,N_1842);
nor U2930 (N_2930,N_1955,N_2040);
and U2931 (N_2931,N_2136,N_2106);
xor U2932 (N_2932,N_2241,N_2051);
nand U2933 (N_2933,N_1908,N_1882);
nand U2934 (N_2934,N_2214,N_2207);
nor U2935 (N_2935,N_1917,N_2119);
nand U2936 (N_2936,N_2198,N_2244);
and U2937 (N_2937,N_1891,N_1953);
nor U2938 (N_2938,N_1919,N_2221);
or U2939 (N_2939,N_2174,N_2370);
nand U2940 (N_2940,N_2347,N_1859);
or U2941 (N_2941,N_2028,N_1922);
nand U2942 (N_2942,N_2309,N_1810);
nand U2943 (N_2943,N_2347,N_2078);
or U2944 (N_2944,N_2058,N_2239);
and U2945 (N_2945,N_1983,N_2297);
nor U2946 (N_2946,N_2302,N_2035);
nor U2947 (N_2947,N_2035,N_1962);
nor U2948 (N_2948,N_1962,N_2330);
nor U2949 (N_2949,N_2106,N_2293);
and U2950 (N_2950,N_1936,N_1900);
and U2951 (N_2951,N_2223,N_2229);
nor U2952 (N_2952,N_2364,N_2352);
xor U2953 (N_2953,N_2256,N_1915);
or U2954 (N_2954,N_1851,N_2058);
nand U2955 (N_2955,N_2247,N_2208);
nand U2956 (N_2956,N_1915,N_1824);
and U2957 (N_2957,N_2089,N_2141);
nor U2958 (N_2958,N_2275,N_2076);
or U2959 (N_2959,N_2305,N_2011);
xnor U2960 (N_2960,N_1906,N_1905);
nand U2961 (N_2961,N_1813,N_1928);
xor U2962 (N_2962,N_2372,N_1996);
or U2963 (N_2963,N_1876,N_1815);
nor U2964 (N_2964,N_1963,N_2387);
nor U2965 (N_2965,N_2195,N_2241);
or U2966 (N_2966,N_2382,N_2197);
nor U2967 (N_2967,N_1854,N_1804);
nand U2968 (N_2968,N_2236,N_2104);
nor U2969 (N_2969,N_1900,N_1952);
and U2970 (N_2970,N_2053,N_2326);
and U2971 (N_2971,N_1832,N_1867);
or U2972 (N_2972,N_1951,N_1804);
or U2973 (N_2973,N_1959,N_2387);
nand U2974 (N_2974,N_2112,N_2358);
or U2975 (N_2975,N_2059,N_1941);
or U2976 (N_2976,N_2092,N_2277);
nor U2977 (N_2977,N_2148,N_1925);
nor U2978 (N_2978,N_1917,N_1853);
nand U2979 (N_2979,N_2387,N_2120);
nor U2980 (N_2980,N_2371,N_1989);
nand U2981 (N_2981,N_2166,N_1859);
and U2982 (N_2982,N_1995,N_2207);
and U2983 (N_2983,N_1952,N_2064);
nand U2984 (N_2984,N_1800,N_2196);
nand U2985 (N_2985,N_2174,N_2232);
nand U2986 (N_2986,N_2381,N_2352);
nor U2987 (N_2987,N_2084,N_2338);
or U2988 (N_2988,N_1803,N_2070);
and U2989 (N_2989,N_2151,N_1976);
nand U2990 (N_2990,N_1899,N_2184);
nand U2991 (N_2991,N_2355,N_1956);
or U2992 (N_2992,N_1957,N_1915);
nor U2993 (N_2993,N_2228,N_2027);
xnor U2994 (N_2994,N_2203,N_2193);
or U2995 (N_2995,N_2204,N_2201);
and U2996 (N_2996,N_2339,N_2002);
nor U2997 (N_2997,N_2315,N_1852);
nor U2998 (N_2998,N_1833,N_2352);
xor U2999 (N_2999,N_2298,N_1977);
nand UO_0 (O_0,N_2460,N_2410);
nand UO_1 (O_1,N_2583,N_2720);
nor UO_2 (O_2,N_2826,N_2512);
nor UO_3 (O_3,N_2744,N_2992);
or UO_4 (O_4,N_2487,N_2730);
nand UO_5 (O_5,N_2932,N_2662);
nor UO_6 (O_6,N_2613,N_2641);
xnor UO_7 (O_7,N_2754,N_2937);
or UO_8 (O_8,N_2848,N_2742);
xnor UO_9 (O_9,N_2882,N_2820);
nor UO_10 (O_10,N_2698,N_2574);
and UO_11 (O_11,N_2614,N_2421);
or UO_12 (O_12,N_2483,N_2941);
and UO_13 (O_13,N_2639,N_2975);
and UO_14 (O_14,N_2624,N_2900);
nand UO_15 (O_15,N_2653,N_2973);
and UO_16 (O_16,N_2616,N_2474);
nand UO_17 (O_17,N_2701,N_2843);
nor UO_18 (O_18,N_2553,N_2737);
and UO_19 (O_19,N_2726,N_2417);
xnor UO_20 (O_20,N_2680,N_2849);
xnor UO_21 (O_21,N_2810,N_2665);
and UO_22 (O_22,N_2850,N_2441);
nand UO_23 (O_23,N_2444,N_2944);
and UO_24 (O_24,N_2567,N_2666);
and UO_25 (O_25,N_2696,N_2447);
or UO_26 (O_26,N_2904,N_2830);
xnor UO_27 (O_27,N_2418,N_2884);
xor UO_28 (O_28,N_2577,N_2437);
or UO_29 (O_29,N_2987,N_2805);
nand UO_30 (O_30,N_2797,N_2840);
or UO_31 (O_31,N_2670,N_2648);
nand UO_32 (O_32,N_2527,N_2606);
nand UO_33 (O_33,N_2546,N_2697);
nand UO_34 (O_34,N_2586,N_2446);
and UO_35 (O_35,N_2981,N_2617);
or UO_36 (O_36,N_2807,N_2828);
and UO_37 (O_37,N_2659,N_2627);
or UO_38 (O_38,N_2886,N_2986);
nand UO_39 (O_39,N_2675,N_2646);
and UO_40 (O_40,N_2596,N_2816);
and UO_41 (O_41,N_2424,N_2642);
or UO_42 (O_42,N_2651,N_2451);
nand UO_43 (O_43,N_2770,N_2762);
nor UO_44 (O_44,N_2456,N_2414);
nand UO_45 (O_45,N_2597,N_2803);
nand UO_46 (O_46,N_2764,N_2504);
nor UO_47 (O_47,N_2619,N_2589);
nand UO_48 (O_48,N_2857,N_2918);
xnor UO_49 (O_49,N_2746,N_2623);
nand UO_50 (O_50,N_2979,N_2528);
or UO_51 (O_51,N_2566,N_2591);
xnor UO_52 (O_52,N_2996,N_2711);
nand UO_53 (O_53,N_2479,N_2573);
and UO_54 (O_54,N_2893,N_2419);
xnor UO_55 (O_55,N_2561,N_2572);
nand UO_56 (O_56,N_2729,N_2459);
xnor UO_57 (O_57,N_2968,N_2916);
xor UO_58 (O_58,N_2773,N_2756);
nor UO_59 (O_59,N_2719,N_2743);
xnor UO_60 (O_60,N_2688,N_2673);
nand UO_61 (O_61,N_2600,N_2988);
xor UO_62 (O_62,N_2721,N_2535);
and UO_63 (O_63,N_2931,N_2819);
nand UO_64 (O_64,N_2611,N_2859);
nor UO_65 (O_65,N_2492,N_2576);
and UO_66 (O_66,N_2440,N_2488);
and UO_67 (O_67,N_2790,N_2838);
xor UO_68 (O_68,N_2707,N_2715);
and UO_69 (O_69,N_2782,N_2883);
nor UO_70 (O_70,N_2407,N_2581);
and UO_71 (O_71,N_2753,N_2485);
xnor UO_72 (O_72,N_2922,N_2984);
or UO_73 (O_73,N_2677,N_2868);
or UO_74 (O_74,N_2661,N_2808);
and UO_75 (O_75,N_2938,N_2925);
nor UO_76 (O_76,N_2693,N_2702);
nor UO_77 (O_77,N_2923,N_2584);
nand UO_78 (O_78,N_2558,N_2632);
nor UO_79 (O_79,N_2818,N_2860);
nand UO_80 (O_80,N_2575,N_2455);
nor UO_81 (O_81,N_2542,N_2888);
and UO_82 (O_82,N_2667,N_2953);
and UO_83 (O_83,N_2794,N_2433);
or UO_84 (O_84,N_2655,N_2491);
nand UO_85 (O_85,N_2590,N_2768);
xor UO_86 (O_86,N_2434,N_2432);
and UO_87 (O_87,N_2679,N_2517);
nand UO_88 (O_88,N_2921,N_2461);
xnor UO_89 (O_89,N_2554,N_2547);
nand UO_90 (O_90,N_2578,N_2962);
xor UO_91 (O_91,N_2842,N_2783);
xnor UO_92 (O_92,N_2776,N_2708);
nor UO_93 (O_93,N_2605,N_2524);
and UO_94 (O_94,N_2947,N_2431);
nor UO_95 (O_95,N_2626,N_2674);
and UO_96 (O_96,N_2462,N_2781);
xor UO_97 (O_97,N_2969,N_2587);
nor UO_98 (O_98,N_2750,N_2656);
or UO_99 (O_99,N_2465,N_2579);
and UO_100 (O_100,N_2891,N_2497);
and UO_101 (O_101,N_2668,N_2519);
xor UO_102 (O_102,N_2873,N_2531);
and UO_103 (O_103,N_2513,N_2847);
and UO_104 (O_104,N_2471,N_2683);
and UO_105 (O_105,N_2602,N_2735);
and UO_106 (O_106,N_2739,N_2878);
nor UO_107 (O_107,N_2714,N_2568);
nand UO_108 (O_108,N_2467,N_2695);
and UO_109 (O_109,N_2423,N_2952);
and UO_110 (O_110,N_2745,N_2644);
and UO_111 (O_111,N_2682,N_2700);
and UO_112 (O_112,N_2454,N_2967);
xor UO_113 (O_113,N_2871,N_2516);
and UO_114 (O_114,N_2425,N_2654);
nor UO_115 (O_115,N_2907,N_2989);
and UO_116 (O_116,N_2920,N_2400);
xnor UO_117 (O_117,N_2959,N_2955);
and UO_118 (O_118,N_2948,N_2951);
or UO_119 (O_119,N_2473,N_2469);
xor UO_120 (O_120,N_2525,N_2974);
and UO_121 (O_121,N_2551,N_2691);
and UO_122 (O_122,N_2747,N_2796);
or UO_123 (O_123,N_2408,N_2569);
xnor UO_124 (O_124,N_2669,N_2518);
xor UO_125 (O_125,N_2834,N_2995);
nor UO_126 (O_126,N_2464,N_2950);
or UO_127 (O_127,N_2502,N_2812);
xor UO_128 (O_128,N_2905,N_2647);
xor UO_129 (O_129,N_2936,N_2480);
and UO_130 (O_130,N_2887,N_2634);
xor UO_131 (O_131,N_2718,N_2486);
and UO_132 (O_132,N_2412,N_2692);
nand UO_133 (O_133,N_2580,N_2404);
nand UO_134 (O_134,N_2401,N_2710);
nand UO_135 (O_135,N_2983,N_2466);
or UO_136 (O_136,N_2875,N_2506);
and UO_137 (O_137,N_2443,N_2870);
nand UO_138 (O_138,N_2548,N_2570);
xnor UO_139 (O_139,N_2724,N_2510);
and UO_140 (O_140,N_2448,N_2601);
or UO_141 (O_141,N_2727,N_2571);
xor UO_142 (O_142,N_2604,N_2536);
nand UO_143 (O_143,N_2761,N_2452);
xor UO_144 (O_144,N_2766,N_2813);
nor UO_145 (O_145,N_2463,N_2684);
nand UO_146 (O_146,N_2458,N_2555);
or UO_147 (O_147,N_2612,N_2949);
and UO_148 (O_148,N_2993,N_2403);
nor UO_149 (O_149,N_2703,N_2978);
nor UO_150 (O_150,N_2935,N_2748);
or UO_151 (O_151,N_2685,N_2736);
xor UO_152 (O_152,N_2833,N_2911);
xor UO_153 (O_153,N_2643,N_2526);
or UO_154 (O_154,N_2765,N_2468);
nand UO_155 (O_155,N_2694,N_2402);
and UO_156 (O_156,N_2846,N_2522);
nor UO_157 (O_157,N_2560,N_2538);
nor UO_158 (O_158,N_2622,N_2476);
and UO_159 (O_159,N_2899,N_2484);
nor UO_160 (O_160,N_2505,N_2549);
and UO_161 (O_161,N_2477,N_2405);
nor UO_162 (O_162,N_2717,N_2759);
nor UO_163 (O_163,N_2752,N_2924);
and UO_164 (O_164,N_2785,N_2411);
nor UO_165 (O_165,N_2521,N_2844);
or UO_166 (O_166,N_2609,N_2852);
nor UO_167 (O_167,N_2652,N_2582);
nand UO_168 (O_168,N_2801,N_2919);
nor UO_169 (O_169,N_2544,N_2789);
and UO_170 (O_170,N_2503,N_2942);
nand UO_171 (O_171,N_2856,N_2442);
nand UO_172 (O_172,N_2982,N_2885);
nor UO_173 (O_173,N_2603,N_2814);
xnor UO_174 (O_174,N_2956,N_2788);
xnor UO_175 (O_175,N_2917,N_2489);
xor UO_176 (O_176,N_2908,N_2636);
nor UO_177 (O_177,N_2998,N_2915);
xor UO_178 (O_178,N_2585,N_2496);
and UO_179 (O_179,N_2775,N_2449);
and UO_180 (O_180,N_2903,N_2594);
nor UO_181 (O_181,N_2734,N_2564);
and UO_182 (O_182,N_2867,N_2645);
and UO_183 (O_183,N_2705,N_2427);
nor UO_184 (O_184,N_2927,N_2610);
and UO_185 (O_185,N_2621,N_2628);
or UO_186 (O_186,N_2879,N_2985);
nand UO_187 (O_187,N_2416,N_2649);
nor UO_188 (O_188,N_2749,N_2738);
and UO_189 (O_189,N_2615,N_2881);
xor UO_190 (O_190,N_2740,N_2533);
nand UO_191 (O_191,N_2787,N_2501);
xor UO_192 (O_192,N_2687,N_2934);
xnor UO_193 (O_193,N_2965,N_2650);
or UO_194 (O_194,N_2890,N_2997);
nor UO_195 (O_195,N_2543,N_2530);
and UO_196 (O_196,N_2663,N_2593);
and UO_197 (O_197,N_2629,N_2926);
or UO_198 (O_198,N_2539,N_2481);
nor UO_199 (O_199,N_2876,N_2631);
nor UO_200 (O_200,N_2990,N_2565);
or UO_201 (O_201,N_2757,N_2913);
nand UO_202 (O_202,N_2409,N_2957);
or UO_203 (O_203,N_2784,N_2709);
nand UO_204 (O_204,N_2798,N_2608);
and UO_205 (O_205,N_2836,N_2430);
or UO_206 (O_206,N_2971,N_2478);
nor UO_207 (O_207,N_2532,N_2865);
nor UO_208 (O_208,N_2943,N_2945);
xnor UO_209 (O_209,N_2827,N_2795);
or UO_210 (O_210,N_2874,N_2660);
and UO_211 (O_211,N_2620,N_2855);
xnor UO_212 (O_212,N_2723,N_2439);
nand UO_213 (O_213,N_2658,N_2495);
nand UO_214 (O_214,N_2450,N_2598);
and UO_215 (O_215,N_2896,N_2704);
and UO_216 (O_216,N_2595,N_2771);
nand UO_217 (O_217,N_2428,N_2777);
xor UO_218 (O_218,N_2638,N_2493);
and UO_219 (O_219,N_2824,N_2854);
nand UO_220 (O_220,N_2681,N_2438);
xor UO_221 (O_221,N_2537,N_2839);
or UO_222 (O_222,N_2509,N_2500);
xnor UO_223 (O_223,N_2457,N_2690);
or UO_224 (O_224,N_2961,N_2767);
nand UO_225 (O_225,N_2960,N_2637);
nand UO_226 (O_226,N_2545,N_2599);
xnor UO_227 (O_227,N_2898,N_2977);
and UO_228 (O_228,N_2625,N_2731);
or UO_229 (O_229,N_2760,N_2792);
and UO_230 (O_230,N_2712,N_2779);
or UO_231 (O_231,N_2832,N_2910);
and UO_232 (O_232,N_2678,N_2453);
nand UO_233 (O_233,N_2515,N_2954);
nand UO_234 (O_234,N_2445,N_2592);
nand UO_235 (O_235,N_2912,N_2413);
xnor UO_236 (O_236,N_2901,N_2906);
nor UO_237 (O_237,N_2494,N_2728);
or UO_238 (O_238,N_2817,N_2563);
nor UO_239 (O_239,N_2939,N_2499);
and UO_240 (O_240,N_2664,N_2804);
xnor UO_241 (O_241,N_2415,N_2894);
and UO_242 (O_242,N_2470,N_2799);
or UO_243 (O_243,N_2802,N_2822);
or UO_244 (O_244,N_2806,N_2507);
or UO_245 (O_245,N_2862,N_2793);
nand UO_246 (O_246,N_2825,N_2933);
and UO_247 (O_247,N_2588,N_2562);
nand UO_248 (O_248,N_2657,N_2841);
xor UO_249 (O_249,N_2902,N_2999);
or UO_250 (O_250,N_2809,N_2972);
nand UO_251 (O_251,N_2877,N_2406);
nor UO_252 (O_252,N_2863,N_2892);
nor UO_253 (O_253,N_2534,N_2895);
nor UO_254 (O_254,N_2672,N_2914);
nor UO_255 (O_255,N_2633,N_2897);
nand UO_256 (O_256,N_2861,N_2699);
nand UO_257 (O_257,N_2436,N_2940);
nand UO_258 (O_258,N_2786,N_2889);
or UO_259 (O_259,N_2800,N_2869);
nand UO_260 (O_260,N_2815,N_2929);
nand UO_261 (O_261,N_2559,N_2845);
nor UO_262 (O_262,N_2607,N_2853);
nand UO_263 (O_263,N_2426,N_2529);
or UO_264 (O_264,N_2640,N_2963);
nand UO_265 (O_265,N_2716,N_2970);
and UO_266 (O_266,N_2811,N_2964);
xnor UO_267 (O_267,N_2864,N_2722);
xnor UO_268 (O_268,N_2420,N_2732);
xnor UO_269 (O_269,N_2552,N_2872);
and UO_270 (O_270,N_2851,N_2994);
nor UO_271 (O_271,N_2958,N_2733);
nor UO_272 (O_272,N_2772,N_2966);
xor UO_273 (O_273,N_2676,N_2909);
nor UO_274 (O_274,N_2557,N_2508);
xnor UO_275 (O_275,N_2866,N_2751);
and UO_276 (O_276,N_2755,N_2778);
and UO_277 (O_277,N_2541,N_2689);
nand UO_278 (O_278,N_2550,N_2829);
or UO_279 (O_279,N_2422,N_2991);
and UO_280 (O_280,N_2429,N_2686);
and UO_281 (O_281,N_2490,N_2763);
nand UO_282 (O_282,N_2930,N_2540);
xnor UO_283 (O_283,N_2498,N_2725);
nand UO_284 (O_284,N_2706,N_2980);
nand UO_285 (O_285,N_2520,N_2858);
or UO_286 (O_286,N_2472,N_2523);
or UO_287 (O_287,N_2831,N_2741);
xor UO_288 (O_288,N_2758,N_2630);
xor UO_289 (O_289,N_2823,N_2671);
nor UO_290 (O_290,N_2511,N_2713);
or UO_291 (O_291,N_2514,N_2976);
nand UO_292 (O_292,N_2774,N_2482);
nand UO_293 (O_293,N_2769,N_2880);
nand UO_294 (O_294,N_2435,N_2837);
or UO_295 (O_295,N_2946,N_2780);
xnor UO_296 (O_296,N_2618,N_2475);
nor UO_297 (O_297,N_2635,N_2835);
xnor UO_298 (O_298,N_2556,N_2791);
nand UO_299 (O_299,N_2928,N_2821);
nand UO_300 (O_300,N_2518,N_2967);
nand UO_301 (O_301,N_2744,N_2991);
xor UO_302 (O_302,N_2674,N_2902);
nor UO_303 (O_303,N_2854,N_2590);
nand UO_304 (O_304,N_2456,N_2959);
nor UO_305 (O_305,N_2823,N_2897);
nand UO_306 (O_306,N_2785,N_2570);
xor UO_307 (O_307,N_2986,N_2947);
xnor UO_308 (O_308,N_2484,N_2905);
nand UO_309 (O_309,N_2448,N_2811);
or UO_310 (O_310,N_2972,N_2885);
nand UO_311 (O_311,N_2617,N_2462);
and UO_312 (O_312,N_2796,N_2639);
xor UO_313 (O_313,N_2547,N_2481);
or UO_314 (O_314,N_2832,N_2430);
xnor UO_315 (O_315,N_2855,N_2962);
xor UO_316 (O_316,N_2988,N_2405);
or UO_317 (O_317,N_2833,N_2661);
xnor UO_318 (O_318,N_2549,N_2808);
and UO_319 (O_319,N_2748,N_2644);
and UO_320 (O_320,N_2821,N_2777);
xor UO_321 (O_321,N_2769,N_2723);
or UO_322 (O_322,N_2427,N_2775);
or UO_323 (O_323,N_2965,N_2625);
and UO_324 (O_324,N_2466,N_2562);
or UO_325 (O_325,N_2686,N_2461);
nand UO_326 (O_326,N_2664,N_2491);
xor UO_327 (O_327,N_2707,N_2432);
or UO_328 (O_328,N_2990,N_2795);
xnor UO_329 (O_329,N_2444,N_2453);
xor UO_330 (O_330,N_2646,N_2558);
and UO_331 (O_331,N_2846,N_2619);
or UO_332 (O_332,N_2707,N_2847);
or UO_333 (O_333,N_2882,N_2488);
nand UO_334 (O_334,N_2706,N_2544);
or UO_335 (O_335,N_2836,N_2998);
nand UO_336 (O_336,N_2631,N_2605);
nor UO_337 (O_337,N_2586,N_2686);
nor UO_338 (O_338,N_2971,N_2558);
and UO_339 (O_339,N_2977,N_2954);
and UO_340 (O_340,N_2552,N_2702);
xor UO_341 (O_341,N_2475,N_2777);
or UO_342 (O_342,N_2417,N_2452);
xor UO_343 (O_343,N_2557,N_2593);
nand UO_344 (O_344,N_2733,N_2966);
xor UO_345 (O_345,N_2820,N_2790);
or UO_346 (O_346,N_2632,N_2486);
nand UO_347 (O_347,N_2586,N_2726);
nor UO_348 (O_348,N_2946,N_2586);
and UO_349 (O_349,N_2624,N_2857);
xor UO_350 (O_350,N_2858,N_2985);
or UO_351 (O_351,N_2503,N_2660);
xor UO_352 (O_352,N_2494,N_2712);
or UO_353 (O_353,N_2920,N_2818);
nor UO_354 (O_354,N_2918,N_2950);
nor UO_355 (O_355,N_2748,N_2463);
xnor UO_356 (O_356,N_2822,N_2473);
or UO_357 (O_357,N_2499,N_2830);
or UO_358 (O_358,N_2991,N_2863);
nand UO_359 (O_359,N_2830,N_2591);
and UO_360 (O_360,N_2427,N_2777);
nand UO_361 (O_361,N_2777,N_2745);
xnor UO_362 (O_362,N_2892,N_2458);
xor UO_363 (O_363,N_2619,N_2471);
or UO_364 (O_364,N_2630,N_2652);
and UO_365 (O_365,N_2634,N_2993);
nand UO_366 (O_366,N_2988,N_2712);
xnor UO_367 (O_367,N_2832,N_2588);
or UO_368 (O_368,N_2659,N_2658);
xor UO_369 (O_369,N_2442,N_2472);
xor UO_370 (O_370,N_2483,N_2725);
and UO_371 (O_371,N_2943,N_2724);
nand UO_372 (O_372,N_2999,N_2855);
nand UO_373 (O_373,N_2539,N_2635);
or UO_374 (O_374,N_2859,N_2772);
nor UO_375 (O_375,N_2414,N_2710);
nor UO_376 (O_376,N_2967,N_2627);
or UO_377 (O_377,N_2611,N_2989);
xnor UO_378 (O_378,N_2916,N_2953);
or UO_379 (O_379,N_2872,N_2589);
or UO_380 (O_380,N_2619,N_2935);
nor UO_381 (O_381,N_2482,N_2849);
nand UO_382 (O_382,N_2892,N_2864);
or UO_383 (O_383,N_2575,N_2743);
or UO_384 (O_384,N_2599,N_2738);
and UO_385 (O_385,N_2971,N_2910);
nand UO_386 (O_386,N_2796,N_2841);
xor UO_387 (O_387,N_2769,N_2450);
or UO_388 (O_388,N_2704,N_2638);
or UO_389 (O_389,N_2892,N_2968);
nand UO_390 (O_390,N_2551,N_2635);
nor UO_391 (O_391,N_2966,N_2472);
nor UO_392 (O_392,N_2678,N_2762);
nand UO_393 (O_393,N_2646,N_2766);
nand UO_394 (O_394,N_2808,N_2686);
xor UO_395 (O_395,N_2874,N_2610);
nor UO_396 (O_396,N_2639,N_2461);
and UO_397 (O_397,N_2820,N_2982);
xnor UO_398 (O_398,N_2580,N_2817);
nor UO_399 (O_399,N_2558,N_2908);
nand UO_400 (O_400,N_2935,N_2959);
or UO_401 (O_401,N_2413,N_2674);
or UO_402 (O_402,N_2673,N_2484);
and UO_403 (O_403,N_2924,N_2436);
nor UO_404 (O_404,N_2766,N_2980);
or UO_405 (O_405,N_2781,N_2734);
or UO_406 (O_406,N_2805,N_2604);
and UO_407 (O_407,N_2523,N_2530);
and UO_408 (O_408,N_2591,N_2813);
nor UO_409 (O_409,N_2841,N_2810);
or UO_410 (O_410,N_2834,N_2448);
xor UO_411 (O_411,N_2416,N_2991);
nand UO_412 (O_412,N_2586,N_2499);
nor UO_413 (O_413,N_2687,N_2953);
nor UO_414 (O_414,N_2891,N_2988);
or UO_415 (O_415,N_2794,N_2896);
xor UO_416 (O_416,N_2757,N_2952);
nor UO_417 (O_417,N_2913,N_2443);
xor UO_418 (O_418,N_2922,N_2787);
nor UO_419 (O_419,N_2885,N_2921);
xor UO_420 (O_420,N_2548,N_2550);
or UO_421 (O_421,N_2670,N_2429);
nand UO_422 (O_422,N_2854,N_2419);
or UO_423 (O_423,N_2867,N_2988);
and UO_424 (O_424,N_2703,N_2492);
or UO_425 (O_425,N_2989,N_2701);
nor UO_426 (O_426,N_2615,N_2523);
xnor UO_427 (O_427,N_2415,N_2677);
nand UO_428 (O_428,N_2971,N_2815);
and UO_429 (O_429,N_2522,N_2587);
xor UO_430 (O_430,N_2420,N_2474);
and UO_431 (O_431,N_2730,N_2738);
nor UO_432 (O_432,N_2666,N_2603);
xnor UO_433 (O_433,N_2551,N_2589);
xor UO_434 (O_434,N_2818,N_2555);
and UO_435 (O_435,N_2601,N_2600);
or UO_436 (O_436,N_2750,N_2971);
and UO_437 (O_437,N_2491,N_2615);
nor UO_438 (O_438,N_2999,N_2791);
nand UO_439 (O_439,N_2499,N_2537);
nand UO_440 (O_440,N_2478,N_2487);
or UO_441 (O_441,N_2439,N_2836);
or UO_442 (O_442,N_2740,N_2511);
xor UO_443 (O_443,N_2825,N_2732);
and UO_444 (O_444,N_2800,N_2753);
nand UO_445 (O_445,N_2672,N_2494);
xor UO_446 (O_446,N_2579,N_2473);
and UO_447 (O_447,N_2951,N_2436);
nand UO_448 (O_448,N_2740,N_2750);
xor UO_449 (O_449,N_2778,N_2548);
xor UO_450 (O_450,N_2932,N_2564);
nand UO_451 (O_451,N_2689,N_2440);
nor UO_452 (O_452,N_2656,N_2747);
or UO_453 (O_453,N_2417,N_2610);
and UO_454 (O_454,N_2552,N_2950);
and UO_455 (O_455,N_2490,N_2463);
xor UO_456 (O_456,N_2945,N_2573);
nand UO_457 (O_457,N_2831,N_2722);
or UO_458 (O_458,N_2964,N_2933);
nor UO_459 (O_459,N_2637,N_2766);
or UO_460 (O_460,N_2720,N_2445);
nand UO_461 (O_461,N_2400,N_2919);
or UO_462 (O_462,N_2891,N_2574);
nor UO_463 (O_463,N_2908,N_2408);
or UO_464 (O_464,N_2757,N_2796);
or UO_465 (O_465,N_2492,N_2433);
nor UO_466 (O_466,N_2725,N_2411);
and UO_467 (O_467,N_2404,N_2738);
or UO_468 (O_468,N_2744,N_2717);
nor UO_469 (O_469,N_2516,N_2676);
nor UO_470 (O_470,N_2526,N_2934);
nand UO_471 (O_471,N_2886,N_2642);
nor UO_472 (O_472,N_2597,N_2551);
xor UO_473 (O_473,N_2584,N_2800);
and UO_474 (O_474,N_2765,N_2432);
nor UO_475 (O_475,N_2520,N_2727);
or UO_476 (O_476,N_2772,N_2610);
or UO_477 (O_477,N_2911,N_2414);
xor UO_478 (O_478,N_2633,N_2760);
nor UO_479 (O_479,N_2813,N_2573);
xnor UO_480 (O_480,N_2471,N_2468);
or UO_481 (O_481,N_2582,N_2609);
nor UO_482 (O_482,N_2537,N_2557);
xnor UO_483 (O_483,N_2951,N_2449);
xor UO_484 (O_484,N_2517,N_2538);
nand UO_485 (O_485,N_2986,N_2581);
nor UO_486 (O_486,N_2819,N_2695);
and UO_487 (O_487,N_2907,N_2600);
xor UO_488 (O_488,N_2411,N_2465);
xnor UO_489 (O_489,N_2660,N_2804);
xnor UO_490 (O_490,N_2640,N_2767);
or UO_491 (O_491,N_2449,N_2468);
nor UO_492 (O_492,N_2931,N_2993);
nor UO_493 (O_493,N_2696,N_2666);
nand UO_494 (O_494,N_2481,N_2799);
xor UO_495 (O_495,N_2522,N_2641);
and UO_496 (O_496,N_2852,N_2503);
and UO_497 (O_497,N_2512,N_2915);
nor UO_498 (O_498,N_2832,N_2724);
nand UO_499 (O_499,N_2533,N_2919);
endmodule