module basic_1500_15000_2000_15_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1051,In_689);
nand U1 (N_1,In_1261,In_163);
xor U2 (N_2,In_363,In_1174);
or U3 (N_3,In_1415,In_41);
xor U4 (N_4,In_59,In_633);
xnor U5 (N_5,In_356,In_207);
xnor U6 (N_6,In_884,In_384);
nand U7 (N_7,In_201,In_1306);
or U8 (N_8,In_327,In_476);
nor U9 (N_9,In_1096,In_979);
or U10 (N_10,In_1316,In_686);
or U11 (N_11,In_974,In_1173);
or U12 (N_12,In_1387,In_1063);
xor U13 (N_13,In_562,In_194);
or U14 (N_14,In_944,In_752);
or U15 (N_15,In_1179,In_604);
and U16 (N_16,In_282,In_129);
xnor U17 (N_17,In_1374,In_116);
nor U18 (N_18,In_1206,In_1113);
and U19 (N_19,In_703,In_1246);
nor U20 (N_20,In_1403,In_925);
nor U21 (N_21,In_1477,In_1241);
nor U22 (N_22,In_205,In_1159);
nor U23 (N_23,In_71,In_948);
or U24 (N_24,In_447,In_533);
nor U25 (N_25,In_671,In_698);
nand U26 (N_26,In_861,In_910);
or U27 (N_27,In_240,In_783);
and U28 (N_28,In_1185,In_203);
nand U29 (N_29,In_836,In_1389);
nor U30 (N_30,In_1048,In_199);
or U31 (N_31,In_584,In_863);
nand U32 (N_32,In_955,In_1473);
and U33 (N_33,In_1238,In_426);
or U34 (N_34,In_1247,In_727);
and U35 (N_35,In_322,In_741);
nand U36 (N_36,In_543,In_1282);
and U37 (N_37,In_168,In_110);
xnor U38 (N_38,In_873,In_1266);
and U39 (N_39,In_311,In_184);
nand U40 (N_40,In_522,In_1050);
nor U41 (N_41,In_957,In_65);
nor U42 (N_42,In_745,In_758);
nand U43 (N_43,In_821,In_552);
or U44 (N_44,In_1423,In_331);
xor U45 (N_45,In_229,In_867);
xor U46 (N_46,In_937,In_467);
nor U47 (N_47,In_1053,In_993);
or U48 (N_48,In_764,In_888);
nand U49 (N_49,In_731,In_1449);
or U50 (N_50,In_1118,In_621);
nand U51 (N_51,In_870,In_411);
xnor U52 (N_52,In_958,In_720);
nand U53 (N_53,In_765,In_872);
or U54 (N_54,In_315,In_811);
nand U55 (N_55,In_923,In_302);
or U56 (N_56,In_1112,In_209);
nand U57 (N_57,In_674,In_1304);
xnor U58 (N_58,In_457,In_669);
nand U59 (N_59,In_1209,In_250);
nand U60 (N_60,In_593,In_1143);
xor U61 (N_61,In_1092,In_135);
or U62 (N_62,In_351,In_1401);
or U63 (N_63,In_657,In_241);
nand U64 (N_64,In_1452,In_337);
nor U65 (N_65,In_1071,In_865);
nor U66 (N_66,In_566,In_1386);
nor U67 (N_67,In_27,In_301);
nor U68 (N_68,In_477,In_653);
xor U69 (N_69,In_936,In_513);
and U70 (N_70,In_378,In_1407);
nand U71 (N_71,In_1091,In_596);
or U72 (N_72,In_625,In_432);
nand U73 (N_73,In_185,In_126);
nand U74 (N_74,In_1313,In_710);
nand U75 (N_75,In_261,In_51);
xor U76 (N_76,In_316,In_1464);
or U77 (N_77,In_749,In_128);
and U78 (N_78,In_733,In_1237);
and U79 (N_79,In_428,In_537);
or U80 (N_80,In_133,In_1084);
nor U81 (N_81,In_1479,In_1256);
nor U82 (N_82,In_1418,In_603);
xor U83 (N_83,In_975,In_855);
or U84 (N_84,In_862,In_670);
and U85 (N_85,In_568,In_355);
xnor U86 (N_86,In_608,In_375);
nor U87 (N_87,In_182,In_935);
nand U88 (N_88,In_1287,In_1055);
nand U89 (N_89,In_453,In_897);
nor U90 (N_90,In_732,In_187);
nor U91 (N_91,In_1229,In_1487);
xnor U92 (N_92,In_28,In_46);
nand U93 (N_93,In_524,In_359);
and U94 (N_94,In_946,In_858);
and U95 (N_95,In_723,In_1163);
or U96 (N_96,In_484,In_298);
nand U97 (N_97,In_730,In_415);
nor U98 (N_98,In_1139,In_407);
and U99 (N_99,In_1029,In_1130);
or U100 (N_100,In_532,In_488);
nor U101 (N_101,In_1413,In_1297);
nand U102 (N_102,In_124,In_228);
nand U103 (N_103,In_797,In_390);
and U104 (N_104,In_306,In_953);
or U105 (N_105,In_1003,In_440);
nor U106 (N_106,In_450,In_1170);
nand U107 (N_107,In_1002,In_553);
or U108 (N_108,In_950,In_58);
nand U109 (N_109,In_112,In_1052);
nand U110 (N_110,In_914,In_1150);
nor U111 (N_111,In_24,In_1450);
xnor U112 (N_112,In_1199,In_677);
and U113 (N_113,In_538,In_788);
or U114 (N_114,In_83,In_183);
xnor U115 (N_115,In_1392,In_586);
or U116 (N_116,In_1280,In_44);
and U117 (N_117,In_416,In_526);
nand U118 (N_118,In_399,In_820);
xnor U119 (N_119,In_414,In_62);
or U120 (N_120,In_857,In_683);
or U121 (N_121,In_1074,In_512);
nand U122 (N_122,In_273,In_1345);
xnor U123 (N_123,In_1484,In_728);
and U124 (N_124,In_1428,In_1176);
and U125 (N_125,In_1172,In_1189);
nor U126 (N_126,In_1146,In_577);
or U127 (N_127,In_1125,In_1250);
xor U128 (N_128,In_238,In_365);
nor U129 (N_129,In_1262,In_853);
nand U130 (N_130,In_1135,In_169);
xnor U131 (N_131,In_118,In_1134);
or U132 (N_132,In_518,In_827);
xor U133 (N_133,In_462,In_13);
and U134 (N_134,In_1362,In_708);
nor U135 (N_135,In_419,In_1033);
and U136 (N_136,In_259,In_368);
nor U137 (N_137,In_983,In_172);
xnor U138 (N_138,In_560,In_1308);
nor U139 (N_139,In_427,In_142);
or U140 (N_140,In_1400,In_1284);
or U141 (N_141,In_502,In_1106);
xnor U142 (N_142,In_381,In_490);
nand U143 (N_143,In_264,In_1167);
and U144 (N_144,In_304,In_812);
nor U145 (N_145,In_707,In_1412);
or U146 (N_146,In_180,In_1405);
or U147 (N_147,In_1375,In_81);
and U148 (N_148,In_808,In_104);
xnor U149 (N_149,In_1359,In_418);
and U150 (N_150,In_1142,In_191);
or U151 (N_151,In_1411,In_1398);
nor U152 (N_152,In_1433,In_511);
or U153 (N_153,In_1079,In_1217);
nand U154 (N_154,In_1164,In_482);
and U155 (N_155,In_206,In_179);
xor U156 (N_156,In_1393,In_1465);
xnor U157 (N_157,In_819,In_451);
xor U158 (N_158,In_449,In_1310);
nand U159 (N_159,In_1495,In_726);
nor U160 (N_160,In_1168,In_646);
or U161 (N_161,In_15,In_1026);
and U162 (N_162,In_1332,In_445);
or U163 (N_163,In_219,In_466);
and U164 (N_164,In_320,In_735);
nor U165 (N_165,In_739,In_523);
nor U166 (N_166,In_786,In_1093);
nor U167 (N_167,In_1388,In_1457);
xnor U168 (N_168,In_1348,In_1046);
xnor U169 (N_169,In_159,In_895);
nor U170 (N_170,In_1488,In_592);
nand U171 (N_171,In_3,In_117);
nor U172 (N_172,In_684,In_988);
or U173 (N_173,In_115,In_1132);
xor U174 (N_174,In_1335,In_297);
nand U175 (N_175,In_270,In_1214);
nand U176 (N_176,In_889,In_770);
and U177 (N_177,In_47,In_377);
xor U178 (N_178,In_400,In_590);
nand U179 (N_179,In_602,In_98);
xor U180 (N_180,In_260,In_310);
nand U181 (N_181,In_1271,In_509);
nand U182 (N_182,In_891,In_1235);
xor U183 (N_183,In_911,In_531);
and U184 (N_184,In_434,In_225);
xnor U185 (N_185,In_1165,In_559);
nand U186 (N_186,In_767,In_892);
nor U187 (N_187,In_262,In_1222);
nand U188 (N_188,In_1458,In_1381);
nand U189 (N_189,In_539,In_913);
nand U190 (N_190,In_1078,In_1082);
nand U191 (N_191,In_848,In_890);
xor U192 (N_192,In_794,In_109);
xnor U193 (N_193,In_1278,In_1267);
or U194 (N_194,In_329,In_204);
xor U195 (N_195,In_1270,In_806);
nor U196 (N_196,In_963,In_1160);
xnor U197 (N_197,In_473,In_1086);
and U198 (N_198,In_747,In_549);
or U199 (N_199,In_1027,In_641);
or U200 (N_200,In_1215,In_705);
nand U201 (N_201,In_660,In_1140);
or U202 (N_202,In_985,In_146);
xnor U203 (N_203,In_175,In_137);
nor U204 (N_204,In_995,In_828);
nor U205 (N_205,In_681,In_284);
xnor U206 (N_206,In_1382,In_515);
xor U207 (N_207,In_1211,In_1137);
and U208 (N_208,In_279,In_442);
or U209 (N_209,In_223,In_272);
nand U210 (N_210,In_1269,In_1309);
nand U211 (N_211,In_551,In_572);
and U212 (N_212,In_254,In_650);
and U213 (N_213,In_1268,In_114);
nor U214 (N_214,In_1305,In_475);
and U215 (N_215,In_1116,In_908);
xor U216 (N_216,In_165,In_1257);
xor U217 (N_217,In_1076,In_875);
nand U218 (N_218,In_479,In_167);
or U219 (N_219,In_245,In_736);
nand U220 (N_220,In_1358,In_1356);
nand U221 (N_221,In_437,In_1144);
nand U222 (N_222,In_155,In_706);
nand U223 (N_223,In_1080,In_1181);
xor U224 (N_224,In_189,In_912);
nor U225 (N_225,In_1236,In_695);
xnor U226 (N_226,In_56,In_69);
xor U227 (N_227,In_694,In_1472);
and U228 (N_228,In_1162,In_265);
nand U229 (N_229,In_942,In_487);
nor U230 (N_230,In_1156,In_1192);
xor U231 (N_231,In_95,In_637);
and U232 (N_232,In_1200,In_692);
and U233 (N_233,In_1087,In_1028);
nor U234 (N_234,In_55,In_973);
or U235 (N_235,In_339,In_1024);
or U236 (N_236,In_1221,In_992);
and U237 (N_237,In_32,In_57);
and U238 (N_238,In_345,In_521);
nor U239 (N_239,In_573,In_599);
xnor U240 (N_240,In_317,In_938);
and U241 (N_241,In_64,In_1083);
xor U242 (N_242,In_998,In_990);
and U243 (N_243,In_930,In_606);
xor U244 (N_244,In_18,In_1126);
nand U245 (N_245,In_215,In_900);
nor U246 (N_246,In_1149,In_251);
nor U247 (N_247,In_790,In_679);
or U248 (N_248,In_1249,In_1120);
or U249 (N_249,In_1276,In_308);
or U250 (N_250,In_130,In_1281);
nor U251 (N_251,In_1239,In_578);
and U252 (N_252,In_1258,In_639);
and U253 (N_253,In_1019,In_1471);
nand U254 (N_254,In_1497,In_1141);
nor U255 (N_255,In_1224,In_61);
xnor U256 (N_256,In_1397,In_1491);
nor U257 (N_257,In_1015,In_1417);
xor U258 (N_258,In_1489,In_931);
xnor U259 (N_259,In_200,In_678);
and U260 (N_260,In_1444,In_546);
nor U261 (N_261,In_1157,In_801);
and U262 (N_262,In_823,In_787);
and U263 (N_263,In_750,In_154);
and U264 (N_264,In_965,In_644);
nand U265 (N_265,In_547,In_171);
nand U266 (N_266,In_1369,In_781);
or U267 (N_267,In_896,In_771);
nand U268 (N_268,In_186,In_854);
nor U269 (N_269,In_101,In_221);
nand U270 (N_270,In_74,In_376);
nand U271 (N_271,In_438,In_1445);
nor U272 (N_272,In_1404,In_334);
xnor U273 (N_273,In_76,In_757);
xor U274 (N_274,In_127,In_247);
and U275 (N_275,In_766,In_1260);
or U276 (N_276,In_1277,In_612);
nor U277 (N_277,In_667,In_1067);
or U278 (N_278,In_564,In_630);
nor U279 (N_279,In_465,In_275);
or U280 (N_280,In_1049,In_1022);
nor U281 (N_281,In_1041,In_594);
and U282 (N_282,In_1363,In_1133);
and U283 (N_283,In_197,In_1303);
and U284 (N_284,In_1161,In_1343);
xnor U285 (N_285,In_545,In_91);
nand U286 (N_286,In_212,In_319);
or U287 (N_287,In_1158,In_902);
xor U288 (N_288,In_555,In_323);
or U289 (N_289,In_105,In_89);
and U290 (N_290,In_1000,In_1429);
or U291 (N_291,In_1391,In_1307);
or U292 (N_292,In_226,In_1216);
and U293 (N_293,In_624,In_932);
or U294 (N_294,In_14,In_1390);
or U295 (N_295,In_655,In_21);
xor U296 (N_296,In_996,In_680);
or U297 (N_297,In_843,In_1432);
nor U298 (N_298,In_682,In_386);
nand U299 (N_299,In_582,In_580);
nor U300 (N_300,In_237,In_1231);
xnor U301 (N_301,In_63,In_360);
nor U302 (N_302,In_978,In_718);
xor U303 (N_303,In_286,In_1439);
nor U304 (N_304,In_609,In_1320);
nand U305 (N_305,In_525,In_759);
and U306 (N_306,In_1294,In_690);
xor U307 (N_307,In_1101,In_409);
xor U308 (N_308,In_534,In_474);
nor U309 (N_309,In_583,In_1493);
or U310 (N_310,In_1115,In_158);
xor U311 (N_311,In_1447,In_470);
nor U312 (N_312,In_234,In_1494);
or U313 (N_313,In_591,In_980);
and U314 (N_314,In_1124,In_951);
nand U315 (N_315,In_1322,In_166);
and U316 (N_316,In_35,In_491);
nor U317 (N_317,In_510,In_1104);
and U318 (N_318,In_1226,In_805);
nand U319 (N_319,In_94,In_659);
xnor U320 (N_320,In_252,In_1330);
nor U321 (N_321,In_1321,In_738);
or U322 (N_322,In_102,In_144);
nor U323 (N_323,In_748,In_792);
nor U324 (N_324,In_1191,In_1204);
nand U325 (N_325,In_406,In_1344);
nor U326 (N_326,In_1153,In_1201);
and U327 (N_327,In_987,In_1427);
nor U328 (N_328,In_688,In_1272);
xnor U329 (N_329,In_1014,In_554);
or U330 (N_330,In_132,In_1107);
or U331 (N_331,In_50,In_394);
xnor U332 (N_332,In_38,In_164);
and U333 (N_333,In_877,In_587);
xor U334 (N_334,In_852,In_8);
or U335 (N_335,In_1286,In_6);
xnor U336 (N_336,In_1383,In_396);
or U337 (N_337,In_1251,In_1207);
nor U338 (N_338,In_1408,In_840);
and U339 (N_339,In_768,In_263);
and U340 (N_340,In_832,In_145);
or U341 (N_341,In_575,In_780);
nor U342 (N_342,In_486,In_926);
nand U343 (N_343,In_530,In_846);
nor U344 (N_344,In_1057,In_236);
and U345 (N_345,In_1196,In_1380);
and U346 (N_346,In_1111,In_1114);
and U347 (N_347,In_1410,In_269);
xor U348 (N_348,In_1230,In_924);
nand U349 (N_349,In_1311,In_99);
xnor U350 (N_350,In_714,In_313);
nand U351 (N_351,In_632,In_498);
and U352 (N_352,In_907,In_244);
and U353 (N_353,In_1443,In_1442);
nand U354 (N_354,In_785,In_88);
and U355 (N_355,In_1486,In_1296);
xnor U356 (N_356,In_638,In_611);
nand U357 (N_357,In_119,In_218);
or U358 (N_358,In_544,In_652);
and U359 (N_359,In_903,In_803);
nand U360 (N_360,In_141,In_333);
xnor U361 (N_361,In_1291,In_446);
xor U362 (N_362,In_901,In_702);
nand U363 (N_363,In_328,In_1148);
or U364 (N_364,In_520,In_841);
nor U365 (N_365,In_1461,In_1421);
xnor U366 (N_366,In_147,In_42);
nor U367 (N_367,In_1169,In_928);
nor U368 (N_368,In_335,In_1166);
xnor U369 (N_369,In_152,In_86);
and U370 (N_370,In_1436,In_826);
nor U371 (N_371,In_960,In_277);
xor U372 (N_372,In_849,In_1333);
nor U373 (N_373,In_404,In_1037);
or U374 (N_374,In_1047,In_1422);
or U375 (N_375,In_149,In_962);
xnor U376 (N_376,In_1045,In_1056);
xor U377 (N_377,In_1102,In_503);
or U378 (N_378,In_468,In_373);
or U379 (N_379,In_494,In_922);
nor U380 (N_380,In_19,In_459);
and U381 (N_381,In_1127,In_70);
xor U382 (N_382,In_984,In_26);
or U383 (N_383,In_1285,In_1193);
nor U384 (N_384,In_1034,In_585);
and U385 (N_385,In_598,In_882);
xor U386 (N_386,In_123,In_981);
nor U387 (N_387,In_1350,In_676);
nor U388 (N_388,In_763,In_281);
or U389 (N_389,In_945,In_318);
xor U390 (N_390,In_886,In_274);
nand U391 (N_391,In_1490,In_1292);
xnor U392 (N_392,In_1463,In_108);
nor U393 (N_393,In_388,In_314);
or U394 (N_394,In_514,In_480);
nor U395 (N_395,In_366,In_700);
nor U396 (N_396,In_654,In_391);
xor U397 (N_397,In_278,In_1240);
and U398 (N_398,In_385,In_1361);
or U399 (N_399,In_1182,In_1299);
xnor U400 (N_400,In_1468,In_1453);
or U401 (N_401,In_290,In_919);
and U402 (N_402,In_813,In_1425);
nor U403 (N_403,In_916,In_699);
and U404 (N_404,In_1470,In_1008);
or U405 (N_405,In_1289,In_367);
nor U406 (N_406,In_1242,In_139);
and U407 (N_407,In_220,In_452);
and U408 (N_408,In_1347,In_174);
nand U409 (N_409,In_113,In_343);
nor U410 (N_410,In_614,In_1036);
and U411 (N_411,In_742,In_1368);
xnor U412 (N_412,In_809,In_222);
nand U413 (N_413,In_616,In_517);
or U414 (N_414,In_970,In_294);
or U415 (N_415,In_565,In_483);
nor U416 (N_416,In_1264,In_340);
nand U417 (N_417,In_605,In_825);
nor U418 (N_418,In_435,In_267);
or U419 (N_419,In_40,In_1);
or U420 (N_420,In_776,In_471);
nor U421 (N_421,In_542,In_190);
and U422 (N_422,In_34,In_967);
xnor U423 (N_423,In_188,In_1326);
nor U424 (N_424,In_791,In_1263);
or U425 (N_425,In_1184,In_711);
and U426 (N_426,In_372,In_561);
or U427 (N_427,In_986,In_325);
nand U428 (N_428,In_496,In_563);
xnor U429 (N_429,In_1248,In_620);
nand U430 (N_430,In_1081,In_389);
nand U431 (N_431,In_838,In_921);
xnor U432 (N_432,In_312,In_224);
xor U433 (N_433,In_1395,In_1043);
xnor U434 (N_434,In_131,In_1259);
and U435 (N_435,In_1180,In_774);
xnor U436 (N_436,In_927,In_431);
nand U437 (N_437,In_613,In_395);
nor U438 (N_438,In_454,In_1040);
or U439 (N_439,In_1012,In_1085);
nor U440 (N_440,In_814,In_800);
or U441 (N_441,In_799,In_276);
or U442 (N_442,In_1075,In_52);
nand U443 (N_443,In_601,In_784);
xnor U444 (N_444,In_666,In_610);
xor U445 (N_445,In_23,In_1317);
nor U446 (N_446,In_16,In_78);
nand U447 (N_447,In_1295,In_715);
or U448 (N_448,In_122,In_999);
nor U449 (N_449,In_125,In_899);
or U450 (N_450,In_934,In_208);
and U451 (N_451,In_227,In_248);
xnor U452 (N_452,In_291,In_460);
xor U453 (N_453,In_1252,In_789);
nor U454 (N_454,In_160,In_1331);
nand U455 (N_455,In_178,In_1440);
nand U456 (N_456,In_1290,In_1435);
and U457 (N_457,In_305,In_619);
nor U458 (N_458,In_421,In_569);
nor U459 (N_459,In_1462,In_10);
and U460 (N_460,In_725,In_810);
or U461 (N_461,In_1077,In_1070);
or U462 (N_462,In_444,In_497);
nor U463 (N_463,In_1123,In_753);
nand U464 (N_464,In_1044,In_734);
nand U465 (N_465,In_433,In_600);
nand U466 (N_466,In_249,In_216);
or U467 (N_467,In_1424,In_737);
or U468 (N_468,In_239,In_939);
nor U469 (N_469,In_1254,In_839);
nor U470 (N_470,In_1406,In_920);
and U471 (N_471,In_1253,In_929);
and U472 (N_472,In_2,In_1223);
and U473 (N_473,In_777,In_1446);
or U474 (N_474,In_242,In_1441);
xnor U475 (N_475,In_1274,In_358);
xor U476 (N_476,In_798,In_280);
xor U477 (N_477,In_1351,In_1469);
nor U478 (N_478,In_341,In_1234);
or U479 (N_479,In_300,In_507);
nand U480 (N_480,In_230,In_9);
or U481 (N_481,In_1129,In_744);
or U482 (N_482,In_818,In_1183);
xor U483 (N_483,In_1336,In_134);
nor U484 (N_484,In_1315,In_346);
nor U485 (N_485,In_150,In_501);
or U486 (N_486,In_1202,In_493);
or U487 (N_487,In_1007,In_1353);
xor U488 (N_488,In_721,In_1365);
or U489 (N_489,In_1346,In_1198);
and U490 (N_490,In_835,In_850);
xnor U491 (N_491,In_425,In_1366);
nor U492 (N_492,In_869,In_1301);
xnor U493 (N_493,In_448,In_1434);
or U494 (N_494,In_364,In_557);
nand U495 (N_495,In_157,In_1419);
and U496 (N_496,In_296,In_943);
or U497 (N_497,In_408,In_1373);
nand U498 (N_498,In_344,In_392);
nand U499 (N_499,In_1352,In_151);
and U500 (N_500,In_1225,In_570);
xor U501 (N_501,In_1061,In_722);
xnor U502 (N_502,In_782,In_634);
nor U503 (N_503,In_342,In_793);
and U504 (N_504,In_266,In_1454);
or U505 (N_505,In_622,In_536);
and U506 (N_506,In_1314,In_1220);
xor U507 (N_507,In_1066,In_1105);
or U508 (N_508,In_627,In_778);
or U509 (N_509,In_1186,In_1094);
and U510 (N_510,In_1228,In_860);
nand U511 (N_511,In_1244,In_629);
or U512 (N_512,In_878,In_658);
nand U513 (N_513,In_231,In_1378);
or U514 (N_514,In_321,In_1448);
nor U515 (N_515,In_370,In_795);
or U516 (N_516,In_90,In_1354);
xnor U517 (N_517,In_1485,In_1175);
nor U518 (N_518,In_898,In_847);
nor U519 (N_519,In_53,In_1467);
or U520 (N_520,In_548,In_79);
or U521 (N_521,In_804,In_1394);
or U522 (N_522,In_640,In_111);
xnor U523 (N_523,In_121,In_656);
nand U524 (N_524,In_968,In_307);
nand U525 (N_525,In_881,In_22);
nor U526 (N_526,In_1496,In_181);
nand U527 (N_527,In_665,In_508);
nand U528 (N_528,In_7,In_1054);
and U529 (N_529,In_326,In_96);
nor U530 (N_530,In_195,In_330);
xnor U531 (N_531,In_309,In_663);
or U532 (N_532,In_1409,In_1152);
or U533 (N_533,In_618,In_1385);
nand U534 (N_534,In_29,In_198);
nor U535 (N_535,In_623,In_1319);
and U536 (N_536,In_1155,In_1357);
or U537 (N_537,In_779,In_1178);
xor U538 (N_538,In_33,In_192);
or U539 (N_539,In_1498,In_161);
nor U540 (N_540,In_1218,In_879);
and U541 (N_541,In_1219,In_574);
xnor U542 (N_542,In_107,In_550);
or U543 (N_543,In_393,In_668);
or U544 (N_544,In_0,In_691);
nand U545 (N_545,In_1478,In_413);
nor U546 (N_546,In_380,In_885);
nand U547 (N_547,In_1420,In_1460);
or U548 (N_548,In_1068,In_977);
and U549 (N_549,In_1431,In_754);
and U550 (N_550,In_478,In_299);
or U551 (N_551,In_1195,In_75);
nor U552 (N_552,In_217,In_92);
and U553 (N_553,In_500,In_196);
or U554 (N_554,In_1456,In_1099);
nand U555 (N_555,In_1009,In_976);
nand U556 (N_556,In_1100,In_685);
nand U557 (N_557,In_816,In_1300);
nand U558 (N_558,In_100,In_1197);
and U559 (N_559,In_636,In_971);
or U560 (N_560,In_834,In_662);
nand U561 (N_561,In_541,In_1039);
or U562 (N_562,In_824,In_120);
and U563 (N_563,In_952,In_1136);
nand U564 (N_564,In_717,In_894);
xor U565 (N_565,In_472,In_1499);
and U566 (N_566,In_422,In_362);
xor U567 (N_567,In_664,In_905);
or U568 (N_568,In_463,In_719);
nor U569 (N_569,In_148,In_429);
nor U570 (N_570,In_235,In_571);
nand U571 (N_571,In_492,In_295);
nor U572 (N_572,In_796,In_1349);
or U573 (N_573,In_535,In_915);
and U574 (N_574,In_243,In_202);
or U575 (N_575,In_1376,In_379);
xor U576 (N_576,In_1227,In_1128);
xor U577 (N_577,In_1103,In_36);
or U578 (N_578,In_519,In_1145);
xor U579 (N_579,In_969,In_845);
nand U580 (N_580,In_73,In_424);
and U581 (N_581,In_283,In_85);
or U582 (N_582,In_1367,In_106);
xnor U583 (N_583,In_410,In_1032);
xor U584 (N_584,In_1030,In_1426);
nor U585 (N_585,In_815,In_822);
or U586 (N_586,In_499,In_1337);
xor U587 (N_587,In_772,In_851);
nand U588 (N_588,In_1131,In_1325);
or U589 (N_589,In_607,In_258);
xnor U590 (N_590,In_1438,In_1414);
xor U591 (N_591,In_1005,In_43);
nor U592 (N_592,In_635,In_704);
nand U593 (N_593,In_1059,In_588);
or U594 (N_594,In_1342,In_138);
or U595 (N_595,In_1065,In_762);
nand U596 (N_596,In_66,In_1119);
and U597 (N_597,In_68,In_353);
or U598 (N_598,In_989,In_1474);
xor U599 (N_599,In_947,In_1302);
or U600 (N_600,In_349,In_994);
or U601 (N_601,In_893,In_1001);
or U602 (N_602,In_193,In_529);
nor U603 (N_603,In_649,In_906);
or U604 (N_604,In_257,In_904);
nor U605 (N_605,In_775,In_831);
nand U606 (N_606,In_597,In_97);
xnor U607 (N_607,In_350,In_506);
and U608 (N_608,In_1098,In_1399);
xnor U609 (N_609,In_12,In_558);
xnor U610 (N_610,In_527,In_1031);
xnor U611 (N_611,In_369,In_39);
xnor U612 (N_612,In_673,In_712);
or U613 (N_613,In_866,In_1122);
or U614 (N_614,In_292,In_1255);
and U615 (N_615,In_402,In_271);
nand U616 (N_616,In_864,In_1312);
nor U617 (N_617,In_615,In_1232);
nor U618 (N_618,In_648,In_60);
nand U619 (N_619,In_1021,In_37);
or U620 (N_620,In_4,In_769);
and U621 (N_621,In_949,In_1492);
xnor U622 (N_622,In_661,In_959);
nor U623 (N_623,In_1370,In_1480);
nand U624 (N_624,In_1069,In_303);
nand U625 (N_625,In_1095,In_1372);
xor U626 (N_626,In_441,In_675);
nand U627 (N_627,In_210,In_348);
and U628 (N_628,In_693,In_1265);
and U629 (N_629,In_842,In_255);
nor U630 (N_630,In_1379,In_1110);
and U631 (N_631,In_232,In_954);
nor U632 (N_632,In_887,In_177);
nor U633 (N_633,In_643,In_1340);
or U634 (N_634,In_1273,In_817);
or U635 (N_635,In_1323,In_417);
and U636 (N_636,In_1203,In_713);
nor U637 (N_637,In_1430,In_1020);
or U638 (N_638,In_972,In_170);
nand U639 (N_639,In_347,In_464);
xnor U640 (N_640,In_1355,In_49);
or U641 (N_641,In_642,In_581);
and U642 (N_642,In_1171,In_398);
and U643 (N_643,In_1451,In_382);
or U644 (N_644,In_1213,In_213);
xor U645 (N_645,In_1038,In_1058);
nand U646 (N_646,In_1088,In_30);
nor U647 (N_647,In_982,In_1212);
nor U648 (N_648,In_352,In_1364);
xor U649 (N_649,In_374,In_1073);
nand U650 (N_650,In_439,In_1339);
nand U651 (N_651,In_1190,In_461);
and U652 (N_652,In_1437,In_1188);
nand U653 (N_653,In_933,In_941);
and U654 (N_654,In_489,In_1396);
and U655 (N_655,In_1466,In_495);
xor U656 (N_656,In_324,In_837);
and U657 (N_657,In_1483,In_833);
or U658 (N_658,In_1329,In_332);
xor U659 (N_659,In_729,In_883);
or U660 (N_660,In_423,In_48);
or U661 (N_661,In_1109,In_1013);
or U662 (N_662,In_1017,In_162);
and U663 (N_663,In_93,In_589);
nand U664 (N_664,In_631,In_45);
and U665 (N_665,In_405,In_709);
xor U666 (N_666,In_505,In_54);
and U667 (N_667,In_336,In_77);
or U668 (N_668,In_387,In_628);
xnor U669 (N_669,In_1318,In_455);
xor U670 (N_670,In_1064,In_761);
and U671 (N_671,In_504,In_595);
nor U672 (N_672,In_25,In_576);
xnor U673 (N_673,In_1205,In_403);
and U674 (N_674,In_868,In_1208);
and U675 (N_675,In_287,In_773);
xor U676 (N_676,In_1018,In_528);
and U677 (N_677,In_1341,In_1117);
and U678 (N_678,In_964,In_961);
nand U679 (N_679,In_397,In_940);
or U680 (N_680,In_1187,In_136);
and U681 (N_681,In_918,In_516);
xor U682 (N_682,In_268,In_966);
and U683 (N_683,In_1210,In_1328);
nor U684 (N_684,In_874,In_697);
nand U685 (N_685,In_1371,In_436);
or U686 (N_686,In_1338,In_84);
nand U687 (N_687,In_756,In_17);
xor U688 (N_688,In_997,In_1090);
and U689 (N_689,In_956,In_371);
or U690 (N_690,In_991,In_143);
and U691 (N_691,In_807,In_1481);
nor U692 (N_692,In_724,In_1006);
xor U693 (N_693,In_456,In_253);
nand U694 (N_694,In_1476,In_1062);
nand U695 (N_695,In_485,In_755);
and U696 (N_696,In_469,In_1023);
nand U697 (N_697,In_1293,In_645);
xor U698 (N_698,In_103,In_412);
xnor U699 (N_699,In_1151,In_696);
xor U700 (N_700,In_1288,In_1154);
nor U701 (N_701,In_1138,In_859);
nand U702 (N_702,In_746,In_256);
or U703 (N_703,In_1016,In_1243);
xor U704 (N_704,In_1482,In_1377);
or U705 (N_705,In_1072,In_1283);
and U706 (N_706,In_687,In_802);
and U707 (N_707,In_288,In_481);
and U708 (N_708,In_856,In_740);
or U709 (N_709,In_917,In_1298);
xor U710 (N_710,In_67,In_357);
and U711 (N_711,In_1011,In_579);
nor U712 (N_712,In_830,In_617);
nor U713 (N_713,In_540,In_626);
or U714 (N_714,In_1177,In_87);
nand U715 (N_715,In_338,In_289);
or U716 (N_716,In_1004,In_401);
and U717 (N_717,In_1360,In_829);
xnor U718 (N_718,In_1416,In_214);
xor U719 (N_719,In_876,In_760);
and U720 (N_720,In_1402,In_156);
nand U721 (N_721,In_1010,In_285);
xnor U722 (N_722,In_20,In_1042);
xor U723 (N_723,In_246,In_567);
nand U724 (N_724,In_701,In_1455);
or U725 (N_725,In_443,In_354);
xor U726 (N_726,In_80,In_1089);
xor U727 (N_727,In_430,In_672);
and U728 (N_728,In_556,In_5);
xnor U729 (N_729,In_909,In_1384);
or U730 (N_730,In_293,In_1327);
xnor U731 (N_731,In_176,In_211);
nor U732 (N_732,In_1475,In_880);
nand U733 (N_733,In_743,In_1233);
nand U734 (N_734,In_1245,In_1324);
and U735 (N_735,In_716,In_361);
and U736 (N_736,In_1035,In_1275);
and U737 (N_737,In_11,In_140);
nand U738 (N_738,In_458,In_173);
and U739 (N_739,In_1334,In_1097);
xnor U740 (N_740,In_751,In_383);
nand U741 (N_741,In_420,In_1279);
nor U742 (N_742,In_1025,In_1147);
nand U743 (N_743,In_72,In_1108);
xor U744 (N_744,In_82,In_844);
and U745 (N_745,In_153,In_1194);
xor U746 (N_746,In_1459,In_1121);
and U747 (N_747,In_647,In_31);
and U748 (N_748,In_651,In_871);
or U749 (N_749,In_233,In_1060);
or U750 (N_750,In_534,In_768);
and U751 (N_751,In_217,In_207);
nand U752 (N_752,In_1016,In_726);
xnor U753 (N_753,In_284,In_1436);
or U754 (N_754,In_457,In_701);
xnor U755 (N_755,In_657,In_22);
nand U756 (N_756,In_1047,In_639);
nand U757 (N_757,In_259,In_691);
nand U758 (N_758,In_1398,In_1006);
nand U759 (N_759,In_889,In_500);
xnor U760 (N_760,In_1117,In_729);
nor U761 (N_761,In_483,In_260);
and U762 (N_762,In_1371,In_1299);
and U763 (N_763,In_308,In_764);
xor U764 (N_764,In_669,In_1223);
and U765 (N_765,In_183,In_1044);
nand U766 (N_766,In_1230,In_757);
nor U767 (N_767,In_140,In_1349);
and U768 (N_768,In_419,In_631);
nor U769 (N_769,In_692,In_737);
xnor U770 (N_770,In_382,In_1164);
nor U771 (N_771,In_44,In_1165);
xor U772 (N_772,In_1404,In_267);
nor U773 (N_773,In_424,In_61);
xor U774 (N_774,In_162,In_67);
or U775 (N_775,In_958,In_473);
nand U776 (N_776,In_367,In_1377);
nand U777 (N_777,In_1185,In_53);
xor U778 (N_778,In_347,In_1060);
or U779 (N_779,In_68,In_1265);
or U780 (N_780,In_941,In_252);
xnor U781 (N_781,In_635,In_901);
nor U782 (N_782,In_348,In_1473);
or U783 (N_783,In_1342,In_634);
nand U784 (N_784,In_1192,In_1050);
xor U785 (N_785,In_1471,In_1058);
xor U786 (N_786,In_1224,In_1120);
nor U787 (N_787,In_477,In_238);
and U788 (N_788,In_459,In_843);
xnor U789 (N_789,In_414,In_1282);
nand U790 (N_790,In_1483,In_572);
and U791 (N_791,In_1450,In_1123);
nand U792 (N_792,In_456,In_208);
xor U793 (N_793,In_509,In_1436);
nor U794 (N_794,In_1240,In_174);
nand U795 (N_795,In_99,In_324);
and U796 (N_796,In_608,In_1219);
xor U797 (N_797,In_1135,In_818);
and U798 (N_798,In_623,In_721);
nor U799 (N_799,In_523,In_1229);
and U800 (N_800,In_613,In_1238);
and U801 (N_801,In_1088,In_911);
xor U802 (N_802,In_850,In_36);
nor U803 (N_803,In_1065,In_692);
nand U804 (N_804,In_145,In_829);
nor U805 (N_805,In_1020,In_566);
or U806 (N_806,In_1262,In_356);
nand U807 (N_807,In_1226,In_862);
nor U808 (N_808,In_575,In_1422);
and U809 (N_809,In_582,In_1097);
or U810 (N_810,In_327,In_421);
nor U811 (N_811,In_487,In_1027);
xor U812 (N_812,In_519,In_312);
xnor U813 (N_813,In_924,In_229);
or U814 (N_814,In_66,In_1083);
or U815 (N_815,In_1168,In_966);
nor U816 (N_816,In_987,In_1220);
xnor U817 (N_817,In_1322,In_715);
and U818 (N_818,In_979,In_487);
xnor U819 (N_819,In_307,In_1268);
nor U820 (N_820,In_1425,In_1298);
nand U821 (N_821,In_1297,In_687);
and U822 (N_822,In_901,In_794);
nor U823 (N_823,In_1226,In_134);
or U824 (N_824,In_1160,In_243);
and U825 (N_825,In_731,In_734);
nor U826 (N_826,In_573,In_769);
nand U827 (N_827,In_456,In_597);
and U828 (N_828,In_1410,In_385);
or U829 (N_829,In_225,In_861);
xor U830 (N_830,In_795,In_1297);
and U831 (N_831,In_1315,In_262);
or U832 (N_832,In_690,In_442);
or U833 (N_833,In_489,In_383);
xnor U834 (N_834,In_1170,In_1004);
or U835 (N_835,In_1121,In_953);
and U836 (N_836,In_1486,In_656);
nand U837 (N_837,In_275,In_208);
nand U838 (N_838,In_818,In_1420);
xor U839 (N_839,In_1439,In_1227);
xor U840 (N_840,In_380,In_482);
nand U841 (N_841,In_1316,In_490);
or U842 (N_842,In_1356,In_264);
and U843 (N_843,In_42,In_1448);
and U844 (N_844,In_285,In_748);
nor U845 (N_845,In_836,In_563);
and U846 (N_846,In_1056,In_865);
and U847 (N_847,In_1499,In_407);
and U848 (N_848,In_1443,In_405);
and U849 (N_849,In_1027,In_1330);
or U850 (N_850,In_1363,In_415);
nand U851 (N_851,In_432,In_762);
xor U852 (N_852,In_374,In_118);
nand U853 (N_853,In_924,In_390);
nor U854 (N_854,In_965,In_800);
and U855 (N_855,In_127,In_1025);
xnor U856 (N_856,In_826,In_895);
xnor U857 (N_857,In_190,In_1472);
and U858 (N_858,In_15,In_1095);
xnor U859 (N_859,In_347,In_68);
or U860 (N_860,In_722,In_665);
nor U861 (N_861,In_179,In_606);
nand U862 (N_862,In_1411,In_748);
or U863 (N_863,In_199,In_1441);
and U864 (N_864,In_344,In_1387);
and U865 (N_865,In_1116,In_682);
or U866 (N_866,In_452,In_1044);
or U867 (N_867,In_1423,In_1360);
and U868 (N_868,In_120,In_333);
nand U869 (N_869,In_964,In_471);
xor U870 (N_870,In_184,In_231);
nand U871 (N_871,In_322,In_349);
nor U872 (N_872,In_1442,In_1088);
and U873 (N_873,In_847,In_1097);
or U874 (N_874,In_21,In_179);
nand U875 (N_875,In_1348,In_766);
xor U876 (N_876,In_1123,In_1020);
xor U877 (N_877,In_400,In_1396);
and U878 (N_878,In_802,In_1467);
xor U879 (N_879,In_620,In_1200);
nor U880 (N_880,In_103,In_74);
nand U881 (N_881,In_1221,In_755);
nand U882 (N_882,In_829,In_711);
nor U883 (N_883,In_457,In_1097);
nor U884 (N_884,In_1107,In_1205);
nor U885 (N_885,In_670,In_957);
xnor U886 (N_886,In_630,In_1089);
nor U887 (N_887,In_1136,In_90);
xor U888 (N_888,In_16,In_595);
xnor U889 (N_889,In_112,In_873);
or U890 (N_890,In_322,In_59);
nor U891 (N_891,In_392,In_1106);
and U892 (N_892,In_1445,In_1289);
xnor U893 (N_893,In_679,In_549);
nand U894 (N_894,In_982,In_803);
xnor U895 (N_895,In_752,In_1214);
xor U896 (N_896,In_1102,In_1007);
nand U897 (N_897,In_1340,In_1395);
or U898 (N_898,In_534,In_1154);
nor U899 (N_899,In_1305,In_320);
or U900 (N_900,In_9,In_915);
nand U901 (N_901,In_472,In_908);
or U902 (N_902,In_989,In_746);
nor U903 (N_903,In_447,In_1119);
xor U904 (N_904,In_335,In_282);
nand U905 (N_905,In_820,In_701);
nor U906 (N_906,In_732,In_606);
nand U907 (N_907,In_746,In_247);
and U908 (N_908,In_322,In_371);
and U909 (N_909,In_231,In_1122);
xor U910 (N_910,In_705,In_19);
nand U911 (N_911,In_1492,In_94);
nor U912 (N_912,In_491,In_1201);
xnor U913 (N_913,In_1384,In_89);
or U914 (N_914,In_166,In_1243);
xnor U915 (N_915,In_183,In_721);
nor U916 (N_916,In_1019,In_1010);
or U917 (N_917,In_363,In_23);
or U918 (N_918,In_1410,In_654);
nor U919 (N_919,In_400,In_82);
or U920 (N_920,In_190,In_1128);
and U921 (N_921,In_17,In_1470);
and U922 (N_922,In_284,In_999);
or U923 (N_923,In_521,In_951);
or U924 (N_924,In_1231,In_716);
nand U925 (N_925,In_1426,In_826);
nor U926 (N_926,In_439,In_287);
and U927 (N_927,In_674,In_1045);
xnor U928 (N_928,In_1415,In_1082);
xnor U929 (N_929,In_547,In_1011);
and U930 (N_930,In_25,In_865);
nand U931 (N_931,In_1331,In_803);
nor U932 (N_932,In_886,In_875);
xnor U933 (N_933,In_646,In_525);
nor U934 (N_934,In_766,In_735);
nand U935 (N_935,In_1402,In_867);
nand U936 (N_936,In_526,In_1287);
or U937 (N_937,In_1080,In_405);
and U938 (N_938,In_1181,In_313);
or U939 (N_939,In_325,In_667);
or U940 (N_940,In_216,In_1297);
or U941 (N_941,In_536,In_1390);
nand U942 (N_942,In_1041,In_35);
nand U943 (N_943,In_578,In_355);
nand U944 (N_944,In_1355,In_867);
nand U945 (N_945,In_324,In_587);
and U946 (N_946,In_222,In_1086);
nand U947 (N_947,In_191,In_563);
xor U948 (N_948,In_823,In_1418);
nor U949 (N_949,In_489,In_268);
or U950 (N_950,In_606,In_1475);
nor U951 (N_951,In_1369,In_1148);
nor U952 (N_952,In_1332,In_806);
and U953 (N_953,In_57,In_633);
and U954 (N_954,In_255,In_814);
or U955 (N_955,In_1319,In_148);
nor U956 (N_956,In_908,In_392);
and U957 (N_957,In_1342,In_767);
nand U958 (N_958,In_948,In_812);
or U959 (N_959,In_121,In_695);
xor U960 (N_960,In_797,In_116);
nand U961 (N_961,In_490,In_752);
and U962 (N_962,In_755,In_1355);
nand U963 (N_963,In_1057,In_622);
or U964 (N_964,In_263,In_464);
nor U965 (N_965,In_776,In_655);
nor U966 (N_966,In_1272,In_27);
and U967 (N_967,In_267,In_521);
xnor U968 (N_968,In_150,In_802);
nor U969 (N_969,In_987,In_1399);
nor U970 (N_970,In_420,In_1262);
and U971 (N_971,In_135,In_1423);
xnor U972 (N_972,In_60,In_233);
nor U973 (N_973,In_1388,In_659);
nor U974 (N_974,In_135,In_711);
nor U975 (N_975,In_1148,In_293);
nand U976 (N_976,In_756,In_43);
nand U977 (N_977,In_187,In_782);
and U978 (N_978,In_772,In_1452);
nor U979 (N_979,In_278,In_37);
nor U980 (N_980,In_367,In_918);
xnor U981 (N_981,In_1150,In_537);
and U982 (N_982,In_1303,In_1408);
nor U983 (N_983,In_136,In_767);
xnor U984 (N_984,In_1373,In_1137);
or U985 (N_985,In_1495,In_1302);
or U986 (N_986,In_87,In_31);
nor U987 (N_987,In_656,In_1134);
or U988 (N_988,In_303,In_452);
and U989 (N_989,In_820,In_1245);
or U990 (N_990,In_1346,In_67);
xor U991 (N_991,In_711,In_288);
or U992 (N_992,In_548,In_610);
nor U993 (N_993,In_1131,In_1455);
nor U994 (N_994,In_263,In_782);
and U995 (N_995,In_286,In_1245);
and U996 (N_996,In_660,In_865);
and U997 (N_997,In_994,In_55);
nor U998 (N_998,In_1050,In_1344);
nor U999 (N_999,In_935,In_143);
nor U1000 (N_1000,N_0,N_465);
xor U1001 (N_1001,N_779,N_770);
and U1002 (N_1002,N_81,N_556);
xnor U1003 (N_1003,N_606,N_402);
and U1004 (N_1004,N_226,N_953);
xor U1005 (N_1005,N_169,N_150);
xnor U1006 (N_1006,N_989,N_324);
nor U1007 (N_1007,N_537,N_462);
nand U1008 (N_1008,N_723,N_731);
xnor U1009 (N_1009,N_333,N_706);
nand U1010 (N_1010,N_860,N_526);
or U1011 (N_1011,N_107,N_819);
or U1012 (N_1012,N_557,N_390);
or U1013 (N_1013,N_604,N_51);
nand U1014 (N_1014,N_547,N_159);
nand U1015 (N_1015,N_354,N_973);
or U1016 (N_1016,N_182,N_196);
or U1017 (N_1017,N_11,N_659);
and U1018 (N_1018,N_689,N_845);
nor U1019 (N_1019,N_21,N_934);
nor U1020 (N_1020,N_135,N_483);
nor U1021 (N_1021,N_175,N_612);
nand U1022 (N_1022,N_65,N_717);
or U1023 (N_1023,N_886,N_593);
nand U1024 (N_1024,N_589,N_710);
xor U1025 (N_1025,N_112,N_539);
nor U1026 (N_1026,N_430,N_345);
nor U1027 (N_1027,N_592,N_910);
or U1028 (N_1028,N_514,N_444);
xor U1029 (N_1029,N_8,N_963);
nor U1030 (N_1030,N_85,N_814);
and U1031 (N_1031,N_715,N_296);
nand U1032 (N_1032,N_249,N_875);
nand U1033 (N_1033,N_15,N_550);
xnor U1034 (N_1034,N_272,N_419);
nand U1035 (N_1035,N_87,N_732);
nand U1036 (N_1036,N_984,N_184);
xnor U1037 (N_1037,N_221,N_40);
nor U1038 (N_1038,N_287,N_610);
nand U1039 (N_1039,N_136,N_358);
and U1040 (N_1040,N_303,N_62);
nor U1041 (N_1041,N_145,N_628);
or U1042 (N_1042,N_362,N_290);
nand U1043 (N_1043,N_903,N_785);
nor U1044 (N_1044,N_985,N_520);
xnor U1045 (N_1045,N_231,N_747);
nor U1046 (N_1046,N_868,N_377);
nand U1047 (N_1047,N_677,N_666);
or U1048 (N_1048,N_437,N_30);
nor U1049 (N_1049,N_309,N_359);
or U1050 (N_1050,N_906,N_554);
nor U1051 (N_1051,N_113,N_896);
xnor U1052 (N_1052,N_394,N_262);
nor U1053 (N_1053,N_928,N_339);
and U1054 (N_1054,N_157,N_801);
xor U1055 (N_1055,N_937,N_316);
xnor U1056 (N_1056,N_281,N_944);
or U1057 (N_1057,N_237,N_713);
or U1058 (N_1058,N_890,N_803);
or U1059 (N_1059,N_168,N_684);
and U1060 (N_1060,N_172,N_337);
xor U1061 (N_1061,N_841,N_477);
nand U1062 (N_1062,N_340,N_240);
nand U1063 (N_1063,N_523,N_307);
and U1064 (N_1064,N_207,N_880);
or U1065 (N_1065,N_117,N_189);
nor U1066 (N_1066,N_314,N_425);
or U1067 (N_1067,N_297,N_108);
xor U1068 (N_1068,N_332,N_180);
nor U1069 (N_1069,N_773,N_688);
xor U1070 (N_1070,N_536,N_218);
nor U1071 (N_1071,N_486,N_644);
xor U1072 (N_1072,N_469,N_538);
and U1073 (N_1073,N_326,N_63);
nand U1074 (N_1074,N_84,N_697);
nand U1075 (N_1075,N_828,N_772);
or U1076 (N_1076,N_96,N_929);
xor U1077 (N_1077,N_698,N_99);
xor U1078 (N_1078,N_975,N_413);
and U1079 (N_1079,N_844,N_19);
and U1080 (N_1080,N_621,N_204);
xor U1081 (N_1081,N_369,N_368);
xor U1082 (N_1082,N_443,N_267);
or U1083 (N_1083,N_692,N_161);
or U1084 (N_1084,N_453,N_230);
xor U1085 (N_1085,N_969,N_508);
xor U1086 (N_1086,N_306,N_948);
nand U1087 (N_1087,N_435,N_280);
nand U1088 (N_1088,N_106,N_711);
and U1089 (N_1089,N_133,N_351);
nand U1090 (N_1090,N_728,N_178);
and U1091 (N_1091,N_160,N_44);
or U1092 (N_1092,N_986,N_146);
nand U1093 (N_1093,N_118,N_490);
or U1094 (N_1094,N_742,N_568);
xnor U1095 (N_1095,N_774,N_859);
and U1096 (N_1096,N_170,N_909);
nand U1097 (N_1097,N_387,N_856);
nor U1098 (N_1098,N_195,N_813);
and U1099 (N_1099,N_636,N_75);
and U1100 (N_1100,N_642,N_385);
or U1101 (N_1101,N_573,N_510);
xor U1102 (N_1102,N_766,N_38);
and U1103 (N_1103,N_433,N_327);
and U1104 (N_1104,N_877,N_727);
xnor U1105 (N_1105,N_116,N_565);
and U1106 (N_1106,N_755,N_43);
nor U1107 (N_1107,N_751,N_241);
nand U1108 (N_1108,N_648,N_591);
nor U1109 (N_1109,N_485,N_939);
and U1110 (N_1110,N_846,N_501);
xnor U1111 (N_1111,N_61,N_791);
nand U1112 (N_1112,N_609,N_972);
nand U1113 (N_1113,N_153,N_676);
xor U1114 (N_1114,N_276,N_349);
nor U1115 (N_1115,N_566,N_397);
nand U1116 (N_1116,N_217,N_293);
and U1117 (N_1117,N_505,N_981);
and U1118 (N_1118,N_509,N_3);
nor U1119 (N_1119,N_367,N_709);
xor U1120 (N_1120,N_29,N_432);
xor U1121 (N_1121,N_4,N_600);
and U1122 (N_1122,N_524,N_251);
nor U1123 (N_1123,N_696,N_53);
nand U1124 (N_1124,N_561,N_708);
nor U1125 (N_1125,N_79,N_750);
xor U1126 (N_1126,N_257,N_882);
or U1127 (N_1127,N_28,N_899);
xnor U1128 (N_1128,N_285,N_756);
and U1129 (N_1129,N_827,N_990);
xnor U1130 (N_1130,N_121,N_590);
nor U1131 (N_1131,N_849,N_424);
xor U1132 (N_1132,N_542,N_391);
nand U1133 (N_1133,N_822,N_323);
nand U1134 (N_1134,N_586,N_529);
or U1135 (N_1135,N_236,N_457);
nand U1136 (N_1136,N_900,N_474);
and U1137 (N_1137,N_414,N_716);
or U1138 (N_1138,N_487,N_873);
nor U1139 (N_1139,N_993,N_553);
xnor U1140 (N_1140,N_871,N_320);
or U1141 (N_1141,N_734,N_122);
or U1142 (N_1142,N_464,N_611);
xnor U1143 (N_1143,N_795,N_833);
xor U1144 (N_1144,N_872,N_321);
nand U1145 (N_1145,N_735,N_86);
and U1146 (N_1146,N_914,N_898);
or U1147 (N_1147,N_942,N_567);
or U1148 (N_1148,N_999,N_506);
nand U1149 (N_1149,N_638,N_317);
or U1150 (N_1150,N_620,N_461);
and U1151 (N_1151,N_344,N_162);
or U1152 (N_1152,N_407,N_881);
xnor U1153 (N_1153,N_515,N_821);
and U1154 (N_1154,N_216,N_493);
or U1155 (N_1155,N_870,N_534);
nand U1156 (N_1156,N_489,N_174);
nor U1157 (N_1157,N_258,N_330);
or U1158 (N_1158,N_192,N_16);
nand U1159 (N_1159,N_607,N_533);
or U1160 (N_1160,N_410,N_625);
or U1161 (N_1161,N_458,N_250);
and U1162 (N_1162,N_507,N_420);
nor U1163 (N_1163,N_163,N_370);
nor U1164 (N_1164,N_102,N_256);
and U1165 (N_1165,N_137,N_201);
or U1166 (N_1166,N_799,N_793);
xor U1167 (N_1167,N_862,N_98);
or U1168 (N_1168,N_90,N_156);
nor U1169 (N_1169,N_718,N_234);
and U1170 (N_1170,N_315,N_748);
nand U1171 (N_1171,N_94,N_781);
nand U1172 (N_1172,N_674,N_603);
nor U1173 (N_1173,N_253,N_70);
nand U1174 (N_1174,N_954,N_782);
or U1175 (N_1175,N_416,N_152);
xor U1176 (N_1176,N_434,N_919);
nor U1177 (N_1177,N_48,N_543);
nand U1178 (N_1178,N_657,N_439);
nor U1179 (N_1179,N_661,N_970);
or U1180 (N_1180,N_587,N_426);
or U1181 (N_1181,N_513,N_166);
xor U1182 (N_1182,N_701,N_863);
nand U1183 (N_1183,N_925,N_843);
nand U1184 (N_1184,N_699,N_380);
or U1185 (N_1185,N_105,N_491);
nor U1186 (N_1186,N_824,N_431);
nand U1187 (N_1187,N_737,N_951);
xor U1188 (N_1188,N_436,N_730);
nand U1189 (N_1189,N_915,N_746);
and U1190 (N_1190,N_632,N_202);
or U1191 (N_1191,N_421,N_653);
or U1192 (N_1192,N_974,N_911);
nand U1193 (N_1193,N_476,N_259);
xnor U1194 (N_1194,N_649,N_960);
nor U1195 (N_1195,N_356,N_670);
nand U1196 (N_1196,N_268,N_572);
xnor U1197 (N_1197,N_254,N_222);
xnor U1198 (N_1198,N_357,N_947);
or U1199 (N_1199,N_197,N_233);
or U1200 (N_1200,N_138,N_940);
nand U1201 (N_1201,N_167,N_245);
nand U1202 (N_1202,N_384,N_941);
xor U1203 (N_1203,N_705,N_594);
xor U1204 (N_1204,N_576,N_68);
nand U1205 (N_1205,N_473,N_831);
or U1206 (N_1206,N_114,N_78);
xor U1207 (N_1207,N_27,N_151);
nand U1208 (N_1208,N_905,N_685);
nor U1209 (N_1209,N_325,N_838);
nand U1210 (N_1210,N_129,N_294);
and U1211 (N_1211,N_408,N_996);
xnor U1212 (N_1212,N_82,N_726);
or U1213 (N_1213,N_190,N_348);
nand U1214 (N_1214,N_298,N_69);
nor U1215 (N_1215,N_322,N_968);
xnor U1216 (N_1216,N_95,N_994);
nand U1217 (N_1217,N_398,N_191);
nor U1218 (N_1218,N_777,N_312);
or U1219 (N_1219,N_456,N_784);
xor U1220 (N_1220,N_88,N_978);
and U1221 (N_1221,N_57,N_527);
or U1222 (N_1222,N_578,N_757);
or U1223 (N_1223,N_37,N_946);
xor U1224 (N_1224,N_155,N_127);
xor U1225 (N_1225,N_866,N_375);
nand U1226 (N_1226,N_209,N_480);
or U1227 (N_1227,N_459,N_46);
nor U1228 (N_1228,N_269,N_2);
and U1229 (N_1229,N_998,N_422);
or U1230 (N_1230,N_14,N_580);
xnor U1231 (N_1231,N_598,N_411);
or U1232 (N_1232,N_763,N_379);
nand U1233 (N_1233,N_551,N_512);
xor U1234 (N_1234,N_311,N_336);
nand U1235 (N_1235,N_468,N_641);
xnor U1236 (N_1236,N_749,N_647);
and U1237 (N_1237,N_992,N_679);
nor U1238 (N_1238,N_805,N_829);
xor U1239 (N_1239,N_203,N_289);
nand U1240 (N_1240,N_401,N_186);
nand U1241 (N_1241,N_400,N_71);
nand U1242 (N_1242,N_36,N_364);
nand U1243 (N_1243,N_719,N_549);
nand U1244 (N_1244,N_879,N_24);
xnor U1245 (N_1245,N_405,N_404);
nand U1246 (N_1246,N_132,N_235);
and U1247 (N_1247,N_694,N_555);
xor U1248 (N_1248,N_788,N_54);
or U1249 (N_1249,N_669,N_807);
or U1250 (N_1250,N_148,N_342);
or U1251 (N_1251,N_373,N_310);
nor U1252 (N_1252,N_761,N_173);
and U1253 (N_1253,N_664,N_855);
or U1254 (N_1254,N_738,N_759);
and U1255 (N_1255,N_584,N_809);
xnor U1256 (N_1256,N_406,N_745);
xnor U1257 (N_1257,N_183,N_577);
xnor U1258 (N_1258,N_273,N_199);
xnor U1259 (N_1259,N_193,N_574);
nand U1260 (N_1260,N_760,N_229);
nor U1261 (N_1261,N_502,N_252);
and U1262 (N_1262,N_255,N_977);
xor U1263 (N_1263,N_517,N_511);
and U1264 (N_1264,N_945,N_979);
nand U1265 (N_1265,N_32,N_17);
or U1266 (N_1266,N_25,N_680);
or U1267 (N_1267,N_56,N_912);
nand U1268 (N_1268,N_101,N_720);
xnor U1269 (N_1269,N_579,N_907);
nor U1270 (N_1270,N_823,N_125);
and U1271 (N_1271,N_494,N_995);
nor U1272 (N_1272,N_18,N_399);
and U1273 (N_1273,N_758,N_614);
nor U1274 (N_1274,N_637,N_961);
and U1275 (N_1275,N_712,N_208);
nor U1276 (N_1276,N_35,N_23);
nor U1277 (N_1277,N_707,N_198);
and U1278 (N_1278,N_671,N_286);
nor U1279 (N_1279,N_335,N_67);
nand U1280 (N_1280,N_215,N_662);
nor U1281 (N_1281,N_930,N_9);
nand U1282 (N_1282,N_278,N_288);
or U1283 (N_1283,N_149,N_481);
or U1284 (N_1284,N_851,N_583);
nor U1285 (N_1285,N_392,N_683);
xnor U1286 (N_1286,N_595,N_22);
nand U1287 (N_1287,N_918,N_936);
nand U1288 (N_1288,N_20,N_672);
xor U1289 (N_1289,N_522,N_894);
or U1290 (N_1290,N_423,N_5);
nand U1291 (N_1291,N_334,N_91);
nand U1292 (N_1292,N_164,N_834);
nand U1293 (N_1293,N_59,N_639);
and U1294 (N_1294,N_646,N_244);
xnor U1295 (N_1295,N_381,N_284);
xor U1296 (N_1296,N_858,N_219);
xor U1297 (N_1297,N_313,N_353);
xor U1298 (N_1298,N_427,N_546);
nand U1299 (N_1299,N_608,N_451);
xnor U1300 (N_1300,N_765,N_588);
and U1301 (N_1301,N_605,N_49);
or U1302 (N_1302,N_528,N_495);
nand U1303 (N_1303,N_270,N_531);
and U1304 (N_1304,N_545,N_214);
or U1305 (N_1305,N_722,N_847);
and U1306 (N_1306,N_319,N_109);
or U1307 (N_1307,N_452,N_675);
nor U1308 (N_1308,N_615,N_33);
nand U1309 (N_1309,N_365,N_123);
or U1310 (N_1310,N_623,N_503);
and U1311 (N_1311,N_652,N_617);
nand U1312 (N_1312,N_352,N_239);
or U1313 (N_1313,N_581,N_966);
xnor U1314 (N_1314,N_787,N_12);
nand U1315 (N_1315,N_158,N_943);
and U1316 (N_1316,N_518,N_300);
nand U1317 (N_1317,N_988,N_724);
xor U1318 (N_1318,N_55,N_857);
nand U1319 (N_1319,N_139,N_864);
or U1320 (N_1320,N_837,N_475);
nand U1321 (N_1321,N_144,N_991);
or U1322 (N_1322,N_635,N_802);
nor U1323 (N_1323,N_962,N_569);
nor U1324 (N_1324,N_171,N_769);
or U1325 (N_1325,N_570,N_34);
and U1326 (N_1326,N_897,N_181);
and U1327 (N_1327,N_564,N_100);
xor U1328 (N_1328,N_955,N_825);
or U1329 (N_1329,N_26,N_640);
xor U1330 (N_1330,N_386,N_304);
xor U1331 (N_1331,N_396,N_403);
and U1332 (N_1332,N_525,N_927);
or U1333 (N_1333,N_764,N_128);
nand U1334 (N_1334,N_200,N_89);
xnor U1335 (N_1335,N_130,N_931);
nor U1336 (N_1336,N_187,N_922);
nand U1337 (N_1337,N_448,N_134);
and U1338 (N_1338,N_780,N_210);
xnor U1339 (N_1339,N_277,N_225);
and U1340 (N_1340,N_840,N_768);
nor U1341 (N_1341,N_976,N_559);
nor U1342 (N_1342,N_908,N_839);
and U1343 (N_1343,N_308,N_884);
or U1344 (N_1344,N_361,N_874);
or U1345 (N_1345,N_582,N_741);
or U1346 (N_1346,N_811,N_622);
nor U1347 (N_1347,N_42,N_889);
nand U1348 (N_1348,N_775,N_869);
nand U1349 (N_1349,N_74,N_496);
nand U1350 (N_1350,N_454,N_935);
nand U1351 (N_1351,N_967,N_497);
or U1352 (N_1352,N_832,N_393);
nand U1353 (N_1353,N_540,N_224);
and U1354 (N_1354,N_261,N_602);
and U1355 (N_1355,N_58,N_887);
nand U1356 (N_1356,N_767,N_783);
or U1357 (N_1357,N_363,N_654);
nor U1358 (N_1358,N_301,N_740);
xor U1359 (N_1359,N_228,N_441);
nand U1360 (N_1360,N_933,N_563);
nor U1361 (N_1361,N_613,N_265);
nand U1362 (N_1362,N_283,N_678);
nor U1363 (N_1363,N_264,N_376);
xor U1364 (N_1364,N_959,N_77);
xnor U1365 (N_1365,N_206,N_143);
nor U1366 (N_1366,N_630,N_292);
xor U1367 (N_1367,N_558,N_532);
nor U1368 (N_1368,N_904,N_227);
nor U1369 (N_1369,N_552,N_371);
nor U1370 (N_1370,N_338,N_263);
nand U1371 (N_1371,N_725,N_836);
nor U1372 (N_1372,N_7,N_388);
and U1373 (N_1373,N_971,N_762);
or U1374 (N_1374,N_665,N_800);
and U1375 (N_1375,N_119,N_687);
nor U1376 (N_1376,N_848,N_893);
xnor U1377 (N_1377,N_140,N_651);
or U1378 (N_1378,N_798,N_956);
and U1379 (N_1379,N_482,N_374);
and U1380 (N_1380,N_560,N_110);
xor U1381 (N_1381,N_445,N_861);
nor U1382 (N_1382,N_796,N_47);
nand U1383 (N_1383,N_350,N_341);
or U1384 (N_1384,N_484,N_519);
nor U1385 (N_1385,N_6,N_13);
and U1386 (N_1386,N_498,N_412);
and U1387 (N_1387,N_471,N_76);
xor U1388 (N_1388,N_39,N_949);
nor U1389 (N_1389,N_810,N_778);
and U1390 (N_1390,N_378,N_729);
xnor U1391 (N_1391,N_347,N_530);
and U1392 (N_1392,N_901,N_704);
or U1393 (N_1393,N_274,N_176);
and U1394 (N_1394,N_295,N_575);
xor U1395 (N_1395,N_460,N_142);
nor U1396 (N_1396,N_417,N_693);
nor U1397 (N_1397,N_562,N_690);
nor U1398 (N_1398,N_804,N_987);
nand U1399 (N_1399,N_700,N_429);
and U1400 (N_1400,N_104,N_479);
or U1401 (N_1401,N_842,N_571);
xnor U1402 (N_1402,N_852,N_818);
nand U1403 (N_1403,N_242,N_521);
xor U1404 (N_1404,N_667,N_921);
nor U1405 (N_1405,N_428,N_926);
or U1406 (N_1406,N_599,N_466);
or U1407 (N_1407,N_329,N_544);
xor U1408 (N_1408,N_126,N_878);
or U1409 (N_1409,N_41,N_205);
or U1410 (N_1410,N_790,N_141);
nor U1411 (N_1411,N_629,N_31);
nand U1412 (N_1412,N_656,N_744);
and U1413 (N_1413,N_721,N_902);
nor U1414 (N_1414,N_753,N_681);
xor U1415 (N_1415,N_920,N_663);
or U1416 (N_1416,N_913,N_279);
nor U1417 (N_1417,N_739,N_409);
nor U1418 (N_1418,N_876,N_695);
and U1419 (N_1419,N_808,N_247);
xnor U1420 (N_1420,N_463,N_771);
nor U1421 (N_1421,N_179,N_535);
or U1422 (N_1422,N_624,N_645);
or U1423 (N_1423,N_888,N_660);
nand U1424 (N_1424,N_786,N_923);
or U1425 (N_1425,N_343,N_754);
nand U1426 (N_1426,N_982,N_147);
xnor U1427 (N_1427,N_854,N_291);
or U1428 (N_1428,N_455,N_643);
nor U1429 (N_1429,N_447,N_305);
and U1430 (N_1430,N_916,N_792);
nor U1431 (N_1431,N_658,N_103);
xnor U1432 (N_1432,N_938,N_446);
and U1433 (N_1433,N_585,N_633);
nand U1434 (N_1434,N_789,N_52);
nand U1435 (N_1435,N_248,N_188);
nand U1436 (N_1436,N_246,N_92);
nor U1437 (N_1437,N_932,N_470);
xor U1438 (N_1438,N_165,N_131);
nor U1439 (N_1439,N_812,N_631);
xor U1440 (N_1440,N_980,N_243);
xor U1441 (N_1441,N_797,N_440);
nor U1442 (N_1442,N_299,N_60);
nor U1443 (N_1443,N_355,N_826);
or U1444 (N_1444,N_650,N_736);
xor U1445 (N_1445,N_302,N_111);
or U1446 (N_1446,N_597,N_395);
and U1447 (N_1447,N_865,N_917);
nand U1448 (N_1448,N_924,N_442);
or U1449 (N_1449,N_504,N_634);
and U1450 (N_1450,N_714,N_817);
nor U1451 (N_1451,N_957,N_952);
and U1452 (N_1452,N_958,N_835);
and U1453 (N_1453,N_212,N_627);
nor U1454 (N_1454,N_282,N_691);
and U1455 (N_1455,N_619,N_418);
nand U1456 (N_1456,N_883,N_478);
or U1457 (N_1457,N_271,N_266);
or U1458 (N_1458,N_72,N_93);
nor U1459 (N_1459,N_382,N_820);
or U1460 (N_1460,N_806,N_815);
nor U1461 (N_1461,N_548,N_346);
xnor U1462 (N_1462,N_83,N_275);
nor U1463 (N_1463,N_850,N_776);
or U1464 (N_1464,N_499,N_673);
xor U1465 (N_1465,N_867,N_500);
nor U1466 (N_1466,N_885,N_64);
nand U1467 (N_1467,N_964,N_626);
nor U1468 (N_1468,N_73,N_115);
and U1469 (N_1469,N_655,N_541);
xnor U1470 (N_1470,N_686,N_360);
nor U1471 (N_1471,N_220,N_472);
nand U1472 (N_1472,N_45,N_50);
nand U1473 (N_1473,N_194,N_668);
xnor U1474 (N_1474,N_816,N_366);
and U1475 (N_1475,N_415,N_983);
nand U1476 (N_1476,N_702,N_703);
xnor U1477 (N_1477,N_80,N_211);
nor U1478 (N_1478,N_177,N_830);
nor U1479 (N_1479,N_10,N_743);
or U1480 (N_1480,N_97,N_492);
and U1481 (N_1481,N_601,N_450);
xnor U1482 (N_1482,N_223,N_213);
nand U1483 (N_1483,N_618,N_185);
nand U1484 (N_1484,N_596,N_232);
xnor U1485 (N_1485,N_154,N_752);
nand U1486 (N_1486,N_449,N_120);
or U1487 (N_1487,N_895,N_260);
nand U1488 (N_1488,N_891,N_853);
or U1489 (N_1489,N_372,N_331);
xor U1490 (N_1490,N_328,N_682);
nor U1491 (N_1491,N_383,N_318);
or U1492 (N_1492,N_892,N_124);
and U1493 (N_1493,N_950,N_616);
xnor U1494 (N_1494,N_997,N_733);
and U1495 (N_1495,N_467,N_66);
and U1496 (N_1496,N_516,N_238);
nand U1497 (N_1497,N_794,N_488);
and U1498 (N_1498,N_438,N_1);
nand U1499 (N_1499,N_965,N_389);
and U1500 (N_1500,N_88,N_760);
nor U1501 (N_1501,N_634,N_651);
or U1502 (N_1502,N_229,N_938);
and U1503 (N_1503,N_42,N_630);
nor U1504 (N_1504,N_284,N_961);
and U1505 (N_1505,N_232,N_28);
and U1506 (N_1506,N_194,N_927);
or U1507 (N_1507,N_501,N_70);
and U1508 (N_1508,N_674,N_396);
and U1509 (N_1509,N_377,N_833);
and U1510 (N_1510,N_629,N_538);
nor U1511 (N_1511,N_66,N_723);
or U1512 (N_1512,N_111,N_26);
nand U1513 (N_1513,N_587,N_2);
xnor U1514 (N_1514,N_944,N_902);
nor U1515 (N_1515,N_866,N_966);
xor U1516 (N_1516,N_833,N_686);
nor U1517 (N_1517,N_372,N_336);
nor U1518 (N_1518,N_893,N_42);
nand U1519 (N_1519,N_287,N_422);
nor U1520 (N_1520,N_258,N_891);
or U1521 (N_1521,N_108,N_271);
xnor U1522 (N_1522,N_745,N_147);
or U1523 (N_1523,N_772,N_983);
nand U1524 (N_1524,N_417,N_646);
xnor U1525 (N_1525,N_221,N_462);
xor U1526 (N_1526,N_546,N_279);
nand U1527 (N_1527,N_306,N_302);
nand U1528 (N_1528,N_998,N_993);
xor U1529 (N_1529,N_386,N_249);
nand U1530 (N_1530,N_787,N_367);
xnor U1531 (N_1531,N_213,N_585);
and U1532 (N_1532,N_832,N_591);
xor U1533 (N_1533,N_326,N_665);
and U1534 (N_1534,N_169,N_696);
or U1535 (N_1535,N_446,N_380);
nor U1536 (N_1536,N_441,N_804);
or U1537 (N_1537,N_338,N_127);
nor U1538 (N_1538,N_585,N_795);
nand U1539 (N_1539,N_34,N_64);
or U1540 (N_1540,N_761,N_499);
or U1541 (N_1541,N_503,N_774);
or U1542 (N_1542,N_301,N_801);
nor U1543 (N_1543,N_554,N_447);
nand U1544 (N_1544,N_647,N_386);
or U1545 (N_1545,N_552,N_416);
nor U1546 (N_1546,N_639,N_272);
or U1547 (N_1547,N_310,N_893);
nand U1548 (N_1548,N_259,N_568);
and U1549 (N_1549,N_700,N_407);
xor U1550 (N_1550,N_248,N_342);
nor U1551 (N_1551,N_563,N_976);
nor U1552 (N_1552,N_648,N_734);
xor U1553 (N_1553,N_880,N_759);
and U1554 (N_1554,N_556,N_338);
or U1555 (N_1555,N_272,N_301);
xor U1556 (N_1556,N_40,N_478);
xor U1557 (N_1557,N_783,N_797);
nor U1558 (N_1558,N_851,N_242);
nand U1559 (N_1559,N_208,N_890);
and U1560 (N_1560,N_348,N_273);
xnor U1561 (N_1561,N_639,N_868);
nor U1562 (N_1562,N_165,N_862);
nand U1563 (N_1563,N_19,N_346);
nand U1564 (N_1564,N_169,N_351);
and U1565 (N_1565,N_816,N_352);
xnor U1566 (N_1566,N_198,N_324);
or U1567 (N_1567,N_776,N_446);
nand U1568 (N_1568,N_456,N_995);
and U1569 (N_1569,N_413,N_763);
and U1570 (N_1570,N_641,N_227);
and U1571 (N_1571,N_717,N_765);
or U1572 (N_1572,N_495,N_12);
nor U1573 (N_1573,N_249,N_677);
nor U1574 (N_1574,N_261,N_498);
or U1575 (N_1575,N_889,N_822);
xor U1576 (N_1576,N_317,N_726);
nor U1577 (N_1577,N_295,N_587);
nor U1578 (N_1578,N_235,N_724);
or U1579 (N_1579,N_368,N_888);
or U1580 (N_1580,N_780,N_109);
nor U1581 (N_1581,N_854,N_522);
xnor U1582 (N_1582,N_610,N_204);
and U1583 (N_1583,N_514,N_687);
nand U1584 (N_1584,N_530,N_519);
or U1585 (N_1585,N_824,N_24);
or U1586 (N_1586,N_868,N_736);
nand U1587 (N_1587,N_912,N_753);
nor U1588 (N_1588,N_941,N_306);
nand U1589 (N_1589,N_79,N_641);
and U1590 (N_1590,N_866,N_42);
and U1591 (N_1591,N_38,N_674);
nor U1592 (N_1592,N_967,N_172);
nor U1593 (N_1593,N_876,N_608);
and U1594 (N_1594,N_337,N_578);
or U1595 (N_1595,N_717,N_760);
or U1596 (N_1596,N_410,N_676);
and U1597 (N_1597,N_997,N_812);
and U1598 (N_1598,N_950,N_22);
nor U1599 (N_1599,N_597,N_38);
nand U1600 (N_1600,N_548,N_79);
xor U1601 (N_1601,N_669,N_657);
or U1602 (N_1602,N_253,N_173);
xnor U1603 (N_1603,N_10,N_835);
nand U1604 (N_1604,N_509,N_418);
nand U1605 (N_1605,N_263,N_953);
nor U1606 (N_1606,N_51,N_610);
nand U1607 (N_1607,N_178,N_55);
nand U1608 (N_1608,N_627,N_205);
xnor U1609 (N_1609,N_795,N_356);
and U1610 (N_1610,N_891,N_63);
or U1611 (N_1611,N_602,N_931);
and U1612 (N_1612,N_357,N_278);
or U1613 (N_1613,N_79,N_918);
and U1614 (N_1614,N_329,N_459);
nor U1615 (N_1615,N_719,N_302);
nor U1616 (N_1616,N_679,N_22);
xnor U1617 (N_1617,N_657,N_307);
xor U1618 (N_1618,N_497,N_712);
xor U1619 (N_1619,N_659,N_749);
xnor U1620 (N_1620,N_834,N_546);
or U1621 (N_1621,N_769,N_369);
nor U1622 (N_1622,N_444,N_858);
nand U1623 (N_1623,N_637,N_948);
nor U1624 (N_1624,N_39,N_794);
nor U1625 (N_1625,N_900,N_545);
nand U1626 (N_1626,N_462,N_821);
nand U1627 (N_1627,N_965,N_370);
nand U1628 (N_1628,N_292,N_150);
nand U1629 (N_1629,N_219,N_780);
nand U1630 (N_1630,N_49,N_827);
and U1631 (N_1631,N_665,N_747);
nand U1632 (N_1632,N_390,N_823);
or U1633 (N_1633,N_872,N_225);
and U1634 (N_1634,N_777,N_732);
xnor U1635 (N_1635,N_241,N_268);
and U1636 (N_1636,N_868,N_902);
nand U1637 (N_1637,N_288,N_426);
and U1638 (N_1638,N_279,N_2);
xor U1639 (N_1639,N_529,N_504);
nor U1640 (N_1640,N_793,N_57);
nor U1641 (N_1641,N_758,N_468);
nor U1642 (N_1642,N_1,N_768);
xnor U1643 (N_1643,N_635,N_141);
and U1644 (N_1644,N_952,N_147);
and U1645 (N_1645,N_639,N_128);
nand U1646 (N_1646,N_878,N_596);
or U1647 (N_1647,N_16,N_230);
or U1648 (N_1648,N_976,N_712);
or U1649 (N_1649,N_64,N_803);
nor U1650 (N_1650,N_961,N_371);
or U1651 (N_1651,N_91,N_890);
xor U1652 (N_1652,N_183,N_223);
nor U1653 (N_1653,N_197,N_928);
or U1654 (N_1654,N_371,N_656);
nor U1655 (N_1655,N_898,N_11);
xor U1656 (N_1656,N_533,N_460);
xnor U1657 (N_1657,N_488,N_197);
and U1658 (N_1658,N_404,N_139);
or U1659 (N_1659,N_988,N_868);
nor U1660 (N_1660,N_773,N_735);
xor U1661 (N_1661,N_269,N_808);
xor U1662 (N_1662,N_178,N_771);
or U1663 (N_1663,N_574,N_175);
xor U1664 (N_1664,N_946,N_72);
nand U1665 (N_1665,N_555,N_786);
and U1666 (N_1666,N_71,N_527);
nand U1667 (N_1667,N_469,N_588);
nand U1668 (N_1668,N_725,N_951);
nand U1669 (N_1669,N_32,N_943);
xnor U1670 (N_1670,N_834,N_55);
and U1671 (N_1671,N_173,N_371);
nand U1672 (N_1672,N_783,N_460);
nor U1673 (N_1673,N_156,N_628);
xor U1674 (N_1674,N_586,N_636);
or U1675 (N_1675,N_256,N_802);
nand U1676 (N_1676,N_12,N_241);
xnor U1677 (N_1677,N_361,N_644);
or U1678 (N_1678,N_682,N_290);
xor U1679 (N_1679,N_171,N_286);
and U1680 (N_1680,N_592,N_216);
nor U1681 (N_1681,N_815,N_60);
or U1682 (N_1682,N_171,N_147);
nand U1683 (N_1683,N_425,N_544);
nor U1684 (N_1684,N_88,N_821);
nor U1685 (N_1685,N_102,N_782);
nor U1686 (N_1686,N_800,N_533);
or U1687 (N_1687,N_123,N_754);
xnor U1688 (N_1688,N_698,N_359);
xor U1689 (N_1689,N_890,N_316);
nor U1690 (N_1690,N_665,N_94);
xnor U1691 (N_1691,N_579,N_165);
nand U1692 (N_1692,N_956,N_860);
nand U1693 (N_1693,N_739,N_736);
and U1694 (N_1694,N_143,N_495);
or U1695 (N_1695,N_900,N_251);
nand U1696 (N_1696,N_258,N_778);
nor U1697 (N_1697,N_84,N_367);
and U1698 (N_1698,N_111,N_764);
and U1699 (N_1699,N_221,N_303);
and U1700 (N_1700,N_102,N_387);
nand U1701 (N_1701,N_810,N_180);
nand U1702 (N_1702,N_244,N_723);
xnor U1703 (N_1703,N_926,N_724);
and U1704 (N_1704,N_44,N_827);
and U1705 (N_1705,N_562,N_649);
or U1706 (N_1706,N_151,N_210);
nand U1707 (N_1707,N_835,N_440);
nor U1708 (N_1708,N_664,N_386);
nor U1709 (N_1709,N_308,N_514);
nor U1710 (N_1710,N_725,N_524);
and U1711 (N_1711,N_481,N_320);
and U1712 (N_1712,N_799,N_730);
xnor U1713 (N_1713,N_609,N_200);
and U1714 (N_1714,N_482,N_666);
nor U1715 (N_1715,N_479,N_868);
nor U1716 (N_1716,N_676,N_201);
nor U1717 (N_1717,N_592,N_768);
nor U1718 (N_1718,N_770,N_202);
nand U1719 (N_1719,N_350,N_177);
nor U1720 (N_1720,N_429,N_312);
or U1721 (N_1721,N_690,N_852);
and U1722 (N_1722,N_521,N_746);
nor U1723 (N_1723,N_52,N_883);
and U1724 (N_1724,N_571,N_653);
xnor U1725 (N_1725,N_783,N_356);
xor U1726 (N_1726,N_823,N_39);
and U1727 (N_1727,N_662,N_992);
or U1728 (N_1728,N_656,N_618);
and U1729 (N_1729,N_281,N_557);
and U1730 (N_1730,N_46,N_60);
xnor U1731 (N_1731,N_431,N_976);
nand U1732 (N_1732,N_510,N_67);
or U1733 (N_1733,N_24,N_204);
nand U1734 (N_1734,N_775,N_80);
or U1735 (N_1735,N_801,N_6);
xor U1736 (N_1736,N_870,N_871);
nor U1737 (N_1737,N_759,N_754);
nand U1738 (N_1738,N_128,N_236);
or U1739 (N_1739,N_481,N_666);
nor U1740 (N_1740,N_511,N_866);
nand U1741 (N_1741,N_225,N_530);
nor U1742 (N_1742,N_769,N_763);
nor U1743 (N_1743,N_722,N_220);
or U1744 (N_1744,N_560,N_420);
and U1745 (N_1745,N_846,N_812);
nand U1746 (N_1746,N_732,N_674);
and U1747 (N_1747,N_431,N_490);
or U1748 (N_1748,N_455,N_759);
or U1749 (N_1749,N_586,N_469);
nor U1750 (N_1750,N_636,N_949);
or U1751 (N_1751,N_341,N_166);
or U1752 (N_1752,N_966,N_266);
and U1753 (N_1753,N_217,N_510);
xor U1754 (N_1754,N_469,N_450);
and U1755 (N_1755,N_391,N_333);
xnor U1756 (N_1756,N_987,N_500);
nor U1757 (N_1757,N_630,N_467);
or U1758 (N_1758,N_558,N_528);
nor U1759 (N_1759,N_79,N_855);
or U1760 (N_1760,N_333,N_544);
xnor U1761 (N_1761,N_146,N_220);
and U1762 (N_1762,N_854,N_312);
nand U1763 (N_1763,N_493,N_618);
or U1764 (N_1764,N_496,N_800);
xor U1765 (N_1765,N_271,N_755);
and U1766 (N_1766,N_715,N_49);
nor U1767 (N_1767,N_184,N_222);
or U1768 (N_1768,N_634,N_80);
nor U1769 (N_1769,N_453,N_266);
or U1770 (N_1770,N_925,N_613);
and U1771 (N_1771,N_356,N_322);
xor U1772 (N_1772,N_514,N_674);
nor U1773 (N_1773,N_160,N_682);
nand U1774 (N_1774,N_287,N_676);
nor U1775 (N_1775,N_575,N_19);
and U1776 (N_1776,N_24,N_997);
and U1777 (N_1777,N_279,N_849);
nor U1778 (N_1778,N_625,N_479);
nand U1779 (N_1779,N_651,N_150);
nor U1780 (N_1780,N_563,N_127);
or U1781 (N_1781,N_224,N_732);
or U1782 (N_1782,N_628,N_399);
xor U1783 (N_1783,N_84,N_712);
xnor U1784 (N_1784,N_774,N_41);
nor U1785 (N_1785,N_234,N_959);
and U1786 (N_1786,N_399,N_591);
nand U1787 (N_1787,N_198,N_171);
and U1788 (N_1788,N_620,N_914);
and U1789 (N_1789,N_160,N_409);
and U1790 (N_1790,N_494,N_23);
xor U1791 (N_1791,N_913,N_222);
xor U1792 (N_1792,N_641,N_823);
or U1793 (N_1793,N_312,N_72);
nand U1794 (N_1794,N_652,N_198);
xor U1795 (N_1795,N_520,N_750);
nand U1796 (N_1796,N_142,N_214);
or U1797 (N_1797,N_373,N_376);
or U1798 (N_1798,N_956,N_179);
nand U1799 (N_1799,N_902,N_934);
or U1800 (N_1800,N_211,N_362);
nand U1801 (N_1801,N_375,N_745);
nand U1802 (N_1802,N_971,N_448);
and U1803 (N_1803,N_506,N_379);
or U1804 (N_1804,N_213,N_35);
nand U1805 (N_1805,N_783,N_69);
and U1806 (N_1806,N_833,N_898);
and U1807 (N_1807,N_422,N_816);
nand U1808 (N_1808,N_206,N_640);
nor U1809 (N_1809,N_473,N_463);
or U1810 (N_1810,N_508,N_609);
nor U1811 (N_1811,N_885,N_200);
nor U1812 (N_1812,N_125,N_935);
nor U1813 (N_1813,N_628,N_415);
or U1814 (N_1814,N_194,N_940);
nor U1815 (N_1815,N_72,N_962);
nand U1816 (N_1816,N_389,N_99);
nand U1817 (N_1817,N_729,N_481);
xnor U1818 (N_1818,N_634,N_303);
nand U1819 (N_1819,N_902,N_706);
and U1820 (N_1820,N_293,N_890);
xor U1821 (N_1821,N_461,N_513);
nor U1822 (N_1822,N_869,N_654);
or U1823 (N_1823,N_748,N_588);
xor U1824 (N_1824,N_773,N_473);
or U1825 (N_1825,N_746,N_273);
and U1826 (N_1826,N_744,N_267);
nand U1827 (N_1827,N_368,N_0);
or U1828 (N_1828,N_59,N_673);
or U1829 (N_1829,N_32,N_796);
nand U1830 (N_1830,N_658,N_557);
nor U1831 (N_1831,N_962,N_825);
or U1832 (N_1832,N_379,N_857);
nand U1833 (N_1833,N_301,N_252);
xor U1834 (N_1834,N_820,N_425);
or U1835 (N_1835,N_553,N_346);
xor U1836 (N_1836,N_792,N_321);
nand U1837 (N_1837,N_710,N_868);
and U1838 (N_1838,N_842,N_497);
nor U1839 (N_1839,N_654,N_355);
nor U1840 (N_1840,N_762,N_849);
nand U1841 (N_1841,N_335,N_905);
nor U1842 (N_1842,N_709,N_251);
nand U1843 (N_1843,N_117,N_528);
nor U1844 (N_1844,N_98,N_93);
or U1845 (N_1845,N_611,N_399);
nor U1846 (N_1846,N_228,N_435);
or U1847 (N_1847,N_111,N_314);
and U1848 (N_1848,N_408,N_872);
or U1849 (N_1849,N_703,N_740);
nor U1850 (N_1850,N_329,N_211);
xor U1851 (N_1851,N_599,N_365);
xnor U1852 (N_1852,N_993,N_577);
xor U1853 (N_1853,N_70,N_278);
and U1854 (N_1854,N_964,N_288);
xor U1855 (N_1855,N_748,N_576);
nor U1856 (N_1856,N_329,N_399);
xnor U1857 (N_1857,N_155,N_380);
or U1858 (N_1858,N_556,N_478);
or U1859 (N_1859,N_539,N_706);
or U1860 (N_1860,N_699,N_611);
or U1861 (N_1861,N_358,N_15);
nand U1862 (N_1862,N_121,N_766);
nand U1863 (N_1863,N_152,N_673);
nor U1864 (N_1864,N_968,N_65);
or U1865 (N_1865,N_994,N_911);
nor U1866 (N_1866,N_378,N_758);
nand U1867 (N_1867,N_776,N_655);
nand U1868 (N_1868,N_90,N_686);
and U1869 (N_1869,N_224,N_390);
xor U1870 (N_1870,N_404,N_266);
or U1871 (N_1871,N_926,N_933);
nand U1872 (N_1872,N_850,N_999);
nor U1873 (N_1873,N_25,N_85);
or U1874 (N_1874,N_133,N_761);
or U1875 (N_1875,N_73,N_468);
or U1876 (N_1876,N_31,N_528);
or U1877 (N_1877,N_524,N_641);
xor U1878 (N_1878,N_761,N_572);
and U1879 (N_1879,N_968,N_451);
nand U1880 (N_1880,N_231,N_47);
nor U1881 (N_1881,N_839,N_268);
nor U1882 (N_1882,N_715,N_225);
or U1883 (N_1883,N_847,N_607);
xor U1884 (N_1884,N_398,N_530);
nand U1885 (N_1885,N_314,N_171);
and U1886 (N_1886,N_262,N_997);
and U1887 (N_1887,N_904,N_887);
nor U1888 (N_1888,N_227,N_482);
nor U1889 (N_1889,N_300,N_647);
and U1890 (N_1890,N_257,N_371);
and U1891 (N_1891,N_420,N_812);
or U1892 (N_1892,N_708,N_266);
and U1893 (N_1893,N_949,N_986);
nor U1894 (N_1894,N_720,N_957);
and U1895 (N_1895,N_147,N_293);
and U1896 (N_1896,N_760,N_749);
or U1897 (N_1897,N_182,N_708);
xor U1898 (N_1898,N_685,N_147);
nand U1899 (N_1899,N_218,N_0);
xor U1900 (N_1900,N_263,N_109);
and U1901 (N_1901,N_844,N_410);
and U1902 (N_1902,N_432,N_190);
nor U1903 (N_1903,N_790,N_800);
nor U1904 (N_1904,N_506,N_562);
nor U1905 (N_1905,N_980,N_207);
xor U1906 (N_1906,N_59,N_590);
nor U1907 (N_1907,N_869,N_915);
xor U1908 (N_1908,N_466,N_278);
nor U1909 (N_1909,N_991,N_228);
nand U1910 (N_1910,N_137,N_62);
xnor U1911 (N_1911,N_899,N_890);
nor U1912 (N_1912,N_170,N_821);
nand U1913 (N_1913,N_422,N_304);
xor U1914 (N_1914,N_731,N_803);
nor U1915 (N_1915,N_442,N_219);
nor U1916 (N_1916,N_99,N_929);
or U1917 (N_1917,N_18,N_175);
nand U1918 (N_1918,N_64,N_486);
or U1919 (N_1919,N_559,N_269);
nor U1920 (N_1920,N_314,N_50);
xnor U1921 (N_1921,N_118,N_248);
nor U1922 (N_1922,N_283,N_938);
and U1923 (N_1923,N_112,N_230);
nand U1924 (N_1924,N_478,N_891);
xnor U1925 (N_1925,N_41,N_381);
or U1926 (N_1926,N_107,N_632);
or U1927 (N_1927,N_876,N_892);
xor U1928 (N_1928,N_742,N_658);
nand U1929 (N_1929,N_618,N_502);
and U1930 (N_1930,N_241,N_773);
or U1931 (N_1931,N_40,N_719);
nand U1932 (N_1932,N_973,N_202);
or U1933 (N_1933,N_896,N_415);
nor U1934 (N_1934,N_196,N_165);
and U1935 (N_1935,N_307,N_212);
nor U1936 (N_1936,N_667,N_147);
nand U1937 (N_1937,N_833,N_26);
and U1938 (N_1938,N_855,N_694);
nand U1939 (N_1939,N_120,N_702);
and U1940 (N_1940,N_717,N_91);
and U1941 (N_1941,N_94,N_986);
and U1942 (N_1942,N_988,N_158);
and U1943 (N_1943,N_63,N_488);
xnor U1944 (N_1944,N_448,N_302);
and U1945 (N_1945,N_320,N_780);
nor U1946 (N_1946,N_367,N_267);
xnor U1947 (N_1947,N_686,N_958);
xnor U1948 (N_1948,N_162,N_950);
nor U1949 (N_1949,N_79,N_578);
nor U1950 (N_1950,N_580,N_475);
xor U1951 (N_1951,N_118,N_398);
nor U1952 (N_1952,N_50,N_0);
and U1953 (N_1953,N_265,N_852);
xor U1954 (N_1954,N_743,N_691);
xnor U1955 (N_1955,N_236,N_899);
and U1956 (N_1956,N_792,N_582);
or U1957 (N_1957,N_689,N_314);
xnor U1958 (N_1958,N_748,N_330);
or U1959 (N_1959,N_18,N_744);
or U1960 (N_1960,N_226,N_419);
or U1961 (N_1961,N_834,N_352);
nand U1962 (N_1962,N_968,N_669);
and U1963 (N_1963,N_650,N_144);
xor U1964 (N_1964,N_654,N_83);
nor U1965 (N_1965,N_87,N_785);
nor U1966 (N_1966,N_584,N_622);
xor U1967 (N_1967,N_804,N_75);
or U1968 (N_1968,N_533,N_212);
and U1969 (N_1969,N_491,N_378);
nor U1970 (N_1970,N_154,N_175);
and U1971 (N_1971,N_852,N_723);
and U1972 (N_1972,N_401,N_226);
nor U1973 (N_1973,N_881,N_375);
xor U1974 (N_1974,N_405,N_285);
or U1975 (N_1975,N_453,N_51);
xnor U1976 (N_1976,N_59,N_346);
nor U1977 (N_1977,N_484,N_97);
nand U1978 (N_1978,N_47,N_966);
xor U1979 (N_1979,N_664,N_357);
xor U1980 (N_1980,N_31,N_536);
xnor U1981 (N_1981,N_158,N_188);
nand U1982 (N_1982,N_10,N_301);
or U1983 (N_1983,N_298,N_144);
and U1984 (N_1984,N_456,N_312);
nand U1985 (N_1985,N_537,N_729);
xnor U1986 (N_1986,N_774,N_769);
xor U1987 (N_1987,N_554,N_43);
nor U1988 (N_1988,N_91,N_828);
or U1989 (N_1989,N_235,N_608);
or U1990 (N_1990,N_598,N_797);
xnor U1991 (N_1991,N_190,N_71);
nand U1992 (N_1992,N_186,N_179);
or U1993 (N_1993,N_175,N_27);
xnor U1994 (N_1994,N_678,N_934);
nor U1995 (N_1995,N_304,N_938);
or U1996 (N_1996,N_462,N_119);
xor U1997 (N_1997,N_476,N_501);
nand U1998 (N_1998,N_791,N_614);
nor U1999 (N_1999,N_455,N_183);
nor U2000 (N_2000,N_1893,N_1325);
xnor U2001 (N_2001,N_1224,N_1473);
nor U2002 (N_2002,N_1243,N_1166);
and U2003 (N_2003,N_1687,N_1212);
nand U2004 (N_2004,N_1927,N_1593);
nor U2005 (N_2005,N_1969,N_1784);
and U2006 (N_2006,N_1836,N_1288);
and U2007 (N_2007,N_1978,N_1804);
and U2008 (N_2008,N_1630,N_1680);
nand U2009 (N_2009,N_1960,N_1356);
nor U2010 (N_2010,N_1386,N_1782);
nand U2011 (N_2011,N_1946,N_1152);
and U2012 (N_2012,N_1575,N_1823);
and U2013 (N_2013,N_1449,N_1013);
nand U2014 (N_2014,N_1874,N_1176);
nor U2015 (N_2015,N_1493,N_1292);
nor U2016 (N_2016,N_1928,N_1581);
nor U2017 (N_2017,N_1659,N_1898);
or U2018 (N_2018,N_1372,N_1636);
nor U2019 (N_2019,N_1350,N_1240);
nor U2020 (N_2020,N_1500,N_1147);
xnor U2021 (N_2021,N_1663,N_1448);
nand U2022 (N_2022,N_1868,N_1091);
nor U2023 (N_2023,N_1711,N_1870);
nor U2024 (N_2024,N_1661,N_1279);
xor U2025 (N_2025,N_1549,N_1304);
or U2026 (N_2026,N_1786,N_1562);
or U2027 (N_2027,N_1457,N_1080);
xnor U2028 (N_2028,N_1787,N_1516);
and U2029 (N_2029,N_1227,N_1496);
xor U2030 (N_2030,N_1184,N_1252);
xor U2031 (N_2031,N_1320,N_1451);
nand U2032 (N_2032,N_1805,N_1869);
nand U2033 (N_2033,N_1750,N_1125);
nor U2034 (N_2034,N_1880,N_1168);
and U2035 (N_2035,N_1317,N_1192);
or U2036 (N_2036,N_1172,N_1190);
or U2037 (N_2037,N_1682,N_1937);
nand U2038 (N_2038,N_1363,N_1040);
and U2039 (N_2039,N_1533,N_1383);
or U2040 (N_2040,N_1268,N_1608);
or U2041 (N_2041,N_1828,N_1128);
nand U2042 (N_2042,N_1289,N_1485);
xnor U2043 (N_2043,N_1681,N_1117);
and U2044 (N_2044,N_1370,N_1482);
nor U2045 (N_2045,N_1997,N_1111);
nand U2046 (N_2046,N_1980,N_1855);
nand U2047 (N_2047,N_1234,N_1050);
nand U2048 (N_2048,N_1708,N_1217);
nor U2049 (N_2049,N_1440,N_1196);
or U2050 (N_2050,N_1657,N_1803);
nand U2051 (N_2051,N_1223,N_1506);
and U2052 (N_2052,N_1300,N_1436);
nand U2053 (N_2053,N_1334,N_1016);
nor U2054 (N_2054,N_1902,N_1469);
or U2055 (N_2055,N_1367,N_1497);
nand U2056 (N_2056,N_1915,N_1468);
nor U2057 (N_2057,N_1036,N_1311);
xor U2058 (N_2058,N_1344,N_1783);
xnor U2059 (N_2059,N_1038,N_1671);
and U2060 (N_2060,N_1364,N_1421);
nor U2061 (N_2061,N_1834,N_1156);
or U2062 (N_2062,N_1812,N_1404);
xor U2063 (N_2063,N_1753,N_1976);
or U2064 (N_2064,N_1751,N_1800);
or U2065 (N_2065,N_1603,N_1480);
nor U2066 (N_2066,N_1492,N_1498);
or U2067 (N_2067,N_1861,N_1071);
xor U2068 (N_2068,N_1972,N_1063);
and U2069 (N_2069,N_1616,N_1802);
or U2070 (N_2070,N_1160,N_1570);
or U2071 (N_2071,N_1715,N_1664);
nand U2072 (N_2072,N_1433,N_1548);
nor U2073 (N_2073,N_1914,N_1863);
and U2074 (N_2074,N_1258,N_1723);
nor U2075 (N_2075,N_1662,N_1261);
nor U2076 (N_2076,N_1707,N_1423);
or U2077 (N_2077,N_1745,N_1435);
or U2078 (N_2078,N_1286,N_1652);
xor U2079 (N_2079,N_1820,N_1860);
nor U2080 (N_2080,N_1271,N_1226);
nor U2081 (N_2081,N_1700,N_1264);
xnor U2082 (N_2082,N_1489,N_1420);
nand U2083 (N_2083,N_1012,N_1845);
nand U2084 (N_2084,N_1442,N_1116);
or U2085 (N_2085,N_1503,N_1504);
and U2086 (N_2086,N_1337,N_1591);
nor U2087 (N_2087,N_1683,N_1043);
xor U2088 (N_2088,N_1505,N_1371);
nand U2089 (N_2089,N_1244,N_1000);
nand U2090 (N_2090,N_1971,N_1573);
nor U2091 (N_2091,N_1280,N_1919);
or U2092 (N_2092,N_1838,N_1495);
nand U2093 (N_2093,N_1411,N_1453);
xor U2094 (N_2094,N_1219,N_1635);
nor U2095 (N_2095,N_1136,N_1284);
and U2096 (N_2096,N_1164,N_1734);
nand U2097 (N_2097,N_1743,N_1952);
xnor U2098 (N_2098,N_1157,N_1522);
nor U2099 (N_2099,N_1672,N_1118);
nor U2100 (N_2100,N_1725,N_1826);
or U2101 (N_2101,N_1621,N_1899);
nor U2102 (N_2102,N_1844,N_1528);
and U2103 (N_2103,N_1677,N_1892);
or U2104 (N_2104,N_1890,N_1739);
nor U2105 (N_2105,N_1619,N_1054);
and U2106 (N_2106,N_1895,N_1816);
nor U2107 (N_2107,N_1084,N_1666);
xor U2108 (N_2108,N_1189,N_1088);
nand U2109 (N_2109,N_1182,N_1001);
or U2110 (N_2110,N_1149,N_1425);
nor U2111 (N_2111,N_1610,N_1897);
nor U2112 (N_2112,N_1207,N_1991);
nand U2113 (N_2113,N_1430,N_1471);
and U2114 (N_2114,N_1346,N_1586);
nand U2115 (N_2115,N_1151,N_1426);
nand U2116 (N_2116,N_1097,N_1428);
nor U2117 (N_2117,N_1384,N_1094);
nand U2118 (N_2118,N_1220,N_1102);
nand U2119 (N_2119,N_1537,N_1958);
or U2120 (N_2120,N_1211,N_1772);
or U2121 (N_2121,N_1110,N_1465);
and U2122 (N_2122,N_1520,N_1085);
nor U2123 (N_2123,N_1534,N_1710);
nor U2124 (N_2124,N_1571,N_1185);
or U2125 (N_2125,N_1079,N_1720);
and U2126 (N_2126,N_1756,N_1565);
xnor U2127 (N_2127,N_1287,N_1273);
nand U2128 (N_2128,N_1068,N_1993);
nand U2129 (N_2129,N_1256,N_1546);
or U2130 (N_2130,N_1312,N_1086);
or U2131 (N_2131,N_1405,N_1073);
or U2132 (N_2132,N_1884,N_1808);
xor U2133 (N_2133,N_1476,N_1229);
xor U2134 (N_2134,N_1736,N_1951);
nor U2135 (N_2135,N_1560,N_1938);
nand U2136 (N_2136,N_1988,N_1278);
nand U2137 (N_2137,N_1995,N_1393);
or U2138 (N_2138,N_1414,N_1840);
xor U2139 (N_2139,N_1254,N_1922);
nand U2140 (N_2140,N_1193,N_1459);
or U2141 (N_2141,N_1759,N_1552);
nor U2142 (N_2142,N_1053,N_1321);
or U2143 (N_2143,N_1566,N_1512);
nand U2144 (N_2144,N_1748,N_1749);
nand U2145 (N_2145,N_1294,N_1467);
and U2146 (N_2146,N_1954,N_1587);
and U2147 (N_2147,N_1934,N_1557);
nand U2148 (N_2148,N_1022,N_1197);
or U2149 (N_2149,N_1859,N_1093);
nand U2150 (N_2150,N_1925,N_1352);
and U2151 (N_2151,N_1600,N_1235);
and U2152 (N_2152,N_1741,N_1777);
nor U2153 (N_2153,N_1615,N_1567);
xnor U2154 (N_2154,N_1719,N_1841);
or U2155 (N_2155,N_1265,N_1732);
xor U2156 (N_2156,N_1961,N_1900);
nor U2157 (N_2157,N_1402,N_1075);
nor U2158 (N_2158,N_1452,N_1413);
xor U2159 (N_2159,N_1391,N_1589);
or U2160 (N_2160,N_1510,N_1018);
or U2161 (N_2161,N_1106,N_1042);
nor U2162 (N_2162,N_1788,N_1134);
and U2163 (N_2163,N_1667,N_1195);
xnor U2164 (N_2164,N_1689,N_1889);
nor U2165 (N_2165,N_1810,N_1024);
and U2166 (N_2166,N_1576,N_1901);
or U2167 (N_2167,N_1947,N_1336);
nand U2168 (N_2168,N_1470,N_1851);
or U2169 (N_2169,N_1472,N_1887);
or U2170 (N_2170,N_1507,N_1545);
or U2171 (N_2171,N_1996,N_1854);
nand U2172 (N_2172,N_1578,N_1762);
nand U2173 (N_2173,N_1964,N_1330);
nand U2174 (N_2174,N_1717,N_1077);
and U2175 (N_2175,N_1742,N_1354);
nand U2176 (N_2176,N_1544,N_1424);
or U2177 (N_2177,N_1701,N_1685);
nand U2178 (N_2178,N_1153,N_1807);
and U2179 (N_2179,N_1021,N_1323);
xnor U2180 (N_2180,N_1441,N_1833);
xor U2181 (N_2181,N_1251,N_1709);
xor U2182 (N_2182,N_1454,N_1237);
nand U2183 (N_2183,N_1642,N_1523);
and U2184 (N_2184,N_1201,N_1095);
or U2185 (N_2185,N_1983,N_1296);
xnor U2186 (N_2186,N_1058,N_1269);
and U2187 (N_2187,N_1963,N_1656);
or U2188 (N_2188,N_1852,N_1796);
or U2189 (N_2189,N_1167,N_1222);
nand U2190 (N_2190,N_1939,N_1674);
and U2191 (N_2191,N_1015,N_1598);
nand U2192 (N_2192,N_1555,N_1526);
or U2193 (N_2193,N_1607,N_1849);
and U2194 (N_2194,N_1886,N_1155);
xor U2195 (N_2195,N_1654,N_1098);
nand U2196 (N_2196,N_1318,N_1005);
or U2197 (N_2197,N_1568,N_1799);
xor U2198 (N_2198,N_1204,N_1401);
or U2199 (N_2199,N_1314,N_1609);
nor U2200 (N_2200,N_1398,N_1596);
nor U2201 (N_2201,N_1403,N_1694);
nor U2202 (N_2202,N_1409,N_1180);
xor U2203 (N_2203,N_1101,N_1640);
xnor U2204 (N_2204,N_1553,N_1582);
nor U2205 (N_2205,N_1691,N_1888);
xnor U2206 (N_2206,N_1767,N_1797);
nor U2207 (N_2207,N_1646,N_1248);
nor U2208 (N_2208,N_1918,N_1366);
or U2209 (N_2209,N_1558,N_1026);
nor U2210 (N_2210,N_1806,N_1940);
xnor U2211 (N_2211,N_1203,N_1766);
or U2212 (N_2212,N_1399,N_1039);
xnor U2213 (N_2213,N_1542,N_1194);
and U2214 (N_2214,N_1577,N_1967);
xnor U2215 (N_2215,N_1023,N_1987);
xor U2216 (N_2216,N_1295,N_1225);
nand U2217 (N_2217,N_1397,N_1910);
nor U2218 (N_2218,N_1062,N_1357);
and U2219 (N_2219,N_1521,N_1198);
or U2220 (N_2220,N_1360,N_1714);
and U2221 (N_2221,N_1067,N_1913);
nor U2222 (N_2222,N_1342,N_1092);
nor U2223 (N_2223,N_1322,N_1529);
nand U2224 (N_2224,N_1059,N_1381);
xor U2225 (N_2225,N_1724,N_1930);
xor U2226 (N_2226,N_1712,N_1141);
and U2227 (N_2227,N_1390,N_1463);
nand U2228 (N_2228,N_1916,N_1290);
xnor U2229 (N_2229,N_1885,N_1965);
nor U2230 (N_2230,N_1032,N_1175);
and U2231 (N_2231,N_1395,N_1232);
nor U2232 (N_2232,N_1090,N_1408);
and U2233 (N_2233,N_1539,N_1066);
and U2234 (N_2234,N_1746,N_1045);
nand U2235 (N_2235,N_1181,N_1985);
xor U2236 (N_2236,N_1324,N_1006);
nand U2237 (N_2237,N_1862,N_1769);
nand U2238 (N_2238,N_1879,N_1733);
nand U2239 (N_2239,N_1641,N_1873);
and U2240 (N_2240,N_1931,N_1121);
or U2241 (N_2241,N_1949,N_1339);
nor U2242 (N_2242,N_1678,N_1475);
nor U2243 (N_2243,N_1263,N_1602);
nand U2244 (N_2244,N_1986,N_1639);
and U2245 (N_2245,N_1331,N_1373);
nor U2246 (N_2246,N_1257,N_1599);
and U2247 (N_2247,N_1998,N_1626);
nand U2248 (N_2248,N_1455,N_1653);
nor U2249 (N_2249,N_1658,N_1754);
and U2250 (N_2250,N_1113,N_1948);
xor U2251 (N_2251,N_1903,N_1298);
nor U2252 (N_2252,N_1353,N_1064);
nand U2253 (N_2253,N_1911,N_1768);
xor U2254 (N_2254,N_1627,N_1213);
xnor U2255 (N_2255,N_1907,N_1396);
or U2256 (N_2256,N_1835,N_1010);
nand U2257 (N_2257,N_1538,N_1781);
nor U2258 (N_2258,N_1942,N_1158);
nor U2259 (N_2259,N_1392,N_1569);
nand U2260 (N_2260,N_1205,N_1973);
nor U2261 (N_2261,N_1518,N_1527);
nand U2262 (N_2262,N_1726,N_1186);
nor U2263 (N_2263,N_1776,N_1981);
and U2264 (N_2264,N_1519,N_1620);
nand U2265 (N_2265,N_1249,N_1530);
xor U2266 (N_2266,N_1301,N_1313);
xor U2267 (N_2267,N_1129,N_1531);
nor U2268 (N_2268,N_1792,N_1675);
nand U2269 (N_2269,N_1069,N_1131);
nor U2270 (N_2270,N_1362,N_1923);
nor U2271 (N_2271,N_1588,N_1200);
nand U2272 (N_2272,N_1340,N_1437);
or U2273 (N_2273,N_1462,N_1209);
nand U2274 (N_2274,N_1597,N_1380);
nor U2275 (N_2275,N_1696,N_1536);
nor U2276 (N_2276,N_1894,N_1305);
xnor U2277 (N_2277,N_1843,N_1326);
and U2278 (N_2278,N_1611,N_1738);
nand U2279 (N_2279,N_1634,N_1905);
nand U2280 (N_2280,N_1072,N_1850);
nand U2281 (N_2281,N_1215,N_1159);
nand U2282 (N_2282,N_1601,N_1135);
nand U2283 (N_2283,N_1379,N_1815);
nand U2284 (N_2284,N_1479,N_1982);
or U2285 (N_2285,N_1028,N_1486);
or U2286 (N_2286,N_1771,N_1169);
and U2287 (N_2287,N_1099,N_1474);
or U2288 (N_2288,N_1375,N_1030);
xor U2289 (N_2289,N_1143,N_1303);
or U2290 (N_2290,N_1962,N_1574);
or U2291 (N_2291,N_1103,N_1580);
nand U2292 (N_2292,N_1950,N_1543);
nor U2293 (N_2293,N_1645,N_1456);
nor U2294 (N_2294,N_1881,N_1780);
or U2295 (N_2295,N_1382,N_1713);
or U2296 (N_2296,N_1896,N_1049);
xor U2297 (N_2297,N_1488,N_1957);
nor U2298 (N_2298,N_1517,N_1761);
and U2299 (N_2299,N_1585,N_1126);
nand U2300 (N_2300,N_1385,N_1458);
and U2301 (N_2301,N_1926,N_1660);
nor U2302 (N_2302,N_1216,N_1262);
nand U2303 (N_2303,N_1124,N_1990);
xnor U2304 (N_2304,N_1082,N_1590);
and U2305 (N_2305,N_1108,N_1718);
nand U2306 (N_2306,N_1348,N_1187);
nor U2307 (N_2307,N_1613,N_1283);
or U2308 (N_2308,N_1883,N_1811);
nand U2309 (N_2309,N_1809,N_1171);
xnor U2310 (N_2310,N_1757,N_1060);
nor U2311 (N_2311,N_1306,N_1764);
and U2312 (N_2312,N_1004,N_1744);
xor U2313 (N_2313,N_1698,N_1008);
nor U2314 (N_2314,N_1297,N_1832);
and U2315 (N_2315,N_1935,N_1089);
or U2316 (N_2316,N_1866,N_1702);
nand U2317 (N_2317,N_1316,N_1774);
or U2318 (N_2318,N_1540,N_1535);
and U2319 (N_2319,N_1007,N_1464);
nor U2320 (N_2320,N_1044,N_1206);
xnor U2321 (N_2321,N_1343,N_1081);
or U2322 (N_2322,N_1550,N_1813);
xor U2323 (N_2323,N_1460,N_1775);
and U2324 (N_2324,N_1994,N_1604);
xnor U2325 (N_2325,N_1145,N_1847);
and U2326 (N_2326,N_1722,N_1992);
and U2327 (N_2327,N_1633,N_1477);
xnor U2328 (N_2328,N_1355,N_1584);
or U2329 (N_2329,N_1105,N_1422);
and U2330 (N_2330,N_1315,N_1842);
xnor U2331 (N_2331,N_1114,N_1140);
and U2332 (N_2332,N_1791,N_1115);
nand U2333 (N_2333,N_1908,N_1891);
or U2334 (N_2334,N_1848,N_1328);
nor U2335 (N_2335,N_1830,N_1984);
and U2336 (N_2336,N_1202,N_1929);
nand U2337 (N_2337,N_1502,N_1867);
nor U2338 (N_2338,N_1014,N_1857);
xnor U2339 (N_2339,N_1728,N_1697);
and U2340 (N_2340,N_1127,N_1078);
and U2341 (N_2341,N_1188,N_1266);
xor U2342 (N_2342,N_1484,N_1831);
nand U2343 (N_2343,N_1394,N_1999);
and U2344 (N_2344,N_1977,N_1882);
or U2345 (N_2345,N_1956,N_1142);
and U2346 (N_2346,N_1137,N_1716);
nor U2347 (N_2347,N_1020,N_1347);
or U2348 (N_2348,N_1174,N_1490);
or U2349 (N_2349,N_1310,N_1563);
and U2350 (N_2350,N_1191,N_1632);
nor U2351 (N_2351,N_1275,N_1670);
and U2352 (N_2352,N_1461,N_1122);
xor U2353 (N_2353,N_1793,N_1647);
xnor U2354 (N_2354,N_1755,N_1406);
nand U2355 (N_2355,N_1332,N_1856);
or U2356 (N_2356,N_1236,N_1335);
xor U2357 (N_2357,N_1376,N_1221);
nor U2358 (N_2358,N_1912,N_1351);
or U2359 (N_2359,N_1438,N_1444);
nand U2360 (N_2360,N_1872,N_1119);
or U2361 (N_2361,N_1242,N_1684);
nor U2362 (N_2362,N_1513,N_1904);
or U2363 (N_2363,N_1302,N_1541);
and U2364 (N_2364,N_1760,N_1214);
or U2365 (N_2365,N_1100,N_1592);
xor U2366 (N_2366,N_1629,N_1747);
nand U2367 (N_2367,N_1239,N_1933);
or U2368 (N_2368,N_1637,N_1649);
or U2369 (N_2369,N_1291,N_1345);
or U2370 (N_2370,N_1144,N_1644);
xnor U2371 (N_2371,N_1735,N_1966);
and U2372 (N_2372,N_1259,N_1763);
nor U2373 (N_2373,N_1876,N_1622);
xor U2374 (N_2374,N_1035,N_1499);
nor U2375 (N_2375,N_1250,N_1794);
or U2376 (N_2376,N_1041,N_1027);
and U2377 (N_2377,N_1359,N_1989);
or U2378 (N_2378,N_1524,N_1758);
nand U2379 (N_2379,N_1612,N_1688);
nor U2380 (N_2380,N_1556,N_1432);
and U2381 (N_2381,N_1051,N_1551);
or U2382 (N_2382,N_1076,N_1170);
and U2383 (N_2383,N_1943,N_1770);
nand U2384 (N_2384,N_1415,N_1429);
nand U2385 (N_2385,N_1827,N_1277);
or U2386 (N_2386,N_1163,N_1276);
and U2387 (N_2387,N_1487,N_1628);
nor U2388 (N_2388,N_1699,N_1029);
nor U2389 (N_2389,N_1165,N_1686);
nor U2390 (N_2390,N_1795,N_1959);
nor U2391 (N_2391,N_1046,N_1614);
nor U2392 (N_2392,N_1148,N_1668);
and U2393 (N_2393,N_1052,N_1975);
or U2394 (N_2394,N_1564,N_1341);
xor U2395 (N_2395,N_1501,N_1270);
nand U2396 (N_2396,N_1445,N_1814);
xnor U2397 (N_2397,N_1162,N_1638);
xor U2398 (N_2398,N_1695,N_1057);
nor U2399 (N_2399,N_1450,N_1002);
or U2400 (N_2400,N_1388,N_1112);
nand U2401 (N_2401,N_1877,N_1218);
and U2402 (N_2402,N_1818,N_1706);
xnor U2403 (N_2403,N_1778,N_1974);
xor U2404 (N_2404,N_1096,N_1245);
nor U2405 (N_2405,N_1074,N_1418);
xnor U2406 (N_2406,N_1779,N_1338);
xor U2407 (N_2407,N_1679,N_1238);
nor U2408 (N_2408,N_1491,N_1412);
or U2409 (N_2409,N_1729,N_1798);
nand U2410 (N_2410,N_1389,N_1154);
xor U2411 (N_2411,N_1864,N_1561);
nor U2412 (N_2412,N_1361,N_1308);
or U2413 (N_2413,N_1511,N_1083);
nor U2414 (N_2414,N_1033,N_1208);
and U2415 (N_2415,N_1494,N_1824);
nor U2416 (N_2416,N_1648,N_1979);
nand U2417 (N_2417,N_1070,N_1478);
xnor U2418 (N_2418,N_1061,N_1150);
and U2419 (N_2419,N_1307,N_1509);
nand U2420 (N_2420,N_1417,N_1594);
and U2421 (N_2421,N_1439,N_1837);
xor U2422 (N_2422,N_1274,N_1087);
nand U2423 (N_2423,N_1572,N_1272);
nor U2424 (N_2424,N_1853,N_1693);
or U2425 (N_2425,N_1309,N_1019);
and U2426 (N_2426,N_1643,N_1909);
and U2427 (N_2427,N_1839,N_1921);
and U2428 (N_2428,N_1427,N_1822);
nand U2429 (N_2429,N_1941,N_1906);
nor U2430 (N_2430,N_1817,N_1179);
xnor U2431 (N_2431,N_1605,N_1241);
xnor U2432 (N_2432,N_1293,N_1819);
and U2433 (N_2433,N_1009,N_1228);
nor U2434 (N_2434,N_1130,N_1120);
and U2435 (N_2435,N_1281,N_1410);
xor U2436 (N_2436,N_1690,N_1559);
or U2437 (N_2437,N_1434,N_1945);
xnor U2438 (N_2438,N_1631,N_1944);
and U2439 (N_2439,N_1765,N_1730);
xor U2440 (N_2440,N_1617,N_1655);
nand U2441 (N_2441,N_1056,N_1673);
and U2442 (N_2442,N_1400,N_1651);
nand U2443 (N_2443,N_1789,N_1737);
nor U2444 (N_2444,N_1358,N_1953);
xnor U2445 (N_2445,N_1055,N_1801);
nand U2446 (N_2446,N_1650,N_1183);
nor U2447 (N_2447,N_1047,N_1230);
nor U2448 (N_2448,N_1865,N_1369);
and U2449 (N_2449,N_1247,N_1407);
nand U2450 (N_2450,N_1936,N_1285);
nand U2451 (N_2451,N_1825,N_1011);
nor U2452 (N_2452,N_1132,N_1731);
nand U2453 (N_2453,N_1785,N_1721);
and U2454 (N_2454,N_1329,N_1178);
or U2455 (N_2455,N_1446,N_1625);
or U2456 (N_2456,N_1665,N_1377);
nor U2457 (N_2457,N_1525,N_1443);
and U2458 (N_2458,N_1970,N_1173);
or U2459 (N_2459,N_1508,N_1017);
xnor U2460 (N_2460,N_1676,N_1327);
and U2461 (N_2461,N_1416,N_1282);
or U2462 (N_2462,N_1003,N_1669);
or U2463 (N_2463,N_1255,N_1333);
nand U2464 (N_2464,N_1579,N_1932);
xnor U2465 (N_2465,N_1703,N_1924);
nand U2466 (N_2466,N_1133,N_1955);
or U2467 (N_2467,N_1319,N_1199);
nand U2468 (N_2468,N_1875,N_1727);
nor U2469 (N_2469,N_1623,N_1107);
xor U2470 (N_2470,N_1048,N_1846);
xor U2471 (N_2471,N_1624,N_1034);
nor U2472 (N_2472,N_1349,N_1246);
xnor U2473 (N_2473,N_1233,N_1037);
xor U2474 (N_2474,N_1920,N_1790);
and U2475 (N_2475,N_1547,N_1365);
nand U2476 (N_2476,N_1583,N_1104);
nor U2477 (N_2477,N_1368,N_1878);
or U2478 (N_2478,N_1031,N_1740);
xor U2479 (N_2479,N_1821,N_1253);
xor U2480 (N_2480,N_1773,N_1532);
or U2481 (N_2481,N_1123,N_1466);
xnor U2482 (N_2482,N_1917,N_1231);
or U2483 (N_2483,N_1705,N_1299);
and U2484 (N_2484,N_1606,N_1419);
nor U2485 (N_2485,N_1554,N_1514);
or U2486 (N_2486,N_1378,N_1374);
or U2487 (N_2487,N_1858,N_1431);
nor U2488 (N_2488,N_1210,N_1260);
or U2489 (N_2489,N_1447,N_1177);
nor U2490 (N_2490,N_1387,N_1139);
nor U2491 (N_2491,N_1481,N_1595);
nor U2492 (N_2492,N_1146,N_1109);
xor U2493 (N_2493,N_1025,N_1871);
and U2494 (N_2494,N_1968,N_1138);
xor U2495 (N_2495,N_1752,N_1704);
or U2496 (N_2496,N_1515,N_1829);
and U2497 (N_2497,N_1267,N_1692);
and U2498 (N_2498,N_1161,N_1483);
or U2499 (N_2499,N_1618,N_1065);
nand U2500 (N_2500,N_1482,N_1113);
nand U2501 (N_2501,N_1179,N_1719);
or U2502 (N_2502,N_1598,N_1597);
nor U2503 (N_2503,N_1369,N_1841);
nand U2504 (N_2504,N_1442,N_1698);
xnor U2505 (N_2505,N_1885,N_1509);
xnor U2506 (N_2506,N_1121,N_1751);
or U2507 (N_2507,N_1121,N_1685);
nor U2508 (N_2508,N_1991,N_1814);
and U2509 (N_2509,N_1084,N_1107);
nand U2510 (N_2510,N_1303,N_1417);
or U2511 (N_2511,N_1479,N_1868);
nor U2512 (N_2512,N_1245,N_1322);
nor U2513 (N_2513,N_1606,N_1241);
or U2514 (N_2514,N_1621,N_1536);
nor U2515 (N_2515,N_1544,N_1076);
nand U2516 (N_2516,N_1638,N_1121);
nor U2517 (N_2517,N_1827,N_1092);
nor U2518 (N_2518,N_1490,N_1706);
nor U2519 (N_2519,N_1427,N_1815);
or U2520 (N_2520,N_1135,N_1959);
and U2521 (N_2521,N_1408,N_1040);
or U2522 (N_2522,N_1196,N_1787);
and U2523 (N_2523,N_1081,N_1135);
and U2524 (N_2524,N_1484,N_1191);
nor U2525 (N_2525,N_1877,N_1799);
nand U2526 (N_2526,N_1251,N_1427);
and U2527 (N_2527,N_1405,N_1987);
nor U2528 (N_2528,N_1921,N_1664);
nand U2529 (N_2529,N_1012,N_1958);
and U2530 (N_2530,N_1992,N_1584);
nand U2531 (N_2531,N_1639,N_1991);
nand U2532 (N_2532,N_1220,N_1104);
and U2533 (N_2533,N_1743,N_1862);
nand U2534 (N_2534,N_1311,N_1876);
nand U2535 (N_2535,N_1835,N_1258);
xor U2536 (N_2536,N_1658,N_1123);
nand U2537 (N_2537,N_1322,N_1490);
nand U2538 (N_2538,N_1248,N_1121);
nor U2539 (N_2539,N_1797,N_1682);
nor U2540 (N_2540,N_1126,N_1245);
xnor U2541 (N_2541,N_1802,N_1680);
and U2542 (N_2542,N_1884,N_1489);
or U2543 (N_2543,N_1497,N_1184);
nor U2544 (N_2544,N_1374,N_1216);
or U2545 (N_2545,N_1181,N_1918);
or U2546 (N_2546,N_1271,N_1443);
xnor U2547 (N_2547,N_1542,N_1685);
nand U2548 (N_2548,N_1919,N_1802);
or U2549 (N_2549,N_1547,N_1061);
nor U2550 (N_2550,N_1674,N_1495);
and U2551 (N_2551,N_1079,N_1445);
nand U2552 (N_2552,N_1172,N_1252);
and U2553 (N_2553,N_1372,N_1425);
nor U2554 (N_2554,N_1746,N_1977);
xor U2555 (N_2555,N_1590,N_1711);
xnor U2556 (N_2556,N_1910,N_1179);
xnor U2557 (N_2557,N_1631,N_1517);
or U2558 (N_2558,N_1356,N_1804);
xnor U2559 (N_2559,N_1148,N_1221);
xor U2560 (N_2560,N_1822,N_1877);
nor U2561 (N_2561,N_1553,N_1297);
and U2562 (N_2562,N_1136,N_1094);
and U2563 (N_2563,N_1868,N_1698);
xnor U2564 (N_2564,N_1212,N_1331);
nor U2565 (N_2565,N_1846,N_1869);
or U2566 (N_2566,N_1012,N_1036);
and U2567 (N_2567,N_1695,N_1131);
or U2568 (N_2568,N_1368,N_1762);
and U2569 (N_2569,N_1975,N_1235);
xnor U2570 (N_2570,N_1827,N_1886);
or U2571 (N_2571,N_1742,N_1131);
or U2572 (N_2572,N_1062,N_1599);
or U2573 (N_2573,N_1499,N_1221);
xnor U2574 (N_2574,N_1607,N_1233);
xor U2575 (N_2575,N_1251,N_1166);
and U2576 (N_2576,N_1417,N_1861);
and U2577 (N_2577,N_1196,N_1352);
and U2578 (N_2578,N_1987,N_1157);
or U2579 (N_2579,N_1591,N_1282);
nor U2580 (N_2580,N_1755,N_1144);
or U2581 (N_2581,N_1872,N_1625);
xor U2582 (N_2582,N_1727,N_1229);
nand U2583 (N_2583,N_1075,N_1812);
or U2584 (N_2584,N_1147,N_1975);
or U2585 (N_2585,N_1150,N_1501);
nor U2586 (N_2586,N_1583,N_1653);
xor U2587 (N_2587,N_1189,N_1350);
xor U2588 (N_2588,N_1369,N_1649);
xnor U2589 (N_2589,N_1855,N_1263);
nor U2590 (N_2590,N_1263,N_1259);
xnor U2591 (N_2591,N_1943,N_1598);
and U2592 (N_2592,N_1504,N_1109);
xor U2593 (N_2593,N_1537,N_1743);
and U2594 (N_2594,N_1797,N_1955);
or U2595 (N_2595,N_1281,N_1656);
nand U2596 (N_2596,N_1773,N_1087);
xnor U2597 (N_2597,N_1164,N_1990);
nor U2598 (N_2598,N_1763,N_1411);
nand U2599 (N_2599,N_1221,N_1179);
nand U2600 (N_2600,N_1190,N_1497);
nor U2601 (N_2601,N_1847,N_1380);
or U2602 (N_2602,N_1595,N_1920);
or U2603 (N_2603,N_1537,N_1700);
nand U2604 (N_2604,N_1561,N_1229);
nand U2605 (N_2605,N_1521,N_1385);
nor U2606 (N_2606,N_1867,N_1100);
nor U2607 (N_2607,N_1276,N_1222);
or U2608 (N_2608,N_1152,N_1246);
or U2609 (N_2609,N_1113,N_1916);
xor U2610 (N_2610,N_1282,N_1090);
and U2611 (N_2611,N_1695,N_1920);
or U2612 (N_2612,N_1965,N_1430);
and U2613 (N_2613,N_1346,N_1437);
nor U2614 (N_2614,N_1796,N_1402);
xor U2615 (N_2615,N_1504,N_1977);
nand U2616 (N_2616,N_1481,N_1620);
nand U2617 (N_2617,N_1278,N_1637);
and U2618 (N_2618,N_1735,N_1158);
xor U2619 (N_2619,N_1096,N_1030);
nor U2620 (N_2620,N_1864,N_1848);
and U2621 (N_2621,N_1043,N_1091);
or U2622 (N_2622,N_1523,N_1044);
nor U2623 (N_2623,N_1396,N_1356);
nand U2624 (N_2624,N_1563,N_1377);
xnor U2625 (N_2625,N_1058,N_1827);
nand U2626 (N_2626,N_1421,N_1967);
nor U2627 (N_2627,N_1980,N_1120);
nand U2628 (N_2628,N_1211,N_1245);
or U2629 (N_2629,N_1797,N_1902);
xor U2630 (N_2630,N_1129,N_1087);
nor U2631 (N_2631,N_1840,N_1235);
or U2632 (N_2632,N_1808,N_1097);
and U2633 (N_2633,N_1738,N_1234);
or U2634 (N_2634,N_1080,N_1791);
xor U2635 (N_2635,N_1499,N_1980);
xor U2636 (N_2636,N_1954,N_1797);
xnor U2637 (N_2637,N_1860,N_1134);
and U2638 (N_2638,N_1194,N_1979);
xor U2639 (N_2639,N_1611,N_1638);
nand U2640 (N_2640,N_1949,N_1236);
nand U2641 (N_2641,N_1378,N_1097);
nand U2642 (N_2642,N_1330,N_1241);
or U2643 (N_2643,N_1371,N_1364);
xor U2644 (N_2644,N_1411,N_1366);
and U2645 (N_2645,N_1408,N_1231);
and U2646 (N_2646,N_1231,N_1869);
nand U2647 (N_2647,N_1826,N_1113);
or U2648 (N_2648,N_1820,N_1611);
and U2649 (N_2649,N_1191,N_1043);
nand U2650 (N_2650,N_1168,N_1109);
xor U2651 (N_2651,N_1926,N_1178);
nand U2652 (N_2652,N_1553,N_1539);
xnor U2653 (N_2653,N_1216,N_1944);
and U2654 (N_2654,N_1010,N_1702);
nor U2655 (N_2655,N_1667,N_1791);
nand U2656 (N_2656,N_1680,N_1908);
xnor U2657 (N_2657,N_1161,N_1665);
nand U2658 (N_2658,N_1295,N_1204);
xor U2659 (N_2659,N_1326,N_1827);
and U2660 (N_2660,N_1547,N_1665);
xor U2661 (N_2661,N_1535,N_1207);
nand U2662 (N_2662,N_1758,N_1273);
or U2663 (N_2663,N_1489,N_1400);
nor U2664 (N_2664,N_1271,N_1902);
and U2665 (N_2665,N_1759,N_1990);
nand U2666 (N_2666,N_1882,N_1512);
or U2667 (N_2667,N_1110,N_1632);
or U2668 (N_2668,N_1857,N_1665);
nand U2669 (N_2669,N_1630,N_1279);
nand U2670 (N_2670,N_1286,N_1491);
nor U2671 (N_2671,N_1726,N_1646);
and U2672 (N_2672,N_1881,N_1242);
or U2673 (N_2673,N_1188,N_1723);
nand U2674 (N_2674,N_1859,N_1358);
and U2675 (N_2675,N_1937,N_1144);
or U2676 (N_2676,N_1288,N_1041);
xnor U2677 (N_2677,N_1611,N_1177);
or U2678 (N_2678,N_1571,N_1707);
and U2679 (N_2679,N_1149,N_1254);
and U2680 (N_2680,N_1328,N_1796);
or U2681 (N_2681,N_1771,N_1548);
nand U2682 (N_2682,N_1816,N_1621);
xor U2683 (N_2683,N_1033,N_1059);
nand U2684 (N_2684,N_1204,N_1624);
nor U2685 (N_2685,N_1794,N_1745);
xor U2686 (N_2686,N_1073,N_1771);
nor U2687 (N_2687,N_1350,N_1811);
nand U2688 (N_2688,N_1132,N_1470);
xnor U2689 (N_2689,N_1732,N_1494);
or U2690 (N_2690,N_1617,N_1450);
and U2691 (N_2691,N_1464,N_1395);
nor U2692 (N_2692,N_1309,N_1000);
and U2693 (N_2693,N_1793,N_1450);
or U2694 (N_2694,N_1815,N_1267);
or U2695 (N_2695,N_1380,N_1659);
xor U2696 (N_2696,N_1188,N_1830);
xor U2697 (N_2697,N_1262,N_1249);
nand U2698 (N_2698,N_1102,N_1197);
nand U2699 (N_2699,N_1652,N_1732);
and U2700 (N_2700,N_1223,N_1898);
or U2701 (N_2701,N_1392,N_1244);
nand U2702 (N_2702,N_1841,N_1097);
nand U2703 (N_2703,N_1552,N_1928);
nand U2704 (N_2704,N_1435,N_1164);
nand U2705 (N_2705,N_1819,N_1864);
and U2706 (N_2706,N_1468,N_1353);
nand U2707 (N_2707,N_1996,N_1693);
and U2708 (N_2708,N_1080,N_1436);
or U2709 (N_2709,N_1729,N_1677);
or U2710 (N_2710,N_1935,N_1739);
nand U2711 (N_2711,N_1196,N_1991);
nand U2712 (N_2712,N_1450,N_1738);
xnor U2713 (N_2713,N_1392,N_1610);
and U2714 (N_2714,N_1397,N_1529);
or U2715 (N_2715,N_1250,N_1523);
xnor U2716 (N_2716,N_1434,N_1780);
nand U2717 (N_2717,N_1716,N_1286);
nand U2718 (N_2718,N_1322,N_1449);
or U2719 (N_2719,N_1602,N_1015);
and U2720 (N_2720,N_1340,N_1944);
nor U2721 (N_2721,N_1788,N_1787);
or U2722 (N_2722,N_1979,N_1201);
or U2723 (N_2723,N_1407,N_1583);
xor U2724 (N_2724,N_1917,N_1133);
nand U2725 (N_2725,N_1522,N_1327);
or U2726 (N_2726,N_1032,N_1325);
and U2727 (N_2727,N_1015,N_1674);
nor U2728 (N_2728,N_1567,N_1950);
or U2729 (N_2729,N_1673,N_1822);
and U2730 (N_2730,N_1100,N_1282);
nand U2731 (N_2731,N_1811,N_1135);
and U2732 (N_2732,N_1490,N_1487);
nand U2733 (N_2733,N_1602,N_1097);
or U2734 (N_2734,N_1504,N_1544);
nand U2735 (N_2735,N_1595,N_1242);
and U2736 (N_2736,N_1827,N_1440);
or U2737 (N_2737,N_1407,N_1587);
or U2738 (N_2738,N_1593,N_1913);
nor U2739 (N_2739,N_1966,N_1588);
and U2740 (N_2740,N_1233,N_1875);
nand U2741 (N_2741,N_1089,N_1277);
and U2742 (N_2742,N_1433,N_1206);
or U2743 (N_2743,N_1314,N_1455);
nor U2744 (N_2744,N_1291,N_1785);
nand U2745 (N_2745,N_1876,N_1246);
nand U2746 (N_2746,N_1447,N_1341);
nand U2747 (N_2747,N_1710,N_1576);
nor U2748 (N_2748,N_1870,N_1529);
nand U2749 (N_2749,N_1200,N_1923);
xor U2750 (N_2750,N_1537,N_1880);
nand U2751 (N_2751,N_1095,N_1216);
nor U2752 (N_2752,N_1462,N_1330);
or U2753 (N_2753,N_1110,N_1945);
nand U2754 (N_2754,N_1256,N_1362);
and U2755 (N_2755,N_1363,N_1798);
and U2756 (N_2756,N_1998,N_1530);
xor U2757 (N_2757,N_1985,N_1049);
and U2758 (N_2758,N_1625,N_1670);
or U2759 (N_2759,N_1093,N_1146);
xor U2760 (N_2760,N_1103,N_1395);
nor U2761 (N_2761,N_1846,N_1052);
nand U2762 (N_2762,N_1482,N_1942);
nand U2763 (N_2763,N_1532,N_1573);
xor U2764 (N_2764,N_1362,N_1237);
xnor U2765 (N_2765,N_1291,N_1718);
and U2766 (N_2766,N_1308,N_1754);
nand U2767 (N_2767,N_1190,N_1694);
and U2768 (N_2768,N_1730,N_1826);
nand U2769 (N_2769,N_1903,N_1649);
nand U2770 (N_2770,N_1766,N_1947);
xnor U2771 (N_2771,N_1004,N_1865);
xor U2772 (N_2772,N_1424,N_1829);
or U2773 (N_2773,N_1108,N_1151);
and U2774 (N_2774,N_1749,N_1548);
nor U2775 (N_2775,N_1160,N_1594);
nand U2776 (N_2776,N_1405,N_1241);
nor U2777 (N_2777,N_1251,N_1361);
and U2778 (N_2778,N_1046,N_1986);
nand U2779 (N_2779,N_1527,N_1051);
or U2780 (N_2780,N_1744,N_1137);
xor U2781 (N_2781,N_1900,N_1905);
nor U2782 (N_2782,N_1878,N_1396);
xnor U2783 (N_2783,N_1593,N_1540);
nand U2784 (N_2784,N_1569,N_1833);
nor U2785 (N_2785,N_1489,N_1781);
xor U2786 (N_2786,N_1475,N_1721);
nor U2787 (N_2787,N_1940,N_1680);
nand U2788 (N_2788,N_1392,N_1145);
nand U2789 (N_2789,N_1657,N_1081);
xor U2790 (N_2790,N_1720,N_1221);
nand U2791 (N_2791,N_1668,N_1155);
or U2792 (N_2792,N_1361,N_1185);
or U2793 (N_2793,N_1642,N_1036);
nor U2794 (N_2794,N_1716,N_1783);
and U2795 (N_2795,N_1780,N_1541);
or U2796 (N_2796,N_1966,N_1511);
xor U2797 (N_2797,N_1077,N_1773);
and U2798 (N_2798,N_1263,N_1322);
xor U2799 (N_2799,N_1539,N_1362);
nor U2800 (N_2800,N_1580,N_1886);
xor U2801 (N_2801,N_1322,N_1618);
nand U2802 (N_2802,N_1037,N_1475);
xnor U2803 (N_2803,N_1715,N_1149);
or U2804 (N_2804,N_1190,N_1025);
nor U2805 (N_2805,N_1578,N_1595);
xor U2806 (N_2806,N_1624,N_1986);
xnor U2807 (N_2807,N_1329,N_1102);
or U2808 (N_2808,N_1346,N_1287);
nand U2809 (N_2809,N_1294,N_1339);
or U2810 (N_2810,N_1788,N_1256);
nor U2811 (N_2811,N_1711,N_1392);
or U2812 (N_2812,N_1627,N_1341);
nor U2813 (N_2813,N_1641,N_1404);
and U2814 (N_2814,N_1643,N_1326);
and U2815 (N_2815,N_1353,N_1262);
nand U2816 (N_2816,N_1259,N_1919);
nor U2817 (N_2817,N_1676,N_1429);
or U2818 (N_2818,N_1112,N_1875);
xor U2819 (N_2819,N_1825,N_1215);
nor U2820 (N_2820,N_1184,N_1568);
and U2821 (N_2821,N_1774,N_1984);
and U2822 (N_2822,N_1618,N_1349);
or U2823 (N_2823,N_1160,N_1408);
nand U2824 (N_2824,N_1587,N_1035);
nor U2825 (N_2825,N_1207,N_1695);
nor U2826 (N_2826,N_1814,N_1801);
or U2827 (N_2827,N_1870,N_1992);
or U2828 (N_2828,N_1290,N_1711);
or U2829 (N_2829,N_1934,N_1823);
nor U2830 (N_2830,N_1041,N_1097);
and U2831 (N_2831,N_1670,N_1574);
xnor U2832 (N_2832,N_1722,N_1431);
nand U2833 (N_2833,N_1861,N_1147);
and U2834 (N_2834,N_1619,N_1424);
nand U2835 (N_2835,N_1466,N_1897);
and U2836 (N_2836,N_1271,N_1573);
nand U2837 (N_2837,N_1194,N_1858);
xnor U2838 (N_2838,N_1358,N_1564);
nand U2839 (N_2839,N_1763,N_1278);
nor U2840 (N_2840,N_1875,N_1771);
xnor U2841 (N_2841,N_1719,N_1194);
nor U2842 (N_2842,N_1646,N_1133);
nand U2843 (N_2843,N_1961,N_1797);
nor U2844 (N_2844,N_1056,N_1844);
or U2845 (N_2845,N_1316,N_1211);
or U2846 (N_2846,N_1479,N_1601);
xnor U2847 (N_2847,N_1698,N_1752);
nor U2848 (N_2848,N_1712,N_1426);
xor U2849 (N_2849,N_1964,N_1146);
or U2850 (N_2850,N_1331,N_1406);
nor U2851 (N_2851,N_1605,N_1146);
xor U2852 (N_2852,N_1683,N_1090);
or U2853 (N_2853,N_1099,N_1244);
or U2854 (N_2854,N_1262,N_1850);
xor U2855 (N_2855,N_1066,N_1623);
or U2856 (N_2856,N_1985,N_1154);
nor U2857 (N_2857,N_1102,N_1231);
nor U2858 (N_2858,N_1538,N_1768);
or U2859 (N_2859,N_1158,N_1922);
nand U2860 (N_2860,N_1321,N_1365);
nor U2861 (N_2861,N_1630,N_1059);
or U2862 (N_2862,N_1637,N_1578);
nor U2863 (N_2863,N_1858,N_1443);
xnor U2864 (N_2864,N_1847,N_1184);
or U2865 (N_2865,N_1529,N_1855);
nand U2866 (N_2866,N_1237,N_1881);
or U2867 (N_2867,N_1351,N_1025);
or U2868 (N_2868,N_1380,N_1570);
xor U2869 (N_2869,N_1083,N_1532);
nand U2870 (N_2870,N_1865,N_1601);
nand U2871 (N_2871,N_1007,N_1542);
and U2872 (N_2872,N_1854,N_1462);
and U2873 (N_2873,N_1222,N_1751);
nand U2874 (N_2874,N_1858,N_1881);
or U2875 (N_2875,N_1627,N_1044);
or U2876 (N_2876,N_1255,N_1282);
xor U2877 (N_2877,N_1169,N_1616);
and U2878 (N_2878,N_1793,N_1054);
nor U2879 (N_2879,N_1967,N_1240);
or U2880 (N_2880,N_1934,N_1582);
nand U2881 (N_2881,N_1479,N_1049);
xnor U2882 (N_2882,N_1304,N_1164);
or U2883 (N_2883,N_1373,N_1966);
nand U2884 (N_2884,N_1323,N_1723);
or U2885 (N_2885,N_1258,N_1812);
nor U2886 (N_2886,N_1210,N_1143);
nand U2887 (N_2887,N_1086,N_1255);
nor U2888 (N_2888,N_1816,N_1963);
xnor U2889 (N_2889,N_1409,N_1355);
nand U2890 (N_2890,N_1690,N_1217);
nor U2891 (N_2891,N_1578,N_1869);
nand U2892 (N_2892,N_1307,N_1140);
or U2893 (N_2893,N_1852,N_1971);
nor U2894 (N_2894,N_1873,N_1379);
nand U2895 (N_2895,N_1906,N_1395);
nand U2896 (N_2896,N_1893,N_1033);
nor U2897 (N_2897,N_1106,N_1419);
or U2898 (N_2898,N_1972,N_1867);
xor U2899 (N_2899,N_1268,N_1920);
nand U2900 (N_2900,N_1329,N_1137);
nand U2901 (N_2901,N_1946,N_1860);
or U2902 (N_2902,N_1724,N_1683);
and U2903 (N_2903,N_1696,N_1442);
or U2904 (N_2904,N_1769,N_1303);
nand U2905 (N_2905,N_1259,N_1705);
and U2906 (N_2906,N_1843,N_1300);
xor U2907 (N_2907,N_1267,N_1584);
nand U2908 (N_2908,N_1752,N_1369);
nand U2909 (N_2909,N_1092,N_1927);
xor U2910 (N_2910,N_1345,N_1728);
and U2911 (N_2911,N_1533,N_1961);
xor U2912 (N_2912,N_1170,N_1119);
or U2913 (N_2913,N_1499,N_1461);
nor U2914 (N_2914,N_1816,N_1449);
or U2915 (N_2915,N_1843,N_1520);
or U2916 (N_2916,N_1373,N_1573);
and U2917 (N_2917,N_1427,N_1217);
or U2918 (N_2918,N_1542,N_1035);
or U2919 (N_2919,N_1937,N_1271);
xor U2920 (N_2920,N_1538,N_1324);
nor U2921 (N_2921,N_1305,N_1847);
or U2922 (N_2922,N_1905,N_1706);
nor U2923 (N_2923,N_1605,N_1727);
xor U2924 (N_2924,N_1190,N_1253);
and U2925 (N_2925,N_1342,N_1946);
nor U2926 (N_2926,N_1982,N_1590);
nor U2927 (N_2927,N_1151,N_1872);
nand U2928 (N_2928,N_1369,N_1664);
and U2929 (N_2929,N_1796,N_1944);
xnor U2930 (N_2930,N_1910,N_1614);
and U2931 (N_2931,N_1844,N_1432);
xor U2932 (N_2932,N_1202,N_1643);
xnor U2933 (N_2933,N_1140,N_1556);
nor U2934 (N_2934,N_1896,N_1304);
or U2935 (N_2935,N_1084,N_1927);
nand U2936 (N_2936,N_1968,N_1706);
xnor U2937 (N_2937,N_1354,N_1687);
nand U2938 (N_2938,N_1382,N_1893);
and U2939 (N_2939,N_1357,N_1889);
and U2940 (N_2940,N_1335,N_1415);
nor U2941 (N_2941,N_1087,N_1247);
xnor U2942 (N_2942,N_1357,N_1610);
xor U2943 (N_2943,N_1934,N_1615);
xor U2944 (N_2944,N_1484,N_1722);
nor U2945 (N_2945,N_1238,N_1626);
nand U2946 (N_2946,N_1701,N_1644);
xor U2947 (N_2947,N_1126,N_1181);
nand U2948 (N_2948,N_1511,N_1791);
or U2949 (N_2949,N_1496,N_1767);
nand U2950 (N_2950,N_1036,N_1758);
and U2951 (N_2951,N_1616,N_1441);
nor U2952 (N_2952,N_1582,N_1590);
xnor U2953 (N_2953,N_1293,N_1967);
and U2954 (N_2954,N_1688,N_1952);
nor U2955 (N_2955,N_1438,N_1113);
xor U2956 (N_2956,N_1331,N_1117);
nand U2957 (N_2957,N_1187,N_1062);
nor U2958 (N_2958,N_1911,N_1742);
or U2959 (N_2959,N_1565,N_1196);
nand U2960 (N_2960,N_1225,N_1698);
and U2961 (N_2961,N_1970,N_1890);
xnor U2962 (N_2962,N_1064,N_1340);
and U2963 (N_2963,N_1103,N_1249);
nor U2964 (N_2964,N_1333,N_1859);
xnor U2965 (N_2965,N_1319,N_1172);
nand U2966 (N_2966,N_1125,N_1131);
or U2967 (N_2967,N_1944,N_1901);
and U2968 (N_2968,N_1473,N_1773);
nor U2969 (N_2969,N_1727,N_1262);
and U2970 (N_2970,N_1554,N_1802);
nand U2971 (N_2971,N_1472,N_1807);
and U2972 (N_2972,N_1444,N_1608);
or U2973 (N_2973,N_1155,N_1389);
and U2974 (N_2974,N_1230,N_1074);
xor U2975 (N_2975,N_1501,N_1334);
nor U2976 (N_2976,N_1325,N_1707);
nor U2977 (N_2977,N_1455,N_1446);
nand U2978 (N_2978,N_1662,N_1314);
and U2979 (N_2979,N_1765,N_1944);
nand U2980 (N_2980,N_1180,N_1535);
nor U2981 (N_2981,N_1061,N_1215);
nor U2982 (N_2982,N_1502,N_1990);
or U2983 (N_2983,N_1937,N_1279);
and U2984 (N_2984,N_1440,N_1636);
nand U2985 (N_2985,N_1783,N_1983);
nor U2986 (N_2986,N_1483,N_1912);
xnor U2987 (N_2987,N_1062,N_1309);
or U2988 (N_2988,N_1223,N_1530);
xnor U2989 (N_2989,N_1252,N_1587);
xor U2990 (N_2990,N_1054,N_1155);
or U2991 (N_2991,N_1999,N_1055);
and U2992 (N_2992,N_1877,N_1038);
nand U2993 (N_2993,N_1864,N_1223);
xnor U2994 (N_2994,N_1947,N_1801);
nand U2995 (N_2995,N_1383,N_1459);
nor U2996 (N_2996,N_1452,N_1462);
or U2997 (N_2997,N_1390,N_1623);
nor U2998 (N_2998,N_1247,N_1376);
or U2999 (N_2999,N_1834,N_1749);
xor U3000 (N_3000,N_2682,N_2955);
nand U3001 (N_3001,N_2315,N_2549);
and U3002 (N_3002,N_2793,N_2543);
nand U3003 (N_3003,N_2102,N_2910);
nand U3004 (N_3004,N_2189,N_2007);
nor U3005 (N_3005,N_2712,N_2835);
and U3006 (N_3006,N_2217,N_2299);
and U3007 (N_3007,N_2055,N_2720);
or U3008 (N_3008,N_2404,N_2454);
xor U3009 (N_3009,N_2537,N_2039);
nand U3010 (N_3010,N_2030,N_2347);
xnor U3011 (N_3011,N_2427,N_2453);
xnor U3012 (N_3012,N_2115,N_2208);
and U3013 (N_3013,N_2624,N_2657);
and U3014 (N_3014,N_2412,N_2701);
xnor U3015 (N_3015,N_2672,N_2261);
nor U3016 (N_3016,N_2795,N_2787);
and U3017 (N_3017,N_2557,N_2178);
nor U3018 (N_3018,N_2942,N_2829);
nand U3019 (N_3019,N_2480,N_2113);
xor U3020 (N_3020,N_2108,N_2279);
nor U3021 (N_3021,N_2839,N_2020);
and U3022 (N_3022,N_2877,N_2396);
or U3023 (N_3023,N_2563,N_2500);
and U3024 (N_3024,N_2226,N_2072);
nor U3025 (N_3025,N_2604,N_2650);
xor U3026 (N_3026,N_2005,N_2886);
or U3027 (N_3027,N_2647,N_2070);
xor U3028 (N_3028,N_2848,N_2861);
or U3029 (N_3029,N_2060,N_2222);
or U3030 (N_3030,N_2174,N_2661);
nand U3031 (N_3031,N_2048,N_2369);
xnor U3032 (N_3032,N_2096,N_2056);
or U3033 (N_3033,N_2742,N_2838);
or U3034 (N_3034,N_2564,N_2365);
or U3035 (N_3035,N_2808,N_2802);
nor U3036 (N_3036,N_2988,N_2502);
and U3037 (N_3037,N_2989,N_2159);
or U3038 (N_3038,N_2263,N_2560);
nand U3039 (N_3039,N_2639,N_2403);
and U3040 (N_3040,N_2739,N_2152);
or U3041 (N_3041,N_2721,N_2642);
and U3042 (N_3042,N_2418,N_2387);
nand U3043 (N_3043,N_2840,N_2129);
nor U3044 (N_3044,N_2173,N_2817);
or U3045 (N_3045,N_2291,N_2874);
nor U3046 (N_3046,N_2180,N_2466);
nand U3047 (N_3047,N_2170,N_2197);
and U3048 (N_3048,N_2059,N_2755);
or U3049 (N_3049,N_2089,N_2851);
xor U3050 (N_3050,N_2336,N_2933);
and U3051 (N_3051,N_2338,N_2087);
and U3052 (N_3052,N_2846,N_2553);
xnor U3053 (N_3053,N_2111,N_2099);
or U3054 (N_3054,N_2779,N_2716);
or U3055 (N_3055,N_2765,N_2429);
nand U3056 (N_3056,N_2295,N_2531);
nor U3057 (N_3057,N_2085,N_2756);
xnor U3058 (N_3058,N_2797,N_2457);
or U3059 (N_3059,N_2745,N_2962);
or U3060 (N_3060,N_2930,N_2456);
or U3061 (N_3061,N_2319,N_2920);
or U3062 (N_3062,N_2722,N_2691);
xor U3063 (N_3063,N_2743,N_2616);
and U3064 (N_3064,N_2138,N_2488);
and U3065 (N_3065,N_2330,N_2784);
nand U3066 (N_3066,N_2011,N_2006);
and U3067 (N_3067,N_2306,N_2651);
xor U3068 (N_3068,N_2442,N_2836);
nor U3069 (N_3069,N_2938,N_2850);
nand U3070 (N_3070,N_2866,N_2535);
nor U3071 (N_3071,N_2934,N_2818);
nand U3072 (N_3072,N_2798,N_2694);
nor U3073 (N_3073,N_2735,N_2061);
and U3074 (N_3074,N_2340,N_2555);
and U3075 (N_3075,N_2234,N_2097);
nand U3076 (N_3076,N_2621,N_2094);
xnor U3077 (N_3077,N_2957,N_2758);
and U3078 (N_3078,N_2332,N_2872);
nor U3079 (N_3079,N_2757,N_2827);
nor U3080 (N_3080,N_2092,N_2337);
nand U3081 (N_3081,N_2717,N_2357);
nand U3082 (N_3082,N_2034,N_2978);
or U3083 (N_3083,N_2820,N_2154);
nor U3084 (N_3084,N_2885,N_2390);
or U3085 (N_3085,N_2550,N_2235);
and U3086 (N_3086,N_2546,N_2090);
nand U3087 (N_3087,N_2402,N_2467);
nor U3088 (N_3088,N_2576,N_2750);
xor U3089 (N_3089,N_2462,N_2527);
or U3090 (N_3090,N_2508,N_2358);
nor U3091 (N_3091,N_2073,N_2852);
nand U3092 (N_3092,N_2037,N_2669);
and U3093 (N_3093,N_2899,N_2249);
and U3094 (N_3094,N_2510,N_2380);
and U3095 (N_3095,N_2495,N_2698);
nor U3096 (N_3096,N_2038,N_2163);
and U3097 (N_3097,N_2386,N_2952);
and U3098 (N_3098,N_2186,N_2881);
nand U3099 (N_3099,N_2477,N_2479);
nand U3100 (N_3100,N_2329,N_2443);
nand U3101 (N_3101,N_2395,N_2935);
xnor U3102 (N_3102,N_2754,N_2972);
nor U3103 (N_3103,N_2946,N_2278);
nand U3104 (N_3104,N_2351,N_2548);
and U3105 (N_3105,N_2282,N_2752);
or U3106 (N_3106,N_2903,N_2663);
nand U3107 (N_3107,N_2632,N_2021);
xor U3108 (N_3108,N_2534,N_2385);
nand U3109 (N_3109,N_2890,N_2507);
nor U3110 (N_3110,N_2803,N_2376);
or U3111 (N_3111,N_2476,N_2411);
or U3112 (N_3112,N_2091,N_2924);
nand U3113 (N_3113,N_2825,N_2211);
or U3114 (N_3114,N_2882,N_2216);
nand U3115 (N_3115,N_2328,N_2871);
xnor U3116 (N_3116,N_2878,N_2305);
and U3117 (N_3117,N_2298,N_2789);
nor U3118 (N_3118,N_2455,N_2210);
xnor U3119 (N_3119,N_2645,N_2100);
or U3120 (N_3120,N_2079,N_2744);
nor U3121 (N_3121,N_2228,N_2759);
and U3122 (N_3122,N_2285,N_2318);
and U3123 (N_3123,N_2796,N_2486);
xor U3124 (N_3124,N_2425,N_2312);
xnor U3125 (N_3125,N_2517,N_2909);
or U3126 (N_3126,N_2383,N_2451);
nor U3127 (N_3127,N_2071,N_2204);
xnor U3128 (N_3128,N_2589,N_2855);
nor U3129 (N_3129,N_2074,N_2146);
and U3130 (N_3130,N_2421,N_2348);
xor U3131 (N_3131,N_2937,N_2002);
nand U3132 (N_3132,N_2482,N_2736);
or U3133 (N_3133,N_2671,N_2975);
and U3134 (N_3134,N_2018,N_2522);
or U3135 (N_3135,N_2898,N_2280);
or U3136 (N_3136,N_2928,N_2891);
nand U3137 (N_3137,N_2794,N_2469);
or U3138 (N_3138,N_2939,N_2856);
nand U3139 (N_3139,N_2049,N_2696);
nand U3140 (N_3140,N_2243,N_2088);
or U3141 (N_3141,N_2252,N_2927);
nor U3142 (N_3142,N_2292,N_2136);
and U3143 (N_3143,N_2904,N_2106);
nand U3144 (N_3144,N_2496,N_2580);
or U3145 (N_3145,N_2405,N_2976);
and U3146 (N_3146,N_2157,N_2653);
nand U3147 (N_3147,N_2008,N_2951);
or U3148 (N_3148,N_2300,N_2044);
or U3149 (N_3149,N_2579,N_2352);
nor U3150 (N_3150,N_2419,N_2431);
or U3151 (N_3151,N_2370,N_2791);
nand U3152 (N_3152,N_2414,N_2017);
xnor U3153 (N_3153,N_2459,N_2738);
nand U3154 (N_3154,N_2491,N_2257);
xnor U3155 (N_3155,N_2926,N_2889);
or U3156 (N_3156,N_2125,N_2967);
xor U3157 (N_3157,N_2316,N_2413);
xor U3158 (N_3158,N_2741,N_2317);
xnor U3159 (N_3159,N_2854,N_2296);
or U3160 (N_3160,N_2268,N_2999);
nand U3161 (N_3161,N_2905,N_2948);
or U3162 (N_3162,N_2936,N_2198);
or U3163 (N_3163,N_2849,N_2618);
nor U3164 (N_3164,N_2516,N_2705);
nand U3165 (N_3165,N_2104,N_2169);
nor U3166 (N_3166,N_2193,N_2110);
xnor U3167 (N_3167,N_2659,N_2001);
or U3168 (N_3168,N_2182,N_2232);
nor U3169 (N_3169,N_2654,N_2445);
and U3170 (N_3170,N_2212,N_2192);
xor U3171 (N_3171,N_2121,N_2393);
nor U3172 (N_3172,N_2966,N_2473);
and U3173 (N_3173,N_2792,N_2906);
or U3174 (N_3174,N_2984,N_2233);
and U3175 (N_3175,N_2655,N_2600);
nand U3176 (N_3176,N_2475,N_2066);
or U3177 (N_3177,N_2202,N_2956);
and U3178 (N_3178,N_2410,N_2275);
or U3179 (N_3179,N_2897,N_2595);
nor U3180 (N_3180,N_2023,N_2266);
or U3181 (N_3181,N_2324,N_2350);
nand U3182 (N_3182,N_2753,N_2126);
and U3183 (N_3183,N_2723,N_2747);
xor U3184 (N_3184,N_2623,N_2371);
nor U3185 (N_3185,N_2139,N_2588);
nor U3186 (N_3186,N_2912,N_2969);
or U3187 (N_3187,N_2730,N_2031);
or U3188 (N_3188,N_2276,N_2824);
nand U3189 (N_3189,N_2697,N_2987);
xor U3190 (N_3190,N_2360,N_2195);
and U3191 (N_3191,N_2775,N_2944);
and U3192 (N_3192,N_2605,N_2540);
nor U3193 (N_3193,N_2494,N_2441);
nand U3194 (N_3194,N_2870,N_2888);
or U3195 (N_3195,N_2346,N_2177);
nor U3196 (N_3196,N_2913,N_2172);
nand U3197 (N_3197,N_2492,N_2424);
nor U3198 (N_3198,N_2433,N_2029);
nor U3199 (N_3199,N_2707,N_2501);
nand U3200 (N_3200,N_2963,N_2751);
xor U3201 (N_3201,N_2270,N_2949);
nand U3202 (N_3202,N_2961,N_2361);
and U3203 (N_3203,N_2950,N_2238);
nor U3204 (N_3204,N_2185,N_2215);
or U3205 (N_3205,N_2065,N_2526);
nor U3206 (N_3206,N_2613,N_2719);
and U3207 (N_3207,N_2118,N_2602);
or U3208 (N_3208,N_2625,N_2641);
xor U3209 (N_3209,N_2101,N_2313);
or U3210 (N_3210,N_2041,N_2907);
or U3211 (N_3211,N_2541,N_2043);
nor U3212 (N_3212,N_2581,N_2981);
or U3213 (N_3213,N_2286,N_2117);
or U3214 (N_3214,N_2098,N_2505);
nand U3215 (N_3215,N_2807,N_2678);
or U3216 (N_3216,N_2985,N_2628);
nand U3217 (N_3217,N_2627,N_2648);
nand U3218 (N_3218,N_2472,N_2076);
nand U3219 (N_3219,N_2590,N_2155);
nand U3220 (N_3220,N_2816,N_2593);
or U3221 (N_3221,N_2223,N_2200);
or U3222 (N_3222,N_2919,N_2958);
nand U3223 (N_3223,N_2801,N_2067);
nand U3224 (N_3224,N_2964,N_2847);
and U3225 (N_3225,N_2686,N_2584);
xnor U3226 (N_3226,N_2863,N_2788);
and U3227 (N_3227,N_2069,N_2040);
and U3228 (N_3228,N_2970,N_2761);
and U3229 (N_3229,N_2301,N_2144);
nor U3230 (N_3230,N_2635,N_2248);
nor U3231 (N_3231,N_2677,N_2996);
nand U3232 (N_3232,N_2504,N_2033);
xor U3233 (N_3233,N_2973,N_2833);
nand U3234 (N_3234,N_2068,N_2407);
nor U3235 (N_3235,N_2596,N_2575);
or U3236 (N_3236,N_2325,N_2729);
xor U3237 (N_3237,N_2607,N_2731);
nand U3238 (N_3238,N_2025,N_2503);
xor U3239 (N_3239,N_2811,N_2810);
xor U3240 (N_3240,N_2690,N_2046);
or U3241 (N_3241,N_2687,N_2470);
xor U3242 (N_3242,N_2941,N_2237);
or U3243 (N_3243,N_2762,N_2760);
nand U3244 (N_3244,N_2241,N_2815);
or U3245 (N_3245,N_2323,N_2577);
and U3246 (N_3246,N_2790,N_2116);
xor U3247 (N_3247,N_2458,N_2450);
or U3248 (N_3248,N_2992,N_2225);
xnor U3249 (N_3249,N_2271,N_2288);
nor U3250 (N_3250,N_2239,N_2597);
nand U3251 (N_3251,N_2436,N_2895);
nand U3252 (N_3252,N_2868,N_2434);
xnor U3253 (N_3253,N_2734,N_2284);
nor U3254 (N_3254,N_2213,N_2900);
nor U3255 (N_3255,N_2084,N_2539);
and U3256 (N_3256,N_2599,N_2132);
xor U3257 (N_3257,N_2063,N_2683);
nand U3258 (N_3258,N_2181,N_2670);
nor U3259 (N_3259,N_2626,N_2649);
or U3260 (N_3260,N_2554,N_2016);
and U3261 (N_3261,N_2047,N_2865);
xnor U3262 (N_3262,N_2447,N_2191);
xor U3263 (N_3263,N_2461,N_2205);
or U3264 (N_3264,N_2499,N_2314);
nand U3265 (N_3265,N_2460,N_2585);
or U3266 (N_3266,N_2977,N_2766);
nor U3267 (N_3267,N_2594,N_2528);
and U3268 (N_3268,N_2331,N_2381);
xor U3269 (N_3269,N_2269,N_2994);
xnor U3270 (N_3270,N_2947,N_2574);
nor U3271 (N_3271,N_2013,N_2769);
or U3272 (N_3272,N_2864,N_2609);
or U3273 (N_3273,N_2774,N_2706);
xor U3274 (N_3274,N_2297,N_2971);
nand U3275 (N_3275,N_2448,N_2051);
xor U3276 (N_3276,N_2902,N_2354);
xnor U3277 (N_3277,N_2026,N_2859);
nand U3278 (N_3278,N_2610,N_2032);
xor U3279 (N_3279,N_2179,N_2326);
nand U3280 (N_3280,N_2133,N_2437);
or U3281 (N_3281,N_2583,N_2770);
and U3282 (N_3282,N_2119,N_2399);
nand U3283 (N_3283,N_2397,N_2559);
or U3284 (N_3284,N_2161,N_2151);
xor U3285 (N_3285,N_2733,N_2053);
and U3286 (N_3286,N_2258,N_2800);
or U3287 (N_3287,N_2438,N_2781);
nor U3288 (N_3288,N_2538,N_2289);
and U3289 (N_3289,N_2805,N_2343);
nor U3290 (N_3290,N_2551,N_2165);
xor U3291 (N_3291,N_2320,N_2614);
nand U3292 (N_3292,N_2294,N_2979);
xnor U3293 (N_3293,N_2545,N_2832);
xnor U3294 (N_3294,N_2416,N_2915);
nand U3295 (N_3295,N_2841,N_2601);
and U3296 (N_3296,N_2876,N_2571);
and U3297 (N_3297,N_2322,N_2175);
or U3298 (N_3298,N_2603,N_2484);
and U3299 (N_3299,N_2862,N_2558);
and U3300 (N_3300,N_2303,N_2509);
xnor U3301 (N_3301,N_2114,N_2130);
nand U3302 (N_3302,N_2965,N_2812);
or U3303 (N_3303,N_2024,N_2831);
xor U3304 (N_3304,N_2894,N_2004);
or U3305 (N_3305,N_2804,N_2646);
or U3306 (N_3306,N_2245,N_2513);
nand U3307 (N_3307,N_2464,N_2171);
nand U3308 (N_3308,N_2783,N_2452);
nand U3309 (N_3309,N_2218,N_2879);
or U3310 (N_3310,N_2821,N_2974);
or U3311 (N_3311,N_2281,N_2489);
or U3312 (N_3312,N_2887,N_2630);
and U3313 (N_3313,N_2107,N_2633);
or U3314 (N_3314,N_2901,N_2867);
or U3315 (N_3315,N_2598,N_2262);
and U3316 (N_3316,N_2362,N_2699);
nand U3317 (N_3317,N_2556,N_2240);
or U3318 (N_3318,N_2893,N_2439);
xor U3319 (N_3319,N_2015,N_2483);
nor U3320 (N_3320,N_2112,N_2570);
nor U3321 (N_3321,N_2430,N_2689);
or U3322 (N_3322,N_2035,N_2644);
or U3323 (N_3323,N_2378,N_2667);
or U3324 (N_3324,N_2382,N_2264);
nor U3325 (N_3325,N_2565,N_2700);
and U3326 (N_3326,N_2188,N_2374);
and U3327 (N_3327,N_2080,N_2547);
nor U3328 (N_3328,N_2704,N_2529);
xnor U3329 (N_3329,N_2147,N_2656);
nor U3330 (N_3330,N_2010,N_2674);
xor U3331 (N_3331,N_2711,N_2207);
xnor U3332 (N_3332,N_2620,N_2446);
and U3333 (N_3333,N_2168,N_2377);
nand U3334 (N_3334,N_2149,N_2858);
xnor U3335 (N_3335,N_2520,N_2493);
xor U3336 (N_3336,N_2081,N_2162);
nand U3337 (N_3337,N_2426,N_2142);
nand U3338 (N_3338,N_2995,N_2637);
xor U3339 (N_3339,N_2629,N_2845);
nand U3340 (N_3340,N_2183,N_2355);
nor U3341 (N_3341,N_2022,N_2150);
or U3342 (N_3342,N_2883,N_2219);
nand U3343 (N_3343,N_2478,N_2267);
or U3344 (N_3344,N_2660,N_2229);
nor U3345 (N_3345,N_2379,N_2463);
or U3346 (N_3346,N_2423,N_2375);
xor U3347 (N_3347,N_2260,N_2843);
xnor U3348 (N_3348,N_2542,N_2544);
or U3349 (N_3349,N_2943,N_2400);
nor U3350 (N_3350,N_2998,N_2619);
nor U3351 (N_3351,N_2283,N_2444);
nor U3352 (N_3352,N_2572,N_2945);
or U3353 (N_3353,N_2873,N_2519);
nand U3354 (N_3354,N_2591,N_2842);
and U3355 (N_3355,N_2880,N_2631);
or U3356 (N_3356,N_2675,N_2058);
nand U3357 (N_3357,N_2922,N_2702);
and U3358 (N_3358,N_2954,N_2201);
and U3359 (N_3359,N_2036,N_2586);
or U3360 (N_3360,N_2715,N_2156);
nor U3361 (N_3361,N_2658,N_2481);
and U3362 (N_3362,N_2506,N_2875);
and U3363 (N_3363,N_2986,N_2401);
or U3364 (N_3364,N_2515,N_2908);
and U3365 (N_3365,N_2339,N_2256);
or U3366 (N_3366,N_2310,N_2932);
nand U3367 (N_3367,N_2042,N_2834);
nor U3368 (N_3368,N_2290,N_2725);
nand U3369 (N_3369,N_2124,N_2911);
xnor U3370 (N_3370,N_2344,N_2273);
or U3371 (N_3371,N_2959,N_2814);
nor U3372 (N_3372,N_2737,N_2160);
xor U3373 (N_3373,N_2676,N_2167);
xor U3374 (N_3374,N_2786,N_2221);
xnor U3375 (N_3375,N_2732,N_2131);
nand U3376 (N_3376,N_2617,N_2771);
xnor U3377 (N_3377,N_2384,N_2103);
or U3378 (N_3378,N_2608,N_2251);
nor U3379 (N_3379,N_2776,N_2611);
nand U3380 (N_3380,N_2334,N_2014);
nor U3381 (N_3381,N_2896,N_2763);
xor U3382 (N_3382,N_2767,N_2826);
or U3383 (N_3383,N_2468,N_2184);
and U3384 (N_3384,N_2123,N_2077);
or U3385 (N_3385,N_2844,N_2253);
nand U3386 (N_3386,N_2000,N_2465);
nand U3387 (N_3387,N_2860,N_2740);
nor U3388 (N_3388,N_2993,N_2302);
nand U3389 (N_3389,N_2749,N_2511);
xnor U3390 (N_3390,N_2746,N_2127);
nand U3391 (N_3391,N_2363,N_2809);
and U3392 (N_3392,N_2220,N_2518);
or U3393 (N_3393,N_2960,N_2695);
and U3394 (N_3394,N_2471,N_2359);
and U3395 (N_3395,N_2709,N_2164);
xnor U3396 (N_3396,N_2140,N_2692);
xor U3397 (N_3397,N_2837,N_2345);
nor U3398 (N_3398,N_2086,N_2892);
nand U3399 (N_3399,N_2388,N_2636);
nand U3400 (N_3400,N_2668,N_2166);
and U3401 (N_3401,N_2569,N_2512);
nand U3402 (N_3402,N_2304,N_2277);
or U3403 (N_3403,N_2724,N_2778);
or U3404 (N_3404,N_2128,N_2095);
and U3405 (N_3405,N_2490,N_2533);
and U3406 (N_3406,N_2366,N_2869);
nand U3407 (N_3407,N_2003,N_2931);
and U3408 (N_3408,N_2684,N_2428);
nand U3409 (N_3409,N_2105,N_2525);
nor U3410 (N_3410,N_2640,N_2940);
xor U3411 (N_3411,N_2398,N_2622);
or U3412 (N_3412,N_2703,N_2780);
and U3413 (N_3413,N_2524,N_2187);
and U3414 (N_3414,N_2373,N_2308);
nand U3415 (N_3415,N_2914,N_2806);
nand U3416 (N_3416,N_2272,N_2372);
nand U3417 (N_3417,N_2082,N_2307);
nand U3418 (N_3418,N_2255,N_2209);
xor U3419 (N_3419,N_2773,N_2009);
nand U3420 (N_3420,N_2349,N_2714);
nor U3421 (N_3421,N_2415,N_2982);
or U3422 (N_3422,N_2828,N_2536);
xnor U3423 (N_3423,N_2148,N_2335);
and U3424 (N_3424,N_2242,N_2497);
nor U3425 (N_3425,N_2199,N_2389);
and U3426 (N_3426,N_2634,N_2681);
or U3427 (N_3427,N_2688,N_2214);
nand U3428 (N_3428,N_2592,N_2799);
or U3429 (N_3429,N_2135,N_2728);
and U3430 (N_3430,N_2028,N_2748);
nor U3431 (N_3431,N_2045,N_2368);
or U3432 (N_3432,N_2582,N_2293);
or U3433 (N_3433,N_2666,N_2230);
xor U3434 (N_3434,N_2109,N_2777);
or U3435 (N_3435,N_2772,N_2680);
nor U3436 (N_3436,N_2054,N_2679);
or U3437 (N_3437,N_2673,N_2568);
or U3438 (N_3438,N_2853,N_2356);
nor U3439 (N_3439,N_2693,N_2078);
nand U3440 (N_3440,N_2997,N_2064);
xor U3441 (N_3441,N_2980,N_2485);
nor U3442 (N_3442,N_2190,N_2196);
xnor U3443 (N_3443,N_2929,N_2785);
xor U3444 (N_3444,N_2923,N_2578);
xnor U3445 (N_3445,N_2925,N_2417);
xor U3446 (N_3446,N_2857,N_2265);
nor U3447 (N_3447,N_2768,N_2246);
or U3448 (N_3448,N_2206,N_2953);
or U3449 (N_3449,N_2141,N_2521);
and U3450 (N_3450,N_2440,N_2093);
nor U3451 (N_3451,N_2983,N_2057);
nand U3452 (N_3452,N_2523,N_2822);
and U3453 (N_3453,N_2236,N_2227);
nand U3454 (N_3454,N_2552,N_2587);
and U3455 (N_3455,N_2342,N_2514);
nor U3456 (N_3456,N_2259,N_2573);
or U3457 (N_3457,N_2408,N_2321);
and U3458 (N_3458,N_2449,N_2250);
nor U3459 (N_3459,N_2561,N_2664);
nor U3460 (N_3460,N_2685,N_2143);
nand U3461 (N_3461,N_2327,N_2422);
nor U3462 (N_3462,N_2819,N_2782);
and U3463 (N_3463,N_2062,N_2391);
xnor U3464 (N_3464,N_2830,N_2341);
and U3465 (N_3465,N_2247,N_2194);
nand U3466 (N_3466,N_2019,N_2176);
xor U3467 (N_3467,N_2432,N_2394);
nand U3468 (N_3468,N_2120,N_2367);
xor U3469 (N_3469,N_2921,N_2083);
and U3470 (N_3470,N_2333,N_2665);
and U3471 (N_3471,N_2075,N_2287);
nor U3472 (N_3472,N_2409,N_2392);
xnor U3473 (N_3473,N_2918,N_2713);
and U3474 (N_3474,N_2052,N_2615);
nand U3475 (N_3475,N_2364,N_2244);
and U3476 (N_3476,N_2612,N_2662);
and U3477 (N_3477,N_2530,N_2153);
xnor U3478 (N_3478,N_2638,N_2567);
nor U3479 (N_3479,N_2309,N_2990);
or U3480 (N_3480,N_2122,N_2562);
nand U3481 (N_3481,N_2487,N_2353);
or U3482 (N_3482,N_2727,N_2726);
nand U3483 (N_3483,N_2420,N_2027);
xnor U3484 (N_3484,N_2231,N_2137);
nor U3485 (N_3485,N_2718,N_2917);
xnor U3486 (N_3486,N_2145,N_2050);
or U3487 (N_3487,N_2710,N_2916);
nand U3488 (N_3488,N_2474,N_2435);
or U3489 (N_3489,N_2254,N_2406);
or U3490 (N_3490,N_2884,N_2823);
xnor U3491 (N_3491,N_2813,N_2012);
and U3492 (N_3492,N_2643,N_2968);
or U3493 (N_3493,N_2158,N_2606);
xnor U3494 (N_3494,N_2708,N_2652);
nand U3495 (N_3495,N_2991,N_2498);
and U3496 (N_3496,N_2532,N_2274);
xor U3497 (N_3497,N_2134,N_2311);
xor U3498 (N_3498,N_2224,N_2764);
nand U3499 (N_3499,N_2566,N_2203);
nor U3500 (N_3500,N_2162,N_2675);
or U3501 (N_3501,N_2237,N_2520);
or U3502 (N_3502,N_2546,N_2403);
or U3503 (N_3503,N_2227,N_2842);
or U3504 (N_3504,N_2564,N_2161);
nor U3505 (N_3505,N_2772,N_2417);
or U3506 (N_3506,N_2656,N_2348);
nor U3507 (N_3507,N_2994,N_2405);
xnor U3508 (N_3508,N_2652,N_2575);
and U3509 (N_3509,N_2825,N_2262);
nor U3510 (N_3510,N_2419,N_2557);
nand U3511 (N_3511,N_2750,N_2474);
xor U3512 (N_3512,N_2734,N_2419);
nand U3513 (N_3513,N_2924,N_2463);
xor U3514 (N_3514,N_2227,N_2047);
nand U3515 (N_3515,N_2119,N_2240);
and U3516 (N_3516,N_2612,N_2927);
or U3517 (N_3517,N_2319,N_2033);
xor U3518 (N_3518,N_2378,N_2213);
xor U3519 (N_3519,N_2718,N_2312);
and U3520 (N_3520,N_2770,N_2552);
xnor U3521 (N_3521,N_2314,N_2483);
or U3522 (N_3522,N_2271,N_2981);
and U3523 (N_3523,N_2850,N_2039);
nor U3524 (N_3524,N_2888,N_2566);
nor U3525 (N_3525,N_2351,N_2236);
xor U3526 (N_3526,N_2226,N_2786);
or U3527 (N_3527,N_2473,N_2203);
nand U3528 (N_3528,N_2146,N_2708);
nand U3529 (N_3529,N_2657,N_2460);
or U3530 (N_3530,N_2792,N_2969);
nor U3531 (N_3531,N_2381,N_2275);
nor U3532 (N_3532,N_2802,N_2939);
xor U3533 (N_3533,N_2911,N_2705);
nand U3534 (N_3534,N_2675,N_2135);
nand U3535 (N_3535,N_2829,N_2187);
nor U3536 (N_3536,N_2417,N_2660);
nor U3537 (N_3537,N_2986,N_2588);
nand U3538 (N_3538,N_2468,N_2661);
nand U3539 (N_3539,N_2483,N_2808);
nand U3540 (N_3540,N_2137,N_2394);
xor U3541 (N_3541,N_2006,N_2567);
or U3542 (N_3542,N_2013,N_2800);
nand U3543 (N_3543,N_2547,N_2062);
and U3544 (N_3544,N_2522,N_2628);
nand U3545 (N_3545,N_2032,N_2359);
nor U3546 (N_3546,N_2287,N_2383);
xor U3547 (N_3547,N_2559,N_2540);
nand U3548 (N_3548,N_2441,N_2553);
xor U3549 (N_3549,N_2186,N_2629);
nand U3550 (N_3550,N_2198,N_2956);
nor U3551 (N_3551,N_2094,N_2865);
nor U3552 (N_3552,N_2871,N_2750);
and U3553 (N_3553,N_2524,N_2395);
nor U3554 (N_3554,N_2846,N_2076);
nor U3555 (N_3555,N_2729,N_2756);
and U3556 (N_3556,N_2715,N_2450);
or U3557 (N_3557,N_2714,N_2441);
or U3558 (N_3558,N_2418,N_2355);
or U3559 (N_3559,N_2048,N_2532);
xor U3560 (N_3560,N_2417,N_2654);
xor U3561 (N_3561,N_2264,N_2763);
and U3562 (N_3562,N_2598,N_2053);
nand U3563 (N_3563,N_2683,N_2527);
nor U3564 (N_3564,N_2693,N_2882);
or U3565 (N_3565,N_2540,N_2657);
and U3566 (N_3566,N_2515,N_2767);
xor U3567 (N_3567,N_2059,N_2313);
nand U3568 (N_3568,N_2638,N_2129);
nor U3569 (N_3569,N_2967,N_2098);
xor U3570 (N_3570,N_2751,N_2004);
xnor U3571 (N_3571,N_2035,N_2804);
nand U3572 (N_3572,N_2109,N_2334);
nor U3573 (N_3573,N_2423,N_2991);
and U3574 (N_3574,N_2574,N_2996);
or U3575 (N_3575,N_2987,N_2436);
nand U3576 (N_3576,N_2307,N_2169);
and U3577 (N_3577,N_2565,N_2018);
or U3578 (N_3578,N_2605,N_2927);
nor U3579 (N_3579,N_2325,N_2631);
and U3580 (N_3580,N_2353,N_2169);
or U3581 (N_3581,N_2151,N_2172);
and U3582 (N_3582,N_2927,N_2892);
or U3583 (N_3583,N_2278,N_2307);
nor U3584 (N_3584,N_2652,N_2924);
xor U3585 (N_3585,N_2765,N_2506);
or U3586 (N_3586,N_2640,N_2855);
nand U3587 (N_3587,N_2739,N_2628);
or U3588 (N_3588,N_2128,N_2944);
or U3589 (N_3589,N_2963,N_2628);
and U3590 (N_3590,N_2223,N_2650);
nor U3591 (N_3591,N_2785,N_2402);
nor U3592 (N_3592,N_2757,N_2164);
nand U3593 (N_3593,N_2514,N_2496);
or U3594 (N_3594,N_2448,N_2694);
nor U3595 (N_3595,N_2465,N_2816);
or U3596 (N_3596,N_2642,N_2578);
nand U3597 (N_3597,N_2337,N_2799);
or U3598 (N_3598,N_2436,N_2759);
nor U3599 (N_3599,N_2229,N_2173);
xor U3600 (N_3600,N_2330,N_2502);
and U3601 (N_3601,N_2048,N_2505);
nand U3602 (N_3602,N_2528,N_2852);
nand U3603 (N_3603,N_2062,N_2879);
and U3604 (N_3604,N_2713,N_2855);
or U3605 (N_3605,N_2264,N_2894);
nor U3606 (N_3606,N_2608,N_2950);
and U3607 (N_3607,N_2064,N_2153);
and U3608 (N_3608,N_2679,N_2959);
and U3609 (N_3609,N_2940,N_2698);
and U3610 (N_3610,N_2448,N_2715);
nor U3611 (N_3611,N_2637,N_2962);
nand U3612 (N_3612,N_2892,N_2279);
xnor U3613 (N_3613,N_2049,N_2369);
nor U3614 (N_3614,N_2346,N_2250);
nand U3615 (N_3615,N_2006,N_2273);
or U3616 (N_3616,N_2512,N_2685);
nand U3617 (N_3617,N_2829,N_2278);
nand U3618 (N_3618,N_2301,N_2217);
and U3619 (N_3619,N_2783,N_2719);
or U3620 (N_3620,N_2050,N_2265);
nand U3621 (N_3621,N_2830,N_2127);
or U3622 (N_3622,N_2835,N_2608);
nor U3623 (N_3623,N_2538,N_2412);
and U3624 (N_3624,N_2109,N_2363);
nor U3625 (N_3625,N_2217,N_2701);
or U3626 (N_3626,N_2256,N_2472);
xor U3627 (N_3627,N_2680,N_2279);
nand U3628 (N_3628,N_2111,N_2477);
or U3629 (N_3629,N_2495,N_2201);
or U3630 (N_3630,N_2957,N_2988);
nand U3631 (N_3631,N_2417,N_2875);
xor U3632 (N_3632,N_2910,N_2601);
nand U3633 (N_3633,N_2019,N_2405);
nor U3634 (N_3634,N_2789,N_2739);
and U3635 (N_3635,N_2355,N_2945);
nor U3636 (N_3636,N_2005,N_2860);
or U3637 (N_3637,N_2478,N_2519);
xor U3638 (N_3638,N_2707,N_2062);
nand U3639 (N_3639,N_2577,N_2710);
nor U3640 (N_3640,N_2808,N_2327);
xor U3641 (N_3641,N_2004,N_2390);
xor U3642 (N_3642,N_2977,N_2489);
or U3643 (N_3643,N_2273,N_2883);
nand U3644 (N_3644,N_2047,N_2099);
xnor U3645 (N_3645,N_2886,N_2702);
and U3646 (N_3646,N_2919,N_2630);
or U3647 (N_3647,N_2642,N_2727);
or U3648 (N_3648,N_2804,N_2042);
or U3649 (N_3649,N_2006,N_2357);
xnor U3650 (N_3650,N_2947,N_2802);
or U3651 (N_3651,N_2731,N_2324);
nand U3652 (N_3652,N_2501,N_2077);
or U3653 (N_3653,N_2976,N_2641);
xnor U3654 (N_3654,N_2803,N_2074);
and U3655 (N_3655,N_2188,N_2078);
nand U3656 (N_3656,N_2554,N_2333);
or U3657 (N_3657,N_2432,N_2425);
nor U3658 (N_3658,N_2366,N_2488);
and U3659 (N_3659,N_2553,N_2690);
nor U3660 (N_3660,N_2514,N_2040);
or U3661 (N_3661,N_2030,N_2965);
nand U3662 (N_3662,N_2779,N_2998);
or U3663 (N_3663,N_2071,N_2496);
nor U3664 (N_3664,N_2407,N_2492);
or U3665 (N_3665,N_2880,N_2070);
or U3666 (N_3666,N_2602,N_2838);
or U3667 (N_3667,N_2335,N_2446);
or U3668 (N_3668,N_2074,N_2229);
nand U3669 (N_3669,N_2633,N_2636);
xnor U3670 (N_3670,N_2810,N_2404);
and U3671 (N_3671,N_2970,N_2650);
nor U3672 (N_3672,N_2523,N_2498);
nor U3673 (N_3673,N_2973,N_2381);
and U3674 (N_3674,N_2688,N_2554);
or U3675 (N_3675,N_2332,N_2681);
and U3676 (N_3676,N_2932,N_2652);
xnor U3677 (N_3677,N_2497,N_2673);
nor U3678 (N_3678,N_2263,N_2666);
xnor U3679 (N_3679,N_2466,N_2646);
xor U3680 (N_3680,N_2972,N_2560);
xor U3681 (N_3681,N_2229,N_2352);
nor U3682 (N_3682,N_2466,N_2047);
and U3683 (N_3683,N_2532,N_2466);
xnor U3684 (N_3684,N_2614,N_2301);
or U3685 (N_3685,N_2992,N_2901);
xnor U3686 (N_3686,N_2932,N_2386);
or U3687 (N_3687,N_2400,N_2505);
nor U3688 (N_3688,N_2454,N_2262);
xnor U3689 (N_3689,N_2755,N_2570);
nor U3690 (N_3690,N_2732,N_2915);
nand U3691 (N_3691,N_2499,N_2815);
nor U3692 (N_3692,N_2883,N_2041);
xnor U3693 (N_3693,N_2571,N_2168);
nand U3694 (N_3694,N_2053,N_2990);
nand U3695 (N_3695,N_2493,N_2042);
nand U3696 (N_3696,N_2384,N_2062);
nand U3697 (N_3697,N_2596,N_2426);
xnor U3698 (N_3698,N_2505,N_2580);
or U3699 (N_3699,N_2708,N_2634);
or U3700 (N_3700,N_2724,N_2277);
xnor U3701 (N_3701,N_2345,N_2214);
and U3702 (N_3702,N_2875,N_2606);
and U3703 (N_3703,N_2860,N_2484);
nor U3704 (N_3704,N_2708,N_2315);
or U3705 (N_3705,N_2558,N_2049);
or U3706 (N_3706,N_2401,N_2831);
nor U3707 (N_3707,N_2905,N_2660);
and U3708 (N_3708,N_2356,N_2219);
or U3709 (N_3709,N_2795,N_2088);
xor U3710 (N_3710,N_2102,N_2436);
or U3711 (N_3711,N_2349,N_2509);
and U3712 (N_3712,N_2110,N_2202);
and U3713 (N_3713,N_2418,N_2419);
nand U3714 (N_3714,N_2135,N_2307);
and U3715 (N_3715,N_2769,N_2275);
nand U3716 (N_3716,N_2653,N_2785);
nor U3717 (N_3717,N_2703,N_2690);
and U3718 (N_3718,N_2054,N_2113);
nand U3719 (N_3719,N_2407,N_2874);
and U3720 (N_3720,N_2212,N_2716);
nand U3721 (N_3721,N_2354,N_2053);
or U3722 (N_3722,N_2973,N_2811);
nand U3723 (N_3723,N_2037,N_2184);
and U3724 (N_3724,N_2651,N_2134);
nand U3725 (N_3725,N_2976,N_2832);
xor U3726 (N_3726,N_2631,N_2516);
xnor U3727 (N_3727,N_2987,N_2579);
nor U3728 (N_3728,N_2373,N_2321);
or U3729 (N_3729,N_2080,N_2178);
or U3730 (N_3730,N_2849,N_2549);
xor U3731 (N_3731,N_2041,N_2186);
nor U3732 (N_3732,N_2301,N_2290);
or U3733 (N_3733,N_2353,N_2238);
xor U3734 (N_3734,N_2800,N_2844);
nand U3735 (N_3735,N_2253,N_2261);
or U3736 (N_3736,N_2947,N_2347);
nand U3737 (N_3737,N_2183,N_2877);
nor U3738 (N_3738,N_2805,N_2945);
xnor U3739 (N_3739,N_2077,N_2805);
or U3740 (N_3740,N_2308,N_2027);
nor U3741 (N_3741,N_2148,N_2889);
xor U3742 (N_3742,N_2249,N_2728);
nor U3743 (N_3743,N_2735,N_2956);
nand U3744 (N_3744,N_2621,N_2919);
xnor U3745 (N_3745,N_2967,N_2372);
and U3746 (N_3746,N_2745,N_2417);
xnor U3747 (N_3747,N_2579,N_2232);
nand U3748 (N_3748,N_2434,N_2917);
xor U3749 (N_3749,N_2638,N_2500);
and U3750 (N_3750,N_2143,N_2387);
nor U3751 (N_3751,N_2425,N_2294);
or U3752 (N_3752,N_2698,N_2934);
or U3753 (N_3753,N_2777,N_2675);
nor U3754 (N_3754,N_2257,N_2337);
nand U3755 (N_3755,N_2403,N_2854);
xor U3756 (N_3756,N_2568,N_2943);
or U3757 (N_3757,N_2284,N_2112);
nor U3758 (N_3758,N_2897,N_2778);
and U3759 (N_3759,N_2921,N_2500);
nor U3760 (N_3760,N_2865,N_2850);
xnor U3761 (N_3761,N_2759,N_2247);
nor U3762 (N_3762,N_2680,N_2342);
xnor U3763 (N_3763,N_2613,N_2036);
nor U3764 (N_3764,N_2860,N_2732);
nand U3765 (N_3765,N_2269,N_2816);
nand U3766 (N_3766,N_2088,N_2655);
nand U3767 (N_3767,N_2994,N_2808);
and U3768 (N_3768,N_2338,N_2531);
and U3769 (N_3769,N_2001,N_2973);
nand U3770 (N_3770,N_2031,N_2781);
nand U3771 (N_3771,N_2048,N_2045);
or U3772 (N_3772,N_2584,N_2740);
nor U3773 (N_3773,N_2815,N_2185);
or U3774 (N_3774,N_2551,N_2630);
nor U3775 (N_3775,N_2895,N_2380);
nor U3776 (N_3776,N_2695,N_2462);
xnor U3777 (N_3777,N_2287,N_2398);
or U3778 (N_3778,N_2353,N_2777);
xor U3779 (N_3779,N_2549,N_2730);
xnor U3780 (N_3780,N_2274,N_2570);
xor U3781 (N_3781,N_2125,N_2817);
nand U3782 (N_3782,N_2391,N_2603);
nand U3783 (N_3783,N_2348,N_2449);
nand U3784 (N_3784,N_2845,N_2460);
nor U3785 (N_3785,N_2349,N_2734);
nand U3786 (N_3786,N_2486,N_2733);
nor U3787 (N_3787,N_2592,N_2705);
and U3788 (N_3788,N_2725,N_2022);
nor U3789 (N_3789,N_2947,N_2378);
or U3790 (N_3790,N_2176,N_2123);
nand U3791 (N_3791,N_2479,N_2153);
xnor U3792 (N_3792,N_2921,N_2472);
xnor U3793 (N_3793,N_2244,N_2360);
and U3794 (N_3794,N_2680,N_2787);
and U3795 (N_3795,N_2174,N_2911);
xnor U3796 (N_3796,N_2112,N_2551);
and U3797 (N_3797,N_2544,N_2744);
and U3798 (N_3798,N_2268,N_2438);
nor U3799 (N_3799,N_2272,N_2484);
nor U3800 (N_3800,N_2774,N_2212);
or U3801 (N_3801,N_2401,N_2549);
nor U3802 (N_3802,N_2022,N_2676);
and U3803 (N_3803,N_2651,N_2026);
xnor U3804 (N_3804,N_2467,N_2279);
nand U3805 (N_3805,N_2016,N_2194);
nand U3806 (N_3806,N_2873,N_2734);
xor U3807 (N_3807,N_2262,N_2623);
xnor U3808 (N_3808,N_2066,N_2807);
and U3809 (N_3809,N_2455,N_2464);
and U3810 (N_3810,N_2076,N_2596);
and U3811 (N_3811,N_2501,N_2168);
or U3812 (N_3812,N_2338,N_2599);
or U3813 (N_3813,N_2818,N_2650);
and U3814 (N_3814,N_2526,N_2347);
and U3815 (N_3815,N_2376,N_2566);
and U3816 (N_3816,N_2994,N_2473);
or U3817 (N_3817,N_2718,N_2538);
nand U3818 (N_3818,N_2242,N_2991);
nor U3819 (N_3819,N_2301,N_2433);
xnor U3820 (N_3820,N_2482,N_2660);
xnor U3821 (N_3821,N_2322,N_2697);
xnor U3822 (N_3822,N_2148,N_2807);
nor U3823 (N_3823,N_2830,N_2501);
or U3824 (N_3824,N_2625,N_2823);
or U3825 (N_3825,N_2746,N_2727);
nor U3826 (N_3826,N_2754,N_2885);
nor U3827 (N_3827,N_2327,N_2223);
nand U3828 (N_3828,N_2724,N_2565);
nor U3829 (N_3829,N_2882,N_2685);
nand U3830 (N_3830,N_2384,N_2155);
nand U3831 (N_3831,N_2528,N_2985);
and U3832 (N_3832,N_2957,N_2230);
nor U3833 (N_3833,N_2825,N_2797);
nor U3834 (N_3834,N_2710,N_2944);
and U3835 (N_3835,N_2958,N_2262);
or U3836 (N_3836,N_2209,N_2626);
and U3837 (N_3837,N_2426,N_2831);
and U3838 (N_3838,N_2114,N_2836);
and U3839 (N_3839,N_2359,N_2962);
or U3840 (N_3840,N_2750,N_2443);
or U3841 (N_3841,N_2263,N_2138);
nor U3842 (N_3842,N_2706,N_2909);
xor U3843 (N_3843,N_2581,N_2508);
xnor U3844 (N_3844,N_2673,N_2897);
or U3845 (N_3845,N_2617,N_2364);
nor U3846 (N_3846,N_2849,N_2734);
xnor U3847 (N_3847,N_2977,N_2759);
nor U3848 (N_3848,N_2623,N_2400);
and U3849 (N_3849,N_2600,N_2204);
nand U3850 (N_3850,N_2114,N_2959);
and U3851 (N_3851,N_2547,N_2382);
xnor U3852 (N_3852,N_2636,N_2221);
and U3853 (N_3853,N_2829,N_2245);
or U3854 (N_3854,N_2439,N_2754);
or U3855 (N_3855,N_2644,N_2982);
xor U3856 (N_3856,N_2670,N_2723);
nand U3857 (N_3857,N_2017,N_2992);
xor U3858 (N_3858,N_2929,N_2008);
nor U3859 (N_3859,N_2973,N_2008);
and U3860 (N_3860,N_2050,N_2656);
nor U3861 (N_3861,N_2589,N_2162);
nor U3862 (N_3862,N_2294,N_2132);
xnor U3863 (N_3863,N_2851,N_2375);
nand U3864 (N_3864,N_2018,N_2117);
xor U3865 (N_3865,N_2352,N_2230);
nor U3866 (N_3866,N_2726,N_2360);
nor U3867 (N_3867,N_2879,N_2603);
nor U3868 (N_3868,N_2634,N_2169);
nor U3869 (N_3869,N_2706,N_2464);
nor U3870 (N_3870,N_2106,N_2861);
nand U3871 (N_3871,N_2904,N_2332);
nor U3872 (N_3872,N_2670,N_2679);
nor U3873 (N_3873,N_2408,N_2556);
or U3874 (N_3874,N_2432,N_2281);
and U3875 (N_3875,N_2744,N_2720);
and U3876 (N_3876,N_2257,N_2648);
or U3877 (N_3877,N_2096,N_2758);
nand U3878 (N_3878,N_2593,N_2120);
nand U3879 (N_3879,N_2269,N_2723);
and U3880 (N_3880,N_2453,N_2817);
xor U3881 (N_3881,N_2136,N_2172);
nand U3882 (N_3882,N_2014,N_2217);
and U3883 (N_3883,N_2547,N_2248);
nor U3884 (N_3884,N_2700,N_2675);
nand U3885 (N_3885,N_2988,N_2921);
nor U3886 (N_3886,N_2353,N_2516);
nor U3887 (N_3887,N_2524,N_2146);
or U3888 (N_3888,N_2281,N_2640);
nand U3889 (N_3889,N_2070,N_2579);
nand U3890 (N_3890,N_2482,N_2026);
and U3891 (N_3891,N_2372,N_2485);
xnor U3892 (N_3892,N_2061,N_2237);
or U3893 (N_3893,N_2643,N_2544);
xnor U3894 (N_3894,N_2649,N_2303);
and U3895 (N_3895,N_2791,N_2306);
or U3896 (N_3896,N_2225,N_2128);
xor U3897 (N_3897,N_2421,N_2806);
nand U3898 (N_3898,N_2722,N_2984);
or U3899 (N_3899,N_2383,N_2388);
xor U3900 (N_3900,N_2102,N_2184);
nand U3901 (N_3901,N_2105,N_2521);
nor U3902 (N_3902,N_2523,N_2003);
and U3903 (N_3903,N_2410,N_2690);
or U3904 (N_3904,N_2649,N_2713);
nand U3905 (N_3905,N_2073,N_2108);
or U3906 (N_3906,N_2813,N_2062);
nand U3907 (N_3907,N_2782,N_2948);
nand U3908 (N_3908,N_2576,N_2833);
nor U3909 (N_3909,N_2884,N_2153);
or U3910 (N_3910,N_2382,N_2778);
or U3911 (N_3911,N_2230,N_2602);
nand U3912 (N_3912,N_2227,N_2233);
nand U3913 (N_3913,N_2451,N_2999);
nor U3914 (N_3914,N_2624,N_2124);
and U3915 (N_3915,N_2464,N_2512);
xnor U3916 (N_3916,N_2966,N_2430);
or U3917 (N_3917,N_2398,N_2584);
and U3918 (N_3918,N_2354,N_2300);
nand U3919 (N_3919,N_2799,N_2617);
and U3920 (N_3920,N_2209,N_2756);
or U3921 (N_3921,N_2573,N_2589);
nor U3922 (N_3922,N_2768,N_2987);
xor U3923 (N_3923,N_2692,N_2434);
or U3924 (N_3924,N_2520,N_2823);
xnor U3925 (N_3925,N_2069,N_2023);
xnor U3926 (N_3926,N_2676,N_2280);
or U3927 (N_3927,N_2222,N_2651);
or U3928 (N_3928,N_2947,N_2254);
xor U3929 (N_3929,N_2759,N_2438);
and U3930 (N_3930,N_2118,N_2156);
and U3931 (N_3931,N_2412,N_2748);
nor U3932 (N_3932,N_2357,N_2344);
or U3933 (N_3933,N_2827,N_2729);
nor U3934 (N_3934,N_2698,N_2066);
nand U3935 (N_3935,N_2654,N_2799);
nand U3936 (N_3936,N_2298,N_2476);
xor U3937 (N_3937,N_2832,N_2869);
nor U3938 (N_3938,N_2224,N_2260);
and U3939 (N_3939,N_2733,N_2119);
nor U3940 (N_3940,N_2829,N_2390);
nor U3941 (N_3941,N_2425,N_2106);
xor U3942 (N_3942,N_2897,N_2458);
and U3943 (N_3943,N_2900,N_2354);
and U3944 (N_3944,N_2645,N_2278);
or U3945 (N_3945,N_2719,N_2279);
nor U3946 (N_3946,N_2691,N_2685);
nor U3947 (N_3947,N_2314,N_2446);
or U3948 (N_3948,N_2699,N_2006);
nand U3949 (N_3949,N_2464,N_2298);
nand U3950 (N_3950,N_2389,N_2192);
xnor U3951 (N_3951,N_2936,N_2068);
nand U3952 (N_3952,N_2126,N_2422);
nand U3953 (N_3953,N_2592,N_2566);
and U3954 (N_3954,N_2455,N_2626);
nand U3955 (N_3955,N_2919,N_2253);
nand U3956 (N_3956,N_2047,N_2304);
xnor U3957 (N_3957,N_2184,N_2063);
nand U3958 (N_3958,N_2549,N_2440);
nor U3959 (N_3959,N_2045,N_2154);
nand U3960 (N_3960,N_2272,N_2596);
and U3961 (N_3961,N_2804,N_2489);
and U3962 (N_3962,N_2581,N_2242);
nor U3963 (N_3963,N_2746,N_2135);
nor U3964 (N_3964,N_2206,N_2386);
xnor U3965 (N_3965,N_2687,N_2682);
xnor U3966 (N_3966,N_2755,N_2847);
nor U3967 (N_3967,N_2639,N_2510);
nor U3968 (N_3968,N_2246,N_2649);
xor U3969 (N_3969,N_2164,N_2420);
and U3970 (N_3970,N_2665,N_2143);
and U3971 (N_3971,N_2343,N_2250);
nor U3972 (N_3972,N_2790,N_2729);
nand U3973 (N_3973,N_2504,N_2247);
or U3974 (N_3974,N_2064,N_2702);
xnor U3975 (N_3975,N_2316,N_2757);
nor U3976 (N_3976,N_2037,N_2756);
nand U3977 (N_3977,N_2199,N_2583);
or U3978 (N_3978,N_2066,N_2160);
and U3979 (N_3979,N_2461,N_2584);
and U3980 (N_3980,N_2624,N_2391);
and U3981 (N_3981,N_2760,N_2273);
xor U3982 (N_3982,N_2223,N_2083);
or U3983 (N_3983,N_2169,N_2425);
or U3984 (N_3984,N_2771,N_2558);
nor U3985 (N_3985,N_2332,N_2213);
and U3986 (N_3986,N_2920,N_2262);
nand U3987 (N_3987,N_2287,N_2806);
nor U3988 (N_3988,N_2996,N_2430);
and U3989 (N_3989,N_2428,N_2564);
nand U3990 (N_3990,N_2923,N_2792);
nor U3991 (N_3991,N_2970,N_2537);
and U3992 (N_3992,N_2603,N_2449);
xnor U3993 (N_3993,N_2939,N_2326);
nor U3994 (N_3994,N_2234,N_2481);
nand U3995 (N_3995,N_2989,N_2977);
xor U3996 (N_3996,N_2750,N_2283);
nand U3997 (N_3997,N_2890,N_2072);
or U3998 (N_3998,N_2826,N_2036);
or U3999 (N_3999,N_2687,N_2458);
or U4000 (N_4000,N_3355,N_3981);
or U4001 (N_4001,N_3433,N_3964);
or U4002 (N_4002,N_3026,N_3604);
and U4003 (N_4003,N_3375,N_3987);
nand U4004 (N_4004,N_3528,N_3037);
nor U4005 (N_4005,N_3845,N_3971);
or U4006 (N_4006,N_3113,N_3295);
xnor U4007 (N_4007,N_3319,N_3051);
nor U4008 (N_4008,N_3048,N_3975);
nand U4009 (N_4009,N_3960,N_3665);
nor U4010 (N_4010,N_3261,N_3818);
xnor U4011 (N_4011,N_3311,N_3111);
and U4012 (N_4012,N_3153,N_3911);
and U4013 (N_4013,N_3614,N_3378);
nand U4014 (N_4014,N_3786,N_3748);
nor U4015 (N_4015,N_3112,N_3650);
nand U4016 (N_4016,N_3227,N_3186);
or U4017 (N_4017,N_3585,N_3451);
nor U4018 (N_4018,N_3538,N_3092);
nor U4019 (N_4019,N_3773,N_3126);
nor U4020 (N_4020,N_3966,N_3948);
or U4021 (N_4021,N_3997,N_3065);
nand U4022 (N_4022,N_3937,N_3656);
or U4023 (N_4023,N_3539,N_3744);
nor U4024 (N_4024,N_3624,N_3146);
nand U4025 (N_4025,N_3853,N_3235);
and U4026 (N_4026,N_3961,N_3769);
or U4027 (N_4027,N_3492,N_3803);
xor U4028 (N_4028,N_3586,N_3014);
xor U4029 (N_4029,N_3380,N_3565);
nand U4030 (N_4030,N_3663,N_3875);
or U4031 (N_4031,N_3495,N_3429);
nor U4032 (N_4032,N_3594,N_3169);
and U4033 (N_4033,N_3731,N_3354);
nand U4034 (N_4034,N_3298,N_3816);
nor U4035 (N_4035,N_3001,N_3088);
nor U4036 (N_4036,N_3511,N_3681);
xnor U4037 (N_4037,N_3794,N_3042);
xnor U4038 (N_4038,N_3920,N_3487);
or U4039 (N_4039,N_3182,N_3030);
and U4040 (N_4040,N_3011,N_3583);
nand U4041 (N_4041,N_3189,N_3788);
xor U4042 (N_4042,N_3757,N_3469);
or U4043 (N_4043,N_3256,N_3637);
or U4044 (N_4044,N_3581,N_3108);
xor U4045 (N_4045,N_3303,N_3062);
nand U4046 (N_4046,N_3313,N_3868);
nand U4047 (N_4047,N_3117,N_3489);
nor U4048 (N_4048,N_3806,N_3310);
xnor U4049 (N_4049,N_3357,N_3172);
nor U4050 (N_4050,N_3903,N_3345);
or U4051 (N_4051,N_3555,N_3279);
nor U4052 (N_4052,N_3363,N_3050);
xor U4053 (N_4053,N_3139,N_3213);
nor U4054 (N_4054,N_3796,N_3337);
or U4055 (N_4055,N_3943,N_3514);
xor U4056 (N_4056,N_3450,N_3952);
or U4057 (N_4057,N_3175,N_3499);
nor U4058 (N_4058,N_3630,N_3567);
nor U4059 (N_4059,N_3304,N_3435);
or U4060 (N_4060,N_3939,N_3106);
and U4061 (N_4061,N_3749,N_3922);
and U4062 (N_4062,N_3084,N_3606);
nor U4063 (N_4063,N_3801,N_3196);
nand U4064 (N_4064,N_3289,N_3554);
nand U4065 (N_4065,N_3183,N_3340);
nand U4066 (N_4066,N_3129,N_3880);
or U4067 (N_4067,N_3927,N_3835);
nand U4068 (N_4068,N_3385,N_3694);
nand U4069 (N_4069,N_3364,N_3655);
and U4070 (N_4070,N_3725,N_3610);
or U4071 (N_4071,N_3959,N_3376);
nor U4072 (N_4072,N_3527,N_3382);
nand U4073 (N_4073,N_3659,N_3817);
nand U4074 (N_4074,N_3645,N_3603);
and U4075 (N_4075,N_3251,N_3431);
xor U4076 (N_4076,N_3432,N_3219);
nand U4077 (N_4077,N_3592,N_3596);
or U4078 (N_4078,N_3359,N_3902);
nand U4079 (N_4079,N_3881,N_3068);
nor U4080 (N_4080,N_3346,N_3910);
nand U4081 (N_4081,N_3210,N_3632);
and U4082 (N_4082,N_3023,N_3244);
nand U4083 (N_4083,N_3043,N_3755);
and U4084 (N_4084,N_3970,N_3674);
and U4085 (N_4085,N_3468,N_3577);
xor U4086 (N_4086,N_3832,N_3841);
nand U4087 (N_4087,N_3163,N_3718);
and U4088 (N_4088,N_3497,N_3621);
nand U4089 (N_4089,N_3504,N_3214);
or U4090 (N_4090,N_3522,N_3033);
nand U4091 (N_4091,N_3523,N_3562);
nand U4092 (N_4092,N_3820,N_3849);
nor U4093 (N_4093,N_3669,N_3609);
or U4094 (N_4094,N_3181,N_3118);
nand U4095 (N_4095,N_3142,N_3616);
or U4096 (N_4096,N_3662,N_3459);
xnor U4097 (N_4097,N_3929,N_3334);
and U4098 (N_4098,N_3737,N_3756);
xor U4099 (N_4099,N_3263,N_3713);
or U4100 (N_4100,N_3206,N_3485);
nand U4101 (N_4101,N_3388,N_3125);
and U4102 (N_4102,N_3253,N_3447);
or U4103 (N_4103,N_3016,N_3283);
xnor U4104 (N_4104,N_3266,N_3984);
or U4105 (N_4105,N_3776,N_3781);
xor U4106 (N_4106,N_3123,N_3983);
nand U4107 (N_4107,N_3184,N_3002);
nor U4108 (N_4108,N_3804,N_3954);
xor U4109 (N_4109,N_3573,N_3735);
nand U4110 (N_4110,N_3063,N_3278);
or U4111 (N_4111,N_3782,N_3208);
nand U4112 (N_4112,N_3484,N_3255);
nand U4113 (N_4113,N_3454,N_3199);
nand U4114 (N_4114,N_3398,N_3942);
and U4115 (N_4115,N_3322,N_3874);
nor U4116 (N_4116,N_3321,N_3453);
or U4117 (N_4117,N_3611,N_3416);
xor U4118 (N_4118,N_3374,N_3353);
and U4119 (N_4119,N_3140,N_3720);
or U4120 (N_4120,N_3526,N_3563);
or U4121 (N_4121,N_3542,N_3272);
or U4122 (N_4122,N_3015,N_3933);
nand U4123 (N_4123,N_3275,N_3480);
xor U4124 (N_4124,N_3286,N_3017);
xor U4125 (N_4125,N_3906,N_3414);
xnor U4126 (N_4126,N_3895,N_3722);
and U4127 (N_4127,N_3209,N_3701);
nor U4128 (N_4128,N_3985,N_3925);
and U4129 (N_4129,N_3391,N_3934);
and U4130 (N_4130,N_3932,N_3884);
nor U4131 (N_4131,N_3540,N_3191);
and U4132 (N_4132,N_3067,N_3162);
xnor U4133 (N_4133,N_3945,N_3684);
xor U4134 (N_4134,N_3423,N_3185);
xnor U4135 (N_4135,N_3056,N_3203);
nand U4136 (N_4136,N_3673,N_3010);
nand U4137 (N_4137,N_3282,N_3246);
xnor U4138 (N_4138,N_3814,N_3928);
nand U4139 (N_4139,N_3605,N_3443);
nor U4140 (N_4140,N_3697,N_3838);
or U4141 (N_4141,N_3369,N_3116);
nand U4142 (N_4142,N_3893,N_3020);
xor U4143 (N_4143,N_3520,N_3530);
xnor U4144 (N_4144,N_3615,N_3348);
nor U4145 (N_4145,N_3025,N_3482);
xor U4146 (N_4146,N_3765,N_3505);
xnor U4147 (N_4147,N_3407,N_3548);
or U4148 (N_4148,N_3897,N_3440);
xor U4149 (N_4149,N_3613,N_3559);
or U4150 (N_4150,N_3836,N_3869);
xor U4151 (N_4151,N_3711,N_3785);
xor U4152 (N_4152,N_3972,N_3031);
nand U4153 (N_4153,N_3418,N_3233);
or U4154 (N_4154,N_3742,N_3270);
nand U4155 (N_4155,N_3865,N_3161);
xnor U4156 (N_4156,N_3561,N_3202);
or U4157 (N_4157,N_3822,N_3783);
nand U4158 (N_4158,N_3992,N_3753);
or U4159 (N_4159,N_3634,N_3517);
or U4160 (N_4160,N_3059,N_3515);
nor U4161 (N_4161,N_3686,N_3029);
or U4162 (N_4162,N_3022,N_3411);
xnor U4163 (N_4163,N_3779,N_3508);
and U4164 (N_4164,N_3807,N_3723);
nor U4165 (N_4165,N_3847,N_3296);
or U4166 (N_4166,N_3390,N_3598);
or U4167 (N_4167,N_3490,N_3507);
nand U4168 (N_4168,N_3844,N_3264);
and U4169 (N_4169,N_3223,N_3541);
or U4170 (N_4170,N_3128,N_3285);
nand U4171 (N_4171,N_3446,N_3076);
or U4172 (N_4172,N_3620,N_3240);
nor U4173 (N_4173,N_3365,N_3758);
and U4174 (N_4174,N_3070,N_3930);
or U4175 (N_4175,N_3165,N_3114);
and U4176 (N_4176,N_3372,N_3915);
nand U4177 (N_4177,N_3081,N_3371);
or U4178 (N_4178,N_3350,N_3940);
xnor U4179 (N_4179,N_3589,N_3766);
or U4180 (N_4180,N_3093,N_3104);
and U4181 (N_4181,N_3591,N_3397);
nand U4182 (N_4182,N_3545,N_3462);
and U4183 (N_4183,N_3052,N_3619);
or U4184 (N_4184,N_3837,N_3087);
nor U4185 (N_4185,N_3236,N_3300);
and U4186 (N_4186,N_3965,N_3077);
nand U4187 (N_4187,N_3623,N_3234);
xnor U4188 (N_4188,N_3245,N_3383);
or U4189 (N_4189,N_3103,N_3908);
nor U4190 (N_4190,N_3276,N_3360);
nor U4191 (N_4191,N_3228,N_3980);
or U4192 (N_4192,N_3299,N_3652);
xnor U4193 (N_4193,N_3819,N_3976);
nand U4194 (N_4194,N_3789,N_3848);
and U4195 (N_4195,N_3341,N_3878);
and U4196 (N_4196,N_3898,N_3339);
xor U4197 (N_4197,N_3316,N_3840);
nand U4198 (N_4198,N_3644,N_3852);
xnor U4199 (N_4199,N_3639,N_3994);
xor U4200 (N_4200,N_3327,N_3373);
xnor U4201 (N_4201,N_3368,N_3590);
and U4202 (N_4202,N_3347,N_3085);
nand U4203 (N_4203,N_3900,N_3225);
nand U4204 (N_4204,N_3524,N_3728);
and U4205 (N_4205,N_3741,N_3699);
nor U4206 (N_4206,N_3419,N_3361);
or U4207 (N_4207,N_3131,N_3580);
or U4208 (N_4208,N_3716,N_3323);
and U4209 (N_4209,N_3366,N_3399);
and U4210 (N_4210,N_3506,N_3705);
or U4211 (N_4211,N_3457,N_3293);
xor U4212 (N_4212,N_3177,N_3536);
xnor U4213 (N_4213,N_3990,N_3094);
nor U4214 (N_4214,N_3473,N_3171);
nor U4215 (N_4215,N_3086,N_3885);
and U4216 (N_4216,N_3254,N_3154);
nand U4217 (N_4217,N_3465,N_3805);
and U4218 (N_4218,N_3207,N_3557);
nand U4219 (N_4219,N_3386,N_3491);
nor U4220 (N_4220,N_3680,N_3216);
nor U4221 (N_4221,N_3257,N_3335);
and U4222 (N_4222,N_3120,N_3102);
or U4223 (N_4223,N_3973,N_3099);
nor U4224 (N_4224,N_3799,N_3892);
or U4225 (N_4225,N_3978,N_3863);
or U4226 (N_4226,N_3122,N_3151);
or U4227 (N_4227,N_3860,N_3008);
nor U4228 (N_4228,N_3879,N_3058);
nor U4229 (N_4229,N_3618,N_3888);
xnor U4230 (N_4230,N_3362,N_3518);
nor U4231 (N_4231,N_3608,N_3115);
and U4232 (N_4232,N_3274,N_3824);
nor U4233 (N_4233,N_3534,N_3124);
nor U4234 (N_4234,N_3325,N_3951);
and U4235 (N_4235,N_3999,N_3287);
or U4236 (N_4236,N_3269,N_3883);
xor U4237 (N_4237,N_3859,N_3096);
nor U4238 (N_4238,N_3670,N_3239);
and U4239 (N_4239,N_3343,N_3483);
nor U4240 (N_4240,N_3509,N_3479);
nor U4241 (N_4241,N_3552,N_3570);
or U4242 (N_4242,N_3501,N_3463);
nor U4243 (N_4243,N_3729,N_3370);
xnor U4244 (N_4244,N_3628,N_3587);
nor U4245 (N_4245,N_3704,N_3963);
nor U4246 (N_4246,N_3698,N_3944);
or U4247 (N_4247,N_3834,N_3212);
nor U4248 (N_4248,N_3715,N_3761);
nor U4249 (N_4249,N_3743,N_3647);
nor U4250 (N_4250,N_3800,N_3247);
and U4251 (N_4251,N_3260,N_3710);
xor U4252 (N_4252,N_3080,N_3547);
or U4253 (N_4253,N_3168,N_3073);
nand U4254 (N_4254,N_3622,N_3935);
nor U4255 (N_4255,N_3467,N_3226);
or U4256 (N_4256,N_3143,N_3958);
xor U4257 (N_4257,N_3338,N_3071);
or U4258 (N_4258,N_3531,N_3019);
nor U4259 (N_4259,N_3053,N_3222);
nor U4260 (N_4260,N_3192,N_3866);
nand U4261 (N_4261,N_3302,N_3923);
or U4262 (N_4262,N_3045,N_3503);
and U4263 (N_4263,N_3689,N_3405);
nor U4264 (N_4264,N_3919,N_3747);
nand U4265 (N_4265,N_3588,N_3061);
or U4266 (N_4266,N_3455,N_3107);
nand U4267 (N_4267,N_3018,N_3460);
nor U4268 (N_4268,N_3809,N_3315);
or U4269 (N_4269,N_3657,N_3119);
and U4270 (N_4270,N_3352,N_3825);
and U4271 (N_4271,N_3317,N_3721);
or U4272 (N_4272,N_3344,N_3329);
nand U4273 (N_4273,N_3166,N_3201);
nor U4274 (N_4274,N_3549,N_3089);
nor U4275 (N_4275,N_3763,N_3535);
nand U4276 (N_4276,N_3082,N_3738);
and U4277 (N_4277,N_3989,N_3791);
and U4278 (N_4278,N_3007,N_3633);
nor U4279 (N_4279,N_3195,N_3851);
nand U4280 (N_4280,N_3601,N_3823);
xor U4281 (N_4281,N_3708,N_3496);
nor U4282 (N_4282,N_3850,N_3798);
nand U4283 (N_4283,N_3510,N_3179);
and U4284 (N_4284,N_3013,N_3696);
nor U4285 (N_4285,N_3069,N_3907);
nand U4286 (N_4286,N_3280,N_3896);
nand U4287 (N_4287,N_3564,N_3533);
xnor U4288 (N_4288,N_3387,N_3294);
nor U4289 (N_4289,N_3733,N_3444);
nand U4290 (N_4290,N_3049,N_3148);
or U4291 (N_4291,N_3617,N_3730);
or U4292 (N_4292,N_3946,N_3947);
and U4293 (N_4293,N_3100,N_3660);
or U4294 (N_4294,N_3241,N_3413);
xnor U4295 (N_4295,N_3475,N_3599);
or U4296 (N_4296,N_3005,N_3072);
or U4297 (N_4297,N_3727,N_3035);
xnor U4298 (N_4298,N_3795,N_3712);
xor U4299 (N_4299,N_3941,N_3318);
nor U4300 (N_4300,N_3190,N_3575);
or U4301 (N_4301,N_3187,N_3150);
or U4302 (N_4302,N_3726,N_3894);
nor U4303 (N_4303,N_3250,N_3105);
or U4304 (N_4304,N_3331,N_3991);
and U4305 (N_4305,N_3631,N_3178);
nor U4306 (N_4306,N_3090,N_3332);
nor U4307 (N_4307,N_3493,N_3595);
nand U4308 (N_4308,N_3424,N_3936);
or U4309 (N_4309,N_3039,N_3764);
and U4310 (N_4310,N_3890,N_3926);
xnor U4311 (N_4311,N_3243,N_3476);
and U4312 (N_4312,N_3231,N_3403);
nand U4313 (N_4313,N_3464,N_3544);
and U4314 (N_4314,N_3995,N_3215);
and U4315 (N_4315,N_3754,N_3145);
xnor U4316 (N_4316,N_3734,N_3034);
nor U4317 (N_4317,N_3717,N_3091);
nor U4318 (N_4318,N_3676,N_3205);
and U4319 (N_4319,N_3430,N_3158);
nor U4320 (N_4320,N_3719,N_3217);
nand U4321 (N_4321,N_3356,N_3427);
xnor U4322 (N_4322,N_3882,N_3982);
xor U4323 (N_4323,N_3974,N_3027);
xor U4324 (N_4324,N_3872,N_3400);
and U4325 (N_4325,N_3078,N_3180);
nor U4326 (N_4326,N_3358,N_3060);
nand U4327 (N_4327,N_3762,N_3760);
and U4328 (N_4328,N_3500,N_3558);
xnor U4329 (N_4329,N_3855,N_3675);
and U4330 (N_4330,N_3924,N_3157);
or U4331 (N_4331,N_3640,N_3532);
or U4332 (N_4332,N_3551,N_3569);
nor U4333 (N_4333,N_3470,N_3351);
or U4334 (N_4334,N_3649,N_3408);
or U4335 (N_4335,N_3312,N_3211);
nand U4336 (N_4336,N_3685,N_3194);
and U4337 (N_4337,N_3095,N_3248);
or U4338 (N_4338,N_3938,N_3229);
and U4339 (N_4339,N_3778,N_3702);
nand U4340 (N_4340,N_3271,N_3775);
nor U4341 (N_4341,N_3658,N_3308);
and U4342 (N_4342,N_3955,N_3164);
xnor U4343 (N_4343,N_3097,N_3170);
or U4344 (N_4344,N_3474,N_3133);
nand U4345 (N_4345,N_3349,N_3284);
nand U4346 (N_4346,N_3324,N_3854);
nor U4347 (N_4347,N_3695,N_3422);
nand U4348 (N_4348,N_3237,N_3367);
xnor U4349 (N_4349,N_3529,N_3913);
or U4350 (N_4350,N_3574,N_3147);
nand U4351 (N_4351,N_3259,N_3305);
and U4352 (N_4352,N_3041,N_3130);
or U4353 (N_4353,N_3320,N_3667);
xnor U4354 (N_4354,N_3826,N_3498);
xnor U4355 (N_4355,N_3486,N_3075);
or U4356 (N_4356,N_3602,N_3404);
xor U4357 (N_4357,N_3739,N_3750);
xor U4358 (N_4358,N_3714,N_3521);
nor U4359 (N_4359,N_3745,N_3481);
and U4360 (N_4360,N_3379,N_3003);
nand U4361 (N_4361,N_3813,N_3771);
nor U4362 (N_4362,N_3571,N_3625);
nand U4363 (N_4363,N_3032,N_3998);
and U4364 (N_4364,N_3342,N_3988);
xor U4365 (N_4365,N_3000,N_3047);
or U4366 (N_4366,N_3384,N_3333);
xor U4367 (N_4367,N_3843,N_3083);
xor U4368 (N_4368,N_3802,N_3876);
or U4369 (N_4369,N_3668,N_3395);
nor U4370 (N_4370,N_3155,N_3905);
and U4371 (N_4371,N_3693,N_3054);
xnor U4372 (N_4372,N_3780,N_3636);
or U4373 (N_4373,N_3292,N_3870);
and U4374 (N_4374,N_3218,N_3230);
nand U4375 (N_4375,N_3004,N_3627);
and U4376 (N_4376,N_3436,N_3193);
and U4377 (N_4377,N_3098,N_3830);
nor U4378 (N_4378,N_3409,N_3471);
and U4379 (N_4379,N_3301,N_3267);
and U4380 (N_4380,N_3550,N_3642);
xor U4381 (N_4381,N_3441,N_3572);
nand U4382 (N_4382,N_3846,N_3160);
nor U4383 (N_4383,N_3525,N_3537);
or U4384 (N_4384,N_3381,N_3024);
and U4385 (N_4385,N_3314,N_3173);
and U4386 (N_4386,N_3415,N_3220);
xor U4387 (N_4387,N_3707,N_3904);
nor U4388 (N_4388,N_3736,N_3873);
or U4389 (N_4389,N_3767,N_3831);
xnor U4390 (N_4390,N_3238,N_3821);
xor U4391 (N_4391,N_3768,N_3137);
xnor U4392 (N_4392,N_3425,N_3687);
xnor U4393 (N_4393,N_3445,N_3774);
nor U4394 (N_4394,N_3977,N_3597);
xor U4395 (N_4395,N_3174,N_3144);
and U4396 (N_4396,N_3957,N_3671);
xor U4397 (N_4397,N_3028,N_3224);
xor U4398 (N_4398,N_3901,N_3437);
or U4399 (N_4399,N_3553,N_3864);
nor U4400 (N_4400,N_3412,N_3740);
xnor U4401 (N_4401,N_3653,N_3576);
nor U4402 (N_4402,N_3967,N_3249);
xnor U4403 (N_4403,N_3629,N_3394);
and U4404 (N_4404,N_3962,N_3159);
and U4405 (N_4405,N_3772,N_3833);
or U4406 (N_4406,N_3953,N_3921);
nor U4407 (N_4407,N_3044,N_3428);
or U4408 (N_4408,N_3221,N_3456);
or U4409 (N_4409,N_3691,N_3519);
nand U4410 (N_4410,N_3461,N_3152);
or U4411 (N_4411,N_3709,N_3265);
or U4412 (N_4412,N_3262,N_3135);
or U4413 (N_4413,N_3829,N_3477);
and U4414 (N_4414,N_3040,N_3654);
or U4415 (N_4415,N_3560,N_3074);
nor U4416 (N_4416,N_3101,N_3986);
nor U4417 (N_4417,N_3887,N_3751);
xnor U4418 (N_4418,N_3328,N_3273);
and U4419 (N_4419,N_3410,N_3664);
xor U4420 (N_4420,N_3889,N_3306);
or U4421 (N_4421,N_3288,N_3827);
xor U4422 (N_4422,N_3336,N_3198);
or U4423 (N_4423,N_3466,N_3607);
nor U4424 (N_4424,N_3808,N_3784);
nor U4425 (N_4425,N_3188,N_3512);
and U4426 (N_4426,N_3679,N_3856);
nand U4427 (N_4427,N_3797,N_3307);
or U4428 (N_4428,N_3886,N_3478);
xnor U4429 (N_4429,N_3330,N_3012);
xnor U4430 (N_4430,N_3472,N_3417);
nand U4431 (N_4431,N_3579,N_3197);
xnor U4432 (N_4432,N_3156,N_3393);
nor U4433 (N_4433,N_3677,N_3449);
and U4434 (N_4434,N_3917,N_3706);
and U4435 (N_4435,N_3121,N_3584);
or U4436 (N_4436,N_3448,N_3309);
or U4437 (N_4437,N_3732,N_3899);
xnor U4438 (N_4438,N_3626,N_3516);
or U4439 (N_4439,N_3666,N_3651);
nand U4440 (N_4440,N_3290,N_3252);
nor U4441 (N_4441,N_3127,N_3600);
nand U4442 (N_4442,N_3232,N_3956);
nand U4443 (N_4443,N_3692,N_3912);
nand U4444 (N_4444,N_3057,N_3683);
nor U4445 (N_4445,N_3167,N_3421);
and U4446 (N_4446,N_3064,N_3700);
or U4447 (N_4447,N_3996,N_3724);
nand U4448 (N_4448,N_3839,N_3055);
nor U4449 (N_4449,N_3858,N_3066);
and U4450 (N_4450,N_3021,N_3993);
nor U4451 (N_4451,N_3661,N_3877);
nor U4452 (N_4452,N_3777,N_3787);
and U4453 (N_4453,N_3009,N_3950);
nor U4454 (N_4454,N_3036,N_3458);
nand U4455 (N_4455,N_3268,N_3006);
or U4456 (N_4456,N_3568,N_3648);
or U4457 (N_4457,N_3812,N_3862);
or U4458 (N_4458,N_3109,N_3377);
or U4459 (N_4459,N_3678,N_3578);
nor U4460 (N_4460,N_3969,N_3909);
and U4461 (N_4461,N_3566,N_3582);
and U4462 (N_4462,N_3703,N_3635);
and U4463 (N_4463,N_3204,N_3857);
nand U4464 (N_4464,N_3326,N_3038);
and U4465 (N_4465,N_3392,N_3914);
or U4466 (N_4466,N_3138,N_3793);
and U4467 (N_4467,N_3752,N_3646);
and U4468 (N_4468,N_3949,N_3079);
and U4469 (N_4469,N_3452,N_3931);
and U4470 (N_4470,N_3277,N_3811);
or U4471 (N_4471,N_3396,N_3442);
and U4472 (N_4472,N_3815,N_3426);
xnor U4473 (N_4473,N_3502,N_3389);
nand U4474 (N_4474,N_3828,N_3149);
or U4475 (N_4475,N_3439,N_3641);
xor U4476 (N_4476,N_3891,N_3401);
or U4477 (N_4477,N_3438,N_3871);
nand U4478 (N_4478,N_3867,N_3494);
nand U4479 (N_4479,N_3688,N_3790);
xor U4480 (N_4480,N_3132,N_3638);
or U4481 (N_4481,N_3546,N_3258);
xnor U4482 (N_4482,N_3291,N_3979);
or U4483 (N_4483,N_3242,N_3682);
and U4484 (N_4484,N_3968,N_3770);
nand U4485 (N_4485,N_3281,N_3046);
xnor U4486 (N_4486,N_3792,N_3406);
and U4487 (N_4487,N_3141,N_3861);
and U4488 (N_4488,N_3746,N_3759);
xor U4489 (N_4489,N_3134,N_3110);
or U4490 (N_4490,N_3402,N_3810);
nand U4491 (N_4491,N_3842,N_3690);
and U4492 (N_4492,N_3672,N_3136);
and U4493 (N_4493,N_3513,N_3488);
and U4494 (N_4494,N_3643,N_3543);
nor U4495 (N_4495,N_3556,N_3612);
nor U4496 (N_4496,N_3593,N_3420);
nand U4497 (N_4497,N_3918,N_3297);
and U4498 (N_4498,N_3916,N_3176);
xnor U4499 (N_4499,N_3200,N_3434);
and U4500 (N_4500,N_3983,N_3253);
xnor U4501 (N_4501,N_3198,N_3750);
or U4502 (N_4502,N_3195,N_3721);
nor U4503 (N_4503,N_3928,N_3424);
nand U4504 (N_4504,N_3975,N_3598);
nand U4505 (N_4505,N_3840,N_3295);
nand U4506 (N_4506,N_3942,N_3430);
nand U4507 (N_4507,N_3105,N_3309);
and U4508 (N_4508,N_3799,N_3016);
nor U4509 (N_4509,N_3745,N_3562);
or U4510 (N_4510,N_3924,N_3667);
nand U4511 (N_4511,N_3013,N_3706);
xnor U4512 (N_4512,N_3592,N_3720);
nand U4513 (N_4513,N_3653,N_3409);
and U4514 (N_4514,N_3654,N_3403);
nand U4515 (N_4515,N_3630,N_3836);
xor U4516 (N_4516,N_3258,N_3203);
or U4517 (N_4517,N_3503,N_3941);
or U4518 (N_4518,N_3454,N_3373);
nand U4519 (N_4519,N_3738,N_3861);
nand U4520 (N_4520,N_3266,N_3227);
or U4521 (N_4521,N_3489,N_3342);
nand U4522 (N_4522,N_3975,N_3726);
nor U4523 (N_4523,N_3832,N_3316);
or U4524 (N_4524,N_3130,N_3021);
xnor U4525 (N_4525,N_3572,N_3081);
nor U4526 (N_4526,N_3279,N_3324);
or U4527 (N_4527,N_3361,N_3939);
xor U4528 (N_4528,N_3465,N_3885);
nand U4529 (N_4529,N_3872,N_3773);
xnor U4530 (N_4530,N_3594,N_3251);
nor U4531 (N_4531,N_3492,N_3572);
or U4532 (N_4532,N_3071,N_3249);
or U4533 (N_4533,N_3495,N_3779);
xor U4534 (N_4534,N_3392,N_3570);
xor U4535 (N_4535,N_3175,N_3580);
and U4536 (N_4536,N_3917,N_3855);
nor U4537 (N_4537,N_3968,N_3536);
nor U4538 (N_4538,N_3757,N_3752);
nand U4539 (N_4539,N_3603,N_3136);
nand U4540 (N_4540,N_3963,N_3808);
xor U4541 (N_4541,N_3230,N_3168);
nor U4542 (N_4542,N_3813,N_3542);
or U4543 (N_4543,N_3828,N_3856);
nor U4544 (N_4544,N_3820,N_3256);
xor U4545 (N_4545,N_3666,N_3528);
and U4546 (N_4546,N_3416,N_3148);
xnor U4547 (N_4547,N_3058,N_3727);
xnor U4548 (N_4548,N_3509,N_3967);
nor U4549 (N_4549,N_3053,N_3908);
xnor U4550 (N_4550,N_3716,N_3435);
xnor U4551 (N_4551,N_3623,N_3925);
and U4552 (N_4552,N_3493,N_3303);
xor U4553 (N_4553,N_3532,N_3981);
nand U4554 (N_4554,N_3478,N_3246);
or U4555 (N_4555,N_3497,N_3168);
or U4556 (N_4556,N_3467,N_3790);
or U4557 (N_4557,N_3699,N_3829);
or U4558 (N_4558,N_3171,N_3210);
and U4559 (N_4559,N_3498,N_3829);
xor U4560 (N_4560,N_3481,N_3746);
and U4561 (N_4561,N_3469,N_3716);
xnor U4562 (N_4562,N_3888,N_3308);
and U4563 (N_4563,N_3563,N_3084);
or U4564 (N_4564,N_3616,N_3582);
nor U4565 (N_4565,N_3197,N_3325);
xnor U4566 (N_4566,N_3341,N_3942);
nand U4567 (N_4567,N_3059,N_3939);
nor U4568 (N_4568,N_3689,N_3950);
xnor U4569 (N_4569,N_3838,N_3552);
xnor U4570 (N_4570,N_3871,N_3429);
and U4571 (N_4571,N_3117,N_3477);
and U4572 (N_4572,N_3430,N_3475);
nand U4573 (N_4573,N_3131,N_3266);
and U4574 (N_4574,N_3480,N_3155);
xor U4575 (N_4575,N_3381,N_3213);
nand U4576 (N_4576,N_3952,N_3334);
nor U4577 (N_4577,N_3661,N_3396);
and U4578 (N_4578,N_3676,N_3024);
or U4579 (N_4579,N_3258,N_3679);
and U4580 (N_4580,N_3631,N_3415);
xnor U4581 (N_4581,N_3963,N_3245);
xor U4582 (N_4582,N_3348,N_3276);
or U4583 (N_4583,N_3945,N_3140);
nand U4584 (N_4584,N_3265,N_3280);
or U4585 (N_4585,N_3123,N_3763);
or U4586 (N_4586,N_3578,N_3403);
or U4587 (N_4587,N_3354,N_3561);
nor U4588 (N_4588,N_3069,N_3008);
nor U4589 (N_4589,N_3943,N_3823);
xor U4590 (N_4590,N_3520,N_3409);
or U4591 (N_4591,N_3326,N_3217);
xnor U4592 (N_4592,N_3999,N_3369);
or U4593 (N_4593,N_3016,N_3206);
xnor U4594 (N_4594,N_3800,N_3655);
nor U4595 (N_4595,N_3571,N_3093);
nand U4596 (N_4596,N_3892,N_3937);
and U4597 (N_4597,N_3387,N_3025);
nand U4598 (N_4598,N_3374,N_3880);
or U4599 (N_4599,N_3240,N_3790);
nand U4600 (N_4600,N_3877,N_3066);
xor U4601 (N_4601,N_3198,N_3783);
or U4602 (N_4602,N_3007,N_3446);
and U4603 (N_4603,N_3491,N_3684);
and U4604 (N_4604,N_3615,N_3650);
or U4605 (N_4605,N_3017,N_3020);
or U4606 (N_4606,N_3920,N_3846);
nor U4607 (N_4607,N_3327,N_3533);
xnor U4608 (N_4608,N_3961,N_3478);
or U4609 (N_4609,N_3769,N_3778);
xor U4610 (N_4610,N_3078,N_3560);
nor U4611 (N_4611,N_3233,N_3665);
or U4612 (N_4612,N_3391,N_3695);
xnor U4613 (N_4613,N_3264,N_3709);
and U4614 (N_4614,N_3617,N_3938);
nor U4615 (N_4615,N_3492,N_3407);
xnor U4616 (N_4616,N_3040,N_3870);
or U4617 (N_4617,N_3397,N_3616);
nor U4618 (N_4618,N_3479,N_3083);
xnor U4619 (N_4619,N_3568,N_3219);
nor U4620 (N_4620,N_3550,N_3207);
or U4621 (N_4621,N_3818,N_3477);
nand U4622 (N_4622,N_3036,N_3722);
or U4623 (N_4623,N_3547,N_3519);
nor U4624 (N_4624,N_3538,N_3809);
or U4625 (N_4625,N_3662,N_3666);
and U4626 (N_4626,N_3332,N_3314);
and U4627 (N_4627,N_3645,N_3182);
or U4628 (N_4628,N_3430,N_3011);
and U4629 (N_4629,N_3607,N_3227);
nand U4630 (N_4630,N_3024,N_3493);
nand U4631 (N_4631,N_3267,N_3052);
and U4632 (N_4632,N_3092,N_3005);
xor U4633 (N_4633,N_3808,N_3653);
nor U4634 (N_4634,N_3009,N_3651);
and U4635 (N_4635,N_3055,N_3536);
nand U4636 (N_4636,N_3769,N_3799);
and U4637 (N_4637,N_3419,N_3427);
nand U4638 (N_4638,N_3086,N_3226);
or U4639 (N_4639,N_3205,N_3169);
xor U4640 (N_4640,N_3447,N_3354);
nand U4641 (N_4641,N_3729,N_3317);
nor U4642 (N_4642,N_3529,N_3345);
and U4643 (N_4643,N_3796,N_3166);
nor U4644 (N_4644,N_3953,N_3900);
nor U4645 (N_4645,N_3911,N_3677);
nor U4646 (N_4646,N_3162,N_3627);
xor U4647 (N_4647,N_3648,N_3528);
and U4648 (N_4648,N_3053,N_3563);
and U4649 (N_4649,N_3377,N_3614);
nand U4650 (N_4650,N_3661,N_3954);
xor U4651 (N_4651,N_3688,N_3671);
nor U4652 (N_4652,N_3935,N_3235);
or U4653 (N_4653,N_3020,N_3924);
and U4654 (N_4654,N_3488,N_3963);
xnor U4655 (N_4655,N_3418,N_3238);
xor U4656 (N_4656,N_3824,N_3212);
xor U4657 (N_4657,N_3943,N_3537);
or U4658 (N_4658,N_3064,N_3542);
xor U4659 (N_4659,N_3665,N_3143);
xor U4660 (N_4660,N_3424,N_3402);
and U4661 (N_4661,N_3086,N_3564);
and U4662 (N_4662,N_3052,N_3827);
or U4663 (N_4663,N_3821,N_3557);
nor U4664 (N_4664,N_3569,N_3733);
and U4665 (N_4665,N_3200,N_3625);
and U4666 (N_4666,N_3587,N_3465);
nand U4667 (N_4667,N_3231,N_3840);
nand U4668 (N_4668,N_3128,N_3863);
nand U4669 (N_4669,N_3561,N_3818);
nand U4670 (N_4670,N_3013,N_3732);
xor U4671 (N_4671,N_3425,N_3233);
nand U4672 (N_4672,N_3524,N_3932);
nand U4673 (N_4673,N_3788,N_3344);
or U4674 (N_4674,N_3950,N_3198);
or U4675 (N_4675,N_3889,N_3195);
nand U4676 (N_4676,N_3998,N_3560);
nand U4677 (N_4677,N_3493,N_3509);
xor U4678 (N_4678,N_3181,N_3993);
and U4679 (N_4679,N_3878,N_3057);
nor U4680 (N_4680,N_3557,N_3873);
nor U4681 (N_4681,N_3385,N_3940);
and U4682 (N_4682,N_3052,N_3704);
nor U4683 (N_4683,N_3490,N_3911);
or U4684 (N_4684,N_3016,N_3554);
xnor U4685 (N_4685,N_3268,N_3510);
xnor U4686 (N_4686,N_3864,N_3417);
xnor U4687 (N_4687,N_3982,N_3761);
or U4688 (N_4688,N_3697,N_3212);
and U4689 (N_4689,N_3854,N_3483);
or U4690 (N_4690,N_3330,N_3841);
nand U4691 (N_4691,N_3701,N_3958);
nor U4692 (N_4692,N_3214,N_3656);
xnor U4693 (N_4693,N_3639,N_3720);
or U4694 (N_4694,N_3666,N_3146);
xor U4695 (N_4695,N_3093,N_3482);
or U4696 (N_4696,N_3042,N_3701);
nor U4697 (N_4697,N_3481,N_3884);
nand U4698 (N_4698,N_3128,N_3660);
xnor U4699 (N_4699,N_3013,N_3256);
and U4700 (N_4700,N_3230,N_3984);
and U4701 (N_4701,N_3459,N_3397);
or U4702 (N_4702,N_3369,N_3386);
nor U4703 (N_4703,N_3715,N_3733);
nand U4704 (N_4704,N_3445,N_3277);
and U4705 (N_4705,N_3379,N_3632);
or U4706 (N_4706,N_3629,N_3380);
and U4707 (N_4707,N_3651,N_3544);
xor U4708 (N_4708,N_3038,N_3771);
and U4709 (N_4709,N_3438,N_3054);
nor U4710 (N_4710,N_3712,N_3062);
and U4711 (N_4711,N_3111,N_3258);
nor U4712 (N_4712,N_3701,N_3957);
nand U4713 (N_4713,N_3049,N_3392);
nor U4714 (N_4714,N_3520,N_3182);
and U4715 (N_4715,N_3985,N_3642);
nand U4716 (N_4716,N_3682,N_3291);
or U4717 (N_4717,N_3377,N_3228);
nor U4718 (N_4718,N_3509,N_3840);
nand U4719 (N_4719,N_3209,N_3930);
xor U4720 (N_4720,N_3564,N_3129);
xnor U4721 (N_4721,N_3952,N_3441);
or U4722 (N_4722,N_3464,N_3138);
nor U4723 (N_4723,N_3053,N_3555);
nand U4724 (N_4724,N_3882,N_3866);
nand U4725 (N_4725,N_3926,N_3076);
nor U4726 (N_4726,N_3109,N_3399);
nand U4727 (N_4727,N_3310,N_3240);
xnor U4728 (N_4728,N_3956,N_3363);
nor U4729 (N_4729,N_3825,N_3367);
nor U4730 (N_4730,N_3411,N_3349);
nand U4731 (N_4731,N_3330,N_3744);
nor U4732 (N_4732,N_3745,N_3963);
xnor U4733 (N_4733,N_3700,N_3214);
and U4734 (N_4734,N_3656,N_3256);
nand U4735 (N_4735,N_3650,N_3015);
or U4736 (N_4736,N_3351,N_3022);
or U4737 (N_4737,N_3132,N_3035);
nor U4738 (N_4738,N_3733,N_3230);
and U4739 (N_4739,N_3610,N_3442);
nand U4740 (N_4740,N_3385,N_3008);
and U4741 (N_4741,N_3531,N_3262);
nand U4742 (N_4742,N_3629,N_3773);
and U4743 (N_4743,N_3847,N_3393);
xor U4744 (N_4744,N_3973,N_3733);
nand U4745 (N_4745,N_3121,N_3439);
nor U4746 (N_4746,N_3088,N_3809);
xnor U4747 (N_4747,N_3532,N_3471);
or U4748 (N_4748,N_3897,N_3019);
nand U4749 (N_4749,N_3601,N_3038);
and U4750 (N_4750,N_3024,N_3296);
xor U4751 (N_4751,N_3297,N_3495);
and U4752 (N_4752,N_3111,N_3809);
and U4753 (N_4753,N_3723,N_3745);
xor U4754 (N_4754,N_3055,N_3968);
nor U4755 (N_4755,N_3688,N_3695);
nor U4756 (N_4756,N_3512,N_3310);
xor U4757 (N_4757,N_3205,N_3716);
xor U4758 (N_4758,N_3398,N_3852);
or U4759 (N_4759,N_3576,N_3920);
or U4760 (N_4760,N_3895,N_3775);
and U4761 (N_4761,N_3716,N_3988);
nand U4762 (N_4762,N_3749,N_3286);
and U4763 (N_4763,N_3639,N_3462);
nor U4764 (N_4764,N_3638,N_3581);
xor U4765 (N_4765,N_3320,N_3882);
nor U4766 (N_4766,N_3343,N_3827);
and U4767 (N_4767,N_3132,N_3462);
nor U4768 (N_4768,N_3138,N_3578);
xor U4769 (N_4769,N_3015,N_3902);
or U4770 (N_4770,N_3871,N_3087);
nand U4771 (N_4771,N_3484,N_3226);
xnor U4772 (N_4772,N_3182,N_3675);
or U4773 (N_4773,N_3017,N_3656);
or U4774 (N_4774,N_3772,N_3809);
xnor U4775 (N_4775,N_3104,N_3408);
nor U4776 (N_4776,N_3617,N_3698);
or U4777 (N_4777,N_3332,N_3542);
xnor U4778 (N_4778,N_3607,N_3005);
and U4779 (N_4779,N_3579,N_3255);
or U4780 (N_4780,N_3352,N_3417);
nor U4781 (N_4781,N_3123,N_3015);
nor U4782 (N_4782,N_3669,N_3708);
nor U4783 (N_4783,N_3041,N_3509);
xnor U4784 (N_4784,N_3885,N_3260);
and U4785 (N_4785,N_3835,N_3786);
nand U4786 (N_4786,N_3467,N_3787);
or U4787 (N_4787,N_3779,N_3859);
nor U4788 (N_4788,N_3611,N_3932);
or U4789 (N_4789,N_3339,N_3423);
nor U4790 (N_4790,N_3976,N_3710);
xnor U4791 (N_4791,N_3308,N_3337);
xor U4792 (N_4792,N_3970,N_3281);
nor U4793 (N_4793,N_3230,N_3716);
or U4794 (N_4794,N_3160,N_3503);
and U4795 (N_4795,N_3780,N_3550);
and U4796 (N_4796,N_3353,N_3930);
xor U4797 (N_4797,N_3062,N_3502);
xor U4798 (N_4798,N_3290,N_3275);
or U4799 (N_4799,N_3738,N_3503);
and U4800 (N_4800,N_3763,N_3311);
or U4801 (N_4801,N_3317,N_3050);
and U4802 (N_4802,N_3653,N_3877);
nor U4803 (N_4803,N_3169,N_3367);
and U4804 (N_4804,N_3871,N_3117);
nor U4805 (N_4805,N_3425,N_3521);
or U4806 (N_4806,N_3768,N_3375);
nor U4807 (N_4807,N_3036,N_3112);
nand U4808 (N_4808,N_3877,N_3614);
xnor U4809 (N_4809,N_3979,N_3755);
and U4810 (N_4810,N_3207,N_3803);
and U4811 (N_4811,N_3993,N_3007);
and U4812 (N_4812,N_3520,N_3085);
and U4813 (N_4813,N_3977,N_3273);
nand U4814 (N_4814,N_3165,N_3864);
nor U4815 (N_4815,N_3403,N_3220);
nand U4816 (N_4816,N_3395,N_3942);
nor U4817 (N_4817,N_3202,N_3962);
nor U4818 (N_4818,N_3126,N_3613);
nor U4819 (N_4819,N_3296,N_3702);
and U4820 (N_4820,N_3441,N_3814);
and U4821 (N_4821,N_3906,N_3784);
nor U4822 (N_4822,N_3288,N_3922);
nor U4823 (N_4823,N_3040,N_3884);
or U4824 (N_4824,N_3797,N_3718);
and U4825 (N_4825,N_3051,N_3292);
or U4826 (N_4826,N_3448,N_3045);
xor U4827 (N_4827,N_3759,N_3771);
and U4828 (N_4828,N_3022,N_3570);
or U4829 (N_4829,N_3373,N_3986);
and U4830 (N_4830,N_3967,N_3871);
and U4831 (N_4831,N_3420,N_3149);
or U4832 (N_4832,N_3865,N_3072);
and U4833 (N_4833,N_3363,N_3118);
nand U4834 (N_4834,N_3969,N_3148);
xor U4835 (N_4835,N_3831,N_3814);
nand U4836 (N_4836,N_3610,N_3998);
nand U4837 (N_4837,N_3182,N_3414);
nand U4838 (N_4838,N_3213,N_3993);
nor U4839 (N_4839,N_3843,N_3321);
and U4840 (N_4840,N_3509,N_3538);
nor U4841 (N_4841,N_3579,N_3220);
or U4842 (N_4842,N_3774,N_3906);
or U4843 (N_4843,N_3167,N_3637);
xor U4844 (N_4844,N_3973,N_3664);
nor U4845 (N_4845,N_3190,N_3049);
nor U4846 (N_4846,N_3390,N_3573);
or U4847 (N_4847,N_3615,N_3482);
nand U4848 (N_4848,N_3986,N_3696);
nor U4849 (N_4849,N_3049,N_3154);
xnor U4850 (N_4850,N_3730,N_3909);
or U4851 (N_4851,N_3976,N_3960);
nor U4852 (N_4852,N_3095,N_3647);
nand U4853 (N_4853,N_3375,N_3922);
xnor U4854 (N_4854,N_3340,N_3736);
or U4855 (N_4855,N_3054,N_3182);
nor U4856 (N_4856,N_3725,N_3765);
nor U4857 (N_4857,N_3791,N_3002);
or U4858 (N_4858,N_3509,N_3253);
and U4859 (N_4859,N_3757,N_3111);
and U4860 (N_4860,N_3303,N_3506);
or U4861 (N_4861,N_3666,N_3891);
xnor U4862 (N_4862,N_3925,N_3184);
nand U4863 (N_4863,N_3491,N_3682);
and U4864 (N_4864,N_3157,N_3103);
xor U4865 (N_4865,N_3707,N_3493);
xnor U4866 (N_4866,N_3588,N_3923);
nand U4867 (N_4867,N_3724,N_3240);
and U4868 (N_4868,N_3129,N_3622);
or U4869 (N_4869,N_3266,N_3463);
nand U4870 (N_4870,N_3118,N_3039);
and U4871 (N_4871,N_3850,N_3062);
nand U4872 (N_4872,N_3331,N_3515);
nor U4873 (N_4873,N_3288,N_3533);
nor U4874 (N_4874,N_3115,N_3682);
and U4875 (N_4875,N_3533,N_3294);
or U4876 (N_4876,N_3794,N_3382);
nor U4877 (N_4877,N_3488,N_3368);
or U4878 (N_4878,N_3113,N_3076);
and U4879 (N_4879,N_3031,N_3497);
xor U4880 (N_4880,N_3362,N_3561);
and U4881 (N_4881,N_3641,N_3504);
and U4882 (N_4882,N_3868,N_3274);
nor U4883 (N_4883,N_3104,N_3495);
nand U4884 (N_4884,N_3943,N_3100);
and U4885 (N_4885,N_3824,N_3191);
and U4886 (N_4886,N_3302,N_3959);
nand U4887 (N_4887,N_3933,N_3487);
xor U4888 (N_4888,N_3916,N_3675);
and U4889 (N_4889,N_3689,N_3166);
xor U4890 (N_4890,N_3991,N_3667);
nand U4891 (N_4891,N_3987,N_3864);
xnor U4892 (N_4892,N_3237,N_3794);
nor U4893 (N_4893,N_3171,N_3492);
xnor U4894 (N_4894,N_3984,N_3283);
nor U4895 (N_4895,N_3932,N_3094);
nand U4896 (N_4896,N_3223,N_3224);
xor U4897 (N_4897,N_3109,N_3898);
and U4898 (N_4898,N_3992,N_3464);
nor U4899 (N_4899,N_3078,N_3357);
nor U4900 (N_4900,N_3690,N_3685);
or U4901 (N_4901,N_3035,N_3576);
xor U4902 (N_4902,N_3906,N_3368);
xor U4903 (N_4903,N_3981,N_3941);
nor U4904 (N_4904,N_3207,N_3180);
and U4905 (N_4905,N_3952,N_3375);
xnor U4906 (N_4906,N_3855,N_3880);
or U4907 (N_4907,N_3423,N_3235);
nand U4908 (N_4908,N_3805,N_3928);
nand U4909 (N_4909,N_3443,N_3584);
or U4910 (N_4910,N_3877,N_3445);
xnor U4911 (N_4911,N_3266,N_3387);
nand U4912 (N_4912,N_3271,N_3594);
xnor U4913 (N_4913,N_3098,N_3786);
and U4914 (N_4914,N_3622,N_3056);
or U4915 (N_4915,N_3646,N_3954);
nand U4916 (N_4916,N_3606,N_3551);
and U4917 (N_4917,N_3273,N_3023);
or U4918 (N_4918,N_3970,N_3511);
and U4919 (N_4919,N_3946,N_3775);
xor U4920 (N_4920,N_3704,N_3291);
or U4921 (N_4921,N_3295,N_3801);
and U4922 (N_4922,N_3695,N_3314);
or U4923 (N_4923,N_3126,N_3083);
or U4924 (N_4924,N_3110,N_3931);
nand U4925 (N_4925,N_3352,N_3155);
or U4926 (N_4926,N_3711,N_3060);
and U4927 (N_4927,N_3101,N_3171);
and U4928 (N_4928,N_3548,N_3826);
and U4929 (N_4929,N_3749,N_3595);
nor U4930 (N_4930,N_3402,N_3627);
xnor U4931 (N_4931,N_3608,N_3754);
or U4932 (N_4932,N_3745,N_3088);
and U4933 (N_4933,N_3662,N_3096);
and U4934 (N_4934,N_3747,N_3776);
nor U4935 (N_4935,N_3807,N_3635);
nand U4936 (N_4936,N_3789,N_3426);
and U4937 (N_4937,N_3372,N_3162);
or U4938 (N_4938,N_3481,N_3886);
and U4939 (N_4939,N_3320,N_3512);
nand U4940 (N_4940,N_3729,N_3415);
nor U4941 (N_4941,N_3705,N_3781);
and U4942 (N_4942,N_3312,N_3599);
nor U4943 (N_4943,N_3010,N_3420);
xnor U4944 (N_4944,N_3179,N_3873);
and U4945 (N_4945,N_3977,N_3299);
nor U4946 (N_4946,N_3340,N_3812);
nand U4947 (N_4947,N_3134,N_3249);
and U4948 (N_4948,N_3242,N_3005);
xor U4949 (N_4949,N_3940,N_3941);
nor U4950 (N_4950,N_3518,N_3736);
or U4951 (N_4951,N_3089,N_3977);
or U4952 (N_4952,N_3156,N_3767);
nand U4953 (N_4953,N_3470,N_3429);
nor U4954 (N_4954,N_3709,N_3627);
and U4955 (N_4955,N_3817,N_3208);
nand U4956 (N_4956,N_3647,N_3770);
xor U4957 (N_4957,N_3553,N_3502);
or U4958 (N_4958,N_3088,N_3773);
nor U4959 (N_4959,N_3464,N_3583);
or U4960 (N_4960,N_3241,N_3424);
xnor U4961 (N_4961,N_3377,N_3209);
or U4962 (N_4962,N_3263,N_3615);
xnor U4963 (N_4963,N_3637,N_3754);
nand U4964 (N_4964,N_3670,N_3627);
xnor U4965 (N_4965,N_3853,N_3101);
nor U4966 (N_4966,N_3038,N_3581);
and U4967 (N_4967,N_3505,N_3415);
and U4968 (N_4968,N_3869,N_3823);
and U4969 (N_4969,N_3557,N_3912);
or U4970 (N_4970,N_3838,N_3167);
nor U4971 (N_4971,N_3928,N_3715);
and U4972 (N_4972,N_3867,N_3537);
and U4973 (N_4973,N_3901,N_3001);
nand U4974 (N_4974,N_3518,N_3122);
nor U4975 (N_4975,N_3399,N_3822);
xor U4976 (N_4976,N_3785,N_3165);
nor U4977 (N_4977,N_3063,N_3504);
xnor U4978 (N_4978,N_3477,N_3338);
nor U4979 (N_4979,N_3311,N_3808);
nand U4980 (N_4980,N_3531,N_3718);
xor U4981 (N_4981,N_3573,N_3579);
and U4982 (N_4982,N_3629,N_3498);
nor U4983 (N_4983,N_3350,N_3141);
nor U4984 (N_4984,N_3995,N_3608);
nor U4985 (N_4985,N_3706,N_3533);
or U4986 (N_4986,N_3867,N_3116);
nand U4987 (N_4987,N_3791,N_3748);
or U4988 (N_4988,N_3428,N_3946);
xor U4989 (N_4989,N_3378,N_3897);
xor U4990 (N_4990,N_3267,N_3172);
and U4991 (N_4991,N_3975,N_3683);
nor U4992 (N_4992,N_3726,N_3817);
nand U4993 (N_4993,N_3648,N_3735);
and U4994 (N_4994,N_3958,N_3760);
nor U4995 (N_4995,N_3280,N_3438);
nand U4996 (N_4996,N_3445,N_3853);
nor U4997 (N_4997,N_3762,N_3664);
nor U4998 (N_4998,N_3338,N_3405);
nand U4999 (N_4999,N_3147,N_3020);
xnor U5000 (N_5000,N_4436,N_4100);
or U5001 (N_5001,N_4619,N_4646);
or U5002 (N_5002,N_4584,N_4187);
or U5003 (N_5003,N_4770,N_4676);
xor U5004 (N_5004,N_4505,N_4501);
nor U5005 (N_5005,N_4420,N_4617);
nor U5006 (N_5006,N_4635,N_4106);
nand U5007 (N_5007,N_4230,N_4224);
nor U5008 (N_5008,N_4331,N_4042);
nand U5009 (N_5009,N_4081,N_4632);
and U5010 (N_5010,N_4105,N_4320);
or U5011 (N_5011,N_4589,N_4748);
or U5012 (N_5012,N_4246,N_4416);
nor U5013 (N_5013,N_4259,N_4338);
nor U5014 (N_5014,N_4704,N_4243);
and U5015 (N_5015,N_4705,N_4842);
or U5016 (N_5016,N_4247,N_4747);
nor U5017 (N_5017,N_4857,N_4658);
nor U5018 (N_5018,N_4924,N_4917);
and U5019 (N_5019,N_4793,N_4322);
xor U5020 (N_5020,N_4387,N_4863);
nor U5021 (N_5021,N_4626,N_4598);
or U5022 (N_5022,N_4260,N_4935);
or U5023 (N_5023,N_4755,N_4452);
xnor U5024 (N_5024,N_4385,N_4319);
xor U5025 (N_5025,N_4353,N_4869);
xnor U5026 (N_5026,N_4440,N_4342);
xnor U5027 (N_5027,N_4184,N_4064);
or U5028 (N_5028,N_4098,N_4824);
nor U5029 (N_5029,N_4914,N_4061);
nand U5030 (N_5030,N_4075,N_4957);
xor U5031 (N_5031,N_4998,N_4838);
or U5032 (N_5032,N_4923,N_4275);
xnor U5033 (N_5033,N_4860,N_4744);
or U5034 (N_5034,N_4932,N_4110);
xor U5035 (N_5035,N_4989,N_4997);
nor U5036 (N_5036,N_4473,N_4135);
nand U5037 (N_5037,N_4879,N_4126);
xor U5038 (N_5038,N_4897,N_4763);
nor U5039 (N_5039,N_4163,N_4173);
or U5040 (N_5040,N_4131,N_4905);
nor U5041 (N_5041,N_4774,N_4432);
nand U5042 (N_5042,N_4345,N_4688);
nand U5043 (N_5043,N_4987,N_4739);
or U5044 (N_5044,N_4164,N_4036);
xor U5045 (N_5045,N_4511,N_4941);
and U5046 (N_5046,N_4426,N_4295);
or U5047 (N_5047,N_4868,N_4616);
xor U5048 (N_5048,N_4800,N_4401);
and U5049 (N_5049,N_4825,N_4277);
or U5050 (N_5050,N_4487,N_4778);
or U5051 (N_5051,N_4009,N_4422);
nor U5052 (N_5052,N_4768,N_4291);
xnor U5053 (N_5053,N_4805,N_4303);
nand U5054 (N_5054,N_4643,N_4142);
and U5055 (N_5055,N_4798,N_4433);
nand U5056 (N_5056,N_4389,N_4166);
or U5057 (N_5057,N_4085,N_4468);
or U5058 (N_5058,N_4380,N_4047);
nor U5059 (N_5059,N_4955,N_4076);
or U5060 (N_5060,N_4661,N_4618);
or U5061 (N_5061,N_4783,N_4527);
nand U5062 (N_5062,N_4453,N_4831);
nand U5063 (N_5063,N_4614,N_4734);
and U5064 (N_5064,N_4370,N_4197);
nor U5065 (N_5065,N_4114,N_4776);
and U5066 (N_5066,N_4912,N_4031);
nor U5067 (N_5067,N_4760,N_4637);
or U5068 (N_5068,N_4486,N_4060);
or U5069 (N_5069,N_4535,N_4881);
and U5070 (N_5070,N_4025,N_4300);
xor U5071 (N_5071,N_4520,N_4029);
and U5072 (N_5072,N_4145,N_4648);
xnor U5073 (N_5073,N_4876,N_4754);
xor U5074 (N_5074,N_4927,N_4143);
nor U5075 (N_5075,N_4507,N_4671);
nor U5076 (N_5076,N_4310,N_4628);
or U5077 (N_5077,N_4968,N_4410);
nand U5078 (N_5078,N_4896,N_4457);
nand U5079 (N_5079,N_4082,N_4785);
and U5080 (N_5080,N_4948,N_4070);
nor U5081 (N_5081,N_4156,N_4318);
nor U5082 (N_5082,N_4299,N_4728);
nor U5083 (N_5083,N_4232,N_4451);
or U5084 (N_5084,N_4610,N_4483);
nand U5085 (N_5085,N_4152,N_4974);
or U5086 (N_5086,N_4804,N_4821);
and U5087 (N_5087,N_4874,N_4133);
nand U5088 (N_5088,N_4194,N_4008);
xnor U5089 (N_5089,N_4059,N_4687);
or U5090 (N_5090,N_4490,N_4719);
nor U5091 (N_5091,N_4978,N_4922);
xnor U5092 (N_5092,N_4642,N_4995);
or U5093 (N_5093,N_4192,N_4561);
nor U5094 (N_5094,N_4673,N_4052);
and U5095 (N_5095,N_4634,N_4523);
nor U5096 (N_5096,N_4678,N_4534);
nor U5097 (N_5097,N_4383,N_4976);
or U5098 (N_5098,N_4962,N_4878);
xnor U5099 (N_5099,N_4652,N_4888);
and U5100 (N_5100,N_4716,N_4111);
nor U5101 (N_5101,N_4693,N_4204);
xnor U5102 (N_5102,N_4553,N_4738);
nor U5103 (N_5103,N_4298,N_4791);
or U5104 (N_5104,N_4159,N_4725);
nand U5105 (N_5105,N_4240,N_4549);
nand U5106 (N_5106,N_4253,N_4139);
or U5107 (N_5107,N_4597,N_4560);
xnor U5108 (N_5108,N_4789,N_4216);
or U5109 (N_5109,N_4373,N_4663);
or U5110 (N_5110,N_4855,N_4093);
or U5111 (N_5111,N_4758,N_4582);
nand U5112 (N_5112,N_4586,N_4362);
and U5113 (N_5113,N_4516,N_4810);
xnor U5114 (N_5114,N_4478,N_4311);
or U5115 (N_5115,N_4335,N_4454);
nor U5116 (N_5116,N_4528,N_4116);
xnor U5117 (N_5117,N_4577,N_4474);
or U5118 (N_5118,N_4154,N_4852);
xnor U5119 (N_5119,N_4390,N_4118);
xnor U5120 (N_5120,N_4236,N_4206);
nor U5121 (N_5121,N_4500,N_4127);
nor U5122 (N_5122,N_4826,N_4980);
and U5123 (N_5123,N_4558,N_4262);
nor U5124 (N_5124,N_4727,N_4792);
or U5125 (N_5125,N_4048,N_4695);
nand U5126 (N_5126,N_4063,N_4956);
nand U5127 (N_5127,N_4714,N_4257);
and U5128 (N_5128,N_4899,N_4833);
nor U5129 (N_5129,N_4394,N_4669);
and U5130 (N_5130,N_4199,N_4344);
and U5131 (N_5131,N_4965,N_4429);
xor U5132 (N_5132,N_4065,N_4496);
xnor U5133 (N_5133,N_4428,N_4330);
xnor U5134 (N_5134,N_4732,N_4514);
nand U5135 (N_5135,N_4808,N_4324);
and U5136 (N_5136,N_4321,N_4435);
and U5137 (N_5137,N_4461,N_4827);
or U5138 (N_5138,N_4019,N_4759);
nor U5139 (N_5139,N_4668,N_4749);
nand U5140 (N_5140,N_4954,N_4532);
xor U5141 (N_5141,N_4915,N_4971);
and U5142 (N_5142,N_4209,N_4254);
nand U5143 (N_5143,N_4228,N_4062);
xnor U5144 (N_5144,N_4032,N_4049);
nor U5145 (N_5145,N_4581,N_4023);
or U5146 (N_5146,N_4456,N_4449);
or U5147 (N_5147,N_4506,N_4641);
nand U5148 (N_5148,N_4423,N_4392);
and U5149 (N_5149,N_4653,N_4724);
nand U5150 (N_5150,N_4891,N_4702);
nor U5151 (N_5151,N_4201,N_4984);
xor U5152 (N_5152,N_4949,N_4574);
or U5153 (N_5153,N_4633,N_4745);
nor U5154 (N_5154,N_4186,N_4684);
and U5155 (N_5155,N_4638,N_4587);
or U5156 (N_5156,N_4710,N_4006);
nand U5157 (N_5157,N_4363,N_4237);
nor U5158 (N_5158,N_4404,N_4244);
or U5159 (N_5159,N_4165,N_4280);
or U5160 (N_5160,N_4567,N_4990);
and U5161 (N_5161,N_4227,N_4659);
or U5162 (N_5162,N_4347,N_4301);
xnor U5163 (N_5163,N_4753,N_4447);
and U5164 (N_5164,N_4285,N_4811);
and U5165 (N_5165,N_4884,N_4323);
nand U5166 (N_5166,N_4602,N_4182);
nand U5167 (N_5167,N_4475,N_4408);
nand U5168 (N_5168,N_4424,N_4736);
nand U5169 (N_5169,N_4266,N_4906);
nand U5170 (N_5170,N_4179,N_4109);
nand U5171 (N_5171,N_4485,N_4212);
nand U5172 (N_5172,N_4622,N_4557);
and U5173 (N_5173,N_4667,N_4446);
xnor U5174 (N_5174,N_4095,N_4292);
or U5175 (N_5175,N_4469,N_4596);
and U5176 (N_5176,N_4620,N_4541);
and U5177 (N_5177,N_4830,N_4007);
nand U5178 (N_5178,N_4928,N_4544);
or U5179 (N_5179,N_4942,N_4217);
xnor U5180 (N_5180,N_4326,N_4657);
and U5181 (N_5181,N_4252,N_4701);
or U5182 (N_5182,N_4125,N_4645);
or U5183 (N_5183,N_4074,N_4866);
or U5184 (N_5184,N_4819,N_4037);
xor U5185 (N_5185,N_4024,N_4802);
nand U5186 (N_5186,N_4806,N_4307);
and U5187 (N_5187,N_4411,N_4122);
nand U5188 (N_5188,N_4913,N_4950);
nor U5189 (N_5189,N_4388,N_4066);
nor U5190 (N_5190,N_4531,N_4418);
nand U5191 (N_5191,N_4592,N_4480);
or U5192 (N_5192,N_4828,N_4892);
xnor U5193 (N_5193,N_4926,N_4621);
nand U5194 (N_5194,N_4844,N_4349);
and U5195 (N_5195,N_4441,N_4375);
or U5196 (N_5196,N_4296,N_4117);
nand U5197 (N_5197,N_4611,N_4103);
and U5198 (N_5198,N_4222,N_4593);
and U5199 (N_5199,N_4940,N_4921);
or U5200 (N_5200,N_4107,N_4071);
xnor U5201 (N_5201,N_4113,N_4251);
nand U5202 (N_5202,N_4672,N_4067);
nor U5203 (N_5203,N_4434,N_4386);
or U5204 (N_5204,N_4439,N_4289);
xor U5205 (N_5205,N_4911,N_4859);
nand U5206 (N_5206,N_4903,N_4689);
and U5207 (N_5207,N_4700,N_4934);
nand U5208 (N_5208,N_4033,N_4276);
xnor U5209 (N_5209,N_4554,N_4279);
nand U5210 (N_5210,N_4972,N_4088);
nor U5211 (N_5211,N_4482,N_4578);
nand U5212 (N_5212,N_4885,N_4011);
xnor U5213 (N_5213,N_4699,N_4900);
or U5214 (N_5214,N_4283,N_4352);
or U5215 (N_5215,N_4250,N_4120);
nand U5216 (N_5216,N_4001,N_4479);
xnor U5217 (N_5217,N_4901,N_4396);
nand U5218 (N_5218,N_4051,N_4214);
and U5219 (N_5219,N_4234,N_4650);
xor U5220 (N_5220,N_4101,N_4910);
or U5221 (N_5221,N_4431,N_4613);
and U5222 (N_5222,N_4889,N_4493);
or U5223 (N_5223,N_4945,N_4499);
xnor U5224 (N_5224,N_4312,N_4545);
xor U5225 (N_5225,N_4639,N_4814);
nand U5226 (N_5226,N_4988,N_4951);
or U5227 (N_5227,N_4415,N_4281);
nand U5228 (N_5228,N_4662,N_4834);
nor U5229 (N_5229,N_4382,N_4438);
nand U5230 (N_5230,N_4952,N_4104);
and U5231 (N_5231,N_4600,N_4686);
nor U5232 (N_5232,N_4590,N_4448);
or U5233 (N_5233,N_4495,N_4297);
xnor U5234 (N_5234,N_4078,N_4681);
xnor U5235 (N_5235,N_4265,N_4369);
nand U5236 (N_5236,N_4517,N_4332);
xnor U5237 (N_5237,N_4378,N_4459);
xnor U5238 (N_5238,N_4132,N_4012);
nand U5239 (N_5239,N_4670,N_4162);
nor U5240 (N_5240,N_4605,N_4835);
or U5241 (N_5241,N_4210,N_4542);
xor U5242 (N_5242,N_4039,N_4666);
xor U5243 (N_5243,N_4178,N_4731);
or U5244 (N_5244,N_4102,N_4513);
or U5245 (N_5245,N_4822,N_4185);
xor U5246 (N_5246,N_4969,N_4358);
or U5247 (N_5247,N_4221,N_4851);
or U5248 (N_5248,N_4895,N_4930);
or U5249 (N_5249,N_4729,N_4953);
and U5250 (N_5250,N_4966,N_4005);
xor U5251 (N_5251,N_4723,N_4003);
nand U5252 (N_5252,N_4556,N_4317);
and U5253 (N_5253,N_4769,N_4366);
or U5254 (N_5254,N_4034,N_4014);
or U5255 (N_5255,N_4263,N_4177);
and U5256 (N_5256,N_4845,N_4053);
nor U5257 (N_5257,N_4815,N_4521);
and U5258 (N_5258,N_4069,N_4720);
nand U5259 (N_5259,N_4525,N_4027);
or U5260 (N_5260,N_4817,N_4916);
nor U5261 (N_5261,N_4991,N_4624);
and U5262 (N_5262,N_4981,N_4837);
nor U5263 (N_5263,N_4271,N_4421);
or U5264 (N_5264,N_4537,N_4765);
nand U5265 (N_5265,N_4208,N_4020);
nor U5266 (N_5266,N_4302,N_4004);
xnor U5267 (N_5267,N_4947,N_4999);
nand U5268 (N_5268,N_4882,N_4211);
and U5269 (N_5269,N_4625,N_4591);
or U5270 (N_5270,N_4337,N_4570);
xor U5271 (N_5271,N_4403,N_4180);
nor U5272 (N_5272,N_4092,N_4807);
xnor U5273 (N_5273,N_4213,N_4551);
and U5274 (N_5274,N_4255,N_4138);
and U5275 (N_5275,N_4465,N_4498);
and U5276 (N_5276,N_4929,N_4346);
xor U5277 (N_5277,N_4356,N_4750);
nor U5278 (N_5278,N_4887,N_4226);
nand U5279 (N_5279,N_4640,N_4683);
and U5280 (N_5280,N_4399,N_4801);
nor U5281 (N_5281,N_4249,N_4413);
xor U5282 (N_5282,N_4559,N_4711);
xnor U5283 (N_5283,N_4707,N_4994);
nor U5284 (N_5284,N_4795,N_4872);
nand U5285 (N_5285,N_4464,N_4141);
nor U5286 (N_5286,N_4809,N_4115);
xor U5287 (N_5287,N_4733,N_4274);
or U5288 (N_5288,N_4608,N_4647);
nor U5289 (N_5289,N_4040,N_4269);
or U5290 (N_5290,N_4463,N_4044);
and U5291 (N_5291,N_4158,N_4609);
nand U5292 (N_5292,N_4364,N_4151);
nor U5293 (N_5293,N_4973,N_4588);
xnor U5294 (N_5294,N_4936,N_4130);
xor U5295 (N_5295,N_4547,N_4960);
and U5296 (N_5296,N_4144,N_4533);
and U5297 (N_5297,N_4000,N_4354);
and U5298 (N_5298,N_4050,N_4183);
nand U5299 (N_5299,N_4746,N_4938);
nand U5300 (N_5300,N_4627,N_4536);
nor U5301 (N_5301,N_4694,N_4843);
and U5302 (N_5302,N_4171,N_4235);
nand U5303 (N_5303,N_4030,N_4775);
or U5304 (N_5304,N_4944,N_4565);
or U5305 (N_5305,N_4623,N_4489);
nand U5306 (N_5306,N_4503,N_4864);
xor U5307 (N_5307,N_4195,N_4594);
or U5308 (N_5308,N_4518,N_4631);
and U5309 (N_5309,N_4709,N_4391);
nor U5310 (N_5310,N_4002,N_4796);
or U5311 (N_5311,N_4225,N_4893);
and U5312 (N_5312,N_4696,N_4170);
or U5313 (N_5313,N_4357,N_4146);
nand U5314 (N_5314,N_4055,N_4191);
nand U5315 (N_5315,N_4787,N_4982);
xor U5316 (N_5316,N_4543,N_4979);
xnor U5317 (N_5317,N_4284,N_4016);
nand U5318 (N_5318,N_4963,N_4540);
and U5319 (N_5319,N_4022,N_4522);
xor U5320 (N_5320,N_4339,N_4782);
or U5321 (N_5321,N_4674,N_4583);
or U5322 (N_5322,N_4038,N_4476);
nand U5323 (N_5323,N_4248,N_4360);
or U5324 (N_5324,N_4494,N_4443);
nand U5325 (N_5325,N_4664,N_4290);
nand U5326 (N_5326,N_4245,N_4772);
or U5327 (N_5327,N_4898,N_4309);
xor U5328 (N_5328,N_4137,N_4797);
or U5329 (N_5329,N_4526,N_4757);
nand U5330 (N_5330,N_4412,N_4351);
xnor U5331 (N_5331,N_4196,N_4068);
or U5332 (N_5332,N_4155,N_4172);
xor U5333 (N_5333,N_4477,N_4649);
or U5334 (N_5334,N_4207,N_4794);
nand U5335 (N_5335,N_4579,N_4367);
or U5336 (N_5336,N_4256,N_4466);
and U5337 (N_5337,N_4530,N_4961);
nand U5338 (N_5338,N_4123,N_4181);
or U5339 (N_5339,N_4333,N_4829);
nand U5340 (N_5340,N_4568,N_4730);
xnor U5341 (N_5341,N_4455,N_4943);
nand U5342 (N_5342,N_4058,N_4328);
nor U5343 (N_5343,N_4350,N_4374);
and U5344 (N_5344,N_4871,N_4629);
xnor U5345 (N_5345,N_4713,N_4381);
or U5346 (N_5346,N_4169,N_4508);
or U5347 (N_5347,N_4336,N_4268);
nor U5348 (N_5348,N_4931,N_4119);
and U5349 (N_5349,N_4959,N_4136);
nor U5350 (N_5350,N_4121,N_4737);
nor U5351 (N_5351,N_4975,N_4045);
or U5352 (N_5352,N_4112,N_4445);
or U5353 (N_5353,N_4902,N_4604);
xor U5354 (N_5354,N_4203,N_4128);
nor U5355 (N_5355,N_4089,N_4218);
nor U5356 (N_5356,N_4017,N_4108);
or U5357 (N_5357,N_4293,N_4419);
and U5358 (N_5358,N_4865,N_4220);
xnor U5359 (N_5359,N_4886,N_4046);
nor U5360 (N_5360,N_4083,N_4086);
xor U5361 (N_5361,N_4504,N_4867);
xor U5362 (N_5362,N_4174,N_4812);
xnor U5363 (N_5363,N_4712,N_4028);
and U5364 (N_5364,N_4890,N_4189);
xor U5365 (N_5365,N_4484,N_4918);
xor U5366 (N_5366,N_4550,N_4147);
or U5367 (N_5367,N_4097,N_4680);
nand U5368 (N_5368,N_4264,N_4985);
nand U5369 (N_5369,N_4883,N_4706);
nand U5370 (N_5370,N_4781,N_4188);
and U5371 (N_5371,N_4278,N_4134);
or U5372 (N_5372,N_4467,N_4355);
or U5373 (N_5373,N_4964,N_4690);
xnor U5374 (N_5374,N_4790,N_4018);
nor U5375 (N_5375,N_4261,N_4677);
or U5376 (N_5376,N_4546,N_4481);
nor U5377 (N_5377,N_4698,N_4992);
or U5378 (N_5378,N_4771,N_4427);
and U5379 (N_5379,N_4569,N_4233);
nand U5380 (N_5380,N_4340,N_4200);
nor U5381 (N_5381,N_4304,N_4853);
and U5382 (N_5382,N_4215,N_4472);
nor U5383 (N_5383,N_4091,N_4970);
nor U5384 (N_5384,N_4512,N_4015);
nand U5385 (N_5385,N_4073,N_4741);
nor U5386 (N_5386,N_4470,N_4656);
nand U5387 (N_5387,N_4909,N_4908);
xnor U5388 (N_5388,N_4555,N_4442);
xor U5389 (N_5389,N_4873,N_4272);
or U5390 (N_5390,N_4847,N_4870);
or U5391 (N_5391,N_4717,N_4703);
or U5392 (N_5392,N_4742,N_4041);
nor U5393 (N_5393,N_4223,N_4846);
nor U5394 (N_5394,N_4376,N_4715);
nor U5395 (N_5395,N_4818,N_4329);
nand U5396 (N_5396,N_4398,N_4856);
xor U5397 (N_5397,N_4365,N_4832);
nor U5398 (N_5398,N_4722,N_4087);
and U5399 (N_5399,N_4840,N_4316);
nor U5400 (N_5400,N_4599,N_4773);
xnor U5401 (N_5401,N_4849,N_4359);
and U5402 (N_5402,N_4761,N_4056);
nand U5403 (N_5403,N_4993,N_4751);
and U5404 (N_5404,N_4270,N_4239);
and U5405 (N_5405,N_4996,N_4655);
nand U5406 (N_5406,N_4444,N_4026);
or U5407 (N_5407,N_4334,N_4077);
or U5408 (N_5408,N_4096,N_4841);
nand U5409 (N_5409,N_4572,N_4820);
and U5410 (N_5410,N_4651,N_4219);
nor U5411 (N_5411,N_4348,N_4777);
and U5412 (N_5412,N_4630,N_4202);
and U5413 (N_5413,N_4509,N_4850);
and U5414 (N_5414,N_4665,N_4607);
xor U5415 (N_5415,N_4090,N_4858);
and U5416 (N_5416,N_4361,N_4967);
nor U5417 (N_5417,N_4437,N_4904);
nor U5418 (N_5418,N_4764,N_4035);
nand U5419 (N_5419,N_4417,N_4176);
xor U5420 (N_5420,N_4958,N_4153);
or U5421 (N_5421,N_4368,N_4685);
nor U5422 (N_5422,N_4595,N_4099);
nand U5423 (N_5423,N_4384,N_4571);
and U5424 (N_5424,N_4371,N_4407);
and U5425 (N_5425,N_4784,N_4314);
nand U5426 (N_5426,N_4393,N_4460);
nand U5427 (N_5427,N_4562,N_4679);
and U5428 (N_5428,N_4799,N_4405);
or U5429 (N_5429,N_4636,N_4175);
and U5430 (N_5430,N_4861,N_4450);
nor U5431 (N_5431,N_4735,N_4552);
and U5432 (N_5432,N_4372,N_4767);
nand U5433 (N_5433,N_4538,N_4124);
or U5434 (N_5434,N_4379,N_4524);
or U5435 (N_5435,N_4306,N_4925);
nor U5436 (N_5436,N_4462,N_4894);
nand U5437 (N_5437,N_4242,N_4157);
or U5438 (N_5438,N_4043,N_4190);
nor U5439 (N_5439,N_4519,N_4205);
and U5440 (N_5440,N_4308,N_4919);
and U5441 (N_5441,N_4875,N_4288);
nand U5442 (N_5442,N_4497,N_4697);
or U5443 (N_5443,N_4341,N_4539);
nor U5444 (N_5444,N_4488,N_4612);
or U5445 (N_5445,N_4548,N_4325);
or U5446 (N_5446,N_4149,N_4400);
xor U5447 (N_5447,N_4691,N_4231);
nand U5448 (N_5448,N_4079,N_4939);
or U5449 (N_5449,N_4766,N_4395);
and U5450 (N_5450,N_4836,N_4933);
nor U5451 (N_5451,N_4946,N_4343);
nor U5452 (N_5452,N_4743,N_4327);
xnor U5453 (N_5453,N_4229,N_4726);
nor U5454 (N_5454,N_4094,N_4057);
xor U5455 (N_5455,N_4072,N_4129);
or U5456 (N_5456,N_4080,N_4021);
and U5457 (N_5457,N_4193,N_4839);
and U5458 (N_5458,N_4780,N_4756);
nand U5459 (N_5459,N_4406,N_4425);
xor U5460 (N_5460,N_4294,N_4813);
nor U5461 (N_5461,N_4258,N_4397);
and U5462 (N_5462,N_4377,N_4282);
nor U5463 (N_5463,N_4471,N_4267);
xnor U5464 (N_5464,N_4660,N_4084);
xnor U5465 (N_5465,N_4977,N_4167);
and U5466 (N_5466,N_4601,N_4675);
and U5467 (N_5467,N_4013,N_4937);
nand U5468 (N_5468,N_4148,N_4907);
xnor U5469 (N_5469,N_4580,N_4315);
and U5470 (N_5470,N_4803,N_4502);
and U5471 (N_5471,N_4161,N_4752);
nand U5472 (N_5472,N_4273,N_4786);
nor U5473 (N_5473,N_4564,N_4877);
and U5474 (N_5474,N_4576,N_4862);
or U5475 (N_5475,N_4241,N_4606);
nand U5476 (N_5476,N_4603,N_4563);
nor U5477 (N_5477,N_4529,N_4654);
and U5478 (N_5478,N_4573,N_4168);
and U5479 (N_5479,N_4880,N_4615);
xor U5480 (N_5480,N_4823,N_4986);
and U5481 (N_5481,N_4788,N_4054);
or U5482 (N_5482,N_4150,N_4854);
nand U5483 (N_5483,N_4238,N_4160);
xor U5484 (N_5484,N_4920,N_4492);
and U5485 (N_5485,N_4692,N_4779);
nand U5486 (N_5486,N_4305,N_4140);
and U5487 (N_5487,N_4287,N_4198);
and U5488 (N_5488,N_4983,N_4313);
nand U5489 (N_5489,N_4402,N_4010);
or U5490 (N_5490,N_4682,N_4644);
or U5491 (N_5491,N_4414,N_4848);
nand U5492 (N_5492,N_4510,N_4430);
nand U5493 (N_5493,N_4718,N_4286);
or U5494 (N_5494,N_4566,N_4515);
nor U5495 (N_5495,N_4721,N_4816);
or U5496 (N_5496,N_4740,N_4491);
xor U5497 (N_5497,N_4409,N_4708);
nand U5498 (N_5498,N_4458,N_4585);
or U5499 (N_5499,N_4762,N_4575);
and U5500 (N_5500,N_4367,N_4043);
nor U5501 (N_5501,N_4804,N_4527);
and U5502 (N_5502,N_4109,N_4599);
nand U5503 (N_5503,N_4679,N_4425);
xor U5504 (N_5504,N_4881,N_4314);
and U5505 (N_5505,N_4958,N_4810);
nor U5506 (N_5506,N_4783,N_4538);
or U5507 (N_5507,N_4923,N_4682);
or U5508 (N_5508,N_4459,N_4274);
and U5509 (N_5509,N_4862,N_4442);
nor U5510 (N_5510,N_4888,N_4563);
and U5511 (N_5511,N_4843,N_4587);
nand U5512 (N_5512,N_4577,N_4345);
or U5513 (N_5513,N_4902,N_4421);
and U5514 (N_5514,N_4669,N_4860);
xor U5515 (N_5515,N_4317,N_4843);
xnor U5516 (N_5516,N_4122,N_4488);
or U5517 (N_5517,N_4375,N_4043);
nand U5518 (N_5518,N_4642,N_4421);
nand U5519 (N_5519,N_4849,N_4246);
nor U5520 (N_5520,N_4260,N_4563);
nand U5521 (N_5521,N_4012,N_4342);
xor U5522 (N_5522,N_4224,N_4326);
nor U5523 (N_5523,N_4064,N_4760);
xnor U5524 (N_5524,N_4743,N_4282);
and U5525 (N_5525,N_4415,N_4150);
nor U5526 (N_5526,N_4341,N_4363);
or U5527 (N_5527,N_4051,N_4067);
nor U5528 (N_5528,N_4068,N_4617);
or U5529 (N_5529,N_4534,N_4406);
or U5530 (N_5530,N_4041,N_4294);
and U5531 (N_5531,N_4389,N_4143);
xor U5532 (N_5532,N_4761,N_4499);
nor U5533 (N_5533,N_4602,N_4305);
and U5534 (N_5534,N_4275,N_4781);
xnor U5535 (N_5535,N_4894,N_4957);
nor U5536 (N_5536,N_4634,N_4198);
and U5537 (N_5537,N_4138,N_4269);
nor U5538 (N_5538,N_4126,N_4353);
nand U5539 (N_5539,N_4340,N_4023);
xnor U5540 (N_5540,N_4264,N_4070);
xor U5541 (N_5541,N_4151,N_4532);
nor U5542 (N_5542,N_4883,N_4663);
nor U5543 (N_5543,N_4273,N_4990);
or U5544 (N_5544,N_4335,N_4318);
and U5545 (N_5545,N_4059,N_4914);
and U5546 (N_5546,N_4733,N_4986);
nand U5547 (N_5547,N_4845,N_4625);
nand U5548 (N_5548,N_4624,N_4460);
nand U5549 (N_5549,N_4004,N_4360);
or U5550 (N_5550,N_4524,N_4169);
nand U5551 (N_5551,N_4915,N_4197);
nand U5552 (N_5552,N_4895,N_4514);
and U5553 (N_5553,N_4034,N_4917);
or U5554 (N_5554,N_4835,N_4610);
or U5555 (N_5555,N_4471,N_4299);
and U5556 (N_5556,N_4822,N_4227);
nor U5557 (N_5557,N_4963,N_4340);
or U5558 (N_5558,N_4110,N_4458);
xnor U5559 (N_5559,N_4264,N_4749);
nor U5560 (N_5560,N_4047,N_4831);
or U5561 (N_5561,N_4910,N_4793);
xnor U5562 (N_5562,N_4660,N_4793);
nand U5563 (N_5563,N_4949,N_4120);
nand U5564 (N_5564,N_4247,N_4654);
or U5565 (N_5565,N_4799,N_4784);
or U5566 (N_5566,N_4696,N_4594);
and U5567 (N_5567,N_4837,N_4412);
nand U5568 (N_5568,N_4500,N_4576);
nand U5569 (N_5569,N_4014,N_4447);
nor U5570 (N_5570,N_4466,N_4144);
or U5571 (N_5571,N_4859,N_4850);
or U5572 (N_5572,N_4555,N_4086);
and U5573 (N_5573,N_4102,N_4256);
xnor U5574 (N_5574,N_4859,N_4890);
or U5575 (N_5575,N_4444,N_4887);
or U5576 (N_5576,N_4180,N_4836);
nor U5577 (N_5577,N_4405,N_4828);
xnor U5578 (N_5578,N_4682,N_4683);
nor U5579 (N_5579,N_4375,N_4145);
and U5580 (N_5580,N_4562,N_4293);
nand U5581 (N_5581,N_4320,N_4538);
or U5582 (N_5582,N_4028,N_4815);
xor U5583 (N_5583,N_4170,N_4506);
and U5584 (N_5584,N_4385,N_4399);
nor U5585 (N_5585,N_4949,N_4284);
or U5586 (N_5586,N_4110,N_4319);
xor U5587 (N_5587,N_4128,N_4463);
nand U5588 (N_5588,N_4012,N_4570);
nor U5589 (N_5589,N_4132,N_4293);
nor U5590 (N_5590,N_4465,N_4472);
or U5591 (N_5591,N_4474,N_4845);
nor U5592 (N_5592,N_4733,N_4923);
and U5593 (N_5593,N_4700,N_4751);
nor U5594 (N_5594,N_4563,N_4130);
and U5595 (N_5595,N_4081,N_4640);
xnor U5596 (N_5596,N_4022,N_4035);
xnor U5597 (N_5597,N_4557,N_4331);
xor U5598 (N_5598,N_4511,N_4710);
or U5599 (N_5599,N_4910,N_4116);
or U5600 (N_5600,N_4763,N_4982);
or U5601 (N_5601,N_4204,N_4927);
xnor U5602 (N_5602,N_4536,N_4006);
and U5603 (N_5603,N_4557,N_4987);
or U5604 (N_5604,N_4443,N_4959);
nand U5605 (N_5605,N_4573,N_4350);
nor U5606 (N_5606,N_4395,N_4626);
or U5607 (N_5607,N_4168,N_4141);
nand U5608 (N_5608,N_4452,N_4921);
and U5609 (N_5609,N_4882,N_4636);
nor U5610 (N_5610,N_4265,N_4358);
nor U5611 (N_5611,N_4948,N_4445);
nor U5612 (N_5612,N_4981,N_4136);
nand U5613 (N_5613,N_4556,N_4174);
or U5614 (N_5614,N_4830,N_4511);
nor U5615 (N_5615,N_4483,N_4798);
nor U5616 (N_5616,N_4345,N_4526);
nand U5617 (N_5617,N_4188,N_4003);
or U5618 (N_5618,N_4790,N_4376);
nor U5619 (N_5619,N_4525,N_4469);
and U5620 (N_5620,N_4331,N_4037);
nor U5621 (N_5621,N_4016,N_4287);
or U5622 (N_5622,N_4177,N_4210);
nor U5623 (N_5623,N_4832,N_4892);
or U5624 (N_5624,N_4710,N_4960);
nor U5625 (N_5625,N_4384,N_4718);
or U5626 (N_5626,N_4256,N_4206);
nand U5627 (N_5627,N_4136,N_4299);
xnor U5628 (N_5628,N_4856,N_4338);
or U5629 (N_5629,N_4243,N_4371);
nor U5630 (N_5630,N_4578,N_4828);
or U5631 (N_5631,N_4724,N_4435);
or U5632 (N_5632,N_4999,N_4256);
and U5633 (N_5633,N_4193,N_4342);
nor U5634 (N_5634,N_4581,N_4032);
and U5635 (N_5635,N_4311,N_4166);
or U5636 (N_5636,N_4334,N_4771);
nor U5637 (N_5637,N_4346,N_4557);
nand U5638 (N_5638,N_4368,N_4778);
or U5639 (N_5639,N_4305,N_4748);
xor U5640 (N_5640,N_4465,N_4936);
nand U5641 (N_5641,N_4470,N_4611);
xor U5642 (N_5642,N_4671,N_4281);
nand U5643 (N_5643,N_4438,N_4563);
and U5644 (N_5644,N_4171,N_4231);
nor U5645 (N_5645,N_4261,N_4864);
or U5646 (N_5646,N_4447,N_4585);
or U5647 (N_5647,N_4404,N_4064);
xor U5648 (N_5648,N_4809,N_4761);
or U5649 (N_5649,N_4590,N_4776);
and U5650 (N_5650,N_4518,N_4906);
nor U5651 (N_5651,N_4080,N_4388);
or U5652 (N_5652,N_4324,N_4515);
or U5653 (N_5653,N_4920,N_4336);
or U5654 (N_5654,N_4371,N_4181);
or U5655 (N_5655,N_4605,N_4921);
nand U5656 (N_5656,N_4060,N_4333);
nor U5657 (N_5657,N_4710,N_4895);
or U5658 (N_5658,N_4386,N_4505);
and U5659 (N_5659,N_4804,N_4321);
nand U5660 (N_5660,N_4244,N_4447);
or U5661 (N_5661,N_4291,N_4713);
nor U5662 (N_5662,N_4688,N_4800);
and U5663 (N_5663,N_4860,N_4153);
nor U5664 (N_5664,N_4465,N_4346);
nand U5665 (N_5665,N_4521,N_4867);
xor U5666 (N_5666,N_4873,N_4383);
or U5667 (N_5667,N_4167,N_4543);
nand U5668 (N_5668,N_4102,N_4344);
nor U5669 (N_5669,N_4516,N_4790);
nand U5670 (N_5670,N_4008,N_4588);
or U5671 (N_5671,N_4609,N_4799);
nor U5672 (N_5672,N_4002,N_4975);
or U5673 (N_5673,N_4957,N_4301);
nor U5674 (N_5674,N_4624,N_4311);
and U5675 (N_5675,N_4606,N_4419);
nand U5676 (N_5676,N_4303,N_4649);
nand U5677 (N_5677,N_4342,N_4575);
and U5678 (N_5678,N_4864,N_4644);
or U5679 (N_5679,N_4694,N_4385);
nor U5680 (N_5680,N_4848,N_4906);
and U5681 (N_5681,N_4968,N_4537);
and U5682 (N_5682,N_4244,N_4262);
nor U5683 (N_5683,N_4224,N_4208);
and U5684 (N_5684,N_4601,N_4038);
xnor U5685 (N_5685,N_4395,N_4179);
nor U5686 (N_5686,N_4764,N_4776);
or U5687 (N_5687,N_4094,N_4739);
xnor U5688 (N_5688,N_4112,N_4906);
nand U5689 (N_5689,N_4678,N_4473);
and U5690 (N_5690,N_4171,N_4775);
nand U5691 (N_5691,N_4760,N_4210);
nor U5692 (N_5692,N_4864,N_4975);
nor U5693 (N_5693,N_4213,N_4157);
xnor U5694 (N_5694,N_4512,N_4866);
nand U5695 (N_5695,N_4290,N_4568);
nor U5696 (N_5696,N_4230,N_4909);
xnor U5697 (N_5697,N_4678,N_4539);
nand U5698 (N_5698,N_4436,N_4851);
and U5699 (N_5699,N_4525,N_4171);
nor U5700 (N_5700,N_4812,N_4158);
nand U5701 (N_5701,N_4935,N_4181);
and U5702 (N_5702,N_4505,N_4876);
nand U5703 (N_5703,N_4288,N_4496);
and U5704 (N_5704,N_4406,N_4469);
or U5705 (N_5705,N_4683,N_4990);
xnor U5706 (N_5706,N_4966,N_4782);
nor U5707 (N_5707,N_4439,N_4344);
nand U5708 (N_5708,N_4177,N_4353);
nand U5709 (N_5709,N_4005,N_4084);
xor U5710 (N_5710,N_4036,N_4686);
or U5711 (N_5711,N_4565,N_4713);
xor U5712 (N_5712,N_4714,N_4882);
xor U5713 (N_5713,N_4969,N_4655);
or U5714 (N_5714,N_4581,N_4027);
xor U5715 (N_5715,N_4392,N_4050);
and U5716 (N_5716,N_4685,N_4402);
nand U5717 (N_5717,N_4648,N_4294);
and U5718 (N_5718,N_4928,N_4921);
or U5719 (N_5719,N_4509,N_4932);
and U5720 (N_5720,N_4781,N_4017);
nand U5721 (N_5721,N_4875,N_4447);
nor U5722 (N_5722,N_4989,N_4171);
or U5723 (N_5723,N_4867,N_4005);
nand U5724 (N_5724,N_4797,N_4891);
xnor U5725 (N_5725,N_4752,N_4334);
xnor U5726 (N_5726,N_4708,N_4377);
or U5727 (N_5727,N_4440,N_4999);
nor U5728 (N_5728,N_4302,N_4357);
and U5729 (N_5729,N_4043,N_4920);
nand U5730 (N_5730,N_4501,N_4091);
nor U5731 (N_5731,N_4291,N_4359);
nor U5732 (N_5732,N_4910,N_4920);
nand U5733 (N_5733,N_4700,N_4828);
or U5734 (N_5734,N_4176,N_4054);
and U5735 (N_5735,N_4207,N_4183);
or U5736 (N_5736,N_4595,N_4327);
nand U5737 (N_5737,N_4060,N_4356);
nand U5738 (N_5738,N_4555,N_4164);
or U5739 (N_5739,N_4859,N_4403);
xnor U5740 (N_5740,N_4892,N_4315);
or U5741 (N_5741,N_4258,N_4190);
and U5742 (N_5742,N_4911,N_4714);
xnor U5743 (N_5743,N_4254,N_4585);
and U5744 (N_5744,N_4816,N_4197);
nor U5745 (N_5745,N_4791,N_4131);
and U5746 (N_5746,N_4613,N_4753);
or U5747 (N_5747,N_4340,N_4639);
or U5748 (N_5748,N_4166,N_4445);
xnor U5749 (N_5749,N_4911,N_4201);
and U5750 (N_5750,N_4814,N_4448);
and U5751 (N_5751,N_4047,N_4852);
nor U5752 (N_5752,N_4290,N_4518);
nor U5753 (N_5753,N_4025,N_4516);
or U5754 (N_5754,N_4855,N_4161);
and U5755 (N_5755,N_4981,N_4552);
nor U5756 (N_5756,N_4777,N_4940);
nand U5757 (N_5757,N_4516,N_4819);
or U5758 (N_5758,N_4238,N_4298);
nand U5759 (N_5759,N_4620,N_4964);
or U5760 (N_5760,N_4194,N_4150);
or U5761 (N_5761,N_4175,N_4566);
nor U5762 (N_5762,N_4158,N_4391);
xnor U5763 (N_5763,N_4412,N_4029);
xnor U5764 (N_5764,N_4074,N_4062);
nand U5765 (N_5765,N_4976,N_4404);
nand U5766 (N_5766,N_4182,N_4388);
or U5767 (N_5767,N_4846,N_4606);
nor U5768 (N_5768,N_4900,N_4169);
or U5769 (N_5769,N_4607,N_4263);
xnor U5770 (N_5770,N_4922,N_4203);
and U5771 (N_5771,N_4964,N_4286);
and U5772 (N_5772,N_4071,N_4633);
xnor U5773 (N_5773,N_4190,N_4361);
or U5774 (N_5774,N_4494,N_4122);
nand U5775 (N_5775,N_4311,N_4458);
nand U5776 (N_5776,N_4371,N_4012);
and U5777 (N_5777,N_4286,N_4735);
nand U5778 (N_5778,N_4361,N_4657);
nand U5779 (N_5779,N_4460,N_4607);
nor U5780 (N_5780,N_4332,N_4537);
nor U5781 (N_5781,N_4053,N_4847);
xor U5782 (N_5782,N_4587,N_4556);
xor U5783 (N_5783,N_4995,N_4549);
and U5784 (N_5784,N_4397,N_4125);
nand U5785 (N_5785,N_4057,N_4966);
and U5786 (N_5786,N_4015,N_4906);
or U5787 (N_5787,N_4948,N_4801);
nand U5788 (N_5788,N_4169,N_4252);
or U5789 (N_5789,N_4693,N_4373);
or U5790 (N_5790,N_4102,N_4689);
and U5791 (N_5791,N_4028,N_4575);
or U5792 (N_5792,N_4354,N_4960);
xnor U5793 (N_5793,N_4563,N_4780);
xnor U5794 (N_5794,N_4759,N_4515);
or U5795 (N_5795,N_4541,N_4152);
xnor U5796 (N_5796,N_4962,N_4070);
or U5797 (N_5797,N_4637,N_4113);
or U5798 (N_5798,N_4690,N_4403);
and U5799 (N_5799,N_4908,N_4439);
nand U5800 (N_5800,N_4916,N_4439);
nor U5801 (N_5801,N_4164,N_4061);
nor U5802 (N_5802,N_4742,N_4589);
nor U5803 (N_5803,N_4048,N_4370);
xnor U5804 (N_5804,N_4833,N_4059);
nor U5805 (N_5805,N_4670,N_4126);
and U5806 (N_5806,N_4196,N_4912);
nor U5807 (N_5807,N_4798,N_4785);
nand U5808 (N_5808,N_4838,N_4958);
or U5809 (N_5809,N_4775,N_4519);
and U5810 (N_5810,N_4276,N_4354);
nor U5811 (N_5811,N_4973,N_4426);
and U5812 (N_5812,N_4202,N_4743);
or U5813 (N_5813,N_4242,N_4392);
xnor U5814 (N_5814,N_4147,N_4677);
or U5815 (N_5815,N_4987,N_4125);
nand U5816 (N_5816,N_4586,N_4189);
and U5817 (N_5817,N_4715,N_4162);
nor U5818 (N_5818,N_4323,N_4017);
nand U5819 (N_5819,N_4480,N_4544);
nor U5820 (N_5820,N_4028,N_4950);
and U5821 (N_5821,N_4455,N_4032);
or U5822 (N_5822,N_4846,N_4097);
nor U5823 (N_5823,N_4817,N_4643);
xnor U5824 (N_5824,N_4309,N_4061);
or U5825 (N_5825,N_4739,N_4153);
and U5826 (N_5826,N_4276,N_4359);
and U5827 (N_5827,N_4594,N_4912);
nor U5828 (N_5828,N_4262,N_4405);
nor U5829 (N_5829,N_4579,N_4500);
and U5830 (N_5830,N_4838,N_4753);
xnor U5831 (N_5831,N_4028,N_4569);
and U5832 (N_5832,N_4319,N_4853);
and U5833 (N_5833,N_4416,N_4925);
nor U5834 (N_5834,N_4652,N_4625);
nor U5835 (N_5835,N_4846,N_4251);
nor U5836 (N_5836,N_4490,N_4620);
nor U5837 (N_5837,N_4044,N_4082);
and U5838 (N_5838,N_4871,N_4565);
or U5839 (N_5839,N_4194,N_4978);
xor U5840 (N_5840,N_4197,N_4952);
and U5841 (N_5841,N_4731,N_4140);
nand U5842 (N_5842,N_4229,N_4463);
and U5843 (N_5843,N_4066,N_4652);
xnor U5844 (N_5844,N_4107,N_4574);
xnor U5845 (N_5845,N_4103,N_4046);
and U5846 (N_5846,N_4222,N_4358);
nand U5847 (N_5847,N_4572,N_4275);
nor U5848 (N_5848,N_4540,N_4621);
xor U5849 (N_5849,N_4422,N_4091);
nand U5850 (N_5850,N_4102,N_4699);
and U5851 (N_5851,N_4859,N_4201);
xor U5852 (N_5852,N_4951,N_4929);
and U5853 (N_5853,N_4682,N_4863);
nor U5854 (N_5854,N_4490,N_4928);
nand U5855 (N_5855,N_4067,N_4246);
nand U5856 (N_5856,N_4217,N_4440);
nor U5857 (N_5857,N_4124,N_4641);
nor U5858 (N_5858,N_4981,N_4297);
or U5859 (N_5859,N_4689,N_4216);
xnor U5860 (N_5860,N_4236,N_4294);
nor U5861 (N_5861,N_4004,N_4258);
or U5862 (N_5862,N_4944,N_4177);
nor U5863 (N_5863,N_4563,N_4090);
or U5864 (N_5864,N_4933,N_4596);
and U5865 (N_5865,N_4163,N_4492);
nand U5866 (N_5866,N_4342,N_4297);
and U5867 (N_5867,N_4088,N_4462);
or U5868 (N_5868,N_4500,N_4205);
nor U5869 (N_5869,N_4886,N_4930);
nor U5870 (N_5870,N_4170,N_4613);
and U5871 (N_5871,N_4512,N_4889);
nor U5872 (N_5872,N_4345,N_4493);
nand U5873 (N_5873,N_4643,N_4314);
nand U5874 (N_5874,N_4617,N_4612);
and U5875 (N_5875,N_4654,N_4924);
xnor U5876 (N_5876,N_4529,N_4751);
and U5877 (N_5877,N_4161,N_4260);
nor U5878 (N_5878,N_4569,N_4168);
xnor U5879 (N_5879,N_4258,N_4976);
or U5880 (N_5880,N_4589,N_4665);
nor U5881 (N_5881,N_4866,N_4868);
nand U5882 (N_5882,N_4054,N_4641);
nand U5883 (N_5883,N_4305,N_4045);
and U5884 (N_5884,N_4841,N_4926);
or U5885 (N_5885,N_4103,N_4330);
xor U5886 (N_5886,N_4060,N_4742);
and U5887 (N_5887,N_4112,N_4951);
nor U5888 (N_5888,N_4731,N_4900);
or U5889 (N_5889,N_4554,N_4292);
nand U5890 (N_5890,N_4722,N_4294);
and U5891 (N_5891,N_4685,N_4006);
nand U5892 (N_5892,N_4807,N_4747);
nor U5893 (N_5893,N_4232,N_4160);
xnor U5894 (N_5894,N_4194,N_4280);
nor U5895 (N_5895,N_4017,N_4760);
nor U5896 (N_5896,N_4024,N_4005);
and U5897 (N_5897,N_4158,N_4385);
or U5898 (N_5898,N_4684,N_4774);
nand U5899 (N_5899,N_4899,N_4794);
nand U5900 (N_5900,N_4532,N_4092);
nand U5901 (N_5901,N_4781,N_4556);
and U5902 (N_5902,N_4972,N_4557);
xor U5903 (N_5903,N_4221,N_4425);
nand U5904 (N_5904,N_4907,N_4280);
and U5905 (N_5905,N_4680,N_4447);
nor U5906 (N_5906,N_4190,N_4980);
or U5907 (N_5907,N_4445,N_4943);
xor U5908 (N_5908,N_4034,N_4985);
or U5909 (N_5909,N_4623,N_4433);
xnor U5910 (N_5910,N_4319,N_4085);
nand U5911 (N_5911,N_4815,N_4771);
and U5912 (N_5912,N_4111,N_4773);
and U5913 (N_5913,N_4443,N_4454);
nor U5914 (N_5914,N_4516,N_4153);
xor U5915 (N_5915,N_4626,N_4655);
nand U5916 (N_5916,N_4605,N_4518);
xnor U5917 (N_5917,N_4084,N_4628);
or U5918 (N_5918,N_4698,N_4503);
xnor U5919 (N_5919,N_4439,N_4090);
xor U5920 (N_5920,N_4203,N_4939);
and U5921 (N_5921,N_4468,N_4404);
and U5922 (N_5922,N_4935,N_4867);
or U5923 (N_5923,N_4857,N_4916);
or U5924 (N_5924,N_4297,N_4016);
nor U5925 (N_5925,N_4171,N_4294);
xor U5926 (N_5926,N_4196,N_4452);
nor U5927 (N_5927,N_4100,N_4538);
nor U5928 (N_5928,N_4880,N_4871);
xor U5929 (N_5929,N_4549,N_4902);
nand U5930 (N_5930,N_4965,N_4228);
and U5931 (N_5931,N_4946,N_4654);
nand U5932 (N_5932,N_4426,N_4726);
or U5933 (N_5933,N_4215,N_4107);
nand U5934 (N_5934,N_4461,N_4801);
nand U5935 (N_5935,N_4981,N_4797);
nor U5936 (N_5936,N_4374,N_4122);
or U5937 (N_5937,N_4079,N_4042);
nand U5938 (N_5938,N_4803,N_4472);
nor U5939 (N_5939,N_4317,N_4658);
and U5940 (N_5940,N_4177,N_4059);
xor U5941 (N_5941,N_4041,N_4392);
and U5942 (N_5942,N_4582,N_4590);
or U5943 (N_5943,N_4215,N_4068);
nor U5944 (N_5944,N_4357,N_4608);
xnor U5945 (N_5945,N_4645,N_4044);
nand U5946 (N_5946,N_4642,N_4268);
and U5947 (N_5947,N_4026,N_4486);
nor U5948 (N_5948,N_4569,N_4269);
nor U5949 (N_5949,N_4212,N_4084);
nand U5950 (N_5950,N_4866,N_4532);
nand U5951 (N_5951,N_4929,N_4700);
xnor U5952 (N_5952,N_4999,N_4778);
or U5953 (N_5953,N_4310,N_4043);
and U5954 (N_5954,N_4899,N_4083);
and U5955 (N_5955,N_4233,N_4129);
xnor U5956 (N_5956,N_4467,N_4257);
and U5957 (N_5957,N_4808,N_4197);
xor U5958 (N_5958,N_4508,N_4288);
and U5959 (N_5959,N_4238,N_4608);
and U5960 (N_5960,N_4002,N_4662);
or U5961 (N_5961,N_4147,N_4810);
xor U5962 (N_5962,N_4040,N_4625);
or U5963 (N_5963,N_4273,N_4468);
nand U5964 (N_5964,N_4243,N_4271);
nand U5965 (N_5965,N_4899,N_4456);
xnor U5966 (N_5966,N_4927,N_4911);
or U5967 (N_5967,N_4840,N_4456);
nand U5968 (N_5968,N_4346,N_4783);
nor U5969 (N_5969,N_4247,N_4338);
or U5970 (N_5970,N_4301,N_4633);
xnor U5971 (N_5971,N_4344,N_4628);
nand U5972 (N_5972,N_4863,N_4990);
nand U5973 (N_5973,N_4422,N_4989);
xor U5974 (N_5974,N_4511,N_4657);
nor U5975 (N_5975,N_4373,N_4548);
xnor U5976 (N_5976,N_4723,N_4089);
or U5977 (N_5977,N_4519,N_4379);
xnor U5978 (N_5978,N_4124,N_4561);
xor U5979 (N_5979,N_4086,N_4817);
nand U5980 (N_5980,N_4507,N_4851);
nand U5981 (N_5981,N_4107,N_4681);
or U5982 (N_5982,N_4829,N_4227);
nand U5983 (N_5983,N_4671,N_4344);
xor U5984 (N_5984,N_4424,N_4669);
and U5985 (N_5985,N_4701,N_4877);
nor U5986 (N_5986,N_4846,N_4897);
nor U5987 (N_5987,N_4555,N_4831);
and U5988 (N_5988,N_4274,N_4562);
or U5989 (N_5989,N_4483,N_4999);
nand U5990 (N_5990,N_4712,N_4120);
xor U5991 (N_5991,N_4825,N_4691);
and U5992 (N_5992,N_4288,N_4497);
nand U5993 (N_5993,N_4256,N_4147);
and U5994 (N_5994,N_4836,N_4629);
and U5995 (N_5995,N_4282,N_4129);
or U5996 (N_5996,N_4883,N_4156);
and U5997 (N_5997,N_4298,N_4623);
and U5998 (N_5998,N_4717,N_4951);
and U5999 (N_5999,N_4988,N_4598);
nor U6000 (N_6000,N_5521,N_5972);
and U6001 (N_6001,N_5742,N_5625);
nand U6002 (N_6002,N_5507,N_5875);
nor U6003 (N_6003,N_5609,N_5828);
and U6004 (N_6004,N_5141,N_5228);
nor U6005 (N_6005,N_5271,N_5378);
nor U6006 (N_6006,N_5598,N_5415);
xor U6007 (N_6007,N_5465,N_5993);
and U6008 (N_6008,N_5599,N_5475);
nor U6009 (N_6009,N_5057,N_5023);
nor U6010 (N_6010,N_5254,N_5160);
and U6011 (N_6011,N_5178,N_5398);
or U6012 (N_6012,N_5355,N_5820);
nor U6013 (N_6013,N_5102,N_5547);
nand U6014 (N_6014,N_5528,N_5269);
and U6015 (N_6015,N_5846,N_5296);
xnor U6016 (N_6016,N_5761,N_5764);
nand U6017 (N_6017,N_5455,N_5476);
nor U6018 (N_6018,N_5444,N_5147);
or U6019 (N_6019,N_5631,N_5028);
xnor U6020 (N_6020,N_5516,N_5853);
or U6021 (N_6021,N_5128,N_5186);
and U6022 (N_6022,N_5816,N_5255);
or U6023 (N_6023,N_5244,N_5669);
nor U6024 (N_6024,N_5084,N_5462);
xnor U6025 (N_6025,N_5637,N_5103);
xor U6026 (N_6026,N_5098,N_5788);
and U6027 (N_6027,N_5422,N_5293);
nand U6028 (N_6028,N_5689,N_5275);
nor U6029 (N_6029,N_5396,N_5333);
and U6030 (N_6030,N_5308,N_5407);
nand U6031 (N_6031,N_5922,N_5077);
and U6032 (N_6032,N_5985,N_5947);
or U6033 (N_6033,N_5750,N_5302);
xor U6034 (N_6034,N_5582,N_5665);
nand U6035 (N_6035,N_5256,N_5388);
or U6036 (N_6036,N_5896,N_5526);
nor U6037 (N_6037,N_5174,N_5496);
nor U6038 (N_6038,N_5871,N_5113);
and U6039 (N_6039,N_5586,N_5723);
nand U6040 (N_6040,N_5849,N_5703);
or U6041 (N_6041,N_5721,N_5978);
or U6042 (N_6042,N_5202,N_5322);
nand U6043 (N_6043,N_5060,N_5889);
xor U6044 (N_6044,N_5590,N_5183);
nor U6045 (N_6045,N_5215,N_5911);
nor U6046 (N_6046,N_5674,N_5320);
nand U6047 (N_6047,N_5424,N_5038);
nand U6048 (N_6048,N_5180,N_5165);
xor U6049 (N_6049,N_5150,N_5205);
and U6050 (N_6050,N_5488,N_5367);
or U6051 (N_6051,N_5633,N_5433);
nand U6052 (N_6052,N_5695,N_5574);
nor U6053 (N_6053,N_5391,N_5067);
and U6054 (N_6054,N_5880,N_5305);
nor U6055 (N_6055,N_5207,N_5680);
xor U6056 (N_6056,N_5681,N_5117);
or U6057 (N_6057,N_5752,N_5482);
and U6058 (N_6058,N_5263,N_5121);
nand U6059 (N_6059,N_5096,N_5048);
nand U6060 (N_6060,N_5604,N_5274);
xnor U6061 (N_6061,N_5670,N_5266);
xnor U6062 (N_6062,N_5214,N_5027);
nor U6063 (N_6063,N_5557,N_5401);
or U6064 (N_6064,N_5942,N_5551);
and U6065 (N_6065,N_5618,N_5058);
and U6066 (N_6066,N_5678,N_5746);
nand U6067 (N_6067,N_5197,N_5236);
or U6068 (N_6068,N_5111,N_5356);
xnor U6069 (N_6069,N_5369,N_5239);
and U6070 (N_6070,N_5312,N_5222);
nand U6071 (N_6071,N_5772,N_5417);
xor U6072 (N_6072,N_5389,N_5134);
xnor U6073 (N_6073,N_5535,N_5017);
nand U6074 (N_6074,N_5890,N_5129);
xnor U6075 (N_6075,N_5710,N_5770);
nand U6076 (N_6076,N_5387,N_5039);
nand U6077 (N_6077,N_5583,N_5522);
and U6078 (N_6078,N_5650,N_5468);
nor U6079 (N_6079,N_5785,N_5954);
nand U6080 (N_6080,N_5285,N_5497);
nand U6081 (N_6081,N_5578,N_5203);
xnor U6082 (N_6082,N_5923,N_5863);
nor U6083 (N_6083,N_5780,N_5216);
xnor U6084 (N_6084,N_5570,N_5511);
nor U6085 (N_6085,N_5635,N_5221);
xnor U6086 (N_6086,N_5445,N_5858);
nand U6087 (N_6087,N_5061,N_5987);
xor U6088 (N_6088,N_5009,N_5399);
nand U6089 (N_6089,N_5775,N_5852);
and U6090 (N_6090,N_5409,N_5519);
and U6091 (N_6091,N_5966,N_5999);
xnor U6092 (N_6092,N_5323,N_5166);
xnor U6093 (N_6093,N_5257,N_5550);
nor U6094 (N_6094,N_5158,N_5553);
and U6095 (N_6095,N_5525,N_5850);
nor U6096 (N_6096,N_5037,N_5666);
nand U6097 (N_6097,N_5301,N_5753);
nand U6098 (N_6098,N_5054,N_5163);
or U6099 (N_6099,N_5608,N_5545);
xor U6100 (N_6100,N_5071,N_5848);
xnor U6101 (N_6101,N_5382,N_5095);
xor U6102 (N_6102,N_5171,N_5684);
nand U6103 (N_6103,N_5493,N_5515);
nor U6104 (N_6104,N_5510,N_5287);
nor U6105 (N_6105,N_5626,N_5247);
nor U6106 (N_6106,N_5963,N_5575);
nor U6107 (N_6107,N_5331,N_5246);
nor U6108 (N_6108,N_5267,N_5139);
xor U6109 (N_6109,N_5512,N_5107);
nor U6110 (N_6110,N_5672,N_5745);
nand U6111 (N_6111,N_5769,N_5800);
or U6112 (N_6112,N_5088,N_5936);
nand U6113 (N_6113,N_5719,N_5938);
or U6114 (N_6114,N_5304,N_5699);
or U6115 (N_6115,N_5019,N_5573);
and U6116 (N_6116,N_5974,N_5961);
xor U6117 (N_6117,N_5649,N_5925);
xnor U6118 (N_6118,N_5075,N_5930);
or U6119 (N_6119,N_5464,N_5135);
nor U6120 (N_6120,N_5825,N_5621);
xor U6121 (N_6121,N_5435,N_5109);
nand U6122 (N_6122,N_5142,N_5513);
and U6123 (N_6123,N_5994,N_5687);
and U6124 (N_6124,N_5926,N_5851);
and U6125 (N_6125,N_5335,N_5073);
nand U6126 (N_6126,N_5600,N_5471);
and U6127 (N_6127,N_5503,N_5085);
and U6128 (N_6128,N_5414,N_5504);
nor U6129 (N_6129,N_5904,N_5835);
nand U6130 (N_6130,N_5339,N_5393);
nor U6131 (N_6131,N_5998,N_5748);
xor U6132 (N_6132,N_5225,N_5238);
nand U6133 (N_6133,N_5831,N_5146);
and U6134 (N_6134,N_5924,N_5363);
or U6135 (N_6135,N_5122,N_5726);
nand U6136 (N_6136,N_5402,N_5562);
or U6137 (N_6137,N_5155,N_5306);
or U6138 (N_6138,N_5405,N_5962);
xor U6139 (N_6139,N_5112,N_5912);
or U6140 (N_6140,N_5212,N_5231);
and U6141 (N_6141,N_5640,N_5892);
nand U6142 (N_6142,N_5997,N_5400);
and U6143 (N_6143,N_5636,N_5549);
nor U6144 (N_6144,N_5241,N_5097);
xor U6145 (N_6145,N_5458,N_5866);
and U6146 (N_6146,N_5771,N_5983);
nand U6147 (N_6147,N_5778,N_5300);
and U6148 (N_6148,N_5470,N_5564);
and U6149 (N_6149,N_5918,N_5052);
and U6150 (N_6150,N_5690,N_5226);
or U6151 (N_6151,N_5260,N_5698);
and U6152 (N_6152,N_5796,N_5877);
nand U6153 (N_6153,N_5701,N_5007);
nand U6154 (N_6154,N_5706,N_5451);
nand U6155 (N_6155,N_5539,N_5090);
and U6156 (N_6156,N_5727,N_5492);
nand U6157 (N_6157,N_5715,N_5679);
and U6158 (N_6158,N_5661,N_5694);
or U6159 (N_6159,N_5676,N_5015);
or U6160 (N_6160,N_5043,N_5478);
nand U6161 (N_6161,N_5316,N_5986);
xor U6162 (N_6162,N_5533,N_5532);
or U6163 (N_6163,N_5830,N_5234);
and U6164 (N_6164,N_5707,N_5131);
nand U6165 (N_6165,N_5350,N_5810);
nand U6166 (N_6166,N_5971,N_5291);
or U6167 (N_6167,N_5915,N_5728);
nor U6168 (N_6168,N_5232,N_5844);
nand U6169 (N_6169,N_5235,N_5928);
and U6170 (N_6170,N_5196,N_5654);
nor U6171 (N_6171,N_5298,N_5423);
nand U6172 (N_6172,N_5783,N_5354);
xnor U6173 (N_6173,N_5299,N_5161);
or U6174 (N_6174,N_5480,N_5991);
nand U6175 (N_6175,N_5591,N_5885);
nand U6176 (N_6176,N_5056,N_5781);
and U6177 (N_6177,N_5001,N_5279);
and U6178 (N_6178,N_5977,N_5798);
nand U6179 (N_6179,N_5760,N_5651);
nor U6180 (N_6180,N_5869,N_5711);
nand U6181 (N_6181,N_5939,N_5086);
xnor U6182 (N_6182,N_5349,N_5328);
xnor U6183 (N_6183,N_5708,N_5091);
or U6184 (N_6184,N_5420,N_5886);
and U6185 (N_6185,N_5273,N_5290);
nand U6186 (N_6186,N_5933,N_5779);
and U6187 (N_6187,N_5377,N_5594);
nor U6188 (N_6188,N_5094,N_5566);
and U6189 (N_6189,N_5580,N_5531);
nand U6190 (N_6190,N_5743,N_5457);
xor U6191 (N_6191,N_5348,N_5499);
nor U6192 (N_6192,N_5395,N_5068);
or U6193 (N_6193,N_5883,N_5452);
and U6194 (N_6194,N_5144,N_5537);
or U6195 (N_6195,N_5408,N_5261);
xor U6196 (N_6196,N_5882,N_5344);
nand U6197 (N_6197,N_5763,N_5448);
nand U6198 (N_6198,N_5530,N_5087);
nor U6199 (N_6199,N_5000,N_5258);
nand U6200 (N_6200,N_5546,N_5603);
nor U6201 (N_6201,N_5127,N_5916);
or U6202 (N_6202,N_5114,N_5065);
and U6203 (N_6203,N_5948,N_5115);
nand U6204 (N_6204,N_5031,N_5992);
nand U6205 (N_6205,N_5156,N_5805);
nand U6206 (N_6206,N_5739,N_5317);
xor U6207 (N_6207,N_5441,N_5861);
and U6208 (N_6208,N_5069,N_5958);
nor U6209 (N_6209,N_5303,N_5657);
xor U6210 (N_6210,N_5380,N_5064);
or U6211 (N_6211,N_5572,N_5149);
or U6212 (N_6212,N_5313,N_5342);
xor U6213 (N_6213,N_5229,N_5286);
nand U6214 (N_6214,N_5804,N_5116);
and U6215 (N_6215,N_5130,N_5988);
xnor U6216 (N_6216,N_5026,N_5093);
and U6217 (N_6217,N_5449,N_5901);
and U6218 (N_6218,N_5979,N_5191);
or U6219 (N_6219,N_5284,N_5766);
xor U6220 (N_6220,N_5453,N_5211);
and U6221 (N_6221,N_5867,N_5264);
and U6222 (N_6222,N_5647,N_5059);
xor U6223 (N_6223,N_5919,N_5645);
nor U6224 (N_6224,N_5747,N_5686);
xor U6225 (N_6225,N_5738,N_5597);
or U6226 (N_6226,N_5995,N_5192);
and U6227 (N_6227,N_5538,N_5252);
and U6228 (N_6228,N_5152,N_5439);
and U6229 (N_6229,N_5104,N_5860);
nor U6230 (N_6230,N_5619,N_5506);
or U6231 (N_6231,N_5730,N_5474);
or U6232 (N_6232,N_5479,N_5815);
nor U6233 (N_6233,N_5555,N_5319);
or U6234 (N_6234,N_5589,N_5934);
and U6235 (N_6235,N_5432,N_5614);
nor U6236 (N_6236,N_5210,N_5485);
nand U6237 (N_6237,N_5277,N_5187);
nor U6238 (N_6238,N_5042,N_5421);
xor U6239 (N_6239,N_5789,N_5249);
nor U6240 (N_6240,N_5253,N_5935);
or U6241 (N_6241,N_5812,N_5632);
xor U6242 (N_6242,N_5945,N_5957);
nor U6243 (N_6243,N_5872,N_5419);
xnor U6244 (N_6244,N_5136,N_5579);
and U6245 (N_6245,N_5782,N_5008);
nor U6246 (N_6246,N_5888,N_5843);
xor U6247 (N_6247,N_5989,N_5491);
and U6248 (N_6248,N_5696,N_5372);
and U6249 (N_6249,N_5472,N_5683);
and U6250 (N_6250,N_5955,N_5824);
nor U6251 (N_6251,N_5898,N_5386);
xor U6252 (N_6252,N_5145,N_5324);
xnor U6253 (N_6253,N_5371,N_5032);
nor U6254 (N_6254,N_5663,N_5700);
or U6255 (N_6255,N_5230,N_5341);
and U6256 (N_6256,N_5737,N_5949);
nor U6257 (N_6257,N_5223,N_5361);
or U6258 (N_6258,N_5964,N_5394);
nor U6259 (N_6259,N_5410,N_5865);
and U6260 (N_6260,N_5219,N_5834);
nand U6261 (N_6261,N_5662,N_5385);
nor U6262 (N_6262,N_5280,N_5213);
xor U6263 (N_6263,N_5240,N_5601);
and U6264 (N_6264,N_5125,N_5829);
or U6265 (N_6265,N_5646,N_5375);
nor U6266 (N_6266,N_5514,N_5897);
xnor U6267 (N_6267,N_5404,N_5741);
xor U6268 (N_6268,N_5906,N_5642);
or U6269 (N_6269,N_5732,N_5460);
xnor U6270 (N_6270,N_5920,N_5554);
and U6271 (N_6271,N_5664,N_5283);
and U6272 (N_6272,N_5776,N_5259);
or U6273 (N_6273,N_5383,N_5195);
nor U6274 (N_6274,N_5046,N_5675);
nand U6275 (N_6275,N_5329,N_5047);
nor U6276 (N_6276,N_5330,N_5101);
xnor U6277 (N_6277,N_5802,N_5688);
or U6278 (N_6278,N_5173,N_5893);
xor U6279 (N_6279,N_5629,N_5425);
nor U6280 (N_6280,N_5940,N_5660);
and U6281 (N_6281,N_5030,N_5864);
nand U6282 (N_6282,N_5790,N_5859);
or U6283 (N_6283,N_5080,N_5245);
or U6284 (N_6284,N_5941,N_5910);
and U6285 (N_6285,N_5157,N_5177);
and U6286 (N_6286,N_5814,N_5327);
and U6287 (N_6287,N_5697,N_5132);
nor U6288 (N_6288,N_5990,N_5821);
nor U6289 (N_6289,N_5801,N_5729);
xor U6290 (N_6290,N_5063,N_5489);
xor U6291 (N_6291,N_5169,N_5819);
nor U6292 (N_6292,N_5833,N_5894);
or U6293 (N_6293,N_5189,N_5012);
nor U6294 (N_6294,N_5029,N_5418);
and U6295 (N_6295,N_5184,N_5913);
xor U6296 (N_6296,N_5365,N_5921);
or U6297 (N_6297,N_5975,N_5845);
xnor U6298 (N_6298,N_5237,N_5416);
nand U6299 (N_6299,N_5929,N_5011);
or U6300 (N_6300,N_5704,N_5352);
xnor U6301 (N_6301,N_5768,N_5944);
nand U6302 (N_6302,N_5596,N_5176);
xor U6303 (N_6303,N_5656,N_5874);
xor U6304 (N_6304,N_5952,N_5841);
xor U6305 (N_6305,N_5517,N_5099);
xnor U6306 (N_6306,N_5803,N_5053);
nand U6307 (N_6307,N_5854,N_5895);
xor U6308 (N_6308,N_5051,N_5784);
nand U6309 (N_6309,N_5022,N_5250);
or U6310 (N_6310,N_5765,N_5368);
xnor U6311 (N_6311,N_5390,N_5908);
nand U6312 (N_6312,N_5643,N_5151);
or U6313 (N_6313,N_5270,N_5374);
nand U6314 (N_6314,N_5630,N_5217);
and U6315 (N_6315,N_5050,N_5120);
nand U6316 (N_6316,N_5667,N_5137);
nand U6317 (N_6317,N_5438,N_5823);
or U6318 (N_6318,N_5878,N_5907);
xnor U6319 (N_6319,N_5403,N_5639);
or U6320 (N_6320,N_5899,N_5552);
and U6321 (N_6321,N_5624,N_5794);
nand U6322 (N_6322,N_5321,N_5276);
nor U6323 (N_6323,N_5502,N_5641);
xnor U6324 (N_6324,N_5456,N_5620);
nand U6325 (N_6325,N_5967,N_5153);
xor U6326 (N_6326,N_5036,N_5175);
nor U6327 (N_6327,N_5932,N_5827);
or U6328 (N_6328,N_5969,N_5837);
nand U6329 (N_6329,N_5126,N_5446);
nor U6330 (N_6330,N_5025,N_5822);
nand U6331 (N_6331,N_5072,N_5959);
nor U6332 (N_6332,N_5079,N_5295);
nor U6333 (N_6333,N_5242,N_5611);
nor U6334 (N_6334,N_5034,N_5541);
nor U6335 (N_6335,N_5351,N_5100);
and U6336 (N_6336,N_5204,N_5358);
nor U6337 (N_6337,N_5498,N_5868);
xor U6338 (N_6338,N_5787,N_5345);
or U6339 (N_6339,N_5292,N_5370);
or U6340 (N_6340,N_5110,N_5634);
and U6341 (N_6341,N_5494,N_5288);
nor U6342 (N_6342,N_5795,N_5725);
or U6343 (N_6343,N_5903,N_5658);
and U6344 (N_6344,N_5200,N_5487);
or U6345 (N_6345,N_5148,N_5227);
xor U6346 (N_6346,N_5140,N_5188);
xor U6347 (N_6347,N_5536,N_5673);
nand U6348 (N_6348,N_5965,N_5713);
and U6349 (N_6349,N_5567,N_5671);
or U6350 (N_6350,N_5759,N_5193);
nor U6351 (N_6351,N_5198,N_5900);
nor U6352 (N_6352,N_5172,N_5450);
nand U6353 (N_6353,N_5722,N_5045);
nor U6354 (N_6354,N_5543,N_5447);
xor U6355 (N_6355,N_5556,N_5756);
xor U6356 (N_6356,N_5876,N_5887);
and U6357 (N_6357,N_5190,N_5762);
or U6358 (N_6358,N_5490,N_5384);
xnor U6359 (N_6359,N_5199,N_5092);
nand U6360 (N_6360,N_5716,N_5870);
nor U6361 (N_6361,N_5343,N_5044);
nor U6362 (N_6362,N_5818,N_5616);
nor U6363 (N_6363,N_5581,N_5278);
nand U6364 (N_6364,N_5524,N_5773);
or U6365 (N_6365,N_5454,N_5495);
nor U6366 (N_6366,N_5839,N_5440);
nor U6367 (N_6367,N_5020,N_5976);
nand U6368 (N_6368,N_5705,N_5248);
or U6369 (N_6369,N_5381,N_5162);
nand U6370 (N_6370,N_5744,N_5527);
or U6371 (N_6371,N_5652,N_5477);
nand U6372 (N_6372,N_5182,N_5791);
nand U6373 (N_6373,N_5082,N_5627);
or U6374 (N_6374,N_5811,N_5607);
nand U6375 (N_6375,N_5340,N_5544);
xor U6376 (N_6376,N_5392,N_5655);
nand U6377 (N_6377,N_5500,N_5311);
nand U6378 (N_6378,N_5006,N_5168);
xnor U6379 (N_6379,N_5337,N_5758);
nand U6380 (N_6380,N_5428,N_5733);
and U6381 (N_6381,N_5584,N_5960);
nand U6382 (N_6382,N_5813,N_5461);
or U6383 (N_6383,N_5638,N_5243);
nand U6384 (N_6384,N_5406,N_5587);
and U6385 (N_6385,N_5055,N_5777);
nand U6386 (N_6386,N_5857,N_5281);
nand U6387 (N_6387,N_5862,N_5879);
nand U6388 (N_6388,N_5891,N_5612);
xor U6389 (N_6389,N_5873,N_5605);
nor U6390 (N_6390,N_5426,N_5397);
and U6391 (N_6391,N_5682,N_5792);
nand U6392 (N_6392,N_5314,N_5167);
nand U6393 (N_6393,N_5508,N_5123);
nor U6394 (N_6394,N_5565,N_5076);
nand U6395 (N_6395,N_5668,N_5569);
nand U6396 (N_6396,N_5617,N_5807);
or U6397 (N_6397,N_5809,N_5459);
and U6398 (N_6398,N_5346,N_5430);
or U6399 (N_6399,N_5797,N_5937);
xor U6400 (N_6400,N_5653,N_5427);
xnor U6401 (N_6401,N_5289,N_5585);
nor U6402 (N_6402,N_5442,N_5836);
and U6403 (N_6403,N_5909,N_5014);
and U6404 (N_6404,N_5981,N_5588);
or U6405 (N_6405,N_5847,N_5373);
nand U6406 (N_6406,N_5035,N_5218);
nor U6407 (N_6407,N_5968,N_5693);
nor U6408 (N_6408,N_5364,N_5786);
and U6409 (N_6409,N_5412,N_5767);
nor U6410 (N_6410,N_5914,N_5606);
or U6411 (N_6411,N_5206,N_5118);
nor U6412 (N_6412,N_5793,N_5540);
nand U6413 (N_6413,N_5265,N_5360);
nand U6414 (N_6414,N_5953,N_5602);
nand U6415 (N_6415,N_5734,N_5548);
xnor U6416 (N_6416,N_5542,N_5749);
or U6417 (N_6417,N_5049,N_5083);
nand U6418 (N_6418,N_5509,N_5179);
and U6419 (N_6419,N_5436,N_5411);
xor U6420 (N_6420,N_5806,N_5709);
xor U6421 (N_6421,N_5613,N_5799);
nand U6422 (N_6422,N_5170,N_5659);
nand U6423 (N_6423,N_5610,N_5362);
nor U6424 (N_6424,N_5010,N_5070);
and U6425 (N_6425,N_5004,N_5951);
xnor U6426 (N_6426,N_5262,N_5041);
xor U6427 (N_6427,N_5297,N_5154);
nand U6428 (N_6428,N_5366,N_5826);
and U6429 (N_6429,N_5062,N_5755);
or U6430 (N_6430,N_5268,N_5013);
and U6431 (N_6431,N_5326,N_5379);
nand U6432 (N_6432,N_5469,N_5520);
or U6433 (N_6433,N_5712,N_5623);
nor U6434 (N_6434,N_5518,N_5956);
and U6435 (N_6435,N_5561,N_5577);
nor U6436 (N_6436,N_5754,N_5692);
xnor U6437 (N_6437,N_5105,N_5691);
xor U6438 (N_6438,N_5576,N_5855);
xnor U6439 (N_6439,N_5124,N_5164);
xnor U6440 (N_6440,N_5318,N_5838);
nor U6441 (N_6441,N_5463,N_5074);
and U6442 (N_6442,N_5950,N_5718);
or U6443 (N_6443,N_5856,N_5534);
nor U6444 (N_6444,N_5560,N_5970);
nand U6445 (N_6445,N_5902,N_5332);
and U6446 (N_6446,N_5159,N_5751);
or U6447 (N_6447,N_5466,N_5481);
or U6448 (N_6448,N_5003,N_5133);
nor U6449 (N_6449,N_5648,N_5840);
nand U6450 (N_6450,N_5194,N_5927);
and U6451 (N_6451,N_5622,N_5568);
nor U6452 (N_6452,N_5307,N_5081);
nor U6453 (N_6453,N_5143,N_5563);
nor U6454 (N_6454,N_5224,N_5353);
nand U6455 (N_6455,N_5434,N_5437);
nand U6456 (N_6456,N_5024,N_5066);
or U6457 (N_6457,N_5905,N_5018);
xnor U6458 (N_6458,N_5917,N_5002);
xnor U6459 (N_6459,N_5282,N_5309);
nand U6460 (N_6460,N_5431,N_5325);
nand U6461 (N_6461,N_5817,N_5016);
and U6462 (N_6462,N_5808,N_5106);
nor U6463 (N_6463,N_5484,N_5593);
xor U6464 (N_6464,N_5571,N_5996);
or U6465 (N_6465,N_5884,N_5220);
or U6466 (N_6466,N_5467,N_5005);
or U6467 (N_6467,N_5842,N_5592);
nor U6468 (N_6468,N_5529,N_5717);
and U6469 (N_6469,N_5443,N_5736);
nand U6470 (N_6470,N_5558,N_5021);
nand U6471 (N_6471,N_5982,N_5078);
xnor U6472 (N_6472,N_5201,N_5724);
nand U6473 (N_6473,N_5731,N_5740);
and U6474 (N_6474,N_5714,N_5931);
and U6475 (N_6475,N_5559,N_5980);
nor U6476 (N_6476,N_5628,N_5338);
nand U6477 (N_6477,N_5483,N_5973);
or U6478 (N_6478,N_5505,N_5943);
xor U6479 (N_6479,N_5233,N_5272);
or U6480 (N_6480,N_5735,N_5251);
and U6481 (N_6481,N_5336,N_5334);
nor U6482 (N_6482,N_5832,N_5685);
xnor U6483 (N_6483,N_5357,N_5310);
or U6484 (N_6484,N_5595,N_5294);
nor U6485 (N_6485,N_5359,N_5757);
nor U6486 (N_6486,N_5523,N_5376);
nand U6487 (N_6487,N_5347,N_5881);
or U6488 (N_6488,N_5185,N_5413);
and U6489 (N_6489,N_5946,N_5089);
nor U6490 (N_6490,N_5119,N_5473);
or U6491 (N_6491,N_5209,N_5033);
nor U6492 (N_6492,N_5774,N_5138);
and U6493 (N_6493,N_5677,N_5429);
nand U6494 (N_6494,N_5181,N_5108);
nor U6495 (N_6495,N_5486,N_5040);
or U6496 (N_6496,N_5720,N_5702);
nand U6497 (N_6497,N_5984,N_5501);
nand U6498 (N_6498,N_5315,N_5615);
or U6499 (N_6499,N_5208,N_5644);
or U6500 (N_6500,N_5254,N_5350);
nand U6501 (N_6501,N_5847,N_5574);
and U6502 (N_6502,N_5095,N_5737);
nand U6503 (N_6503,N_5087,N_5724);
nand U6504 (N_6504,N_5876,N_5175);
or U6505 (N_6505,N_5395,N_5830);
or U6506 (N_6506,N_5972,N_5383);
nor U6507 (N_6507,N_5096,N_5350);
nand U6508 (N_6508,N_5363,N_5167);
xor U6509 (N_6509,N_5227,N_5080);
or U6510 (N_6510,N_5884,N_5418);
and U6511 (N_6511,N_5341,N_5845);
nand U6512 (N_6512,N_5658,N_5679);
or U6513 (N_6513,N_5544,N_5311);
nor U6514 (N_6514,N_5432,N_5276);
nand U6515 (N_6515,N_5196,N_5548);
nand U6516 (N_6516,N_5275,N_5619);
and U6517 (N_6517,N_5082,N_5534);
nand U6518 (N_6518,N_5347,N_5459);
nor U6519 (N_6519,N_5640,N_5730);
nor U6520 (N_6520,N_5431,N_5216);
or U6521 (N_6521,N_5356,N_5832);
nand U6522 (N_6522,N_5123,N_5942);
xnor U6523 (N_6523,N_5467,N_5421);
nand U6524 (N_6524,N_5378,N_5471);
nand U6525 (N_6525,N_5319,N_5888);
or U6526 (N_6526,N_5040,N_5944);
xnor U6527 (N_6527,N_5155,N_5843);
xor U6528 (N_6528,N_5628,N_5461);
or U6529 (N_6529,N_5834,N_5361);
or U6530 (N_6530,N_5012,N_5947);
xor U6531 (N_6531,N_5384,N_5650);
or U6532 (N_6532,N_5283,N_5745);
nand U6533 (N_6533,N_5523,N_5460);
or U6534 (N_6534,N_5051,N_5117);
xnor U6535 (N_6535,N_5548,N_5671);
and U6536 (N_6536,N_5871,N_5553);
and U6537 (N_6537,N_5528,N_5939);
nor U6538 (N_6538,N_5298,N_5691);
nor U6539 (N_6539,N_5620,N_5186);
xor U6540 (N_6540,N_5193,N_5259);
nand U6541 (N_6541,N_5211,N_5664);
or U6542 (N_6542,N_5684,N_5303);
or U6543 (N_6543,N_5718,N_5122);
and U6544 (N_6544,N_5912,N_5426);
or U6545 (N_6545,N_5537,N_5495);
or U6546 (N_6546,N_5527,N_5993);
nand U6547 (N_6547,N_5010,N_5066);
nor U6548 (N_6548,N_5378,N_5910);
nor U6549 (N_6549,N_5912,N_5783);
or U6550 (N_6550,N_5146,N_5925);
nand U6551 (N_6551,N_5928,N_5119);
nor U6552 (N_6552,N_5548,N_5644);
or U6553 (N_6553,N_5785,N_5147);
nand U6554 (N_6554,N_5566,N_5469);
nand U6555 (N_6555,N_5356,N_5554);
nor U6556 (N_6556,N_5617,N_5183);
xnor U6557 (N_6557,N_5450,N_5091);
and U6558 (N_6558,N_5430,N_5498);
nor U6559 (N_6559,N_5845,N_5899);
nor U6560 (N_6560,N_5591,N_5524);
nand U6561 (N_6561,N_5204,N_5873);
or U6562 (N_6562,N_5617,N_5265);
or U6563 (N_6563,N_5718,N_5044);
and U6564 (N_6564,N_5505,N_5090);
nor U6565 (N_6565,N_5773,N_5588);
or U6566 (N_6566,N_5059,N_5586);
and U6567 (N_6567,N_5816,N_5425);
xor U6568 (N_6568,N_5523,N_5996);
nand U6569 (N_6569,N_5646,N_5001);
xnor U6570 (N_6570,N_5688,N_5743);
nor U6571 (N_6571,N_5881,N_5012);
and U6572 (N_6572,N_5628,N_5894);
or U6573 (N_6573,N_5113,N_5177);
xor U6574 (N_6574,N_5007,N_5298);
and U6575 (N_6575,N_5415,N_5067);
and U6576 (N_6576,N_5410,N_5106);
and U6577 (N_6577,N_5929,N_5813);
nor U6578 (N_6578,N_5505,N_5864);
or U6579 (N_6579,N_5359,N_5600);
nor U6580 (N_6580,N_5906,N_5865);
and U6581 (N_6581,N_5790,N_5614);
nand U6582 (N_6582,N_5764,N_5443);
nand U6583 (N_6583,N_5008,N_5910);
xor U6584 (N_6584,N_5421,N_5453);
or U6585 (N_6585,N_5741,N_5324);
or U6586 (N_6586,N_5878,N_5104);
nor U6587 (N_6587,N_5406,N_5740);
nor U6588 (N_6588,N_5466,N_5711);
or U6589 (N_6589,N_5970,N_5198);
nand U6590 (N_6590,N_5860,N_5135);
or U6591 (N_6591,N_5509,N_5954);
nor U6592 (N_6592,N_5783,N_5011);
nand U6593 (N_6593,N_5710,N_5576);
or U6594 (N_6594,N_5626,N_5692);
xnor U6595 (N_6595,N_5892,N_5466);
xor U6596 (N_6596,N_5272,N_5586);
xnor U6597 (N_6597,N_5970,N_5825);
and U6598 (N_6598,N_5028,N_5819);
and U6599 (N_6599,N_5028,N_5252);
and U6600 (N_6600,N_5153,N_5472);
nor U6601 (N_6601,N_5303,N_5333);
xor U6602 (N_6602,N_5063,N_5213);
nor U6603 (N_6603,N_5368,N_5562);
nor U6604 (N_6604,N_5990,N_5501);
nor U6605 (N_6605,N_5503,N_5240);
or U6606 (N_6606,N_5176,N_5192);
nor U6607 (N_6607,N_5186,N_5273);
nand U6608 (N_6608,N_5329,N_5250);
nor U6609 (N_6609,N_5570,N_5991);
nand U6610 (N_6610,N_5672,N_5630);
and U6611 (N_6611,N_5902,N_5899);
nor U6612 (N_6612,N_5296,N_5698);
and U6613 (N_6613,N_5686,N_5197);
nor U6614 (N_6614,N_5537,N_5397);
and U6615 (N_6615,N_5660,N_5174);
or U6616 (N_6616,N_5636,N_5290);
or U6617 (N_6617,N_5964,N_5650);
or U6618 (N_6618,N_5782,N_5912);
nand U6619 (N_6619,N_5458,N_5298);
nand U6620 (N_6620,N_5865,N_5871);
or U6621 (N_6621,N_5917,N_5759);
or U6622 (N_6622,N_5730,N_5834);
and U6623 (N_6623,N_5068,N_5926);
or U6624 (N_6624,N_5118,N_5038);
nand U6625 (N_6625,N_5067,N_5596);
nor U6626 (N_6626,N_5741,N_5244);
xnor U6627 (N_6627,N_5784,N_5231);
nor U6628 (N_6628,N_5365,N_5609);
or U6629 (N_6629,N_5807,N_5030);
and U6630 (N_6630,N_5662,N_5043);
or U6631 (N_6631,N_5598,N_5447);
nor U6632 (N_6632,N_5911,N_5060);
nor U6633 (N_6633,N_5661,N_5646);
or U6634 (N_6634,N_5644,N_5429);
or U6635 (N_6635,N_5173,N_5187);
nand U6636 (N_6636,N_5858,N_5722);
or U6637 (N_6637,N_5562,N_5040);
or U6638 (N_6638,N_5958,N_5965);
xnor U6639 (N_6639,N_5412,N_5705);
and U6640 (N_6640,N_5544,N_5124);
nor U6641 (N_6641,N_5884,N_5605);
nand U6642 (N_6642,N_5963,N_5170);
and U6643 (N_6643,N_5147,N_5236);
or U6644 (N_6644,N_5738,N_5778);
nand U6645 (N_6645,N_5355,N_5562);
nand U6646 (N_6646,N_5687,N_5806);
xnor U6647 (N_6647,N_5804,N_5571);
and U6648 (N_6648,N_5217,N_5801);
or U6649 (N_6649,N_5766,N_5817);
and U6650 (N_6650,N_5476,N_5156);
nor U6651 (N_6651,N_5075,N_5239);
nor U6652 (N_6652,N_5542,N_5142);
nor U6653 (N_6653,N_5619,N_5571);
nor U6654 (N_6654,N_5819,N_5912);
nor U6655 (N_6655,N_5307,N_5778);
nand U6656 (N_6656,N_5226,N_5820);
or U6657 (N_6657,N_5543,N_5455);
xor U6658 (N_6658,N_5288,N_5322);
and U6659 (N_6659,N_5558,N_5787);
nand U6660 (N_6660,N_5073,N_5720);
xor U6661 (N_6661,N_5666,N_5167);
nor U6662 (N_6662,N_5732,N_5476);
or U6663 (N_6663,N_5281,N_5952);
nor U6664 (N_6664,N_5663,N_5314);
or U6665 (N_6665,N_5892,N_5034);
or U6666 (N_6666,N_5796,N_5513);
xor U6667 (N_6667,N_5673,N_5580);
or U6668 (N_6668,N_5679,N_5581);
or U6669 (N_6669,N_5199,N_5503);
and U6670 (N_6670,N_5173,N_5706);
nand U6671 (N_6671,N_5194,N_5542);
and U6672 (N_6672,N_5362,N_5869);
nand U6673 (N_6673,N_5009,N_5594);
or U6674 (N_6674,N_5929,N_5230);
and U6675 (N_6675,N_5996,N_5093);
nand U6676 (N_6676,N_5092,N_5574);
xor U6677 (N_6677,N_5484,N_5036);
or U6678 (N_6678,N_5498,N_5758);
or U6679 (N_6679,N_5612,N_5229);
or U6680 (N_6680,N_5387,N_5073);
or U6681 (N_6681,N_5684,N_5743);
nand U6682 (N_6682,N_5949,N_5162);
nand U6683 (N_6683,N_5034,N_5578);
xnor U6684 (N_6684,N_5781,N_5629);
nand U6685 (N_6685,N_5397,N_5700);
and U6686 (N_6686,N_5118,N_5755);
or U6687 (N_6687,N_5262,N_5102);
nand U6688 (N_6688,N_5241,N_5032);
and U6689 (N_6689,N_5910,N_5673);
or U6690 (N_6690,N_5988,N_5101);
or U6691 (N_6691,N_5064,N_5250);
or U6692 (N_6692,N_5997,N_5676);
nor U6693 (N_6693,N_5220,N_5540);
xnor U6694 (N_6694,N_5090,N_5093);
and U6695 (N_6695,N_5039,N_5172);
nor U6696 (N_6696,N_5808,N_5348);
xnor U6697 (N_6697,N_5762,N_5043);
and U6698 (N_6698,N_5000,N_5588);
nor U6699 (N_6699,N_5557,N_5083);
nand U6700 (N_6700,N_5249,N_5005);
and U6701 (N_6701,N_5218,N_5196);
nor U6702 (N_6702,N_5517,N_5899);
and U6703 (N_6703,N_5907,N_5914);
or U6704 (N_6704,N_5097,N_5619);
or U6705 (N_6705,N_5632,N_5101);
or U6706 (N_6706,N_5850,N_5133);
nor U6707 (N_6707,N_5968,N_5158);
xnor U6708 (N_6708,N_5393,N_5268);
or U6709 (N_6709,N_5343,N_5253);
nand U6710 (N_6710,N_5979,N_5448);
nor U6711 (N_6711,N_5207,N_5248);
or U6712 (N_6712,N_5315,N_5374);
nor U6713 (N_6713,N_5270,N_5189);
and U6714 (N_6714,N_5888,N_5800);
nand U6715 (N_6715,N_5089,N_5738);
xor U6716 (N_6716,N_5312,N_5098);
xor U6717 (N_6717,N_5582,N_5974);
nand U6718 (N_6718,N_5061,N_5088);
and U6719 (N_6719,N_5876,N_5181);
nor U6720 (N_6720,N_5655,N_5554);
or U6721 (N_6721,N_5221,N_5186);
and U6722 (N_6722,N_5833,N_5795);
or U6723 (N_6723,N_5573,N_5270);
nor U6724 (N_6724,N_5085,N_5884);
or U6725 (N_6725,N_5807,N_5666);
nor U6726 (N_6726,N_5366,N_5443);
nor U6727 (N_6727,N_5306,N_5157);
and U6728 (N_6728,N_5091,N_5997);
nor U6729 (N_6729,N_5864,N_5317);
or U6730 (N_6730,N_5429,N_5456);
nand U6731 (N_6731,N_5596,N_5364);
xor U6732 (N_6732,N_5423,N_5911);
xor U6733 (N_6733,N_5927,N_5101);
nor U6734 (N_6734,N_5544,N_5870);
nand U6735 (N_6735,N_5507,N_5453);
nand U6736 (N_6736,N_5628,N_5585);
nor U6737 (N_6737,N_5883,N_5517);
xnor U6738 (N_6738,N_5007,N_5084);
xor U6739 (N_6739,N_5434,N_5461);
nand U6740 (N_6740,N_5020,N_5208);
or U6741 (N_6741,N_5718,N_5898);
xor U6742 (N_6742,N_5226,N_5961);
nand U6743 (N_6743,N_5714,N_5322);
and U6744 (N_6744,N_5152,N_5923);
nand U6745 (N_6745,N_5351,N_5920);
and U6746 (N_6746,N_5830,N_5698);
nor U6747 (N_6747,N_5868,N_5168);
or U6748 (N_6748,N_5571,N_5194);
nand U6749 (N_6749,N_5281,N_5410);
xor U6750 (N_6750,N_5686,N_5860);
nand U6751 (N_6751,N_5013,N_5995);
or U6752 (N_6752,N_5816,N_5364);
and U6753 (N_6753,N_5183,N_5154);
or U6754 (N_6754,N_5193,N_5403);
and U6755 (N_6755,N_5486,N_5329);
or U6756 (N_6756,N_5103,N_5163);
nand U6757 (N_6757,N_5366,N_5301);
and U6758 (N_6758,N_5037,N_5574);
nand U6759 (N_6759,N_5504,N_5186);
xor U6760 (N_6760,N_5385,N_5356);
or U6761 (N_6761,N_5812,N_5097);
nor U6762 (N_6762,N_5359,N_5159);
or U6763 (N_6763,N_5034,N_5949);
or U6764 (N_6764,N_5339,N_5664);
and U6765 (N_6765,N_5821,N_5195);
nand U6766 (N_6766,N_5842,N_5372);
nand U6767 (N_6767,N_5975,N_5911);
nand U6768 (N_6768,N_5884,N_5032);
nor U6769 (N_6769,N_5959,N_5518);
or U6770 (N_6770,N_5791,N_5203);
nor U6771 (N_6771,N_5554,N_5592);
xnor U6772 (N_6772,N_5076,N_5051);
xor U6773 (N_6773,N_5316,N_5007);
or U6774 (N_6774,N_5706,N_5975);
and U6775 (N_6775,N_5805,N_5343);
xor U6776 (N_6776,N_5587,N_5658);
xor U6777 (N_6777,N_5354,N_5843);
or U6778 (N_6778,N_5780,N_5903);
nand U6779 (N_6779,N_5785,N_5869);
nor U6780 (N_6780,N_5025,N_5320);
nand U6781 (N_6781,N_5820,N_5386);
nor U6782 (N_6782,N_5429,N_5579);
and U6783 (N_6783,N_5148,N_5535);
xor U6784 (N_6784,N_5763,N_5299);
nand U6785 (N_6785,N_5267,N_5754);
or U6786 (N_6786,N_5178,N_5563);
or U6787 (N_6787,N_5287,N_5616);
and U6788 (N_6788,N_5256,N_5636);
and U6789 (N_6789,N_5685,N_5081);
nor U6790 (N_6790,N_5305,N_5868);
nand U6791 (N_6791,N_5008,N_5539);
or U6792 (N_6792,N_5272,N_5590);
nand U6793 (N_6793,N_5581,N_5929);
or U6794 (N_6794,N_5022,N_5210);
nor U6795 (N_6795,N_5037,N_5036);
and U6796 (N_6796,N_5920,N_5795);
and U6797 (N_6797,N_5426,N_5147);
or U6798 (N_6798,N_5029,N_5201);
or U6799 (N_6799,N_5187,N_5180);
and U6800 (N_6800,N_5412,N_5693);
or U6801 (N_6801,N_5081,N_5699);
and U6802 (N_6802,N_5488,N_5769);
nand U6803 (N_6803,N_5166,N_5264);
and U6804 (N_6804,N_5114,N_5486);
xor U6805 (N_6805,N_5791,N_5073);
nand U6806 (N_6806,N_5155,N_5137);
and U6807 (N_6807,N_5208,N_5366);
nor U6808 (N_6808,N_5054,N_5641);
and U6809 (N_6809,N_5279,N_5118);
nand U6810 (N_6810,N_5072,N_5716);
and U6811 (N_6811,N_5605,N_5278);
or U6812 (N_6812,N_5410,N_5671);
or U6813 (N_6813,N_5867,N_5484);
nand U6814 (N_6814,N_5805,N_5947);
xnor U6815 (N_6815,N_5525,N_5644);
or U6816 (N_6816,N_5723,N_5219);
xor U6817 (N_6817,N_5841,N_5446);
xnor U6818 (N_6818,N_5889,N_5068);
xor U6819 (N_6819,N_5501,N_5222);
nor U6820 (N_6820,N_5299,N_5877);
nor U6821 (N_6821,N_5530,N_5105);
nor U6822 (N_6822,N_5457,N_5705);
xor U6823 (N_6823,N_5041,N_5748);
xor U6824 (N_6824,N_5758,N_5846);
or U6825 (N_6825,N_5592,N_5211);
nor U6826 (N_6826,N_5583,N_5428);
nor U6827 (N_6827,N_5421,N_5603);
nor U6828 (N_6828,N_5218,N_5970);
nand U6829 (N_6829,N_5301,N_5774);
nand U6830 (N_6830,N_5852,N_5166);
and U6831 (N_6831,N_5888,N_5621);
nand U6832 (N_6832,N_5816,N_5509);
and U6833 (N_6833,N_5639,N_5222);
xnor U6834 (N_6834,N_5904,N_5823);
nor U6835 (N_6835,N_5043,N_5920);
nand U6836 (N_6836,N_5908,N_5466);
nand U6837 (N_6837,N_5338,N_5815);
nand U6838 (N_6838,N_5091,N_5216);
xor U6839 (N_6839,N_5382,N_5870);
or U6840 (N_6840,N_5548,N_5241);
and U6841 (N_6841,N_5243,N_5904);
or U6842 (N_6842,N_5112,N_5379);
nor U6843 (N_6843,N_5629,N_5779);
nand U6844 (N_6844,N_5656,N_5691);
nor U6845 (N_6845,N_5744,N_5254);
xnor U6846 (N_6846,N_5178,N_5920);
and U6847 (N_6847,N_5546,N_5960);
nand U6848 (N_6848,N_5535,N_5394);
or U6849 (N_6849,N_5909,N_5972);
nand U6850 (N_6850,N_5430,N_5371);
xnor U6851 (N_6851,N_5091,N_5948);
or U6852 (N_6852,N_5518,N_5626);
xnor U6853 (N_6853,N_5241,N_5372);
nand U6854 (N_6854,N_5924,N_5477);
nor U6855 (N_6855,N_5752,N_5076);
or U6856 (N_6856,N_5397,N_5942);
nor U6857 (N_6857,N_5951,N_5204);
nand U6858 (N_6858,N_5885,N_5429);
xor U6859 (N_6859,N_5460,N_5194);
nor U6860 (N_6860,N_5855,N_5813);
nor U6861 (N_6861,N_5673,N_5091);
xnor U6862 (N_6862,N_5474,N_5941);
xor U6863 (N_6863,N_5247,N_5733);
or U6864 (N_6864,N_5705,N_5830);
and U6865 (N_6865,N_5398,N_5188);
or U6866 (N_6866,N_5247,N_5829);
or U6867 (N_6867,N_5862,N_5577);
or U6868 (N_6868,N_5855,N_5920);
or U6869 (N_6869,N_5125,N_5359);
xor U6870 (N_6870,N_5509,N_5932);
and U6871 (N_6871,N_5561,N_5452);
nand U6872 (N_6872,N_5013,N_5033);
and U6873 (N_6873,N_5366,N_5374);
and U6874 (N_6874,N_5871,N_5726);
nor U6875 (N_6875,N_5021,N_5952);
or U6876 (N_6876,N_5938,N_5494);
xnor U6877 (N_6877,N_5007,N_5982);
nor U6878 (N_6878,N_5149,N_5525);
nor U6879 (N_6879,N_5557,N_5972);
xnor U6880 (N_6880,N_5935,N_5919);
nor U6881 (N_6881,N_5700,N_5145);
nand U6882 (N_6882,N_5527,N_5529);
nand U6883 (N_6883,N_5786,N_5432);
and U6884 (N_6884,N_5405,N_5459);
and U6885 (N_6885,N_5734,N_5322);
xor U6886 (N_6886,N_5200,N_5440);
and U6887 (N_6887,N_5750,N_5998);
or U6888 (N_6888,N_5091,N_5620);
xor U6889 (N_6889,N_5268,N_5396);
or U6890 (N_6890,N_5019,N_5557);
nand U6891 (N_6891,N_5400,N_5214);
and U6892 (N_6892,N_5391,N_5992);
xor U6893 (N_6893,N_5211,N_5980);
or U6894 (N_6894,N_5410,N_5919);
nand U6895 (N_6895,N_5432,N_5695);
or U6896 (N_6896,N_5537,N_5808);
xnor U6897 (N_6897,N_5718,N_5435);
nand U6898 (N_6898,N_5779,N_5787);
nor U6899 (N_6899,N_5484,N_5516);
nand U6900 (N_6900,N_5561,N_5027);
or U6901 (N_6901,N_5039,N_5482);
and U6902 (N_6902,N_5072,N_5001);
nor U6903 (N_6903,N_5324,N_5136);
xor U6904 (N_6904,N_5043,N_5509);
xnor U6905 (N_6905,N_5068,N_5954);
and U6906 (N_6906,N_5281,N_5290);
xnor U6907 (N_6907,N_5485,N_5681);
xor U6908 (N_6908,N_5189,N_5039);
or U6909 (N_6909,N_5303,N_5719);
and U6910 (N_6910,N_5676,N_5937);
nor U6911 (N_6911,N_5125,N_5647);
nand U6912 (N_6912,N_5929,N_5577);
and U6913 (N_6913,N_5068,N_5498);
and U6914 (N_6914,N_5846,N_5941);
and U6915 (N_6915,N_5755,N_5313);
nand U6916 (N_6916,N_5039,N_5942);
and U6917 (N_6917,N_5721,N_5777);
nor U6918 (N_6918,N_5494,N_5157);
xor U6919 (N_6919,N_5616,N_5232);
nor U6920 (N_6920,N_5053,N_5293);
xor U6921 (N_6921,N_5950,N_5507);
nor U6922 (N_6922,N_5566,N_5218);
nand U6923 (N_6923,N_5322,N_5603);
or U6924 (N_6924,N_5518,N_5194);
xnor U6925 (N_6925,N_5688,N_5726);
nor U6926 (N_6926,N_5338,N_5988);
nand U6927 (N_6927,N_5630,N_5487);
nor U6928 (N_6928,N_5779,N_5581);
xor U6929 (N_6929,N_5510,N_5317);
or U6930 (N_6930,N_5176,N_5893);
nand U6931 (N_6931,N_5121,N_5510);
or U6932 (N_6932,N_5799,N_5858);
and U6933 (N_6933,N_5574,N_5056);
and U6934 (N_6934,N_5669,N_5315);
and U6935 (N_6935,N_5282,N_5437);
nor U6936 (N_6936,N_5075,N_5272);
and U6937 (N_6937,N_5702,N_5754);
or U6938 (N_6938,N_5956,N_5562);
nor U6939 (N_6939,N_5277,N_5791);
and U6940 (N_6940,N_5607,N_5170);
nand U6941 (N_6941,N_5465,N_5047);
nor U6942 (N_6942,N_5433,N_5301);
or U6943 (N_6943,N_5818,N_5964);
nor U6944 (N_6944,N_5023,N_5611);
and U6945 (N_6945,N_5941,N_5953);
and U6946 (N_6946,N_5256,N_5378);
and U6947 (N_6947,N_5491,N_5021);
xnor U6948 (N_6948,N_5906,N_5444);
xnor U6949 (N_6949,N_5512,N_5864);
xor U6950 (N_6950,N_5833,N_5964);
and U6951 (N_6951,N_5881,N_5696);
xor U6952 (N_6952,N_5244,N_5606);
and U6953 (N_6953,N_5602,N_5807);
xor U6954 (N_6954,N_5612,N_5134);
and U6955 (N_6955,N_5265,N_5098);
xnor U6956 (N_6956,N_5025,N_5383);
and U6957 (N_6957,N_5608,N_5116);
and U6958 (N_6958,N_5533,N_5362);
nor U6959 (N_6959,N_5564,N_5834);
and U6960 (N_6960,N_5453,N_5929);
and U6961 (N_6961,N_5961,N_5583);
xnor U6962 (N_6962,N_5455,N_5496);
nor U6963 (N_6963,N_5428,N_5818);
nor U6964 (N_6964,N_5915,N_5637);
nand U6965 (N_6965,N_5904,N_5283);
xnor U6966 (N_6966,N_5673,N_5077);
xnor U6967 (N_6967,N_5776,N_5105);
and U6968 (N_6968,N_5100,N_5008);
nor U6969 (N_6969,N_5620,N_5073);
and U6970 (N_6970,N_5841,N_5449);
or U6971 (N_6971,N_5404,N_5104);
nor U6972 (N_6972,N_5670,N_5044);
nand U6973 (N_6973,N_5488,N_5126);
and U6974 (N_6974,N_5408,N_5154);
nand U6975 (N_6975,N_5579,N_5982);
nor U6976 (N_6976,N_5308,N_5863);
xor U6977 (N_6977,N_5965,N_5079);
nor U6978 (N_6978,N_5727,N_5894);
xor U6979 (N_6979,N_5999,N_5092);
or U6980 (N_6980,N_5864,N_5306);
xor U6981 (N_6981,N_5173,N_5103);
or U6982 (N_6982,N_5064,N_5133);
or U6983 (N_6983,N_5824,N_5023);
nand U6984 (N_6984,N_5659,N_5911);
nor U6985 (N_6985,N_5970,N_5401);
and U6986 (N_6986,N_5315,N_5085);
and U6987 (N_6987,N_5773,N_5291);
or U6988 (N_6988,N_5162,N_5611);
nand U6989 (N_6989,N_5877,N_5318);
and U6990 (N_6990,N_5197,N_5238);
nand U6991 (N_6991,N_5609,N_5498);
xnor U6992 (N_6992,N_5622,N_5117);
xnor U6993 (N_6993,N_5013,N_5411);
and U6994 (N_6994,N_5174,N_5446);
and U6995 (N_6995,N_5509,N_5774);
nand U6996 (N_6996,N_5839,N_5233);
nand U6997 (N_6997,N_5419,N_5905);
or U6998 (N_6998,N_5878,N_5179);
and U6999 (N_6999,N_5439,N_5181);
and U7000 (N_7000,N_6216,N_6988);
or U7001 (N_7001,N_6624,N_6153);
nor U7002 (N_7002,N_6774,N_6525);
nor U7003 (N_7003,N_6682,N_6690);
xnor U7004 (N_7004,N_6821,N_6009);
nand U7005 (N_7005,N_6407,N_6401);
xor U7006 (N_7006,N_6882,N_6843);
xnor U7007 (N_7007,N_6379,N_6274);
nand U7008 (N_7008,N_6116,N_6177);
and U7009 (N_7009,N_6260,N_6822);
or U7010 (N_7010,N_6374,N_6916);
or U7011 (N_7011,N_6780,N_6669);
nand U7012 (N_7012,N_6458,N_6312);
nand U7013 (N_7013,N_6889,N_6434);
and U7014 (N_7014,N_6880,N_6508);
xnor U7015 (N_7015,N_6006,N_6213);
nor U7016 (N_7016,N_6787,N_6511);
and U7017 (N_7017,N_6278,N_6926);
nor U7018 (N_7018,N_6048,N_6777);
or U7019 (N_7019,N_6020,N_6903);
nand U7020 (N_7020,N_6380,N_6874);
xnor U7021 (N_7021,N_6793,N_6686);
or U7022 (N_7022,N_6151,N_6581);
or U7023 (N_7023,N_6107,N_6616);
nor U7024 (N_7024,N_6991,N_6764);
xor U7025 (N_7025,N_6681,N_6322);
or U7026 (N_7026,N_6363,N_6655);
nand U7027 (N_7027,N_6255,N_6629);
xor U7028 (N_7028,N_6329,N_6314);
and U7029 (N_7029,N_6394,N_6258);
nand U7030 (N_7030,N_6659,N_6931);
and U7031 (N_7031,N_6033,N_6792);
and U7032 (N_7032,N_6077,N_6014);
and U7033 (N_7033,N_6444,N_6289);
xor U7034 (N_7034,N_6190,N_6085);
xnor U7035 (N_7035,N_6310,N_6680);
nor U7036 (N_7036,N_6735,N_6226);
nor U7037 (N_7037,N_6097,N_6593);
nor U7038 (N_7038,N_6157,N_6052);
and U7039 (N_7039,N_6248,N_6356);
nor U7040 (N_7040,N_6575,N_6744);
xor U7041 (N_7041,N_6221,N_6202);
nor U7042 (N_7042,N_6058,N_6553);
xnor U7043 (N_7043,N_6638,N_6142);
and U7044 (N_7044,N_6748,N_6244);
or U7045 (N_7045,N_6045,N_6555);
nand U7046 (N_7046,N_6257,N_6209);
and U7047 (N_7047,N_6261,N_6080);
and U7048 (N_7048,N_6711,N_6715);
xor U7049 (N_7049,N_6489,N_6622);
and U7050 (N_7050,N_6670,N_6129);
nand U7051 (N_7051,N_6073,N_6398);
and U7052 (N_7052,N_6658,N_6105);
nand U7053 (N_7053,N_6873,N_6164);
nand U7054 (N_7054,N_6396,N_6038);
xnor U7055 (N_7055,N_6527,N_6950);
or U7056 (N_7056,N_6013,N_6666);
nor U7057 (N_7057,N_6391,N_6371);
or U7058 (N_7058,N_6280,N_6929);
nand U7059 (N_7059,N_6617,N_6357);
and U7060 (N_7060,N_6090,N_6019);
and U7061 (N_7061,N_6850,N_6640);
nor U7062 (N_7062,N_6533,N_6932);
xor U7063 (N_7063,N_6016,N_6698);
xnor U7064 (N_7064,N_6072,N_6369);
and U7065 (N_7065,N_6896,N_6423);
or U7066 (N_7066,N_6302,N_6942);
nand U7067 (N_7067,N_6361,N_6187);
nor U7068 (N_7068,N_6217,N_6778);
xnor U7069 (N_7069,N_6567,N_6246);
nand U7070 (N_7070,N_6951,N_6225);
xnor U7071 (N_7071,N_6566,N_6456);
and U7072 (N_7072,N_6119,N_6952);
and U7073 (N_7073,N_6347,N_6413);
or U7074 (N_7074,N_6293,N_6849);
and U7075 (N_7075,N_6124,N_6415);
nand U7076 (N_7076,N_6721,N_6879);
xor U7077 (N_7077,N_6471,N_6049);
nand U7078 (N_7078,N_6832,N_6806);
and U7079 (N_7079,N_6002,N_6776);
nand U7080 (N_7080,N_6061,N_6336);
or U7081 (N_7081,N_6410,N_6986);
xnor U7082 (N_7082,N_6166,N_6488);
nor U7083 (N_7083,N_6234,N_6265);
xnor U7084 (N_7084,N_6355,N_6925);
xnor U7085 (N_7085,N_6263,N_6718);
and U7086 (N_7086,N_6344,N_6325);
or U7087 (N_7087,N_6276,N_6192);
or U7088 (N_7088,N_6240,N_6892);
xnor U7089 (N_7089,N_6865,N_6397);
xor U7090 (N_7090,N_6102,N_6904);
nand U7091 (N_7091,N_6037,N_6341);
and U7092 (N_7092,N_6271,N_6877);
and U7093 (N_7093,N_6936,N_6803);
and U7094 (N_7094,N_6883,N_6043);
xor U7095 (N_7095,N_6921,N_6333);
xor U7096 (N_7096,N_6633,N_6165);
xor U7097 (N_7097,N_6494,N_6007);
nand U7098 (N_7098,N_6156,N_6436);
xor U7099 (N_7099,N_6122,N_6772);
nor U7100 (N_7100,N_6027,N_6709);
nand U7101 (N_7101,N_6411,N_6685);
xor U7102 (N_7102,N_6501,N_6502);
nor U7103 (N_7103,N_6684,N_6961);
or U7104 (N_7104,N_6219,N_6580);
xor U7105 (N_7105,N_6449,N_6392);
or U7106 (N_7106,N_6702,N_6220);
nand U7107 (N_7107,N_6466,N_6955);
nor U7108 (N_7108,N_6717,N_6439);
nor U7109 (N_7109,N_6180,N_6370);
or U7110 (N_7110,N_6453,N_6826);
and U7111 (N_7111,N_6734,N_6573);
or U7112 (N_7112,N_6464,N_6656);
nand U7113 (N_7113,N_6830,N_6603);
nand U7114 (N_7114,N_6938,N_6706);
nor U7115 (N_7115,N_6982,N_6763);
nor U7116 (N_7116,N_6040,N_6492);
xor U7117 (N_7117,N_6923,N_6206);
nand U7118 (N_7118,N_6163,N_6661);
xor U7119 (N_7119,N_6330,N_6383);
nand U7120 (N_7120,N_6095,N_6476);
or U7121 (N_7121,N_6798,N_6340);
nand U7122 (N_7122,N_6524,N_6848);
nand U7123 (N_7123,N_6055,N_6389);
nor U7124 (N_7124,N_6677,N_6704);
nand U7125 (N_7125,N_6059,N_6399);
and U7126 (N_7126,N_6403,N_6412);
or U7127 (N_7127,N_6065,N_6765);
nand U7128 (N_7128,N_6599,N_6132);
and U7129 (N_7129,N_6388,N_6611);
nor U7130 (N_7130,N_6429,N_6993);
and U7131 (N_7131,N_6239,N_6420);
xnor U7132 (N_7132,N_6900,N_6868);
xor U7133 (N_7133,N_6762,N_6922);
nor U7134 (N_7134,N_6432,N_6249);
xnor U7135 (N_7135,N_6319,N_6044);
xor U7136 (N_7136,N_6247,N_6195);
and U7137 (N_7137,N_6967,N_6521);
nand U7138 (N_7138,N_6859,N_6724);
or U7139 (N_7139,N_6651,N_6558);
and U7140 (N_7140,N_6468,N_6948);
nand U7141 (N_7141,N_6784,N_6997);
and U7142 (N_7142,N_6625,N_6299);
xnor U7143 (N_7143,N_6446,N_6409);
nor U7144 (N_7144,N_6954,N_6242);
nand U7145 (N_7145,N_6005,N_6963);
nor U7146 (N_7146,N_6920,N_6106);
nor U7147 (N_7147,N_6548,N_6632);
and U7148 (N_7148,N_6649,N_6816);
nor U7149 (N_7149,N_6838,N_6086);
nand U7150 (N_7150,N_6496,N_6979);
xor U7151 (N_7151,N_6245,N_6876);
nor U7152 (N_7152,N_6123,N_6770);
nor U7153 (N_7153,N_6985,N_6585);
or U7154 (N_7154,N_6968,N_6243);
or U7155 (N_7155,N_6273,N_6384);
or U7156 (N_7156,N_6750,N_6545);
nor U7157 (N_7157,N_6079,N_6256);
xor U7158 (N_7158,N_6214,N_6550);
and U7159 (N_7159,N_6001,N_6634);
xor U7160 (N_7160,N_6918,N_6224);
or U7161 (N_7161,N_6154,N_6886);
nor U7162 (N_7162,N_6069,N_6066);
xnor U7163 (N_7163,N_6729,N_6189);
xnor U7164 (N_7164,N_6976,N_6109);
or U7165 (N_7165,N_6506,N_6168);
nand U7166 (N_7166,N_6200,N_6732);
nand U7167 (N_7167,N_6707,N_6099);
or U7168 (N_7168,N_6373,N_6474);
nand U7169 (N_7169,N_6408,N_6746);
xor U7170 (N_7170,N_6455,N_6120);
nand U7171 (N_7171,N_6913,N_6212);
and U7172 (N_7172,N_6771,N_6056);
nor U7173 (N_7173,N_6930,N_6198);
nor U7174 (N_7174,N_6435,N_6962);
or U7175 (N_7175,N_6939,N_6463);
or U7176 (N_7176,N_6554,N_6515);
nand U7177 (N_7177,N_6811,N_6440);
and U7178 (N_7178,N_6825,N_6068);
and U7179 (N_7179,N_6133,N_6313);
nor U7180 (N_7180,N_6775,N_6783);
nand U7181 (N_7181,N_6687,N_6927);
and U7182 (N_7182,N_6241,N_6761);
nor U7183 (N_7183,N_6691,N_6676);
nor U7184 (N_7184,N_6740,N_6606);
nor U7185 (N_7185,N_6473,N_6644);
xor U7186 (N_7186,N_6688,N_6251);
nand U7187 (N_7187,N_6737,N_6141);
or U7188 (N_7188,N_6703,N_6710);
or U7189 (N_7189,N_6531,N_6499);
or U7190 (N_7190,N_6509,N_6098);
xor U7191 (N_7191,N_6878,N_6364);
nand U7192 (N_7192,N_6884,N_6089);
xor U7193 (N_7193,N_6812,N_6532);
nor U7194 (N_7194,N_6957,N_6117);
nor U7195 (N_7195,N_6025,N_6281);
nand U7196 (N_7196,N_6268,N_6990);
and U7197 (N_7197,N_6570,N_6722);
nand U7198 (N_7198,N_6568,N_6094);
nand U7199 (N_7199,N_6262,N_6478);
nand U7200 (N_7200,N_6272,N_6201);
nand U7201 (N_7201,N_6945,N_6084);
or U7202 (N_7202,N_6238,N_6529);
nor U7203 (N_7203,N_6184,N_6155);
or U7204 (N_7204,N_6088,N_6287);
xor U7205 (N_7205,N_6022,N_6317);
nand U7206 (N_7206,N_6186,N_6510);
xor U7207 (N_7207,N_6395,N_6442);
or U7208 (N_7208,N_6375,N_6070);
or U7209 (N_7209,N_6181,N_6078);
or U7210 (N_7210,N_6730,N_6110);
nand U7211 (N_7211,N_6600,N_6414);
xnor U7212 (N_7212,N_6801,N_6888);
or U7213 (N_7213,N_6259,N_6517);
xnor U7214 (N_7214,N_6614,N_6911);
and U7215 (N_7215,N_6588,N_6191);
nand U7216 (N_7216,N_6311,N_6475);
xnor U7217 (N_7217,N_6067,N_6026);
or U7218 (N_7218,N_6528,N_6004);
and U7219 (N_7219,N_6326,N_6618);
nor U7220 (N_7220,N_6030,N_6743);
or U7221 (N_7221,N_6572,N_6895);
nand U7222 (N_7222,N_6814,N_6577);
nand U7223 (N_7223,N_6233,N_6958);
and U7224 (N_7224,N_6091,N_6790);
xnor U7225 (N_7225,N_6269,N_6108);
or U7226 (N_7226,N_6791,N_6467);
nor U7227 (N_7227,N_6665,N_6788);
or U7228 (N_7228,N_6867,N_6021);
nand U7229 (N_7229,N_6254,N_6708);
xor U7230 (N_7230,N_6893,N_6586);
nor U7231 (N_7231,N_6779,N_6796);
nor U7232 (N_7232,N_6980,N_6881);
xor U7233 (N_7233,N_6320,N_6235);
or U7234 (N_7234,N_6683,N_6060);
nand U7235 (N_7235,N_6228,N_6368);
and U7236 (N_7236,N_6047,N_6470);
nor U7237 (N_7237,N_6689,N_6343);
and U7238 (N_7238,N_6978,N_6653);
nor U7239 (N_7239,N_6654,N_6479);
and U7240 (N_7240,N_6359,N_6785);
or U7241 (N_7241,N_6844,N_6457);
xor U7242 (N_7242,N_6114,N_6137);
nand U7243 (N_7243,N_6753,N_6424);
or U7244 (N_7244,N_6719,N_6188);
nor U7245 (N_7245,N_6053,N_6367);
xnor U7246 (N_7246,N_6174,N_6899);
nor U7247 (N_7247,N_6348,N_6824);
or U7248 (N_7248,N_6933,N_6767);
nor U7249 (N_7249,N_6615,N_6998);
nor U7250 (N_7250,N_6973,N_6802);
and U7251 (N_7251,N_6366,N_6300);
nand U7252 (N_7252,N_6747,N_6643);
nor U7253 (N_7253,N_6549,N_6196);
nor U7254 (N_7254,N_6076,N_6754);
nor U7255 (N_7255,N_6134,N_6335);
xnor U7256 (N_7256,N_6178,N_6840);
and U7257 (N_7257,N_6530,N_6378);
and U7258 (N_7258,N_6605,N_6277);
or U7259 (N_7259,N_6041,N_6639);
nor U7260 (N_7260,N_6342,N_6182);
xnor U7261 (N_7261,N_6716,N_6935);
nand U7262 (N_7262,N_6820,N_6046);
nor U7263 (N_7263,N_6578,N_6267);
or U7264 (N_7264,N_6306,N_6286);
or U7265 (N_7265,N_6204,N_6619);
nand U7266 (N_7266,N_6063,N_6620);
and U7267 (N_7267,N_6159,N_6769);
xor U7268 (N_7268,N_6175,N_6284);
and U7269 (N_7269,N_6146,N_6885);
xor U7270 (N_7270,N_6327,N_6294);
nor U7271 (N_7271,N_6766,N_6839);
or U7272 (N_7272,N_6742,N_6352);
and U7273 (N_7273,N_6773,N_6081);
and U7274 (N_7274,N_6828,N_6660);
and U7275 (N_7275,N_6346,N_6890);
or U7276 (N_7276,N_6183,N_6334);
and U7277 (N_7277,N_6128,N_6757);
nand U7278 (N_7278,N_6984,N_6662);
nand U7279 (N_7279,N_6297,N_6516);
nor U7280 (N_7280,N_6836,N_6008);
xor U7281 (N_7281,N_6694,N_6800);
nor U7282 (N_7282,N_6668,N_6050);
xor U7283 (N_7283,N_6908,N_6140);
nand U7284 (N_7284,N_6387,N_6862);
nand U7285 (N_7285,N_6914,N_6970);
xor U7286 (N_7286,N_6635,N_6738);
xor U7287 (N_7287,N_6485,N_6894);
nand U7288 (N_7288,N_6641,N_6860);
nand U7289 (N_7289,N_6111,N_6768);
or U7290 (N_7290,N_6152,N_6941);
or U7291 (N_7291,N_6460,N_6833);
and U7292 (N_7292,N_6372,N_6465);
nor U7293 (N_7293,N_6237,N_6318);
nor U7294 (N_7294,N_6115,N_6520);
nor U7295 (N_7295,N_6541,N_6934);
and U7296 (N_7296,N_6835,N_6514);
nand U7297 (N_7297,N_6275,N_6127);
and U7298 (N_7298,N_6584,N_6810);
and U7299 (N_7299,N_6418,N_6917);
and U7300 (N_7300,N_6544,N_6331);
nand U7301 (N_7301,N_6171,N_6569);
xor U7302 (N_7302,N_6571,N_6760);
nand U7303 (N_7303,N_6697,N_6448);
or U7304 (N_7304,N_6552,N_6621);
xnor U7305 (N_7305,N_6345,N_6282);
nand U7306 (N_7306,N_6087,N_6113);
or U7307 (N_7307,N_6207,N_6487);
xnor U7308 (N_7308,N_6491,N_6462);
nor U7309 (N_7309,N_6504,N_6288);
and U7310 (N_7310,N_6960,N_6304);
and U7311 (N_7311,N_6270,N_6279);
nor U7312 (N_7312,N_6583,N_6169);
nand U7313 (N_7313,N_6559,N_6445);
nor U7314 (N_7314,N_6587,N_6875);
nor U7315 (N_7315,N_6185,N_6869);
nor U7316 (N_7316,N_6406,N_6992);
xnor U7317 (N_7317,N_6574,N_6675);
xor U7318 (N_7318,N_6227,N_6323);
or U7319 (N_7319,N_6292,N_6562);
and U7320 (N_7320,N_6536,N_6236);
nor U7321 (N_7321,N_6498,N_6560);
or U7322 (N_7322,N_6147,N_6362);
nor U7323 (N_7323,N_6136,N_6351);
nand U7324 (N_7324,N_6609,N_6266);
nand U7325 (N_7325,N_6402,N_6781);
nand U7326 (N_7326,N_6598,N_6540);
xnor U7327 (N_7327,N_6608,N_6438);
and U7328 (N_7328,N_6645,N_6430);
nand U7329 (N_7329,N_6752,N_6664);
nand U7330 (N_7330,N_6173,N_6607);
or U7331 (N_7331,N_6349,N_6546);
or U7332 (N_7332,N_6104,N_6493);
nor U7333 (N_7333,N_6425,N_6461);
and U7334 (N_7334,N_6199,N_6477);
nor U7335 (N_7335,N_6321,N_6017);
nor U7336 (N_7336,N_6695,N_6138);
nand U7337 (N_7337,N_6483,N_6229);
and U7338 (N_7338,N_6901,N_6029);
nor U7339 (N_7339,N_6995,N_6328);
and U7340 (N_7340,N_6543,N_6906);
nor U7341 (N_7341,N_6308,N_6969);
or U7342 (N_7342,N_6112,N_6035);
or U7343 (N_7343,N_6381,N_6039);
xnor U7344 (N_7344,N_6999,N_6845);
nor U7345 (N_7345,N_6135,N_6427);
and U7346 (N_7346,N_6160,N_6481);
or U7347 (N_7347,N_6179,N_6145);
and U7348 (N_7348,N_6720,N_6861);
nor U7349 (N_7349,N_6829,N_6539);
nor U7350 (N_7350,N_6672,N_6628);
nor U7351 (N_7351,N_6994,N_6512);
and U7352 (N_7352,N_6563,N_6853);
nand U7353 (N_7353,N_6139,N_6441);
xnor U7354 (N_7354,N_6291,N_6513);
nor U7355 (N_7355,N_6071,N_6852);
nand U7356 (N_7356,N_6534,N_6851);
and U7357 (N_7357,N_6360,N_6338);
or U7358 (N_7358,N_6647,N_6426);
nor U7359 (N_7359,N_6981,N_6428);
xor U7360 (N_7360,N_6795,N_6484);
or U7361 (N_7361,N_6551,N_6597);
or U7362 (N_7362,N_6222,N_6285);
xnor U7363 (N_7363,N_6400,N_6290);
or U7364 (N_7364,N_6472,N_6096);
nor U7365 (N_7365,N_6674,N_6696);
nand U7366 (N_7366,N_6393,N_6579);
nor U7367 (N_7367,N_6758,N_6522);
and U7368 (N_7368,N_6149,N_6699);
nand U7369 (N_7369,N_6443,N_6459);
or U7370 (N_7370,N_6405,N_6714);
nor U7371 (N_7371,N_6057,N_6648);
xnor U7372 (N_7372,N_6121,N_6054);
or U7373 (N_7373,N_6870,N_6382);
and U7374 (N_7374,N_6556,N_6203);
and U7375 (N_7375,N_6834,N_6871);
and U7376 (N_7376,N_6042,N_6943);
nand U7377 (N_7377,N_6678,N_6032);
xor U7378 (N_7378,N_6503,N_6975);
xnor U7379 (N_7379,N_6637,N_6486);
nor U7380 (N_7380,N_6819,N_6416);
and U7381 (N_7381,N_6167,N_6592);
nor U7382 (N_7382,N_6526,N_6725);
nand U7383 (N_7383,N_6799,N_6495);
xnor U7384 (N_7384,N_6944,N_6947);
or U7385 (N_7385,N_6673,N_6910);
and U7386 (N_7386,N_6626,N_6417);
nand U7387 (N_7387,N_6339,N_6846);
xor U7388 (N_7388,N_6211,N_6295);
nand U7389 (N_7389,N_6612,N_6028);
xor U7390 (N_7390,N_6193,N_6176);
nor U7391 (N_7391,N_6296,N_6101);
nor U7392 (N_7392,N_6505,N_6253);
or U7393 (N_7393,N_6298,N_6162);
nor U7394 (N_7394,N_6727,N_6807);
and U7395 (N_7395,N_6497,N_6010);
xor U7396 (N_7396,N_6898,N_6602);
nand U7397 (N_7397,N_6723,N_6928);
and U7398 (N_7398,N_6130,N_6949);
nor U7399 (N_7399,N_6959,N_6646);
or U7400 (N_7400,N_6582,N_6301);
xor U7401 (N_7401,N_6051,N_6808);
xnor U7402 (N_7402,N_6858,N_6977);
nor U7403 (N_7403,N_6946,N_6663);
nor U7404 (N_7404,N_6856,N_6604);
and U7405 (N_7405,N_6897,N_6671);
xnor U7406 (N_7406,N_6011,N_6857);
and U7407 (N_7407,N_6631,N_6837);
nand U7408 (N_7408,N_6657,N_6500);
xnor U7409 (N_7409,N_6194,N_6789);
and U7410 (N_7410,N_6170,N_6376);
and U7411 (N_7411,N_6422,N_6636);
and U7412 (N_7412,N_6855,N_6118);
and U7413 (N_7413,N_6842,N_6018);
or U7414 (N_7414,N_6751,N_6786);
and U7415 (N_7415,N_6891,N_6613);
and U7416 (N_7416,N_6365,N_6252);
xnor U7417 (N_7417,N_6749,N_6082);
nand U7418 (N_7418,N_6452,N_6794);
and U7419 (N_7419,N_6332,N_6755);
nor U7420 (N_7420,N_6797,N_6972);
xnor U7421 (N_7421,N_6215,N_6940);
nor U7422 (N_7422,N_6125,N_6966);
nor U7423 (N_7423,N_6538,N_6523);
nor U7424 (N_7424,N_6827,N_6003);
and U7425 (N_7425,N_6131,N_6953);
nor U7426 (N_7426,N_6823,N_6983);
nor U7427 (N_7427,N_6482,N_6337);
nor U7428 (N_7428,N_6305,N_6887);
nor U7429 (N_7429,N_6358,N_6565);
nor U7430 (N_7430,N_6208,N_6804);
nor U7431 (N_7431,N_6692,N_6863);
nand U7432 (N_7432,N_6907,N_6652);
xnor U7433 (N_7433,N_6283,N_6205);
or U7434 (N_7434,N_6736,N_6700);
nand U7435 (N_7435,N_6385,N_6576);
and U7436 (N_7436,N_6817,N_6012);
or U7437 (N_7437,N_6150,N_6610);
and U7438 (N_7438,N_6447,N_6756);
xor U7439 (N_7439,N_6377,N_6809);
xor U7440 (N_7440,N_6679,N_6507);
xnor U7441 (N_7441,N_6956,N_6596);
xor U7442 (N_7442,N_6728,N_6075);
xor U7443 (N_7443,N_6590,N_6642);
or U7444 (N_7444,N_6143,N_6712);
or U7445 (N_7445,N_6433,N_6595);
nor U7446 (N_7446,N_6739,N_6996);
nor U7447 (N_7447,N_6519,N_6854);
or U7448 (N_7448,N_6542,N_6557);
nor U7449 (N_7449,N_6564,N_6390);
and U7450 (N_7450,N_6036,N_6701);
nand U7451 (N_7451,N_6782,N_6872);
nand U7452 (N_7452,N_6451,N_6223);
or U7453 (N_7453,N_6083,N_6915);
xor U7454 (N_7454,N_6015,N_6103);
or U7455 (N_7455,N_6623,N_6480);
and U7456 (N_7456,N_6264,N_6126);
xor U7457 (N_7457,N_6404,N_6912);
nand U7458 (N_7458,N_6831,N_6594);
nor U7459 (N_7459,N_6431,N_6074);
and U7460 (N_7460,N_6987,N_6547);
or U7461 (N_7461,N_6158,N_6902);
xnor U7462 (N_7462,N_6627,N_6024);
and U7463 (N_7463,N_6232,N_6454);
nor U7464 (N_7464,N_6841,N_6197);
nor U7465 (N_7465,N_6231,N_6210);
and U7466 (N_7466,N_6630,N_6230);
and U7467 (N_7467,N_6353,N_6450);
nor U7468 (N_7468,N_6092,N_6589);
xor U7469 (N_7469,N_6093,N_6805);
nor U7470 (N_7470,N_6726,N_6437);
and U7471 (N_7471,N_6866,N_6535);
and U7472 (N_7472,N_6303,N_6847);
xor U7473 (N_7473,N_6469,N_6815);
nor U7474 (N_7474,N_6419,N_6818);
nand U7475 (N_7475,N_6965,N_6971);
xor U7476 (N_7476,N_6759,N_6741);
xor U7477 (N_7477,N_6144,N_6490);
and U7478 (N_7478,N_6031,N_6350);
and U7479 (N_7479,N_6905,N_6601);
nor U7480 (N_7480,N_6937,N_6315);
and U7481 (N_7481,N_6964,N_6667);
and U7482 (N_7482,N_6421,N_6518);
nor U7483 (N_7483,N_6316,N_6324);
nor U7484 (N_7484,N_6000,N_6693);
nor U7485 (N_7485,N_6537,N_6713);
and U7486 (N_7486,N_6650,N_6561);
and U7487 (N_7487,N_6250,N_6733);
xnor U7488 (N_7488,N_6909,N_6148);
nor U7489 (N_7489,N_6386,N_6974);
xnor U7490 (N_7490,N_6218,N_6023);
nand U7491 (N_7491,N_6924,N_6100);
or U7492 (N_7492,N_6919,N_6034);
or U7493 (N_7493,N_6813,N_6064);
or U7494 (N_7494,N_6989,N_6591);
nor U7495 (N_7495,N_6705,N_6731);
xnor U7496 (N_7496,N_6864,N_6745);
nor U7497 (N_7497,N_6307,N_6172);
nand U7498 (N_7498,N_6161,N_6062);
nor U7499 (N_7499,N_6309,N_6354);
nand U7500 (N_7500,N_6304,N_6674);
xnor U7501 (N_7501,N_6262,N_6382);
or U7502 (N_7502,N_6767,N_6969);
nand U7503 (N_7503,N_6900,N_6861);
nor U7504 (N_7504,N_6648,N_6262);
nand U7505 (N_7505,N_6912,N_6932);
nand U7506 (N_7506,N_6826,N_6491);
and U7507 (N_7507,N_6226,N_6002);
and U7508 (N_7508,N_6039,N_6943);
xor U7509 (N_7509,N_6394,N_6509);
nand U7510 (N_7510,N_6984,N_6492);
nand U7511 (N_7511,N_6698,N_6696);
nand U7512 (N_7512,N_6987,N_6570);
xor U7513 (N_7513,N_6164,N_6415);
and U7514 (N_7514,N_6346,N_6856);
nor U7515 (N_7515,N_6864,N_6475);
and U7516 (N_7516,N_6526,N_6286);
nor U7517 (N_7517,N_6121,N_6918);
xnor U7518 (N_7518,N_6831,N_6029);
and U7519 (N_7519,N_6822,N_6684);
xnor U7520 (N_7520,N_6498,N_6851);
nor U7521 (N_7521,N_6360,N_6453);
nor U7522 (N_7522,N_6333,N_6925);
nor U7523 (N_7523,N_6516,N_6757);
nor U7524 (N_7524,N_6618,N_6976);
xor U7525 (N_7525,N_6017,N_6156);
nor U7526 (N_7526,N_6090,N_6878);
and U7527 (N_7527,N_6716,N_6751);
or U7528 (N_7528,N_6010,N_6007);
xnor U7529 (N_7529,N_6007,N_6342);
xor U7530 (N_7530,N_6752,N_6482);
and U7531 (N_7531,N_6118,N_6852);
nand U7532 (N_7532,N_6844,N_6474);
or U7533 (N_7533,N_6260,N_6645);
nor U7534 (N_7534,N_6996,N_6905);
xor U7535 (N_7535,N_6402,N_6228);
and U7536 (N_7536,N_6630,N_6152);
and U7537 (N_7537,N_6038,N_6137);
nor U7538 (N_7538,N_6472,N_6843);
nand U7539 (N_7539,N_6967,N_6598);
nand U7540 (N_7540,N_6747,N_6745);
nor U7541 (N_7541,N_6781,N_6309);
and U7542 (N_7542,N_6576,N_6750);
nor U7543 (N_7543,N_6057,N_6079);
or U7544 (N_7544,N_6831,N_6339);
xor U7545 (N_7545,N_6802,N_6314);
xnor U7546 (N_7546,N_6762,N_6325);
or U7547 (N_7547,N_6397,N_6375);
nand U7548 (N_7548,N_6746,N_6259);
nor U7549 (N_7549,N_6528,N_6972);
xnor U7550 (N_7550,N_6953,N_6971);
xnor U7551 (N_7551,N_6802,N_6197);
xor U7552 (N_7552,N_6715,N_6788);
xor U7553 (N_7553,N_6949,N_6307);
and U7554 (N_7554,N_6652,N_6279);
nor U7555 (N_7555,N_6876,N_6081);
nand U7556 (N_7556,N_6055,N_6155);
and U7557 (N_7557,N_6385,N_6706);
and U7558 (N_7558,N_6492,N_6647);
nand U7559 (N_7559,N_6149,N_6971);
nand U7560 (N_7560,N_6271,N_6689);
nor U7561 (N_7561,N_6616,N_6035);
nand U7562 (N_7562,N_6243,N_6136);
nor U7563 (N_7563,N_6156,N_6938);
or U7564 (N_7564,N_6332,N_6236);
xor U7565 (N_7565,N_6835,N_6149);
xnor U7566 (N_7566,N_6298,N_6207);
xor U7567 (N_7567,N_6058,N_6313);
xnor U7568 (N_7568,N_6936,N_6601);
nor U7569 (N_7569,N_6890,N_6018);
xor U7570 (N_7570,N_6974,N_6787);
and U7571 (N_7571,N_6924,N_6593);
nor U7572 (N_7572,N_6552,N_6636);
nand U7573 (N_7573,N_6522,N_6025);
or U7574 (N_7574,N_6887,N_6643);
nor U7575 (N_7575,N_6538,N_6054);
and U7576 (N_7576,N_6343,N_6315);
or U7577 (N_7577,N_6288,N_6281);
or U7578 (N_7578,N_6197,N_6224);
or U7579 (N_7579,N_6178,N_6740);
or U7580 (N_7580,N_6756,N_6937);
or U7581 (N_7581,N_6341,N_6647);
xnor U7582 (N_7582,N_6658,N_6218);
and U7583 (N_7583,N_6518,N_6679);
nand U7584 (N_7584,N_6028,N_6615);
xnor U7585 (N_7585,N_6636,N_6957);
nand U7586 (N_7586,N_6197,N_6981);
xor U7587 (N_7587,N_6553,N_6502);
nor U7588 (N_7588,N_6924,N_6975);
and U7589 (N_7589,N_6818,N_6761);
nor U7590 (N_7590,N_6453,N_6825);
or U7591 (N_7591,N_6031,N_6341);
and U7592 (N_7592,N_6659,N_6261);
xor U7593 (N_7593,N_6240,N_6295);
or U7594 (N_7594,N_6466,N_6316);
and U7595 (N_7595,N_6598,N_6050);
nand U7596 (N_7596,N_6453,N_6838);
nand U7597 (N_7597,N_6703,N_6711);
nor U7598 (N_7598,N_6329,N_6210);
or U7599 (N_7599,N_6660,N_6584);
or U7600 (N_7600,N_6241,N_6024);
xnor U7601 (N_7601,N_6183,N_6851);
xor U7602 (N_7602,N_6391,N_6402);
and U7603 (N_7603,N_6235,N_6565);
nand U7604 (N_7604,N_6865,N_6923);
and U7605 (N_7605,N_6887,N_6409);
nor U7606 (N_7606,N_6322,N_6741);
or U7607 (N_7607,N_6460,N_6380);
nor U7608 (N_7608,N_6577,N_6659);
xnor U7609 (N_7609,N_6943,N_6189);
and U7610 (N_7610,N_6129,N_6868);
xnor U7611 (N_7611,N_6764,N_6001);
or U7612 (N_7612,N_6452,N_6976);
nor U7613 (N_7613,N_6764,N_6061);
xnor U7614 (N_7614,N_6076,N_6336);
nor U7615 (N_7615,N_6609,N_6642);
nand U7616 (N_7616,N_6202,N_6010);
nor U7617 (N_7617,N_6514,N_6261);
or U7618 (N_7618,N_6687,N_6587);
and U7619 (N_7619,N_6401,N_6257);
nand U7620 (N_7620,N_6474,N_6104);
nand U7621 (N_7621,N_6958,N_6830);
nor U7622 (N_7622,N_6303,N_6434);
nand U7623 (N_7623,N_6779,N_6981);
or U7624 (N_7624,N_6282,N_6667);
or U7625 (N_7625,N_6698,N_6748);
nand U7626 (N_7626,N_6794,N_6786);
and U7627 (N_7627,N_6139,N_6542);
nor U7628 (N_7628,N_6831,N_6524);
nor U7629 (N_7629,N_6278,N_6343);
xnor U7630 (N_7630,N_6639,N_6391);
and U7631 (N_7631,N_6193,N_6398);
or U7632 (N_7632,N_6770,N_6939);
and U7633 (N_7633,N_6677,N_6060);
or U7634 (N_7634,N_6159,N_6768);
and U7635 (N_7635,N_6460,N_6204);
nand U7636 (N_7636,N_6411,N_6070);
nor U7637 (N_7637,N_6338,N_6000);
nor U7638 (N_7638,N_6021,N_6628);
nand U7639 (N_7639,N_6360,N_6315);
nand U7640 (N_7640,N_6001,N_6067);
and U7641 (N_7641,N_6521,N_6517);
nor U7642 (N_7642,N_6722,N_6141);
nand U7643 (N_7643,N_6342,N_6157);
nand U7644 (N_7644,N_6562,N_6560);
nor U7645 (N_7645,N_6165,N_6046);
nand U7646 (N_7646,N_6738,N_6121);
nor U7647 (N_7647,N_6765,N_6261);
nand U7648 (N_7648,N_6748,N_6573);
and U7649 (N_7649,N_6835,N_6960);
or U7650 (N_7650,N_6391,N_6720);
nand U7651 (N_7651,N_6887,N_6357);
nor U7652 (N_7652,N_6645,N_6916);
and U7653 (N_7653,N_6723,N_6583);
xnor U7654 (N_7654,N_6526,N_6182);
nor U7655 (N_7655,N_6273,N_6471);
and U7656 (N_7656,N_6529,N_6442);
nor U7657 (N_7657,N_6512,N_6444);
or U7658 (N_7658,N_6624,N_6575);
or U7659 (N_7659,N_6972,N_6839);
nor U7660 (N_7660,N_6854,N_6284);
nor U7661 (N_7661,N_6491,N_6084);
xor U7662 (N_7662,N_6750,N_6862);
or U7663 (N_7663,N_6625,N_6534);
or U7664 (N_7664,N_6465,N_6552);
xnor U7665 (N_7665,N_6867,N_6255);
or U7666 (N_7666,N_6748,N_6344);
or U7667 (N_7667,N_6394,N_6634);
or U7668 (N_7668,N_6745,N_6719);
nor U7669 (N_7669,N_6950,N_6836);
and U7670 (N_7670,N_6837,N_6803);
xnor U7671 (N_7671,N_6151,N_6828);
and U7672 (N_7672,N_6000,N_6011);
and U7673 (N_7673,N_6813,N_6414);
and U7674 (N_7674,N_6688,N_6350);
or U7675 (N_7675,N_6841,N_6745);
nand U7676 (N_7676,N_6472,N_6768);
and U7677 (N_7677,N_6528,N_6225);
and U7678 (N_7678,N_6027,N_6869);
xor U7679 (N_7679,N_6774,N_6808);
nor U7680 (N_7680,N_6635,N_6888);
xor U7681 (N_7681,N_6043,N_6451);
xnor U7682 (N_7682,N_6758,N_6321);
or U7683 (N_7683,N_6256,N_6239);
xor U7684 (N_7684,N_6383,N_6398);
nand U7685 (N_7685,N_6113,N_6232);
xnor U7686 (N_7686,N_6637,N_6405);
nor U7687 (N_7687,N_6793,N_6841);
or U7688 (N_7688,N_6799,N_6611);
xor U7689 (N_7689,N_6211,N_6737);
nand U7690 (N_7690,N_6007,N_6328);
xor U7691 (N_7691,N_6330,N_6333);
nor U7692 (N_7692,N_6145,N_6187);
xor U7693 (N_7693,N_6687,N_6301);
nand U7694 (N_7694,N_6379,N_6015);
xnor U7695 (N_7695,N_6578,N_6033);
xnor U7696 (N_7696,N_6005,N_6972);
nand U7697 (N_7697,N_6120,N_6032);
xnor U7698 (N_7698,N_6465,N_6139);
and U7699 (N_7699,N_6200,N_6316);
nor U7700 (N_7700,N_6999,N_6389);
xnor U7701 (N_7701,N_6193,N_6352);
xnor U7702 (N_7702,N_6395,N_6440);
nor U7703 (N_7703,N_6042,N_6072);
and U7704 (N_7704,N_6777,N_6066);
xor U7705 (N_7705,N_6410,N_6201);
and U7706 (N_7706,N_6983,N_6030);
or U7707 (N_7707,N_6308,N_6725);
nor U7708 (N_7708,N_6914,N_6043);
nand U7709 (N_7709,N_6675,N_6532);
nand U7710 (N_7710,N_6332,N_6470);
or U7711 (N_7711,N_6651,N_6798);
nor U7712 (N_7712,N_6274,N_6324);
xor U7713 (N_7713,N_6569,N_6415);
or U7714 (N_7714,N_6722,N_6087);
xor U7715 (N_7715,N_6897,N_6232);
nand U7716 (N_7716,N_6223,N_6356);
nand U7717 (N_7717,N_6288,N_6427);
or U7718 (N_7718,N_6707,N_6190);
xnor U7719 (N_7719,N_6885,N_6967);
xnor U7720 (N_7720,N_6960,N_6288);
nor U7721 (N_7721,N_6186,N_6045);
or U7722 (N_7722,N_6333,N_6430);
or U7723 (N_7723,N_6973,N_6433);
and U7724 (N_7724,N_6556,N_6025);
nand U7725 (N_7725,N_6915,N_6581);
or U7726 (N_7726,N_6648,N_6748);
xnor U7727 (N_7727,N_6430,N_6620);
and U7728 (N_7728,N_6824,N_6541);
xnor U7729 (N_7729,N_6052,N_6571);
nor U7730 (N_7730,N_6209,N_6143);
xnor U7731 (N_7731,N_6072,N_6341);
and U7732 (N_7732,N_6794,N_6433);
nand U7733 (N_7733,N_6576,N_6504);
nor U7734 (N_7734,N_6764,N_6356);
nand U7735 (N_7735,N_6026,N_6507);
or U7736 (N_7736,N_6611,N_6383);
nor U7737 (N_7737,N_6036,N_6578);
xor U7738 (N_7738,N_6346,N_6441);
nor U7739 (N_7739,N_6404,N_6651);
and U7740 (N_7740,N_6499,N_6849);
nor U7741 (N_7741,N_6014,N_6756);
and U7742 (N_7742,N_6270,N_6096);
and U7743 (N_7743,N_6418,N_6767);
or U7744 (N_7744,N_6657,N_6008);
nand U7745 (N_7745,N_6773,N_6186);
and U7746 (N_7746,N_6309,N_6601);
nor U7747 (N_7747,N_6047,N_6579);
or U7748 (N_7748,N_6508,N_6974);
or U7749 (N_7749,N_6414,N_6269);
nand U7750 (N_7750,N_6098,N_6121);
or U7751 (N_7751,N_6047,N_6812);
and U7752 (N_7752,N_6328,N_6047);
xnor U7753 (N_7753,N_6403,N_6964);
nor U7754 (N_7754,N_6810,N_6602);
nand U7755 (N_7755,N_6934,N_6874);
or U7756 (N_7756,N_6332,N_6887);
xor U7757 (N_7757,N_6474,N_6171);
xor U7758 (N_7758,N_6011,N_6279);
xor U7759 (N_7759,N_6155,N_6628);
nand U7760 (N_7760,N_6527,N_6257);
or U7761 (N_7761,N_6552,N_6756);
xnor U7762 (N_7762,N_6726,N_6459);
nor U7763 (N_7763,N_6884,N_6198);
xor U7764 (N_7764,N_6215,N_6800);
nand U7765 (N_7765,N_6113,N_6923);
nand U7766 (N_7766,N_6053,N_6578);
or U7767 (N_7767,N_6184,N_6649);
and U7768 (N_7768,N_6039,N_6675);
nand U7769 (N_7769,N_6226,N_6214);
xor U7770 (N_7770,N_6566,N_6187);
nor U7771 (N_7771,N_6685,N_6083);
and U7772 (N_7772,N_6945,N_6211);
and U7773 (N_7773,N_6581,N_6506);
and U7774 (N_7774,N_6219,N_6868);
xor U7775 (N_7775,N_6579,N_6820);
and U7776 (N_7776,N_6319,N_6051);
or U7777 (N_7777,N_6803,N_6669);
nand U7778 (N_7778,N_6837,N_6594);
or U7779 (N_7779,N_6703,N_6160);
xor U7780 (N_7780,N_6127,N_6398);
or U7781 (N_7781,N_6193,N_6274);
and U7782 (N_7782,N_6130,N_6266);
nor U7783 (N_7783,N_6499,N_6503);
or U7784 (N_7784,N_6911,N_6113);
nand U7785 (N_7785,N_6895,N_6674);
or U7786 (N_7786,N_6311,N_6233);
nand U7787 (N_7787,N_6992,N_6749);
or U7788 (N_7788,N_6559,N_6522);
and U7789 (N_7789,N_6235,N_6939);
nor U7790 (N_7790,N_6245,N_6243);
nand U7791 (N_7791,N_6762,N_6916);
or U7792 (N_7792,N_6214,N_6046);
xor U7793 (N_7793,N_6976,N_6818);
nand U7794 (N_7794,N_6418,N_6199);
nand U7795 (N_7795,N_6915,N_6784);
nor U7796 (N_7796,N_6195,N_6227);
or U7797 (N_7797,N_6526,N_6440);
nor U7798 (N_7798,N_6243,N_6896);
or U7799 (N_7799,N_6192,N_6536);
and U7800 (N_7800,N_6247,N_6425);
nand U7801 (N_7801,N_6135,N_6433);
xor U7802 (N_7802,N_6297,N_6589);
nor U7803 (N_7803,N_6593,N_6361);
and U7804 (N_7804,N_6725,N_6304);
nor U7805 (N_7805,N_6746,N_6883);
nor U7806 (N_7806,N_6835,N_6321);
nand U7807 (N_7807,N_6972,N_6629);
nand U7808 (N_7808,N_6477,N_6038);
or U7809 (N_7809,N_6054,N_6526);
nand U7810 (N_7810,N_6036,N_6032);
and U7811 (N_7811,N_6063,N_6534);
nor U7812 (N_7812,N_6348,N_6045);
or U7813 (N_7813,N_6651,N_6940);
xnor U7814 (N_7814,N_6643,N_6199);
and U7815 (N_7815,N_6374,N_6456);
or U7816 (N_7816,N_6638,N_6101);
xor U7817 (N_7817,N_6954,N_6477);
nand U7818 (N_7818,N_6913,N_6105);
or U7819 (N_7819,N_6341,N_6506);
nor U7820 (N_7820,N_6802,N_6000);
nand U7821 (N_7821,N_6388,N_6989);
nor U7822 (N_7822,N_6281,N_6165);
nor U7823 (N_7823,N_6342,N_6765);
and U7824 (N_7824,N_6347,N_6669);
and U7825 (N_7825,N_6790,N_6631);
xnor U7826 (N_7826,N_6495,N_6885);
nand U7827 (N_7827,N_6385,N_6093);
nand U7828 (N_7828,N_6888,N_6984);
or U7829 (N_7829,N_6165,N_6910);
xnor U7830 (N_7830,N_6998,N_6943);
nand U7831 (N_7831,N_6138,N_6169);
xor U7832 (N_7832,N_6170,N_6308);
or U7833 (N_7833,N_6067,N_6587);
and U7834 (N_7834,N_6255,N_6956);
nor U7835 (N_7835,N_6109,N_6765);
or U7836 (N_7836,N_6670,N_6810);
xor U7837 (N_7837,N_6785,N_6213);
or U7838 (N_7838,N_6300,N_6538);
nor U7839 (N_7839,N_6122,N_6891);
and U7840 (N_7840,N_6094,N_6606);
or U7841 (N_7841,N_6461,N_6627);
or U7842 (N_7842,N_6172,N_6194);
nand U7843 (N_7843,N_6291,N_6409);
or U7844 (N_7844,N_6289,N_6775);
and U7845 (N_7845,N_6537,N_6732);
and U7846 (N_7846,N_6240,N_6431);
or U7847 (N_7847,N_6542,N_6194);
nand U7848 (N_7848,N_6567,N_6579);
and U7849 (N_7849,N_6507,N_6553);
xnor U7850 (N_7850,N_6830,N_6198);
and U7851 (N_7851,N_6022,N_6020);
xor U7852 (N_7852,N_6978,N_6981);
and U7853 (N_7853,N_6646,N_6701);
nand U7854 (N_7854,N_6254,N_6342);
and U7855 (N_7855,N_6427,N_6310);
nand U7856 (N_7856,N_6662,N_6991);
nor U7857 (N_7857,N_6022,N_6302);
nand U7858 (N_7858,N_6624,N_6154);
and U7859 (N_7859,N_6995,N_6275);
nand U7860 (N_7860,N_6223,N_6703);
xnor U7861 (N_7861,N_6305,N_6480);
nor U7862 (N_7862,N_6788,N_6500);
xnor U7863 (N_7863,N_6552,N_6597);
xor U7864 (N_7864,N_6739,N_6207);
nand U7865 (N_7865,N_6061,N_6022);
and U7866 (N_7866,N_6537,N_6688);
nand U7867 (N_7867,N_6435,N_6447);
xnor U7868 (N_7868,N_6876,N_6534);
and U7869 (N_7869,N_6940,N_6720);
nor U7870 (N_7870,N_6243,N_6146);
xor U7871 (N_7871,N_6628,N_6978);
nand U7872 (N_7872,N_6196,N_6245);
or U7873 (N_7873,N_6672,N_6906);
nor U7874 (N_7874,N_6166,N_6000);
nor U7875 (N_7875,N_6887,N_6666);
nand U7876 (N_7876,N_6758,N_6902);
nand U7877 (N_7877,N_6130,N_6197);
and U7878 (N_7878,N_6595,N_6913);
and U7879 (N_7879,N_6396,N_6725);
or U7880 (N_7880,N_6891,N_6672);
or U7881 (N_7881,N_6665,N_6307);
nor U7882 (N_7882,N_6714,N_6075);
or U7883 (N_7883,N_6439,N_6940);
and U7884 (N_7884,N_6158,N_6446);
and U7885 (N_7885,N_6344,N_6011);
nand U7886 (N_7886,N_6159,N_6277);
and U7887 (N_7887,N_6599,N_6854);
and U7888 (N_7888,N_6436,N_6904);
nand U7889 (N_7889,N_6850,N_6308);
nand U7890 (N_7890,N_6231,N_6874);
nor U7891 (N_7891,N_6767,N_6754);
or U7892 (N_7892,N_6761,N_6059);
and U7893 (N_7893,N_6698,N_6722);
xnor U7894 (N_7894,N_6731,N_6715);
xor U7895 (N_7895,N_6075,N_6927);
and U7896 (N_7896,N_6706,N_6898);
or U7897 (N_7897,N_6155,N_6000);
xnor U7898 (N_7898,N_6559,N_6472);
or U7899 (N_7899,N_6873,N_6671);
and U7900 (N_7900,N_6116,N_6548);
and U7901 (N_7901,N_6271,N_6069);
or U7902 (N_7902,N_6472,N_6743);
and U7903 (N_7903,N_6941,N_6268);
xnor U7904 (N_7904,N_6142,N_6651);
xnor U7905 (N_7905,N_6964,N_6490);
nand U7906 (N_7906,N_6510,N_6817);
or U7907 (N_7907,N_6655,N_6227);
nor U7908 (N_7908,N_6072,N_6211);
or U7909 (N_7909,N_6613,N_6470);
and U7910 (N_7910,N_6948,N_6259);
nor U7911 (N_7911,N_6901,N_6683);
or U7912 (N_7912,N_6363,N_6526);
nor U7913 (N_7913,N_6440,N_6281);
nand U7914 (N_7914,N_6706,N_6088);
xnor U7915 (N_7915,N_6477,N_6804);
or U7916 (N_7916,N_6199,N_6363);
nand U7917 (N_7917,N_6598,N_6604);
nor U7918 (N_7918,N_6052,N_6738);
nand U7919 (N_7919,N_6651,N_6445);
and U7920 (N_7920,N_6345,N_6776);
nand U7921 (N_7921,N_6740,N_6933);
nand U7922 (N_7922,N_6786,N_6410);
xnor U7923 (N_7923,N_6843,N_6967);
nand U7924 (N_7924,N_6251,N_6739);
xor U7925 (N_7925,N_6001,N_6129);
nand U7926 (N_7926,N_6997,N_6885);
and U7927 (N_7927,N_6952,N_6002);
nand U7928 (N_7928,N_6438,N_6243);
or U7929 (N_7929,N_6283,N_6892);
nor U7930 (N_7930,N_6731,N_6215);
or U7931 (N_7931,N_6825,N_6370);
nand U7932 (N_7932,N_6585,N_6399);
xor U7933 (N_7933,N_6886,N_6847);
nor U7934 (N_7934,N_6436,N_6339);
nand U7935 (N_7935,N_6044,N_6411);
or U7936 (N_7936,N_6937,N_6132);
and U7937 (N_7937,N_6451,N_6335);
and U7938 (N_7938,N_6241,N_6698);
or U7939 (N_7939,N_6881,N_6763);
nor U7940 (N_7940,N_6316,N_6719);
or U7941 (N_7941,N_6269,N_6771);
and U7942 (N_7942,N_6833,N_6597);
and U7943 (N_7943,N_6455,N_6718);
nor U7944 (N_7944,N_6016,N_6097);
or U7945 (N_7945,N_6427,N_6583);
xor U7946 (N_7946,N_6609,N_6008);
or U7947 (N_7947,N_6321,N_6490);
and U7948 (N_7948,N_6660,N_6741);
and U7949 (N_7949,N_6741,N_6856);
or U7950 (N_7950,N_6770,N_6594);
or U7951 (N_7951,N_6887,N_6892);
nand U7952 (N_7952,N_6005,N_6362);
xnor U7953 (N_7953,N_6305,N_6780);
or U7954 (N_7954,N_6848,N_6422);
nor U7955 (N_7955,N_6061,N_6425);
nor U7956 (N_7956,N_6459,N_6892);
and U7957 (N_7957,N_6645,N_6031);
nor U7958 (N_7958,N_6119,N_6633);
and U7959 (N_7959,N_6763,N_6661);
and U7960 (N_7960,N_6039,N_6237);
nand U7961 (N_7961,N_6517,N_6681);
or U7962 (N_7962,N_6691,N_6826);
nor U7963 (N_7963,N_6581,N_6170);
and U7964 (N_7964,N_6029,N_6894);
nor U7965 (N_7965,N_6781,N_6927);
nor U7966 (N_7966,N_6755,N_6930);
and U7967 (N_7967,N_6269,N_6743);
and U7968 (N_7968,N_6069,N_6233);
and U7969 (N_7969,N_6616,N_6962);
or U7970 (N_7970,N_6921,N_6724);
nand U7971 (N_7971,N_6382,N_6070);
nor U7972 (N_7972,N_6601,N_6264);
nand U7973 (N_7973,N_6683,N_6368);
xor U7974 (N_7974,N_6632,N_6220);
or U7975 (N_7975,N_6305,N_6174);
nor U7976 (N_7976,N_6130,N_6437);
nor U7977 (N_7977,N_6263,N_6569);
xor U7978 (N_7978,N_6112,N_6737);
and U7979 (N_7979,N_6552,N_6555);
nand U7980 (N_7980,N_6602,N_6592);
xor U7981 (N_7981,N_6133,N_6956);
and U7982 (N_7982,N_6245,N_6155);
nand U7983 (N_7983,N_6957,N_6896);
xor U7984 (N_7984,N_6183,N_6088);
and U7985 (N_7985,N_6131,N_6406);
nor U7986 (N_7986,N_6083,N_6155);
and U7987 (N_7987,N_6591,N_6341);
and U7988 (N_7988,N_6770,N_6746);
xor U7989 (N_7989,N_6288,N_6487);
xor U7990 (N_7990,N_6500,N_6930);
xor U7991 (N_7991,N_6207,N_6292);
nor U7992 (N_7992,N_6981,N_6281);
and U7993 (N_7993,N_6321,N_6571);
xnor U7994 (N_7994,N_6740,N_6637);
nor U7995 (N_7995,N_6538,N_6812);
and U7996 (N_7996,N_6924,N_6366);
nor U7997 (N_7997,N_6481,N_6465);
nand U7998 (N_7998,N_6140,N_6552);
and U7999 (N_7999,N_6276,N_6755);
nor U8000 (N_8000,N_7213,N_7200);
xor U8001 (N_8001,N_7344,N_7948);
or U8002 (N_8002,N_7264,N_7936);
nor U8003 (N_8003,N_7730,N_7028);
or U8004 (N_8004,N_7336,N_7727);
and U8005 (N_8005,N_7412,N_7013);
xor U8006 (N_8006,N_7233,N_7031);
and U8007 (N_8007,N_7614,N_7268);
and U8008 (N_8008,N_7751,N_7868);
nand U8009 (N_8009,N_7760,N_7805);
and U8010 (N_8010,N_7899,N_7556);
or U8011 (N_8011,N_7754,N_7974);
or U8012 (N_8012,N_7650,N_7257);
nor U8013 (N_8013,N_7922,N_7806);
xnor U8014 (N_8014,N_7318,N_7005);
and U8015 (N_8015,N_7267,N_7039);
or U8016 (N_8016,N_7712,N_7226);
and U8017 (N_8017,N_7792,N_7341);
xnor U8018 (N_8018,N_7865,N_7400);
or U8019 (N_8019,N_7354,N_7174);
and U8020 (N_8020,N_7181,N_7687);
nor U8021 (N_8021,N_7006,N_7225);
or U8022 (N_8022,N_7721,N_7443);
and U8023 (N_8023,N_7686,N_7821);
xnor U8024 (N_8024,N_7581,N_7552);
nor U8025 (N_8025,N_7563,N_7555);
nor U8026 (N_8026,N_7889,N_7606);
xor U8027 (N_8027,N_7757,N_7572);
nand U8028 (N_8028,N_7017,N_7693);
nand U8029 (N_8029,N_7585,N_7111);
xnor U8030 (N_8030,N_7077,N_7998);
xnor U8031 (N_8031,N_7176,N_7208);
and U8032 (N_8032,N_7060,N_7363);
xnor U8033 (N_8033,N_7676,N_7682);
or U8034 (N_8034,N_7625,N_7883);
xor U8035 (N_8035,N_7022,N_7837);
xor U8036 (N_8036,N_7755,N_7628);
or U8037 (N_8037,N_7371,N_7718);
nand U8038 (N_8038,N_7924,N_7553);
or U8039 (N_8039,N_7912,N_7360);
nor U8040 (N_8040,N_7421,N_7397);
or U8041 (N_8041,N_7826,N_7423);
nand U8042 (N_8042,N_7689,N_7918);
nor U8043 (N_8043,N_7781,N_7876);
nand U8044 (N_8044,N_7498,N_7593);
and U8045 (N_8045,N_7231,N_7603);
nand U8046 (N_8046,N_7660,N_7128);
nand U8047 (N_8047,N_7582,N_7476);
or U8048 (N_8048,N_7189,N_7833);
nor U8049 (N_8049,N_7367,N_7444);
xor U8050 (N_8050,N_7294,N_7595);
and U8051 (N_8051,N_7938,N_7795);
or U8052 (N_8052,N_7641,N_7507);
and U8053 (N_8053,N_7254,N_7223);
xor U8054 (N_8054,N_7265,N_7583);
xnor U8055 (N_8055,N_7588,N_7932);
nor U8056 (N_8056,N_7089,N_7199);
nand U8057 (N_8057,N_7368,N_7631);
nor U8058 (N_8058,N_7056,N_7277);
nor U8059 (N_8059,N_7157,N_7505);
xnor U8060 (N_8060,N_7736,N_7870);
or U8061 (N_8061,N_7527,N_7976);
or U8062 (N_8062,N_7418,N_7433);
xor U8063 (N_8063,N_7680,N_7475);
nand U8064 (N_8064,N_7081,N_7486);
xor U8065 (N_8065,N_7009,N_7000);
nor U8066 (N_8066,N_7049,N_7352);
nor U8067 (N_8067,N_7840,N_7280);
or U8068 (N_8068,N_7731,N_7129);
nand U8069 (N_8069,N_7801,N_7304);
nor U8070 (N_8070,N_7518,N_7732);
nor U8071 (N_8071,N_7988,N_7608);
and U8072 (N_8072,N_7076,N_7432);
and U8073 (N_8073,N_7916,N_7927);
and U8074 (N_8074,N_7725,N_7671);
or U8075 (N_8075,N_7282,N_7414);
and U8076 (N_8076,N_7420,N_7182);
and U8077 (N_8077,N_7714,N_7402);
nand U8078 (N_8078,N_7985,N_7422);
xnor U8079 (N_8079,N_7255,N_7955);
nand U8080 (N_8080,N_7707,N_7458);
and U8081 (N_8081,N_7487,N_7205);
nor U8082 (N_8082,N_7121,N_7695);
and U8083 (N_8083,N_7424,N_7470);
nor U8084 (N_8084,N_7219,N_7087);
xnor U8085 (N_8085,N_7417,N_7733);
xnor U8086 (N_8086,N_7366,N_7279);
and U8087 (N_8087,N_7055,N_7888);
nor U8088 (N_8088,N_7559,N_7679);
nand U8089 (N_8089,N_7549,N_7197);
nor U8090 (N_8090,N_7163,N_7093);
or U8091 (N_8091,N_7361,N_7147);
nand U8092 (N_8092,N_7990,N_7744);
nor U8093 (N_8093,N_7235,N_7848);
and U8094 (N_8094,N_7669,N_7289);
nand U8095 (N_8095,N_7873,N_7831);
or U8096 (N_8096,N_7465,N_7243);
nand U8097 (N_8097,N_7229,N_7961);
and U8098 (N_8098,N_7619,N_7075);
and U8099 (N_8099,N_7320,N_7867);
xnor U8100 (N_8100,N_7038,N_7774);
nor U8101 (N_8101,N_7393,N_7069);
nor U8102 (N_8102,N_7646,N_7701);
or U8103 (N_8103,N_7431,N_7372);
nor U8104 (N_8104,N_7584,N_7763);
nand U8105 (N_8105,N_7632,N_7083);
nor U8106 (N_8106,N_7617,N_7364);
nand U8107 (N_8107,N_7537,N_7053);
nor U8108 (N_8108,N_7849,N_7872);
nand U8109 (N_8109,N_7466,N_7058);
and U8110 (N_8110,N_7193,N_7705);
xnor U8111 (N_8111,N_7657,N_7313);
xor U8112 (N_8112,N_7376,N_7050);
and U8113 (N_8113,N_7312,N_7230);
xor U8114 (N_8114,N_7566,N_7975);
nand U8115 (N_8115,N_7984,N_7885);
nand U8116 (N_8116,N_7716,N_7856);
xor U8117 (N_8117,N_7790,N_7810);
xor U8118 (N_8118,N_7239,N_7569);
xor U8119 (N_8119,N_7604,N_7943);
nand U8120 (N_8120,N_7911,N_7258);
nand U8121 (N_8121,N_7812,N_7309);
nand U8122 (N_8122,N_7340,N_7272);
or U8123 (N_8123,N_7863,N_7112);
and U8124 (N_8124,N_7994,N_7579);
nor U8125 (N_8125,N_7652,N_7426);
xor U8126 (N_8126,N_7045,N_7962);
or U8127 (N_8127,N_7770,N_7122);
or U8128 (N_8128,N_7131,N_7110);
or U8129 (N_8129,N_7134,N_7074);
or U8130 (N_8130,N_7797,N_7630);
nand U8131 (N_8131,N_7036,N_7180);
or U8132 (N_8132,N_7471,N_7434);
or U8133 (N_8133,N_7085,N_7452);
or U8134 (N_8134,N_7843,N_7905);
or U8135 (N_8135,N_7859,N_7541);
xor U8136 (N_8136,N_7966,N_7827);
or U8137 (N_8137,N_7381,N_7117);
or U8138 (N_8138,N_7665,N_7184);
and U8139 (N_8139,N_7123,N_7140);
xor U8140 (N_8140,N_7807,N_7202);
or U8141 (N_8141,N_7884,N_7993);
or U8142 (N_8142,N_7203,N_7970);
nor U8143 (N_8143,N_7623,N_7079);
xnor U8144 (N_8144,N_7285,N_7830);
xor U8145 (N_8145,N_7250,N_7501);
xor U8146 (N_8146,N_7311,N_7410);
xor U8147 (N_8147,N_7002,N_7096);
nor U8148 (N_8148,N_7910,N_7535);
and U8149 (N_8149,N_7793,N_7351);
or U8150 (N_8150,N_7405,N_7611);
nor U8151 (N_8151,N_7963,N_7347);
and U8152 (N_8152,N_7438,N_7370);
xor U8153 (N_8153,N_7626,N_7035);
nor U8154 (N_8154,N_7777,N_7253);
xor U8155 (N_8155,N_7783,N_7146);
and U8156 (N_8156,N_7153,N_7078);
or U8157 (N_8157,N_7775,N_7717);
nand U8158 (N_8158,N_7214,N_7594);
xor U8159 (N_8159,N_7335,N_7880);
and U8160 (N_8160,N_7857,N_7847);
and U8161 (N_8161,N_7871,N_7310);
nand U8162 (N_8162,N_7427,N_7896);
nand U8163 (N_8163,N_7558,N_7448);
nor U8164 (N_8164,N_7598,N_7930);
nand U8165 (N_8165,N_7789,N_7404);
and U8166 (N_8166,N_7548,N_7064);
nand U8167 (N_8167,N_7511,N_7674);
nor U8168 (N_8168,N_7043,N_7490);
nor U8169 (N_8169,N_7365,N_7454);
nand U8170 (N_8170,N_7305,N_7528);
nor U8171 (N_8171,N_7495,N_7972);
and U8172 (N_8172,N_7479,N_7105);
xor U8173 (N_8173,N_7903,N_7408);
or U8174 (N_8174,N_7429,N_7869);
or U8175 (N_8175,N_7605,N_7252);
nand U8176 (N_8176,N_7383,N_7862);
or U8177 (N_8177,N_7769,N_7602);
or U8178 (N_8178,N_7021,N_7949);
xnor U8179 (N_8179,N_7879,N_7092);
nand U8180 (N_8180,N_7908,N_7349);
or U8181 (N_8181,N_7014,N_7296);
nand U8182 (N_8182,N_7771,N_7044);
or U8183 (N_8183,N_7287,N_7828);
xnor U8184 (N_8184,N_7920,N_7459);
xnor U8185 (N_8185,N_7251,N_7767);
nand U8186 (N_8186,N_7386,N_7001);
and U8187 (N_8187,N_7485,N_7571);
and U8188 (N_8188,N_7729,N_7544);
nand U8189 (N_8189,N_7708,N_7629);
nor U8190 (N_8190,N_7143,N_7195);
nand U8191 (N_8191,N_7356,N_7067);
nand U8192 (N_8192,N_7670,N_7357);
nand U8193 (N_8193,N_7151,N_7655);
or U8194 (N_8194,N_7982,N_7804);
xor U8195 (N_8195,N_7683,N_7168);
and U8196 (N_8196,N_7692,N_7166);
xor U8197 (N_8197,N_7915,N_7207);
nor U8198 (N_8198,N_7520,N_7832);
nand U8199 (N_8199,N_7720,N_7530);
nand U8200 (N_8200,N_7453,N_7973);
or U8201 (N_8201,N_7206,N_7185);
nor U8202 (N_8202,N_7428,N_7165);
xor U8203 (N_8203,N_7198,N_7467);
nor U8204 (N_8204,N_7483,N_7834);
or U8205 (N_8205,N_7981,N_7723);
or U8206 (N_8206,N_7461,N_7664);
nor U8207 (N_8207,N_7543,N_7644);
and U8208 (N_8208,N_7090,N_7124);
xnor U8209 (N_8209,N_7722,N_7314);
nand U8210 (N_8210,N_7517,N_7942);
nand U8211 (N_8211,N_7515,N_7413);
nand U8212 (N_8212,N_7618,N_7817);
nor U8213 (N_8213,N_7242,N_7024);
nand U8214 (N_8214,N_7224,N_7977);
nor U8215 (N_8215,N_7749,N_7882);
nor U8216 (N_8216,N_7983,N_7167);
nor U8217 (N_8217,N_7169,N_7564);
xnor U8218 (N_8218,N_7492,N_7577);
xnor U8219 (N_8219,N_7667,N_7474);
and U8220 (N_8220,N_7647,N_7950);
xnor U8221 (N_8221,N_7338,N_7878);
and U8222 (N_8222,N_7132,N_7048);
and U8223 (N_8223,N_7419,N_7100);
and U8224 (N_8224,N_7462,N_7108);
nand U8225 (N_8225,N_7854,N_7523);
xnor U8226 (N_8226,N_7190,N_7678);
nor U8227 (N_8227,N_7261,N_7234);
nand U8228 (N_8228,N_7324,N_7150);
xnor U8229 (N_8229,N_7904,N_7109);
xor U8230 (N_8230,N_7160,N_7097);
and U8231 (N_8231,N_7675,N_7525);
and U8232 (N_8232,N_7656,N_7509);
xor U8233 (N_8233,N_7946,N_7355);
xor U8234 (N_8234,N_7640,N_7791);
nor U8235 (N_8235,N_7968,N_7599);
nor U8236 (N_8236,N_7449,N_7302);
xnor U8237 (N_8237,N_7724,N_7874);
or U8238 (N_8238,N_7216,N_7457);
or U8239 (N_8239,N_7508,N_7416);
and U8240 (N_8240,N_7020,N_7245);
nor U8241 (N_8241,N_7481,N_7497);
nor U8242 (N_8242,N_7196,N_7964);
nand U8243 (N_8243,N_7928,N_7957);
xor U8244 (N_8244,N_7597,N_7934);
nand U8245 (N_8245,N_7561,N_7415);
and U8246 (N_8246,N_7526,N_7846);
or U8247 (N_8247,N_7348,N_7425);
xnor U8248 (N_8248,N_7937,N_7987);
or U8249 (N_8249,N_7947,N_7115);
or U8250 (N_8250,N_7685,N_7177);
and U8251 (N_8251,N_7596,N_7892);
xnor U8252 (N_8252,N_7071,N_7398);
xor U8253 (N_8253,N_7116,N_7662);
nand U8254 (N_8254,N_7468,N_7748);
nand U8255 (N_8255,N_7740,N_7694);
or U8256 (N_8256,N_7299,N_7306);
or U8257 (N_8257,N_7591,N_7909);
or U8258 (N_8258,N_7375,N_7220);
and U8259 (N_8259,N_7482,N_7780);
nor U8260 (N_8260,N_7504,N_7574);
xnor U8261 (N_8261,N_7025,N_7088);
nand U8262 (N_8262,N_7183,N_7902);
and U8263 (N_8263,N_7969,N_7350);
and U8264 (N_8264,N_7991,N_7127);
nand U8265 (N_8265,N_7330,N_7342);
nor U8266 (N_8266,N_7395,N_7051);
nor U8267 (N_8267,N_7886,N_7620);
nor U8268 (N_8268,N_7401,N_7329);
xnor U8269 (N_8269,N_7814,N_7709);
and U8270 (N_8270,N_7389,N_7297);
and U8271 (N_8271,N_7666,N_7753);
and U8272 (N_8272,N_7275,N_7362);
xnor U8273 (N_8273,N_7634,N_7900);
nor U8274 (N_8274,N_7283,N_7489);
nor U8275 (N_8275,N_7808,N_7041);
nor U8276 (N_8276,N_7951,N_7046);
nand U8277 (N_8277,N_7392,N_7472);
and U8278 (N_8278,N_7411,N_7845);
xnor U8279 (N_8279,N_7399,N_7906);
xnor U8280 (N_8280,N_7798,N_7500);
nand U8281 (N_8281,N_7741,N_7534);
and U8282 (N_8282,N_7945,N_7374);
and U8283 (N_8283,N_7057,N_7824);
xor U8284 (N_8284,N_7822,N_7894);
nand U8285 (N_8285,N_7012,N_7378);
nor U8286 (N_8286,N_7688,N_7575);
xor U8287 (N_8287,N_7278,N_7815);
nand U8288 (N_8288,N_7086,N_7825);
nand U8289 (N_8289,N_7496,N_7697);
or U8290 (N_8290,N_7866,N_7861);
xor U8291 (N_8291,N_7719,N_7855);
and U8292 (N_8292,N_7547,N_7691);
xnor U8293 (N_8293,N_7142,N_7803);
nand U8294 (N_8294,N_7735,N_7241);
and U8295 (N_8295,N_7782,N_7293);
nor U8296 (N_8296,N_7616,N_7385);
and U8297 (N_8297,N_7568,N_7015);
nor U8298 (N_8298,N_7322,N_7276);
nand U8299 (N_8299,N_7066,N_7651);
and U8300 (N_8300,N_7334,N_7711);
or U8301 (N_8301,N_7502,N_7271);
xnor U8302 (N_8302,N_7642,N_7004);
or U8303 (N_8303,N_7333,N_7034);
nor U8304 (N_8304,N_7439,N_7442);
xor U8305 (N_8305,N_7301,N_7171);
nand U8306 (N_8306,N_7484,N_7514);
xnor U8307 (N_8307,N_7155,N_7997);
nand U8308 (N_8308,N_7159,N_7139);
and U8309 (N_8309,N_7784,N_7463);
nor U8310 (N_8310,N_7152,N_7923);
nor U8311 (N_8311,N_7194,N_7103);
xnor U8312 (N_8312,N_7811,N_7690);
and U8313 (N_8313,N_7407,N_7018);
nand U8314 (N_8314,N_7645,N_7033);
and U8315 (N_8315,N_7510,N_7288);
nor U8316 (N_8316,N_7823,N_7145);
xnor U8317 (N_8317,N_7844,N_7546);
xnor U8318 (N_8318,N_7677,N_7084);
and U8319 (N_8319,N_7321,N_7533);
xor U8320 (N_8320,N_7772,N_7622);
xor U8321 (N_8321,N_7217,N_7073);
and U8322 (N_8322,N_7958,N_7126);
or U8323 (N_8323,N_7643,N_7170);
or U8324 (N_8324,N_7281,N_7842);
nor U8325 (N_8325,N_7391,N_7764);
nor U8326 (N_8326,N_7512,N_7455);
xor U8327 (N_8327,N_7102,N_7654);
nand U8328 (N_8328,N_7480,N_7238);
nand U8329 (N_8329,N_7125,N_7358);
nor U8330 (N_8330,N_7939,N_7699);
xor U8331 (N_8331,N_7901,N_7996);
nand U8332 (N_8332,N_7491,N_7668);
xor U8333 (N_8333,N_7788,N_7460);
xor U8334 (N_8334,N_7221,N_7637);
or U8335 (N_8335,N_7661,N_7373);
nand U8336 (N_8336,N_7186,N_7187);
or U8337 (N_8337,N_7858,N_7681);
nor U8338 (N_8338,N_7328,N_7726);
nand U8339 (N_8339,N_7099,N_7298);
xnor U8340 (N_8340,N_7030,N_7130);
nor U8341 (N_8341,N_7737,N_7891);
nor U8342 (N_8342,N_7308,N_7094);
and U8343 (N_8343,N_7802,N_7047);
and U8344 (N_8344,N_7388,N_7118);
and U8345 (N_8345,N_7343,N_7477);
nor U8346 (N_8346,N_7540,N_7698);
and U8347 (N_8347,N_7488,N_7759);
xnor U8348 (N_8348,N_7451,N_7913);
nand U8349 (N_8349,N_7291,N_7895);
nand U8350 (N_8350,N_7881,N_7337);
or U8351 (N_8351,N_7259,N_7851);
nor U8352 (N_8352,N_7766,N_7332);
nand U8353 (N_8353,N_7567,N_7829);
nand U8354 (N_8354,N_7149,N_7853);
xnor U8355 (N_8355,N_7580,N_7052);
xnor U8356 (N_8356,N_7440,N_7960);
xnor U8357 (N_8357,N_7746,N_7779);
nand U8358 (N_8358,N_7023,N_7464);
xor U8359 (N_8359,N_7369,N_7156);
or U8360 (N_8360,N_7138,N_7326);
nand U8361 (N_8361,N_7104,N_7787);
xor U8362 (N_8362,N_7765,N_7536);
nor U8363 (N_8363,N_7435,N_7327);
or U8364 (N_8364,N_7761,N_7172);
nand U8365 (N_8365,N_7739,N_7237);
nor U8366 (N_8366,N_7545,N_7260);
xnor U8367 (N_8367,N_7919,N_7713);
or U8368 (N_8368,N_7954,N_7917);
or U8369 (N_8369,N_7228,N_7612);
nand U8370 (N_8370,N_7494,N_7841);
nand U8371 (N_8371,N_7246,N_7852);
nor U8372 (N_8372,N_7550,N_7215);
nand U8373 (N_8373,N_7560,N_7072);
xor U8374 (N_8374,N_7813,N_7800);
or U8375 (N_8375,N_7624,N_7154);
nand U8376 (N_8376,N_7926,N_7995);
nand U8377 (N_8377,N_7148,N_7010);
or U8378 (N_8378,N_7008,N_7119);
xnor U8379 (N_8379,N_7380,N_7286);
xor U8380 (N_8380,N_7345,N_7532);
or U8381 (N_8381,N_7702,N_7839);
nor U8382 (N_8382,N_7026,N_7240);
nor U8383 (N_8383,N_7897,N_7639);
or U8384 (N_8384,N_7953,N_7430);
or U8385 (N_8385,N_7274,N_7587);
xnor U8386 (N_8386,N_7967,N_7437);
xnor U8387 (N_8387,N_7519,N_7893);
nor U8388 (N_8388,N_7396,N_7971);
nor U8389 (N_8389,N_7672,N_7752);
nand U8390 (N_8390,N_7270,N_7820);
nor U8391 (N_8391,N_7758,N_7211);
xnor U8392 (N_8392,N_7648,N_7210);
nor U8393 (N_8393,N_7027,N_7522);
or U8394 (N_8394,N_7263,N_7120);
xor U8395 (N_8395,N_7794,N_7204);
or U8396 (N_8396,N_7609,N_7877);
and U8397 (N_8397,N_7607,N_7658);
and U8398 (N_8398,N_7379,N_7011);
nor U8399 (N_8399,N_7315,N_7570);
and U8400 (N_8400,N_7082,N_7638);
or U8401 (N_8401,N_7353,N_7450);
nor U8402 (N_8402,N_7222,N_7921);
nand U8403 (N_8403,N_7135,N_7499);
and U8404 (N_8404,N_7173,N_7319);
and U8405 (N_8405,N_7161,N_7256);
and U8406 (N_8406,N_7158,N_7290);
and U8407 (N_8407,N_7710,N_7019);
xnor U8408 (N_8408,N_7809,N_7836);
and U8409 (N_8409,N_7133,N_7236);
and U8410 (N_8410,N_7557,N_7042);
nand U8411 (N_8411,N_7107,N_7621);
xnor U8412 (N_8412,N_7095,N_7387);
nand U8413 (N_8413,N_7786,N_7091);
xor U8414 (N_8414,N_7706,N_7040);
xor U8415 (N_8415,N_7303,N_7065);
and U8416 (N_8416,N_7521,N_7113);
xnor U8417 (N_8417,N_7359,N_7931);
nor U8418 (N_8418,N_7538,N_7377);
nor U8419 (N_8419,N_7218,N_7244);
nor U8420 (N_8420,N_7554,N_7295);
xor U8421 (N_8421,N_7406,N_7300);
and U8422 (N_8422,N_7663,N_7745);
xnor U8423 (N_8423,N_7586,N_7601);
nand U8424 (N_8424,N_7999,N_7673);
and U8425 (N_8425,N_7633,N_7696);
nor U8426 (N_8426,N_7636,N_7684);
xnor U8427 (N_8427,N_7860,N_7284);
and U8428 (N_8428,N_7940,N_7980);
or U8429 (N_8429,N_7441,N_7390);
xor U8430 (N_8430,N_7653,N_7610);
or U8431 (N_8431,N_7956,N_7576);
xor U8432 (N_8432,N_7925,N_7978);
and U8433 (N_8433,N_7573,N_7890);
and U8434 (N_8434,N_7192,N_7212);
and U8435 (N_8435,N_7191,N_7627);
nand U8436 (N_8436,N_7513,N_7747);
nand U8437 (N_8437,N_7469,N_7162);
and U8438 (N_8438,N_7835,N_7819);
or U8439 (N_8439,N_7589,N_7952);
and U8440 (N_8440,N_7478,N_7164);
or U8441 (N_8441,N_7944,N_7756);
xnor U8442 (N_8442,N_7898,N_7054);
and U8443 (N_8443,N_7635,N_7933);
nand U8444 (N_8444,N_7382,N_7273);
nor U8445 (N_8445,N_7503,N_7551);
xnor U8446 (N_8446,N_7773,N_7317);
and U8447 (N_8447,N_7307,N_7175);
nand U8448 (N_8448,N_7070,N_7838);
and U8449 (N_8449,N_7201,N_7114);
nor U8450 (N_8450,N_7292,N_7816);
nand U8451 (N_8451,N_7531,N_7456);
and U8452 (N_8452,N_7700,N_7059);
xor U8453 (N_8453,N_7445,N_7394);
nand U8454 (N_8454,N_7715,N_7742);
nor U8455 (N_8455,N_7037,N_7738);
or U8456 (N_8456,N_7704,N_7703);
nand U8457 (N_8457,N_7232,N_7935);
or U8458 (N_8458,N_7144,N_7136);
xor U8459 (N_8459,N_7785,N_7959);
xor U8460 (N_8460,N_7864,N_7269);
and U8461 (N_8461,N_7179,N_7098);
xnor U8462 (N_8462,N_7529,N_7516);
or U8463 (N_8463,N_7063,N_7178);
nand U8464 (N_8464,N_7248,N_7106);
or U8465 (N_8465,N_7965,N_7796);
nand U8466 (N_8466,N_7316,N_7101);
and U8467 (N_8467,N_7323,N_7649);
or U8468 (N_8468,N_7062,N_7776);
and U8469 (N_8469,N_7778,N_7346);
nor U8470 (N_8470,N_7542,N_7068);
nor U8471 (N_8471,N_7209,N_7590);
nor U8472 (N_8472,N_7565,N_7613);
nor U8473 (N_8473,N_7615,N_7907);
nor U8474 (N_8474,N_7734,N_7941);
and U8475 (N_8475,N_7029,N_7850);
xnor U8476 (N_8476,N_7247,N_7061);
and U8477 (N_8477,N_7929,N_7914);
nor U8478 (N_8478,N_7818,N_7768);
nand U8479 (N_8479,N_7562,N_7003);
nand U8480 (N_8480,N_7659,N_7080);
xor U8481 (N_8481,N_7524,N_7578);
or U8482 (N_8482,N_7506,N_7137);
xnor U8483 (N_8483,N_7331,N_7600);
nor U8484 (N_8484,N_7592,N_7799);
xnor U8485 (N_8485,N_7989,N_7141);
nor U8486 (N_8486,N_7325,N_7227);
or U8487 (N_8487,N_7266,N_7875);
nand U8488 (N_8488,N_7403,N_7016);
xor U8489 (N_8489,N_7979,N_7728);
and U8490 (N_8490,N_7188,N_7007);
and U8491 (N_8491,N_7986,N_7493);
and U8492 (N_8492,N_7887,N_7339);
or U8493 (N_8493,N_7447,N_7539);
xnor U8494 (N_8494,N_7446,N_7409);
xor U8495 (N_8495,N_7743,N_7436);
and U8496 (N_8496,N_7384,N_7473);
and U8497 (N_8497,N_7032,N_7750);
nand U8498 (N_8498,N_7262,N_7249);
or U8499 (N_8499,N_7992,N_7762);
nand U8500 (N_8500,N_7803,N_7895);
xor U8501 (N_8501,N_7556,N_7739);
or U8502 (N_8502,N_7443,N_7637);
and U8503 (N_8503,N_7256,N_7614);
nor U8504 (N_8504,N_7310,N_7603);
or U8505 (N_8505,N_7341,N_7920);
nand U8506 (N_8506,N_7188,N_7707);
xnor U8507 (N_8507,N_7050,N_7923);
nor U8508 (N_8508,N_7538,N_7490);
and U8509 (N_8509,N_7473,N_7542);
nand U8510 (N_8510,N_7742,N_7398);
or U8511 (N_8511,N_7224,N_7740);
nand U8512 (N_8512,N_7913,N_7761);
or U8513 (N_8513,N_7532,N_7509);
nand U8514 (N_8514,N_7092,N_7040);
and U8515 (N_8515,N_7757,N_7115);
nand U8516 (N_8516,N_7476,N_7050);
nand U8517 (N_8517,N_7661,N_7663);
nand U8518 (N_8518,N_7450,N_7143);
and U8519 (N_8519,N_7504,N_7111);
nand U8520 (N_8520,N_7544,N_7888);
nor U8521 (N_8521,N_7007,N_7178);
nand U8522 (N_8522,N_7021,N_7860);
nor U8523 (N_8523,N_7837,N_7637);
or U8524 (N_8524,N_7978,N_7247);
nor U8525 (N_8525,N_7120,N_7492);
nand U8526 (N_8526,N_7512,N_7846);
nor U8527 (N_8527,N_7843,N_7864);
xnor U8528 (N_8528,N_7145,N_7431);
xnor U8529 (N_8529,N_7218,N_7449);
nor U8530 (N_8530,N_7403,N_7837);
nand U8531 (N_8531,N_7134,N_7664);
nand U8532 (N_8532,N_7686,N_7600);
and U8533 (N_8533,N_7773,N_7808);
xnor U8534 (N_8534,N_7444,N_7044);
xnor U8535 (N_8535,N_7395,N_7042);
or U8536 (N_8536,N_7444,N_7815);
nand U8537 (N_8537,N_7467,N_7558);
nand U8538 (N_8538,N_7769,N_7723);
xnor U8539 (N_8539,N_7334,N_7263);
xnor U8540 (N_8540,N_7498,N_7517);
nor U8541 (N_8541,N_7635,N_7593);
nand U8542 (N_8542,N_7565,N_7978);
xnor U8543 (N_8543,N_7754,N_7051);
nand U8544 (N_8544,N_7811,N_7645);
or U8545 (N_8545,N_7981,N_7108);
nor U8546 (N_8546,N_7993,N_7950);
xor U8547 (N_8547,N_7377,N_7110);
and U8548 (N_8548,N_7336,N_7245);
nor U8549 (N_8549,N_7941,N_7646);
nand U8550 (N_8550,N_7158,N_7922);
nor U8551 (N_8551,N_7801,N_7731);
or U8552 (N_8552,N_7215,N_7819);
or U8553 (N_8553,N_7048,N_7343);
nand U8554 (N_8554,N_7713,N_7870);
or U8555 (N_8555,N_7393,N_7212);
and U8556 (N_8556,N_7306,N_7225);
nor U8557 (N_8557,N_7254,N_7255);
nand U8558 (N_8558,N_7755,N_7608);
and U8559 (N_8559,N_7705,N_7920);
nor U8560 (N_8560,N_7241,N_7401);
nand U8561 (N_8561,N_7106,N_7107);
xor U8562 (N_8562,N_7815,N_7588);
xor U8563 (N_8563,N_7995,N_7683);
nor U8564 (N_8564,N_7754,N_7100);
xor U8565 (N_8565,N_7099,N_7844);
and U8566 (N_8566,N_7175,N_7540);
and U8567 (N_8567,N_7203,N_7671);
and U8568 (N_8568,N_7193,N_7231);
and U8569 (N_8569,N_7469,N_7363);
or U8570 (N_8570,N_7706,N_7633);
and U8571 (N_8571,N_7100,N_7867);
xor U8572 (N_8572,N_7387,N_7744);
and U8573 (N_8573,N_7720,N_7983);
xor U8574 (N_8574,N_7590,N_7490);
xor U8575 (N_8575,N_7820,N_7589);
nor U8576 (N_8576,N_7726,N_7411);
nand U8577 (N_8577,N_7348,N_7593);
nor U8578 (N_8578,N_7206,N_7464);
nand U8579 (N_8579,N_7511,N_7636);
and U8580 (N_8580,N_7533,N_7358);
and U8581 (N_8581,N_7521,N_7967);
or U8582 (N_8582,N_7725,N_7564);
and U8583 (N_8583,N_7209,N_7415);
nand U8584 (N_8584,N_7841,N_7206);
or U8585 (N_8585,N_7808,N_7246);
or U8586 (N_8586,N_7552,N_7853);
or U8587 (N_8587,N_7109,N_7111);
nor U8588 (N_8588,N_7408,N_7073);
or U8589 (N_8589,N_7496,N_7787);
xnor U8590 (N_8590,N_7278,N_7717);
and U8591 (N_8591,N_7880,N_7331);
xor U8592 (N_8592,N_7871,N_7054);
nor U8593 (N_8593,N_7031,N_7760);
xnor U8594 (N_8594,N_7733,N_7175);
nand U8595 (N_8595,N_7637,N_7318);
xor U8596 (N_8596,N_7163,N_7907);
nor U8597 (N_8597,N_7827,N_7703);
nand U8598 (N_8598,N_7400,N_7489);
nand U8599 (N_8599,N_7324,N_7752);
nor U8600 (N_8600,N_7318,N_7861);
xnor U8601 (N_8601,N_7634,N_7066);
xor U8602 (N_8602,N_7194,N_7994);
nor U8603 (N_8603,N_7285,N_7543);
nand U8604 (N_8604,N_7509,N_7843);
nor U8605 (N_8605,N_7220,N_7768);
nand U8606 (N_8606,N_7905,N_7105);
and U8607 (N_8607,N_7252,N_7171);
and U8608 (N_8608,N_7219,N_7438);
and U8609 (N_8609,N_7524,N_7446);
nor U8610 (N_8610,N_7320,N_7467);
nand U8611 (N_8611,N_7554,N_7005);
nor U8612 (N_8612,N_7489,N_7480);
nor U8613 (N_8613,N_7153,N_7265);
nand U8614 (N_8614,N_7347,N_7560);
or U8615 (N_8615,N_7718,N_7990);
and U8616 (N_8616,N_7576,N_7933);
xor U8617 (N_8617,N_7951,N_7643);
and U8618 (N_8618,N_7322,N_7526);
nand U8619 (N_8619,N_7332,N_7158);
nor U8620 (N_8620,N_7613,N_7287);
nand U8621 (N_8621,N_7860,N_7601);
and U8622 (N_8622,N_7764,N_7004);
nand U8623 (N_8623,N_7698,N_7876);
nand U8624 (N_8624,N_7634,N_7025);
xnor U8625 (N_8625,N_7362,N_7450);
xor U8626 (N_8626,N_7573,N_7007);
nand U8627 (N_8627,N_7488,N_7096);
and U8628 (N_8628,N_7991,N_7887);
or U8629 (N_8629,N_7353,N_7890);
nor U8630 (N_8630,N_7259,N_7241);
or U8631 (N_8631,N_7278,N_7272);
nand U8632 (N_8632,N_7647,N_7338);
xnor U8633 (N_8633,N_7445,N_7188);
nand U8634 (N_8634,N_7624,N_7243);
xor U8635 (N_8635,N_7085,N_7857);
nor U8636 (N_8636,N_7388,N_7002);
or U8637 (N_8637,N_7452,N_7927);
nor U8638 (N_8638,N_7315,N_7159);
or U8639 (N_8639,N_7342,N_7801);
nand U8640 (N_8640,N_7370,N_7491);
xor U8641 (N_8641,N_7344,N_7463);
nor U8642 (N_8642,N_7444,N_7500);
nor U8643 (N_8643,N_7037,N_7775);
and U8644 (N_8644,N_7568,N_7569);
nand U8645 (N_8645,N_7282,N_7538);
nand U8646 (N_8646,N_7592,N_7170);
xnor U8647 (N_8647,N_7437,N_7739);
or U8648 (N_8648,N_7671,N_7570);
xnor U8649 (N_8649,N_7517,N_7741);
nand U8650 (N_8650,N_7137,N_7544);
or U8651 (N_8651,N_7159,N_7000);
nand U8652 (N_8652,N_7364,N_7288);
nand U8653 (N_8653,N_7539,N_7140);
nor U8654 (N_8654,N_7153,N_7792);
or U8655 (N_8655,N_7603,N_7003);
or U8656 (N_8656,N_7487,N_7464);
nand U8657 (N_8657,N_7450,N_7825);
nor U8658 (N_8658,N_7501,N_7675);
nand U8659 (N_8659,N_7308,N_7472);
or U8660 (N_8660,N_7594,N_7017);
nand U8661 (N_8661,N_7723,N_7936);
and U8662 (N_8662,N_7336,N_7490);
xor U8663 (N_8663,N_7183,N_7649);
or U8664 (N_8664,N_7184,N_7250);
nor U8665 (N_8665,N_7722,N_7415);
or U8666 (N_8666,N_7864,N_7233);
xor U8667 (N_8667,N_7142,N_7251);
nand U8668 (N_8668,N_7303,N_7078);
nor U8669 (N_8669,N_7222,N_7805);
nand U8670 (N_8670,N_7620,N_7263);
and U8671 (N_8671,N_7110,N_7752);
or U8672 (N_8672,N_7241,N_7469);
and U8673 (N_8673,N_7253,N_7706);
or U8674 (N_8674,N_7273,N_7898);
nand U8675 (N_8675,N_7751,N_7917);
or U8676 (N_8676,N_7124,N_7899);
or U8677 (N_8677,N_7306,N_7544);
nand U8678 (N_8678,N_7156,N_7295);
nor U8679 (N_8679,N_7938,N_7136);
or U8680 (N_8680,N_7922,N_7174);
xor U8681 (N_8681,N_7807,N_7288);
or U8682 (N_8682,N_7870,N_7918);
nand U8683 (N_8683,N_7541,N_7942);
nor U8684 (N_8684,N_7842,N_7718);
nor U8685 (N_8685,N_7821,N_7999);
nor U8686 (N_8686,N_7258,N_7599);
xor U8687 (N_8687,N_7325,N_7130);
and U8688 (N_8688,N_7511,N_7815);
xnor U8689 (N_8689,N_7147,N_7942);
and U8690 (N_8690,N_7287,N_7166);
or U8691 (N_8691,N_7672,N_7324);
nand U8692 (N_8692,N_7614,N_7865);
nand U8693 (N_8693,N_7070,N_7395);
or U8694 (N_8694,N_7956,N_7716);
and U8695 (N_8695,N_7881,N_7463);
or U8696 (N_8696,N_7327,N_7423);
or U8697 (N_8697,N_7583,N_7848);
and U8698 (N_8698,N_7136,N_7281);
nor U8699 (N_8699,N_7635,N_7229);
nor U8700 (N_8700,N_7435,N_7574);
and U8701 (N_8701,N_7458,N_7569);
and U8702 (N_8702,N_7413,N_7977);
and U8703 (N_8703,N_7759,N_7476);
xnor U8704 (N_8704,N_7900,N_7620);
nor U8705 (N_8705,N_7868,N_7916);
nand U8706 (N_8706,N_7400,N_7737);
or U8707 (N_8707,N_7485,N_7332);
nand U8708 (N_8708,N_7323,N_7339);
xnor U8709 (N_8709,N_7176,N_7428);
or U8710 (N_8710,N_7192,N_7664);
and U8711 (N_8711,N_7547,N_7389);
and U8712 (N_8712,N_7120,N_7305);
or U8713 (N_8713,N_7495,N_7397);
nand U8714 (N_8714,N_7859,N_7354);
or U8715 (N_8715,N_7258,N_7546);
or U8716 (N_8716,N_7724,N_7332);
and U8717 (N_8717,N_7294,N_7254);
nand U8718 (N_8718,N_7402,N_7077);
xnor U8719 (N_8719,N_7931,N_7905);
xor U8720 (N_8720,N_7960,N_7095);
and U8721 (N_8721,N_7530,N_7633);
or U8722 (N_8722,N_7823,N_7084);
nand U8723 (N_8723,N_7839,N_7363);
nand U8724 (N_8724,N_7127,N_7272);
and U8725 (N_8725,N_7133,N_7561);
nor U8726 (N_8726,N_7794,N_7982);
and U8727 (N_8727,N_7707,N_7089);
and U8728 (N_8728,N_7121,N_7848);
nand U8729 (N_8729,N_7286,N_7428);
and U8730 (N_8730,N_7652,N_7401);
or U8731 (N_8731,N_7835,N_7648);
and U8732 (N_8732,N_7490,N_7376);
nand U8733 (N_8733,N_7361,N_7525);
and U8734 (N_8734,N_7720,N_7911);
and U8735 (N_8735,N_7107,N_7955);
nand U8736 (N_8736,N_7977,N_7982);
nand U8737 (N_8737,N_7471,N_7161);
nand U8738 (N_8738,N_7596,N_7714);
xnor U8739 (N_8739,N_7047,N_7897);
nor U8740 (N_8740,N_7553,N_7745);
nand U8741 (N_8741,N_7473,N_7821);
xor U8742 (N_8742,N_7756,N_7493);
nand U8743 (N_8743,N_7549,N_7032);
xor U8744 (N_8744,N_7936,N_7168);
xnor U8745 (N_8745,N_7018,N_7468);
nor U8746 (N_8746,N_7831,N_7083);
or U8747 (N_8747,N_7629,N_7294);
nand U8748 (N_8748,N_7925,N_7091);
or U8749 (N_8749,N_7751,N_7370);
xor U8750 (N_8750,N_7566,N_7983);
or U8751 (N_8751,N_7711,N_7168);
or U8752 (N_8752,N_7298,N_7017);
nor U8753 (N_8753,N_7979,N_7829);
xnor U8754 (N_8754,N_7392,N_7106);
or U8755 (N_8755,N_7175,N_7035);
and U8756 (N_8756,N_7468,N_7103);
nor U8757 (N_8757,N_7795,N_7321);
nor U8758 (N_8758,N_7658,N_7517);
nand U8759 (N_8759,N_7627,N_7920);
nand U8760 (N_8760,N_7155,N_7525);
and U8761 (N_8761,N_7147,N_7473);
xnor U8762 (N_8762,N_7840,N_7972);
nand U8763 (N_8763,N_7350,N_7886);
and U8764 (N_8764,N_7868,N_7671);
and U8765 (N_8765,N_7950,N_7031);
nand U8766 (N_8766,N_7463,N_7102);
nand U8767 (N_8767,N_7340,N_7251);
nand U8768 (N_8768,N_7697,N_7247);
nand U8769 (N_8769,N_7474,N_7804);
nor U8770 (N_8770,N_7885,N_7253);
or U8771 (N_8771,N_7007,N_7146);
or U8772 (N_8772,N_7589,N_7146);
xnor U8773 (N_8773,N_7360,N_7387);
nand U8774 (N_8774,N_7447,N_7167);
and U8775 (N_8775,N_7119,N_7325);
and U8776 (N_8776,N_7335,N_7219);
xnor U8777 (N_8777,N_7220,N_7822);
xor U8778 (N_8778,N_7753,N_7726);
nand U8779 (N_8779,N_7145,N_7670);
nor U8780 (N_8780,N_7223,N_7589);
nand U8781 (N_8781,N_7706,N_7030);
and U8782 (N_8782,N_7020,N_7634);
nor U8783 (N_8783,N_7027,N_7156);
or U8784 (N_8784,N_7805,N_7741);
and U8785 (N_8785,N_7904,N_7519);
or U8786 (N_8786,N_7097,N_7710);
nand U8787 (N_8787,N_7179,N_7692);
or U8788 (N_8788,N_7665,N_7430);
xor U8789 (N_8789,N_7251,N_7064);
or U8790 (N_8790,N_7118,N_7044);
or U8791 (N_8791,N_7511,N_7837);
or U8792 (N_8792,N_7371,N_7943);
and U8793 (N_8793,N_7988,N_7751);
or U8794 (N_8794,N_7718,N_7793);
nor U8795 (N_8795,N_7725,N_7437);
nor U8796 (N_8796,N_7821,N_7148);
nor U8797 (N_8797,N_7651,N_7388);
or U8798 (N_8798,N_7953,N_7807);
xor U8799 (N_8799,N_7951,N_7989);
and U8800 (N_8800,N_7806,N_7998);
xor U8801 (N_8801,N_7246,N_7926);
xor U8802 (N_8802,N_7328,N_7403);
xor U8803 (N_8803,N_7816,N_7681);
or U8804 (N_8804,N_7887,N_7040);
xor U8805 (N_8805,N_7082,N_7762);
xnor U8806 (N_8806,N_7956,N_7872);
and U8807 (N_8807,N_7453,N_7678);
and U8808 (N_8808,N_7086,N_7144);
nand U8809 (N_8809,N_7009,N_7966);
nor U8810 (N_8810,N_7733,N_7914);
or U8811 (N_8811,N_7918,N_7796);
and U8812 (N_8812,N_7527,N_7421);
or U8813 (N_8813,N_7221,N_7749);
or U8814 (N_8814,N_7766,N_7470);
nor U8815 (N_8815,N_7723,N_7386);
xnor U8816 (N_8816,N_7814,N_7963);
xor U8817 (N_8817,N_7959,N_7966);
nand U8818 (N_8818,N_7740,N_7373);
nor U8819 (N_8819,N_7860,N_7417);
nand U8820 (N_8820,N_7350,N_7932);
or U8821 (N_8821,N_7021,N_7448);
or U8822 (N_8822,N_7555,N_7763);
and U8823 (N_8823,N_7048,N_7476);
and U8824 (N_8824,N_7615,N_7869);
and U8825 (N_8825,N_7495,N_7062);
or U8826 (N_8826,N_7550,N_7273);
nand U8827 (N_8827,N_7480,N_7428);
xnor U8828 (N_8828,N_7637,N_7700);
or U8829 (N_8829,N_7020,N_7688);
nand U8830 (N_8830,N_7739,N_7138);
or U8831 (N_8831,N_7523,N_7502);
nand U8832 (N_8832,N_7059,N_7767);
nand U8833 (N_8833,N_7599,N_7821);
and U8834 (N_8834,N_7324,N_7925);
nand U8835 (N_8835,N_7732,N_7296);
nand U8836 (N_8836,N_7376,N_7850);
nand U8837 (N_8837,N_7453,N_7414);
xnor U8838 (N_8838,N_7885,N_7538);
and U8839 (N_8839,N_7931,N_7072);
xnor U8840 (N_8840,N_7696,N_7827);
xor U8841 (N_8841,N_7524,N_7912);
nand U8842 (N_8842,N_7570,N_7470);
nand U8843 (N_8843,N_7791,N_7397);
xor U8844 (N_8844,N_7976,N_7453);
and U8845 (N_8845,N_7690,N_7013);
nor U8846 (N_8846,N_7531,N_7445);
and U8847 (N_8847,N_7485,N_7711);
nor U8848 (N_8848,N_7588,N_7227);
xnor U8849 (N_8849,N_7263,N_7724);
nor U8850 (N_8850,N_7872,N_7163);
nand U8851 (N_8851,N_7495,N_7757);
nor U8852 (N_8852,N_7913,N_7845);
or U8853 (N_8853,N_7148,N_7189);
nand U8854 (N_8854,N_7763,N_7038);
nand U8855 (N_8855,N_7883,N_7881);
nand U8856 (N_8856,N_7830,N_7824);
and U8857 (N_8857,N_7058,N_7293);
nor U8858 (N_8858,N_7171,N_7286);
and U8859 (N_8859,N_7061,N_7444);
xor U8860 (N_8860,N_7409,N_7988);
nor U8861 (N_8861,N_7764,N_7343);
and U8862 (N_8862,N_7632,N_7974);
nand U8863 (N_8863,N_7910,N_7625);
xor U8864 (N_8864,N_7975,N_7538);
nand U8865 (N_8865,N_7456,N_7541);
xnor U8866 (N_8866,N_7342,N_7833);
xor U8867 (N_8867,N_7527,N_7747);
or U8868 (N_8868,N_7692,N_7156);
and U8869 (N_8869,N_7729,N_7796);
xor U8870 (N_8870,N_7101,N_7494);
nor U8871 (N_8871,N_7002,N_7714);
and U8872 (N_8872,N_7853,N_7112);
and U8873 (N_8873,N_7381,N_7639);
xnor U8874 (N_8874,N_7157,N_7635);
and U8875 (N_8875,N_7769,N_7076);
nor U8876 (N_8876,N_7905,N_7083);
nor U8877 (N_8877,N_7372,N_7352);
and U8878 (N_8878,N_7117,N_7071);
nand U8879 (N_8879,N_7173,N_7329);
nand U8880 (N_8880,N_7347,N_7863);
nand U8881 (N_8881,N_7811,N_7978);
and U8882 (N_8882,N_7471,N_7512);
xor U8883 (N_8883,N_7032,N_7637);
or U8884 (N_8884,N_7461,N_7066);
xor U8885 (N_8885,N_7884,N_7317);
or U8886 (N_8886,N_7067,N_7335);
nand U8887 (N_8887,N_7819,N_7525);
and U8888 (N_8888,N_7761,N_7073);
xnor U8889 (N_8889,N_7560,N_7813);
or U8890 (N_8890,N_7620,N_7471);
nand U8891 (N_8891,N_7598,N_7596);
and U8892 (N_8892,N_7482,N_7574);
nand U8893 (N_8893,N_7012,N_7329);
or U8894 (N_8894,N_7995,N_7780);
xor U8895 (N_8895,N_7793,N_7522);
xor U8896 (N_8896,N_7646,N_7399);
and U8897 (N_8897,N_7266,N_7163);
nor U8898 (N_8898,N_7864,N_7787);
xnor U8899 (N_8899,N_7733,N_7453);
nand U8900 (N_8900,N_7044,N_7562);
nor U8901 (N_8901,N_7473,N_7611);
nand U8902 (N_8902,N_7868,N_7276);
nand U8903 (N_8903,N_7854,N_7621);
nor U8904 (N_8904,N_7797,N_7233);
nor U8905 (N_8905,N_7410,N_7389);
nand U8906 (N_8906,N_7428,N_7833);
nand U8907 (N_8907,N_7028,N_7505);
and U8908 (N_8908,N_7656,N_7671);
and U8909 (N_8909,N_7216,N_7080);
nand U8910 (N_8910,N_7777,N_7632);
xor U8911 (N_8911,N_7983,N_7381);
xor U8912 (N_8912,N_7256,N_7078);
or U8913 (N_8913,N_7059,N_7364);
and U8914 (N_8914,N_7244,N_7658);
nor U8915 (N_8915,N_7365,N_7190);
or U8916 (N_8916,N_7913,N_7532);
xor U8917 (N_8917,N_7194,N_7526);
or U8918 (N_8918,N_7695,N_7160);
nand U8919 (N_8919,N_7053,N_7979);
xor U8920 (N_8920,N_7509,N_7029);
or U8921 (N_8921,N_7738,N_7027);
xor U8922 (N_8922,N_7716,N_7618);
or U8923 (N_8923,N_7036,N_7120);
xor U8924 (N_8924,N_7387,N_7533);
xnor U8925 (N_8925,N_7086,N_7740);
nor U8926 (N_8926,N_7743,N_7164);
or U8927 (N_8927,N_7823,N_7262);
nand U8928 (N_8928,N_7204,N_7258);
nand U8929 (N_8929,N_7030,N_7995);
or U8930 (N_8930,N_7890,N_7012);
xor U8931 (N_8931,N_7214,N_7332);
and U8932 (N_8932,N_7152,N_7894);
xnor U8933 (N_8933,N_7435,N_7422);
or U8934 (N_8934,N_7380,N_7738);
or U8935 (N_8935,N_7461,N_7965);
nand U8936 (N_8936,N_7170,N_7255);
nand U8937 (N_8937,N_7065,N_7335);
and U8938 (N_8938,N_7691,N_7983);
nand U8939 (N_8939,N_7826,N_7188);
and U8940 (N_8940,N_7517,N_7416);
or U8941 (N_8941,N_7792,N_7376);
and U8942 (N_8942,N_7238,N_7118);
nand U8943 (N_8943,N_7689,N_7433);
and U8944 (N_8944,N_7563,N_7261);
or U8945 (N_8945,N_7664,N_7738);
nand U8946 (N_8946,N_7007,N_7304);
xnor U8947 (N_8947,N_7875,N_7900);
xnor U8948 (N_8948,N_7351,N_7804);
nor U8949 (N_8949,N_7216,N_7517);
xor U8950 (N_8950,N_7246,N_7233);
xor U8951 (N_8951,N_7028,N_7413);
nand U8952 (N_8952,N_7270,N_7812);
nor U8953 (N_8953,N_7678,N_7015);
xnor U8954 (N_8954,N_7460,N_7873);
or U8955 (N_8955,N_7721,N_7356);
nand U8956 (N_8956,N_7676,N_7865);
or U8957 (N_8957,N_7971,N_7704);
and U8958 (N_8958,N_7293,N_7855);
nor U8959 (N_8959,N_7160,N_7961);
nor U8960 (N_8960,N_7159,N_7927);
or U8961 (N_8961,N_7635,N_7543);
and U8962 (N_8962,N_7132,N_7837);
and U8963 (N_8963,N_7173,N_7559);
nand U8964 (N_8964,N_7056,N_7216);
or U8965 (N_8965,N_7006,N_7638);
nand U8966 (N_8966,N_7089,N_7512);
nor U8967 (N_8967,N_7193,N_7229);
or U8968 (N_8968,N_7475,N_7076);
xor U8969 (N_8969,N_7407,N_7391);
xnor U8970 (N_8970,N_7685,N_7459);
nor U8971 (N_8971,N_7649,N_7252);
xor U8972 (N_8972,N_7717,N_7263);
xnor U8973 (N_8973,N_7446,N_7103);
nand U8974 (N_8974,N_7152,N_7355);
xnor U8975 (N_8975,N_7786,N_7643);
or U8976 (N_8976,N_7779,N_7183);
xnor U8977 (N_8977,N_7648,N_7274);
and U8978 (N_8978,N_7450,N_7503);
and U8979 (N_8979,N_7525,N_7121);
and U8980 (N_8980,N_7439,N_7199);
or U8981 (N_8981,N_7449,N_7981);
nand U8982 (N_8982,N_7795,N_7156);
xnor U8983 (N_8983,N_7363,N_7207);
nand U8984 (N_8984,N_7181,N_7453);
nand U8985 (N_8985,N_7884,N_7995);
and U8986 (N_8986,N_7542,N_7816);
nand U8987 (N_8987,N_7993,N_7535);
and U8988 (N_8988,N_7607,N_7958);
xor U8989 (N_8989,N_7248,N_7861);
or U8990 (N_8990,N_7613,N_7347);
and U8991 (N_8991,N_7641,N_7175);
xor U8992 (N_8992,N_7867,N_7282);
xor U8993 (N_8993,N_7641,N_7818);
and U8994 (N_8994,N_7718,N_7886);
xnor U8995 (N_8995,N_7609,N_7401);
and U8996 (N_8996,N_7936,N_7696);
nand U8997 (N_8997,N_7150,N_7947);
or U8998 (N_8998,N_7322,N_7960);
nor U8999 (N_8999,N_7361,N_7997);
xor U9000 (N_9000,N_8129,N_8342);
and U9001 (N_9001,N_8800,N_8251);
xor U9002 (N_9002,N_8906,N_8227);
nor U9003 (N_9003,N_8156,N_8645);
nor U9004 (N_9004,N_8330,N_8795);
nand U9005 (N_9005,N_8865,N_8676);
nand U9006 (N_9006,N_8025,N_8709);
or U9007 (N_9007,N_8395,N_8169);
nor U9008 (N_9008,N_8353,N_8858);
or U9009 (N_9009,N_8873,N_8933);
nor U9010 (N_9010,N_8638,N_8988);
nand U9011 (N_9011,N_8293,N_8606);
and U9012 (N_9012,N_8076,N_8135);
and U9013 (N_9013,N_8429,N_8028);
nor U9014 (N_9014,N_8287,N_8325);
xnor U9015 (N_9015,N_8947,N_8979);
nor U9016 (N_9016,N_8364,N_8171);
or U9017 (N_9017,N_8633,N_8414);
and U9018 (N_9018,N_8813,N_8178);
xor U9019 (N_9019,N_8419,N_8211);
xnor U9020 (N_9020,N_8210,N_8204);
nor U9021 (N_9021,N_8372,N_8486);
nand U9022 (N_9022,N_8432,N_8721);
nor U9023 (N_9023,N_8876,N_8538);
and U9024 (N_9024,N_8540,N_8860);
nor U9025 (N_9025,N_8086,N_8762);
or U9026 (N_9026,N_8331,N_8966);
nand U9027 (N_9027,N_8376,N_8650);
xnor U9028 (N_9028,N_8807,N_8201);
xnor U9029 (N_9029,N_8090,N_8791);
xor U9030 (N_9030,N_8617,N_8984);
nor U9031 (N_9031,N_8277,N_8627);
or U9032 (N_9032,N_8195,N_8886);
xnor U9033 (N_9033,N_8921,N_8336);
nor U9034 (N_9034,N_8073,N_8403);
and U9035 (N_9035,N_8112,N_8066);
nor U9036 (N_9036,N_8216,N_8501);
xor U9037 (N_9037,N_8790,N_8867);
nand U9038 (N_9038,N_8233,N_8767);
nor U9039 (N_9039,N_8522,N_8665);
and U9040 (N_9040,N_8231,N_8475);
xor U9041 (N_9041,N_8639,N_8685);
and U9042 (N_9042,N_8044,N_8549);
or U9043 (N_9043,N_8880,N_8085);
nand U9044 (N_9044,N_8386,N_8026);
nand U9045 (N_9045,N_8447,N_8595);
nand U9046 (N_9046,N_8013,N_8409);
nor U9047 (N_9047,N_8387,N_8763);
xor U9048 (N_9048,N_8582,N_8610);
nor U9049 (N_9049,N_8358,N_8920);
nor U9050 (N_9050,N_8508,N_8956);
nor U9051 (N_9051,N_8958,N_8547);
nor U9052 (N_9052,N_8713,N_8055);
or U9053 (N_9053,N_8731,N_8864);
nor U9054 (N_9054,N_8320,N_8900);
or U9055 (N_9055,N_8029,N_8101);
nor U9056 (N_9056,N_8955,N_8453);
and U9057 (N_9057,N_8374,N_8838);
and U9058 (N_9058,N_8276,N_8872);
and U9059 (N_9059,N_8989,N_8881);
nand U9060 (N_9060,N_8302,N_8602);
nand U9061 (N_9061,N_8964,N_8689);
and U9062 (N_9062,N_8912,N_8438);
and U9063 (N_9063,N_8518,N_8953);
xor U9064 (N_9064,N_8192,N_8868);
nor U9065 (N_9065,N_8114,N_8467);
or U9066 (N_9066,N_8603,N_8637);
and U9067 (N_9067,N_8674,N_8075);
and U9068 (N_9068,N_8539,N_8994);
nand U9069 (N_9069,N_8690,N_8841);
nor U9070 (N_9070,N_8328,N_8670);
nand U9071 (N_9071,N_8244,N_8707);
and U9072 (N_9072,N_8629,N_8533);
nand U9073 (N_9073,N_8837,N_8012);
and U9074 (N_9074,N_8095,N_8162);
and U9075 (N_9075,N_8586,N_8235);
or U9076 (N_9076,N_8407,N_8983);
nor U9077 (N_9077,N_8365,N_8067);
or U9078 (N_9078,N_8283,N_8879);
nor U9079 (N_9079,N_8628,N_8529);
or U9080 (N_9080,N_8772,N_8400);
nand U9081 (N_9081,N_8161,N_8976);
xnor U9082 (N_9082,N_8749,N_8843);
and U9083 (N_9083,N_8613,N_8271);
nor U9084 (N_9084,N_8489,N_8108);
nand U9085 (N_9085,N_8787,N_8669);
nor U9086 (N_9086,N_8016,N_8371);
or U9087 (N_9087,N_8959,N_8064);
nand U9088 (N_9088,N_8279,N_8788);
and U9089 (N_9089,N_8350,N_8315);
or U9090 (N_9090,N_8659,N_8744);
or U9091 (N_9091,N_8185,N_8347);
xnor U9092 (N_9092,N_8521,N_8011);
xnor U9093 (N_9093,N_8461,N_8575);
xnor U9094 (N_9094,N_8046,N_8745);
nand U9095 (N_9095,N_8198,N_8808);
and U9096 (N_9096,N_8498,N_8573);
and U9097 (N_9097,N_8250,N_8113);
and U9098 (N_9098,N_8775,N_8840);
nor U9099 (N_9099,N_8370,N_8809);
or U9100 (N_9100,N_8783,N_8708);
and U9101 (N_9101,N_8243,N_8612);
nor U9102 (N_9102,N_8491,N_8854);
nor U9103 (N_9103,N_8381,N_8001);
nand U9104 (N_9104,N_8159,N_8764);
and U9105 (N_9105,N_8693,N_8033);
or U9106 (N_9106,N_8971,N_8799);
nor U9107 (N_9107,N_8601,N_8862);
nor U9108 (N_9108,N_8150,N_8155);
xnor U9109 (N_9109,N_8779,N_8590);
xnor U9110 (N_9110,N_8926,N_8703);
nand U9111 (N_9111,N_8784,N_8759);
xnor U9112 (N_9112,N_8362,N_8607);
nor U9113 (N_9113,N_8644,N_8986);
nor U9114 (N_9114,N_8380,N_8004);
nor U9115 (N_9115,N_8847,N_8558);
xnor U9116 (N_9116,N_8750,N_8660);
xnor U9117 (N_9117,N_8014,N_8769);
nor U9118 (N_9118,N_8136,N_8985);
nor U9119 (N_9119,N_8304,N_8999);
and U9120 (N_9120,N_8062,N_8094);
nand U9121 (N_9121,N_8544,N_8511);
nand U9122 (N_9122,N_8507,N_8925);
or U9123 (N_9123,N_8175,N_8939);
and U9124 (N_9124,N_8431,N_8294);
nand U9125 (N_9125,N_8584,N_8478);
and U9126 (N_9126,N_8017,N_8272);
and U9127 (N_9127,N_8904,N_8401);
xor U9128 (N_9128,N_8126,N_8899);
and U9129 (N_9129,N_8487,N_8883);
or U9130 (N_9130,N_8123,N_8099);
xor U9131 (N_9131,N_8527,N_8484);
and U9132 (N_9132,N_8074,N_8399);
nand U9133 (N_9133,N_8146,N_8232);
xor U9134 (N_9134,N_8154,N_8087);
nor U9135 (N_9135,N_8036,N_8766);
xor U9136 (N_9136,N_8457,N_8394);
nand U9137 (N_9137,N_8059,N_8007);
nor U9138 (N_9138,N_8619,N_8804);
nor U9139 (N_9139,N_8483,N_8176);
nor U9140 (N_9140,N_8677,N_8416);
nor U9141 (N_9141,N_8887,N_8560);
nand U9142 (N_9142,N_8557,N_8445);
and U9143 (N_9143,N_8249,N_8226);
nand U9144 (N_9144,N_8631,N_8571);
and U9145 (N_9145,N_8542,N_8830);
xor U9146 (N_9146,N_8133,N_8088);
nand U9147 (N_9147,N_8642,N_8888);
nand U9148 (N_9148,N_8857,N_8781);
nor U9149 (N_9149,N_8335,N_8568);
xnor U9150 (N_9150,N_8065,N_8839);
nor U9151 (N_9151,N_8000,N_8165);
or U9152 (N_9152,N_8842,N_8463);
or U9153 (N_9153,N_8494,N_8168);
or U9154 (N_9154,N_8962,N_8577);
nand U9155 (N_9155,N_8318,N_8658);
nand U9156 (N_9156,N_8875,N_8563);
and U9157 (N_9157,N_8802,N_8069);
nor U9158 (N_9158,N_8877,N_8497);
nor U9159 (N_9159,N_8084,N_8182);
nor U9160 (N_9160,N_8488,N_8885);
nor U9161 (N_9161,N_8715,N_8117);
nand U9162 (N_9162,N_8071,N_8092);
or U9163 (N_9163,N_8667,N_8292);
and U9164 (N_9164,N_8082,N_8928);
and U9165 (N_9165,N_8417,N_8149);
nor U9166 (N_9166,N_8034,N_8106);
and U9167 (N_9167,N_8931,N_8058);
nand U9168 (N_9168,N_8600,N_8754);
nor U9169 (N_9169,N_8093,N_8716);
and U9170 (N_9170,N_8091,N_8728);
and U9171 (N_9171,N_8041,N_8428);
or U9172 (N_9172,N_8053,N_8555);
nor U9173 (N_9173,N_8897,N_8411);
nor U9174 (N_9174,N_8493,N_8479);
and U9175 (N_9175,N_8961,N_8869);
and U9176 (N_9176,N_8581,N_8214);
and U9177 (N_9177,N_8756,N_8684);
nand U9178 (N_9178,N_8177,N_8228);
and U9179 (N_9179,N_8596,N_8485);
and U9180 (N_9180,N_8385,N_8189);
or U9181 (N_9181,N_8780,N_8776);
nor U9182 (N_9182,N_8285,N_8910);
or U9183 (N_9183,N_8995,N_8193);
and U9184 (N_9184,N_8977,N_8474);
nand U9185 (N_9185,N_8472,N_8327);
or U9186 (N_9186,N_8505,N_8768);
nor U9187 (N_9187,N_8770,N_8104);
nand U9188 (N_9188,N_8143,N_8822);
or U9189 (N_9189,N_8337,N_8043);
nor U9190 (N_9190,N_8663,N_8755);
and U9191 (N_9191,N_8927,N_8805);
nand U9192 (N_9192,N_8183,N_8050);
xor U9193 (N_9193,N_8882,N_8245);
nor U9194 (N_9194,N_8230,N_8393);
or U9195 (N_9195,N_8918,N_8500);
and U9196 (N_9196,N_8859,N_8435);
xor U9197 (N_9197,N_8240,N_8343);
nor U9198 (N_9198,N_8944,N_8620);
or U9199 (N_9199,N_8433,N_8426);
nand U9200 (N_9200,N_8891,N_8777);
xor U9201 (N_9201,N_8943,N_8290);
nor U9202 (N_9202,N_8427,N_8615);
nor U9203 (N_9203,N_8579,N_8412);
nand U9204 (N_9204,N_8138,N_8229);
or U9205 (N_9205,N_8758,N_8535);
nand U9206 (N_9206,N_8105,N_8309);
xnor U9207 (N_9207,N_8710,N_8031);
or U9208 (N_9208,N_8032,N_8911);
and U9209 (N_9209,N_8641,N_8923);
xnor U9210 (N_9210,N_8566,N_8446);
and U9211 (N_9211,N_8625,N_8616);
xor U9212 (N_9212,N_8991,N_8391);
xor U9213 (N_9213,N_8730,N_8102);
nand U9214 (N_9214,N_8884,N_8960);
xnor U9215 (N_9215,N_8389,N_8167);
nand U9216 (N_9216,N_8711,N_8048);
or U9217 (N_9217,N_8696,N_8384);
and U9218 (N_9218,N_8828,N_8992);
xor U9219 (N_9219,N_8653,N_8422);
nor U9220 (N_9220,N_8778,N_8406);
or U9221 (N_9221,N_8760,N_8274);
nor U9222 (N_9222,N_8469,N_8465);
xor U9223 (N_9223,N_8786,N_8743);
xor U9224 (N_9224,N_8718,N_8848);
xnor U9225 (N_9225,N_8827,N_8098);
and U9226 (N_9226,N_8765,N_8806);
xnor U9227 (N_9227,N_8720,N_8691);
nor U9228 (N_9228,N_8423,N_8367);
nand U9229 (N_9229,N_8821,N_8975);
or U9230 (N_9230,N_8128,N_8726);
and U9231 (N_9231,N_8270,N_8333);
or U9232 (N_9232,N_8151,N_8222);
nor U9233 (N_9233,N_8009,N_8019);
nor U9234 (N_9234,N_8661,N_8903);
nor U9235 (N_9235,N_8456,N_8045);
nand U9236 (N_9236,N_8115,N_8424);
nor U9237 (N_9237,N_8952,N_8556);
nor U9238 (N_9238,N_8578,N_8338);
nand U9239 (N_9239,N_8717,N_8972);
nand U9240 (N_9240,N_8042,N_8852);
nand U9241 (N_9241,N_8378,N_8158);
nand U9242 (N_9242,N_8512,N_8224);
nand U9243 (N_9243,N_8207,N_8930);
xnor U9244 (N_9244,N_8725,N_8588);
nand U9245 (N_9245,N_8190,N_8565);
nand U9246 (N_9246,N_8825,N_8634);
xor U9247 (N_9247,N_8425,N_8773);
nand U9248 (N_9248,N_8916,N_8499);
and U9249 (N_9249,N_8241,N_8893);
or U9250 (N_9250,N_8597,N_8818);
xnor U9251 (N_9251,N_8941,N_8974);
or U9252 (N_9252,N_8314,N_8870);
nand U9253 (N_9253,N_8934,N_8164);
nand U9254 (N_9254,N_8570,N_8405);
nand U9255 (N_9255,N_8967,N_8968);
nand U9256 (N_9256,N_8184,N_8180);
or U9257 (N_9257,N_8205,N_8649);
nor U9258 (N_9258,N_8079,N_8397);
nor U9259 (N_9259,N_8534,N_8832);
or U9260 (N_9260,N_8462,N_8281);
xor U9261 (N_9261,N_8702,N_8587);
xnor U9262 (N_9262,N_8477,N_8450);
or U9263 (N_9263,N_8077,N_8626);
nand U9264 (N_9264,N_8894,N_8257);
xnor U9265 (N_9265,N_8267,N_8408);
xnor U9266 (N_9266,N_8664,N_8945);
or U9267 (N_9267,N_8246,N_8030);
nor U9268 (N_9268,N_8377,N_8915);
nor U9269 (N_9269,N_8608,N_8219);
nor U9270 (N_9270,N_8289,N_8970);
and U9271 (N_9271,N_8221,N_8360);
and U9272 (N_9272,N_8973,N_8348);
and U9273 (N_9273,N_8448,N_8040);
or U9274 (N_9274,N_8686,N_8439);
xor U9275 (N_9275,N_8797,N_8291);
and U9276 (N_9276,N_8890,N_8951);
nand U9277 (N_9277,N_8153,N_8080);
and U9278 (N_9278,N_8459,N_8509);
nand U9279 (N_9279,N_8266,N_8675);
nor U9280 (N_9280,N_8829,N_8134);
or U9281 (N_9281,N_8752,N_8413);
or U9282 (N_9282,N_8127,N_8441);
nand U9283 (N_9283,N_8727,N_8142);
nand U9284 (N_9284,N_8567,N_8390);
xnor U9285 (N_9285,N_8819,N_8208);
nor U9286 (N_9286,N_8037,N_8679);
and U9287 (N_9287,N_8311,N_8170);
and U9288 (N_9288,N_8206,N_8152);
or U9289 (N_9289,N_8735,N_8648);
and U9290 (N_9290,N_8023,N_8349);
nor U9291 (N_9291,N_8254,N_8212);
nor U9292 (N_9292,N_8357,N_8576);
nor U9293 (N_9293,N_8516,N_8609);
xnor U9294 (N_9294,N_8652,N_8256);
and U9295 (N_9295,N_8611,N_8495);
xnor U9296 (N_9296,N_8217,N_8237);
nand U9297 (N_9297,N_8305,N_8678);
nand U9298 (N_9298,N_8049,N_8593);
nor U9299 (N_9299,N_8396,N_8470);
and U9300 (N_9300,N_8751,N_8449);
or U9301 (N_9301,N_8308,N_8197);
nand U9302 (N_9302,N_8202,N_8295);
and U9303 (N_9303,N_8130,N_8363);
nand U9304 (N_9304,N_8255,N_8740);
xnor U9305 (N_9305,N_8836,N_8898);
or U9306 (N_9306,N_8585,N_8794);
xor U9307 (N_9307,N_8681,N_8286);
xor U9308 (N_9308,N_8078,N_8954);
nand U9309 (N_9309,N_8402,N_8174);
and U9310 (N_9310,N_8741,N_8356);
nand U9311 (N_9311,N_8793,N_8589);
and U9312 (N_9312,N_8545,N_8896);
xnor U9313 (N_9313,N_8996,N_8673);
nor U9314 (N_9314,N_8940,N_8273);
nor U9315 (N_9315,N_8199,N_8932);
xnor U9316 (N_9316,N_8196,N_8215);
nor U9317 (N_9317,N_8866,N_8810);
and U9318 (N_9318,N_8096,N_8275);
nand U9319 (N_9319,N_8662,N_8655);
or U9320 (N_9320,N_8490,N_8604);
or U9321 (N_9321,N_8103,N_8181);
or U9322 (N_9322,N_8020,N_8451);
or U9323 (N_9323,N_8420,N_8742);
nand U9324 (N_9324,N_8345,N_8100);
nand U9325 (N_9325,N_8166,N_8632);
nor U9326 (N_9326,N_8253,N_8666);
nand U9327 (N_9327,N_8147,N_8591);
or U9328 (N_9328,N_8824,N_8907);
and U9329 (N_9329,N_8543,N_8341);
nand U9330 (N_9330,N_8324,N_8938);
nand U9331 (N_9331,N_8110,N_8194);
or U9332 (N_9332,N_8909,N_8440);
or U9333 (N_9333,N_8120,N_8307);
or U9334 (N_9334,N_8460,N_8935);
or U9335 (N_9335,N_8415,N_8496);
nand U9336 (N_9336,N_8209,N_8316);
or U9337 (N_9337,N_8801,N_8580);
and U9338 (N_9338,N_8057,N_8892);
xor U9339 (N_9339,N_8109,N_8379);
nor U9340 (N_9340,N_8695,N_8383);
nor U9341 (N_9341,N_8024,N_8520);
or U9342 (N_9342,N_8905,N_8352);
xnor U9343 (N_9343,N_8035,N_8895);
and U9344 (N_9344,N_8122,N_8340);
and U9345 (N_9345,N_8874,N_8265);
nand U9346 (N_9346,N_8346,N_8969);
and U9347 (N_9347,N_8814,N_8853);
xor U9348 (N_9348,N_8990,N_8692);
and U9349 (N_9349,N_8361,N_8220);
nor U9350 (N_9350,N_8811,N_8223);
nor U9351 (N_9351,N_8630,N_8284);
xnor U9352 (N_9352,N_8998,N_8553);
nor U9353 (N_9353,N_8248,N_8430);
nor U9354 (N_9354,N_8278,N_8089);
or U9355 (N_9355,N_8319,N_8442);
nand U9356 (N_9356,N_8753,N_8418);
nand U9357 (N_9357,N_8525,N_8502);
or U9358 (N_9358,N_8021,N_8982);
and U9359 (N_9359,N_8981,N_8052);
or U9360 (N_9360,N_8599,N_8317);
nand U9361 (N_9361,N_8313,N_8282);
xnor U9362 (N_9362,N_8704,N_8083);
nor U9363 (N_9363,N_8005,N_8722);
nand U9364 (N_9364,N_8515,N_8366);
or U9365 (N_9365,N_8213,N_8236);
and U9366 (N_9366,N_8061,N_8738);
xnor U9367 (N_9367,N_8785,N_8592);
xor U9368 (N_9368,N_8038,N_8569);
xor U9369 (N_9369,N_8845,N_8803);
nand U9370 (N_9370,N_8551,N_8913);
and U9371 (N_9371,N_8949,N_8444);
or U9372 (N_9372,N_8334,N_8643);
nor U9373 (N_9373,N_8747,N_8561);
xor U9374 (N_9374,N_8705,N_8145);
or U9375 (N_9375,N_8056,N_8654);
nand U9376 (N_9376,N_8144,N_8303);
nand U9377 (N_9377,N_8562,N_8826);
or U9378 (N_9378,N_8919,N_8310);
nor U9379 (N_9379,N_8160,N_8421);
nor U9380 (N_9380,N_8519,N_8264);
xnor U9381 (N_9381,N_8564,N_8437);
or U9382 (N_9382,N_8140,N_8339);
or U9383 (N_9383,N_8258,N_8594);
and U9384 (N_9384,N_8734,N_8536);
nand U9385 (N_9385,N_8355,N_8119);
or U9386 (N_9386,N_8950,N_8682);
nor U9387 (N_9387,N_8132,N_8846);
and U9388 (N_9388,N_8761,N_8225);
xnor U9389 (N_9389,N_8300,N_8299);
nand U9390 (N_9390,N_8635,N_8163);
nor U9391 (N_9391,N_8404,N_8510);
or U9392 (N_9392,N_8574,N_8528);
nand U9393 (N_9393,N_8382,N_8537);
nor U9394 (N_9394,N_8321,N_8124);
nor U9395 (N_9395,N_8514,N_8622);
nor U9396 (N_9396,N_8018,N_8443);
nand U9397 (N_9397,N_8701,N_8621);
nor U9398 (N_9398,N_8097,N_8729);
nor U9399 (N_9399,N_8946,N_8908);
nor U9400 (N_9400,N_8259,N_8683);
nor U9401 (N_9401,N_8815,N_8288);
nor U9402 (N_9402,N_8323,N_8157);
and U9403 (N_9403,N_8480,N_8957);
or U9404 (N_9404,N_8902,N_8850);
nand U9405 (N_9405,N_8937,N_8978);
or U9406 (N_9406,N_8546,N_8924);
nand U9407 (N_9407,N_8605,N_8027);
xor U9408 (N_9408,N_8746,N_8398);
xor U9409 (N_9409,N_8523,N_8242);
xnor U9410 (N_9410,N_8359,N_8531);
and U9411 (N_9411,N_8002,N_8388);
or U9412 (N_9412,N_8118,N_8252);
and U9413 (N_9413,N_8482,N_8774);
nand U9414 (N_9414,N_8929,N_8455);
nor U9415 (N_9415,N_8833,N_8070);
nor U9416 (N_9416,N_8789,N_8218);
or U9417 (N_9417,N_8186,N_8733);
or U9418 (N_9418,N_8736,N_8618);
or U9419 (N_9419,N_8513,N_8392);
xor U9420 (N_9420,N_8306,N_8039);
xor U9421 (N_9421,N_8541,N_8647);
nand U9422 (N_9422,N_8997,N_8917);
xor U9423 (N_9423,N_8107,N_8834);
nor U9424 (N_9424,N_8188,N_8980);
nor U9425 (N_9425,N_8262,N_8671);
xnor U9426 (N_9426,N_8532,N_8624);
or U9427 (N_9427,N_8548,N_8796);
and U9428 (N_9428,N_8798,N_8326);
nor U9429 (N_9429,N_8003,N_8694);
xnor U9430 (N_9430,N_8583,N_8476);
and U9431 (N_9431,N_8373,N_8247);
nand U9432 (N_9432,N_8623,N_8914);
or U9433 (N_9433,N_8817,N_8139);
xnor U9434 (N_9434,N_8739,N_8072);
and U9435 (N_9435,N_8369,N_8737);
xnor U9436 (N_9436,N_8238,N_8125);
nor U9437 (N_9437,N_8855,N_8481);
xor U9438 (N_9438,N_8301,N_8471);
nor U9439 (N_9439,N_8724,N_8719);
nand U9440 (N_9440,N_8260,N_8816);
xor U9441 (N_9441,N_8015,N_8269);
and U9442 (N_9442,N_8172,N_8111);
xnor U9443 (N_9443,N_8680,N_8047);
or U9444 (N_9444,N_8524,N_8706);
xor U9445 (N_9445,N_8473,N_8006);
nand U9446 (N_9446,N_8116,N_8861);
nand U9447 (N_9447,N_8060,N_8849);
nor U9448 (N_9448,N_8871,N_8368);
or U9449 (N_9449,N_8081,N_8503);
xor U9450 (N_9450,N_8782,N_8010);
nor U9451 (N_9451,N_8344,N_8552);
nor U9452 (N_9452,N_8699,N_8901);
or U9453 (N_9453,N_8851,N_8436);
or U9454 (N_9454,N_8878,N_8640);
nor U9455 (N_9455,N_8121,N_8863);
nand U9456 (N_9456,N_8452,N_8835);
and U9457 (N_9457,N_8141,N_8068);
and U9458 (N_9458,N_8714,N_8191);
and U9459 (N_9459,N_8200,N_8942);
nor U9460 (N_9460,N_8332,N_8454);
nand U9461 (N_9461,N_8434,N_8131);
and U9462 (N_9462,N_8239,N_8820);
and U9463 (N_9463,N_8234,N_8008);
nand U9464 (N_9464,N_8844,N_8297);
nor U9465 (N_9465,N_8051,N_8572);
or U9466 (N_9466,N_8987,N_8757);
nand U9467 (N_9467,N_8856,N_8963);
nor U9468 (N_9468,N_8598,N_8771);
and U9469 (N_9469,N_8936,N_8922);
nand U9470 (N_9470,N_8530,N_8732);
and U9471 (N_9471,N_8322,N_8329);
nand U9472 (N_9472,N_8054,N_8646);
or U9473 (N_9473,N_8672,N_8697);
or U9474 (N_9474,N_8550,N_8698);
xor U9475 (N_9475,N_8268,N_8137);
or U9476 (N_9476,N_8263,N_8312);
nor U9477 (N_9477,N_8464,N_8526);
or U9478 (N_9478,N_8298,N_8812);
nand U9479 (N_9479,N_8280,N_8657);
and U9480 (N_9480,N_8656,N_8375);
xor U9481 (N_9481,N_8517,N_8410);
xor U9482 (N_9482,N_8354,N_8636);
nand U9483 (N_9483,N_8468,N_8492);
nand U9484 (N_9484,N_8554,N_8261);
or U9485 (N_9485,N_8187,N_8993);
or U9486 (N_9486,N_8614,N_8688);
xnor U9487 (N_9487,N_8179,N_8022);
or U9488 (N_9488,N_8687,N_8948);
or U9489 (N_9489,N_8296,N_8351);
xor U9490 (N_9490,N_8965,N_8506);
nand U9491 (N_9491,N_8700,N_8063);
or U9492 (N_9492,N_8559,N_8748);
xnor U9493 (N_9493,N_8466,N_8831);
xnor U9494 (N_9494,N_8823,N_8723);
nand U9495 (N_9495,N_8668,N_8203);
nand U9496 (N_9496,N_8504,N_8148);
nor U9497 (N_9497,N_8712,N_8889);
or U9498 (N_9498,N_8792,N_8173);
or U9499 (N_9499,N_8651,N_8458);
xnor U9500 (N_9500,N_8613,N_8619);
xnor U9501 (N_9501,N_8747,N_8669);
or U9502 (N_9502,N_8530,N_8857);
nand U9503 (N_9503,N_8291,N_8539);
or U9504 (N_9504,N_8731,N_8453);
xnor U9505 (N_9505,N_8831,N_8223);
and U9506 (N_9506,N_8982,N_8799);
nand U9507 (N_9507,N_8837,N_8466);
and U9508 (N_9508,N_8289,N_8416);
xor U9509 (N_9509,N_8892,N_8769);
or U9510 (N_9510,N_8250,N_8639);
xor U9511 (N_9511,N_8089,N_8096);
or U9512 (N_9512,N_8526,N_8729);
and U9513 (N_9513,N_8513,N_8327);
nor U9514 (N_9514,N_8863,N_8328);
xor U9515 (N_9515,N_8255,N_8281);
nor U9516 (N_9516,N_8066,N_8082);
or U9517 (N_9517,N_8908,N_8263);
nand U9518 (N_9518,N_8723,N_8338);
and U9519 (N_9519,N_8590,N_8271);
and U9520 (N_9520,N_8193,N_8573);
or U9521 (N_9521,N_8326,N_8882);
nand U9522 (N_9522,N_8203,N_8828);
or U9523 (N_9523,N_8477,N_8022);
xor U9524 (N_9524,N_8599,N_8844);
nand U9525 (N_9525,N_8723,N_8828);
and U9526 (N_9526,N_8202,N_8181);
nor U9527 (N_9527,N_8959,N_8526);
or U9528 (N_9528,N_8284,N_8620);
or U9529 (N_9529,N_8933,N_8927);
xnor U9530 (N_9530,N_8440,N_8483);
nor U9531 (N_9531,N_8471,N_8041);
or U9532 (N_9532,N_8917,N_8603);
xor U9533 (N_9533,N_8274,N_8608);
and U9534 (N_9534,N_8954,N_8718);
nor U9535 (N_9535,N_8607,N_8372);
and U9536 (N_9536,N_8686,N_8054);
nand U9537 (N_9537,N_8366,N_8632);
or U9538 (N_9538,N_8790,N_8888);
or U9539 (N_9539,N_8423,N_8316);
nor U9540 (N_9540,N_8427,N_8696);
xnor U9541 (N_9541,N_8979,N_8409);
and U9542 (N_9542,N_8335,N_8311);
nand U9543 (N_9543,N_8452,N_8750);
nand U9544 (N_9544,N_8314,N_8335);
nor U9545 (N_9545,N_8014,N_8515);
nor U9546 (N_9546,N_8743,N_8712);
and U9547 (N_9547,N_8344,N_8393);
and U9548 (N_9548,N_8828,N_8632);
nor U9549 (N_9549,N_8277,N_8385);
xor U9550 (N_9550,N_8628,N_8417);
xnor U9551 (N_9551,N_8736,N_8756);
xor U9552 (N_9552,N_8146,N_8239);
xor U9553 (N_9553,N_8294,N_8150);
nand U9554 (N_9554,N_8197,N_8157);
xor U9555 (N_9555,N_8129,N_8453);
nand U9556 (N_9556,N_8677,N_8982);
nor U9557 (N_9557,N_8613,N_8559);
xnor U9558 (N_9558,N_8543,N_8306);
or U9559 (N_9559,N_8680,N_8096);
xnor U9560 (N_9560,N_8148,N_8900);
or U9561 (N_9561,N_8935,N_8477);
and U9562 (N_9562,N_8948,N_8218);
or U9563 (N_9563,N_8221,N_8167);
xnor U9564 (N_9564,N_8761,N_8428);
and U9565 (N_9565,N_8949,N_8303);
nand U9566 (N_9566,N_8558,N_8629);
and U9567 (N_9567,N_8451,N_8741);
and U9568 (N_9568,N_8910,N_8657);
nand U9569 (N_9569,N_8512,N_8509);
nor U9570 (N_9570,N_8502,N_8715);
nor U9571 (N_9571,N_8187,N_8470);
xor U9572 (N_9572,N_8151,N_8944);
and U9573 (N_9573,N_8844,N_8506);
xnor U9574 (N_9574,N_8078,N_8796);
nand U9575 (N_9575,N_8802,N_8915);
or U9576 (N_9576,N_8640,N_8361);
xnor U9577 (N_9577,N_8257,N_8429);
and U9578 (N_9578,N_8738,N_8644);
nand U9579 (N_9579,N_8173,N_8417);
and U9580 (N_9580,N_8182,N_8190);
nor U9581 (N_9581,N_8434,N_8165);
xor U9582 (N_9582,N_8832,N_8741);
nor U9583 (N_9583,N_8845,N_8753);
xnor U9584 (N_9584,N_8485,N_8869);
and U9585 (N_9585,N_8098,N_8177);
nand U9586 (N_9586,N_8951,N_8547);
nand U9587 (N_9587,N_8322,N_8038);
nor U9588 (N_9588,N_8172,N_8493);
or U9589 (N_9589,N_8407,N_8995);
or U9590 (N_9590,N_8922,N_8094);
and U9591 (N_9591,N_8367,N_8964);
nand U9592 (N_9592,N_8553,N_8954);
and U9593 (N_9593,N_8377,N_8012);
and U9594 (N_9594,N_8346,N_8533);
nor U9595 (N_9595,N_8434,N_8085);
xor U9596 (N_9596,N_8742,N_8944);
nor U9597 (N_9597,N_8655,N_8562);
nor U9598 (N_9598,N_8310,N_8040);
xor U9599 (N_9599,N_8140,N_8251);
xnor U9600 (N_9600,N_8123,N_8985);
nor U9601 (N_9601,N_8243,N_8797);
nor U9602 (N_9602,N_8979,N_8346);
and U9603 (N_9603,N_8442,N_8577);
or U9604 (N_9604,N_8191,N_8696);
or U9605 (N_9605,N_8886,N_8208);
and U9606 (N_9606,N_8279,N_8748);
xor U9607 (N_9607,N_8075,N_8899);
or U9608 (N_9608,N_8569,N_8056);
or U9609 (N_9609,N_8710,N_8985);
or U9610 (N_9610,N_8737,N_8262);
nand U9611 (N_9611,N_8112,N_8778);
nor U9612 (N_9612,N_8698,N_8280);
nor U9613 (N_9613,N_8409,N_8167);
xor U9614 (N_9614,N_8403,N_8844);
or U9615 (N_9615,N_8769,N_8797);
and U9616 (N_9616,N_8647,N_8383);
nand U9617 (N_9617,N_8843,N_8036);
nor U9618 (N_9618,N_8449,N_8622);
xnor U9619 (N_9619,N_8620,N_8085);
and U9620 (N_9620,N_8195,N_8413);
xnor U9621 (N_9621,N_8146,N_8561);
or U9622 (N_9622,N_8299,N_8952);
nand U9623 (N_9623,N_8005,N_8460);
nand U9624 (N_9624,N_8947,N_8378);
xnor U9625 (N_9625,N_8782,N_8610);
nor U9626 (N_9626,N_8847,N_8778);
nand U9627 (N_9627,N_8966,N_8437);
xnor U9628 (N_9628,N_8117,N_8126);
xnor U9629 (N_9629,N_8761,N_8661);
xnor U9630 (N_9630,N_8574,N_8442);
nor U9631 (N_9631,N_8558,N_8072);
nand U9632 (N_9632,N_8275,N_8778);
xnor U9633 (N_9633,N_8678,N_8702);
xnor U9634 (N_9634,N_8050,N_8293);
or U9635 (N_9635,N_8387,N_8457);
nor U9636 (N_9636,N_8911,N_8812);
xor U9637 (N_9637,N_8937,N_8257);
xor U9638 (N_9638,N_8350,N_8302);
or U9639 (N_9639,N_8374,N_8341);
or U9640 (N_9640,N_8921,N_8456);
xnor U9641 (N_9641,N_8931,N_8054);
nor U9642 (N_9642,N_8505,N_8085);
nand U9643 (N_9643,N_8063,N_8371);
xnor U9644 (N_9644,N_8319,N_8572);
or U9645 (N_9645,N_8826,N_8263);
nor U9646 (N_9646,N_8312,N_8385);
and U9647 (N_9647,N_8012,N_8501);
nand U9648 (N_9648,N_8583,N_8496);
nor U9649 (N_9649,N_8551,N_8716);
and U9650 (N_9650,N_8134,N_8033);
nor U9651 (N_9651,N_8275,N_8793);
or U9652 (N_9652,N_8641,N_8099);
and U9653 (N_9653,N_8950,N_8469);
xor U9654 (N_9654,N_8389,N_8758);
and U9655 (N_9655,N_8852,N_8561);
xnor U9656 (N_9656,N_8501,N_8677);
and U9657 (N_9657,N_8752,N_8340);
nor U9658 (N_9658,N_8439,N_8917);
nor U9659 (N_9659,N_8580,N_8698);
or U9660 (N_9660,N_8038,N_8916);
xor U9661 (N_9661,N_8037,N_8112);
nor U9662 (N_9662,N_8268,N_8503);
nor U9663 (N_9663,N_8802,N_8241);
nand U9664 (N_9664,N_8740,N_8774);
and U9665 (N_9665,N_8445,N_8742);
or U9666 (N_9666,N_8449,N_8864);
nand U9667 (N_9667,N_8703,N_8315);
nor U9668 (N_9668,N_8750,N_8645);
and U9669 (N_9669,N_8431,N_8043);
nand U9670 (N_9670,N_8991,N_8100);
or U9671 (N_9671,N_8962,N_8796);
and U9672 (N_9672,N_8368,N_8514);
or U9673 (N_9673,N_8345,N_8222);
nor U9674 (N_9674,N_8144,N_8013);
xnor U9675 (N_9675,N_8532,N_8895);
nor U9676 (N_9676,N_8114,N_8629);
or U9677 (N_9677,N_8652,N_8793);
xnor U9678 (N_9678,N_8531,N_8430);
and U9679 (N_9679,N_8154,N_8602);
xnor U9680 (N_9680,N_8434,N_8028);
or U9681 (N_9681,N_8745,N_8732);
xnor U9682 (N_9682,N_8941,N_8852);
nand U9683 (N_9683,N_8796,N_8154);
and U9684 (N_9684,N_8013,N_8641);
or U9685 (N_9685,N_8164,N_8131);
nor U9686 (N_9686,N_8054,N_8911);
and U9687 (N_9687,N_8461,N_8749);
or U9688 (N_9688,N_8883,N_8795);
nor U9689 (N_9689,N_8019,N_8071);
or U9690 (N_9690,N_8822,N_8039);
xnor U9691 (N_9691,N_8935,N_8260);
or U9692 (N_9692,N_8191,N_8762);
nand U9693 (N_9693,N_8513,N_8785);
nor U9694 (N_9694,N_8083,N_8632);
and U9695 (N_9695,N_8165,N_8260);
xnor U9696 (N_9696,N_8339,N_8550);
nand U9697 (N_9697,N_8620,N_8480);
or U9698 (N_9698,N_8057,N_8243);
and U9699 (N_9699,N_8934,N_8551);
and U9700 (N_9700,N_8502,N_8681);
or U9701 (N_9701,N_8164,N_8161);
nor U9702 (N_9702,N_8442,N_8712);
and U9703 (N_9703,N_8555,N_8881);
nand U9704 (N_9704,N_8736,N_8371);
nand U9705 (N_9705,N_8982,N_8121);
nand U9706 (N_9706,N_8793,N_8913);
nand U9707 (N_9707,N_8215,N_8253);
and U9708 (N_9708,N_8353,N_8904);
nand U9709 (N_9709,N_8706,N_8743);
nand U9710 (N_9710,N_8077,N_8185);
and U9711 (N_9711,N_8550,N_8655);
xor U9712 (N_9712,N_8496,N_8228);
xnor U9713 (N_9713,N_8179,N_8359);
nand U9714 (N_9714,N_8949,N_8792);
nand U9715 (N_9715,N_8988,N_8736);
or U9716 (N_9716,N_8304,N_8293);
nand U9717 (N_9717,N_8610,N_8325);
nor U9718 (N_9718,N_8756,N_8760);
and U9719 (N_9719,N_8988,N_8141);
or U9720 (N_9720,N_8151,N_8522);
or U9721 (N_9721,N_8437,N_8468);
and U9722 (N_9722,N_8157,N_8892);
xnor U9723 (N_9723,N_8042,N_8634);
xor U9724 (N_9724,N_8398,N_8347);
nand U9725 (N_9725,N_8794,N_8661);
nor U9726 (N_9726,N_8728,N_8157);
xnor U9727 (N_9727,N_8538,N_8197);
xnor U9728 (N_9728,N_8432,N_8338);
nor U9729 (N_9729,N_8798,N_8055);
and U9730 (N_9730,N_8294,N_8592);
nor U9731 (N_9731,N_8573,N_8247);
xor U9732 (N_9732,N_8293,N_8343);
xor U9733 (N_9733,N_8919,N_8800);
or U9734 (N_9734,N_8109,N_8192);
nand U9735 (N_9735,N_8091,N_8510);
xnor U9736 (N_9736,N_8785,N_8228);
xor U9737 (N_9737,N_8859,N_8665);
and U9738 (N_9738,N_8367,N_8074);
and U9739 (N_9739,N_8751,N_8771);
xnor U9740 (N_9740,N_8929,N_8767);
nor U9741 (N_9741,N_8576,N_8293);
or U9742 (N_9742,N_8287,N_8457);
nand U9743 (N_9743,N_8245,N_8576);
xnor U9744 (N_9744,N_8735,N_8681);
nand U9745 (N_9745,N_8949,N_8186);
or U9746 (N_9746,N_8687,N_8886);
and U9747 (N_9747,N_8331,N_8691);
or U9748 (N_9748,N_8650,N_8595);
nand U9749 (N_9749,N_8073,N_8392);
and U9750 (N_9750,N_8321,N_8634);
or U9751 (N_9751,N_8620,N_8834);
or U9752 (N_9752,N_8710,N_8094);
and U9753 (N_9753,N_8492,N_8342);
nand U9754 (N_9754,N_8206,N_8928);
or U9755 (N_9755,N_8808,N_8660);
and U9756 (N_9756,N_8365,N_8129);
and U9757 (N_9757,N_8815,N_8657);
and U9758 (N_9758,N_8811,N_8681);
and U9759 (N_9759,N_8779,N_8801);
or U9760 (N_9760,N_8073,N_8539);
nor U9761 (N_9761,N_8723,N_8363);
or U9762 (N_9762,N_8846,N_8560);
xnor U9763 (N_9763,N_8380,N_8816);
nand U9764 (N_9764,N_8163,N_8676);
nor U9765 (N_9765,N_8158,N_8090);
nand U9766 (N_9766,N_8846,N_8374);
or U9767 (N_9767,N_8481,N_8889);
nand U9768 (N_9768,N_8229,N_8401);
nor U9769 (N_9769,N_8736,N_8255);
nand U9770 (N_9770,N_8723,N_8135);
and U9771 (N_9771,N_8624,N_8401);
or U9772 (N_9772,N_8796,N_8993);
nand U9773 (N_9773,N_8035,N_8752);
and U9774 (N_9774,N_8523,N_8514);
nand U9775 (N_9775,N_8696,N_8133);
nand U9776 (N_9776,N_8859,N_8730);
nor U9777 (N_9777,N_8493,N_8831);
and U9778 (N_9778,N_8602,N_8957);
or U9779 (N_9779,N_8258,N_8350);
xor U9780 (N_9780,N_8145,N_8671);
nor U9781 (N_9781,N_8031,N_8986);
nor U9782 (N_9782,N_8124,N_8487);
nor U9783 (N_9783,N_8811,N_8161);
xnor U9784 (N_9784,N_8750,N_8039);
and U9785 (N_9785,N_8743,N_8349);
xor U9786 (N_9786,N_8100,N_8903);
nor U9787 (N_9787,N_8828,N_8015);
and U9788 (N_9788,N_8969,N_8147);
and U9789 (N_9789,N_8863,N_8276);
xor U9790 (N_9790,N_8482,N_8755);
and U9791 (N_9791,N_8254,N_8708);
xnor U9792 (N_9792,N_8152,N_8997);
nand U9793 (N_9793,N_8772,N_8364);
or U9794 (N_9794,N_8911,N_8339);
and U9795 (N_9795,N_8215,N_8703);
xnor U9796 (N_9796,N_8627,N_8718);
xor U9797 (N_9797,N_8152,N_8179);
nor U9798 (N_9798,N_8851,N_8515);
nor U9799 (N_9799,N_8037,N_8233);
nor U9800 (N_9800,N_8230,N_8558);
or U9801 (N_9801,N_8711,N_8187);
or U9802 (N_9802,N_8357,N_8805);
and U9803 (N_9803,N_8082,N_8908);
nand U9804 (N_9804,N_8512,N_8853);
or U9805 (N_9805,N_8667,N_8775);
and U9806 (N_9806,N_8589,N_8593);
or U9807 (N_9807,N_8591,N_8629);
nor U9808 (N_9808,N_8451,N_8909);
xor U9809 (N_9809,N_8269,N_8201);
and U9810 (N_9810,N_8754,N_8789);
nor U9811 (N_9811,N_8251,N_8050);
xor U9812 (N_9812,N_8131,N_8851);
or U9813 (N_9813,N_8753,N_8836);
nand U9814 (N_9814,N_8648,N_8261);
and U9815 (N_9815,N_8605,N_8595);
nor U9816 (N_9816,N_8063,N_8255);
and U9817 (N_9817,N_8701,N_8371);
and U9818 (N_9818,N_8150,N_8646);
xnor U9819 (N_9819,N_8122,N_8647);
nor U9820 (N_9820,N_8475,N_8866);
and U9821 (N_9821,N_8648,N_8389);
nor U9822 (N_9822,N_8087,N_8024);
nor U9823 (N_9823,N_8008,N_8950);
and U9824 (N_9824,N_8877,N_8181);
xnor U9825 (N_9825,N_8446,N_8964);
and U9826 (N_9826,N_8030,N_8728);
and U9827 (N_9827,N_8261,N_8910);
and U9828 (N_9828,N_8334,N_8102);
nand U9829 (N_9829,N_8863,N_8304);
nand U9830 (N_9830,N_8863,N_8425);
nand U9831 (N_9831,N_8182,N_8967);
nand U9832 (N_9832,N_8177,N_8401);
or U9833 (N_9833,N_8366,N_8425);
nand U9834 (N_9834,N_8182,N_8879);
xnor U9835 (N_9835,N_8985,N_8370);
and U9836 (N_9836,N_8709,N_8339);
or U9837 (N_9837,N_8809,N_8619);
or U9838 (N_9838,N_8568,N_8140);
or U9839 (N_9839,N_8127,N_8137);
nand U9840 (N_9840,N_8034,N_8775);
and U9841 (N_9841,N_8761,N_8454);
xnor U9842 (N_9842,N_8479,N_8002);
xnor U9843 (N_9843,N_8040,N_8461);
or U9844 (N_9844,N_8345,N_8470);
nand U9845 (N_9845,N_8646,N_8267);
or U9846 (N_9846,N_8396,N_8145);
and U9847 (N_9847,N_8030,N_8410);
or U9848 (N_9848,N_8107,N_8986);
nor U9849 (N_9849,N_8215,N_8767);
nor U9850 (N_9850,N_8177,N_8179);
nand U9851 (N_9851,N_8712,N_8019);
nor U9852 (N_9852,N_8408,N_8241);
or U9853 (N_9853,N_8589,N_8493);
and U9854 (N_9854,N_8471,N_8414);
or U9855 (N_9855,N_8684,N_8693);
nand U9856 (N_9856,N_8196,N_8355);
and U9857 (N_9857,N_8806,N_8056);
nand U9858 (N_9858,N_8268,N_8723);
nor U9859 (N_9859,N_8480,N_8925);
nor U9860 (N_9860,N_8098,N_8240);
nand U9861 (N_9861,N_8332,N_8342);
xnor U9862 (N_9862,N_8037,N_8256);
xor U9863 (N_9863,N_8695,N_8018);
nand U9864 (N_9864,N_8087,N_8863);
and U9865 (N_9865,N_8861,N_8324);
nor U9866 (N_9866,N_8347,N_8441);
nor U9867 (N_9867,N_8300,N_8420);
xor U9868 (N_9868,N_8745,N_8784);
nand U9869 (N_9869,N_8077,N_8886);
nand U9870 (N_9870,N_8255,N_8252);
and U9871 (N_9871,N_8980,N_8433);
xnor U9872 (N_9872,N_8022,N_8167);
and U9873 (N_9873,N_8513,N_8571);
and U9874 (N_9874,N_8592,N_8070);
or U9875 (N_9875,N_8916,N_8268);
and U9876 (N_9876,N_8060,N_8104);
or U9877 (N_9877,N_8315,N_8988);
nor U9878 (N_9878,N_8621,N_8152);
xnor U9879 (N_9879,N_8209,N_8108);
or U9880 (N_9880,N_8745,N_8903);
or U9881 (N_9881,N_8462,N_8490);
nor U9882 (N_9882,N_8022,N_8496);
nand U9883 (N_9883,N_8437,N_8742);
and U9884 (N_9884,N_8960,N_8651);
or U9885 (N_9885,N_8856,N_8340);
or U9886 (N_9886,N_8228,N_8136);
nand U9887 (N_9887,N_8082,N_8531);
xor U9888 (N_9888,N_8415,N_8450);
or U9889 (N_9889,N_8773,N_8404);
nor U9890 (N_9890,N_8665,N_8433);
or U9891 (N_9891,N_8425,N_8873);
xor U9892 (N_9892,N_8303,N_8123);
nand U9893 (N_9893,N_8661,N_8992);
xnor U9894 (N_9894,N_8911,N_8993);
or U9895 (N_9895,N_8315,N_8911);
nor U9896 (N_9896,N_8729,N_8838);
nand U9897 (N_9897,N_8533,N_8785);
nand U9898 (N_9898,N_8649,N_8725);
and U9899 (N_9899,N_8772,N_8988);
nor U9900 (N_9900,N_8292,N_8285);
and U9901 (N_9901,N_8234,N_8807);
and U9902 (N_9902,N_8801,N_8666);
or U9903 (N_9903,N_8136,N_8722);
nand U9904 (N_9904,N_8735,N_8137);
nand U9905 (N_9905,N_8951,N_8359);
xor U9906 (N_9906,N_8950,N_8327);
or U9907 (N_9907,N_8918,N_8294);
nand U9908 (N_9908,N_8761,N_8152);
xor U9909 (N_9909,N_8625,N_8706);
xor U9910 (N_9910,N_8834,N_8398);
or U9911 (N_9911,N_8166,N_8741);
and U9912 (N_9912,N_8960,N_8756);
and U9913 (N_9913,N_8530,N_8869);
nand U9914 (N_9914,N_8186,N_8312);
xor U9915 (N_9915,N_8267,N_8000);
xnor U9916 (N_9916,N_8971,N_8801);
nand U9917 (N_9917,N_8245,N_8163);
and U9918 (N_9918,N_8848,N_8349);
or U9919 (N_9919,N_8983,N_8228);
nor U9920 (N_9920,N_8210,N_8469);
and U9921 (N_9921,N_8569,N_8753);
or U9922 (N_9922,N_8102,N_8332);
nand U9923 (N_9923,N_8916,N_8596);
or U9924 (N_9924,N_8569,N_8361);
nand U9925 (N_9925,N_8244,N_8545);
nand U9926 (N_9926,N_8300,N_8153);
nor U9927 (N_9927,N_8185,N_8854);
nand U9928 (N_9928,N_8602,N_8191);
xnor U9929 (N_9929,N_8042,N_8272);
nand U9930 (N_9930,N_8483,N_8342);
nand U9931 (N_9931,N_8459,N_8435);
or U9932 (N_9932,N_8142,N_8281);
nor U9933 (N_9933,N_8210,N_8507);
nand U9934 (N_9934,N_8468,N_8192);
or U9935 (N_9935,N_8687,N_8814);
or U9936 (N_9936,N_8281,N_8832);
nand U9937 (N_9937,N_8840,N_8251);
and U9938 (N_9938,N_8072,N_8311);
and U9939 (N_9939,N_8940,N_8200);
nand U9940 (N_9940,N_8050,N_8792);
or U9941 (N_9941,N_8006,N_8009);
nor U9942 (N_9942,N_8303,N_8043);
nor U9943 (N_9943,N_8309,N_8846);
nand U9944 (N_9944,N_8141,N_8779);
nand U9945 (N_9945,N_8431,N_8655);
nor U9946 (N_9946,N_8565,N_8366);
or U9947 (N_9947,N_8772,N_8648);
xnor U9948 (N_9948,N_8927,N_8042);
and U9949 (N_9949,N_8925,N_8259);
nor U9950 (N_9950,N_8252,N_8658);
or U9951 (N_9951,N_8465,N_8613);
or U9952 (N_9952,N_8395,N_8880);
nor U9953 (N_9953,N_8519,N_8071);
or U9954 (N_9954,N_8782,N_8190);
xor U9955 (N_9955,N_8142,N_8008);
and U9956 (N_9956,N_8358,N_8002);
nor U9957 (N_9957,N_8628,N_8821);
nand U9958 (N_9958,N_8572,N_8926);
xnor U9959 (N_9959,N_8558,N_8874);
and U9960 (N_9960,N_8122,N_8082);
and U9961 (N_9961,N_8997,N_8546);
nand U9962 (N_9962,N_8505,N_8308);
or U9963 (N_9963,N_8534,N_8971);
or U9964 (N_9964,N_8670,N_8957);
or U9965 (N_9965,N_8013,N_8876);
xor U9966 (N_9966,N_8718,N_8783);
nand U9967 (N_9967,N_8074,N_8808);
xnor U9968 (N_9968,N_8560,N_8152);
nand U9969 (N_9969,N_8442,N_8010);
and U9970 (N_9970,N_8907,N_8650);
nand U9971 (N_9971,N_8294,N_8704);
nand U9972 (N_9972,N_8886,N_8026);
and U9973 (N_9973,N_8865,N_8550);
and U9974 (N_9974,N_8237,N_8758);
and U9975 (N_9975,N_8539,N_8943);
nand U9976 (N_9976,N_8993,N_8520);
or U9977 (N_9977,N_8342,N_8631);
nand U9978 (N_9978,N_8914,N_8351);
nand U9979 (N_9979,N_8404,N_8137);
nand U9980 (N_9980,N_8706,N_8166);
xnor U9981 (N_9981,N_8984,N_8073);
nor U9982 (N_9982,N_8115,N_8217);
or U9983 (N_9983,N_8920,N_8405);
nand U9984 (N_9984,N_8193,N_8500);
xor U9985 (N_9985,N_8827,N_8093);
or U9986 (N_9986,N_8506,N_8505);
nor U9987 (N_9987,N_8029,N_8459);
or U9988 (N_9988,N_8829,N_8328);
or U9989 (N_9989,N_8415,N_8523);
nand U9990 (N_9990,N_8063,N_8650);
or U9991 (N_9991,N_8614,N_8951);
nand U9992 (N_9992,N_8925,N_8824);
or U9993 (N_9993,N_8803,N_8056);
xor U9994 (N_9994,N_8646,N_8723);
or U9995 (N_9995,N_8606,N_8452);
and U9996 (N_9996,N_8498,N_8292);
or U9997 (N_9997,N_8174,N_8646);
xor U9998 (N_9998,N_8442,N_8029);
xnor U9999 (N_9999,N_8558,N_8577);
nand U10000 (N_10000,N_9225,N_9296);
nand U10001 (N_10001,N_9328,N_9791);
and U10002 (N_10002,N_9977,N_9330);
xor U10003 (N_10003,N_9906,N_9024);
xnor U10004 (N_10004,N_9232,N_9574);
or U10005 (N_10005,N_9316,N_9251);
nor U10006 (N_10006,N_9882,N_9040);
nor U10007 (N_10007,N_9527,N_9540);
nor U10008 (N_10008,N_9255,N_9928);
xor U10009 (N_10009,N_9089,N_9781);
nand U10010 (N_10010,N_9116,N_9027);
and U10011 (N_10011,N_9837,N_9698);
nor U10012 (N_10012,N_9431,N_9656);
xnor U10013 (N_10013,N_9158,N_9041);
or U10014 (N_10014,N_9471,N_9575);
nand U10015 (N_10015,N_9507,N_9515);
or U10016 (N_10016,N_9810,N_9758);
nand U10017 (N_10017,N_9353,N_9614);
nand U10018 (N_10018,N_9848,N_9772);
and U10019 (N_10019,N_9458,N_9520);
xor U10020 (N_10020,N_9556,N_9270);
and U10021 (N_10021,N_9466,N_9121);
nand U10022 (N_10022,N_9864,N_9892);
xnor U10023 (N_10023,N_9504,N_9418);
and U10024 (N_10024,N_9413,N_9243);
nor U10025 (N_10025,N_9385,N_9736);
or U10026 (N_10026,N_9167,N_9635);
nor U10027 (N_10027,N_9339,N_9198);
and U10028 (N_10028,N_9846,N_9669);
xor U10029 (N_10029,N_9469,N_9467);
xnor U10030 (N_10030,N_9546,N_9072);
xor U10031 (N_10031,N_9788,N_9051);
nor U10032 (N_10032,N_9658,N_9675);
and U10033 (N_10033,N_9919,N_9541);
xor U10034 (N_10034,N_9048,N_9094);
nor U10035 (N_10035,N_9548,N_9025);
and U10036 (N_10036,N_9529,N_9082);
or U10037 (N_10037,N_9833,N_9213);
and U10038 (N_10038,N_9861,N_9902);
or U10039 (N_10039,N_9602,N_9986);
and U10040 (N_10040,N_9755,N_9484);
xor U10041 (N_10041,N_9227,N_9276);
xnor U10042 (N_10042,N_9445,N_9064);
nor U10043 (N_10043,N_9887,N_9254);
xnor U10044 (N_10044,N_9248,N_9775);
or U10045 (N_10045,N_9049,N_9081);
and U10046 (N_10046,N_9827,N_9065);
or U10047 (N_10047,N_9766,N_9134);
xor U10048 (N_10048,N_9015,N_9921);
or U10049 (N_10049,N_9624,N_9849);
or U10050 (N_10050,N_9436,N_9008);
nand U10051 (N_10051,N_9370,N_9073);
nor U10052 (N_10052,N_9007,N_9274);
nor U10053 (N_10053,N_9231,N_9731);
and U10054 (N_10054,N_9976,N_9118);
or U10055 (N_10055,N_9311,N_9267);
or U10056 (N_10056,N_9320,N_9351);
nor U10057 (N_10057,N_9149,N_9982);
nor U10058 (N_10058,N_9376,N_9787);
and U10059 (N_10059,N_9526,N_9355);
xnor U10060 (N_10060,N_9971,N_9918);
nor U10061 (N_10061,N_9217,N_9647);
xnor U10062 (N_10062,N_9240,N_9528);
and U10063 (N_10063,N_9443,N_9704);
xnor U10064 (N_10064,N_9125,N_9641);
xnor U10065 (N_10065,N_9760,N_9841);
nor U10066 (N_10066,N_9818,N_9741);
nor U10067 (N_10067,N_9927,N_9824);
or U10068 (N_10068,N_9776,N_9830);
or U10069 (N_10069,N_9416,N_9714);
and U10070 (N_10070,N_9703,N_9613);
nand U10071 (N_10071,N_9984,N_9797);
or U10072 (N_10072,N_9054,N_9949);
or U10073 (N_10073,N_9510,N_9067);
nor U10074 (N_10074,N_9636,N_9952);
or U10075 (N_10075,N_9807,N_9399);
xnor U10076 (N_10076,N_9439,N_9811);
and U10077 (N_10077,N_9071,N_9002);
and U10078 (N_10078,N_9687,N_9185);
and U10079 (N_10079,N_9196,N_9990);
xor U10080 (N_10080,N_9281,N_9260);
or U10081 (N_10081,N_9972,N_9562);
nor U10082 (N_10082,N_9131,N_9293);
and U10083 (N_10083,N_9543,N_9674);
and U10084 (N_10084,N_9107,N_9324);
or U10085 (N_10085,N_9172,N_9177);
nor U10086 (N_10086,N_9113,N_9665);
nor U10087 (N_10087,N_9211,N_9866);
xnor U10088 (N_10088,N_9135,N_9059);
nand U10089 (N_10089,N_9045,N_9893);
and U10090 (N_10090,N_9907,N_9783);
nand U10091 (N_10091,N_9657,N_9419);
xor U10092 (N_10092,N_9875,N_9224);
or U10093 (N_10093,N_9967,N_9676);
or U10094 (N_10094,N_9259,N_9909);
nor U10095 (N_10095,N_9444,N_9537);
nor U10096 (N_10096,N_9937,N_9105);
xor U10097 (N_10097,N_9905,N_9076);
nor U10098 (N_10098,N_9568,N_9934);
xnor U10099 (N_10099,N_9156,N_9442);
xor U10100 (N_10100,N_9499,N_9924);
xor U10101 (N_10101,N_9843,N_9680);
nor U10102 (N_10102,N_9662,N_9401);
xnor U10103 (N_10103,N_9237,N_9447);
nand U10104 (N_10104,N_9157,N_9142);
or U10105 (N_10105,N_9070,N_9479);
xor U10106 (N_10106,N_9367,N_9743);
xnor U10107 (N_10107,N_9085,N_9075);
or U10108 (N_10108,N_9190,N_9119);
nor U10109 (N_10109,N_9314,N_9753);
nand U10110 (N_10110,N_9572,N_9816);
nor U10111 (N_10111,N_9285,N_9997);
and U10112 (N_10112,N_9757,N_9554);
xnor U10113 (N_10113,N_9795,N_9481);
xnor U10114 (N_10114,N_9179,N_9470);
or U10115 (N_10115,N_9212,N_9994);
nor U10116 (N_10116,N_9363,N_9505);
or U10117 (N_10117,N_9622,N_9873);
nor U10118 (N_10118,N_9749,N_9813);
xor U10119 (N_10119,N_9646,N_9335);
xnor U10120 (N_10120,N_9780,N_9516);
or U10121 (N_10121,N_9343,N_9784);
or U10122 (N_10122,N_9970,N_9701);
xor U10123 (N_10123,N_9078,N_9410);
or U10124 (N_10124,N_9751,N_9607);
nor U10125 (N_10125,N_9062,N_9136);
nor U10126 (N_10126,N_9171,N_9258);
nor U10127 (N_10127,N_9836,N_9181);
nor U10128 (N_10128,N_9069,N_9186);
nor U10129 (N_10129,N_9911,N_9029);
and U10130 (N_10130,N_9290,N_9677);
nor U10131 (N_10131,N_9139,N_9835);
and U10132 (N_10132,N_9277,N_9730);
and U10133 (N_10133,N_9241,N_9345);
or U10134 (N_10134,N_9310,N_9295);
and U10135 (N_10135,N_9037,N_9869);
xnor U10136 (N_10136,N_9803,N_9618);
nand U10137 (N_10137,N_9796,N_9464);
nand U10138 (N_10138,N_9299,N_9151);
and U10139 (N_10139,N_9583,N_9995);
and U10140 (N_10140,N_9492,N_9140);
nor U10141 (N_10141,N_9739,N_9438);
nand U10142 (N_10142,N_9518,N_9182);
nand U10143 (N_10143,N_9493,N_9154);
or U10144 (N_10144,N_9983,N_9216);
xor U10145 (N_10145,N_9723,N_9621);
or U10146 (N_10146,N_9943,N_9959);
nand U10147 (N_10147,N_9592,N_9111);
nor U10148 (N_10148,N_9397,N_9903);
xor U10149 (N_10149,N_9551,N_9782);
nand U10150 (N_10150,N_9000,N_9815);
or U10151 (N_10151,N_9940,N_9579);
or U10152 (N_10152,N_9508,N_9735);
and U10153 (N_10153,N_9238,N_9603);
xnor U10154 (N_10154,N_9951,N_9838);
xnor U10155 (N_10155,N_9742,N_9457);
nor U10156 (N_10156,N_9322,N_9844);
nor U10157 (N_10157,N_9896,N_9326);
nand U10158 (N_10158,N_9895,N_9889);
and U10159 (N_10159,N_9999,N_9226);
or U10160 (N_10160,N_9106,N_9975);
nand U10161 (N_10161,N_9596,N_9455);
nor U10162 (N_10162,N_9900,N_9981);
and U10163 (N_10163,N_9850,N_9619);
nand U10164 (N_10164,N_9663,N_9099);
nor U10165 (N_10165,N_9331,N_9679);
nor U10166 (N_10166,N_9506,N_9272);
and U10167 (N_10167,N_9495,N_9294);
nand U10168 (N_10168,N_9672,N_9947);
or U10169 (N_10169,N_9050,N_9686);
xnor U10170 (N_10170,N_9020,N_9262);
xor U10171 (N_10171,N_9871,N_9659);
nor U10172 (N_10172,N_9601,N_9567);
and U10173 (N_10173,N_9261,N_9319);
nor U10174 (N_10174,N_9644,N_9503);
xnor U10175 (N_10175,N_9017,N_9372);
xnor U10176 (N_10176,N_9898,N_9283);
and U10177 (N_10177,N_9950,N_9058);
nor U10178 (N_10178,N_9690,N_9033);
nor U10179 (N_10179,N_9756,N_9408);
or U10180 (N_10180,N_9544,N_9832);
xnor U10181 (N_10181,N_9490,N_9184);
and U10182 (N_10182,N_9246,N_9194);
nand U10183 (N_10183,N_9615,N_9195);
nor U10184 (N_10184,N_9138,N_9709);
xor U10185 (N_10185,N_9923,N_9586);
nand U10186 (N_10186,N_9587,N_9778);
nand U10187 (N_10187,N_9192,N_9153);
nand U10188 (N_10188,N_9862,N_9096);
nand U10189 (N_10189,N_9650,N_9103);
nor U10190 (N_10190,N_9150,N_9573);
nor U10191 (N_10191,N_9717,N_9980);
or U10192 (N_10192,N_9944,N_9307);
nor U10193 (N_10193,N_9253,N_9683);
xor U10194 (N_10194,N_9074,N_9651);
xor U10195 (N_10195,N_9378,N_9394);
or U10196 (N_10196,N_9178,N_9130);
and U10197 (N_10197,N_9055,N_9303);
xor U10198 (N_10198,N_9321,N_9565);
and U10199 (N_10199,N_9767,N_9910);
xor U10200 (N_10200,N_9633,N_9129);
and U10201 (N_10201,N_9645,N_9915);
or U10202 (N_10202,N_9496,N_9398);
nor U10203 (N_10203,N_9801,N_9202);
and U10204 (N_10204,N_9170,N_9966);
nand U10205 (N_10205,N_9205,N_9117);
nand U10206 (N_10206,N_9329,N_9908);
nand U10207 (N_10207,N_9373,N_9080);
xor U10208 (N_10208,N_9411,N_9423);
or U10209 (N_10209,N_9093,N_9057);
xor U10210 (N_10210,N_9221,N_9332);
xnor U10211 (N_10211,N_9762,N_9920);
nor U10212 (N_10212,N_9545,N_9812);
xnor U10213 (N_10213,N_9948,N_9061);
nor U10214 (N_10214,N_9460,N_9207);
xor U10215 (N_10215,N_9426,N_9462);
xnor U10216 (N_10216,N_9761,N_9247);
nor U10217 (N_10217,N_9652,N_9273);
nand U10218 (N_10218,N_9885,N_9218);
nor U10219 (N_10219,N_9208,N_9932);
xor U10220 (N_10220,N_9375,N_9682);
nand U10221 (N_10221,N_9806,N_9711);
xor U10222 (N_10222,N_9817,N_9894);
nor U10223 (N_10223,N_9819,N_9786);
or U10224 (N_10224,N_9432,N_9509);
nand U10225 (N_10225,N_9785,N_9234);
nand U10226 (N_10226,N_9530,N_9604);
xor U10227 (N_10227,N_9859,N_9989);
nand U10228 (N_10228,N_9356,N_9448);
and U10229 (N_10229,N_9733,N_9901);
xnor U10230 (N_10230,N_9597,N_9039);
or U10231 (N_10231,N_9800,N_9387);
nand U10232 (N_10232,N_9748,N_9009);
xor U10233 (N_10233,N_9831,N_9114);
nor U10234 (N_10234,N_9144,N_9660);
xor U10235 (N_10235,N_9346,N_9298);
or U10236 (N_10236,N_9744,N_9630);
or U10237 (N_10237,N_9790,N_9349);
nand U10238 (N_10238,N_9974,N_9593);
or U10239 (N_10239,N_9834,N_9616);
nor U10240 (N_10240,N_9088,N_9474);
or U10241 (N_10241,N_9044,N_9511);
and U10242 (N_10242,N_9998,N_9699);
xnor U10243 (N_10243,N_9222,N_9478);
xor U10244 (N_10244,N_9374,N_9124);
or U10245 (N_10245,N_9654,N_9560);
nand U10246 (N_10246,N_9890,N_9609);
or U10247 (N_10247,N_9960,N_9168);
nand U10248 (N_10248,N_9809,N_9858);
or U10249 (N_10249,N_9632,N_9878);
and U10250 (N_10250,N_9482,N_9688);
or U10251 (N_10251,N_9229,N_9019);
or U10252 (N_10252,N_9500,N_9032);
xor U10253 (N_10253,N_9095,N_9720);
and U10254 (N_10254,N_9501,N_9488);
xor U10255 (N_10255,N_9422,N_9611);
nand U10256 (N_10256,N_9104,N_9086);
or U10257 (N_10257,N_9388,N_9162);
xnor U10258 (N_10258,N_9256,N_9664);
nor U10259 (N_10259,N_9774,N_9166);
nand U10260 (N_10260,N_9823,N_9822);
nand U10261 (N_10261,N_9056,N_9588);
or U10262 (N_10262,N_9769,N_9958);
nor U10263 (N_10263,N_9670,N_9963);
nor U10264 (N_10264,N_9368,N_9421);
nand U10265 (N_10265,N_9415,N_9014);
nor U10266 (N_10266,N_9066,N_9305);
and U10267 (N_10267,N_9429,N_9292);
and U10268 (N_10268,N_9768,N_9594);
nand U10269 (N_10269,N_9606,N_9922);
nand U10270 (N_10270,N_9771,N_9128);
nand U10271 (N_10271,N_9855,N_9233);
nor U10272 (N_10272,N_9425,N_9220);
or U10273 (N_10273,N_9013,N_9147);
xor U10274 (N_10274,N_9323,N_9668);
nand U10275 (N_10275,N_9494,N_9288);
nor U10276 (N_10276,N_9726,N_9673);
xor U10277 (N_10277,N_9979,N_9524);
nor U10278 (N_10278,N_9236,N_9141);
xor U10279 (N_10279,N_9721,N_9863);
xor U10280 (N_10280,N_9163,N_9209);
or U10281 (N_10281,N_9384,N_9489);
nand U10282 (N_10282,N_9872,N_9318);
nand U10283 (N_10283,N_9563,N_9021);
or U10284 (N_10284,N_9595,N_9053);
nand U10285 (N_10285,N_9987,N_9765);
xnor U10286 (N_10286,N_9880,N_9638);
and U10287 (N_10287,N_9684,N_9502);
nor U10288 (N_10288,N_9393,N_9468);
or U10289 (N_10289,N_9333,N_9235);
or U10290 (N_10290,N_9325,N_9228);
xor U10291 (N_10291,N_9916,N_9612);
xor U10292 (N_10292,N_9734,N_9098);
or U10293 (N_10293,N_9389,N_9941);
xnor U10294 (N_10294,N_9969,N_9030);
or U10295 (N_10295,N_9991,N_9773);
or U10296 (N_10296,N_9681,N_9090);
nand U10297 (N_10297,N_9517,N_9004);
nand U10298 (N_10298,N_9034,N_9886);
xor U10299 (N_10299,N_9068,N_9725);
nor U10300 (N_10300,N_9291,N_9165);
xor U10301 (N_10301,N_9533,N_9309);
and U10302 (N_10302,N_9404,N_9437);
nor U10303 (N_10303,N_9557,N_9868);
xor U10304 (N_10304,N_9542,N_9018);
nand U10305 (N_10305,N_9347,N_9708);
or U10306 (N_10306,N_9454,N_9821);
nand U10307 (N_10307,N_9779,N_9535);
nand U10308 (N_10308,N_9719,N_9661);
nand U10309 (N_10309,N_9804,N_9264);
or U10310 (N_10310,N_9434,N_9203);
nand U10311 (N_10311,N_9038,N_9965);
or U10312 (N_10312,N_9610,N_9957);
nor U10313 (N_10313,N_9337,N_9707);
nor U10314 (N_10314,N_9145,N_9391);
xor U10315 (N_10315,N_9297,N_9176);
or U10316 (N_10316,N_9110,N_9856);
or U10317 (N_10317,N_9555,N_9655);
nand U10318 (N_10318,N_9132,N_9348);
or U10319 (N_10319,N_9417,N_9480);
nand U10320 (N_10320,N_9204,N_9101);
nor U10321 (N_10321,N_9364,N_9929);
xnor U10322 (N_10322,N_9798,N_9097);
nor U10323 (N_10323,N_9271,N_9476);
xnor U10324 (N_10324,N_9244,N_9327);
and U10325 (N_10325,N_9414,N_9705);
nand U10326 (N_10326,N_9175,N_9148);
nand U10327 (N_10327,N_9746,N_9289);
nor U10328 (N_10328,N_9465,N_9840);
and U10329 (N_10329,N_9477,N_9935);
xnor U10330 (N_10330,N_9354,N_9420);
and U10331 (N_10331,N_9463,N_9534);
nor U10332 (N_10332,N_9475,N_9108);
or U10333 (N_10333,N_9022,N_9945);
and U10334 (N_10334,N_9441,N_9631);
and U10335 (N_10335,N_9881,N_9301);
and U10336 (N_10336,N_9100,N_9589);
and U10337 (N_10337,N_9667,N_9286);
xnor U10338 (N_10338,N_9453,N_9634);
and U10339 (N_10339,N_9031,N_9279);
nand U10340 (N_10340,N_9122,N_9189);
nand U10341 (N_10341,N_9899,N_9193);
nor U10342 (N_10342,N_9052,N_9829);
and U10343 (N_10343,N_9956,N_9115);
nor U10344 (N_10344,N_9706,N_9814);
nor U10345 (N_10345,N_9628,N_9284);
and U10346 (N_10346,N_9777,N_9407);
or U10347 (N_10347,N_9358,N_9275);
xnor U10348 (N_10348,N_9642,N_9973);
nor U10349 (N_10349,N_9390,N_9728);
nor U10350 (N_10350,N_9252,N_9161);
xor U10351 (N_10351,N_9732,N_9729);
nand U10352 (N_10352,N_9914,N_9599);
or U10353 (N_10353,N_9497,N_9164);
and U10354 (N_10354,N_9870,N_9581);
or U10355 (N_10355,N_9483,N_9173);
and U10356 (N_10356,N_9759,N_9199);
nor U10357 (N_10357,N_9913,N_9942);
nor U10358 (N_10358,N_9625,N_9036);
nor U10359 (N_10359,N_9825,N_9491);
and U10360 (N_10360,N_9854,N_9763);
nor U10361 (N_10361,N_9191,N_9933);
and U10362 (N_10362,N_9450,N_9715);
or U10363 (N_10363,N_9396,N_9359);
and U10364 (N_10364,N_9188,N_9580);
nand U10365 (N_10365,N_9847,N_9722);
and U10366 (N_10366,N_9342,N_9649);
xor U10367 (N_10367,N_9793,N_9485);
nor U10368 (N_10368,N_9584,N_9737);
or U10369 (N_10369,N_9245,N_9521);
or U10370 (N_10370,N_9452,N_9269);
and U10371 (N_10371,N_9754,N_9865);
nor U10372 (N_10372,N_9341,N_9925);
and U10373 (N_10373,N_9702,N_9338);
nor U10374 (N_10374,N_9406,N_9005);
or U10375 (N_10375,N_9312,N_9879);
xor U10376 (N_10376,N_9127,N_9472);
nand U10377 (N_10377,N_9627,N_9539);
and U10378 (N_10378,N_9187,N_9888);
and U10379 (N_10379,N_9126,N_9904);
xor U10380 (N_10380,N_9564,N_9694);
nand U10381 (N_10381,N_9084,N_9424);
xor U10382 (N_10382,N_9678,N_9514);
or U10383 (N_10383,N_9696,N_9561);
and U10384 (N_10384,N_9371,N_9160);
nor U10385 (N_10385,N_9532,N_9087);
nor U10386 (N_10386,N_9802,N_9109);
and U10387 (N_10387,N_9978,N_9026);
and U10388 (N_10388,N_9745,N_9201);
or U10389 (N_10389,N_9042,N_9845);
xnor U10390 (N_10390,N_9639,N_9938);
nand U10391 (N_10391,N_9697,N_9666);
xnor U10392 (N_10392,N_9366,N_9412);
and U10393 (N_10393,N_9740,N_9553);
nand U10394 (N_10394,N_9180,N_9152);
nor U10395 (N_10395,N_9459,N_9547);
and U10396 (N_10396,N_9369,N_9671);
xnor U10397 (N_10397,N_9964,N_9608);
nor U10398 (N_10398,N_9003,N_9379);
or U10399 (N_10399,N_9805,N_9427);
or U10400 (N_10400,N_9770,N_9917);
nand U10401 (N_10401,N_9523,N_9752);
xnor U10402 (N_10402,N_9522,N_9936);
nand U10403 (N_10403,N_9011,N_9433);
nor U10404 (N_10404,N_9092,N_9473);
and U10405 (N_10405,N_9536,N_9716);
and U10406 (N_10406,N_9315,N_9381);
nor U10407 (N_10407,N_9449,N_9570);
and U10408 (N_10408,N_9693,N_9302);
nand U10409 (N_10409,N_9155,N_9446);
nor U10410 (N_10410,N_9883,N_9566);
xnor U10411 (N_10411,N_9623,N_9197);
or U10412 (N_10412,N_9112,N_9392);
nor U10413 (N_10413,N_9955,N_9456);
nor U10414 (N_10414,N_9308,N_9874);
and U10415 (N_10415,N_9794,N_9828);
nor U10416 (N_10416,N_9266,N_9043);
nand U10417 (N_10417,N_9598,N_9313);
nand U10418 (N_10418,N_9549,N_9877);
and U10419 (N_10419,N_9278,N_9257);
nand U10420 (N_10420,N_9689,N_9079);
nand U10421 (N_10421,N_9591,N_9724);
nand U10422 (N_10422,N_9028,N_9605);
nor U10423 (N_10423,N_9931,N_9306);
nand U10424 (N_10424,N_9461,N_9077);
or U10425 (N_10425,N_9219,N_9265);
and U10426 (N_10426,N_9640,N_9395);
or U10427 (N_10427,N_9996,N_9402);
or U10428 (N_10428,N_9710,N_9451);
nor U10429 (N_10429,N_9695,N_9712);
nor U10430 (N_10430,N_9023,N_9992);
and U10431 (N_10431,N_9558,N_9361);
and U10432 (N_10432,N_9993,N_9046);
nand U10433 (N_10433,N_9946,N_9486);
or U10434 (N_10434,N_9853,N_9006);
xor U10435 (N_10435,N_9578,N_9852);
and U10436 (N_10436,N_9851,N_9344);
nand U10437 (N_10437,N_9961,N_9282);
or U10438 (N_10438,N_9538,N_9692);
and U10439 (N_10439,N_9200,N_9300);
or U10440 (N_10440,N_9626,N_9571);
nand U10441 (N_10441,N_9365,N_9939);
xnor U10442 (N_10442,N_9362,N_9409);
and U10443 (N_10443,N_9239,N_9531);
nand U10444 (N_10444,N_9513,N_9120);
xor U10445 (N_10445,N_9789,N_9867);
or U10446 (N_10446,N_9820,N_9146);
nand U10447 (N_10447,N_9988,N_9214);
nor U10448 (N_10448,N_9249,N_9250);
nand U10449 (N_10449,N_9738,N_9876);
nor U10450 (N_10450,N_9102,N_9001);
nand U10451 (N_10451,N_9063,N_9242);
nand U10452 (N_10452,N_9317,N_9713);
xor U10453 (N_10453,N_9091,N_9386);
xnor U10454 (N_10454,N_9577,N_9060);
or U10455 (N_10455,N_9792,N_9377);
nand U10456 (N_10456,N_9569,N_9435);
nor U10457 (N_10457,N_9487,N_9585);
nand U10458 (N_10458,N_9440,N_9691);
nand U10459 (N_10459,N_9047,N_9400);
nor U10460 (N_10460,N_9304,N_9643);
or U10461 (N_10461,N_9498,N_9839);
nand U10462 (N_10462,N_9857,N_9930);
and U10463 (N_10463,N_9159,N_9210);
or U10464 (N_10464,N_9512,N_9428);
or U10465 (N_10465,N_9747,N_9268);
and U10466 (N_10466,N_9137,N_9183);
or U10467 (N_10467,N_9912,N_9897);
or U10468 (N_10468,N_9653,N_9016);
xor U10469 (N_10469,N_9525,N_9143);
xnor U10470 (N_10470,N_9430,N_9336);
xnor U10471 (N_10471,N_9519,N_9287);
xor U10472 (N_10472,N_9263,N_9764);
or U10473 (N_10473,N_9559,N_9083);
nor U10474 (N_10474,N_9334,N_9340);
xnor U10475 (N_10475,N_9962,N_9133);
nand U10476 (N_10476,N_9954,N_9637);
nor U10477 (N_10477,N_9700,N_9685);
nor U10478 (N_10478,N_9382,N_9953);
and U10479 (N_10479,N_9884,N_9010);
or U10480 (N_10480,N_9620,N_9123);
nor U10481 (N_10481,N_9576,N_9215);
xnor U10482 (N_10482,N_9403,N_9552);
nor U10483 (N_10483,N_9206,N_9550);
nor U10484 (N_10484,N_9380,N_9582);
nor U10485 (N_10485,N_9405,N_9590);
or U10486 (N_10486,N_9808,N_9230);
and U10487 (N_10487,N_9842,N_9750);
nand U10488 (N_10488,N_9727,N_9352);
or U10489 (N_10489,N_9718,N_9860);
and U10490 (N_10490,N_9360,N_9280);
nand U10491 (N_10491,N_9169,N_9600);
xnor U10492 (N_10492,N_9357,N_9891);
and U10493 (N_10493,N_9968,N_9383);
xnor U10494 (N_10494,N_9223,N_9350);
and U10495 (N_10495,N_9617,N_9799);
xor U10496 (N_10496,N_9174,N_9629);
and U10497 (N_10497,N_9648,N_9035);
nand U10498 (N_10498,N_9826,N_9012);
nand U10499 (N_10499,N_9926,N_9985);
or U10500 (N_10500,N_9846,N_9387);
nand U10501 (N_10501,N_9999,N_9576);
nor U10502 (N_10502,N_9298,N_9826);
xnor U10503 (N_10503,N_9859,N_9226);
nand U10504 (N_10504,N_9308,N_9899);
and U10505 (N_10505,N_9736,N_9061);
and U10506 (N_10506,N_9566,N_9643);
nor U10507 (N_10507,N_9555,N_9108);
and U10508 (N_10508,N_9600,N_9597);
and U10509 (N_10509,N_9187,N_9770);
or U10510 (N_10510,N_9181,N_9696);
and U10511 (N_10511,N_9959,N_9134);
and U10512 (N_10512,N_9360,N_9240);
or U10513 (N_10513,N_9582,N_9012);
nand U10514 (N_10514,N_9843,N_9970);
or U10515 (N_10515,N_9318,N_9111);
nor U10516 (N_10516,N_9856,N_9080);
nand U10517 (N_10517,N_9120,N_9471);
nor U10518 (N_10518,N_9767,N_9319);
and U10519 (N_10519,N_9975,N_9808);
and U10520 (N_10520,N_9671,N_9335);
xnor U10521 (N_10521,N_9392,N_9440);
nand U10522 (N_10522,N_9968,N_9036);
xnor U10523 (N_10523,N_9775,N_9243);
nand U10524 (N_10524,N_9535,N_9391);
xnor U10525 (N_10525,N_9838,N_9602);
nor U10526 (N_10526,N_9395,N_9515);
nand U10527 (N_10527,N_9962,N_9155);
xnor U10528 (N_10528,N_9645,N_9573);
nand U10529 (N_10529,N_9360,N_9982);
nor U10530 (N_10530,N_9562,N_9433);
xnor U10531 (N_10531,N_9383,N_9536);
and U10532 (N_10532,N_9827,N_9031);
nor U10533 (N_10533,N_9800,N_9132);
and U10534 (N_10534,N_9469,N_9919);
nand U10535 (N_10535,N_9746,N_9941);
and U10536 (N_10536,N_9552,N_9316);
nor U10537 (N_10537,N_9912,N_9575);
nor U10538 (N_10538,N_9342,N_9326);
and U10539 (N_10539,N_9824,N_9074);
nor U10540 (N_10540,N_9057,N_9800);
and U10541 (N_10541,N_9475,N_9546);
xnor U10542 (N_10542,N_9393,N_9591);
nor U10543 (N_10543,N_9677,N_9353);
nand U10544 (N_10544,N_9182,N_9034);
or U10545 (N_10545,N_9620,N_9451);
nor U10546 (N_10546,N_9856,N_9712);
nor U10547 (N_10547,N_9827,N_9829);
xor U10548 (N_10548,N_9033,N_9694);
nand U10549 (N_10549,N_9238,N_9034);
or U10550 (N_10550,N_9797,N_9582);
nand U10551 (N_10551,N_9171,N_9488);
xor U10552 (N_10552,N_9593,N_9415);
xnor U10553 (N_10553,N_9162,N_9934);
and U10554 (N_10554,N_9794,N_9322);
nor U10555 (N_10555,N_9514,N_9453);
or U10556 (N_10556,N_9416,N_9822);
and U10557 (N_10557,N_9842,N_9159);
and U10558 (N_10558,N_9514,N_9827);
nand U10559 (N_10559,N_9925,N_9982);
nand U10560 (N_10560,N_9743,N_9155);
xnor U10561 (N_10561,N_9458,N_9485);
xnor U10562 (N_10562,N_9552,N_9540);
or U10563 (N_10563,N_9964,N_9966);
nand U10564 (N_10564,N_9797,N_9618);
nand U10565 (N_10565,N_9276,N_9818);
nor U10566 (N_10566,N_9911,N_9778);
xor U10567 (N_10567,N_9328,N_9613);
xor U10568 (N_10568,N_9416,N_9385);
or U10569 (N_10569,N_9573,N_9043);
and U10570 (N_10570,N_9705,N_9949);
or U10571 (N_10571,N_9594,N_9238);
xor U10572 (N_10572,N_9812,N_9909);
nand U10573 (N_10573,N_9355,N_9924);
and U10574 (N_10574,N_9481,N_9678);
nor U10575 (N_10575,N_9823,N_9047);
or U10576 (N_10576,N_9129,N_9813);
or U10577 (N_10577,N_9811,N_9905);
nor U10578 (N_10578,N_9161,N_9701);
or U10579 (N_10579,N_9696,N_9253);
and U10580 (N_10580,N_9321,N_9867);
nand U10581 (N_10581,N_9721,N_9288);
nor U10582 (N_10582,N_9124,N_9426);
and U10583 (N_10583,N_9736,N_9381);
and U10584 (N_10584,N_9977,N_9565);
and U10585 (N_10585,N_9507,N_9829);
and U10586 (N_10586,N_9665,N_9653);
nand U10587 (N_10587,N_9327,N_9739);
xnor U10588 (N_10588,N_9875,N_9256);
or U10589 (N_10589,N_9739,N_9177);
and U10590 (N_10590,N_9006,N_9862);
xor U10591 (N_10591,N_9043,N_9346);
nand U10592 (N_10592,N_9396,N_9469);
and U10593 (N_10593,N_9361,N_9963);
or U10594 (N_10594,N_9409,N_9561);
xor U10595 (N_10595,N_9259,N_9881);
nand U10596 (N_10596,N_9027,N_9207);
or U10597 (N_10597,N_9682,N_9387);
and U10598 (N_10598,N_9667,N_9482);
xor U10599 (N_10599,N_9086,N_9636);
xnor U10600 (N_10600,N_9982,N_9823);
and U10601 (N_10601,N_9448,N_9671);
and U10602 (N_10602,N_9182,N_9571);
xnor U10603 (N_10603,N_9866,N_9273);
nor U10604 (N_10604,N_9518,N_9681);
nor U10605 (N_10605,N_9670,N_9686);
nor U10606 (N_10606,N_9174,N_9245);
nor U10607 (N_10607,N_9864,N_9295);
nor U10608 (N_10608,N_9919,N_9640);
and U10609 (N_10609,N_9264,N_9909);
or U10610 (N_10610,N_9728,N_9065);
xor U10611 (N_10611,N_9059,N_9520);
xor U10612 (N_10612,N_9270,N_9875);
or U10613 (N_10613,N_9758,N_9155);
xnor U10614 (N_10614,N_9378,N_9153);
or U10615 (N_10615,N_9697,N_9660);
xnor U10616 (N_10616,N_9300,N_9174);
nand U10617 (N_10617,N_9213,N_9215);
xor U10618 (N_10618,N_9480,N_9753);
or U10619 (N_10619,N_9159,N_9419);
xor U10620 (N_10620,N_9590,N_9431);
xnor U10621 (N_10621,N_9911,N_9933);
xnor U10622 (N_10622,N_9728,N_9290);
nand U10623 (N_10623,N_9926,N_9822);
xor U10624 (N_10624,N_9072,N_9238);
nor U10625 (N_10625,N_9812,N_9378);
nand U10626 (N_10626,N_9218,N_9557);
xor U10627 (N_10627,N_9196,N_9341);
xnor U10628 (N_10628,N_9178,N_9664);
or U10629 (N_10629,N_9877,N_9545);
and U10630 (N_10630,N_9206,N_9766);
and U10631 (N_10631,N_9814,N_9624);
nand U10632 (N_10632,N_9842,N_9281);
xnor U10633 (N_10633,N_9059,N_9863);
nand U10634 (N_10634,N_9604,N_9945);
and U10635 (N_10635,N_9530,N_9348);
nor U10636 (N_10636,N_9385,N_9971);
nand U10637 (N_10637,N_9180,N_9794);
and U10638 (N_10638,N_9444,N_9133);
nor U10639 (N_10639,N_9038,N_9031);
and U10640 (N_10640,N_9834,N_9500);
and U10641 (N_10641,N_9881,N_9655);
nand U10642 (N_10642,N_9802,N_9148);
nand U10643 (N_10643,N_9520,N_9769);
xor U10644 (N_10644,N_9809,N_9612);
or U10645 (N_10645,N_9265,N_9704);
nand U10646 (N_10646,N_9287,N_9227);
nand U10647 (N_10647,N_9743,N_9947);
xnor U10648 (N_10648,N_9411,N_9942);
xnor U10649 (N_10649,N_9652,N_9849);
nand U10650 (N_10650,N_9586,N_9452);
xnor U10651 (N_10651,N_9620,N_9948);
nand U10652 (N_10652,N_9487,N_9513);
nor U10653 (N_10653,N_9239,N_9830);
or U10654 (N_10654,N_9854,N_9277);
xor U10655 (N_10655,N_9808,N_9357);
or U10656 (N_10656,N_9551,N_9768);
and U10657 (N_10657,N_9878,N_9019);
or U10658 (N_10658,N_9926,N_9537);
or U10659 (N_10659,N_9394,N_9899);
nor U10660 (N_10660,N_9205,N_9320);
or U10661 (N_10661,N_9523,N_9721);
and U10662 (N_10662,N_9096,N_9082);
nor U10663 (N_10663,N_9421,N_9492);
or U10664 (N_10664,N_9973,N_9121);
nand U10665 (N_10665,N_9008,N_9822);
nand U10666 (N_10666,N_9878,N_9664);
xor U10667 (N_10667,N_9679,N_9034);
nand U10668 (N_10668,N_9596,N_9910);
xnor U10669 (N_10669,N_9645,N_9095);
and U10670 (N_10670,N_9347,N_9345);
and U10671 (N_10671,N_9409,N_9137);
and U10672 (N_10672,N_9711,N_9957);
nand U10673 (N_10673,N_9127,N_9073);
or U10674 (N_10674,N_9403,N_9130);
or U10675 (N_10675,N_9720,N_9743);
xnor U10676 (N_10676,N_9810,N_9502);
and U10677 (N_10677,N_9952,N_9598);
nand U10678 (N_10678,N_9846,N_9356);
nor U10679 (N_10679,N_9301,N_9610);
nor U10680 (N_10680,N_9050,N_9508);
and U10681 (N_10681,N_9563,N_9856);
and U10682 (N_10682,N_9425,N_9884);
xnor U10683 (N_10683,N_9785,N_9676);
xnor U10684 (N_10684,N_9927,N_9121);
or U10685 (N_10685,N_9252,N_9756);
nand U10686 (N_10686,N_9224,N_9087);
or U10687 (N_10687,N_9067,N_9687);
nor U10688 (N_10688,N_9246,N_9271);
and U10689 (N_10689,N_9017,N_9613);
and U10690 (N_10690,N_9085,N_9129);
or U10691 (N_10691,N_9037,N_9772);
nand U10692 (N_10692,N_9951,N_9177);
nand U10693 (N_10693,N_9417,N_9796);
nand U10694 (N_10694,N_9121,N_9939);
nand U10695 (N_10695,N_9751,N_9851);
xnor U10696 (N_10696,N_9310,N_9094);
nor U10697 (N_10697,N_9092,N_9594);
nor U10698 (N_10698,N_9798,N_9515);
nor U10699 (N_10699,N_9674,N_9248);
xnor U10700 (N_10700,N_9341,N_9565);
xnor U10701 (N_10701,N_9355,N_9913);
or U10702 (N_10702,N_9378,N_9237);
and U10703 (N_10703,N_9101,N_9967);
nor U10704 (N_10704,N_9209,N_9706);
nor U10705 (N_10705,N_9029,N_9673);
xor U10706 (N_10706,N_9763,N_9607);
nand U10707 (N_10707,N_9291,N_9933);
nand U10708 (N_10708,N_9480,N_9588);
nand U10709 (N_10709,N_9533,N_9728);
or U10710 (N_10710,N_9669,N_9460);
and U10711 (N_10711,N_9949,N_9819);
or U10712 (N_10712,N_9287,N_9056);
xor U10713 (N_10713,N_9996,N_9409);
nor U10714 (N_10714,N_9712,N_9177);
nor U10715 (N_10715,N_9828,N_9713);
nor U10716 (N_10716,N_9518,N_9435);
or U10717 (N_10717,N_9835,N_9181);
nand U10718 (N_10718,N_9612,N_9248);
nor U10719 (N_10719,N_9816,N_9843);
nor U10720 (N_10720,N_9972,N_9508);
nor U10721 (N_10721,N_9514,N_9273);
nor U10722 (N_10722,N_9171,N_9281);
nor U10723 (N_10723,N_9892,N_9838);
nor U10724 (N_10724,N_9128,N_9239);
nand U10725 (N_10725,N_9996,N_9891);
xor U10726 (N_10726,N_9444,N_9236);
nand U10727 (N_10727,N_9486,N_9756);
xnor U10728 (N_10728,N_9263,N_9186);
nand U10729 (N_10729,N_9303,N_9940);
nor U10730 (N_10730,N_9717,N_9668);
nor U10731 (N_10731,N_9349,N_9008);
and U10732 (N_10732,N_9834,N_9488);
xnor U10733 (N_10733,N_9273,N_9192);
xor U10734 (N_10734,N_9302,N_9442);
or U10735 (N_10735,N_9671,N_9911);
nor U10736 (N_10736,N_9079,N_9833);
or U10737 (N_10737,N_9025,N_9337);
and U10738 (N_10738,N_9479,N_9454);
or U10739 (N_10739,N_9616,N_9245);
or U10740 (N_10740,N_9251,N_9369);
or U10741 (N_10741,N_9125,N_9657);
or U10742 (N_10742,N_9726,N_9417);
xnor U10743 (N_10743,N_9107,N_9308);
and U10744 (N_10744,N_9773,N_9579);
and U10745 (N_10745,N_9416,N_9529);
nand U10746 (N_10746,N_9640,N_9898);
xor U10747 (N_10747,N_9227,N_9613);
and U10748 (N_10748,N_9489,N_9417);
nor U10749 (N_10749,N_9917,N_9007);
xnor U10750 (N_10750,N_9595,N_9681);
or U10751 (N_10751,N_9996,N_9340);
or U10752 (N_10752,N_9831,N_9187);
or U10753 (N_10753,N_9157,N_9372);
xor U10754 (N_10754,N_9714,N_9711);
and U10755 (N_10755,N_9060,N_9094);
or U10756 (N_10756,N_9431,N_9374);
and U10757 (N_10757,N_9356,N_9609);
nand U10758 (N_10758,N_9604,N_9458);
xnor U10759 (N_10759,N_9684,N_9055);
nand U10760 (N_10760,N_9193,N_9090);
nor U10761 (N_10761,N_9223,N_9200);
nor U10762 (N_10762,N_9292,N_9892);
nor U10763 (N_10763,N_9528,N_9239);
xor U10764 (N_10764,N_9842,N_9861);
and U10765 (N_10765,N_9191,N_9921);
nand U10766 (N_10766,N_9203,N_9145);
and U10767 (N_10767,N_9563,N_9090);
or U10768 (N_10768,N_9855,N_9364);
and U10769 (N_10769,N_9872,N_9548);
nor U10770 (N_10770,N_9291,N_9195);
nor U10771 (N_10771,N_9265,N_9853);
xnor U10772 (N_10772,N_9863,N_9793);
and U10773 (N_10773,N_9730,N_9502);
or U10774 (N_10774,N_9446,N_9652);
nor U10775 (N_10775,N_9023,N_9529);
nor U10776 (N_10776,N_9981,N_9495);
and U10777 (N_10777,N_9920,N_9600);
and U10778 (N_10778,N_9292,N_9559);
or U10779 (N_10779,N_9584,N_9799);
nand U10780 (N_10780,N_9541,N_9267);
xor U10781 (N_10781,N_9906,N_9263);
nand U10782 (N_10782,N_9458,N_9957);
or U10783 (N_10783,N_9039,N_9657);
xor U10784 (N_10784,N_9982,N_9313);
nor U10785 (N_10785,N_9784,N_9191);
nand U10786 (N_10786,N_9740,N_9826);
or U10787 (N_10787,N_9244,N_9537);
and U10788 (N_10788,N_9117,N_9718);
nand U10789 (N_10789,N_9853,N_9460);
or U10790 (N_10790,N_9765,N_9603);
and U10791 (N_10791,N_9821,N_9606);
nor U10792 (N_10792,N_9583,N_9323);
nand U10793 (N_10793,N_9822,N_9854);
or U10794 (N_10794,N_9840,N_9246);
nand U10795 (N_10795,N_9477,N_9322);
nor U10796 (N_10796,N_9258,N_9844);
and U10797 (N_10797,N_9388,N_9486);
nor U10798 (N_10798,N_9699,N_9854);
and U10799 (N_10799,N_9103,N_9811);
nand U10800 (N_10800,N_9713,N_9734);
or U10801 (N_10801,N_9857,N_9964);
or U10802 (N_10802,N_9678,N_9781);
and U10803 (N_10803,N_9624,N_9506);
xor U10804 (N_10804,N_9857,N_9694);
and U10805 (N_10805,N_9040,N_9025);
xor U10806 (N_10806,N_9395,N_9884);
or U10807 (N_10807,N_9373,N_9169);
xnor U10808 (N_10808,N_9012,N_9698);
nand U10809 (N_10809,N_9472,N_9389);
or U10810 (N_10810,N_9344,N_9321);
nand U10811 (N_10811,N_9812,N_9213);
xor U10812 (N_10812,N_9662,N_9788);
nor U10813 (N_10813,N_9514,N_9620);
and U10814 (N_10814,N_9914,N_9515);
or U10815 (N_10815,N_9339,N_9470);
nor U10816 (N_10816,N_9453,N_9861);
nand U10817 (N_10817,N_9266,N_9740);
nor U10818 (N_10818,N_9010,N_9554);
nand U10819 (N_10819,N_9325,N_9639);
or U10820 (N_10820,N_9729,N_9219);
nor U10821 (N_10821,N_9513,N_9231);
and U10822 (N_10822,N_9074,N_9414);
and U10823 (N_10823,N_9909,N_9353);
nor U10824 (N_10824,N_9762,N_9411);
nand U10825 (N_10825,N_9552,N_9785);
nor U10826 (N_10826,N_9972,N_9913);
and U10827 (N_10827,N_9975,N_9976);
xor U10828 (N_10828,N_9233,N_9154);
or U10829 (N_10829,N_9992,N_9801);
nand U10830 (N_10830,N_9753,N_9882);
nand U10831 (N_10831,N_9026,N_9084);
xor U10832 (N_10832,N_9459,N_9957);
or U10833 (N_10833,N_9850,N_9736);
nand U10834 (N_10834,N_9582,N_9327);
xor U10835 (N_10835,N_9118,N_9242);
and U10836 (N_10836,N_9838,N_9656);
nand U10837 (N_10837,N_9926,N_9883);
nor U10838 (N_10838,N_9926,N_9820);
xnor U10839 (N_10839,N_9519,N_9195);
xor U10840 (N_10840,N_9122,N_9391);
and U10841 (N_10841,N_9108,N_9990);
nor U10842 (N_10842,N_9939,N_9512);
and U10843 (N_10843,N_9780,N_9101);
and U10844 (N_10844,N_9203,N_9437);
nand U10845 (N_10845,N_9527,N_9920);
or U10846 (N_10846,N_9979,N_9472);
and U10847 (N_10847,N_9657,N_9662);
xnor U10848 (N_10848,N_9050,N_9272);
nand U10849 (N_10849,N_9998,N_9068);
or U10850 (N_10850,N_9059,N_9352);
nand U10851 (N_10851,N_9886,N_9864);
nor U10852 (N_10852,N_9803,N_9216);
and U10853 (N_10853,N_9117,N_9258);
nor U10854 (N_10854,N_9982,N_9845);
and U10855 (N_10855,N_9583,N_9594);
nor U10856 (N_10856,N_9564,N_9437);
and U10857 (N_10857,N_9220,N_9369);
nor U10858 (N_10858,N_9876,N_9488);
nor U10859 (N_10859,N_9851,N_9208);
and U10860 (N_10860,N_9859,N_9719);
xnor U10861 (N_10861,N_9711,N_9888);
xor U10862 (N_10862,N_9935,N_9659);
xor U10863 (N_10863,N_9421,N_9789);
and U10864 (N_10864,N_9192,N_9115);
and U10865 (N_10865,N_9628,N_9873);
nor U10866 (N_10866,N_9483,N_9674);
or U10867 (N_10867,N_9294,N_9578);
nand U10868 (N_10868,N_9794,N_9942);
or U10869 (N_10869,N_9499,N_9351);
nor U10870 (N_10870,N_9447,N_9783);
nor U10871 (N_10871,N_9815,N_9795);
or U10872 (N_10872,N_9771,N_9304);
or U10873 (N_10873,N_9875,N_9624);
or U10874 (N_10874,N_9858,N_9121);
or U10875 (N_10875,N_9865,N_9201);
nand U10876 (N_10876,N_9707,N_9904);
nand U10877 (N_10877,N_9813,N_9544);
or U10878 (N_10878,N_9561,N_9640);
nand U10879 (N_10879,N_9531,N_9134);
nand U10880 (N_10880,N_9476,N_9419);
and U10881 (N_10881,N_9665,N_9250);
or U10882 (N_10882,N_9643,N_9469);
nand U10883 (N_10883,N_9246,N_9912);
and U10884 (N_10884,N_9339,N_9170);
and U10885 (N_10885,N_9066,N_9533);
nand U10886 (N_10886,N_9082,N_9118);
nor U10887 (N_10887,N_9528,N_9324);
nand U10888 (N_10888,N_9021,N_9873);
and U10889 (N_10889,N_9005,N_9418);
or U10890 (N_10890,N_9389,N_9682);
nor U10891 (N_10891,N_9254,N_9462);
nand U10892 (N_10892,N_9825,N_9175);
or U10893 (N_10893,N_9064,N_9386);
nand U10894 (N_10894,N_9102,N_9291);
nor U10895 (N_10895,N_9804,N_9408);
nor U10896 (N_10896,N_9048,N_9013);
nand U10897 (N_10897,N_9782,N_9893);
and U10898 (N_10898,N_9732,N_9439);
nor U10899 (N_10899,N_9002,N_9175);
nand U10900 (N_10900,N_9111,N_9070);
and U10901 (N_10901,N_9024,N_9257);
and U10902 (N_10902,N_9457,N_9694);
nor U10903 (N_10903,N_9271,N_9604);
xnor U10904 (N_10904,N_9021,N_9822);
or U10905 (N_10905,N_9567,N_9468);
xor U10906 (N_10906,N_9742,N_9893);
xor U10907 (N_10907,N_9186,N_9043);
xnor U10908 (N_10908,N_9906,N_9923);
xnor U10909 (N_10909,N_9800,N_9461);
nor U10910 (N_10910,N_9392,N_9506);
and U10911 (N_10911,N_9188,N_9419);
nor U10912 (N_10912,N_9032,N_9382);
or U10913 (N_10913,N_9680,N_9961);
or U10914 (N_10914,N_9779,N_9218);
or U10915 (N_10915,N_9668,N_9300);
nor U10916 (N_10916,N_9389,N_9046);
nor U10917 (N_10917,N_9060,N_9148);
and U10918 (N_10918,N_9030,N_9447);
and U10919 (N_10919,N_9511,N_9836);
nor U10920 (N_10920,N_9357,N_9655);
xnor U10921 (N_10921,N_9155,N_9376);
and U10922 (N_10922,N_9669,N_9133);
xor U10923 (N_10923,N_9665,N_9492);
nand U10924 (N_10924,N_9189,N_9933);
nand U10925 (N_10925,N_9451,N_9914);
nor U10926 (N_10926,N_9374,N_9372);
nor U10927 (N_10927,N_9255,N_9493);
or U10928 (N_10928,N_9292,N_9169);
nand U10929 (N_10929,N_9174,N_9981);
xnor U10930 (N_10930,N_9797,N_9872);
and U10931 (N_10931,N_9176,N_9825);
nor U10932 (N_10932,N_9860,N_9544);
and U10933 (N_10933,N_9121,N_9959);
nor U10934 (N_10934,N_9823,N_9311);
or U10935 (N_10935,N_9562,N_9684);
and U10936 (N_10936,N_9816,N_9997);
xor U10937 (N_10937,N_9684,N_9210);
and U10938 (N_10938,N_9636,N_9479);
xnor U10939 (N_10939,N_9447,N_9395);
or U10940 (N_10940,N_9252,N_9785);
or U10941 (N_10941,N_9030,N_9304);
and U10942 (N_10942,N_9868,N_9880);
or U10943 (N_10943,N_9633,N_9917);
nor U10944 (N_10944,N_9149,N_9819);
or U10945 (N_10945,N_9482,N_9395);
or U10946 (N_10946,N_9394,N_9205);
or U10947 (N_10947,N_9258,N_9001);
nor U10948 (N_10948,N_9119,N_9338);
or U10949 (N_10949,N_9023,N_9436);
nand U10950 (N_10950,N_9106,N_9631);
xor U10951 (N_10951,N_9662,N_9883);
nand U10952 (N_10952,N_9058,N_9737);
and U10953 (N_10953,N_9089,N_9581);
xor U10954 (N_10954,N_9570,N_9648);
and U10955 (N_10955,N_9695,N_9906);
nand U10956 (N_10956,N_9362,N_9084);
xor U10957 (N_10957,N_9962,N_9225);
xnor U10958 (N_10958,N_9970,N_9104);
or U10959 (N_10959,N_9948,N_9607);
or U10960 (N_10960,N_9765,N_9766);
xnor U10961 (N_10961,N_9378,N_9741);
nor U10962 (N_10962,N_9247,N_9108);
or U10963 (N_10963,N_9772,N_9004);
nor U10964 (N_10964,N_9582,N_9755);
xnor U10965 (N_10965,N_9736,N_9671);
xor U10966 (N_10966,N_9991,N_9475);
nor U10967 (N_10967,N_9241,N_9705);
and U10968 (N_10968,N_9665,N_9333);
nand U10969 (N_10969,N_9863,N_9351);
or U10970 (N_10970,N_9247,N_9599);
or U10971 (N_10971,N_9497,N_9262);
and U10972 (N_10972,N_9046,N_9803);
nor U10973 (N_10973,N_9786,N_9320);
and U10974 (N_10974,N_9610,N_9232);
xnor U10975 (N_10975,N_9383,N_9466);
xnor U10976 (N_10976,N_9462,N_9555);
nor U10977 (N_10977,N_9817,N_9046);
nand U10978 (N_10978,N_9494,N_9023);
nand U10979 (N_10979,N_9284,N_9025);
and U10980 (N_10980,N_9516,N_9642);
nor U10981 (N_10981,N_9500,N_9973);
nor U10982 (N_10982,N_9616,N_9922);
nand U10983 (N_10983,N_9587,N_9378);
xnor U10984 (N_10984,N_9511,N_9010);
nor U10985 (N_10985,N_9493,N_9366);
nor U10986 (N_10986,N_9032,N_9259);
and U10987 (N_10987,N_9218,N_9915);
xor U10988 (N_10988,N_9402,N_9243);
nor U10989 (N_10989,N_9677,N_9088);
nand U10990 (N_10990,N_9999,N_9671);
nor U10991 (N_10991,N_9366,N_9621);
nor U10992 (N_10992,N_9327,N_9942);
and U10993 (N_10993,N_9132,N_9668);
nand U10994 (N_10994,N_9241,N_9360);
nand U10995 (N_10995,N_9996,N_9742);
or U10996 (N_10996,N_9828,N_9279);
xor U10997 (N_10997,N_9210,N_9282);
and U10998 (N_10998,N_9354,N_9953);
or U10999 (N_10999,N_9843,N_9674);
and U11000 (N_11000,N_10057,N_10331);
nor U11001 (N_11001,N_10223,N_10807);
nand U11002 (N_11002,N_10943,N_10843);
and U11003 (N_11003,N_10966,N_10599);
xnor U11004 (N_11004,N_10798,N_10508);
or U11005 (N_11005,N_10381,N_10565);
xnor U11006 (N_11006,N_10694,N_10671);
or U11007 (N_11007,N_10292,N_10022);
nor U11008 (N_11008,N_10789,N_10075);
nand U11009 (N_11009,N_10492,N_10835);
nand U11010 (N_11010,N_10093,N_10400);
nor U11011 (N_11011,N_10338,N_10881);
xor U11012 (N_11012,N_10720,N_10315);
nand U11013 (N_11013,N_10870,N_10577);
nor U11014 (N_11014,N_10306,N_10275);
or U11015 (N_11015,N_10156,N_10008);
or U11016 (N_11016,N_10249,N_10396);
xor U11017 (N_11017,N_10619,N_10610);
or U11018 (N_11018,N_10510,N_10889);
and U11019 (N_11019,N_10735,N_10959);
nor U11020 (N_11020,N_10438,N_10218);
or U11021 (N_11021,N_10403,N_10245);
nand U11022 (N_11022,N_10945,N_10727);
nor U11023 (N_11023,N_10733,N_10590);
xor U11024 (N_11024,N_10490,N_10330);
nand U11025 (N_11025,N_10576,N_10939);
nor U11026 (N_11026,N_10775,N_10482);
or U11027 (N_11027,N_10131,N_10595);
nor U11028 (N_11028,N_10630,N_10253);
xnor U11029 (N_11029,N_10056,N_10813);
or U11030 (N_11030,N_10410,N_10903);
or U11031 (N_11031,N_10571,N_10445);
xnor U11032 (N_11032,N_10462,N_10802);
and U11033 (N_11033,N_10913,N_10326);
xnor U11034 (N_11034,N_10845,N_10844);
and U11035 (N_11035,N_10295,N_10277);
or U11036 (N_11036,N_10758,N_10201);
and U11037 (N_11037,N_10192,N_10161);
xnor U11038 (N_11038,N_10616,N_10070);
nand U11039 (N_11039,N_10950,N_10661);
nor U11040 (N_11040,N_10264,N_10494);
or U11041 (N_11041,N_10646,N_10987);
nor U11042 (N_11042,N_10202,N_10804);
or U11043 (N_11043,N_10214,N_10271);
or U11044 (N_11044,N_10140,N_10256);
nor U11045 (N_11045,N_10650,N_10074);
or U11046 (N_11046,N_10088,N_10918);
nand U11047 (N_11047,N_10355,N_10561);
nand U11048 (N_11048,N_10533,N_10626);
or U11049 (N_11049,N_10284,N_10467);
or U11050 (N_11050,N_10760,N_10675);
and U11051 (N_11051,N_10439,N_10560);
nor U11052 (N_11052,N_10696,N_10999);
or U11053 (N_11053,N_10027,N_10091);
and U11054 (N_11054,N_10316,N_10783);
and U11055 (N_11055,N_10266,N_10923);
or U11056 (N_11056,N_10236,N_10772);
nand U11057 (N_11057,N_10904,N_10437);
nor U11058 (N_11058,N_10877,N_10511);
nand U11059 (N_11059,N_10717,N_10633);
or U11060 (N_11060,N_10838,N_10528);
and U11061 (N_11061,N_10773,N_10833);
nand U11062 (N_11062,N_10397,N_10198);
and U11063 (N_11063,N_10384,N_10208);
and U11064 (N_11064,N_10247,N_10108);
xor U11065 (N_11065,N_10183,N_10715);
nor U11066 (N_11066,N_10151,N_10374);
nand U11067 (N_11067,N_10710,N_10159);
xnor U11068 (N_11068,N_10888,N_10433);
and U11069 (N_11069,N_10468,N_10573);
xnor U11070 (N_11070,N_10029,N_10390);
nor U11071 (N_11071,N_10980,N_10244);
and U11072 (N_11072,N_10669,N_10363);
xnor U11073 (N_11073,N_10509,N_10102);
or U11074 (N_11074,N_10246,N_10185);
nor U11075 (N_11075,N_10113,N_10221);
xnor U11076 (N_11076,N_10178,N_10143);
nor U11077 (N_11077,N_10642,N_10354);
nand U11078 (N_11078,N_10288,N_10603);
and U11079 (N_11079,N_10976,N_10181);
xnor U11080 (N_11080,N_10972,N_10078);
or U11081 (N_11081,N_10932,N_10432);
nand U11082 (N_11082,N_10926,N_10891);
or U11083 (N_11083,N_10705,N_10825);
and U11084 (N_11084,N_10228,N_10435);
and U11085 (N_11085,N_10507,N_10971);
and U11086 (N_11086,N_10790,N_10726);
and U11087 (N_11087,N_10150,N_10379);
nand U11088 (N_11088,N_10006,N_10216);
nor U11089 (N_11089,N_10128,N_10352);
xor U11090 (N_11090,N_10578,N_10177);
xor U11091 (N_11091,N_10062,N_10165);
nand U11092 (N_11092,N_10522,N_10491);
nor U11093 (N_11093,N_10232,N_10752);
or U11094 (N_11094,N_10430,N_10529);
or U11095 (N_11095,N_10520,N_10171);
and U11096 (N_11096,N_10089,N_10551);
and U11097 (N_11097,N_10541,N_10919);
nor U11098 (N_11098,N_10855,N_10552);
nand U11099 (N_11099,N_10739,N_10031);
or U11100 (N_11100,N_10584,N_10200);
nor U11101 (N_11101,N_10423,N_10624);
and U11102 (N_11102,N_10883,N_10470);
nor U11103 (N_11103,N_10392,N_10729);
or U11104 (N_11104,N_10530,N_10377);
nand U11105 (N_11105,N_10686,N_10534);
and U11106 (N_11106,N_10519,N_10536);
nand U11107 (N_11107,N_10080,N_10863);
nand U11108 (N_11108,N_10979,N_10900);
or U11109 (N_11109,N_10187,N_10110);
or U11110 (N_11110,N_10645,N_10957);
and U11111 (N_11111,N_10780,N_10428);
and U11112 (N_11112,N_10369,N_10385);
or U11113 (N_11113,N_10254,N_10978);
nor U11114 (N_11114,N_10587,N_10606);
or U11115 (N_11115,N_10938,N_10149);
and U11116 (N_11116,N_10071,N_10389);
and U11117 (N_11117,N_10871,N_10231);
nand U11118 (N_11118,N_10851,N_10698);
nand U11119 (N_11119,N_10521,N_10010);
or U11120 (N_11120,N_10543,N_10882);
or U11121 (N_11121,N_10378,N_10087);
or U11122 (N_11122,N_10142,N_10914);
nor U11123 (N_11123,N_10960,N_10417);
nand U11124 (N_11124,N_10670,N_10864);
xnor U11125 (N_11125,N_10865,N_10836);
and U11126 (N_11126,N_10505,N_10180);
xnor U11127 (N_11127,N_10073,N_10398);
nor U11128 (N_11128,N_10513,N_10688);
nand U11129 (N_11129,N_10699,N_10302);
and U11130 (N_11130,N_10317,N_10693);
nor U11131 (N_11131,N_10328,N_10082);
and U11132 (N_11132,N_10801,N_10342);
and U11133 (N_11133,N_10592,N_10407);
xnor U11134 (N_11134,N_10209,N_10860);
xnor U11135 (N_11135,N_10337,N_10810);
or U11136 (N_11136,N_10689,N_10568);
or U11137 (N_11137,N_10600,N_10627);
xnor U11138 (N_11138,N_10408,N_10213);
and U11139 (N_11139,N_10340,N_10554);
xnor U11140 (N_11140,N_10371,N_10781);
and U11141 (N_11141,N_10105,N_10365);
nand U11142 (N_11142,N_10125,N_10963);
xnor U11143 (N_11143,N_10964,N_10173);
and U11144 (N_11144,N_10459,N_10373);
xnor U11145 (N_11145,N_10443,N_10740);
nor U11146 (N_11146,N_10596,N_10096);
or U11147 (N_11147,N_10925,N_10771);
nor U11148 (N_11148,N_10479,N_10949);
and U11149 (N_11149,N_10765,N_10709);
or U11150 (N_11150,N_10820,N_10147);
nand U11151 (N_11151,N_10424,N_10158);
and U11152 (N_11152,N_10063,N_10997);
or U11153 (N_11153,N_10255,N_10719);
nand U11154 (N_11154,N_10233,N_10313);
nor U11155 (N_11155,N_10906,N_10803);
xnor U11156 (N_11156,N_10629,N_10970);
and U11157 (N_11157,N_10792,N_10872);
xor U11158 (N_11158,N_10039,N_10191);
nand U11159 (N_11159,N_10953,N_10297);
nor U11160 (N_11160,N_10644,N_10665);
nand U11161 (N_11161,N_10793,N_10867);
xor U11162 (N_11162,N_10283,N_10962);
nor U11163 (N_11163,N_10955,N_10602);
nor U11164 (N_11164,N_10251,N_10805);
xnor U11165 (N_11165,N_10120,N_10744);
nand U11166 (N_11166,N_10589,N_10653);
nor U11167 (N_11167,N_10898,N_10707);
and U11168 (N_11168,N_10811,N_10609);
or U11169 (N_11169,N_10655,N_10098);
and U11170 (N_11170,N_10224,N_10037);
or U11171 (N_11171,N_10144,N_10920);
or U11172 (N_11172,N_10751,N_10040);
nor U11173 (N_11173,N_10893,N_10493);
nand U11174 (N_11174,N_10672,N_10455);
xnor U11175 (N_11175,N_10935,N_10054);
xnor U11176 (N_11176,N_10380,N_10025);
xnor U11177 (N_11177,N_10267,N_10270);
nor U11178 (N_11178,N_10262,N_10123);
or U11179 (N_11179,N_10307,N_10303);
xor U11180 (N_11180,N_10831,N_10639);
and U11181 (N_11181,N_10512,N_10287);
nor U11182 (N_11182,N_10614,N_10721);
nor U11183 (N_11183,N_10387,N_10975);
nand U11184 (N_11184,N_10166,N_10931);
and U11185 (N_11185,N_10003,N_10930);
xnor U11186 (N_11186,N_10077,N_10796);
nand U11187 (N_11187,N_10876,N_10204);
xor U11188 (N_11188,N_10759,N_10514);
xor U11189 (N_11189,N_10023,N_10856);
nand U11190 (N_11190,N_10104,N_10222);
nand U11191 (N_11191,N_10212,N_10857);
nand U11192 (N_11192,N_10357,N_10821);
or U11193 (N_11193,N_10032,N_10167);
nor U11194 (N_11194,N_10084,N_10958);
or U11195 (N_11195,N_10299,N_10118);
and U11196 (N_11196,N_10273,N_10632);
and U11197 (N_11197,N_10094,N_10446);
and U11198 (N_11198,N_10687,N_10263);
nand U11199 (N_11199,N_10059,N_10436);
and U11200 (N_11200,N_10924,N_10984);
and U11201 (N_11201,N_10358,N_10902);
nand U11202 (N_11202,N_10853,N_10878);
nand U11203 (N_11203,N_10763,N_10948);
and U11204 (N_11204,N_10890,N_10818);
nor U11205 (N_11205,N_10974,N_10572);
and U11206 (N_11206,N_10656,N_10683);
nor U11207 (N_11207,N_10591,N_10806);
nor U11208 (N_11208,N_10874,N_10449);
nor U11209 (N_11209,N_10637,N_10830);
nor U11210 (N_11210,N_10476,N_10196);
nand U11211 (N_11211,N_10829,N_10993);
and U11212 (N_11212,N_10557,N_10034);
or U11213 (N_11213,N_10314,N_10002);
xnor U11214 (N_11214,N_10359,N_10296);
or U11215 (N_11215,N_10393,N_10137);
nand U11216 (N_11216,N_10947,N_10635);
and U11217 (N_11217,N_10362,N_10915);
nand U11218 (N_11218,N_10608,N_10356);
nand U11219 (N_11219,N_10463,N_10553);
nand U11220 (N_11220,N_10329,N_10441);
nor U11221 (N_11221,N_10788,N_10986);
and U11222 (N_11222,N_10109,N_10910);
or U11223 (N_11223,N_10237,N_10638);
or U11224 (N_11224,N_10366,N_10794);
and U11225 (N_11225,N_10179,N_10946);
nor U11226 (N_11226,N_10164,N_10723);
or U11227 (N_11227,N_10647,N_10823);
xnor U11228 (N_11228,N_10722,N_10927);
and U11229 (N_11229,N_10260,N_10017);
nor U11230 (N_11230,N_10812,N_10009);
nand U11231 (N_11231,N_10444,N_10549);
nand U11232 (N_11232,N_10532,N_10701);
nor U11233 (N_11233,N_10897,N_10827);
xnor U11234 (N_11234,N_10956,N_10086);
nand U11235 (N_11235,N_10992,N_10097);
or U11236 (N_11236,N_10848,N_10839);
nor U11237 (N_11237,N_10879,N_10658);
or U11238 (N_11238,N_10481,N_10767);
or U11239 (N_11239,N_10779,N_10038);
xor U11240 (N_11240,N_10524,N_10382);
or U11241 (N_11241,N_10737,N_10907);
and U11242 (N_11242,N_10988,N_10716);
nand U11243 (N_11243,N_10967,N_10570);
and U11244 (N_11244,N_10585,N_10319);
and U11245 (N_11245,N_10990,N_10160);
nor U11246 (N_11246,N_10840,N_10119);
and U11247 (N_11247,N_10239,N_10757);
nor U11248 (N_11248,N_10341,N_10562);
nor U11249 (N_11249,N_10996,N_10269);
or U11250 (N_11250,N_10613,N_10426);
nand U11251 (N_11251,N_10092,N_10474);
nand U11252 (N_11252,N_10115,N_10598);
or U11253 (N_11253,N_10345,N_10995);
nor U11254 (N_11254,N_10282,N_10103);
or U11255 (N_11255,N_10126,N_10045);
nor U11256 (N_11256,N_10730,N_10951);
xor U11257 (N_11257,N_10268,N_10048);
xnor U11258 (N_11258,N_10667,N_10004);
nand U11259 (N_11259,N_10461,N_10861);
nor U11260 (N_11260,N_10538,N_10257);
xnor U11261 (N_11261,N_10155,N_10581);
xor U11262 (N_11262,N_10170,N_10132);
xor U11263 (N_11263,N_10989,N_10484);
nand U11264 (N_11264,N_10336,N_10193);
xnor U11265 (N_11265,N_10375,N_10674);
and U11266 (N_11266,N_10005,N_10916);
or U11267 (N_11267,N_10873,N_10692);
nor U11268 (N_11268,N_10220,N_10184);
nor U11269 (N_11269,N_10024,N_10607);
xor U11270 (N_11270,N_10046,N_10605);
and U11271 (N_11271,N_10697,N_10517);
or U11272 (N_11272,N_10242,N_10425);
nor U11273 (N_11273,N_10289,N_10936);
and U11274 (N_11274,N_10406,N_10518);
and U11275 (N_11275,N_10998,N_10207);
xor U11276 (N_11276,N_10769,N_10133);
and U11277 (N_11277,N_10011,N_10574);
nand U11278 (N_11278,N_10537,N_10346);
nor U11279 (N_11279,N_10708,N_10069);
or U11280 (N_11280,N_10725,N_10899);
and U11281 (N_11281,N_10047,N_10654);
or U11282 (N_11282,N_10298,N_10895);
xnor U11283 (N_11283,N_10594,N_10621);
nand U11284 (N_11284,N_10977,N_10418);
nand U11285 (N_11285,N_10162,N_10368);
and U11286 (N_11286,N_10318,N_10203);
nor U11287 (N_11287,N_10300,N_10413);
or U11288 (N_11288,N_10286,N_10168);
xnor U11289 (N_11289,N_10555,N_10217);
or U11290 (N_11290,N_10388,N_10350);
or U11291 (N_11291,N_10559,N_10703);
nor U11292 (N_11292,N_10422,N_10064);
nor U11293 (N_11293,N_10886,N_10896);
xor U11294 (N_11294,N_10643,N_10186);
or U11295 (N_11295,N_10146,N_10272);
xor U11296 (N_11296,N_10421,N_10019);
nand U11297 (N_11297,N_10101,N_10335);
nand U11298 (N_11298,N_10364,N_10485);
or U11299 (N_11299,N_10824,N_10367);
xor U11300 (N_11300,N_10542,N_10593);
and U11301 (N_11301,N_10226,N_10007);
or U11302 (N_11302,N_10745,N_10000);
and U11303 (N_11303,N_10814,N_10312);
and U11304 (N_11304,N_10498,N_10841);
or U11305 (N_11305,N_10129,N_10782);
or U11306 (N_11306,N_10205,N_10199);
or U11307 (N_11307,N_10145,N_10016);
nor U11308 (N_11308,N_10588,N_10660);
nor U11309 (N_11309,N_10500,N_10741);
and U11310 (N_11310,N_10718,N_10416);
and U11311 (N_11311,N_10933,N_10107);
nand U11312 (N_11312,N_10457,N_10210);
or U11313 (N_11313,N_10136,N_10100);
and U11314 (N_11314,N_10651,N_10415);
xor U11315 (N_11315,N_10234,N_10525);
or U11316 (N_11316,N_10837,N_10291);
and U11317 (N_11317,N_10501,N_10981);
nor U11318 (N_11318,N_10442,N_10376);
nand U11319 (N_11319,N_10784,N_10447);
nand U11320 (N_11320,N_10545,N_10473);
or U11321 (N_11321,N_10305,N_10440);
and U11322 (N_11322,N_10968,N_10394);
and U11323 (N_11323,N_10453,N_10973);
and U11324 (N_11324,N_10361,N_10405);
or U11325 (N_11325,N_10130,N_10952);
and U11326 (N_11326,N_10250,N_10321);
xnor U11327 (N_11327,N_10750,N_10323);
xnor U11328 (N_11328,N_10539,N_10404);
nand U11329 (N_11329,N_10051,N_10747);
and U11330 (N_11330,N_10912,N_10666);
nand U11331 (N_11331,N_10465,N_10535);
nand U11332 (N_11332,N_10580,N_10499);
xnor U11333 (N_11333,N_10736,N_10612);
nand U11334 (N_11334,N_10795,N_10122);
nand U11335 (N_11335,N_10567,N_10905);
nor U11336 (N_11336,N_10526,N_10035);
or U11337 (N_11337,N_10333,N_10157);
or U11338 (N_11338,N_10049,N_10911);
xor U11339 (N_11339,N_10175,N_10043);
nand U11340 (N_11340,N_10564,N_10869);
or U11341 (N_11341,N_10940,N_10219);
nand U11342 (N_11342,N_10420,N_10954);
nand U11343 (N_11343,N_10664,N_10657);
and U11344 (N_11344,N_10649,N_10480);
nor U11345 (N_11345,N_10106,N_10116);
or U11346 (N_11346,N_10339,N_10431);
and U11347 (N_11347,N_10994,N_10351);
xor U11348 (N_11348,N_10402,N_10922);
xor U11349 (N_11349,N_10134,N_10875);
xnor U11350 (N_11350,N_10597,N_10348);
nand U11351 (N_11351,N_10859,N_10309);
or U11352 (N_11352,N_10885,N_10248);
nor U11353 (N_11353,N_10785,N_10182);
xor U11354 (N_11354,N_10227,N_10847);
or U11355 (N_11355,N_10460,N_10141);
xnor U11356 (N_11356,N_10391,N_10067);
and U11357 (N_11357,N_10755,N_10053);
and U11358 (N_11358,N_10172,N_10189);
xnor U11359 (N_11359,N_10152,N_10799);
nand U11360 (N_11360,N_10884,N_10659);
nor U11361 (N_11361,N_10527,N_10235);
or U11362 (N_11362,N_10566,N_10929);
nand U11363 (N_11363,N_10112,N_10061);
nand U11364 (N_11364,N_10732,N_10343);
or U11365 (N_11365,N_10349,N_10502);
xnor U11366 (N_11366,N_10058,N_10471);
xor U11367 (N_11367,N_10301,N_10076);
nor U11368 (N_11368,N_10546,N_10060);
and U11369 (N_11369,N_10617,N_10866);
nand U11370 (N_11370,N_10206,N_10983);
or U11371 (N_11371,N_10095,N_10036);
xnor U11372 (N_11372,N_10917,N_10325);
and U11373 (N_11373,N_10072,N_10768);
nor U11374 (N_11374,N_10488,N_10832);
xor U11375 (N_11375,N_10754,N_10791);
and U11376 (N_11376,N_10776,N_10748);
nor U11377 (N_11377,N_10258,N_10909);
or U11378 (N_11378,N_10969,N_10815);
and U11379 (N_11379,N_10743,N_10135);
xor U11380 (N_11380,N_10714,N_10961);
nor U11381 (N_11381,N_10809,N_10575);
nand U11382 (N_11382,N_10079,N_10464);
and U11383 (N_11383,N_10887,N_10153);
nand U11384 (N_11384,N_10679,N_10372);
and U11385 (N_11385,N_10618,N_10695);
xnor U11386 (N_11386,N_10921,N_10241);
or U11387 (N_11387,N_10414,N_10290);
nor U11388 (N_11388,N_10894,N_10676);
or U11389 (N_11389,N_10711,N_10991);
nand U11390 (N_11390,N_10044,N_10706);
and U11391 (N_11391,N_10691,N_10252);
and U11392 (N_11392,N_10928,N_10569);
nor U11393 (N_11393,N_10579,N_10764);
nor U11394 (N_11394,N_10834,N_10489);
and U11395 (N_11395,N_10742,N_10817);
and U11396 (N_11396,N_10451,N_10756);
nand U11397 (N_11397,N_10483,N_10409);
xnor U11398 (N_11398,N_10556,N_10028);
xnor U11399 (N_11399,N_10148,N_10169);
nand U11400 (N_11400,N_10127,N_10344);
nor U11401 (N_11401,N_10456,N_10360);
and U11402 (N_11402,N_10276,N_10544);
nand U11403 (N_11403,N_10506,N_10327);
and U11404 (N_11404,N_10117,N_10050);
nor U11405 (N_11405,N_10322,N_10448);
and U11406 (N_11406,N_10429,N_10753);
xnor U11407 (N_11407,N_10800,N_10586);
nor U11408 (N_11408,N_10176,N_10475);
or U11409 (N_11409,N_10066,N_10582);
xnor U11410 (N_11410,N_10901,N_10819);
or U11411 (N_11411,N_10515,N_10215);
nand U11412 (N_11412,N_10636,N_10041);
nand U11413 (N_11413,N_10188,N_10868);
nor U11414 (N_11414,N_10749,N_10477);
and U11415 (N_11415,N_10280,N_10826);
or U11416 (N_11416,N_10469,N_10563);
or U11417 (N_11417,N_10770,N_10583);
nand U11418 (N_11418,N_10419,N_10353);
nand U11419 (N_11419,N_10001,N_10965);
nor U11420 (N_11420,N_10293,N_10620);
and U11421 (N_11421,N_10862,N_10540);
xnor U11422 (N_11422,N_10678,N_10816);
xnor U11423 (N_11423,N_10450,N_10828);
or U11424 (N_11424,N_10854,N_10685);
nor U11425 (N_11425,N_10728,N_10503);
nor U11426 (N_11426,N_10982,N_10842);
xnor U11427 (N_11427,N_10281,N_10713);
or U11428 (N_11428,N_10395,N_10662);
or U11429 (N_11429,N_10850,N_10766);
or U11430 (N_11430,N_10121,N_10849);
xnor U11431 (N_11431,N_10332,N_10194);
nand U11432 (N_11432,N_10648,N_10261);
nor U11433 (N_11433,N_10230,N_10304);
nor U11434 (N_11434,N_10677,N_10611);
xor U11435 (N_11435,N_10383,N_10684);
nand U11436 (N_11436,N_10099,N_10808);
or U11437 (N_11437,N_10195,N_10531);
nor U11438 (N_11438,N_10020,N_10265);
xor U11439 (N_11439,N_10163,N_10496);
and U11440 (N_11440,N_10673,N_10347);
or U11441 (N_11441,N_10274,N_10787);
and U11442 (N_11442,N_10240,N_10012);
or U11443 (N_11443,N_10454,N_10731);
or U11444 (N_11444,N_10704,N_10640);
or U11445 (N_11445,N_10604,N_10033);
nand U11446 (N_11446,N_10174,N_10777);
nand U11447 (N_11447,N_10504,N_10712);
nor U11448 (N_11448,N_10229,N_10052);
nor U11449 (N_11449,N_10497,N_10937);
or U11450 (N_11450,N_10941,N_10934);
xor U11451 (N_11451,N_10324,N_10279);
xor U11452 (N_11452,N_10623,N_10495);
xnor U11453 (N_11453,N_10680,N_10797);
or U11454 (N_11454,N_10015,N_10682);
xor U11455 (N_11455,N_10628,N_10786);
and U11456 (N_11456,N_10399,N_10278);
or U11457 (N_11457,N_10478,N_10197);
nand U11458 (N_11458,N_10139,N_10558);
nand U11459 (N_11459,N_10746,N_10652);
or U11460 (N_11460,N_10294,N_10021);
nor U11461 (N_11461,N_10370,N_10065);
and U11462 (N_11462,N_10880,N_10452);
xor U11463 (N_11463,N_10550,N_10310);
or U11464 (N_11464,N_10401,N_10663);
and U11465 (N_11465,N_10516,N_10014);
nand U11466 (N_11466,N_10822,N_10625);
nor U11467 (N_11467,N_10668,N_10013);
nand U11468 (N_11468,N_10427,N_10487);
nor U11469 (N_11469,N_10386,N_10285);
xor U11470 (N_11470,N_10852,N_10681);
xor U11471 (N_11471,N_10858,N_10311);
xor U11472 (N_11472,N_10090,N_10111);
xor U11473 (N_11473,N_10466,N_10190);
xnor U11474 (N_11474,N_10738,N_10238);
or U11475 (N_11475,N_10547,N_10124);
nand U11476 (N_11476,N_10085,N_10486);
and U11477 (N_11477,N_10690,N_10412);
nand U11478 (N_11478,N_10846,N_10154);
xnor U11479 (N_11479,N_10114,N_10548);
or U11480 (N_11480,N_10778,N_10942);
and U11481 (N_11481,N_10774,N_10761);
nor U11482 (N_11482,N_10225,N_10944);
or U11483 (N_11483,N_10138,N_10985);
or U11484 (N_11484,N_10083,N_10615);
nand U11485 (N_11485,N_10068,N_10641);
xnor U11486 (N_11486,N_10601,N_10042);
nor U11487 (N_11487,N_10308,N_10762);
xnor U11488 (N_11488,N_10523,N_10081);
and U11489 (N_11489,N_10030,N_10634);
nor U11490 (N_11490,N_10700,N_10434);
or U11491 (N_11491,N_10211,N_10702);
or U11492 (N_11492,N_10734,N_10018);
xor U11493 (N_11493,N_10026,N_10908);
or U11494 (N_11494,N_10243,N_10458);
nor U11495 (N_11495,N_10892,N_10622);
xnor U11496 (N_11496,N_10411,N_10724);
nor U11497 (N_11497,N_10334,N_10631);
nand U11498 (N_11498,N_10055,N_10320);
nand U11499 (N_11499,N_10259,N_10472);
xnor U11500 (N_11500,N_10159,N_10117);
nand U11501 (N_11501,N_10189,N_10910);
nor U11502 (N_11502,N_10088,N_10934);
nor U11503 (N_11503,N_10391,N_10506);
nor U11504 (N_11504,N_10826,N_10609);
nand U11505 (N_11505,N_10822,N_10848);
nand U11506 (N_11506,N_10201,N_10998);
xnor U11507 (N_11507,N_10045,N_10741);
xnor U11508 (N_11508,N_10085,N_10871);
and U11509 (N_11509,N_10363,N_10306);
xor U11510 (N_11510,N_10837,N_10598);
and U11511 (N_11511,N_10709,N_10088);
nand U11512 (N_11512,N_10149,N_10411);
or U11513 (N_11513,N_10144,N_10673);
or U11514 (N_11514,N_10539,N_10752);
nor U11515 (N_11515,N_10822,N_10576);
and U11516 (N_11516,N_10946,N_10403);
and U11517 (N_11517,N_10730,N_10230);
xnor U11518 (N_11518,N_10872,N_10189);
or U11519 (N_11519,N_10809,N_10876);
and U11520 (N_11520,N_10884,N_10954);
and U11521 (N_11521,N_10252,N_10514);
and U11522 (N_11522,N_10009,N_10703);
or U11523 (N_11523,N_10786,N_10918);
nor U11524 (N_11524,N_10710,N_10067);
nor U11525 (N_11525,N_10400,N_10166);
nand U11526 (N_11526,N_10168,N_10520);
nor U11527 (N_11527,N_10291,N_10838);
xnor U11528 (N_11528,N_10627,N_10982);
nand U11529 (N_11529,N_10046,N_10071);
or U11530 (N_11530,N_10052,N_10498);
nand U11531 (N_11531,N_10613,N_10286);
and U11532 (N_11532,N_10097,N_10054);
xnor U11533 (N_11533,N_10997,N_10102);
and U11534 (N_11534,N_10107,N_10941);
or U11535 (N_11535,N_10452,N_10385);
nor U11536 (N_11536,N_10523,N_10371);
nor U11537 (N_11537,N_10391,N_10843);
and U11538 (N_11538,N_10279,N_10603);
and U11539 (N_11539,N_10074,N_10694);
or U11540 (N_11540,N_10112,N_10948);
nor U11541 (N_11541,N_10506,N_10354);
nand U11542 (N_11542,N_10388,N_10139);
and U11543 (N_11543,N_10110,N_10512);
nand U11544 (N_11544,N_10360,N_10266);
nor U11545 (N_11545,N_10771,N_10589);
and U11546 (N_11546,N_10051,N_10970);
nand U11547 (N_11547,N_10129,N_10563);
nand U11548 (N_11548,N_10927,N_10034);
nor U11549 (N_11549,N_10002,N_10605);
xor U11550 (N_11550,N_10463,N_10655);
xnor U11551 (N_11551,N_10457,N_10610);
or U11552 (N_11552,N_10974,N_10888);
or U11553 (N_11553,N_10999,N_10284);
and U11554 (N_11554,N_10375,N_10900);
xnor U11555 (N_11555,N_10194,N_10279);
nand U11556 (N_11556,N_10673,N_10019);
nor U11557 (N_11557,N_10102,N_10715);
or U11558 (N_11558,N_10682,N_10157);
or U11559 (N_11559,N_10050,N_10870);
and U11560 (N_11560,N_10867,N_10035);
nor U11561 (N_11561,N_10968,N_10566);
and U11562 (N_11562,N_10807,N_10513);
nor U11563 (N_11563,N_10254,N_10356);
or U11564 (N_11564,N_10518,N_10530);
nor U11565 (N_11565,N_10358,N_10927);
or U11566 (N_11566,N_10259,N_10192);
xor U11567 (N_11567,N_10747,N_10219);
nor U11568 (N_11568,N_10522,N_10306);
and U11569 (N_11569,N_10722,N_10096);
nor U11570 (N_11570,N_10407,N_10259);
or U11571 (N_11571,N_10435,N_10735);
nand U11572 (N_11572,N_10529,N_10698);
nand U11573 (N_11573,N_10238,N_10423);
nor U11574 (N_11574,N_10485,N_10646);
nand U11575 (N_11575,N_10050,N_10490);
and U11576 (N_11576,N_10935,N_10640);
xor U11577 (N_11577,N_10683,N_10064);
or U11578 (N_11578,N_10659,N_10051);
or U11579 (N_11579,N_10531,N_10631);
nand U11580 (N_11580,N_10589,N_10893);
and U11581 (N_11581,N_10454,N_10743);
xnor U11582 (N_11582,N_10402,N_10521);
and U11583 (N_11583,N_10589,N_10236);
and U11584 (N_11584,N_10716,N_10398);
or U11585 (N_11585,N_10941,N_10719);
or U11586 (N_11586,N_10977,N_10616);
and U11587 (N_11587,N_10743,N_10702);
or U11588 (N_11588,N_10852,N_10250);
nor U11589 (N_11589,N_10802,N_10579);
xnor U11590 (N_11590,N_10274,N_10696);
nand U11591 (N_11591,N_10792,N_10141);
and U11592 (N_11592,N_10197,N_10943);
and U11593 (N_11593,N_10458,N_10235);
nand U11594 (N_11594,N_10067,N_10021);
xnor U11595 (N_11595,N_10017,N_10331);
or U11596 (N_11596,N_10386,N_10502);
or U11597 (N_11597,N_10228,N_10136);
or U11598 (N_11598,N_10433,N_10409);
xnor U11599 (N_11599,N_10570,N_10406);
and U11600 (N_11600,N_10576,N_10633);
and U11601 (N_11601,N_10419,N_10722);
xnor U11602 (N_11602,N_10609,N_10705);
nand U11603 (N_11603,N_10044,N_10411);
nand U11604 (N_11604,N_10006,N_10549);
nor U11605 (N_11605,N_10510,N_10434);
or U11606 (N_11606,N_10979,N_10444);
xnor U11607 (N_11607,N_10807,N_10876);
nand U11608 (N_11608,N_10955,N_10961);
nor U11609 (N_11609,N_10094,N_10591);
xor U11610 (N_11610,N_10785,N_10094);
nand U11611 (N_11611,N_10107,N_10750);
or U11612 (N_11612,N_10950,N_10159);
and U11613 (N_11613,N_10926,N_10624);
nor U11614 (N_11614,N_10757,N_10306);
or U11615 (N_11615,N_10304,N_10547);
or U11616 (N_11616,N_10243,N_10250);
xor U11617 (N_11617,N_10146,N_10720);
or U11618 (N_11618,N_10260,N_10642);
nor U11619 (N_11619,N_10436,N_10024);
xnor U11620 (N_11620,N_10423,N_10723);
or U11621 (N_11621,N_10628,N_10111);
xnor U11622 (N_11622,N_10494,N_10262);
xnor U11623 (N_11623,N_10902,N_10948);
xor U11624 (N_11624,N_10529,N_10884);
and U11625 (N_11625,N_10699,N_10105);
nor U11626 (N_11626,N_10679,N_10146);
nand U11627 (N_11627,N_10402,N_10934);
nand U11628 (N_11628,N_10799,N_10248);
or U11629 (N_11629,N_10692,N_10969);
nand U11630 (N_11630,N_10334,N_10340);
and U11631 (N_11631,N_10051,N_10814);
or U11632 (N_11632,N_10104,N_10466);
or U11633 (N_11633,N_10984,N_10896);
or U11634 (N_11634,N_10213,N_10000);
xor U11635 (N_11635,N_10240,N_10950);
nand U11636 (N_11636,N_10979,N_10863);
or U11637 (N_11637,N_10402,N_10130);
and U11638 (N_11638,N_10412,N_10135);
nand U11639 (N_11639,N_10949,N_10079);
nand U11640 (N_11640,N_10051,N_10987);
or U11641 (N_11641,N_10343,N_10185);
xor U11642 (N_11642,N_10428,N_10568);
or U11643 (N_11643,N_10949,N_10091);
nor U11644 (N_11644,N_10756,N_10008);
and U11645 (N_11645,N_10533,N_10539);
nand U11646 (N_11646,N_10486,N_10086);
nor U11647 (N_11647,N_10849,N_10104);
nor U11648 (N_11648,N_10553,N_10808);
and U11649 (N_11649,N_10378,N_10070);
nand U11650 (N_11650,N_10944,N_10932);
or U11651 (N_11651,N_10502,N_10444);
xor U11652 (N_11652,N_10456,N_10218);
or U11653 (N_11653,N_10688,N_10360);
xor U11654 (N_11654,N_10308,N_10038);
nor U11655 (N_11655,N_10894,N_10532);
or U11656 (N_11656,N_10874,N_10191);
and U11657 (N_11657,N_10504,N_10237);
or U11658 (N_11658,N_10717,N_10900);
and U11659 (N_11659,N_10935,N_10410);
and U11660 (N_11660,N_10819,N_10005);
nand U11661 (N_11661,N_10966,N_10266);
and U11662 (N_11662,N_10465,N_10323);
nand U11663 (N_11663,N_10444,N_10410);
nor U11664 (N_11664,N_10967,N_10349);
or U11665 (N_11665,N_10977,N_10854);
and U11666 (N_11666,N_10550,N_10578);
nand U11667 (N_11667,N_10853,N_10432);
xor U11668 (N_11668,N_10270,N_10035);
nand U11669 (N_11669,N_10040,N_10149);
nor U11670 (N_11670,N_10955,N_10513);
nor U11671 (N_11671,N_10028,N_10090);
xor U11672 (N_11672,N_10260,N_10987);
nor U11673 (N_11673,N_10505,N_10562);
xor U11674 (N_11674,N_10008,N_10223);
nand U11675 (N_11675,N_10356,N_10942);
or U11676 (N_11676,N_10716,N_10247);
and U11677 (N_11677,N_10477,N_10695);
or U11678 (N_11678,N_10974,N_10182);
and U11679 (N_11679,N_10980,N_10650);
or U11680 (N_11680,N_10587,N_10842);
and U11681 (N_11681,N_10756,N_10696);
or U11682 (N_11682,N_10414,N_10309);
nand U11683 (N_11683,N_10581,N_10027);
xnor U11684 (N_11684,N_10439,N_10298);
or U11685 (N_11685,N_10139,N_10028);
xnor U11686 (N_11686,N_10405,N_10794);
and U11687 (N_11687,N_10609,N_10301);
xnor U11688 (N_11688,N_10000,N_10479);
or U11689 (N_11689,N_10590,N_10683);
xor U11690 (N_11690,N_10508,N_10109);
xnor U11691 (N_11691,N_10273,N_10824);
xnor U11692 (N_11692,N_10043,N_10448);
nor U11693 (N_11693,N_10086,N_10461);
xor U11694 (N_11694,N_10310,N_10747);
or U11695 (N_11695,N_10307,N_10041);
nand U11696 (N_11696,N_10641,N_10205);
xor U11697 (N_11697,N_10031,N_10014);
or U11698 (N_11698,N_10756,N_10723);
xnor U11699 (N_11699,N_10695,N_10729);
xnor U11700 (N_11700,N_10820,N_10797);
nor U11701 (N_11701,N_10791,N_10563);
and U11702 (N_11702,N_10276,N_10669);
nor U11703 (N_11703,N_10469,N_10902);
or U11704 (N_11704,N_10942,N_10601);
and U11705 (N_11705,N_10861,N_10592);
nor U11706 (N_11706,N_10739,N_10184);
xor U11707 (N_11707,N_10757,N_10975);
nand U11708 (N_11708,N_10772,N_10976);
nor U11709 (N_11709,N_10723,N_10492);
nand U11710 (N_11710,N_10144,N_10399);
nand U11711 (N_11711,N_10769,N_10863);
and U11712 (N_11712,N_10870,N_10901);
and U11713 (N_11713,N_10294,N_10180);
xor U11714 (N_11714,N_10601,N_10143);
xnor U11715 (N_11715,N_10418,N_10274);
or U11716 (N_11716,N_10929,N_10439);
nor U11717 (N_11717,N_10815,N_10022);
nor U11718 (N_11718,N_10545,N_10397);
xor U11719 (N_11719,N_10301,N_10859);
or U11720 (N_11720,N_10936,N_10443);
xor U11721 (N_11721,N_10641,N_10662);
or U11722 (N_11722,N_10710,N_10728);
xnor U11723 (N_11723,N_10580,N_10768);
nand U11724 (N_11724,N_10452,N_10066);
nand U11725 (N_11725,N_10665,N_10714);
nand U11726 (N_11726,N_10538,N_10605);
nor U11727 (N_11727,N_10083,N_10324);
nor U11728 (N_11728,N_10882,N_10474);
and U11729 (N_11729,N_10748,N_10205);
nor U11730 (N_11730,N_10481,N_10304);
nor U11731 (N_11731,N_10091,N_10817);
and U11732 (N_11732,N_10201,N_10288);
or U11733 (N_11733,N_10861,N_10625);
and U11734 (N_11734,N_10221,N_10810);
or U11735 (N_11735,N_10510,N_10974);
and U11736 (N_11736,N_10099,N_10125);
nor U11737 (N_11737,N_10956,N_10976);
or U11738 (N_11738,N_10503,N_10757);
xnor U11739 (N_11739,N_10639,N_10144);
xor U11740 (N_11740,N_10425,N_10719);
xor U11741 (N_11741,N_10850,N_10958);
nor U11742 (N_11742,N_10754,N_10536);
and U11743 (N_11743,N_10290,N_10451);
xnor U11744 (N_11744,N_10564,N_10787);
and U11745 (N_11745,N_10054,N_10477);
nor U11746 (N_11746,N_10953,N_10666);
nand U11747 (N_11747,N_10947,N_10080);
or U11748 (N_11748,N_10429,N_10769);
nand U11749 (N_11749,N_10434,N_10535);
nand U11750 (N_11750,N_10125,N_10311);
and U11751 (N_11751,N_10399,N_10073);
or U11752 (N_11752,N_10510,N_10847);
xor U11753 (N_11753,N_10172,N_10486);
xnor U11754 (N_11754,N_10593,N_10346);
xor U11755 (N_11755,N_10679,N_10085);
nor U11756 (N_11756,N_10641,N_10953);
nor U11757 (N_11757,N_10523,N_10952);
nand U11758 (N_11758,N_10060,N_10671);
xor U11759 (N_11759,N_10296,N_10797);
and U11760 (N_11760,N_10285,N_10972);
nand U11761 (N_11761,N_10589,N_10986);
nand U11762 (N_11762,N_10597,N_10982);
or U11763 (N_11763,N_10265,N_10562);
and U11764 (N_11764,N_10322,N_10924);
nor U11765 (N_11765,N_10090,N_10228);
nor U11766 (N_11766,N_10007,N_10766);
nand U11767 (N_11767,N_10933,N_10718);
and U11768 (N_11768,N_10336,N_10050);
xor U11769 (N_11769,N_10668,N_10850);
or U11770 (N_11770,N_10183,N_10343);
or U11771 (N_11771,N_10646,N_10072);
xor U11772 (N_11772,N_10338,N_10422);
nor U11773 (N_11773,N_10855,N_10451);
and U11774 (N_11774,N_10254,N_10920);
and U11775 (N_11775,N_10548,N_10996);
nand U11776 (N_11776,N_10412,N_10361);
nand U11777 (N_11777,N_10847,N_10591);
nor U11778 (N_11778,N_10858,N_10288);
xnor U11779 (N_11779,N_10726,N_10418);
nand U11780 (N_11780,N_10422,N_10850);
and U11781 (N_11781,N_10368,N_10828);
or U11782 (N_11782,N_10834,N_10687);
xnor U11783 (N_11783,N_10930,N_10149);
and U11784 (N_11784,N_10867,N_10344);
xor U11785 (N_11785,N_10830,N_10871);
xor U11786 (N_11786,N_10054,N_10827);
nand U11787 (N_11787,N_10679,N_10884);
or U11788 (N_11788,N_10816,N_10083);
nor U11789 (N_11789,N_10871,N_10513);
or U11790 (N_11790,N_10251,N_10827);
nand U11791 (N_11791,N_10941,N_10465);
xor U11792 (N_11792,N_10336,N_10100);
and U11793 (N_11793,N_10715,N_10435);
or U11794 (N_11794,N_10186,N_10611);
or U11795 (N_11795,N_10737,N_10336);
or U11796 (N_11796,N_10379,N_10911);
or U11797 (N_11797,N_10708,N_10247);
nand U11798 (N_11798,N_10790,N_10409);
nand U11799 (N_11799,N_10565,N_10850);
or U11800 (N_11800,N_10031,N_10891);
and U11801 (N_11801,N_10205,N_10347);
and U11802 (N_11802,N_10127,N_10643);
or U11803 (N_11803,N_10952,N_10777);
nor U11804 (N_11804,N_10222,N_10353);
nand U11805 (N_11805,N_10010,N_10394);
and U11806 (N_11806,N_10105,N_10668);
or U11807 (N_11807,N_10417,N_10938);
and U11808 (N_11808,N_10058,N_10115);
xnor U11809 (N_11809,N_10177,N_10182);
xnor U11810 (N_11810,N_10311,N_10536);
and U11811 (N_11811,N_10259,N_10528);
or U11812 (N_11812,N_10382,N_10023);
nand U11813 (N_11813,N_10005,N_10899);
and U11814 (N_11814,N_10327,N_10130);
or U11815 (N_11815,N_10337,N_10728);
and U11816 (N_11816,N_10682,N_10079);
nor U11817 (N_11817,N_10532,N_10655);
or U11818 (N_11818,N_10673,N_10109);
and U11819 (N_11819,N_10887,N_10132);
nor U11820 (N_11820,N_10345,N_10346);
or U11821 (N_11821,N_10941,N_10502);
and U11822 (N_11822,N_10162,N_10864);
xnor U11823 (N_11823,N_10150,N_10655);
or U11824 (N_11824,N_10597,N_10873);
or U11825 (N_11825,N_10754,N_10117);
nand U11826 (N_11826,N_10988,N_10412);
or U11827 (N_11827,N_10360,N_10376);
nand U11828 (N_11828,N_10945,N_10868);
nor U11829 (N_11829,N_10117,N_10099);
xnor U11830 (N_11830,N_10885,N_10602);
xor U11831 (N_11831,N_10337,N_10197);
and U11832 (N_11832,N_10748,N_10083);
and U11833 (N_11833,N_10890,N_10879);
or U11834 (N_11834,N_10381,N_10458);
nor U11835 (N_11835,N_10931,N_10354);
nor U11836 (N_11836,N_10958,N_10350);
xor U11837 (N_11837,N_10115,N_10695);
nor U11838 (N_11838,N_10987,N_10542);
or U11839 (N_11839,N_10812,N_10565);
or U11840 (N_11840,N_10256,N_10348);
and U11841 (N_11841,N_10270,N_10618);
or U11842 (N_11842,N_10929,N_10174);
nand U11843 (N_11843,N_10801,N_10309);
or U11844 (N_11844,N_10976,N_10606);
nor U11845 (N_11845,N_10595,N_10977);
and U11846 (N_11846,N_10157,N_10873);
or U11847 (N_11847,N_10857,N_10444);
or U11848 (N_11848,N_10045,N_10177);
or U11849 (N_11849,N_10472,N_10148);
and U11850 (N_11850,N_10868,N_10985);
nor U11851 (N_11851,N_10639,N_10348);
and U11852 (N_11852,N_10424,N_10015);
and U11853 (N_11853,N_10730,N_10958);
and U11854 (N_11854,N_10573,N_10125);
nor U11855 (N_11855,N_10718,N_10802);
nand U11856 (N_11856,N_10048,N_10579);
nor U11857 (N_11857,N_10985,N_10318);
and U11858 (N_11858,N_10977,N_10536);
xor U11859 (N_11859,N_10916,N_10993);
and U11860 (N_11860,N_10924,N_10196);
and U11861 (N_11861,N_10992,N_10330);
nor U11862 (N_11862,N_10944,N_10729);
or U11863 (N_11863,N_10804,N_10289);
nand U11864 (N_11864,N_10467,N_10145);
xnor U11865 (N_11865,N_10498,N_10339);
nand U11866 (N_11866,N_10290,N_10819);
and U11867 (N_11867,N_10804,N_10626);
and U11868 (N_11868,N_10804,N_10914);
nand U11869 (N_11869,N_10319,N_10627);
and U11870 (N_11870,N_10699,N_10843);
xnor U11871 (N_11871,N_10231,N_10676);
and U11872 (N_11872,N_10707,N_10213);
xnor U11873 (N_11873,N_10564,N_10118);
nand U11874 (N_11874,N_10828,N_10542);
or U11875 (N_11875,N_10979,N_10092);
nand U11876 (N_11876,N_10865,N_10693);
and U11877 (N_11877,N_10954,N_10731);
xnor U11878 (N_11878,N_10528,N_10763);
nor U11879 (N_11879,N_10043,N_10926);
xor U11880 (N_11880,N_10999,N_10034);
and U11881 (N_11881,N_10905,N_10372);
nand U11882 (N_11882,N_10091,N_10967);
xor U11883 (N_11883,N_10364,N_10208);
nand U11884 (N_11884,N_10132,N_10499);
and U11885 (N_11885,N_10885,N_10772);
and U11886 (N_11886,N_10391,N_10903);
or U11887 (N_11887,N_10455,N_10174);
or U11888 (N_11888,N_10799,N_10341);
nor U11889 (N_11889,N_10978,N_10781);
nor U11890 (N_11890,N_10797,N_10996);
xor U11891 (N_11891,N_10883,N_10593);
or U11892 (N_11892,N_10016,N_10408);
nand U11893 (N_11893,N_10801,N_10739);
nor U11894 (N_11894,N_10331,N_10581);
nand U11895 (N_11895,N_10688,N_10365);
xnor U11896 (N_11896,N_10431,N_10250);
nand U11897 (N_11897,N_10900,N_10690);
nor U11898 (N_11898,N_10778,N_10902);
xor U11899 (N_11899,N_10786,N_10616);
and U11900 (N_11900,N_10880,N_10204);
nor U11901 (N_11901,N_10298,N_10511);
nor U11902 (N_11902,N_10213,N_10727);
nor U11903 (N_11903,N_10489,N_10016);
nor U11904 (N_11904,N_10914,N_10115);
or U11905 (N_11905,N_10598,N_10951);
nand U11906 (N_11906,N_10128,N_10489);
nor U11907 (N_11907,N_10998,N_10462);
nand U11908 (N_11908,N_10265,N_10332);
nor U11909 (N_11909,N_10057,N_10904);
nand U11910 (N_11910,N_10647,N_10947);
nor U11911 (N_11911,N_10397,N_10861);
nor U11912 (N_11912,N_10858,N_10761);
and U11913 (N_11913,N_10753,N_10810);
or U11914 (N_11914,N_10492,N_10936);
or U11915 (N_11915,N_10806,N_10895);
or U11916 (N_11916,N_10466,N_10841);
nand U11917 (N_11917,N_10017,N_10785);
or U11918 (N_11918,N_10384,N_10165);
xor U11919 (N_11919,N_10014,N_10109);
or U11920 (N_11920,N_10028,N_10905);
nor U11921 (N_11921,N_10587,N_10554);
nor U11922 (N_11922,N_10013,N_10701);
and U11923 (N_11923,N_10438,N_10956);
and U11924 (N_11924,N_10594,N_10760);
and U11925 (N_11925,N_10905,N_10690);
nand U11926 (N_11926,N_10045,N_10505);
nand U11927 (N_11927,N_10122,N_10128);
xnor U11928 (N_11928,N_10374,N_10735);
and U11929 (N_11929,N_10164,N_10435);
or U11930 (N_11930,N_10299,N_10016);
or U11931 (N_11931,N_10611,N_10010);
or U11932 (N_11932,N_10149,N_10618);
and U11933 (N_11933,N_10562,N_10437);
nand U11934 (N_11934,N_10761,N_10699);
and U11935 (N_11935,N_10766,N_10291);
nand U11936 (N_11936,N_10268,N_10399);
or U11937 (N_11937,N_10064,N_10398);
xor U11938 (N_11938,N_10791,N_10349);
or U11939 (N_11939,N_10311,N_10034);
nand U11940 (N_11940,N_10486,N_10523);
xnor U11941 (N_11941,N_10050,N_10769);
or U11942 (N_11942,N_10769,N_10586);
and U11943 (N_11943,N_10457,N_10622);
nor U11944 (N_11944,N_10389,N_10941);
or U11945 (N_11945,N_10447,N_10947);
or U11946 (N_11946,N_10459,N_10956);
xnor U11947 (N_11947,N_10586,N_10049);
nor U11948 (N_11948,N_10965,N_10248);
xor U11949 (N_11949,N_10227,N_10427);
xnor U11950 (N_11950,N_10096,N_10230);
nor U11951 (N_11951,N_10375,N_10596);
nand U11952 (N_11952,N_10187,N_10721);
nand U11953 (N_11953,N_10632,N_10605);
nor U11954 (N_11954,N_10526,N_10568);
and U11955 (N_11955,N_10954,N_10155);
nor U11956 (N_11956,N_10821,N_10766);
nand U11957 (N_11957,N_10227,N_10223);
or U11958 (N_11958,N_10843,N_10671);
nor U11959 (N_11959,N_10817,N_10944);
nand U11960 (N_11960,N_10795,N_10228);
xnor U11961 (N_11961,N_10085,N_10939);
nor U11962 (N_11962,N_10399,N_10229);
or U11963 (N_11963,N_10274,N_10029);
and U11964 (N_11964,N_10755,N_10763);
and U11965 (N_11965,N_10044,N_10623);
nor U11966 (N_11966,N_10899,N_10321);
nor U11967 (N_11967,N_10358,N_10907);
xnor U11968 (N_11968,N_10449,N_10952);
xnor U11969 (N_11969,N_10642,N_10312);
and U11970 (N_11970,N_10410,N_10267);
nor U11971 (N_11971,N_10445,N_10885);
nor U11972 (N_11972,N_10927,N_10942);
or U11973 (N_11973,N_10120,N_10915);
xor U11974 (N_11974,N_10236,N_10587);
and U11975 (N_11975,N_10894,N_10749);
and U11976 (N_11976,N_10421,N_10481);
and U11977 (N_11977,N_10565,N_10708);
or U11978 (N_11978,N_10745,N_10059);
or U11979 (N_11979,N_10465,N_10840);
and U11980 (N_11980,N_10803,N_10071);
nor U11981 (N_11981,N_10904,N_10538);
and U11982 (N_11982,N_10333,N_10673);
xor U11983 (N_11983,N_10429,N_10758);
and U11984 (N_11984,N_10914,N_10543);
and U11985 (N_11985,N_10921,N_10171);
nand U11986 (N_11986,N_10758,N_10632);
xnor U11987 (N_11987,N_10603,N_10639);
xor U11988 (N_11988,N_10648,N_10100);
nor U11989 (N_11989,N_10519,N_10728);
or U11990 (N_11990,N_10398,N_10728);
and U11991 (N_11991,N_10004,N_10123);
nor U11992 (N_11992,N_10310,N_10725);
or U11993 (N_11993,N_10171,N_10585);
nand U11994 (N_11994,N_10078,N_10692);
or U11995 (N_11995,N_10908,N_10627);
nand U11996 (N_11996,N_10552,N_10143);
nand U11997 (N_11997,N_10934,N_10147);
xnor U11998 (N_11998,N_10818,N_10244);
xor U11999 (N_11999,N_10163,N_10970);
or U12000 (N_12000,N_11904,N_11396);
nand U12001 (N_12001,N_11392,N_11019);
nor U12002 (N_12002,N_11277,N_11365);
xor U12003 (N_12003,N_11841,N_11423);
nand U12004 (N_12004,N_11501,N_11881);
xnor U12005 (N_12005,N_11370,N_11249);
xnor U12006 (N_12006,N_11749,N_11390);
or U12007 (N_12007,N_11140,N_11728);
xor U12008 (N_12008,N_11522,N_11516);
nor U12009 (N_12009,N_11264,N_11210);
nor U12010 (N_12010,N_11422,N_11435);
nor U12011 (N_12011,N_11513,N_11860);
or U12012 (N_12012,N_11171,N_11156);
nand U12013 (N_12013,N_11052,N_11153);
and U12014 (N_12014,N_11934,N_11341);
nor U12015 (N_12015,N_11371,N_11295);
and U12016 (N_12016,N_11291,N_11543);
nand U12017 (N_12017,N_11544,N_11023);
nor U12018 (N_12018,N_11048,N_11686);
nand U12019 (N_12019,N_11761,N_11968);
and U12020 (N_12020,N_11481,N_11046);
or U12021 (N_12021,N_11692,N_11244);
nand U12022 (N_12022,N_11381,N_11322);
or U12023 (N_12023,N_11476,N_11213);
and U12024 (N_12024,N_11228,N_11755);
and U12025 (N_12025,N_11503,N_11983);
nand U12026 (N_12026,N_11980,N_11175);
nor U12027 (N_12027,N_11671,N_11633);
xnor U12028 (N_12028,N_11094,N_11553);
nor U12029 (N_12029,N_11283,N_11606);
or U12030 (N_12030,N_11074,N_11225);
nor U12031 (N_12031,N_11152,N_11824);
and U12032 (N_12032,N_11650,N_11573);
or U12033 (N_12033,N_11147,N_11697);
or U12034 (N_12034,N_11710,N_11206);
and U12035 (N_12035,N_11644,N_11666);
nand U12036 (N_12036,N_11621,N_11623);
nand U12037 (N_12037,N_11729,N_11781);
nand U12038 (N_12038,N_11072,N_11012);
or U12039 (N_12039,N_11131,N_11431);
and U12040 (N_12040,N_11694,N_11866);
xor U12041 (N_12041,N_11955,N_11412);
or U12042 (N_12042,N_11090,N_11745);
xor U12043 (N_12043,N_11065,N_11886);
xnor U12044 (N_12044,N_11461,N_11652);
nand U12045 (N_12045,N_11071,N_11007);
xor U12046 (N_12046,N_11184,N_11062);
nor U12047 (N_12047,N_11816,N_11843);
and U12048 (N_12048,N_11819,N_11995);
xor U12049 (N_12049,N_11488,N_11174);
or U12050 (N_12050,N_11654,N_11948);
xnor U12051 (N_12051,N_11681,N_11827);
xnor U12052 (N_12052,N_11580,N_11750);
and U12053 (N_12053,N_11105,N_11526);
and U12054 (N_12054,N_11849,N_11159);
and U12055 (N_12055,N_11639,N_11077);
or U12056 (N_12056,N_11957,N_11196);
nand U12057 (N_12057,N_11847,N_11844);
nand U12058 (N_12058,N_11601,N_11890);
nand U12059 (N_12059,N_11818,N_11255);
nand U12060 (N_12060,N_11906,N_11135);
xnor U12061 (N_12061,N_11429,N_11495);
and U12062 (N_12062,N_11375,N_11776);
nand U12063 (N_12063,N_11059,N_11055);
or U12064 (N_12064,N_11106,N_11610);
xor U12065 (N_12065,N_11188,N_11253);
xor U12066 (N_12066,N_11937,N_11293);
nand U12067 (N_12067,N_11638,N_11514);
nor U12068 (N_12068,N_11970,N_11212);
nand U12069 (N_12069,N_11701,N_11192);
nor U12070 (N_12070,N_11604,N_11400);
xnor U12071 (N_12071,N_11076,N_11383);
xor U12072 (N_12072,N_11663,N_11767);
or U12073 (N_12073,N_11418,N_11913);
nor U12074 (N_12074,N_11411,N_11700);
and U12075 (N_12075,N_11347,N_11587);
nand U12076 (N_12076,N_11098,N_11765);
nand U12077 (N_12077,N_11442,N_11630);
nand U12078 (N_12078,N_11768,N_11256);
nand U12079 (N_12079,N_11441,N_11737);
and U12080 (N_12080,N_11067,N_11005);
or U12081 (N_12081,N_11891,N_11466);
or U12082 (N_12082,N_11304,N_11313);
or U12083 (N_12083,N_11204,N_11637);
or U12084 (N_12084,N_11545,N_11393);
nor U12085 (N_12085,N_11112,N_11326);
nand U12086 (N_12086,N_11763,N_11292);
and U12087 (N_12087,N_11812,N_11199);
or U12088 (N_12088,N_11714,N_11143);
nand U12089 (N_12089,N_11389,N_11925);
xnor U12090 (N_12090,N_11817,N_11532);
and U12091 (N_12091,N_11363,N_11811);
xnor U12092 (N_12092,N_11667,N_11507);
or U12093 (N_12093,N_11519,N_11099);
or U12094 (N_12094,N_11864,N_11360);
and U12095 (N_12095,N_11732,N_11372);
nand U12096 (N_12096,N_11270,N_11856);
and U12097 (N_12097,N_11111,N_11884);
nor U12098 (N_12098,N_11661,N_11744);
nor U12099 (N_12099,N_11003,N_11069);
nand U12100 (N_12100,N_11051,N_11807);
nand U12101 (N_12101,N_11879,N_11454);
nor U12102 (N_12102,N_11629,N_11136);
xor U12103 (N_12103,N_11785,N_11677);
nor U12104 (N_12104,N_11848,N_11956);
nand U12105 (N_12105,N_11774,N_11992);
and U12106 (N_12106,N_11551,N_11464);
xor U12107 (N_12107,N_11696,N_11274);
nor U12108 (N_12108,N_11352,N_11434);
nand U12109 (N_12109,N_11234,N_11288);
or U12110 (N_12110,N_11335,N_11539);
xnor U12111 (N_12111,N_11218,N_11096);
or U12112 (N_12112,N_11440,N_11875);
nor U12113 (N_12113,N_11182,N_11222);
xor U12114 (N_12114,N_11374,N_11211);
or U12115 (N_12115,N_11521,N_11822);
or U12116 (N_12116,N_11149,N_11989);
nor U12117 (N_12117,N_11399,N_11655);
xor U12118 (N_12118,N_11057,N_11808);
nand U12119 (N_12119,N_11905,N_11323);
and U12120 (N_12120,N_11286,N_11971);
nand U12121 (N_12121,N_11706,N_11780);
and U12122 (N_12122,N_11660,N_11517);
xnor U12123 (N_12123,N_11320,N_11004);
xnor U12124 (N_12124,N_11518,N_11314);
nand U12125 (N_12125,N_11034,N_11718);
nand U12126 (N_12126,N_11345,N_11452);
nor U12127 (N_12127,N_11089,N_11586);
and U12128 (N_12128,N_11416,N_11474);
nand U12129 (N_12129,N_11297,N_11746);
xnor U12130 (N_12130,N_11275,N_11061);
nor U12131 (N_12131,N_11085,N_11520);
nor U12132 (N_12132,N_11132,N_11611);
nand U12133 (N_12133,N_11547,N_11317);
nor U12134 (N_12134,N_11598,N_11427);
and U12135 (N_12135,N_11252,N_11803);
xnor U12136 (N_12136,N_11865,N_11709);
xnor U12137 (N_12137,N_11670,N_11590);
or U12138 (N_12138,N_11082,N_11945);
nand U12139 (N_12139,N_11355,N_11397);
xor U12140 (N_12140,N_11603,N_11350);
nor U12141 (N_12141,N_11877,N_11569);
nand U12142 (N_12142,N_11908,N_11845);
xnor U12143 (N_12143,N_11432,N_11962);
xor U12144 (N_12144,N_11013,N_11723);
nand U12145 (N_12145,N_11353,N_11494);
nor U12146 (N_12146,N_11585,N_11713);
and U12147 (N_12147,N_11280,N_11373);
nand U12148 (N_12148,N_11279,N_11402);
nand U12149 (N_12149,N_11009,N_11973);
or U12150 (N_12150,N_11535,N_11690);
or U12151 (N_12151,N_11794,N_11006);
nand U12152 (N_12152,N_11473,N_11640);
nand U12153 (N_12153,N_11678,N_11820);
or U12154 (N_12154,N_11505,N_11008);
or U12155 (N_12155,N_11066,N_11240);
nor U12156 (N_12156,N_11760,N_11506);
or U12157 (N_12157,N_11570,N_11348);
or U12158 (N_12158,N_11556,N_11648);
or U12159 (N_12159,N_11359,N_11364);
xor U12160 (N_12160,N_11385,N_11682);
nor U12161 (N_12161,N_11200,N_11762);
and U12162 (N_12162,N_11231,N_11462);
nor U12163 (N_12163,N_11510,N_11748);
nand U12164 (N_12164,N_11950,N_11178);
and U12165 (N_12165,N_11530,N_11772);
xnor U12166 (N_12166,N_11444,N_11001);
xor U12167 (N_12167,N_11308,N_11162);
nand U12168 (N_12168,N_11540,N_11405);
and U12169 (N_12169,N_11502,N_11436);
or U12170 (N_12170,N_11991,N_11617);
nor U12171 (N_12171,N_11080,N_11467);
xor U12172 (N_12172,N_11997,N_11753);
xor U12173 (N_12173,N_11026,N_11565);
nor U12174 (N_12174,N_11888,N_11882);
or U12175 (N_12175,N_11276,N_11528);
and U12176 (N_12176,N_11407,N_11340);
and U12177 (N_12177,N_11806,N_11979);
xnor U12178 (N_12178,N_11672,N_11408);
xnor U12179 (N_12179,N_11025,N_11311);
or U12180 (N_12180,N_11500,N_11107);
xnor U12181 (N_12181,N_11898,N_11215);
or U12182 (N_12182,N_11475,N_11959);
and U12183 (N_12183,N_11887,N_11766);
nand U12184 (N_12184,N_11897,N_11302);
nor U12185 (N_12185,N_11870,N_11717);
xnor U12186 (N_12186,N_11593,N_11041);
nor U12187 (N_12187,N_11227,N_11736);
or U12188 (N_12188,N_11837,N_11727);
xnor U12189 (N_12189,N_11421,N_11493);
and U12190 (N_12190,N_11413,N_11840);
nand U12191 (N_12191,N_11477,N_11688);
and U12192 (N_12192,N_11981,N_11949);
xnor U12193 (N_12193,N_11424,N_11160);
nor U12194 (N_12194,N_11202,N_11627);
nand U12195 (N_12195,N_11896,N_11928);
nor U12196 (N_12196,N_11060,N_11047);
and U12197 (N_12197,N_11480,N_11880);
nor U12198 (N_12198,N_11636,N_11299);
and U12199 (N_12199,N_11243,N_11619);
or U12200 (N_12200,N_11775,N_11595);
nor U12201 (N_12201,N_11779,N_11095);
xor U12202 (N_12202,N_11926,N_11635);
nand U12203 (N_12203,N_11977,N_11027);
xor U12204 (N_12204,N_11582,N_11369);
nand U12205 (N_12205,N_11226,N_11922);
xnor U12206 (N_12206,N_11662,N_11120);
nand U12207 (N_12207,N_11576,N_11419);
and U12208 (N_12208,N_11835,N_11091);
nor U12209 (N_12209,N_11558,N_11310);
xor U12210 (N_12210,N_11002,N_11319);
or U12211 (N_12211,N_11523,N_11771);
xor U12212 (N_12212,N_11271,N_11911);
and U12213 (N_12213,N_11910,N_11932);
and U12214 (N_12214,N_11119,N_11457);
and U12215 (N_12215,N_11037,N_11715);
xor U12216 (N_12216,N_11260,N_11491);
and U12217 (N_12217,N_11205,N_11823);
xnor U12218 (N_12218,N_11658,N_11919);
nand U12219 (N_12219,N_11221,N_11078);
nor U12220 (N_12220,N_11784,N_11267);
nor U12221 (N_12221,N_11613,N_11600);
nand U12222 (N_12222,N_11577,N_11914);
xnor U12223 (N_12223,N_11883,N_11108);
nor U12224 (N_12224,N_11263,N_11698);
nor U12225 (N_12225,N_11043,N_11938);
nor U12226 (N_12226,N_11975,N_11834);
or U12227 (N_12227,N_11233,N_11097);
or U12228 (N_12228,N_11010,N_11687);
or U12229 (N_12229,N_11838,N_11954);
nor U12230 (N_12230,N_11562,N_11764);
or U12231 (N_12231,N_11022,N_11490);
xor U12232 (N_12232,N_11425,N_11958);
or U12233 (N_12233,N_11825,N_11557);
nand U12234 (N_12234,N_11689,N_11306);
nor U12235 (N_12235,N_11575,N_11708);
or U12236 (N_12236,N_11318,N_11414);
nor U12237 (N_12237,N_11315,N_11596);
nand U12238 (N_12238,N_11088,N_11028);
nand U12239 (N_12239,N_11974,N_11376);
xor U12240 (N_12240,N_11861,N_11965);
nor U12241 (N_12241,N_11073,N_11115);
xnor U12242 (N_12242,N_11272,N_11739);
xor U12243 (N_12243,N_11668,N_11449);
or U12244 (N_12244,N_11081,N_11567);
and U12245 (N_12245,N_11641,N_11921);
nand U12246 (N_12246,N_11216,N_11117);
nor U12247 (N_12247,N_11550,N_11170);
and U12248 (N_12248,N_11038,N_11130);
or U12249 (N_12249,N_11391,N_11792);
and U12250 (N_12250,N_11525,N_11529);
and U12251 (N_12251,N_11536,N_11871);
nand U12252 (N_12252,N_11448,N_11238);
nor U12253 (N_12253,N_11857,N_11118);
nand U12254 (N_12254,N_11999,N_11332);
nand U12255 (N_12255,N_11730,N_11832);
or U12256 (N_12256,N_11181,N_11207);
or U12257 (N_12257,N_11087,N_11742);
nor U12258 (N_12258,N_11931,N_11325);
nand U12259 (N_12259,N_11907,N_11947);
xor U12260 (N_12260,N_11472,N_11484);
nor U12261 (N_12261,N_11952,N_11588);
or U12262 (N_12262,N_11103,N_11125);
or U12263 (N_12263,N_11770,N_11581);
nor U12264 (N_12264,N_11235,N_11296);
nor U12265 (N_12265,N_11334,N_11802);
nor U12266 (N_12266,N_11796,N_11453);
nand U12267 (N_12267,N_11936,N_11224);
xnor U12268 (N_12268,N_11612,N_11508);
nor U12269 (N_12269,N_11996,N_11161);
nor U12270 (N_12270,N_11266,N_11036);
or U12271 (N_12271,N_11110,N_11799);
or U12272 (N_12272,N_11011,N_11787);
nand U12273 (N_12273,N_11994,N_11592);
nand U12274 (N_12274,N_11858,N_11646);
nor U12275 (N_12275,N_11607,N_11721);
or U12276 (N_12276,N_11560,N_11554);
xnor U12277 (N_12277,N_11342,N_11281);
or U12278 (N_12278,N_11786,N_11380);
or U12279 (N_12279,N_11574,N_11123);
xor U12280 (N_12280,N_11836,N_11109);
xor U12281 (N_12281,N_11614,N_11659);
and U12282 (N_12282,N_11814,N_11647);
nor U12283 (N_12283,N_11972,N_11797);
and U12284 (N_12284,N_11031,N_11683);
and U12285 (N_12285,N_11138,N_11236);
and U12286 (N_12286,N_11489,N_11093);
nor U12287 (N_12287,N_11116,N_11417);
nand U12288 (N_12288,N_11564,N_11289);
nand U12289 (N_12289,N_11458,N_11428);
and U12290 (N_12290,N_11021,N_11433);
nor U12291 (N_12291,N_11839,N_11833);
nor U12292 (N_12292,N_11790,N_11531);
nand U12293 (N_12293,N_11214,N_11220);
nor U12294 (N_12294,N_11312,N_11862);
nand U12295 (N_12295,N_11743,N_11899);
and U12296 (N_12296,N_11773,N_11893);
nand U12297 (N_12297,N_11450,N_11533);
xor U12298 (N_12298,N_11854,N_11190);
and U12299 (N_12299,N_11944,N_11079);
nand U12300 (N_12300,N_11704,N_11316);
and U12301 (N_12301,N_11113,N_11969);
or U12302 (N_12302,N_11851,N_11933);
or U12303 (N_12303,N_11254,N_11685);
xnor U12304 (N_12304,N_11759,N_11791);
nand U12305 (N_12305,N_11201,N_11900);
nor U12306 (N_12306,N_11157,N_11331);
nand U12307 (N_12307,N_11684,N_11702);
or U12308 (N_12308,N_11859,N_11250);
nor U12309 (N_12309,N_11483,N_11426);
xor U12310 (N_12310,N_11869,N_11287);
nand U12311 (N_12311,N_11187,N_11795);
xor U12312 (N_12312,N_11404,N_11628);
and U12313 (N_12313,N_11083,N_11198);
nor U12314 (N_12314,N_11141,N_11720);
nand U12315 (N_12315,N_11127,N_11946);
xnor U12316 (N_12316,N_11468,N_11626);
nor U12317 (N_12317,N_11942,N_11406);
and U12318 (N_12318,N_11189,N_11245);
nand U12319 (N_12319,N_11014,N_11145);
nand U12320 (N_12320,N_11534,N_11804);
nor U12321 (N_12321,N_11142,N_11665);
nor U12322 (N_12322,N_11030,N_11387);
nand U12323 (N_12323,N_11492,N_11978);
nor U12324 (N_12324,N_11185,N_11165);
and U12325 (N_12325,N_11752,N_11191);
and U12326 (N_12326,N_11622,N_11219);
and U12327 (N_12327,N_11039,N_11456);
and U12328 (N_12328,N_11268,N_11121);
or U12329 (N_12329,N_11563,N_11487);
or U12330 (N_12330,N_11339,N_11368);
or U12331 (N_12331,N_11699,N_11015);
or U12332 (N_12332,N_11179,N_11571);
or U12333 (N_12333,N_11265,N_11258);
or U12334 (N_12334,N_11032,N_11168);
nand U12335 (N_12335,N_11054,N_11033);
nor U12336 (N_12336,N_11769,N_11976);
or U12337 (N_12337,N_11470,N_11800);
xnor U12338 (N_12338,N_11197,N_11597);
xor U12339 (N_12339,N_11566,N_11757);
nor U12340 (N_12340,N_11894,N_11482);
nor U12341 (N_12341,N_11608,N_11478);
xnor U12342 (N_12342,N_11620,N_11902);
nor U12343 (N_12343,N_11209,N_11583);
and U12344 (N_12344,N_11122,N_11469);
nor U12345 (N_12345,N_11830,N_11541);
nor U12346 (N_12346,N_11068,N_11084);
or U12347 (N_12347,N_11850,N_11398);
or U12348 (N_12348,N_11045,N_11324);
nor U12349 (N_12349,N_11777,N_11632);
nor U12350 (N_12350,N_11337,N_11552);
and U12351 (N_12351,N_11208,N_11829);
or U12352 (N_12352,N_11878,N_11180);
and U12353 (N_12353,N_11446,N_11711);
or U12354 (N_12354,N_11016,N_11303);
xor U12355 (N_12355,N_11437,N_11656);
nor U12356 (N_12356,N_11605,N_11951);
xnor U12357 (N_12357,N_11512,N_11333);
xor U12358 (N_12358,N_11537,N_11943);
nor U12359 (N_12359,N_11726,N_11579);
or U12360 (N_12360,N_11895,N_11939);
nor U12361 (N_12361,N_11146,N_11674);
and U12362 (N_12362,N_11964,N_11863);
or U12363 (N_12363,N_11195,N_11307);
or U12364 (N_12364,N_11327,N_11247);
nor U12365 (N_12365,N_11029,N_11504);
or U12366 (N_12366,N_11042,N_11993);
nand U12367 (N_12367,N_11044,N_11460);
nor U12368 (N_12368,N_11070,N_11542);
nor U12369 (N_12369,N_11357,N_11852);
and U12370 (N_12370,N_11193,N_11309);
nand U12371 (N_12371,N_11987,N_11889);
and U12372 (N_12372,N_11163,N_11259);
or U12373 (N_12373,N_11438,N_11568);
nor U12374 (N_12374,N_11058,N_11150);
xor U12375 (N_12375,N_11751,N_11024);
xnor U12376 (N_12376,N_11035,N_11986);
nor U12377 (N_12377,N_11395,N_11548);
xor U12378 (N_12378,N_11716,N_11915);
and U12379 (N_12379,N_11966,N_11624);
nand U12380 (N_12380,N_11415,N_11876);
nand U12381 (N_12381,N_11410,N_11102);
or U12382 (N_12382,N_11695,N_11378);
and U12383 (N_12383,N_11124,N_11705);
xnor U12384 (N_12384,N_11733,N_11599);
and U12385 (N_12385,N_11329,N_11524);
and U12386 (N_12386,N_11305,N_11230);
nor U12387 (N_12387,N_11909,N_11798);
nand U12388 (N_12388,N_11384,N_11455);
nand U12389 (N_12389,N_11086,N_11128);
or U12390 (N_12390,N_11155,N_11050);
and U12391 (N_12391,N_11868,N_11712);
nand U12392 (N_12392,N_11676,N_11758);
or U12393 (N_12393,N_11815,N_11126);
or U12394 (N_12394,N_11953,N_11903);
xor U12395 (N_12395,N_11923,N_11242);
or U12396 (N_12396,N_11912,N_11101);
and U12397 (N_12397,N_11885,N_11379);
and U12398 (N_12398,N_11782,N_11167);
nand U12399 (N_12399,N_11831,N_11420);
nand U12400 (N_12400,N_11445,N_11982);
and U12401 (N_12401,N_11778,N_11801);
nand U12402 (N_12402,N_11874,N_11217);
nand U12403 (N_12403,N_11176,N_11669);
xnor U12404 (N_12404,N_11394,N_11064);
nor U12405 (N_12405,N_11338,N_11929);
and U12406 (N_12406,N_11328,N_11261);
nand U12407 (N_12407,N_11589,N_11194);
nand U12408 (N_12408,N_11559,N_11485);
or U12409 (N_12409,N_11988,N_11754);
xor U12410 (N_12410,N_11443,N_11591);
nor U12411 (N_12411,N_11645,N_11618);
nand U12412 (N_12412,N_11336,N_11251);
and U12413 (N_12413,N_11354,N_11499);
nor U12414 (N_12414,N_11056,N_11134);
nor U12415 (N_12415,N_11680,N_11651);
nand U12416 (N_12416,N_11092,N_11967);
nor U12417 (N_12417,N_11821,N_11223);
xnor U12418 (N_12418,N_11901,N_11382);
nand U12419 (N_12419,N_11386,N_11430);
xnor U12420 (N_12420,N_11738,N_11463);
or U12421 (N_12421,N_11990,N_11451);
nor U12422 (N_12422,N_11649,N_11151);
nor U12423 (N_12423,N_11330,N_11740);
nor U12424 (N_12424,N_11924,N_11248);
and U12425 (N_12425,N_11731,N_11496);
or U12426 (N_12426,N_11344,N_11960);
and U12427 (N_12427,N_11285,N_11805);
and U12428 (N_12428,N_11961,N_11351);
nand U12429 (N_12429,N_11810,N_11789);
and U12430 (N_12430,N_11144,N_11000);
or U12431 (N_12431,N_11063,N_11643);
nor U12432 (N_12432,N_11040,N_11447);
and U12433 (N_12433,N_11515,N_11918);
xor U12434 (N_12434,N_11498,N_11439);
nor U12435 (N_12435,N_11657,N_11246);
xor U12436 (N_12436,N_11538,N_11783);
nor U12437 (N_12437,N_11735,N_11154);
or U12438 (N_12438,N_11239,N_11177);
nor U12439 (N_12439,N_11625,N_11602);
nand U12440 (N_12440,N_11927,N_11020);
nand U12441 (N_12441,N_11358,N_11693);
nor U12442 (N_12442,N_11139,N_11935);
nor U12443 (N_12443,N_11941,N_11133);
and U12444 (N_12444,N_11963,N_11017);
and U12445 (N_12445,N_11471,N_11367);
and U12446 (N_12446,N_11300,N_11561);
xor U12447 (N_12447,N_11719,N_11294);
nor U12448 (N_12448,N_11703,N_11409);
and U12449 (N_12449,N_11486,N_11511);
nand U12450 (N_12450,N_11616,N_11826);
nor U12451 (N_12451,N_11609,N_11675);
xor U12452 (N_12452,N_11346,N_11572);
or U12453 (N_12453,N_11388,N_11366);
nor U12454 (N_12454,N_11349,N_11241);
and U12455 (N_12455,N_11053,N_11497);
or U12456 (N_12456,N_11229,N_11075);
and U12457 (N_12457,N_11377,N_11361);
nor U12458 (N_12458,N_11273,N_11828);
xnor U12459 (N_12459,N_11724,N_11916);
and U12460 (N_12460,N_11257,N_11892);
nor U12461 (N_12461,N_11756,N_11853);
or U12462 (N_12462,N_11104,N_11984);
xor U12463 (N_12463,N_11290,N_11940);
nand U12464 (N_12464,N_11114,N_11403);
nor U12465 (N_12465,N_11362,N_11809);
and U12466 (N_12466,N_11148,N_11164);
xor U12467 (N_12467,N_11584,N_11998);
or U12468 (N_12468,N_11278,N_11269);
or U12469 (N_12469,N_11401,N_11343);
nor U12470 (N_12470,N_11166,N_11100);
xnor U12471 (N_12471,N_11262,N_11747);
and U12472 (N_12472,N_11846,N_11734);
xor U12473 (N_12473,N_11555,N_11129);
nor U12474 (N_12474,N_11183,N_11203);
or U12475 (N_12475,N_11642,N_11594);
and U12476 (N_12476,N_11298,N_11546);
and U12477 (N_12477,N_11186,N_11578);
or U12478 (N_12478,N_11527,N_11930);
nand U12479 (N_12479,N_11172,N_11301);
or U12480 (N_12480,N_11232,N_11725);
and U12481 (N_12481,N_11985,N_11158);
and U12482 (N_12482,N_11788,N_11169);
nor U12483 (N_12483,N_11634,N_11867);
nor U12484 (N_12484,N_11855,N_11679);
xor U12485 (N_12485,N_11631,N_11653);
nand U12486 (N_12486,N_11741,N_11793);
xnor U12487 (N_12487,N_11673,N_11479);
nor U12488 (N_12488,N_11237,N_11284);
xnor U12489 (N_12489,N_11018,N_11873);
and U12490 (N_12490,N_11664,N_11920);
nand U12491 (N_12491,N_11465,N_11282);
or U12492 (N_12492,N_11321,N_11917);
nor U12493 (N_12493,N_11356,N_11722);
xor U12494 (N_12494,N_11459,N_11615);
nand U12495 (N_12495,N_11691,N_11173);
and U12496 (N_12496,N_11813,N_11872);
xor U12497 (N_12497,N_11549,N_11707);
or U12498 (N_12498,N_11509,N_11049);
or U12499 (N_12499,N_11137,N_11842);
and U12500 (N_12500,N_11105,N_11326);
and U12501 (N_12501,N_11594,N_11739);
or U12502 (N_12502,N_11499,N_11494);
nand U12503 (N_12503,N_11228,N_11083);
or U12504 (N_12504,N_11632,N_11056);
nor U12505 (N_12505,N_11773,N_11916);
nand U12506 (N_12506,N_11420,N_11062);
or U12507 (N_12507,N_11737,N_11819);
nor U12508 (N_12508,N_11987,N_11717);
and U12509 (N_12509,N_11674,N_11100);
nor U12510 (N_12510,N_11087,N_11472);
nor U12511 (N_12511,N_11917,N_11682);
or U12512 (N_12512,N_11896,N_11438);
xor U12513 (N_12513,N_11880,N_11580);
xor U12514 (N_12514,N_11186,N_11369);
nand U12515 (N_12515,N_11384,N_11792);
nand U12516 (N_12516,N_11008,N_11640);
xor U12517 (N_12517,N_11596,N_11662);
xor U12518 (N_12518,N_11438,N_11457);
nor U12519 (N_12519,N_11505,N_11390);
nand U12520 (N_12520,N_11851,N_11481);
and U12521 (N_12521,N_11930,N_11170);
nand U12522 (N_12522,N_11375,N_11909);
and U12523 (N_12523,N_11003,N_11078);
nor U12524 (N_12524,N_11948,N_11594);
and U12525 (N_12525,N_11234,N_11036);
and U12526 (N_12526,N_11447,N_11307);
xnor U12527 (N_12527,N_11470,N_11022);
nand U12528 (N_12528,N_11627,N_11241);
xnor U12529 (N_12529,N_11231,N_11530);
and U12530 (N_12530,N_11953,N_11753);
nand U12531 (N_12531,N_11495,N_11207);
nand U12532 (N_12532,N_11115,N_11863);
nand U12533 (N_12533,N_11424,N_11243);
nand U12534 (N_12534,N_11974,N_11296);
or U12535 (N_12535,N_11543,N_11925);
nor U12536 (N_12536,N_11243,N_11441);
or U12537 (N_12537,N_11919,N_11105);
xor U12538 (N_12538,N_11421,N_11511);
xor U12539 (N_12539,N_11553,N_11378);
or U12540 (N_12540,N_11776,N_11479);
nand U12541 (N_12541,N_11805,N_11343);
or U12542 (N_12542,N_11096,N_11906);
xnor U12543 (N_12543,N_11717,N_11690);
nand U12544 (N_12544,N_11261,N_11436);
nand U12545 (N_12545,N_11114,N_11524);
or U12546 (N_12546,N_11164,N_11365);
xor U12547 (N_12547,N_11846,N_11943);
xnor U12548 (N_12548,N_11859,N_11875);
xnor U12549 (N_12549,N_11005,N_11506);
or U12550 (N_12550,N_11722,N_11504);
or U12551 (N_12551,N_11231,N_11985);
xnor U12552 (N_12552,N_11056,N_11099);
or U12553 (N_12553,N_11803,N_11005);
and U12554 (N_12554,N_11972,N_11142);
xnor U12555 (N_12555,N_11065,N_11939);
nor U12556 (N_12556,N_11607,N_11988);
or U12557 (N_12557,N_11882,N_11970);
and U12558 (N_12558,N_11185,N_11229);
nand U12559 (N_12559,N_11827,N_11578);
or U12560 (N_12560,N_11500,N_11076);
and U12561 (N_12561,N_11066,N_11126);
nand U12562 (N_12562,N_11755,N_11408);
or U12563 (N_12563,N_11178,N_11327);
or U12564 (N_12564,N_11833,N_11943);
or U12565 (N_12565,N_11392,N_11205);
and U12566 (N_12566,N_11476,N_11761);
nand U12567 (N_12567,N_11228,N_11968);
or U12568 (N_12568,N_11789,N_11231);
nand U12569 (N_12569,N_11407,N_11477);
xnor U12570 (N_12570,N_11651,N_11677);
or U12571 (N_12571,N_11712,N_11324);
nor U12572 (N_12572,N_11838,N_11408);
nor U12573 (N_12573,N_11099,N_11202);
and U12574 (N_12574,N_11547,N_11286);
nor U12575 (N_12575,N_11614,N_11780);
nor U12576 (N_12576,N_11208,N_11562);
nor U12577 (N_12577,N_11116,N_11475);
nand U12578 (N_12578,N_11490,N_11137);
nand U12579 (N_12579,N_11754,N_11052);
nand U12580 (N_12580,N_11316,N_11519);
nor U12581 (N_12581,N_11419,N_11136);
nand U12582 (N_12582,N_11466,N_11001);
nand U12583 (N_12583,N_11206,N_11489);
nand U12584 (N_12584,N_11282,N_11473);
or U12585 (N_12585,N_11858,N_11429);
nand U12586 (N_12586,N_11612,N_11391);
nand U12587 (N_12587,N_11565,N_11438);
or U12588 (N_12588,N_11388,N_11594);
nand U12589 (N_12589,N_11073,N_11950);
nand U12590 (N_12590,N_11847,N_11138);
nor U12591 (N_12591,N_11368,N_11630);
xor U12592 (N_12592,N_11318,N_11366);
xnor U12593 (N_12593,N_11267,N_11292);
and U12594 (N_12594,N_11353,N_11900);
nor U12595 (N_12595,N_11616,N_11061);
and U12596 (N_12596,N_11929,N_11063);
nand U12597 (N_12597,N_11856,N_11016);
nor U12598 (N_12598,N_11079,N_11766);
nor U12599 (N_12599,N_11769,N_11710);
or U12600 (N_12600,N_11275,N_11409);
xnor U12601 (N_12601,N_11303,N_11936);
xnor U12602 (N_12602,N_11728,N_11726);
nor U12603 (N_12603,N_11289,N_11720);
nand U12604 (N_12604,N_11717,N_11463);
nand U12605 (N_12605,N_11107,N_11887);
and U12606 (N_12606,N_11946,N_11002);
and U12607 (N_12607,N_11720,N_11717);
xnor U12608 (N_12608,N_11637,N_11909);
and U12609 (N_12609,N_11874,N_11315);
and U12610 (N_12610,N_11364,N_11638);
nand U12611 (N_12611,N_11142,N_11146);
xnor U12612 (N_12612,N_11149,N_11906);
and U12613 (N_12613,N_11866,N_11376);
nor U12614 (N_12614,N_11190,N_11369);
and U12615 (N_12615,N_11363,N_11401);
nand U12616 (N_12616,N_11372,N_11146);
xnor U12617 (N_12617,N_11418,N_11020);
or U12618 (N_12618,N_11355,N_11502);
xnor U12619 (N_12619,N_11253,N_11940);
nand U12620 (N_12620,N_11107,N_11606);
nor U12621 (N_12621,N_11148,N_11842);
xnor U12622 (N_12622,N_11572,N_11381);
nor U12623 (N_12623,N_11832,N_11206);
nand U12624 (N_12624,N_11769,N_11248);
or U12625 (N_12625,N_11879,N_11094);
or U12626 (N_12626,N_11868,N_11313);
and U12627 (N_12627,N_11942,N_11219);
and U12628 (N_12628,N_11762,N_11300);
nor U12629 (N_12629,N_11734,N_11456);
xor U12630 (N_12630,N_11308,N_11728);
and U12631 (N_12631,N_11187,N_11938);
nor U12632 (N_12632,N_11457,N_11468);
and U12633 (N_12633,N_11318,N_11319);
xnor U12634 (N_12634,N_11414,N_11262);
or U12635 (N_12635,N_11598,N_11400);
nor U12636 (N_12636,N_11156,N_11779);
nor U12637 (N_12637,N_11395,N_11050);
xor U12638 (N_12638,N_11844,N_11973);
nand U12639 (N_12639,N_11208,N_11006);
nor U12640 (N_12640,N_11605,N_11249);
xnor U12641 (N_12641,N_11687,N_11490);
nor U12642 (N_12642,N_11402,N_11979);
nor U12643 (N_12643,N_11955,N_11202);
and U12644 (N_12644,N_11497,N_11795);
and U12645 (N_12645,N_11874,N_11344);
and U12646 (N_12646,N_11100,N_11603);
nand U12647 (N_12647,N_11011,N_11412);
xor U12648 (N_12648,N_11563,N_11408);
nand U12649 (N_12649,N_11786,N_11834);
xor U12650 (N_12650,N_11132,N_11986);
and U12651 (N_12651,N_11783,N_11209);
or U12652 (N_12652,N_11576,N_11183);
and U12653 (N_12653,N_11104,N_11414);
or U12654 (N_12654,N_11792,N_11747);
nor U12655 (N_12655,N_11067,N_11186);
or U12656 (N_12656,N_11724,N_11342);
or U12657 (N_12657,N_11913,N_11152);
xor U12658 (N_12658,N_11868,N_11711);
xnor U12659 (N_12659,N_11497,N_11141);
and U12660 (N_12660,N_11860,N_11669);
or U12661 (N_12661,N_11247,N_11363);
or U12662 (N_12662,N_11263,N_11481);
or U12663 (N_12663,N_11027,N_11940);
or U12664 (N_12664,N_11078,N_11663);
nor U12665 (N_12665,N_11540,N_11682);
or U12666 (N_12666,N_11565,N_11132);
or U12667 (N_12667,N_11480,N_11830);
nand U12668 (N_12668,N_11157,N_11381);
nor U12669 (N_12669,N_11637,N_11970);
nor U12670 (N_12670,N_11651,N_11866);
nor U12671 (N_12671,N_11103,N_11042);
and U12672 (N_12672,N_11483,N_11577);
nand U12673 (N_12673,N_11449,N_11544);
and U12674 (N_12674,N_11259,N_11687);
nand U12675 (N_12675,N_11958,N_11413);
or U12676 (N_12676,N_11882,N_11197);
or U12677 (N_12677,N_11701,N_11101);
and U12678 (N_12678,N_11518,N_11564);
xnor U12679 (N_12679,N_11521,N_11687);
or U12680 (N_12680,N_11335,N_11338);
and U12681 (N_12681,N_11022,N_11458);
and U12682 (N_12682,N_11059,N_11642);
or U12683 (N_12683,N_11158,N_11113);
xnor U12684 (N_12684,N_11426,N_11318);
and U12685 (N_12685,N_11819,N_11722);
or U12686 (N_12686,N_11364,N_11974);
nor U12687 (N_12687,N_11652,N_11340);
nand U12688 (N_12688,N_11681,N_11782);
xor U12689 (N_12689,N_11933,N_11319);
nand U12690 (N_12690,N_11834,N_11078);
nor U12691 (N_12691,N_11795,N_11397);
xor U12692 (N_12692,N_11449,N_11008);
or U12693 (N_12693,N_11819,N_11554);
or U12694 (N_12694,N_11800,N_11476);
xnor U12695 (N_12695,N_11853,N_11017);
nand U12696 (N_12696,N_11136,N_11801);
nand U12697 (N_12697,N_11816,N_11773);
xor U12698 (N_12698,N_11371,N_11776);
nor U12699 (N_12699,N_11417,N_11276);
nand U12700 (N_12700,N_11028,N_11471);
nor U12701 (N_12701,N_11335,N_11987);
nand U12702 (N_12702,N_11779,N_11031);
nand U12703 (N_12703,N_11174,N_11621);
or U12704 (N_12704,N_11412,N_11185);
xnor U12705 (N_12705,N_11348,N_11560);
and U12706 (N_12706,N_11508,N_11976);
xnor U12707 (N_12707,N_11371,N_11893);
nor U12708 (N_12708,N_11589,N_11628);
xor U12709 (N_12709,N_11612,N_11361);
xor U12710 (N_12710,N_11942,N_11527);
xor U12711 (N_12711,N_11016,N_11414);
nor U12712 (N_12712,N_11608,N_11649);
nor U12713 (N_12713,N_11010,N_11905);
xor U12714 (N_12714,N_11179,N_11292);
nand U12715 (N_12715,N_11779,N_11453);
nor U12716 (N_12716,N_11008,N_11756);
or U12717 (N_12717,N_11641,N_11599);
and U12718 (N_12718,N_11858,N_11234);
or U12719 (N_12719,N_11352,N_11213);
or U12720 (N_12720,N_11240,N_11721);
nand U12721 (N_12721,N_11983,N_11168);
xor U12722 (N_12722,N_11656,N_11599);
xnor U12723 (N_12723,N_11211,N_11553);
nor U12724 (N_12724,N_11899,N_11117);
and U12725 (N_12725,N_11794,N_11396);
nor U12726 (N_12726,N_11324,N_11290);
xnor U12727 (N_12727,N_11181,N_11789);
nor U12728 (N_12728,N_11933,N_11357);
or U12729 (N_12729,N_11915,N_11743);
and U12730 (N_12730,N_11796,N_11515);
xor U12731 (N_12731,N_11634,N_11636);
or U12732 (N_12732,N_11260,N_11429);
or U12733 (N_12733,N_11005,N_11384);
nor U12734 (N_12734,N_11529,N_11808);
nand U12735 (N_12735,N_11332,N_11633);
nand U12736 (N_12736,N_11945,N_11723);
or U12737 (N_12737,N_11514,N_11298);
xor U12738 (N_12738,N_11903,N_11598);
nand U12739 (N_12739,N_11873,N_11567);
and U12740 (N_12740,N_11503,N_11750);
and U12741 (N_12741,N_11834,N_11688);
nor U12742 (N_12742,N_11576,N_11650);
or U12743 (N_12743,N_11008,N_11703);
and U12744 (N_12744,N_11856,N_11706);
or U12745 (N_12745,N_11858,N_11873);
nand U12746 (N_12746,N_11005,N_11174);
xnor U12747 (N_12747,N_11877,N_11413);
xor U12748 (N_12748,N_11097,N_11098);
nor U12749 (N_12749,N_11126,N_11496);
nor U12750 (N_12750,N_11372,N_11200);
and U12751 (N_12751,N_11150,N_11030);
nand U12752 (N_12752,N_11760,N_11383);
nor U12753 (N_12753,N_11012,N_11922);
xor U12754 (N_12754,N_11158,N_11911);
nor U12755 (N_12755,N_11611,N_11838);
nor U12756 (N_12756,N_11415,N_11783);
nand U12757 (N_12757,N_11506,N_11143);
nor U12758 (N_12758,N_11194,N_11110);
nor U12759 (N_12759,N_11041,N_11837);
nor U12760 (N_12760,N_11057,N_11112);
nor U12761 (N_12761,N_11361,N_11153);
or U12762 (N_12762,N_11300,N_11527);
or U12763 (N_12763,N_11994,N_11645);
and U12764 (N_12764,N_11232,N_11365);
nor U12765 (N_12765,N_11468,N_11807);
nand U12766 (N_12766,N_11788,N_11499);
nand U12767 (N_12767,N_11526,N_11565);
nor U12768 (N_12768,N_11120,N_11939);
xor U12769 (N_12769,N_11867,N_11633);
xor U12770 (N_12770,N_11947,N_11078);
nor U12771 (N_12771,N_11794,N_11968);
xor U12772 (N_12772,N_11516,N_11011);
xnor U12773 (N_12773,N_11483,N_11874);
xnor U12774 (N_12774,N_11427,N_11693);
or U12775 (N_12775,N_11856,N_11320);
nand U12776 (N_12776,N_11953,N_11664);
and U12777 (N_12777,N_11277,N_11928);
xnor U12778 (N_12778,N_11750,N_11891);
and U12779 (N_12779,N_11031,N_11871);
nand U12780 (N_12780,N_11038,N_11986);
nand U12781 (N_12781,N_11682,N_11118);
xnor U12782 (N_12782,N_11222,N_11571);
and U12783 (N_12783,N_11464,N_11172);
and U12784 (N_12784,N_11696,N_11852);
and U12785 (N_12785,N_11538,N_11062);
xor U12786 (N_12786,N_11997,N_11403);
and U12787 (N_12787,N_11458,N_11089);
and U12788 (N_12788,N_11572,N_11011);
nand U12789 (N_12789,N_11153,N_11588);
nor U12790 (N_12790,N_11631,N_11725);
xor U12791 (N_12791,N_11777,N_11320);
xnor U12792 (N_12792,N_11429,N_11237);
nor U12793 (N_12793,N_11665,N_11075);
nor U12794 (N_12794,N_11201,N_11260);
and U12795 (N_12795,N_11558,N_11399);
xnor U12796 (N_12796,N_11146,N_11286);
and U12797 (N_12797,N_11771,N_11316);
nor U12798 (N_12798,N_11522,N_11931);
or U12799 (N_12799,N_11332,N_11051);
nand U12800 (N_12800,N_11887,N_11247);
or U12801 (N_12801,N_11511,N_11209);
nand U12802 (N_12802,N_11451,N_11087);
or U12803 (N_12803,N_11281,N_11780);
nor U12804 (N_12804,N_11742,N_11615);
and U12805 (N_12805,N_11530,N_11458);
nand U12806 (N_12806,N_11670,N_11584);
nand U12807 (N_12807,N_11023,N_11439);
nor U12808 (N_12808,N_11165,N_11124);
nand U12809 (N_12809,N_11569,N_11188);
and U12810 (N_12810,N_11565,N_11680);
xor U12811 (N_12811,N_11520,N_11988);
or U12812 (N_12812,N_11250,N_11808);
nand U12813 (N_12813,N_11204,N_11993);
nand U12814 (N_12814,N_11672,N_11605);
and U12815 (N_12815,N_11286,N_11611);
or U12816 (N_12816,N_11361,N_11023);
nand U12817 (N_12817,N_11776,N_11322);
or U12818 (N_12818,N_11126,N_11951);
xnor U12819 (N_12819,N_11738,N_11392);
nor U12820 (N_12820,N_11402,N_11557);
or U12821 (N_12821,N_11860,N_11613);
nor U12822 (N_12822,N_11436,N_11196);
nor U12823 (N_12823,N_11952,N_11383);
nor U12824 (N_12824,N_11599,N_11111);
nor U12825 (N_12825,N_11260,N_11864);
xnor U12826 (N_12826,N_11712,N_11801);
or U12827 (N_12827,N_11486,N_11436);
and U12828 (N_12828,N_11488,N_11506);
nor U12829 (N_12829,N_11518,N_11288);
nand U12830 (N_12830,N_11201,N_11108);
xnor U12831 (N_12831,N_11227,N_11155);
nand U12832 (N_12832,N_11553,N_11459);
and U12833 (N_12833,N_11446,N_11673);
or U12834 (N_12834,N_11995,N_11905);
and U12835 (N_12835,N_11405,N_11802);
or U12836 (N_12836,N_11192,N_11525);
nand U12837 (N_12837,N_11562,N_11707);
nand U12838 (N_12838,N_11864,N_11076);
xnor U12839 (N_12839,N_11350,N_11973);
xor U12840 (N_12840,N_11366,N_11618);
xnor U12841 (N_12841,N_11013,N_11171);
xnor U12842 (N_12842,N_11305,N_11176);
or U12843 (N_12843,N_11459,N_11991);
or U12844 (N_12844,N_11335,N_11325);
nand U12845 (N_12845,N_11557,N_11693);
xnor U12846 (N_12846,N_11973,N_11418);
nor U12847 (N_12847,N_11367,N_11394);
xor U12848 (N_12848,N_11261,N_11823);
or U12849 (N_12849,N_11095,N_11771);
or U12850 (N_12850,N_11525,N_11487);
or U12851 (N_12851,N_11131,N_11964);
and U12852 (N_12852,N_11174,N_11233);
xnor U12853 (N_12853,N_11309,N_11713);
nor U12854 (N_12854,N_11393,N_11305);
nor U12855 (N_12855,N_11159,N_11275);
xnor U12856 (N_12856,N_11619,N_11308);
and U12857 (N_12857,N_11298,N_11573);
and U12858 (N_12858,N_11576,N_11995);
or U12859 (N_12859,N_11475,N_11727);
xor U12860 (N_12860,N_11859,N_11485);
and U12861 (N_12861,N_11763,N_11199);
xnor U12862 (N_12862,N_11041,N_11897);
nor U12863 (N_12863,N_11094,N_11014);
or U12864 (N_12864,N_11620,N_11032);
and U12865 (N_12865,N_11273,N_11762);
nand U12866 (N_12866,N_11225,N_11224);
or U12867 (N_12867,N_11020,N_11513);
nand U12868 (N_12868,N_11098,N_11551);
nor U12869 (N_12869,N_11807,N_11893);
nand U12870 (N_12870,N_11557,N_11263);
and U12871 (N_12871,N_11924,N_11922);
xnor U12872 (N_12872,N_11600,N_11408);
nand U12873 (N_12873,N_11690,N_11718);
nor U12874 (N_12874,N_11481,N_11115);
nor U12875 (N_12875,N_11867,N_11860);
xnor U12876 (N_12876,N_11481,N_11189);
and U12877 (N_12877,N_11461,N_11196);
xnor U12878 (N_12878,N_11644,N_11214);
nand U12879 (N_12879,N_11764,N_11972);
and U12880 (N_12880,N_11471,N_11619);
xnor U12881 (N_12881,N_11061,N_11396);
nor U12882 (N_12882,N_11923,N_11872);
or U12883 (N_12883,N_11868,N_11092);
xor U12884 (N_12884,N_11654,N_11365);
nor U12885 (N_12885,N_11913,N_11332);
or U12886 (N_12886,N_11737,N_11239);
xnor U12887 (N_12887,N_11488,N_11231);
xnor U12888 (N_12888,N_11764,N_11674);
or U12889 (N_12889,N_11570,N_11288);
nand U12890 (N_12890,N_11640,N_11683);
nor U12891 (N_12891,N_11628,N_11689);
xor U12892 (N_12892,N_11951,N_11442);
and U12893 (N_12893,N_11399,N_11783);
or U12894 (N_12894,N_11199,N_11048);
nand U12895 (N_12895,N_11887,N_11663);
nor U12896 (N_12896,N_11384,N_11185);
xnor U12897 (N_12897,N_11527,N_11958);
and U12898 (N_12898,N_11528,N_11127);
or U12899 (N_12899,N_11882,N_11382);
and U12900 (N_12900,N_11345,N_11897);
nand U12901 (N_12901,N_11236,N_11736);
xnor U12902 (N_12902,N_11982,N_11697);
and U12903 (N_12903,N_11071,N_11093);
or U12904 (N_12904,N_11194,N_11103);
nor U12905 (N_12905,N_11968,N_11953);
and U12906 (N_12906,N_11205,N_11034);
xnor U12907 (N_12907,N_11309,N_11291);
nand U12908 (N_12908,N_11762,N_11592);
or U12909 (N_12909,N_11559,N_11923);
and U12910 (N_12910,N_11047,N_11363);
xor U12911 (N_12911,N_11128,N_11661);
and U12912 (N_12912,N_11288,N_11976);
nand U12913 (N_12913,N_11933,N_11964);
or U12914 (N_12914,N_11475,N_11382);
or U12915 (N_12915,N_11947,N_11705);
xor U12916 (N_12916,N_11641,N_11203);
nor U12917 (N_12917,N_11643,N_11857);
or U12918 (N_12918,N_11277,N_11710);
nand U12919 (N_12919,N_11349,N_11410);
xnor U12920 (N_12920,N_11970,N_11607);
xor U12921 (N_12921,N_11174,N_11086);
nor U12922 (N_12922,N_11294,N_11118);
nor U12923 (N_12923,N_11004,N_11370);
or U12924 (N_12924,N_11045,N_11555);
xor U12925 (N_12925,N_11726,N_11671);
and U12926 (N_12926,N_11846,N_11880);
nor U12927 (N_12927,N_11332,N_11805);
or U12928 (N_12928,N_11928,N_11394);
or U12929 (N_12929,N_11634,N_11535);
nor U12930 (N_12930,N_11112,N_11156);
xnor U12931 (N_12931,N_11281,N_11845);
xor U12932 (N_12932,N_11783,N_11701);
nand U12933 (N_12933,N_11130,N_11302);
nand U12934 (N_12934,N_11264,N_11931);
and U12935 (N_12935,N_11266,N_11859);
xor U12936 (N_12936,N_11868,N_11174);
nor U12937 (N_12937,N_11943,N_11594);
nand U12938 (N_12938,N_11810,N_11262);
nand U12939 (N_12939,N_11483,N_11934);
xnor U12940 (N_12940,N_11363,N_11559);
nor U12941 (N_12941,N_11055,N_11722);
xnor U12942 (N_12942,N_11297,N_11604);
and U12943 (N_12943,N_11936,N_11279);
xnor U12944 (N_12944,N_11863,N_11796);
or U12945 (N_12945,N_11382,N_11510);
xor U12946 (N_12946,N_11356,N_11431);
or U12947 (N_12947,N_11199,N_11486);
xnor U12948 (N_12948,N_11518,N_11254);
and U12949 (N_12949,N_11444,N_11135);
xnor U12950 (N_12950,N_11962,N_11593);
and U12951 (N_12951,N_11692,N_11033);
xor U12952 (N_12952,N_11651,N_11872);
xnor U12953 (N_12953,N_11657,N_11816);
or U12954 (N_12954,N_11964,N_11689);
xnor U12955 (N_12955,N_11000,N_11068);
nand U12956 (N_12956,N_11360,N_11243);
or U12957 (N_12957,N_11965,N_11369);
xor U12958 (N_12958,N_11084,N_11447);
and U12959 (N_12959,N_11372,N_11128);
and U12960 (N_12960,N_11564,N_11623);
nand U12961 (N_12961,N_11570,N_11690);
or U12962 (N_12962,N_11119,N_11145);
nor U12963 (N_12963,N_11812,N_11513);
or U12964 (N_12964,N_11432,N_11422);
and U12965 (N_12965,N_11221,N_11943);
nand U12966 (N_12966,N_11495,N_11892);
xor U12967 (N_12967,N_11210,N_11430);
or U12968 (N_12968,N_11065,N_11395);
nor U12969 (N_12969,N_11359,N_11218);
nor U12970 (N_12970,N_11090,N_11439);
xnor U12971 (N_12971,N_11212,N_11083);
nor U12972 (N_12972,N_11657,N_11859);
xor U12973 (N_12973,N_11311,N_11225);
xnor U12974 (N_12974,N_11128,N_11827);
or U12975 (N_12975,N_11986,N_11168);
xor U12976 (N_12976,N_11595,N_11273);
and U12977 (N_12977,N_11063,N_11284);
or U12978 (N_12978,N_11544,N_11212);
or U12979 (N_12979,N_11587,N_11480);
nand U12980 (N_12980,N_11289,N_11888);
nor U12981 (N_12981,N_11162,N_11062);
xor U12982 (N_12982,N_11184,N_11388);
xor U12983 (N_12983,N_11224,N_11963);
nand U12984 (N_12984,N_11844,N_11663);
or U12985 (N_12985,N_11334,N_11542);
nor U12986 (N_12986,N_11256,N_11619);
nor U12987 (N_12987,N_11959,N_11433);
nand U12988 (N_12988,N_11956,N_11985);
nand U12989 (N_12989,N_11386,N_11875);
nor U12990 (N_12990,N_11040,N_11268);
or U12991 (N_12991,N_11770,N_11691);
nor U12992 (N_12992,N_11193,N_11457);
nor U12993 (N_12993,N_11599,N_11438);
or U12994 (N_12994,N_11707,N_11921);
and U12995 (N_12995,N_11068,N_11748);
nand U12996 (N_12996,N_11128,N_11287);
and U12997 (N_12997,N_11010,N_11365);
or U12998 (N_12998,N_11173,N_11571);
or U12999 (N_12999,N_11206,N_11321);
or U13000 (N_13000,N_12808,N_12324);
xnor U13001 (N_13001,N_12529,N_12336);
nor U13002 (N_13002,N_12475,N_12456);
nor U13003 (N_13003,N_12392,N_12589);
and U13004 (N_13004,N_12240,N_12765);
nor U13005 (N_13005,N_12120,N_12809);
or U13006 (N_13006,N_12648,N_12119);
and U13007 (N_13007,N_12834,N_12368);
or U13008 (N_13008,N_12212,N_12201);
nor U13009 (N_13009,N_12527,N_12069);
and U13010 (N_13010,N_12362,N_12867);
nand U13011 (N_13011,N_12854,N_12578);
nand U13012 (N_13012,N_12043,N_12881);
nand U13013 (N_13013,N_12477,N_12889);
nor U13014 (N_13014,N_12391,N_12180);
nor U13015 (N_13015,N_12737,N_12520);
nor U13016 (N_13016,N_12424,N_12715);
xor U13017 (N_13017,N_12916,N_12186);
or U13018 (N_13018,N_12663,N_12866);
and U13019 (N_13019,N_12402,N_12455);
and U13020 (N_13020,N_12683,N_12703);
and U13021 (N_13021,N_12813,N_12577);
nand U13022 (N_13022,N_12123,N_12969);
nand U13023 (N_13023,N_12932,N_12443);
nand U13024 (N_13024,N_12080,N_12386);
nor U13025 (N_13025,N_12526,N_12025);
and U13026 (N_13026,N_12507,N_12549);
nand U13027 (N_13027,N_12206,N_12413);
or U13028 (N_13028,N_12372,N_12490);
xor U13029 (N_13029,N_12097,N_12758);
nand U13030 (N_13030,N_12159,N_12143);
nor U13031 (N_13031,N_12269,N_12566);
or U13032 (N_13032,N_12951,N_12978);
nand U13033 (N_13033,N_12640,N_12914);
and U13034 (N_13034,N_12014,N_12593);
and U13035 (N_13035,N_12620,N_12795);
nor U13036 (N_13036,N_12208,N_12875);
nand U13037 (N_13037,N_12845,N_12855);
or U13038 (N_13038,N_12244,N_12209);
and U13039 (N_13039,N_12289,N_12861);
or U13040 (N_13040,N_12060,N_12117);
nand U13041 (N_13041,N_12639,N_12325);
nand U13042 (N_13042,N_12283,N_12258);
and U13043 (N_13043,N_12374,N_12636);
or U13044 (N_13044,N_12231,N_12411);
nand U13045 (N_13045,N_12706,N_12385);
nor U13046 (N_13046,N_12452,N_12887);
nor U13047 (N_13047,N_12781,N_12766);
and U13048 (N_13048,N_12264,N_12418);
nand U13049 (N_13049,N_12001,N_12437);
and U13050 (N_13050,N_12613,N_12905);
and U13051 (N_13051,N_12751,N_12771);
nand U13052 (N_13052,N_12516,N_12225);
and U13053 (N_13053,N_12864,N_12545);
nor U13054 (N_13054,N_12759,N_12846);
and U13055 (N_13055,N_12695,N_12536);
or U13056 (N_13056,N_12806,N_12515);
or U13057 (N_13057,N_12174,N_12879);
xnor U13058 (N_13058,N_12668,N_12612);
xnor U13059 (N_13059,N_12811,N_12518);
xnor U13060 (N_13060,N_12434,N_12246);
nor U13061 (N_13061,N_12361,N_12915);
and U13062 (N_13062,N_12632,N_12053);
nand U13063 (N_13063,N_12860,N_12601);
or U13064 (N_13064,N_12830,N_12277);
nor U13065 (N_13065,N_12743,N_12128);
xor U13066 (N_13066,N_12262,N_12882);
and U13067 (N_13067,N_12450,N_12054);
nand U13068 (N_13068,N_12422,N_12344);
or U13069 (N_13069,N_12736,N_12740);
nor U13070 (N_13070,N_12934,N_12702);
xor U13071 (N_13071,N_12484,N_12175);
and U13072 (N_13072,N_12606,N_12833);
nor U13073 (N_13073,N_12532,N_12233);
nor U13074 (N_13074,N_12780,N_12533);
nand U13075 (N_13075,N_12318,N_12787);
nor U13076 (N_13076,N_12221,N_12366);
or U13077 (N_13077,N_12219,N_12114);
or U13078 (N_13078,N_12523,N_12598);
or U13079 (N_13079,N_12343,N_12460);
nand U13080 (N_13080,N_12965,N_12608);
xnor U13081 (N_13081,N_12410,N_12548);
xnor U13082 (N_13082,N_12415,N_12302);
and U13083 (N_13083,N_12597,N_12397);
and U13084 (N_13084,N_12627,N_12018);
nand U13085 (N_13085,N_12552,N_12837);
or U13086 (N_13086,N_12818,N_12735);
xnor U13087 (N_13087,N_12382,N_12457);
and U13088 (N_13088,N_12857,N_12746);
nand U13089 (N_13089,N_12616,N_12692);
nor U13090 (N_13090,N_12952,N_12425);
xor U13091 (N_13091,N_12282,N_12429);
nand U13092 (N_13092,N_12888,N_12925);
and U13093 (N_13093,N_12234,N_12885);
xor U13094 (N_13094,N_12676,N_12851);
nor U13095 (N_13095,N_12033,N_12739);
nor U13096 (N_13096,N_12802,N_12842);
and U13097 (N_13097,N_12169,N_12057);
and U13098 (N_13098,N_12728,N_12084);
and U13099 (N_13099,N_12870,N_12367);
or U13100 (N_13100,N_12699,N_12665);
nor U13101 (N_13101,N_12290,N_12610);
xor U13102 (N_13102,N_12989,N_12364);
nand U13103 (N_13103,N_12317,N_12957);
nor U13104 (N_13104,N_12022,N_12605);
nor U13105 (N_13105,N_12034,N_12819);
nand U13106 (N_13106,N_12750,N_12296);
xor U13107 (N_13107,N_12850,N_12971);
or U13108 (N_13108,N_12690,N_12824);
or U13109 (N_13109,N_12253,N_12044);
or U13110 (N_13110,N_12694,N_12094);
nand U13111 (N_13111,N_12917,N_12782);
and U13112 (N_13112,N_12675,N_12964);
and U13113 (N_13113,N_12602,N_12198);
and U13114 (N_13114,N_12954,N_12155);
or U13115 (N_13115,N_12546,N_12300);
xor U13116 (N_13116,N_12310,N_12312);
nand U13117 (N_13117,N_12346,N_12112);
and U13118 (N_13118,N_12307,N_12028);
or U13119 (N_13119,N_12604,N_12946);
and U13120 (N_13120,N_12685,N_12229);
and U13121 (N_13121,N_12775,N_12512);
and U13122 (N_13122,N_12817,N_12628);
nand U13123 (N_13123,N_12567,N_12150);
and U13124 (N_13124,N_12328,N_12899);
xnor U13125 (N_13125,N_12907,N_12862);
and U13126 (N_13126,N_12708,N_12918);
xor U13127 (N_13127,N_12510,N_12213);
xor U13128 (N_13128,N_12394,N_12251);
and U13129 (N_13129,N_12810,N_12467);
and U13130 (N_13130,N_12711,N_12256);
or U13131 (N_13131,N_12752,N_12431);
nand U13132 (N_13132,N_12327,N_12294);
nor U13133 (N_13133,N_12586,N_12458);
nand U13134 (N_13134,N_12634,N_12511);
or U13135 (N_13135,N_12748,N_12508);
and U13136 (N_13136,N_12331,N_12333);
nor U13137 (N_13137,N_12408,N_12961);
or U13138 (N_13138,N_12853,N_12365);
nor U13139 (N_13139,N_12375,N_12357);
xnor U13140 (N_13140,N_12962,N_12565);
nand U13141 (N_13141,N_12009,N_12556);
xnor U13142 (N_13142,N_12933,N_12956);
nand U13143 (N_13143,N_12931,N_12731);
nor U13144 (N_13144,N_12579,N_12188);
xor U13145 (N_13145,N_12684,N_12705);
and U13146 (N_13146,N_12136,N_12129);
or U13147 (N_13147,N_12066,N_12430);
nand U13148 (N_13148,N_12807,N_12921);
nand U13149 (N_13149,N_12544,N_12770);
or U13150 (N_13150,N_12741,N_12911);
nand U13151 (N_13151,N_12662,N_12189);
nand U13152 (N_13152,N_12109,N_12164);
nor U13153 (N_13153,N_12015,N_12255);
xor U13154 (N_13154,N_12894,N_12814);
nor U13155 (N_13155,N_12358,N_12997);
xnor U13156 (N_13156,N_12877,N_12591);
or U13157 (N_13157,N_12047,N_12412);
nand U13158 (N_13158,N_12733,N_12330);
and U13159 (N_13159,N_12267,N_12400);
nor U13160 (N_13160,N_12643,N_12998);
nand U13161 (N_13161,N_12263,N_12531);
nor U13162 (N_13162,N_12826,N_12700);
or U13163 (N_13163,N_12535,N_12626);
and U13164 (N_13164,N_12927,N_12377);
nand U13165 (N_13165,N_12192,N_12827);
and U13166 (N_13166,N_12509,N_12645);
nor U13167 (N_13167,N_12287,N_12607);
nor U13168 (N_13168,N_12704,N_12351);
nand U13169 (N_13169,N_12995,N_12557);
xor U13170 (N_13170,N_12165,N_12359);
xor U13171 (N_13171,N_12134,N_12744);
xnor U13172 (N_13172,N_12769,N_12674);
or U13173 (N_13173,N_12030,N_12204);
or U13174 (N_13174,N_12023,N_12760);
nand U13175 (N_13175,N_12100,N_12801);
and U13176 (N_13176,N_12168,N_12090);
nor U13177 (N_13177,N_12268,N_12580);
xor U13178 (N_13178,N_12913,N_12970);
xor U13179 (N_13179,N_12145,N_12761);
nand U13180 (N_13180,N_12207,N_12172);
nor U13181 (N_13181,N_12503,N_12539);
nand U13182 (N_13182,N_12470,N_12012);
nor U13183 (N_13183,N_12754,N_12401);
xnor U13184 (N_13184,N_12609,N_12250);
nor U13185 (N_13185,N_12494,N_12592);
xnor U13186 (N_13186,N_12187,N_12461);
nor U13187 (N_13187,N_12305,N_12039);
and U13188 (N_13188,N_12976,N_12874);
and U13189 (N_13189,N_12082,N_12716);
and U13190 (N_13190,N_12211,N_12311);
or U13191 (N_13191,N_12275,N_12682);
xnor U13192 (N_13192,N_12149,N_12999);
nand U13193 (N_13193,N_12950,N_12537);
nor U13194 (N_13194,N_12163,N_12876);
nand U13195 (N_13195,N_12166,N_12061);
xor U13196 (N_13196,N_12642,N_12319);
or U13197 (N_13197,N_12462,N_12466);
nand U13198 (N_13198,N_12659,N_12492);
xnor U13199 (N_13199,N_12451,N_12326);
or U13200 (N_13200,N_12156,N_12936);
xor U13201 (N_13201,N_12661,N_12032);
nand U13202 (N_13202,N_12079,N_12767);
and U13203 (N_13203,N_12215,N_12791);
and U13204 (N_13204,N_12341,N_12924);
or U13205 (N_13205,N_12599,N_12352);
or U13206 (N_13206,N_12796,N_12836);
nand U13207 (N_13207,N_12261,N_12587);
nor U13208 (N_13208,N_12922,N_12856);
nor U13209 (N_13209,N_12170,N_12983);
nor U13210 (N_13210,N_12726,N_12930);
or U13211 (N_13211,N_12181,N_12617);
xor U13212 (N_13212,N_12785,N_12232);
xor U13213 (N_13213,N_12140,N_12349);
xnor U13214 (N_13214,N_12757,N_12502);
xor U13215 (N_13215,N_12554,N_12297);
xnor U13216 (N_13216,N_12935,N_12217);
nand U13217 (N_13217,N_12110,N_12235);
xnor U13218 (N_13218,N_12220,N_12649);
nand U13219 (N_13219,N_12948,N_12384);
nor U13220 (N_13220,N_12265,N_12072);
or U13221 (N_13221,N_12776,N_12293);
xor U13222 (N_13222,N_12393,N_12485);
and U13223 (N_13223,N_12495,N_12438);
nand U13224 (N_13224,N_12010,N_12210);
or U13225 (N_13225,N_12959,N_12650);
and U13226 (N_13226,N_12644,N_12421);
or U13227 (N_13227,N_12398,N_12897);
or U13228 (N_13228,N_12623,N_12555);
xnor U13229 (N_13229,N_12445,N_12839);
nor U13230 (N_13230,N_12065,N_12340);
xor U13231 (N_13231,N_12274,N_12202);
nand U13232 (N_13232,N_12026,N_12142);
xor U13233 (N_13233,N_12658,N_12329);
or U13234 (N_13234,N_12360,N_12019);
or U13235 (N_13235,N_12476,N_12588);
xor U13236 (N_13236,N_12670,N_12928);
nor U13237 (N_13237,N_12416,N_12073);
and U13238 (N_13238,N_12064,N_12713);
nand U13239 (N_13239,N_12800,N_12603);
xor U13240 (N_13240,N_12056,N_12525);
nor U13241 (N_13241,N_12104,N_12178);
xnor U13242 (N_13242,N_12342,N_12519);
xor U13243 (N_13243,N_12852,N_12841);
nand U13244 (N_13244,N_12228,N_12666);
and U13245 (N_13245,N_12717,N_12063);
nand U13246 (N_13246,N_12257,N_12468);
nand U13247 (N_13247,N_12505,N_12254);
or U13248 (N_13248,N_12653,N_12582);
or U13249 (N_13249,N_12500,N_12572);
and U13250 (N_13250,N_12637,N_12448);
xor U13251 (N_13251,N_12943,N_12825);
nand U13252 (N_13252,N_12444,N_12903);
nor U13253 (N_13253,N_12173,N_12847);
and U13254 (N_13254,N_12541,N_12832);
nand U13255 (N_13255,N_12303,N_12067);
nor U13256 (N_13256,N_12171,N_12153);
xnor U13257 (N_13257,N_12869,N_12029);
or U13258 (N_13258,N_12972,N_12974);
nor U13259 (N_13259,N_12276,N_12020);
and U13260 (N_13260,N_12772,N_12304);
and U13261 (N_13261,N_12904,N_12195);
nor U13262 (N_13262,N_12160,N_12900);
or U13263 (N_13263,N_12162,N_12147);
or U13264 (N_13264,N_12322,N_12611);
nand U13265 (N_13265,N_12161,N_12988);
nor U13266 (N_13266,N_12655,N_12929);
or U13267 (N_13267,N_12794,N_12177);
nor U13268 (N_13268,N_12724,N_12944);
and U13269 (N_13269,N_12436,N_12105);
xnor U13270 (N_13270,N_12024,N_12280);
and U13271 (N_13271,N_12805,N_12560);
xor U13272 (N_13272,N_12878,N_12687);
or U13273 (N_13273,N_12121,N_12301);
nand U13274 (N_13274,N_12259,N_12947);
and U13275 (N_13275,N_12883,N_12530);
or U13276 (N_13276,N_12630,N_12986);
nand U13277 (N_13277,N_12131,N_12977);
nor U13278 (N_13278,N_12619,N_12369);
nor U13279 (N_13279,N_12486,N_12439);
and U13280 (N_13280,N_12309,N_12348);
xor U13281 (N_13281,N_12844,N_12493);
nor U13282 (N_13282,N_12218,N_12270);
nor U13283 (N_13283,N_12118,N_12449);
or U13284 (N_13284,N_12081,N_12464);
and U13285 (N_13285,N_12405,N_12199);
or U13286 (N_13286,N_12406,N_12098);
nand U13287 (N_13287,N_12838,N_12214);
nor U13288 (N_13288,N_12350,N_12614);
nor U13289 (N_13289,N_12576,N_12901);
and U13290 (N_13290,N_12420,N_12812);
nor U13291 (N_13291,N_12473,N_12584);
and U13292 (N_13292,N_12513,N_12822);
xor U13293 (N_13293,N_12710,N_12562);
xnor U13294 (N_13294,N_12966,N_12453);
xor U13295 (N_13295,N_12454,N_12568);
nand U13296 (N_13296,N_12926,N_12816);
nor U13297 (N_13297,N_12729,N_12055);
and U13298 (N_13298,N_12828,N_12730);
nand U13299 (N_13299,N_12671,N_12945);
nand U13300 (N_13300,N_12815,N_12427);
nor U13301 (N_13301,N_12559,N_12522);
and U13302 (N_13302,N_12720,N_12709);
nor U13303 (N_13303,N_12396,N_12285);
and U13304 (N_13304,N_12077,N_12074);
or U13305 (N_13305,N_12790,N_12224);
nand U13306 (N_13306,N_12481,N_12600);
and U13307 (N_13307,N_12629,N_12409);
and U13308 (N_13308,N_12778,N_12127);
or U13309 (N_13309,N_12742,N_12446);
and U13310 (N_13310,N_12011,N_12433);
nor U13311 (N_13311,N_12553,N_12036);
xor U13312 (N_13312,N_12059,N_12040);
or U13313 (N_13313,N_12558,N_12087);
nand U13314 (N_13314,N_12126,N_12745);
xor U13315 (N_13315,N_12656,N_12435);
nand U13316 (N_13316,N_12474,N_12107);
xor U13317 (N_13317,N_12279,N_12316);
nor U13318 (N_13318,N_12241,N_12281);
nand U13319 (N_13319,N_12058,N_12363);
xnor U13320 (N_13320,N_12483,N_12697);
nor U13321 (N_13321,N_12547,N_12390);
or U13322 (N_13322,N_12334,N_12543);
and U13323 (N_13323,N_12804,N_12227);
and U13324 (N_13324,N_12902,N_12823);
xor U13325 (N_13325,N_12898,N_12320);
nor U13326 (N_13326,N_12919,N_12376);
xor U13327 (N_13327,N_12383,N_12859);
or U13328 (N_13328,N_12756,N_12506);
nand U13329 (N_13329,N_12631,N_12291);
nand U13330 (N_13330,N_12236,N_12091);
nand U13331 (N_13331,N_12006,N_12083);
nand U13332 (N_13332,N_12803,N_12633);
nor U13333 (N_13333,N_12792,N_12696);
and U13334 (N_13334,N_12873,N_12093);
or U13335 (N_13335,N_12762,N_12501);
nand U13336 (N_13336,N_12677,N_12245);
xnor U13337 (N_13337,N_12089,N_12868);
nand U13338 (N_13338,N_12498,N_12292);
nor U13339 (N_13339,N_12447,N_12981);
and U13340 (N_13340,N_12008,N_12306);
nand U13341 (N_13341,N_12102,N_12353);
or U13342 (N_13342,N_12380,N_12693);
xnor U13343 (N_13343,N_12779,N_12990);
nand U13344 (N_13344,N_12561,N_12863);
or U13345 (N_13345,N_12564,N_12940);
and U13346 (N_13346,N_12797,N_12982);
nor U13347 (N_13347,N_12768,N_12985);
nand U13348 (N_13348,N_12497,N_12428);
nand U13349 (N_13349,N_12890,N_12323);
and U13350 (N_13350,N_12622,N_12313);
and U13351 (N_13351,N_12223,N_12892);
xnor U13352 (N_13352,N_12426,N_12299);
xnor U13353 (N_13353,N_12725,N_12909);
xor U13354 (N_13354,N_12441,N_12893);
nor U13355 (N_13355,N_12820,N_12356);
or U13356 (N_13356,N_12938,N_12960);
or U13357 (N_13357,N_12749,N_12680);
or U13358 (N_13358,N_12371,N_12955);
or U13359 (N_13359,N_12139,N_12106);
xnor U13360 (N_13360,N_12821,N_12239);
xor U13361 (N_13361,N_12575,N_12563);
or U13362 (N_13362,N_12871,N_12840);
nor U13363 (N_13363,N_12088,N_12355);
nor U13364 (N_13364,N_12278,N_12242);
nand U13365 (N_13365,N_12078,N_12243);
and U13366 (N_13366,N_12773,N_12583);
xnor U13367 (N_13367,N_12858,N_12647);
or U13368 (N_13368,N_12734,N_12664);
xnor U13369 (N_13369,N_12099,N_12271);
or U13370 (N_13370,N_12108,N_12176);
and U13371 (N_13371,N_12783,N_12273);
nor U13372 (N_13372,N_12538,N_12086);
or U13373 (N_13373,N_12230,N_12184);
and U13374 (N_13374,N_12574,N_12585);
or U13375 (N_13375,N_12167,N_12542);
nand U13376 (N_13376,N_12286,N_12122);
xnor U13377 (N_13377,N_12284,N_12046);
or U13378 (N_13378,N_12252,N_12963);
nor U13379 (N_13379,N_12701,N_12672);
xnor U13380 (N_13380,N_12691,N_12521);
xor U13381 (N_13381,N_12399,N_12968);
xnor U13382 (N_13382,N_12003,N_12266);
or U13383 (N_13383,N_12641,N_12910);
xnor U13384 (N_13384,N_12714,N_12980);
or U13385 (N_13385,N_12595,N_12111);
nor U13386 (N_13386,N_12774,N_12138);
xor U13387 (N_13387,N_12789,N_12132);
xor U13388 (N_13388,N_12017,N_12237);
and U13389 (N_13389,N_12906,N_12660);
nor U13390 (N_13390,N_12551,N_12514);
and U13391 (N_13391,N_12095,N_12569);
nand U13392 (N_13392,N_12625,N_12013);
nand U13393 (N_13393,N_12688,N_12499);
xor U13394 (N_13394,N_12335,N_12183);
nand U13395 (N_13395,N_12152,N_12148);
xor U13396 (N_13396,N_12200,N_12295);
nand U13397 (N_13397,N_12389,N_12075);
or U13398 (N_13398,N_12332,N_12248);
xor U13399 (N_13399,N_12994,N_12482);
nand U13400 (N_13400,N_12115,N_12953);
nand U13401 (N_13401,N_12719,N_12615);
nor U13402 (N_13402,N_12987,N_12041);
nor U13403 (N_13403,N_12478,N_12459);
nand U13404 (N_13404,N_12070,N_12315);
nand U13405 (N_13405,N_12829,N_12373);
or U13406 (N_13406,N_12667,N_12216);
nand U13407 (N_13407,N_12414,N_12196);
nand U13408 (N_13408,N_12124,N_12755);
nor U13409 (N_13409,N_12763,N_12101);
and U13410 (N_13410,N_12949,N_12596);
and U13411 (N_13411,N_12777,N_12732);
xnor U13412 (N_13412,N_12581,N_12045);
xor U13413 (N_13413,N_12116,N_12096);
xnor U13414 (N_13414,N_12423,N_12848);
or U13415 (N_13415,N_12657,N_12113);
or U13416 (N_13416,N_12669,N_12339);
xnor U13417 (N_13417,N_12590,N_12381);
and U13418 (N_13418,N_12249,N_12432);
xor U13419 (N_13419,N_12646,N_12071);
xnor U13420 (N_13420,N_12050,N_12937);
xnor U13421 (N_13421,N_12260,N_12417);
and U13422 (N_13422,N_12942,N_12480);
nand U13423 (N_13423,N_12517,N_12378);
nand U13424 (N_13424,N_12179,N_12487);
nor U13425 (N_13425,N_12678,N_12764);
or U13426 (N_13426,N_12920,N_12321);
or U13427 (N_13427,N_12347,N_12753);
nand U13428 (N_13428,N_12052,N_12786);
or U13429 (N_13429,N_12345,N_12723);
nor U13430 (N_13430,N_12465,N_12489);
nor U13431 (N_13431,N_12068,N_12896);
xnor U13432 (N_13432,N_12440,N_12958);
nand U13433 (N_13433,N_12967,N_12379);
and U13434 (N_13434,N_12395,N_12638);
xnor U13435 (N_13435,N_12404,N_12652);
and U13436 (N_13436,N_12226,N_12442);
and U13437 (N_13437,N_12048,N_12689);
nand U13438 (N_13438,N_12338,N_12722);
nand U13439 (N_13439,N_12496,N_12133);
nand U13440 (N_13440,N_12085,N_12738);
nor U13441 (N_13441,N_12912,N_12941);
xnor U13442 (N_13442,N_12718,N_12471);
nor U13443 (N_13443,N_12747,N_12038);
or U13444 (N_13444,N_12370,N_12337);
xnor U13445 (N_13445,N_12624,N_12472);
or U13446 (N_13446,N_12387,N_12016);
xnor U13447 (N_13447,N_12651,N_12193);
and U13448 (N_13448,N_12573,N_12996);
nand U13449 (N_13449,N_12843,N_12314);
nand U13450 (N_13450,N_12141,N_12308);
nand U13451 (N_13451,N_12403,N_12004);
or U13452 (N_13452,N_12021,N_12788);
nor U13453 (N_13453,N_12727,N_12037);
or U13454 (N_13454,N_12707,N_12158);
or U13455 (N_13455,N_12419,N_12000);
nand U13456 (N_13456,N_12272,N_12298);
xor U13457 (N_13457,N_12005,N_12190);
and U13458 (N_13458,N_12534,N_12135);
nor U13459 (N_13459,N_12654,N_12712);
or U13460 (N_13460,N_12540,N_12621);
nor U13461 (N_13461,N_12679,N_12051);
and U13462 (N_13462,N_12130,N_12407);
or U13463 (N_13463,N_12479,N_12923);
xnor U13464 (N_13464,N_12027,N_12035);
or U13465 (N_13465,N_12092,N_12469);
or U13466 (N_13466,N_12002,N_12144);
and U13467 (N_13467,N_12007,N_12125);
and U13468 (N_13468,N_12488,N_12076);
nand U13469 (N_13469,N_12137,N_12197);
nand U13470 (N_13470,N_12835,N_12686);
nor U13471 (N_13471,N_12884,N_12872);
and U13472 (N_13472,N_12182,N_12524);
nor U13473 (N_13473,N_12984,N_12205);
nor U13474 (N_13474,N_12993,N_12886);
and U13475 (N_13475,N_12062,N_12528);
nand U13476 (N_13476,N_12238,N_12354);
and U13477 (N_13477,N_12042,N_12222);
nand U13478 (N_13478,N_12895,N_12504);
or U13479 (N_13479,N_12865,N_12203);
or U13480 (N_13480,N_12288,N_12154);
nand U13481 (N_13481,N_12191,N_12939);
nor U13482 (N_13482,N_12831,N_12681);
nor U13483 (N_13483,N_12991,N_12463);
nor U13484 (N_13484,N_12049,N_12146);
nand U13485 (N_13485,N_12793,N_12571);
nand U13486 (N_13486,N_12784,N_12618);
and U13487 (N_13487,N_12799,N_12031);
nand U13488 (N_13488,N_12151,N_12491);
or U13489 (N_13489,N_12388,N_12973);
nand U13490 (N_13490,N_12635,N_12992);
or U13491 (N_13491,N_12698,N_12550);
nand U13492 (N_13492,N_12721,N_12247);
xnor U13493 (N_13493,N_12157,N_12798);
nand U13494 (N_13494,N_12570,N_12975);
and U13495 (N_13495,N_12891,N_12103);
or U13496 (N_13496,N_12194,N_12880);
or U13497 (N_13497,N_12849,N_12673);
nor U13498 (N_13498,N_12979,N_12908);
xnor U13499 (N_13499,N_12185,N_12594);
xor U13500 (N_13500,N_12974,N_12952);
nand U13501 (N_13501,N_12600,N_12126);
or U13502 (N_13502,N_12909,N_12158);
nor U13503 (N_13503,N_12034,N_12272);
nor U13504 (N_13504,N_12029,N_12987);
or U13505 (N_13505,N_12470,N_12933);
and U13506 (N_13506,N_12715,N_12106);
xnor U13507 (N_13507,N_12008,N_12275);
nand U13508 (N_13508,N_12418,N_12011);
nand U13509 (N_13509,N_12138,N_12501);
and U13510 (N_13510,N_12957,N_12747);
xnor U13511 (N_13511,N_12008,N_12748);
xnor U13512 (N_13512,N_12039,N_12230);
nand U13513 (N_13513,N_12680,N_12215);
and U13514 (N_13514,N_12182,N_12597);
and U13515 (N_13515,N_12747,N_12244);
xnor U13516 (N_13516,N_12324,N_12181);
nand U13517 (N_13517,N_12995,N_12610);
xor U13518 (N_13518,N_12569,N_12504);
nand U13519 (N_13519,N_12668,N_12366);
nand U13520 (N_13520,N_12473,N_12770);
and U13521 (N_13521,N_12649,N_12702);
or U13522 (N_13522,N_12875,N_12688);
and U13523 (N_13523,N_12553,N_12215);
xnor U13524 (N_13524,N_12701,N_12029);
xnor U13525 (N_13525,N_12981,N_12307);
nor U13526 (N_13526,N_12494,N_12500);
nor U13527 (N_13527,N_12292,N_12976);
nand U13528 (N_13528,N_12134,N_12119);
and U13529 (N_13529,N_12303,N_12649);
nor U13530 (N_13530,N_12174,N_12692);
and U13531 (N_13531,N_12328,N_12453);
or U13532 (N_13532,N_12022,N_12977);
xor U13533 (N_13533,N_12140,N_12667);
nor U13534 (N_13534,N_12190,N_12156);
and U13535 (N_13535,N_12771,N_12234);
and U13536 (N_13536,N_12237,N_12978);
and U13537 (N_13537,N_12362,N_12130);
or U13538 (N_13538,N_12888,N_12422);
xnor U13539 (N_13539,N_12583,N_12528);
and U13540 (N_13540,N_12387,N_12499);
or U13541 (N_13541,N_12731,N_12805);
and U13542 (N_13542,N_12246,N_12792);
or U13543 (N_13543,N_12046,N_12009);
nor U13544 (N_13544,N_12287,N_12316);
or U13545 (N_13545,N_12961,N_12627);
or U13546 (N_13546,N_12385,N_12896);
nor U13547 (N_13547,N_12125,N_12946);
and U13548 (N_13548,N_12667,N_12417);
xor U13549 (N_13549,N_12145,N_12559);
xor U13550 (N_13550,N_12156,N_12333);
or U13551 (N_13551,N_12051,N_12219);
and U13552 (N_13552,N_12491,N_12674);
and U13553 (N_13553,N_12067,N_12485);
nand U13554 (N_13554,N_12292,N_12913);
xnor U13555 (N_13555,N_12741,N_12369);
or U13556 (N_13556,N_12229,N_12984);
or U13557 (N_13557,N_12698,N_12795);
nor U13558 (N_13558,N_12485,N_12010);
nand U13559 (N_13559,N_12665,N_12562);
nor U13560 (N_13560,N_12826,N_12895);
or U13561 (N_13561,N_12425,N_12406);
and U13562 (N_13562,N_12254,N_12601);
or U13563 (N_13563,N_12257,N_12541);
nor U13564 (N_13564,N_12232,N_12659);
and U13565 (N_13565,N_12598,N_12190);
nand U13566 (N_13566,N_12464,N_12782);
and U13567 (N_13567,N_12287,N_12921);
and U13568 (N_13568,N_12145,N_12966);
nor U13569 (N_13569,N_12486,N_12357);
nand U13570 (N_13570,N_12163,N_12333);
or U13571 (N_13571,N_12412,N_12674);
and U13572 (N_13572,N_12632,N_12922);
nand U13573 (N_13573,N_12552,N_12788);
xnor U13574 (N_13574,N_12659,N_12899);
nor U13575 (N_13575,N_12330,N_12264);
nand U13576 (N_13576,N_12723,N_12761);
and U13577 (N_13577,N_12688,N_12817);
or U13578 (N_13578,N_12909,N_12385);
or U13579 (N_13579,N_12234,N_12031);
nor U13580 (N_13580,N_12817,N_12691);
nor U13581 (N_13581,N_12138,N_12654);
or U13582 (N_13582,N_12521,N_12339);
and U13583 (N_13583,N_12238,N_12887);
xnor U13584 (N_13584,N_12163,N_12592);
xnor U13585 (N_13585,N_12763,N_12888);
xnor U13586 (N_13586,N_12967,N_12784);
and U13587 (N_13587,N_12611,N_12716);
nor U13588 (N_13588,N_12623,N_12062);
xnor U13589 (N_13589,N_12971,N_12960);
nand U13590 (N_13590,N_12788,N_12456);
and U13591 (N_13591,N_12709,N_12649);
or U13592 (N_13592,N_12369,N_12425);
xnor U13593 (N_13593,N_12696,N_12153);
xnor U13594 (N_13594,N_12538,N_12362);
and U13595 (N_13595,N_12975,N_12323);
and U13596 (N_13596,N_12759,N_12402);
and U13597 (N_13597,N_12673,N_12667);
nand U13598 (N_13598,N_12998,N_12330);
nor U13599 (N_13599,N_12487,N_12306);
xnor U13600 (N_13600,N_12446,N_12390);
and U13601 (N_13601,N_12146,N_12942);
xor U13602 (N_13602,N_12963,N_12303);
or U13603 (N_13603,N_12103,N_12893);
nor U13604 (N_13604,N_12969,N_12417);
and U13605 (N_13605,N_12121,N_12574);
nor U13606 (N_13606,N_12243,N_12638);
or U13607 (N_13607,N_12985,N_12108);
nand U13608 (N_13608,N_12092,N_12361);
xnor U13609 (N_13609,N_12152,N_12244);
or U13610 (N_13610,N_12583,N_12307);
and U13611 (N_13611,N_12476,N_12842);
nand U13612 (N_13612,N_12679,N_12267);
or U13613 (N_13613,N_12342,N_12433);
and U13614 (N_13614,N_12156,N_12748);
or U13615 (N_13615,N_12975,N_12982);
nand U13616 (N_13616,N_12879,N_12385);
xnor U13617 (N_13617,N_12197,N_12254);
and U13618 (N_13618,N_12599,N_12721);
nor U13619 (N_13619,N_12547,N_12640);
nand U13620 (N_13620,N_12029,N_12631);
nor U13621 (N_13621,N_12168,N_12255);
xnor U13622 (N_13622,N_12105,N_12899);
or U13623 (N_13623,N_12432,N_12699);
or U13624 (N_13624,N_12542,N_12435);
or U13625 (N_13625,N_12996,N_12627);
or U13626 (N_13626,N_12499,N_12069);
nand U13627 (N_13627,N_12930,N_12733);
xor U13628 (N_13628,N_12929,N_12514);
and U13629 (N_13629,N_12567,N_12103);
and U13630 (N_13630,N_12446,N_12245);
or U13631 (N_13631,N_12190,N_12519);
and U13632 (N_13632,N_12309,N_12295);
xor U13633 (N_13633,N_12582,N_12210);
and U13634 (N_13634,N_12031,N_12870);
and U13635 (N_13635,N_12639,N_12185);
and U13636 (N_13636,N_12542,N_12751);
xor U13637 (N_13637,N_12973,N_12679);
xor U13638 (N_13638,N_12123,N_12718);
nor U13639 (N_13639,N_12352,N_12776);
xor U13640 (N_13640,N_12770,N_12749);
xor U13641 (N_13641,N_12854,N_12044);
xor U13642 (N_13642,N_12476,N_12984);
nor U13643 (N_13643,N_12087,N_12219);
nor U13644 (N_13644,N_12693,N_12630);
nor U13645 (N_13645,N_12094,N_12345);
nand U13646 (N_13646,N_12840,N_12638);
and U13647 (N_13647,N_12554,N_12180);
xnor U13648 (N_13648,N_12167,N_12287);
nand U13649 (N_13649,N_12390,N_12380);
and U13650 (N_13650,N_12985,N_12172);
or U13651 (N_13651,N_12747,N_12349);
nor U13652 (N_13652,N_12741,N_12349);
nand U13653 (N_13653,N_12088,N_12798);
or U13654 (N_13654,N_12927,N_12647);
nand U13655 (N_13655,N_12155,N_12554);
nor U13656 (N_13656,N_12475,N_12658);
nand U13657 (N_13657,N_12739,N_12865);
and U13658 (N_13658,N_12874,N_12563);
or U13659 (N_13659,N_12267,N_12248);
xor U13660 (N_13660,N_12841,N_12757);
xnor U13661 (N_13661,N_12281,N_12271);
nor U13662 (N_13662,N_12355,N_12758);
nor U13663 (N_13663,N_12982,N_12183);
nor U13664 (N_13664,N_12331,N_12566);
xnor U13665 (N_13665,N_12379,N_12490);
nor U13666 (N_13666,N_12204,N_12175);
nand U13667 (N_13667,N_12051,N_12283);
xor U13668 (N_13668,N_12386,N_12729);
nor U13669 (N_13669,N_12063,N_12623);
nand U13670 (N_13670,N_12442,N_12669);
nand U13671 (N_13671,N_12413,N_12604);
nor U13672 (N_13672,N_12080,N_12040);
nor U13673 (N_13673,N_12539,N_12583);
nand U13674 (N_13674,N_12359,N_12087);
xor U13675 (N_13675,N_12563,N_12627);
nor U13676 (N_13676,N_12928,N_12986);
xnor U13677 (N_13677,N_12858,N_12130);
or U13678 (N_13678,N_12758,N_12892);
and U13679 (N_13679,N_12134,N_12450);
nor U13680 (N_13680,N_12021,N_12276);
nand U13681 (N_13681,N_12427,N_12732);
nor U13682 (N_13682,N_12877,N_12085);
and U13683 (N_13683,N_12144,N_12694);
nor U13684 (N_13684,N_12591,N_12461);
nand U13685 (N_13685,N_12940,N_12840);
nor U13686 (N_13686,N_12462,N_12690);
xor U13687 (N_13687,N_12143,N_12255);
and U13688 (N_13688,N_12094,N_12350);
or U13689 (N_13689,N_12597,N_12446);
xor U13690 (N_13690,N_12382,N_12136);
and U13691 (N_13691,N_12256,N_12051);
and U13692 (N_13692,N_12921,N_12680);
nor U13693 (N_13693,N_12869,N_12582);
nand U13694 (N_13694,N_12049,N_12837);
or U13695 (N_13695,N_12048,N_12598);
and U13696 (N_13696,N_12186,N_12628);
nand U13697 (N_13697,N_12395,N_12145);
nor U13698 (N_13698,N_12926,N_12326);
and U13699 (N_13699,N_12576,N_12764);
or U13700 (N_13700,N_12578,N_12690);
nand U13701 (N_13701,N_12881,N_12819);
xnor U13702 (N_13702,N_12925,N_12326);
and U13703 (N_13703,N_12150,N_12781);
or U13704 (N_13704,N_12569,N_12747);
and U13705 (N_13705,N_12311,N_12677);
xnor U13706 (N_13706,N_12348,N_12593);
xnor U13707 (N_13707,N_12439,N_12813);
nor U13708 (N_13708,N_12292,N_12579);
and U13709 (N_13709,N_12280,N_12584);
nor U13710 (N_13710,N_12908,N_12627);
or U13711 (N_13711,N_12136,N_12981);
xnor U13712 (N_13712,N_12476,N_12629);
or U13713 (N_13713,N_12987,N_12780);
nand U13714 (N_13714,N_12771,N_12530);
xor U13715 (N_13715,N_12762,N_12006);
or U13716 (N_13716,N_12609,N_12969);
and U13717 (N_13717,N_12960,N_12252);
nor U13718 (N_13718,N_12631,N_12526);
xnor U13719 (N_13719,N_12355,N_12502);
or U13720 (N_13720,N_12282,N_12211);
nand U13721 (N_13721,N_12435,N_12672);
nor U13722 (N_13722,N_12716,N_12753);
nor U13723 (N_13723,N_12050,N_12636);
nand U13724 (N_13724,N_12449,N_12765);
or U13725 (N_13725,N_12269,N_12495);
xor U13726 (N_13726,N_12033,N_12751);
or U13727 (N_13727,N_12645,N_12957);
nor U13728 (N_13728,N_12958,N_12025);
xor U13729 (N_13729,N_12431,N_12782);
nand U13730 (N_13730,N_12858,N_12172);
and U13731 (N_13731,N_12012,N_12782);
or U13732 (N_13732,N_12804,N_12130);
xor U13733 (N_13733,N_12289,N_12244);
nand U13734 (N_13734,N_12053,N_12737);
and U13735 (N_13735,N_12658,N_12651);
or U13736 (N_13736,N_12436,N_12283);
xnor U13737 (N_13737,N_12823,N_12216);
nor U13738 (N_13738,N_12704,N_12202);
nand U13739 (N_13739,N_12021,N_12054);
nor U13740 (N_13740,N_12977,N_12477);
or U13741 (N_13741,N_12681,N_12859);
nor U13742 (N_13742,N_12975,N_12475);
nand U13743 (N_13743,N_12599,N_12647);
and U13744 (N_13744,N_12075,N_12273);
xor U13745 (N_13745,N_12070,N_12005);
nor U13746 (N_13746,N_12036,N_12715);
or U13747 (N_13747,N_12967,N_12328);
xor U13748 (N_13748,N_12497,N_12464);
and U13749 (N_13749,N_12935,N_12165);
xnor U13750 (N_13750,N_12672,N_12137);
xor U13751 (N_13751,N_12587,N_12211);
nand U13752 (N_13752,N_12112,N_12236);
or U13753 (N_13753,N_12186,N_12537);
or U13754 (N_13754,N_12034,N_12432);
and U13755 (N_13755,N_12382,N_12729);
xnor U13756 (N_13756,N_12857,N_12455);
and U13757 (N_13757,N_12699,N_12430);
or U13758 (N_13758,N_12131,N_12749);
and U13759 (N_13759,N_12482,N_12794);
nor U13760 (N_13760,N_12107,N_12368);
and U13761 (N_13761,N_12289,N_12524);
and U13762 (N_13762,N_12509,N_12607);
or U13763 (N_13763,N_12607,N_12237);
and U13764 (N_13764,N_12260,N_12361);
nor U13765 (N_13765,N_12389,N_12871);
and U13766 (N_13766,N_12136,N_12896);
xor U13767 (N_13767,N_12625,N_12431);
nand U13768 (N_13768,N_12266,N_12770);
or U13769 (N_13769,N_12491,N_12853);
and U13770 (N_13770,N_12488,N_12657);
xnor U13771 (N_13771,N_12343,N_12254);
nor U13772 (N_13772,N_12761,N_12116);
xor U13773 (N_13773,N_12774,N_12400);
xor U13774 (N_13774,N_12144,N_12403);
nand U13775 (N_13775,N_12909,N_12436);
nor U13776 (N_13776,N_12302,N_12543);
and U13777 (N_13777,N_12631,N_12762);
nor U13778 (N_13778,N_12164,N_12612);
xnor U13779 (N_13779,N_12337,N_12612);
xor U13780 (N_13780,N_12212,N_12152);
and U13781 (N_13781,N_12289,N_12657);
nand U13782 (N_13782,N_12282,N_12549);
or U13783 (N_13783,N_12293,N_12463);
or U13784 (N_13784,N_12223,N_12962);
xnor U13785 (N_13785,N_12053,N_12202);
and U13786 (N_13786,N_12728,N_12212);
nor U13787 (N_13787,N_12062,N_12742);
xor U13788 (N_13788,N_12730,N_12582);
nand U13789 (N_13789,N_12765,N_12174);
and U13790 (N_13790,N_12903,N_12820);
or U13791 (N_13791,N_12145,N_12396);
nor U13792 (N_13792,N_12934,N_12088);
and U13793 (N_13793,N_12346,N_12525);
or U13794 (N_13794,N_12937,N_12248);
nand U13795 (N_13795,N_12978,N_12281);
nand U13796 (N_13796,N_12397,N_12796);
xnor U13797 (N_13797,N_12453,N_12947);
nand U13798 (N_13798,N_12400,N_12320);
xnor U13799 (N_13799,N_12351,N_12934);
and U13800 (N_13800,N_12145,N_12306);
nor U13801 (N_13801,N_12875,N_12862);
and U13802 (N_13802,N_12596,N_12601);
or U13803 (N_13803,N_12326,N_12757);
nor U13804 (N_13804,N_12344,N_12618);
nand U13805 (N_13805,N_12769,N_12545);
xnor U13806 (N_13806,N_12231,N_12045);
or U13807 (N_13807,N_12686,N_12400);
or U13808 (N_13808,N_12798,N_12665);
and U13809 (N_13809,N_12164,N_12161);
and U13810 (N_13810,N_12793,N_12899);
nor U13811 (N_13811,N_12288,N_12929);
and U13812 (N_13812,N_12905,N_12158);
and U13813 (N_13813,N_12456,N_12568);
or U13814 (N_13814,N_12867,N_12574);
nor U13815 (N_13815,N_12023,N_12646);
nand U13816 (N_13816,N_12493,N_12391);
xor U13817 (N_13817,N_12790,N_12620);
xnor U13818 (N_13818,N_12824,N_12640);
nand U13819 (N_13819,N_12541,N_12965);
or U13820 (N_13820,N_12291,N_12988);
and U13821 (N_13821,N_12190,N_12907);
xor U13822 (N_13822,N_12240,N_12746);
nor U13823 (N_13823,N_12583,N_12219);
or U13824 (N_13824,N_12572,N_12028);
and U13825 (N_13825,N_12955,N_12820);
nor U13826 (N_13826,N_12649,N_12004);
xor U13827 (N_13827,N_12438,N_12927);
xnor U13828 (N_13828,N_12117,N_12819);
or U13829 (N_13829,N_12790,N_12849);
or U13830 (N_13830,N_12450,N_12089);
nor U13831 (N_13831,N_12897,N_12079);
xor U13832 (N_13832,N_12239,N_12534);
nor U13833 (N_13833,N_12379,N_12003);
nor U13834 (N_13834,N_12056,N_12504);
xor U13835 (N_13835,N_12141,N_12526);
and U13836 (N_13836,N_12341,N_12296);
or U13837 (N_13837,N_12449,N_12592);
nand U13838 (N_13838,N_12388,N_12306);
xor U13839 (N_13839,N_12634,N_12543);
or U13840 (N_13840,N_12837,N_12141);
nand U13841 (N_13841,N_12836,N_12736);
xor U13842 (N_13842,N_12425,N_12230);
xnor U13843 (N_13843,N_12100,N_12991);
and U13844 (N_13844,N_12889,N_12319);
nand U13845 (N_13845,N_12253,N_12716);
or U13846 (N_13846,N_12025,N_12705);
nor U13847 (N_13847,N_12347,N_12018);
nor U13848 (N_13848,N_12060,N_12521);
nand U13849 (N_13849,N_12571,N_12117);
or U13850 (N_13850,N_12152,N_12758);
or U13851 (N_13851,N_12776,N_12242);
xor U13852 (N_13852,N_12579,N_12897);
nand U13853 (N_13853,N_12889,N_12293);
and U13854 (N_13854,N_12310,N_12019);
nor U13855 (N_13855,N_12992,N_12616);
and U13856 (N_13856,N_12539,N_12683);
or U13857 (N_13857,N_12191,N_12677);
or U13858 (N_13858,N_12929,N_12387);
and U13859 (N_13859,N_12230,N_12075);
nor U13860 (N_13860,N_12208,N_12128);
nand U13861 (N_13861,N_12756,N_12848);
xnor U13862 (N_13862,N_12207,N_12010);
xor U13863 (N_13863,N_12949,N_12726);
nand U13864 (N_13864,N_12103,N_12377);
nor U13865 (N_13865,N_12778,N_12091);
or U13866 (N_13866,N_12441,N_12034);
and U13867 (N_13867,N_12626,N_12519);
nor U13868 (N_13868,N_12107,N_12437);
nor U13869 (N_13869,N_12418,N_12408);
nor U13870 (N_13870,N_12722,N_12246);
nand U13871 (N_13871,N_12225,N_12333);
nand U13872 (N_13872,N_12563,N_12569);
xnor U13873 (N_13873,N_12470,N_12556);
nor U13874 (N_13874,N_12245,N_12127);
nand U13875 (N_13875,N_12546,N_12363);
nand U13876 (N_13876,N_12655,N_12591);
and U13877 (N_13877,N_12566,N_12014);
xnor U13878 (N_13878,N_12074,N_12860);
xor U13879 (N_13879,N_12841,N_12861);
and U13880 (N_13880,N_12506,N_12982);
nand U13881 (N_13881,N_12819,N_12266);
nand U13882 (N_13882,N_12610,N_12400);
or U13883 (N_13883,N_12071,N_12611);
or U13884 (N_13884,N_12953,N_12449);
or U13885 (N_13885,N_12241,N_12772);
nor U13886 (N_13886,N_12882,N_12608);
nor U13887 (N_13887,N_12754,N_12202);
nand U13888 (N_13888,N_12971,N_12745);
and U13889 (N_13889,N_12718,N_12715);
and U13890 (N_13890,N_12438,N_12777);
or U13891 (N_13891,N_12792,N_12897);
or U13892 (N_13892,N_12424,N_12176);
and U13893 (N_13893,N_12803,N_12915);
or U13894 (N_13894,N_12169,N_12173);
or U13895 (N_13895,N_12135,N_12760);
nand U13896 (N_13896,N_12536,N_12973);
and U13897 (N_13897,N_12062,N_12357);
nor U13898 (N_13898,N_12589,N_12140);
xor U13899 (N_13899,N_12276,N_12300);
or U13900 (N_13900,N_12922,N_12927);
nor U13901 (N_13901,N_12559,N_12076);
nand U13902 (N_13902,N_12630,N_12205);
nand U13903 (N_13903,N_12523,N_12473);
nand U13904 (N_13904,N_12418,N_12401);
xnor U13905 (N_13905,N_12523,N_12213);
and U13906 (N_13906,N_12227,N_12695);
or U13907 (N_13907,N_12276,N_12214);
nand U13908 (N_13908,N_12629,N_12348);
xnor U13909 (N_13909,N_12752,N_12478);
and U13910 (N_13910,N_12281,N_12114);
nand U13911 (N_13911,N_12627,N_12168);
xnor U13912 (N_13912,N_12794,N_12711);
nor U13913 (N_13913,N_12916,N_12150);
nor U13914 (N_13914,N_12016,N_12694);
nand U13915 (N_13915,N_12816,N_12075);
and U13916 (N_13916,N_12924,N_12552);
or U13917 (N_13917,N_12786,N_12554);
and U13918 (N_13918,N_12847,N_12587);
or U13919 (N_13919,N_12383,N_12845);
nand U13920 (N_13920,N_12676,N_12525);
or U13921 (N_13921,N_12567,N_12380);
nor U13922 (N_13922,N_12909,N_12591);
nand U13923 (N_13923,N_12546,N_12926);
nand U13924 (N_13924,N_12661,N_12691);
or U13925 (N_13925,N_12267,N_12608);
nor U13926 (N_13926,N_12302,N_12871);
or U13927 (N_13927,N_12445,N_12734);
nor U13928 (N_13928,N_12616,N_12470);
xnor U13929 (N_13929,N_12187,N_12315);
nor U13930 (N_13930,N_12219,N_12602);
and U13931 (N_13931,N_12657,N_12812);
xor U13932 (N_13932,N_12361,N_12704);
xnor U13933 (N_13933,N_12924,N_12496);
nor U13934 (N_13934,N_12637,N_12936);
xnor U13935 (N_13935,N_12527,N_12062);
nand U13936 (N_13936,N_12691,N_12766);
and U13937 (N_13937,N_12468,N_12395);
xnor U13938 (N_13938,N_12415,N_12538);
or U13939 (N_13939,N_12126,N_12581);
nor U13940 (N_13940,N_12220,N_12350);
and U13941 (N_13941,N_12492,N_12336);
or U13942 (N_13942,N_12740,N_12415);
xnor U13943 (N_13943,N_12427,N_12669);
xor U13944 (N_13944,N_12375,N_12562);
nand U13945 (N_13945,N_12515,N_12810);
xnor U13946 (N_13946,N_12235,N_12035);
nor U13947 (N_13947,N_12583,N_12408);
nand U13948 (N_13948,N_12925,N_12528);
nor U13949 (N_13949,N_12222,N_12865);
nor U13950 (N_13950,N_12441,N_12987);
or U13951 (N_13951,N_12966,N_12669);
xor U13952 (N_13952,N_12092,N_12071);
or U13953 (N_13953,N_12241,N_12875);
xor U13954 (N_13954,N_12328,N_12908);
nor U13955 (N_13955,N_12215,N_12538);
or U13956 (N_13956,N_12729,N_12475);
xnor U13957 (N_13957,N_12219,N_12307);
nand U13958 (N_13958,N_12493,N_12191);
xor U13959 (N_13959,N_12478,N_12123);
xor U13960 (N_13960,N_12351,N_12738);
nor U13961 (N_13961,N_12808,N_12237);
or U13962 (N_13962,N_12549,N_12026);
xnor U13963 (N_13963,N_12725,N_12066);
or U13964 (N_13964,N_12768,N_12001);
xnor U13965 (N_13965,N_12870,N_12401);
xor U13966 (N_13966,N_12090,N_12300);
and U13967 (N_13967,N_12301,N_12848);
nand U13968 (N_13968,N_12683,N_12869);
or U13969 (N_13969,N_12147,N_12781);
nor U13970 (N_13970,N_12014,N_12792);
or U13971 (N_13971,N_12458,N_12971);
xnor U13972 (N_13972,N_12220,N_12957);
or U13973 (N_13973,N_12563,N_12118);
xor U13974 (N_13974,N_12371,N_12824);
or U13975 (N_13975,N_12922,N_12061);
or U13976 (N_13976,N_12295,N_12795);
or U13977 (N_13977,N_12472,N_12543);
or U13978 (N_13978,N_12111,N_12656);
or U13979 (N_13979,N_12647,N_12759);
xor U13980 (N_13980,N_12275,N_12043);
nor U13981 (N_13981,N_12082,N_12272);
xnor U13982 (N_13982,N_12464,N_12390);
or U13983 (N_13983,N_12962,N_12805);
xor U13984 (N_13984,N_12124,N_12237);
or U13985 (N_13985,N_12563,N_12195);
nor U13986 (N_13986,N_12500,N_12052);
or U13987 (N_13987,N_12883,N_12046);
nand U13988 (N_13988,N_12861,N_12152);
or U13989 (N_13989,N_12608,N_12891);
and U13990 (N_13990,N_12462,N_12578);
or U13991 (N_13991,N_12251,N_12424);
xor U13992 (N_13992,N_12628,N_12964);
nand U13993 (N_13993,N_12267,N_12297);
xnor U13994 (N_13994,N_12983,N_12369);
and U13995 (N_13995,N_12369,N_12090);
nand U13996 (N_13996,N_12129,N_12412);
and U13997 (N_13997,N_12856,N_12102);
nor U13998 (N_13998,N_12578,N_12788);
nor U13999 (N_13999,N_12118,N_12042);
and U14000 (N_14000,N_13405,N_13624);
xor U14001 (N_14001,N_13814,N_13218);
and U14002 (N_14002,N_13102,N_13398);
nor U14003 (N_14003,N_13255,N_13902);
and U14004 (N_14004,N_13990,N_13812);
and U14005 (N_14005,N_13552,N_13256);
nor U14006 (N_14006,N_13784,N_13728);
xnor U14007 (N_14007,N_13300,N_13030);
or U14008 (N_14008,N_13717,N_13440);
nand U14009 (N_14009,N_13925,N_13937);
nor U14010 (N_14010,N_13198,N_13646);
and U14011 (N_14011,N_13779,N_13827);
or U14012 (N_14012,N_13560,N_13819);
and U14013 (N_14013,N_13244,N_13838);
nor U14014 (N_14014,N_13752,N_13631);
nand U14015 (N_14015,N_13714,N_13417);
and U14016 (N_14016,N_13229,N_13416);
nor U14017 (N_14017,N_13315,N_13150);
nor U14018 (N_14018,N_13588,N_13831);
and U14019 (N_14019,N_13343,N_13359);
and U14020 (N_14020,N_13409,N_13032);
nand U14021 (N_14021,N_13329,N_13679);
and U14022 (N_14022,N_13822,N_13780);
xnor U14023 (N_14023,N_13133,N_13605);
xnor U14024 (N_14024,N_13017,N_13651);
and U14025 (N_14025,N_13104,N_13850);
or U14026 (N_14026,N_13788,N_13458);
nand U14027 (N_14027,N_13490,N_13826);
nor U14028 (N_14028,N_13573,N_13285);
or U14029 (N_14029,N_13834,N_13567);
or U14030 (N_14030,N_13432,N_13634);
xnor U14031 (N_14031,N_13092,N_13845);
nor U14032 (N_14032,N_13393,N_13379);
nor U14033 (N_14033,N_13557,N_13371);
or U14034 (N_14034,N_13574,N_13444);
or U14035 (N_14035,N_13114,N_13389);
xor U14036 (N_14036,N_13586,N_13072);
xor U14037 (N_14037,N_13709,N_13337);
nor U14038 (N_14038,N_13543,N_13145);
xnor U14039 (N_14039,N_13601,N_13074);
nand U14040 (N_14040,N_13140,N_13429);
nor U14041 (N_14041,N_13487,N_13418);
xnor U14042 (N_14042,N_13587,N_13642);
or U14043 (N_14043,N_13493,N_13810);
or U14044 (N_14044,N_13469,N_13043);
nor U14045 (N_14045,N_13233,N_13764);
xnor U14046 (N_14046,N_13719,N_13744);
nand U14047 (N_14047,N_13356,N_13823);
or U14048 (N_14048,N_13217,N_13886);
and U14049 (N_14049,N_13540,N_13962);
nand U14050 (N_14050,N_13852,N_13840);
and U14051 (N_14051,N_13210,N_13473);
nand U14052 (N_14052,N_13112,N_13097);
nand U14053 (N_14053,N_13530,N_13245);
nor U14054 (N_14054,N_13282,N_13946);
and U14055 (N_14055,N_13160,N_13996);
or U14056 (N_14056,N_13724,N_13031);
xnor U14057 (N_14057,N_13848,N_13449);
xor U14058 (N_14058,N_13873,N_13686);
and U14059 (N_14059,N_13038,N_13224);
or U14060 (N_14060,N_13524,N_13802);
or U14061 (N_14061,N_13123,N_13690);
and U14062 (N_14062,N_13190,N_13638);
and U14063 (N_14063,N_13309,N_13931);
xor U14064 (N_14064,N_13240,N_13948);
and U14065 (N_14065,N_13563,N_13428);
xor U14066 (N_14066,N_13051,N_13893);
and U14067 (N_14067,N_13101,N_13766);
and U14068 (N_14068,N_13919,N_13743);
and U14069 (N_14069,N_13018,N_13555);
xnor U14070 (N_14070,N_13325,N_13580);
nor U14071 (N_14071,N_13401,N_13556);
nand U14072 (N_14072,N_13126,N_13078);
nor U14073 (N_14073,N_13130,N_13363);
and U14074 (N_14074,N_13507,N_13547);
xnor U14075 (N_14075,N_13169,N_13159);
nor U14076 (N_14076,N_13212,N_13463);
nand U14077 (N_14077,N_13495,N_13526);
xor U14078 (N_14078,N_13163,N_13375);
or U14079 (N_14079,N_13773,N_13386);
nand U14080 (N_14080,N_13600,N_13307);
and U14081 (N_14081,N_13277,N_13414);
nand U14082 (N_14082,N_13022,N_13564);
nand U14083 (N_14083,N_13331,N_13930);
nand U14084 (N_14084,N_13790,N_13041);
nor U14085 (N_14085,N_13312,N_13305);
xor U14086 (N_14086,N_13462,N_13774);
xnor U14087 (N_14087,N_13747,N_13756);
nand U14088 (N_14088,N_13448,N_13647);
or U14089 (N_14089,N_13966,N_13640);
nand U14090 (N_14090,N_13385,N_13185);
xor U14091 (N_14091,N_13954,N_13980);
nand U14092 (N_14092,N_13945,N_13614);
nor U14093 (N_14093,N_13258,N_13820);
or U14094 (N_14094,N_13734,N_13311);
xor U14095 (N_14095,N_13982,N_13914);
xnor U14096 (N_14096,N_13264,N_13194);
xnor U14097 (N_14097,N_13942,N_13815);
nand U14098 (N_14098,N_13003,N_13099);
xnor U14099 (N_14099,N_13085,N_13967);
nor U14100 (N_14100,N_13167,N_13915);
or U14101 (N_14101,N_13299,N_13770);
nor U14102 (N_14102,N_13147,N_13139);
and U14103 (N_14103,N_13377,N_13518);
xnor U14104 (N_14104,N_13116,N_13857);
xnor U14105 (N_14105,N_13583,N_13204);
or U14106 (N_14106,N_13579,N_13122);
nand U14107 (N_14107,N_13777,N_13090);
nor U14108 (N_14108,N_13173,N_13411);
and U14109 (N_14109,N_13232,N_13381);
or U14110 (N_14110,N_13438,N_13510);
nand U14111 (N_14111,N_13986,N_13738);
or U14112 (N_14112,N_13193,N_13981);
or U14113 (N_14113,N_13464,N_13641);
nand U14114 (N_14114,N_13644,N_13711);
xor U14115 (N_14115,N_13228,N_13636);
xnor U14116 (N_14116,N_13720,N_13682);
and U14117 (N_14117,N_13266,N_13175);
nor U14118 (N_14118,N_13094,N_13191);
nand U14119 (N_14119,N_13816,N_13751);
nor U14120 (N_14120,N_13082,N_13357);
and U14121 (N_14121,N_13007,N_13786);
and U14122 (N_14122,N_13885,N_13800);
xnor U14123 (N_14123,N_13361,N_13909);
or U14124 (N_14124,N_13179,N_13327);
xnor U14125 (N_14125,N_13408,N_13271);
and U14126 (N_14126,N_13853,N_13799);
and U14127 (N_14127,N_13161,N_13792);
and U14128 (N_14128,N_13274,N_13538);
nor U14129 (N_14129,N_13685,N_13154);
xnor U14130 (N_14130,N_13058,N_13241);
nand U14131 (N_14131,N_13451,N_13506);
xor U14132 (N_14132,N_13195,N_13333);
or U14133 (N_14133,N_13248,N_13671);
nand U14134 (N_14134,N_13054,N_13984);
xor U14135 (N_14135,N_13750,N_13913);
and U14136 (N_14136,N_13172,N_13301);
nand U14137 (N_14137,N_13297,N_13721);
or U14138 (N_14138,N_13177,N_13550);
xor U14139 (N_14139,N_13753,N_13716);
xor U14140 (N_14140,N_13863,N_13358);
nor U14141 (N_14141,N_13968,N_13924);
xor U14142 (N_14142,N_13960,N_13339);
or U14143 (N_14143,N_13544,N_13424);
xnor U14144 (N_14144,N_13267,N_13000);
xnor U14145 (N_14145,N_13045,N_13211);
nand U14146 (N_14146,N_13652,N_13088);
nand U14147 (N_14147,N_13137,N_13558);
nand U14148 (N_14148,N_13336,N_13594);
nand U14149 (N_14149,N_13283,N_13119);
nand U14150 (N_14150,N_13070,N_13459);
nor U14151 (N_14151,N_13132,N_13349);
nor U14152 (N_14152,N_13434,N_13355);
or U14153 (N_14153,N_13667,N_13015);
or U14154 (N_14154,N_13795,N_13578);
nand U14155 (N_14155,N_13370,N_13425);
nor U14156 (N_14156,N_13781,N_13055);
or U14157 (N_14157,N_13040,N_13561);
and U14158 (N_14158,N_13403,N_13707);
nor U14159 (N_14159,N_13236,N_13235);
xor U14160 (N_14160,N_13596,N_13471);
nor U14161 (N_14161,N_13142,N_13771);
nor U14162 (N_14162,N_13314,N_13859);
or U14163 (N_14163,N_13860,N_13376);
and U14164 (N_14164,N_13263,N_13659);
xnor U14165 (N_14165,N_13275,N_13303);
or U14166 (N_14166,N_13033,N_13197);
xor U14167 (N_14167,N_13323,N_13608);
nor U14168 (N_14168,N_13854,N_13681);
xor U14169 (N_14169,N_13989,N_13821);
nand U14170 (N_14170,N_13320,N_13519);
nand U14171 (N_14171,N_13988,N_13949);
nand U14172 (N_14172,N_13192,N_13882);
nand U14173 (N_14173,N_13353,N_13202);
nand U14174 (N_14174,N_13562,N_13662);
nand U14175 (N_14175,N_13023,N_13864);
and U14176 (N_14176,N_13061,N_13699);
nor U14177 (N_14177,N_13247,N_13618);
or U14178 (N_14178,N_13991,N_13598);
nor U14179 (N_14179,N_13551,N_13566);
nand U14180 (N_14180,N_13899,N_13318);
and U14181 (N_14181,N_13936,N_13665);
nor U14182 (N_14182,N_13835,N_13604);
nand U14183 (N_14183,N_13021,N_13250);
or U14184 (N_14184,N_13892,N_13654);
nand U14185 (N_14185,N_13461,N_13929);
and U14186 (N_14186,N_13328,N_13528);
xor U14187 (N_14187,N_13502,N_13725);
nor U14188 (N_14188,N_13867,N_13687);
or U14189 (N_14189,N_13481,N_13941);
xnor U14190 (N_14190,N_13014,N_13237);
or U14191 (N_14191,N_13599,N_13215);
nor U14192 (N_14192,N_13581,N_13657);
nor U14193 (N_14193,N_13384,N_13158);
and U14194 (N_14194,N_13152,N_13399);
and U14195 (N_14195,N_13829,N_13998);
or U14196 (N_14196,N_13727,N_13365);
xor U14197 (N_14197,N_13019,N_13900);
nand U14198 (N_14198,N_13674,N_13201);
nand U14199 (N_14199,N_13862,N_13520);
or U14200 (N_14200,N_13071,N_13171);
xor U14201 (N_14201,N_13317,N_13778);
xor U14202 (N_14202,N_13024,N_13109);
or U14203 (N_14203,N_13722,N_13541);
xor U14204 (N_14204,N_13239,N_13073);
nor U14205 (N_14205,N_13304,N_13057);
nand U14206 (N_14206,N_13100,N_13916);
xnor U14207 (N_14207,N_13442,N_13794);
and U14208 (N_14208,N_13700,N_13056);
nor U14209 (N_14209,N_13372,N_13858);
nand U14210 (N_14210,N_13613,N_13973);
nand U14211 (N_14211,N_13680,N_13825);
nand U14212 (N_14212,N_13912,N_13748);
nor U14213 (N_14213,N_13011,N_13002);
and U14214 (N_14214,N_13576,N_13844);
and U14215 (N_14215,N_13476,N_13230);
nor U14216 (N_14216,N_13742,N_13754);
nor U14217 (N_14217,N_13008,N_13855);
or U14218 (N_14218,N_13896,N_13467);
nor U14219 (N_14219,N_13910,N_13953);
or U14220 (N_14220,N_13141,N_13422);
and U14221 (N_14221,N_13847,N_13162);
nor U14222 (N_14222,N_13592,N_13944);
nand U14223 (N_14223,N_13697,N_13483);
nand U14224 (N_14224,N_13410,N_13692);
nor U14225 (N_14225,N_13723,N_13918);
or U14226 (N_14226,N_13115,N_13895);
and U14227 (N_14227,N_13549,N_13841);
nand U14228 (N_14228,N_13940,N_13437);
nand U14229 (N_14229,N_13977,N_13883);
nor U14230 (N_14230,N_13635,N_13392);
xor U14231 (N_14231,N_13997,N_13517);
nor U14232 (N_14232,N_13068,N_13935);
or U14233 (N_14233,N_13622,N_13803);
nor U14234 (N_14234,N_13620,N_13443);
xnor U14235 (N_14235,N_13589,N_13118);
xor U14236 (N_14236,N_13808,N_13166);
xnor U14237 (N_14237,N_13898,N_13740);
nand U14238 (N_14238,N_13288,N_13289);
xnor U14239 (N_14239,N_13035,N_13334);
or U14240 (N_14240,N_13851,N_13933);
nor U14241 (N_14241,N_13807,N_13768);
or U14242 (N_14242,N_13943,N_13219);
and U14243 (N_14243,N_13108,N_13785);
xnor U14244 (N_14244,N_13231,N_13254);
nand U14245 (N_14245,N_13673,N_13208);
and U14246 (N_14246,N_13972,N_13184);
nand U14247 (N_14247,N_13668,N_13222);
nand U14248 (N_14248,N_13485,N_13249);
and U14249 (N_14249,N_13259,N_13298);
nor U14250 (N_14250,N_13234,N_13261);
or U14251 (N_14251,N_13131,N_13262);
xor U14252 (N_14252,N_13064,N_13875);
and U14253 (N_14253,N_13479,N_13971);
xor U14254 (N_14254,N_13806,N_13837);
nand U14255 (N_14255,N_13096,N_13701);
nand U14256 (N_14256,N_13421,N_13253);
xnor U14257 (N_14257,N_13110,N_13607);
xor U14258 (N_14258,N_13650,N_13324);
xnor U14259 (N_14259,N_13344,N_13509);
nor U14260 (N_14260,N_13767,N_13001);
or U14261 (N_14261,N_13146,N_13335);
nor U14262 (N_14262,N_13715,N_13143);
nor U14263 (N_14263,N_13029,N_13067);
xor U14264 (N_14264,N_13597,N_13891);
or U14265 (N_14265,N_13870,N_13272);
and U14266 (N_14266,N_13059,N_13436);
or U14267 (N_14267,N_13155,N_13952);
and U14268 (N_14268,N_13128,N_13787);
xor U14269 (N_14269,N_13028,N_13515);
and U14270 (N_14270,N_13284,N_13525);
and U14271 (N_14271,N_13593,N_13904);
or U14272 (N_14272,N_13951,N_13400);
or U14273 (N_14273,N_13670,N_13527);
nand U14274 (N_14274,N_13664,N_13920);
and U14275 (N_14275,N_13712,N_13629);
xor U14276 (N_14276,N_13616,N_13731);
nand U14277 (N_14277,N_13373,N_13390);
nor U14278 (N_14278,N_13151,N_13639);
and U14279 (N_14279,N_13117,N_13164);
nor U14280 (N_14280,N_13843,N_13322);
and U14281 (N_14281,N_13426,N_13265);
or U14282 (N_14282,N_13498,N_13447);
xor U14283 (N_14283,N_13702,N_13165);
or U14284 (N_14284,N_13060,N_13983);
nand U14285 (N_14285,N_13503,N_13332);
xnor U14286 (N_14286,N_13772,N_13969);
xor U14287 (N_14287,N_13590,N_13223);
or U14288 (N_14288,N_13508,N_13955);
nand U14289 (N_14289,N_13121,N_13663);
or U14290 (N_14290,N_13310,N_13735);
or U14291 (N_14291,N_13625,N_13149);
nor U14292 (N_14292,N_13086,N_13098);
and U14293 (N_14293,N_13660,N_13737);
nand U14294 (N_14294,N_13733,N_13397);
nor U14295 (N_14295,N_13374,N_13042);
xnor U14296 (N_14296,N_13729,N_13813);
or U14297 (N_14297,N_13052,N_13678);
nand U14298 (N_14298,N_13565,N_13793);
nand U14299 (N_14299,N_13181,N_13050);
or U14300 (N_14300,N_13637,N_13153);
nand U14301 (N_14301,N_13348,N_13611);
or U14302 (N_14302,N_13290,N_13545);
or U14303 (N_14303,N_13120,N_13452);
nand U14304 (N_14304,N_13950,N_13089);
xor U14305 (N_14305,N_13757,N_13534);
or U14306 (N_14306,N_13345,N_13186);
nor U14307 (N_14307,N_13269,N_13975);
nand U14308 (N_14308,N_13460,N_13480);
and U14309 (N_14309,N_13791,N_13559);
and U14310 (N_14310,N_13404,N_13965);
and U14311 (N_14311,N_13496,N_13182);
or U14312 (N_14312,N_13619,N_13884);
and U14313 (N_14313,N_13796,N_13762);
nand U14314 (N_14314,N_13938,N_13268);
and U14315 (N_14315,N_13313,N_13763);
or U14316 (N_14316,N_13466,N_13474);
nand U14317 (N_14317,N_13456,N_13615);
nor U14318 (N_14318,N_13170,N_13279);
nand U14319 (N_14319,N_13316,N_13396);
xnor U14320 (N_14320,N_13959,N_13658);
xnor U14321 (N_14321,N_13431,N_13251);
nand U14322 (N_14322,N_13472,N_13174);
or U14323 (N_14323,N_13603,N_13649);
xor U14324 (N_14324,N_13927,N_13554);
or U14325 (N_14325,N_13630,N_13350);
nand U14326 (N_14326,N_13492,N_13075);
or U14327 (N_14327,N_13465,N_13698);
nor U14328 (N_14328,N_13828,N_13849);
xor U14329 (N_14329,N_13505,N_13994);
and U14330 (N_14330,N_13252,N_13039);
nand U14331 (N_14331,N_13872,N_13183);
nor U14332 (N_14332,N_13575,N_13522);
xnor U14333 (N_14333,N_13278,N_13688);
and U14334 (N_14334,N_13693,N_13643);
nand U14335 (N_14335,N_13963,N_13087);
nand U14336 (N_14336,N_13200,N_13546);
or U14337 (N_14337,N_13691,N_13797);
nor U14338 (N_14338,N_13718,N_13846);
nand U14339 (N_14339,N_13203,N_13106);
or U14340 (N_14340,N_13542,N_13677);
nand U14341 (N_14341,N_13292,N_13427);
nor U14342 (N_14342,N_13364,N_13016);
or U14343 (N_14343,N_13572,N_13260);
and U14344 (N_14344,N_13280,N_13354);
nor U14345 (N_14345,N_13113,N_13513);
nand U14346 (N_14346,N_13342,N_13887);
or U14347 (N_14347,N_13653,N_13696);
or U14348 (N_14348,N_13214,N_13970);
xnor U14349 (N_14349,N_13395,N_13486);
nand U14350 (N_14350,N_13005,N_13623);
or U14351 (N_14351,N_13077,N_13661);
xnor U14352 (N_14352,N_13293,N_13168);
nor U14353 (N_14353,N_13226,N_13413);
nand U14354 (N_14354,N_13013,N_13928);
or U14355 (N_14355,N_13666,N_13585);
xnor U14356 (N_14356,N_13842,N_13066);
or U14357 (N_14357,N_13306,N_13958);
xor U14358 (N_14358,N_13512,N_13897);
xnor U14359 (N_14359,N_13482,N_13360);
or U14360 (N_14360,N_13454,N_13911);
xnor U14361 (N_14361,N_13025,N_13695);
and U14362 (N_14362,N_13648,N_13338);
and U14363 (N_14363,N_13062,N_13987);
xnor U14364 (N_14364,N_13521,N_13220);
nor U14365 (N_14365,N_13632,N_13433);
nor U14366 (N_14366,N_13111,N_13020);
nor U14367 (N_14367,N_13934,N_13514);
nor U14368 (N_14368,N_13286,N_13758);
nor U14369 (N_14369,N_13818,N_13869);
and U14370 (N_14370,N_13532,N_13871);
and U14371 (N_14371,N_13083,N_13484);
nand U14372 (N_14372,N_13368,N_13273);
xnor U14373 (N_14373,N_13656,N_13138);
or U14374 (N_14374,N_13610,N_13048);
nor U14375 (N_14375,N_13415,N_13612);
xor U14376 (N_14376,N_13488,N_13207);
nor U14377 (N_14377,N_13387,N_13741);
nor U14378 (N_14378,N_13866,N_13609);
nand U14379 (N_14379,N_13319,N_13209);
or U14380 (N_14380,N_13591,N_13511);
xnor U14381 (N_14381,N_13817,N_13531);
xor U14382 (N_14382,N_13330,N_13995);
nand U14383 (N_14383,N_13009,N_13776);
and U14384 (N_14384,N_13633,N_13435);
xor U14385 (N_14385,N_13811,N_13881);
or U14386 (N_14386,N_13889,N_13136);
and U14387 (N_14387,N_13759,N_13156);
or U14388 (N_14388,N_13351,N_13257);
nor U14389 (N_14389,N_13703,N_13388);
nand U14390 (N_14390,N_13270,N_13765);
nand U14391 (N_14391,N_13880,N_13105);
nand U14392 (N_14392,N_13407,N_13044);
or U14393 (N_14393,N_13125,N_13903);
nor U14394 (N_14394,N_13346,N_13010);
nand U14395 (N_14395,N_13830,N_13383);
or U14396 (N_14396,N_13749,N_13939);
nand U14397 (N_14397,N_13710,N_13901);
nand U14398 (N_14398,N_13124,N_13499);
nor U14399 (N_14399,N_13675,N_13453);
nor U14400 (N_14400,N_13504,N_13441);
nor U14401 (N_14401,N_13475,N_13302);
xnor U14402 (N_14402,N_13905,N_13961);
and U14403 (N_14403,N_13922,N_13923);
xor U14404 (N_14404,N_13584,N_13063);
xnor U14405 (N_14405,N_13992,N_13523);
nor U14406 (N_14406,N_13127,N_13242);
nor U14407 (N_14407,N_13246,N_13683);
nand U14408 (N_14408,N_13689,N_13917);
xnor U14409 (N_14409,N_13672,N_13888);
or U14410 (N_14410,N_13533,N_13216);
or U14411 (N_14411,N_13107,N_13095);
nor U14412 (N_14412,N_13964,N_13180);
and U14413 (N_14413,N_13536,N_13369);
xnor U14414 (N_14414,N_13804,N_13225);
xor U14415 (N_14415,N_13295,N_13084);
xnor U14416 (N_14416,N_13694,N_13004);
nand U14417 (N_14417,N_13455,N_13206);
and U14418 (N_14418,N_13908,N_13420);
xor U14419 (N_14419,N_13362,N_13189);
xnor U14420 (N_14420,N_13877,N_13570);
nand U14421 (N_14421,N_13926,N_13582);
nand U14422 (N_14422,N_13947,N_13080);
or U14423 (N_14423,N_13046,N_13382);
nand U14424 (N_14424,N_13730,N_13529);
nor U14425 (N_14425,N_13477,N_13548);
and U14426 (N_14426,N_13243,N_13760);
xnor U14427 (N_14427,N_13706,N_13367);
xor U14428 (N_14428,N_13494,N_13876);
and U14429 (N_14429,N_13489,N_13539);
nor U14430 (N_14430,N_13921,N_13148);
and U14431 (N_14431,N_13782,N_13705);
xor U14432 (N_14432,N_13205,N_13769);
xor U14433 (N_14433,N_13053,N_13340);
xor U14434 (N_14434,N_13500,N_13805);
nor U14435 (N_14435,N_13874,N_13079);
nor U14436 (N_14436,N_13157,N_13856);
and U14437 (N_14437,N_13378,N_13419);
xnor U14438 (N_14438,N_13430,N_13134);
and U14439 (N_14439,N_13976,N_13034);
and U14440 (N_14440,N_13238,N_13621);
nand U14441 (N_14441,N_13006,N_13412);
nand U14442 (N_14442,N_13308,N_13497);
nand U14443 (N_14443,N_13221,N_13669);
and U14444 (N_14444,N_13932,N_13868);
nand U14445 (N_14445,N_13617,N_13626);
nor U14446 (N_14446,N_13176,N_13595);
nand U14447 (N_14447,N_13076,N_13296);
nor U14448 (N_14448,N_13979,N_13468);
nor U14449 (N_14449,N_13091,N_13457);
xor U14450 (N_14450,N_13103,N_13326);
and U14451 (N_14451,N_13294,N_13394);
nor U14452 (N_14452,N_13978,N_13366);
and U14453 (N_14453,N_13798,N_13739);
and U14454 (N_14454,N_13999,N_13341);
xor U14455 (N_14455,N_13832,N_13281);
xnor U14456 (N_14456,N_13890,N_13065);
nand U14457 (N_14457,N_13879,N_13745);
and U14458 (N_14458,N_13450,N_13516);
and U14459 (N_14459,N_13291,N_13645);
or U14460 (N_14460,N_13577,N_13036);
and U14461 (N_14461,N_13439,N_13606);
nor U14462 (N_14462,N_13655,N_13713);
nand U14463 (N_14463,N_13861,N_13956);
or U14464 (N_14464,N_13833,N_13789);
xor U14465 (N_14465,N_13213,N_13839);
or U14466 (N_14466,N_13708,N_13824);
xnor U14467 (N_14467,N_13775,N_13732);
xnor U14468 (N_14468,N_13446,N_13704);
and U14469 (N_14469,N_13470,N_13049);
nand U14470 (N_14470,N_13878,N_13391);
and U14471 (N_14471,N_13093,N_13627);
nor U14472 (N_14472,N_13135,N_13402);
nor U14473 (N_14473,N_13676,N_13276);
and U14474 (N_14474,N_13809,N_13227);
nand U14475 (N_14475,N_13907,N_13628);
xnor U14476 (N_14476,N_13571,N_13906);
or U14477 (N_14477,N_13726,N_13761);
and U14478 (N_14478,N_13491,N_13985);
nor U14479 (N_14479,N_13026,N_13037);
xor U14480 (N_14480,N_13069,N_13801);
and U14481 (N_14481,N_13352,N_13321);
xor U14482 (N_14482,N_13196,N_13012);
nand U14483 (N_14483,N_13957,N_13553);
xor U14484 (N_14484,N_13746,N_13537);
nor U14485 (N_14485,N_13027,N_13501);
or U14486 (N_14486,N_13993,N_13287);
nand U14487 (N_14487,N_13684,N_13755);
nand U14488 (N_14488,N_13736,N_13423);
or U14489 (N_14489,N_13568,N_13380);
or U14490 (N_14490,N_13144,N_13602);
xnor U14491 (N_14491,N_13535,N_13081);
xnor U14492 (N_14492,N_13129,N_13478);
or U14493 (N_14493,N_13445,N_13199);
xor U14494 (N_14494,N_13974,N_13836);
nor U14495 (N_14495,N_13178,N_13188);
or U14496 (N_14496,N_13406,N_13047);
nand U14497 (N_14497,N_13783,N_13569);
xor U14498 (N_14498,N_13347,N_13894);
or U14499 (N_14499,N_13865,N_13187);
and U14500 (N_14500,N_13669,N_13536);
xnor U14501 (N_14501,N_13121,N_13972);
or U14502 (N_14502,N_13482,N_13309);
nand U14503 (N_14503,N_13205,N_13179);
and U14504 (N_14504,N_13063,N_13695);
or U14505 (N_14505,N_13026,N_13646);
and U14506 (N_14506,N_13376,N_13464);
nand U14507 (N_14507,N_13781,N_13969);
nand U14508 (N_14508,N_13636,N_13777);
and U14509 (N_14509,N_13832,N_13075);
and U14510 (N_14510,N_13048,N_13372);
or U14511 (N_14511,N_13342,N_13170);
or U14512 (N_14512,N_13876,N_13485);
xnor U14513 (N_14513,N_13913,N_13017);
nor U14514 (N_14514,N_13555,N_13297);
and U14515 (N_14515,N_13921,N_13737);
or U14516 (N_14516,N_13076,N_13380);
or U14517 (N_14517,N_13126,N_13819);
xnor U14518 (N_14518,N_13062,N_13767);
nor U14519 (N_14519,N_13430,N_13488);
and U14520 (N_14520,N_13884,N_13516);
and U14521 (N_14521,N_13113,N_13011);
or U14522 (N_14522,N_13664,N_13588);
or U14523 (N_14523,N_13454,N_13414);
xor U14524 (N_14524,N_13671,N_13354);
or U14525 (N_14525,N_13936,N_13856);
and U14526 (N_14526,N_13369,N_13016);
or U14527 (N_14527,N_13359,N_13387);
or U14528 (N_14528,N_13316,N_13052);
xnor U14529 (N_14529,N_13728,N_13465);
nor U14530 (N_14530,N_13196,N_13299);
or U14531 (N_14531,N_13972,N_13660);
nor U14532 (N_14532,N_13017,N_13113);
and U14533 (N_14533,N_13739,N_13378);
or U14534 (N_14534,N_13578,N_13100);
nor U14535 (N_14535,N_13768,N_13210);
nand U14536 (N_14536,N_13713,N_13009);
or U14537 (N_14537,N_13325,N_13426);
nor U14538 (N_14538,N_13928,N_13079);
xnor U14539 (N_14539,N_13354,N_13999);
nor U14540 (N_14540,N_13900,N_13155);
xnor U14541 (N_14541,N_13902,N_13114);
xnor U14542 (N_14542,N_13812,N_13892);
xor U14543 (N_14543,N_13315,N_13116);
or U14544 (N_14544,N_13688,N_13148);
or U14545 (N_14545,N_13140,N_13700);
and U14546 (N_14546,N_13235,N_13147);
nor U14547 (N_14547,N_13453,N_13025);
nor U14548 (N_14548,N_13161,N_13510);
or U14549 (N_14549,N_13590,N_13738);
nand U14550 (N_14550,N_13461,N_13097);
and U14551 (N_14551,N_13999,N_13560);
nand U14552 (N_14552,N_13874,N_13338);
or U14553 (N_14553,N_13180,N_13230);
nand U14554 (N_14554,N_13267,N_13208);
or U14555 (N_14555,N_13417,N_13215);
nor U14556 (N_14556,N_13470,N_13356);
nand U14557 (N_14557,N_13493,N_13004);
and U14558 (N_14558,N_13126,N_13452);
nand U14559 (N_14559,N_13413,N_13219);
nor U14560 (N_14560,N_13423,N_13639);
and U14561 (N_14561,N_13406,N_13627);
xor U14562 (N_14562,N_13207,N_13192);
and U14563 (N_14563,N_13511,N_13876);
xor U14564 (N_14564,N_13437,N_13655);
and U14565 (N_14565,N_13261,N_13706);
xnor U14566 (N_14566,N_13436,N_13806);
xor U14567 (N_14567,N_13369,N_13123);
xor U14568 (N_14568,N_13005,N_13211);
and U14569 (N_14569,N_13055,N_13498);
and U14570 (N_14570,N_13480,N_13075);
nand U14571 (N_14571,N_13817,N_13616);
nand U14572 (N_14572,N_13387,N_13928);
nand U14573 (N_14573,N_13035,N_13141);
xnor U14574 (N_14574,N_13841,N_13421);
nor U14575 (N_14575,N_13330,N_13367);
nor U14576 (N_14576,N_13050,N_13083);
nand U14577 (N_14577,N_13333,N_13182);
and U14578 (N_14578,N_13832,N_13275);
nor U14579 (N_14579,N_13972,N_13938);
or U14580 (N_14580,N_13137,N_13977);
xnor U14581 (N_14581,N_13740,N_13656);
xor U14582 (N_14582,N_13640,N_13996);
nand U14583 (N_14583,N_13180,N_13136);
or U14584 (N_14584,N_13165,N_13303);
or U14585 (N_14585,N_13613,N_13740);
and U14586 (N_14586,N_13216,N_13182);
or U14587 (N_14587,N_13369,N_13210);
xnor U14588 (N_14588,N_13176,N_13334);
xnor U14589 (N_14589,N_13288,N_13415);
and U14590 (N_14590,N_13874,N_13862);
or U14591 (N_14591,N_13433,N_13614);
and U14592 (N_14592,N_13609,N_13400);
xor U14593 (N_14593,N_13696,N_13812);
nor U14594 (N_14594,N_13852,N_13347);
nor U14595 (N_14595,N_13311,N_13291);
nand U14596 (N_14596,N_13832,N_13679);
nand U14597 (N_14597,N_13279,N_13442);
or U14598 (N_14598,N_13088,N_13312);
or U14599 (N_14599,N_13335,N_13745);
or U14600 (N_14600,N_13811,N_13831);
or U14601 (N_14601,N_13433,N_13309);
or U14602 (N_14602,N_13550,N_13459);
nand U14603 (N_14603,N_13389,N_13667);
or U14604 (N_14604,N_13913,N_13299);
nor U14605 (N_14605,N_13761,N_13003);
or U14606 (N_14606,N_13328,N_13608);
nor U14607 (N_14607,N_13210,N_13593);
nor U14608 (N_14608,N_13729,N_13606);
nand U14609 (N_14609,N_13551,N_13807);
xor U14610 (N_14610,N_13254,N_13554);
and U14611 (N_14611,N_13947,N_13135);
xor U14612 (N_14612,N_13943,N_13193);
nor U14613 (N_14613,N_13637,N_13464);
or U14614 (N_14614,N_13051,N_13527);
xnor U14615 (N_14615,N_13290,N_13883);
and U14616 (N_14616,N_13441,N_13304);
nor U14617 (N_14617,N_13730,N_13233);
and U14618 (N_14618,N_13646,N_13469);
nand U14619 (N_14619,N_13727,N_13728);
xor U14620 (N_14620,N_13692,N_13171);
xnor U14621 (N_14621,N_13018,N_13502);
and U14622 (N_14622,N_13872,N_13210);
xor U14623 (N_14623,N_13304,N_13230);
xnor U14624 (N_14624,N_13997,N_13139);
nand U14625 (N_14625,N_13513,N_13951);
nor U14626 (N_14626,N_13853,N_13091);
and U14627 (N_14627,N_13665,N_13557);
or U14628 (N_14628,N_13253,N_13399);
and U14629 (N_14629,N_13580,N_13772);
and U14630 (N_14630,N_13066,N_13816);
xor U14631 (N_14631,N_13580,N_13143);
nor U14632 (N_14632,N_13276,N_13236);
nor U14633 (N_14633,N_13416,N_13221);
nor U14634 (N_14634,N_13127,N_13694);
and U14635 (N_14635,N_13632,N_13044);
and U14636 (N_14636,N_13839,N_13082);
nand U14637 (N_14637,N_13559,N_13646);
xor U14638 (N_14638,N_13723,N_13397);
xor U14639 (N_14639,N_13619,N_13076);
and U14640 (N_14640,N_13698,N_13370);
or U14641 (N_14641,N_13395,N_13666);
nor U14642 (N_14642,N_13229,N_13034);
nand U14643 (N_14643,N_13816,N_13525);
nand U14644 (N_14644,N_13455,N_13550);
and U14645 (N_14645,N_13242,N_13440);
nor U14646 (N_14646,N_13211,N_13417);
nand U14647 (N_14647,N_13579,N_13824);
xor U14648 (N_14648,N_13061,N_13826);
or U14649 (N_14649,N_13273,N_13930);
or U14650 (N_14650,N_13465,N_13264);
nor U14651 (N_14651,N_13605,N_13475);
xor U14652 (N_14652,N_13888,N_13679);
or U14653 (N_14653,N_13468,N_13497);
and U14654 (N_14654,N_13498,N_13207);
nand U14655 (N_14655,N_13586,N_13209);
and U14656 (N_14656,N_13251,N_13338);
xnor U14657 (N_14657,N_13435,N_13743);
nor U14658 (N_14658,N_13887,N_13794);
and U14659 (N_14659,N_13435,N_13774);
nor U14660 (N_14660,N_13592,N_13011);
and U14661 (N_14661,N_13125,N_13582);
nand U14662 (N_14662,N_13563,N_13323);
or U14663 (N_14663,N_13613,N_13419);
nand U14664 (N_14664,N_13907,N_13305);
or U14665 (N_14665,N_13798,N_13499);
or U14666 (N_14666,N_13069,N_13873);
and U14667 (N_14667,N_13997,N_13969);
xnor U14668 (N_14668,N_13371,N_13692);
nor U14669 (N_14669,N_13221,N_13066);
nor U14670 (N_14670,N_13341,N_13617);
and U14671 (N_14671,N_13477,N_13211);
or U14672 (N_14672,N_13239,N_13522);
xor U14673 (N_14673,N_13856,N_13994);
nor U14674 (N_14674,N_13004,N_13458);
or U14675 (N_14675,N_13057,N_13466);
or U14676 (N_14676,N_13861,N_13081);
or U14677 (N_14677,N_13004,N_13253);
or U14678 (N_14678,N_13593,N_13379);
or U14679 (N_14679,N_13769,N_13931);
and U14680 (N_14680,N_13247,N_13435);
and U14681 (N_14681,N_13070,N_13296);
nor U14682 (N_14682,N_13830,N_13459);
and U14683 (N_14683,N_13491,N_13212);
nor U14684 (N_14684,N_13072,N_13357);
nand U14685 (N_14685,N_13642,N_13373);
nor U14686 (N_14686,N_13240,N_13663);
or U14687 (N_14687,N_13552,N_13399);
or U14688 (N_14688,N_13023,N_13498);
and U14689 (N_14689,N_13685,N_13367);
nor U14690 (N_14690,N_13791,N_13669);
or U14691 (N_14691,N_13718,N_13711);
xnor U14692 (N_14692,N_13216,N_13715);
xnor U14693 (N_14693,N_13642,N_13707);
nand U14694 (N_14694,N_13936,N_13360);
nor U14695 (N_14695,N_13513,N_13703);
and U14696 (N_14696,N_13320,N_13829);
or U14697 (N_14697,N_13708,N_13209);
nand U14698 (N_14698,N_13608,N_13992);
nand U14699 (N_14699,N_13866,N_13970);
and U14700 (N_14700,N_13744,N_13451);
and U14701 (N_14701,N_13546,N_13872);
xnor U14702 (N_14702,N_13425,N_13918);
or U14703 (N_14703,N_13179,N_13174);
nor U14704 (N_14704,N_13239,N_13291);
xor U14705 (N_14705,N_13634,N_13209);
nand U14706 (N_14706,N_13104,N_13345);
or U14707 (N_14707,N_13308,N_13916);
or U14708 (N_14708,N_13762,N_13160);
nor U14709 (N_14709,N_13373,N_13213);
nand U14710 (N_14710,N_13395,N_13040);
or U14711 (N_14711,N_13758,N_13486);
nor U14712 (N_14712,N_13087,N_13332);
nor U14713 (N_14713,N_13718,N_13698);
or U14714 (N_14714,N_13374,N_13495);
xnor U14715 (N_14715,N_13772,N_13785);
nor U14716 (N_14716,N_13485,N_13710);
and U14717 (N_14717,N_13325,N_13298);
and U14718 (N_14718,N_13728,N_13783);
nor U14719 (N_14719,N_13669,N_13689);
nor U14720 (N_14720,N_13987,N_13216);
nor U14721 (N_14721,N_13079,N_13432);
or U14722 (N_14722,N_13152,N_13826);
or U14723 (N_14723,N_13522,N_13115);
and U14724 (N_14724,N_13556,N_13282);
xor U14725 (N_14725,N_13329,N_13343);
or U14726 (N_14726,N_13880,N_13688);
and U14727 (N_14727,N_13986,N_13971);
xor U14728 (N_14728,N_13810,N_13756);
nor U14729 (N_14729,N_13586,N_13575);
and U14730 (N_14730,N_13382,N_13783);
nand U14731 (N_14731,N_13237,N_13376);
and U14732 (N_14732,N_13423,N_13720);
xor U14733 (N_14733,N_13941,N_13921);
xor U14734 (N_14734,N_13043,N_13465);
or U14735 (N_14735,N_13435,N_13333);
nand U14736 (N_14736,N_13093,N_13920);
or U14737 (N_14737,N_13421,N_13859);
or U14738 (N_14738,N_13719,N_13902);
nor U14739 (N_14739,N_13973,N_13887);
nand U14740 (N_14740,N_13364,N_13257);
or U14741 (N_14741,N_13217,N_13914);
nor U14742 (N_14742,N_13687,N_13723);
xnor U14743 (N_14743,N_13135,N_13734);
and U14744 (N_14744,N_13261,N_13647);
or U14745 (N_14745,N_13731,N_13160);
or U14746 (N_14746,N_13172,N_13173);
xor U14747 (N_14747,N_13327,N_13266);
xor U14748 (N_14748,N_13694,N_13367);
and U14749 (N_14749,N_13882,N_13944);
xor U14750 (N_14750,N_13973,N_13180);
or U14751 (N_14751,N_13380,N_13394);
nand U14752 (N_14752,N_13043,N_13991);
nor U14753 (N_14753,N_13113,N_13942);
xnor U14754 (N_14754,N_13338,N_13893);
xor U14755 (N_14755,N_13603,N_13568);
xor U14756 (N_14756,N_13231,N_13521);
and U14757 (N_14757,N_13423,N_13818);
and U14758 (N_14758,N_13313,N_13127);
or U14759 (N_14759,N_13154,N_13149);
xor U14760 (N_14760,N_13372,N_13289);
xor U14761 (N_14761,N_13799,N_13232);
nor U14762 (N_14762,N_13724,N_13935);
and U14763 (N_14763,N_13698,N_13574);
and U14764 (N_14764,N_13691,N_13776);
nand U14765 (N_14765,N_13200,N_13494);
nor U14766 (N_14766,N_13385,N_13440);
and U14767 (N_14767,N_13135,N_13796);
nand U14768 (N_14768,N_13561,N_13832);
or U14769 (N_14769,N_13967,N_13146);
and U14770 (N_14770,N_13884,N_13471);
or U14771 (N_14771,N_13262,N_13209);
xor U14772 (N_14772,N_13301,N_13654);
or U14773 (N_14773,N_13180,N_13132);
xor U14774 (N_14774,N_13079,N_13970);
or U14775 (N_14775,N_13524,N_13044);
or U14776 (N_14776,N_13157,N_13562);
nand U14777 (N_14777,N_13744,N_13015);
nand U14778 (N_14778,N_13209,N_13231);
or U14779 (N_14779,N_13265,N_13852);
and U14780 (N_14780,N_13763,N_13649);
or U14781 (N_14781,N_13553,N_13475);
or U14782 (N_14782,N_13717,N_13484);
nand U14783 (N_14783,N_13051,N_13968);
nand U14784 (N_14784,N_13218,N_13960);
nor U14785 (N_14785,N_13338,N_13339);
nand U14786 (N_14786,N_13847,N_13350);
nand U14787 (N_14787,N_13896,N_13965);
nor U14788 (N_14788,N_13687,N_13470);
nand U14789 (N_14789,N_13502,N_13553);
or U14790 (N_14790,N_13132,N_13593);
xor U14791 (N_14791,N_13665,N_13649);
xnor U14792 (N_14792,N_13168,N_13472);
xor U14793 (N_14793,N_13730,N_13637);
nor U14794 (N_14794,N_13754,N_13239);
and U14795 (N_14795,N_13860,N_13029);
xor U14796 (N_14796,N_13365,N_13224);
and U14797 (N_14797,N_13258,N_13093);
nand U14798 (N_14798,N_13096,N_13982);
nor U14799 (N_14799,N_13312,N_13407);
and U14800 (N_14800,N_13501,N_13473);
nand U14801 (N_14801,N_13648,N_13515);
and U14802 (N_14802,N_13545,N_13047);
and U14803 (N_14803,N_13251,N_13976);
nand U14804 (N_14804,N_13142,N_13633);
nor U14805 (N_14805,N_13972,N_13865);
or U14806 (N_14806,N_13604,N_13221);
and U14807 (N_14807,N_13225,N_13243);
nor U14808 (N_14808,N_13596,N_13302);
and U14809 (N_14809,N_13970,N_13891);
xor U14810 (N_14810,N_13359,N_13508);
xnor U14811 (N_14811,N_13818,N_13520);
xnor U14812 (N_14812,N_13057,N_13376);
xnor U14813 (N_14813,N_13020,N_13755);
and U14814 (N_14814,N_13803,N_13544);
nand U14815 (N_14815,N_13284,N_13620);
xnor U14816 (N_14816,N_13723,N_13439);
xor U14817 (N_14817,N_13592,N_13660);
or U14818 (N_14818,N_13176,N_13239);
nor U14819 (N_14819,N_13253,N_13843);
nand U14820 (N_14820,N_13063,N_13725);
nand U14821 (N_14821,N_13332,N_13640);
or U14822 (N_14822,N_13368,N_13776);
nor U14823 (N_14823,N_13366,N_13630);
nand U14824 (N_14824,N_13183,N_13826);
nor U14825 (N_14825,N_13758,N_13470);
xor U14826 (N_14826,N_13415,N_13233);
nor U14827 (N_14827,N_13942,N_13743);
or U14828 (N_14828,N_13227,N_13456);
xor U14829 (N_14829,N_13338,N_13359);
and U14830 (N_14830,N_13540,N_13213);
or U14831 (N_14831,N_13062,N_13905);
nand U14832 (N_14832,N_13433,N_13034);
nand U14833 (N_14833,N_13778,N_13342);
nand U14834 (N_14834,N_13215,N_13413);
xnor U14835 (N_14835,N_13581,N_13742);
xor U14836 (N_14836,N_13669,N_13625);
xor U14837 (N_14837,N_13793,N_13231);
nor U14838 (N_14838,N_13640,N_13620);
xor U14839 (N_14839,N_13303,N_13428);
or U14840 (N_14840,N_13671,N_13005);
nand U14841 (N_14841,N_13769,N_13944);
and U14842 (N_14842,N_13598,N_13757);
nor U14843 (N_14843,N_13043,N_13467);
xor U14844 (N_14844,N_13505,N_13682);
nand U14845 (N_14845,N_13128,N_13249);
nor U14846 (N_14846,N_13962,N_13952);
or U14847 (N_14847,N_13129,N_13945);
nor U14848 (N_14848,N_13601,N_13280);
nor U14849 (N_14849,N_13689,N_13036);
and U14850 (N_14850,N_13439,N_13253);
xor U14851 (N_14851,N_13902,N_13651);
and U14852 (N_14852,N_13445,N_13924);
or U14853 (N_14853,N_13706,N_13288);
nor U14854 (N_14854,N_13728,N_13127);
or U14855 (N_14855,N_13457,N_13815);
xor U14856 (N_14856,N_13493,N_13488);
or U14857 (N_14857,N_13681,N_13990);
nand U14858 (N_14858,N_13858,N_13920);
or U14859 (N_14859,N_13124,N_13445);
or U14860 (N_14860,N_13129,N_13461);
nor U14861 (N_14861,N_13171,N_13912);
or U14862 (N_14862,N_13693,N_13794);
nand U14863 (N_14863,N_13694,N_13671);
xor U14864 (N_14864,N_13858,N_13341);
or U14865 (N_14865,N_13259,N_13196);
nor U14866 (N_14866,N_13029,N_13269);
and U14867 (N_14867,N_13676,N_13151);
nand U14868 (N_14868,N_13750,N_13388);
nor U14869 (N_14869,N_13744,N_13811);
nor U14870 (N_14870,N_13332,N_13439);
nand U14871 (N_14871,N_13838,N_13650);
or U14872 (N_14872,N_13293,N_13409);
or U14873 (N_14873,N_13857,N_13115);
nand U14874 (N_14874,N_13316,N_13125);
or U14875 (N_14875,N_13696,N_13976);
nand U14876 (N_14876,N_13256,N_13412);
nor U14877 (N_14877,N_13107,N_13768);
nand U14878 (N_14878,N_13819,N_13037);
nand U14879 (N_14879,N_13957,N_13164);
and U14880 (N_14880,N_13728,N_13138);
nor U14881 (N_14881,N_13134,N_13464);
or U14882 (N_14882,N_13607,N_13609);
nor U14883 (N_14883,N_13935,N_13388);
nand U14884 (N_14884,N_13202,N_13611);
nor U14885 (N_14885,N_13588,N_13850);
or U14886 (N_14886,N_13757,N_13591);
nor U14887 (N_14887,N_13362,N_13392);
and U14888 (N_14888,N_13389,N_13558);
and U14889 (N_14889,N_13414,N_13741);
nand U14890 (N_14890,N_13909,N_13290);
nand U14891 (N_14891,N_13336,N_13268);
xor U14892 (N_14892,N_13028,N_13661);
xnor U14893 (N_14893,N_13716,N_13078);
xnor U14894 (N_14894,N_13805,N_13425);
nand U14895 (N_14895,N_13336,N_13486);
or U14896 (N_14896,N_13093,N_13217);
and U14897 (N_14897,N_13714,N_13879);
xor U14898 (N_14898,N_13574,N_13338);
or U14899 (N_14899,N_13593,N_13267);
nor U14900 (N_14900,N_13743,N_13053);
xnor U14901 (N_14901,N_13010,N_13935);
nand U14902 (N_14902,N_13009,N_13359);
xnor U14903 (N_14903,N_13513,N_13103);
xnor U14904 (N_14904,N_13500,N_13671);
nor U14905 (N_14905,N_13010,N_13005);
xor U14906 (N_14906,N_13175,N_13879);
or U14907 (N_14907,N_13264,N_13231);
or U14908 (N_14908,N_13995,N_13516);
or U14909 (N_14909,N_13147,N_13961);
nand U14910 (N_14910,N_13001,N_13251);
xnor U14911 (N_14911,N_13496,N_13387);
nand U14912 (N_14912,N_13741,N_13585);
nand U14913 (N_14913,N_13906,N_13468);
and U14914 (N_14914,N_13603,N_13685);
xor U14915 (N_14915,N_13943,N_13160);
nand U14916 (N_14916,N_13421,N_13014);
or U14917 (N_14917,N_13711,N_13766);
nand U14918 (N_14918,N_13094,N_13464);
nor U14919 (N_14919,N_13076,N_13815);
nor U14920 (N_14920,N_13751,N_13745);
or U14921 (N_14921,N_13766,N_13650);
xor U14922 (N_14922,N_13095,N_13377);
nor U14923 (N_14923,N_13145,N_13926);
nand U14924 (N_14924,N_13471,N_13629);
nor U14925 (N_14925,N_13059,N_13134);
xnor U14926 (N_14926,N_13789,N_13323);
or U14927 (N_14927,N_13347,N_13635);
and U14928 (N_14928,N_13679,N_13021);
nand U14929 (N_14929,N_13631,N_13518);
and U14930 (N_14930,N_13842,N_13018);
nand U14931 (N_14931,N_13418,N_13466);
xor U14932 (N_14932,N_13485,N_13259);
xnor U14933 (N_14933,N_13748,N_13492);
nor U14934 (N_14934,N_13420,N_13801);
or U14935 (N_14935,N_13152,N_13386);
nand U14936 (N_14936,N_13467,N_13215);
nor U14937 (N_14937,N_13663,N_13066);
nor U14938 (N_14938,N_13673,N_13228);
xor U14939 (N_14939,N_13333,N_13902);
and U14940 (N_14940,N_13057,N_13154);
or U14941 (N_14941,N_13557,N_13571);
and U14942 (N_14942,N_13021,N_13314);
or U14943 (N_14943,N_13543,N_13945);
and U14944 (N_14944,N_13473,N_13834);
and U14945 (N_14945,N_13541,N_13392);
nand U14946 (N_14946,N_13305,N_13044);
nor U14947 (N_14947,N_13631,N_13927);
xnor U14948 (N_14948,N_13942,N_13545);
nand U14949 (N_14949,N_13180,N_13769);
nor U14950 (N_14950,N_13689,N_13457);
and U14951 (N_14951,N_13929,N_13795);
or U14952 (N_14952,N_13390,N_13045);
nand U14953 (N_14953,N_13828,N_13752);
xnor U14954 (N_14954,N_13423,N_13831);
xor U14955 (N_14955,N_13432,N_13760);
or U14956 (N_14956,N_13984,N_13661);
or U14957 (N_14957,N_13460,N_13993);
xor U14958 (N_14958,N_13191,N_13647);
and U14959 (N_14959,N_13875,N_13494);
and U14960 (N_14960,N_13964,N_13225);
nor U14961 (N_14961,N_13694,N_13209);
nor U14962 (N_14962,N_13763,N_13073);
nand U14963 (N_14963,N_13231,N_13110);
and U14964 (N_14964,N_13311,N_13574);
nand U14965 (N_14965,N_13229,N_13282);
and U14966 (N_14966,N_13670,N_13329);
or U14967 (N_14967,N_13932,N_13857);
and U14968 (N_14968,N_13524,N_13335);
nor U14969 (N_14969,N_13023,N_13984);
and U14970 (N_14970,N_13330,N_13820);
and U14971 (N_14971,N_13389,N_13355);
and U14972 (N_14972,N_13056,N_13647);
and U14973 (N_14973,N_13003,N_13609);
and U14974 (N_14974,N_13402,N_13603);
xor U14975 (N_14975,N_13578,N_13654);
nor U14976 (N_14976,N_13304,N_13159);
nor U14977 (N_14977,N_13806,N_13376);
xor U14978 (N_14978,N_13619,N_13990);
nand U14979 (N_14979,N_13051,N_13922);
and U14980 (N_14980,N_13765,N_13536);
nor U14981 (N_14981,N_13895,N_13766);
and U14982 (N_14982,N_13519,N_13650);
nand U14983 (N_14983,N_13086,N_13909);
nor U14984 (N_14984,N_13923,N_13328);
and U14985 (N_14985,N_13649,N_13052);
nor U14986 (N_14986,N_13131,N_13859);
or U14987 (N_14987,N_13283,N_13132);
xor U14988 (N_14988,N_13319,N_13146);
and U14989 (N_14989,N_13969,N_13519);
nand U14990 (N_14990,N_13620,N_13924);
xor U14991 (N_14991,N_13140,N_13458);
xor U14992 (N_14992,N_13488,N_13104);
nand U14993 (N_14993,N_13282,N_13834);
and U14994 (N_14994,N_13094,N_13680);
and U14995 (N_14995,N_13528,N_13447);
nand U14996 (N_14996,N_13688,N_13081);
or U14997 (N_14997,N_13162,N_13529);
and U14998 (N_14998,N_13909,N_13230);
xor U14999 (N_14999,N_13655,N_13154);
and UO_0 (O_0,N_14828,N_14423);
nand UO_1 (O_1,N_14303,N_14752);
and UO_2 (O_2,N_14511,N_14967);
or UO_3 (O_3,N_14005,N_14591);
nor UO_4 (O_4,N_14589,N_14021);
and UO_5 (O_5,N_14566,N_14837);
nand UO_6 (O_6,N_14121,N_14137);
or UO_7 (O_7,N_14973,N_14314);
and UO_8 (O_8,N_14624,N_14559);
and UO_9 (O_9,N_14125,N_14133);
nor UO_10 (O_10,N_14236,N_14852);
nand UO_11 (O_11,N_14263,N_14335);
or UO_12 (O_12,N_14681,N_14092);
nand UO_13 (O_13,N_14848,N_14705);
nor UO_14 (O_14,N_14817,N_14963);
and UO_15 (O_15,N_14603,N_14155);
and UO_16 (O_16,N_14082,N_14222);
nor UO_17 (O_17,N_14711,N_14795);
or UO_18 (O_18,N_14994,N_14905);
and UO_19 (O_19,N_14651,N_14202);
nor UO_20 (O_20,N_14728,N_14023);
nor UO_21 (O_21,N_14912,N_14615);
nand UO_22 (O_22,N_14299,N_14324);
nand UO_23 (O_23,N_14838,N_14929);
nand UO_24 (O_24,N_14351,N_14506);
nand UO_25 (O_25,N_14399,N_14840);
and UO_26 (O_26,N_14085,N_14977);
xnor UO_27 (O_27,N_14238,N_14773);
xnor UO_28 (O_28,N_14461,N_14881);
nor UO_29 (O_29,N_14820,N_14574);
nand UO_30 (O_30,N_14485,N_14856);
or UO_31 (O_31,N_14671,N_14394);
xor UO_32 (O_32,N_14001,N_14302);
or UO_33 (O_33,N_14464,N_14971);
nand UO_34 (O_34,N_14906,N_14153);
or UO_35 (O_35,N_14459,N_14784);
and UO_36 (O_36,N_14446,N_14040);
xor UO_37 (O_37,N_14886,N_14327);
or UO_38 (O_38,N_14611,N_14357);
and UO_39 (O_39,N_14514,N_14478);
xor UO_40 (O_40,N_14969,N_14330);
and UO_41 (O_41,N_14715,N_14990);
xnor UO_42 (O_42,N_14173,N_14252);
and UO_43 (O_43,N_14738,N_14080);
xnor UO_44 (O_44,N_14420,N_14943);
or UO_45 (O_45,N_14777,N_14122);
or UO_46 (O_46,N_14344,N_14933);
nand UO_47 (O_47,N_14630,N_14916);
or UO_48 (O_48,N_14207,N_14689);
and UO_49 (O_49,N_14985,N_14783);
or UO_50 (O_50,N_14099,N_14223);
nand UO_51 (O_51,N_14073,N_14551);
and UO_52 (O_52,N_14751,N_14970);
and UO_53 (O_53,N_14575,N_14813);
and UO_54 (O_54,N_14918,N_14050);
or UO_55 (O_55,N_14988,N_14789);
xnor UO_56 (O_56,N_14634,N_14909);
nand UO_57 (O_57,N_14201,N_14758);
or UO_58 (O_58,N_14667,N_14588);
xnor UO_59 (O_59,N_14393,N_14444);
or UO_60 (O_60,N_14741,N_14458);
xor UO_61 (O_61,N_14234,N_14825);
xnor UO_62 (O_62,N_14814,N_14958);
or UO_63 (O_63,N_14554,N_14801);
nand UO_64 (O_64,N_14849,N_14417);
or UO_65 (O_65,N_14867,N_14205);
xnor UO_66 (O_66,N_14673,N_14522);
nand UO_67 (O_67,N_14161,N_14247);
or UO_68 (O_68,N_14437,N_14029);
nor UO_69 (O_69,N_14118,N_14046);
nor UO_70 (O_70,N_14489,N_14313);
or UO_71 (O_71,N_14187,N_14170);
nand UO_72 (O_72,N_14992,N_14112);
and UO_73 (O_73,N_14389,N_14614);
and UO_74 (O_74,N_14142,N_14077);
nand UO_75 (O_75,N_14024,N_14791);
or UO_76 (O_76,N_14650,N_14543);
xor UO_77 (O_77,N_14680,N_14128);
or UO_78 (O_78,N_14516,N_14719);
and UO_79 (O_79,N_14355,N_14225);
nor UO_80 (O_80,N_14013,N_14665);
xnor UO_81 (O_81,N_14494,N_14524);
or UO_82 (O_82,N_14669,N_14707);
nand UO_83 (O_83,N_14286,N_14796);
xnor UO_84 (O_84,N_14954,N_14877);
or UO_85 (O_85,N_14915,N_14310);
or UO_86 (O_86,N_14835,N_14701);
nand UO_87 (O_87,N_14925,N_14536);
and UO_88 (O_88,N_14894,N_14372);
or UO_89 (O_89,N_14298,N_14332);
xor UO_90 (O_90,N_14887,N_14800);
and UO_91 (O_91,N_14336,N_14815);
and UO_92 (O_92,N_14616,N_14192);
nor UO_93 (O_93,N_14189,N_14991);
or UO_94 (O_94,N_14025,N_14333);
or UO_95 (O_95,N_14226,N_14065);
or UO_96 (O_96,N_14316,N_14757);
or UO_97 (O_97,N_14291,N_14150);
xor UO_98 (O_98,N_14476,N_14974);
and UO_99 (O_99,N_14523,N_14340);
xor UO_100 (O_100,N_14410,N_14938);
xor UO_101 (O_101,N_14172,N_14471);
or UO_102 (O_102,N_14966,N_14870);
and UO_103 (O_103,N_14913,N_14384);
nor UO_104 (O_104,N_14910,N_14851);
nor UO_105 (O_105,N_14888,N_14358);
nor UO_106 (O_106,N_14095,N_14003);
xnor UO_107 (O_107,N_14660,N_14527);
nor UO_108 (O_108,N_14637,N_14167);
nor UO_109 (O_109,N_14467,N_14460);
xor UO_110 (O_110,N_14736,N_14058);
and UO_111 (O_111,N_14812,N_14889);
nor UO_112 (O_112,N_14253,N_14334);
nand UO_113 (O_113,N_14104,N_14296);
and UO_114 (O_114,N_14697,N_14433);
xnor UO_115 (O_115,N_14196,N_14127);
nor UO_116 (O_116,N_14064,N_14180);
and UO_117 (O_117,N_14203,N_14490);
and UO_118 (O_118,N_14972,N_14030);
nor UO_119 (O_119,N_14627,N_14592);
xor UO_120 (O_120,N_14034,N_14920);
nand UO_121 (O_121,N_14447,N_14059);
nand UO_122 (O_122,N_14568,N_14737);
and UO_123 (O_123,N_14135,N_14934);
or UO_124 (O_124,N_14367,N_14157);
and UO_125 (O_125,N_14275,N_14045);
nor UO_126 (O_126,N_14590,N_14011);
nor UO_127 (O_127,N_14750,N_14288);
nand UO_128 (O_128,N_14465,N_14239);
nor UO_129 (O_129,N_14079,N_14558);
or UO_130 (O_130,N_14139,N_14858);
nor UO_131 (O_131,N_14708,N_14006);
xor UO_132 (O_132,N_14868,N_14638);
and UO_133 (O_133,N_14824,N_14859);
or UO_134 (O_134,N_14100,N_14890);
nor UO_135 (O_135,N_14106,N_14942);
nor UO_136 (O_136,N_14895,N_14232);
nand UO_137 (O_137,N_14165,N_14980);
xnor UO_138 (O_138,N_14169,N_14578);
or UO_139 (O_139,N_14841,N_14087);
xnor UO_140 (O_140,N_14645,N_14989);
or UO_141 (O_141,N_14331,N_14781);
and UO_142 (O_142,N_14027,N_14556);
nor UO_143 (O_143,N_14349,N_14936);
or UO_144 (O_144,N_14347,N_14141);
nor UO_145 (O_145,N_14427,N_14503);
or UO_146 (O_146,N_14487,N_14484);
xnor UO_147 (O_147,N_14609,N_14756);
and UO_148 (O_148,N_14350,N_14571);
or UO_149 (O_149,N_14152,N_14595);
or UO_150 (O_150,N_14644,N_14287);
xor UO_151 (O_151,N_14731,N_14164);
or UO_152 (O_152,N_14513,N_14216);
and UO_153 (O_153,N_14083,N_14520);
xor UO_154 (O_154,N_14656,N_14594);
and UO_155 (O_155,N_14924,N_14517);
and UO_156 (O_156,N_14402,N_14754);
nand UO_157 (O_157,N_14981,N_14404);
or UO_158 (O_158,N_14553,N_14329);
nand UO_159 (O_159,N_14265,N_14790);
and UO_160 (O_160,N_14063,N_14995);
or UO_161 (O_161,N_14387,N_14612);
or UO_162 (O_162,N_14844,N_14200);
and UO_163 (O_163,N_14537,N_14692);
nor UO_164 (O_164,N_14195,N_14385);
nand UO_165 (O_165,N_14462,N_14109);
xnor UO_166 (O_166,N_14259,N_14096);
and UO_167 (O_167,N_14770,N_14110);
nand UO_168 (O_168,N_14463,N_14111);
nand UO_169 (O_169,N_14720,N_14986);
xor UO_170 (O_170,N_14941,N_14231);
xnor UO_171 (O_171,N_14923,N_14492);
and UO_172 (O_172,N_14706,N_14346);
nand UO_173 (O_173,N_14414,N_14020);
nor UO_174 (O_174,N_14032,N_14049);
xnor UO_175 (O_175,N_14381,N_14832);
or UO_176 (O_176,N_14722,N_14326);
or UO_177 (O_177,N_14140,N_14809);
nand UO_178 (O_178,N_14581,N_14531);
or UO_179 (O_179,N_14015,N_14560);
nor UO_180 (O_180,N_14745,N_14022);
nand UO_181 (O_181,N_14277,N_14961);
nor UO_182 (O_182,N_14069,N_14505);
nor UO_183 (O_183,N_14528,N_14897);
and UO_184 (O_184,N_14090,N_14663);
nor UO_185 (O_185,N_14501,N_14655);
nand UO_186 (O_186,N_14177,N_14597);
nand UO_187 (O_187,N_14899,N_14533);
or UO_188 (O_188,N_14519,N_14424);
xor UO_189 (O_189,N_14338,N_14763);
xnor UO_190 (O_190,N_14017,N_14450);
or UO_191 (O_191,N_14301,N_14369);
nand UO_192 (O_192,N_14957,N_14124);
nand UO_193 (O_193,N_14497,N_14997);
nand UO_194 (O_194,N_14148,N_14400);
or UO_195 (O_195,N_14278,N_14678);
or UO_196 (O_196,N_14717,N_14526);
xor UO_197 (O_197,N_14308,N_14475);
and UO_198 (O_198,N_14539,N_14793);
xor UO_199 (O_199,N_14816,N_14755);
or UO_200 (O_200,N_14432,N_14871);
xor UO_201 (O_201,N_14390,N_14686);
or UO_202 (O_202,N_14089,N_14541);
xnor UO_203 (O_203,N_14654,N_14270);
xnor UO_204 (O_204,N_14659,N_14545);
xnor UO_205 (O_205,N_14716,N_14166);
and UO_206 (O_206,N_14397,N_14392);
xor UO_207 (O_207,N_14186,N_14018);
nor UO_208 (O_208,N_14917,N_14819);
nand UO_209 (O_209,N_14230,N_14472);
xnor UO_210 (O_210,N_14696,N_14401);
xnor UO_211 (O_211,N_14690,N_14855);
and UO_212 (O_212,N_14250,N_14102);
and UO_213 (O_213,N_14193,N_14829);
nand UO_214 (O_214,N_14538,N_14268);
xor UO_215 (O_215,N_14939,N_14983);
or UO_216 (O_216,N_14808,N_14262);
nand UO_217 (O_217,N_14734,N_14078);
nor UO_218 (O_218,N_14411,N_14438);
nor UO_219 (O_219,N_14944,N_14764);
or UO_220 (O_220,N_14418,N_14721);
or UO_221 (O_221,N_14607,N_14081);
nand UO_222 (O_222,N_14904,N_14640);
nand UO_223 (O_223,N_14723,N_14321);
nand UO_224 (O_224,N_14576,N_14875);
or UO_225 (O_225,N_14546,N_14653);
nor UO_226 (O_226,N_14892,N_14235);
xor UO_227 (O_227,N_14159,N_14993);
or UO_228 (O_228,N_14702,N_14976);
xor UO_229 (O_229,N_14317,N_14361);
and UO_230 (O_230,N_14061,N_14469);
nand UO_231 (O_231,N_14434,N_14026);
xor UO_232 (O_232,N_14617,N_14984);
or UO_233 (O_233,N_14138,N_14204);
and UO_234 (O_234,N_14220,N_14348);
and UO_235 (O_235,N_14451,N_14911);
nand UO_236 (O_236,N_14448,N_14132);
and UO_237 (O_237,N_14552,N_14097);
and UO_238 (O_238,N_14675,N_14632);
nor UO_239 (O_239,N_14184,N_14147);
xnor UO_240 (O_240,N_14219,N_14283);
nor UO_241 (O_241,N_14311,N_14328);
nand UO_242 (O_242,N_14436,N_14626);
or UO_243 (O_243,N_14368,N_14873);
nand UO_244 (O_244,N_14785,N_14246);
nor UO_245 (O_245,N_14926,N_14666);
and UO_246 (O_246,N_14171,N_14646);
and UO_247 (O_247,N_14779,N_14668);
xnor UO_248 (O_248,N_14260,N_14098);
nor UO_249 (O_249,N_14922,N_14579);
nor UO_250 (O_250,N_14282,N_14766);
nor UO_251 (O_251,N_14502,N_14782);
nand UO_252 (O_252,N_14685,N_14342);
and UO_253 (O_253,N_14710,N_14228);
nor UO_254 (O_254,N_14012,N_14956);
and UO_255 (O_255,N_14426,N_14691);
xnor UO_256 (O_256,N_14562,N_14573);
nand UO_257 (O_257,N_14709,N_14000);
or UO_258 (O_258,N_14318,N_14953);
nand UO_259 (O_259,N_14601,N_14880);
or UO_260 (O_260,N_14371,N_14643);
or UO_261 (O_261,N_14786,N_14162);
nor UO_262 (O_262,N_14068,N_14035);
nand UO_263 (O_263,N_14679,N_14339);
and UO_264 (O_264,N_14799,N_14126);
nor UO_265 (O_265,N_14237,N_14276);
or UO_266 (O_266,N_14735,N_14215);
nor UO_267 (O_267,N_14951,N_14618);
or UO_268 (O_268,N_14094,N_14453);
and UO_269 (O_269,N_14352,N_14493);
nor UO_270 (O_270,N_14261,N_14674);
xor UO_271 (O_271,N_14622,N_14805);
nand UO_272 (O_272,N_14360,N_14439);
nand UO_273 (O_273,N_14807,N_14670);
nand UO_274 (O_274,N_14481,N_14179);
xnor UO_275 (O_275,N_14629,N_14740);
and UO_276 (O_276,N_14628,N_14120);
nand UO_277 (O_277,N_14131,N_14256);
or UO_278 (O_278,N_14529,N_14876);
and UO_279 (O_279,N_14928,N_14341);
or UO_280 (O_280,N_14038,N_14119);
or UO_281 (O_281,N_14857,N_14584);
or UO_282 (O_282,N_14635,N_14657);
and UO_283 (O_283,N_14608,N_14792);
nor UO_284 (O_284,N_14733,N_14610);
nor UO_285 (O_285,N_14606,N_14435);
nor UO_286 (O_286,N_14714,N_14285);
and UO_287 (O_287,N_14496,N_14946);
or UO_288 (O_288,N_14176,N_14687);
and UO_289 (O_289,N_14949,N_14076);
nand UO_290 (O_290,N_14930,N_14091);
nand UO_291 (O_291,N_14056,N_14445);
nand UO_292 (O_292,N_14778,N_14831);
or UO_293 (O_293,N_14621,N_14712);
xor UO_294 (O_294,N_14882,N_14323);
xnor UO_295 (O_295,N_14775,N_14364);
nand UO_296 (O_296,N_14549,N_14443);
nand UO_297 (O_297,N_14412,N_14479);
and UO_298 (O_298,N_14500,N_14491);
and UO_299 (O_299,N_14123,N_14572);
xnor UO_300 (O_300,N_14821,N_14739);
nand UO_301 (O_301,N_14431,N_14072);
and UO_302 (O_302,N_14319,N_14188);
or UO_303 (O_303,N_14486,N_14343);
or UO_304 (O_304,N_14642,N_14315);
xor UO_305 (O_305,N_14213,N_14101);
nand UO_306 (O_306,N_14744,N_14525);
nor UO_307 (O_307,N_14010,N_14267);
nor UO_308 (O_308,N_14470,N_14093);
or UO_309 (O_309,N_14473,N_14143);
nand UO_310 (O_310,N_14619,N_14955);
or UO_311 (O_311,N_14688,N_14704);
nand UO_312 (O_312,N_14408,N_14377);
nor UO_313 (O_313,N_14113,N_14175);
xor UO_314 (O_314,N_14482,N_14375);
nor UO_315 (O_315,N_14613,N_14521);
nand UO_316 (O_316,N_14586,N_14662);
or UO_317 (O_317,N_14833,N_14293);
nor UO_318 (O_318,N_14499,N_14066);
xnor UO_319 (O_319,N_14547,N_14210);
or UO_320 (O_320,N_14863,N_14466);
nor UO_321 (O_321,N_14214,N_14598);
nand UO_322 (O_322,N_14468,N_14419);
nand UO_323 (O_323,N_14830,N_14583);
nor UO_324 (O_324,N_14599,N_14885);
nand UO_325 (O_325,N_14620,N_14280);
and UO_326 (O_326,N_14718,N_14879);
and UO_327 (O_327,N_14295,N_14051);
or UO_328 (O_328,N_14605,N_14593);
or UO_329 (O_329,N_14962,N_14998);
nor UO_330 (O_330,N_14508,N_14070);
and UO_331 (O_331,N_14163,N_14945);
nand UO_332 (O_332,N_14067,N_14037);
or UO_333 (O_333,N_14103,N_14019);
nor UO_334 (O_334,N_14518,N_14370);
and UO_335 (O_335,N_14409,N_14429);
and UO_336 (O_336,N_14014,N_14016);
xnor UO_337 (O_337,N_14221,N_14818);
and UO_338 (O_338,N_14156,N_14564);
nor UO_339 (O_339,N_14724,N_14388);
and UO_340 (O_340,N_14893,N_14732);
nor UO_341 (O_341,N_14160,N_14209);
and UO_342 (O_342,N_14114,N_14194);
xnor UO_343 (O_343,N_14356,N_14191);
and UO_344 (O_344,N_14683,N_14028);
or UO_345 (O_345,N_14307,N_14797);
nor UO_346 (O_346,N_14765,N_14407);
nand UO_347 (O_347,N_14774,N_14866);
xor UO_348 (O_348,N_14289,N_14822);
and UO_349 (O_349,N_14198,N_14474);
nand UO_350 (O_350,N_14281,N_14378);
nor UO_351 (O_351,N_14698,N_14570);
xnor UO_352 (O_352,N_14585,N_14794);
nor UO_353 (O_353,N_14212,N_14596);
nand UO_354 (O_354,N_14940,N_14788);
and UO_355 (O_355,N_14415,N_14044);
or UO_356 (O_356,N_14241,N_14703);
or UO_357 (O_357,N_14254,N_14057);
xnor UO_358 (O_358,N_14864,N_14636);
or UO_359 (O_359,N_14884,N_14504);
and UO_360 (O_360,N_14396,N_14896);
xnor UO_361 (O_361,N_14548,N_14294);
nor UO_362 (O_362,N_14279,N_14891);
nand UO_363 (O_363,N_14725,N_14353);
nand UO_364 (O_364,N_14206,N_14682);
and UO_365 (O_365,N_14480,N_14759);
xnor UO_366 (O_366,N_14053,N_14987);
nor UO_367 (O_367,N_14004,N_14146);
and UO_368 (O_368,N_14290,N_14495);
nor UO_369 (O_369,N_14380,N_14509);
xnor UO_370 (O_370,N_14649,N_14174);
nor UO_371 (O_371,N_14363,N_14227);
nor UO_372 (O_372,N_14031,N_14305);
and UO_373 (O_373,N_14425,N_14391);
or UO_374 (O_374,N_14823,N_14836);
or UO_375 (O_375,N_14129,N_14117);
or UO_376 (O_376,N_14772,N_14395);
xnor UO_377 (O_377,N_14908,N_14631);
xor UO_378 (O_378,N_14847,N_14009);
xnor UO_379 (O_379,N_14154,N_14055);
nor UO_380 (O_380,N_14602,N_14727);
or UO_381 (O_381,N_14567,N_14359);
xnor UO_382 (O_382,N_14872,N_14577);
or UO_383 (O_383,N_14780,N_14441);
xor UO_384 (O_384,N_14676,N_14224);
and UO_385 (O_385,N_14582,N_14379);
and UO_386 (O_386,N_14047,N_14964);
xnor UO_387 (O_387,N_14271,N_14258);
and UO_388 (O_388,N_14914,N_14623);
nor UO_389 (O_389,N_14312,N_14272);
or UO_390 (O_390,N_14749,N_14999);
nand UO_391 (O_391,N_14534,N_14178);
xor UO_392 (O_392,N_14145,N_14699);
xor UO_393 (O_393,N_14322,N_14742);
nand UO_394 (O_394,N_14243,N_14217);
and UO_395 (O_395,N_14771,N_14105);
and UO_396 (O_396,N_14677,N_14442);
xnor UO_397 (O_397,N_14641,N_14136);
nor UO_398 (O_398,N_14244,N_14366);
and UO_399 (O_399,N_14900,N_14919);
xor UO_400 (O_400,N_14413,N_14743);
xnor UO_401 (O_401,N_14968,N_14309);
nand UO_402 (O_402,N_14060,N_14802);
nor UO_403 (O_403,N_14798,N_14947);
nor UO_404 (O_404,N_14862,N_14182);
xor UO_405 (O_405,N_14292,N_14729);
nor UO_406 (O_406,N_14753,N_14664);
nor UO_407 (O_407,N_14373,N_14456);
or UO_408 (O_408,N_14477,N_14440);
or UO_409 (O_409,N_14008,N_14249);
xnor UO_410 (O_410,N_14761,N_14747);
and UO_411 (O_411,N_14108,N_14002);
nand UO_412 (O_412,N_14647,N_14530);
or UO_413 (O_413,N_14787,N_14255);
nor UO_414 (O_414,N_14297,N_14269);
xor UO_415 (O_415,N_14700,N_14218);
nor UO_416 (O_416,N_14996,N_14007);
nand UO_417 (O_417,N_14039,N_14806);
and UO_418 (O_418,N_14483,N_14902);
nor UO_419 (O_419,N_14033,N_14853);
xor UO_420 (O_420,N_14965,N_14544);
nor UO_421 (O_421,N_14850,N_14211);
nand UO_422 (O_422,N_14587,N_14898);
xor UO_423 (O_423,N_14810,N_14421);
and UO_424 (O_424,N_14158,N_14107);
or UO_425 (O_425,N_14839,N_14600);
and UO_426 (O_426,N_14042,N_14684);
nand UO_427 (O_427,N_14694,N_14982);
nor UO_428 (O_428,N_14846,N_14134);
xor UO_429 (O_429,N_14569,N_14406);
xor UO_430 (O_430,N_14937,N_14826);
nand UO_431 (O_431,N_14510,N_14532);
nand UO_432 (O_432,N_14075,N_14454);
nand UO_433 (O_433,N_14565,N_14403);
and UO_434 (O_434,N_14257,N_14488);
xor UO_435 (O_435,N_14398,N_14935);
or UO_436 (O_436,N_14116,N_14374);
nand UO_437 (O_437,N_14284,N_14563);
xnor UO_438 (O_438,N_14190,N_14811);
nand UO_439 (O_439,N_14803,N_14768);
and UO_440 (O_440,N_14325,N_14507);
or UO_441 (O_441,N_14769,N_14405);
xnor UO_442 (O_442,N_14903,N_14776);
or UO_443 (O_443,N_14274,N_14197);
or UO_444 (O_444,N_14760,N_14625);
or UO_445 (O_445,N_14199,N_14430);
and UO_446 (O_446,N_14185,N_14036);
and UO_447 (O_447,N_14455,N_14959);
xnor UO_448 (O_448,N_14652,N_14376);
nor UO_449 (O_449,N_14883,N_14748);
and UO_450 (O_450,N_14251,N_14535);
nand UO_451 (O_451,N_14762,N_14550);
nand UO_452 (O_452,N_14062,N_14130);
xor UO_453 (O_453,N_14428,N_14952);
and UO_454 (O_454,N_14248,N_14555);
nand UO_455 (O_455,N_14557,N_14452);
nor UO_456 (O_456,N_14345,N_14960);
nand UO_457 (O_457,N_14827,N_14658);
or UO_458 (O_458,N_14726,N_14767);
nor UO_459 (O_459,N_14515,N_14907);
xor UO_460 (O_460,N_14975,N_14845);
nor UO_461 (O_461,N_14661,N_14713);
xor UO_462 (O_462,N_14927,N_14245);
and UO_463 (O_463,N_14383,N_14842);
xnor UO_464 (O_464,N_14874,N_14233);
nor UO_465 (O_465,N_14052,N_14921);
nor UO_466 (O_466,N_14266,N_14208);
or UO_467 (O_467,N_14693,N_14639);
nand UO_468 (O_468,N_14978,N_14168);
nor UO_469 (O_469,N_14306,N_14416);
nand UO_470 (O_470,N_14746,N_14948);
xnor UO_471 (O_471,N_14834,N_14672);
and UO_472 (O_472,N_14865,N_14604);
nand UO_473 (O_473,N_14043,N_14386);
and UO_474 (O_474,N_14542,N_14074);
and UO_475 (O_475,N_14861,N_14901);
and UO_476 (O_476,N_14860,N_14695);
xnor UO_477 (O_477,N_14449,N_14144);
nor UO_478 (O_478,N_14151,N_14457);
or UO_479 (O_479,N_14086,N_14540);
nor UO_480 (O_480,N_14804,N_14242);
nand UO_481 (O_481,N_14354,N_14648);
xnor UO_482 (O_482,N_14273,N_14084);
or UO_483 (O_483,N_14300,N_14115);
and UO_484 (O_484,N_14181,N_14337);
xnor UO_485 (O_485,N_14041,N_14362);
nand UO_486 (O_486,N_14320,N_14878);
and UO_487 (O_487,N_14240,N_14843);
or UO_488 (O_488,N_14365,N_14054);
or UO_489 (O_489,N_14498,N_14149);
nor UO_490 (O_490,N_14382,N_14229);
or UO_491 (O_491,N_14048,N_14931);
nor UO_492 (O_492,N_14512,N_14979);
nor UO_493 (O_493,N_14088,N_14304);
xnor UO_494 (O_494,N_14854,N_14422);
xnor UO_495 (O_495,N_14561,N_14264);
or UO_496 (O_496,N_14950,N_14869);
xor UO_497 (O_497,N_14932,N_14183);
or UO_498 (O_498,N_14633,N_14580);
xor UO_499 (O_499,N_14730,N_14071);
or UO_500 (O_500,N_14040,N_14987);
xnor UO_501 (O_501,N_14201,N_14348);
and UO_502 (O_502,N_14865,N_14084);
or UO_503 (O_503,N_14334,N_14317);
and UO_504 (O_504,N_14464,N_14369);
nor UO_505 (O_505,N_14832,N_14800);
xor UO_506 (O_506,N_14825,N_14380);
nand UO_507 (O_507,N_14396,N_14868);
nand UO_508 (O_508,N_14776,N_14997);
or UO_509 (O_509,N_14011,N_14484);
nor UO_510 (O_510,N_14036,N_14435);
nand UO_511 (O_511,N_14803,N_14065);
xnor UO_512 (O_512,N_14241,N_14062);
nor UO_513 (O_513,N_14622,N_14628);
nor UO_514 (O_514,N_14745,N_14030);
nor UO_515 (O_515,N_14310,N_14967);
or UO_516 (O_516,N_14478,N_14704);
or UO_517 (O_517,N_14507,N_14182);
or UO_518 (O_518,N_14634,N_14826);
nand UO_519 (O_519,N_14877,N_14393);
and UO_520 (O_520,N_14223,N_14649);
and UO_521 (O_521,N_14069,N_14496);
nand UO_522 (O_522,N_14029,N_14849);
or UO_523 (O_523,N_14598,N_14028);
and UO_524 (O_524,N_14472,N_14964);
nor UO_525 (O_525,N_14093,N_14593);
or UO_526 (O_526,N_14314,N_14193);
xor UO_527 (O_527,N_14862,N_14157);
nand UO_528 (O_528,N_14599,N_14036);
nor UO_529 (O_529,N_14908,N_14055);
nand UO_530 (O_530,N_14436,N_14719);
xor UO_531 (O_531,N_14962,N_14280);
or UO_532 (O_532,N_14481,N_14202);
xor UO_533 (O_533,N_14597,N_14695);
nor UO_534 (O_534,N_14763,N_14952);
xor UO_535 (O_535,N_14656,N_14086);
and UO_536 (O_536,N_14459,N_14326);
and UO_537 (O_537,N_14935,N_14663);
nand UO_538 (O_538,N_14264,N_14349);
and UO_539 (O_539,N_14954,N_14615);
and UO_540 (O_540,N_14675,N_14144);
nand UO_541 (O_541,N_14317,N_14789);
nor UO_542 (O_542,N_14453,N_14989);
and UO_543 (O_543,N_14569,N_14250);
and UO_544 (O_544,N_14653,N_14948);
xnor UO_545 (O_545,N_14075,N_14439);
and UO_546 (O_546,N_14360,N_14705);
xnor UO_547 (O_547,N_14924,N_14897);
or UO_548 (O_548,N_14536,N_14449);
xnor UO_549 (O_549,N_14927,N_14216);
nor UO_550 (O_550,N_14401,N_14954);
or UO_551 (O_551,N_14258,N_14052);
nor UO_552 (O_552,N_14154,N_14283);
xor UO_553 (O_553,N_14233,N_14248);
and UO_554 (O_554,N_14591,N_14278);
nand UO_555 (O_555,N_14418,N_14029);
or UO_556 (O_556,N_14831,N_14477);
xnor UO_557 (O_557,N_14128,N_14883);
nor UO_558 (O_558,N_14525,N_14153);
or UO_559 (O_559,N_14646,N_14730);
and UO_560 (O_560,N_14327,N_14569);
and UO_561 (O_561,N_14534,N_14129);
and UO_562 (O_562,N_14093,N_14981);
nand UO_563 (O_563,N_14213,N_14559);
nor UO_564 (O_564,N_14294,N_14613);
xnor UO_565 (O_565,N_14000,N_14703);
or UO_566 (O_566,N_14462,N_14705);
and UO_567 (O_567,N_14192,N_14283);
nand UO_568 (O_568,N_14412,N_14563);
nor UO_569 (O_569,N_14545,N_14546);
nor UO_570 (O_570,N_14983,N_14929);
or UO_571 (O_571,N_14847,N_14855);
xnor UO_572 (O_572,N_14297,N_14261);
nor UO_573 (O_573,N_14224,N_14272);
nor UO_574 (O_574,N_14453,N_14403);
nor UO_575 (O_575,N_14973,N_14047);
nor UO_576 (O_576,N_14259,N_14137);
nand UO_577 (O_577,N_14515,N_14791);
nor UO_578 (O_578,N_14673,N_14922);
nand UO_579 (O_579,N_14914,N_14017);
nand UO_580 (O_580,N_14700,N_14785);
or UO_581 (O_581,N_14040,N_14825);
nand UO_582 (O_582,N_14037,N_14775);
nor UO_583 (O_583,N_14414,N_14990);
or UO_584 (O_584,N_14573,N_14574);
nor UO_585 (O_585,N_14095,N_14838);
nand UO_586 (O_586,N_14854,N_14047);
and UO_587 (O_587,N_14970,N_14176);
xor UO_588 (O_588,N_14372,N_14490);
xnor UO_589 (O_589,N_14238,N_14287);
and UO_590 (O_590,N_14571,N_14312);
and UO_591 (O_591,N_14061,N_14515);
nand UO_592 (O_592,N_14905,N_14326);
and UO_593 (O_593,N_14303,N_14677);
xnor UO_594 (O_594,N_14936,N_14869);
nand UO_595 (O_595,N_14452,N_14034);
xor UO_596 (O_596,N_14229,N_14550);
nand UO_597 (O_597,N_14069,N_14094);
and UO_598 (O_598,N_14855,N_14197);
or UO_599 (O_599,N_14748,N_14317);
or UO_600 (O_600,N_14802,N_14457);
nor UO_601 (O_601,N_14568,N_14409);
nor UO_602 (O_602,N_14181,N_14468);
xor UO_603 (O_603,N_14469,N_14589);
nor UO_604 (O_604,N_14796,N_14747);
and UO_605 (O_605,N_14759,N_14487);
or UO_606 (O_606,N_14495,N_14221);
xor UO_607 (O_607,N_14075,N_14850);
or UO_608 (O_608,N_14833,N_14277);
nand UO_609 (O_609,N_14961,N_14216);
or UO_610 (O_610,N_14215,N_14128);
and UO_611 (O_611,N_14397,N_14587);
nand UO_612 (O_612,N_14412,N_14072);
and UO_613 (O_613,N_14730,N_14604);
xnor UO_614 (O_614,N_14715,N_14161);
xnor UO_615 (O_615,N_14050,N_14997);
nor UO_616 (O_616,N_14149,N_14088);
and UO_617 (O_617,N_14849,N_14756);
or UO_618 (O_618,N_14985,N_14356);
or UO_619 (O_619,N_14007,N_14547);
nand UO_620 (O_620,N_14414,N_14842);
and UO_621 (O_621,N_14928,N_14315);
or UO_622 (O_622,N_14519,N_14984);
or UO_623 (O_623,N_14074,N_14917);
and UO_624 (O_624,N_14490,N_14988);
xor UO_625 (O_625,N_14214,N_14615);
xor UO_626 (O_626,N_14423,N_14129);
nand UO_627 (O_627,N_14249,N_14516);
or UO_628 (O_628,N_14516,N_14117);
nand UO_629 (O_629,N_14361,N_14669);
nand UO_630 (O_630,N_14679,N_14976);
nor UO_631 (O_631,N_14081,N_14590);
nand UO_632 (O_632,N_14978,N_14995);
nor UO_633 (O_633,N_14510,N_14638);
nand UO_634 (O_634,N_14013,N_14374);
nand UO_635 (O_635,N_14401,N_14145);
xor UO_636 (O_636,N_14821,N_14126);
xor UO_637 (O_637,N_14334,N_14969);
nand UO_638 (O_638,N_14819,N_14755);
xor UO_639 (O_639,N_14909,N_14312);
and UO_640 (O_640,N_14785,N_14670);
nor UO_641 (O_641,N_14010,N_14813);
xor UO_642 (O_642,N_14800,N_14770);
or UO_643 (O_643,N_14756,N_14764);
or UO_644 (O_644,N_14207,N_14406);
nor UO_645 (O_645,N_14559,N_14199);
xnor UO_646 (O_646,N_14575,N_14626);
xor UO_647 (O_647,N_14761,N_14515);
and UO_648 (O_648,N_14847,N_14076);
nand UO_649 (O_649,N_14400,N_14247);
xor UO_650 (O_650,N_14874,N_14340);
nand UO_651 (O_651,N_14217,N_14804);
nand UO_652 (O_652,N_14296,N_14249);
xnor UO_653 (O_653,N_14754,N_14289);
nor UO_654 (O_654,N_14002,N_14525);
xnor UO_655 (O_655,N_14011,N_14702);
nor UO_656 (O_656,N_14903,N_14444);
xnor UO_657 (O_657,N_14982,N_14658);
xnor UO_658 (O_658,N_14707,N_14222);
or UO_659 (O_659,N_14461,N_14962);
or UO_660 (O_660,N_14610,N_14572);
nand UO_661 (O_661,N_14134,N_14776);
or UO_662 (O_662,N_14884,N_14110);
xnor UO_663 (O_663,N_14130,N_14518);
nand UO_664 (O_664,N_14469,N_14872);
nor UO_665 (O_665,N_14194,N_14168);
xor UO_666 (O_666,N_14277,N_14629);
nor UO_667 (O_667,N_14929,N_14026);
and UO_668 (O_668,N_14240,N_14395);
and UO_669 (O_669,N_14585,N_14201);
or UO_670 (O_670,N_14963,N_14683);
or UO_671 (O_671,N_14157,N_14549);
and UO_672 (O_672,N_14743,N_14855);
nor UO_673 (O_673,N_14469,N_14448);
nor UO_674 (O_674,N_14927,N_14145);
nand UO_675 (O_675,N_14269,N_14314);
and UO_676 (O_676,N_14897,N_14237);
or UO_677 (O_677,N_14126,N_14308);
or UO_678 (O_678,N_14645,N_14222);
nor UO_679 (O_679,N_14556,N_14891);
or UO_680 (O_680,N_14620,N_14656);
xor UO_681 (O_681,N_14086,N_14676);
or UO_682 (O_682,N_14193,N_14489);
nand UO_683 (O_683,N_14658,N_14529);
nor UO_684 (O_684,N_14017,N_14115);
nor UO_685 (O_685,N_14462,N_14092);
nor UO_686 (O_686,N_14381,N_14314);
nor UO_687 (O_687,N_14168,N_14320);
and UO_688 (O_688,N_14704,N_14839);
and UO_689 (O_689,N_14177,N_14875);
nor UO_690 (O_690,N_14692,N_14620);
nor UO_691 (O_691,N_14094,N_14763);
and UO_692 (O_692,N_14045,N_14044);
and UO_693 (O_693,N_14366,N_14973);
and UO_694 (O_694,N_14845,N_14392);
or UO_695 (O_695,N_14324,N_14368);
and UO_696 (O_696,N_14750,N_14257);
nor UO_697 (O_697,N_14894,N_14923);
and UO_698 (O_698,N_14896,N_14979);
xor UO_699 (O_699,N_14686,N_14779);
or UO_700 (O_700,N_14788,N_14957);
xnor UO_701 (O_701,N_14603,N_14235);
nor UO_702 (O_702,N_14768,N_14328);
or UO_703 (O_703,N_14607,N_14401);
or UO_704 (O_704,N_14506,N_14462);
nand UO_705 (O_705,N_14888,N_14882);
nand UO_706 (O_706,N_14418,N_14566);
nor UO_707 (O_707,N_14811,N_14289);
and UO_708 (O_708,N_14988,N_14593);
nor UO_709 (O_709,N_14119,N_14238);
nor UO_710 (O_710,N_14116,N_14524);
nand UO_711 (O_711,N_14787,N_14446);
xnor UO_712 (O_712,N_14999,N_14007);
xnor UO_713 (O_713,N_14099,N_14280);
nor UO_714 (O_714,N_14998,N_14652);
xnor UO_715 (O_715,N_14291,N_14792);
nor UO_716 (O_716,N_14549,N_14219);
xor UO_717 (O_717,N_14905,N_14555);
nor UO_718 (O_718,N_14822,N_14567);
xor UO_719 (O_719,N_14419,N_14488);
nand UO_720 (O_720,N_14835,N_14401);
and UO_721 (O_721,N_14869,N_14817);
and UO_722 (O_722,N_14019,N_14520);
and UO_723 (O_723,N_14728,N_14064);
and UO_724 (O_724,N_14555,N_14579);
xnor UO_725 (O_725,N_14994,N_14225);
or UO_726 (O_726,N_14546,N_14652);
nor UO_727 (O_727,N_14683,N_14728);
nand UO_728 (O_728,N_14612,N_14238);
or UO_729 (O_729,N_14491,N_14023);
and UO_730 (O_730,N_14055,N_14291);
nor UO_731 (O_731,N_14493,N_14334);
nor UO_732 (O_732,N_14766,N_14226);
nand UO_733 (O_733,N_14141,N_14006);
nand UO_734 (O_734,N_14301,N_14297);
nand UO_735 (O_735,N_14127,N_14920);
nor UO_736 (O_736,N_14224,N_14821);
xnor UO_737 (O_737,N_14228,N_14167);
nor UO_738 (O_738,N_14784,N_14594);
xnor UO_739 (O_739,N_14349,N_14661);
xnor UO_740 (O_740,N_14764,N_14493);
nand UO_741 (O_741,N_14352,N_14000);
and UO_742 (O_742,N_14867,N_14031);
nand UO_743 (O_743,N_14974,N_14960);
nand UO_744 (O_744,N_14423,N_14300);
and UO_745 (O_745,N_14568,N_14510);
and UO_746 (O_746,N_14254,N_14899);
and UO_747 (O_747,N_14462,N_14722);
or UO_748 (O_748,N_14140,N_14093);
xor UO_749 (O_749,N_14831,N_14434);
nor UO_750 (O_750,N_14333,N_14867);
or UO_751 (O_751,N_14989,N_14278);
or UO_752 (O_752,N_14428,N_14707);
nor UO_753 (O_753,N_14274,N_14689);
and UO_754 (O_754,N_14363,N_14519);
xor UO_755 (O_755,N_14005,N_14413);
xor UO_756 (O_756,N_14765,N_14215);
nor UO_757 (O_757,N_14059,N_14100);
xnor UO_758 (O_758,N_14498,N_14403);
nand UO_759 (O_759,N_14512,N_14651);
xnor UO_760 (O_760,N_14922,N_14857);
nor UO_761 (O_761,N_14530,N_14484);
or UO_762 (O_762,N_14841,N_14723);
and UO_763 (O_763,N_14376,N_14063);
xnor UO_764 (O_764,N_14598,N_14001);
xor UO_765 (O_765,N_14635,N_14717);
and UO_766 (O_766,N_14301,N_14266);
xor UO_767 (O_767,N_14943,N_14340);
or UO_768 (O_768,N_14142,N_14381);
or UO_769 (O_769,N_14198,N_14764);
and UO_770 (O_770,N_14922,N_14441);
xor UO_771 (O_771,N_14227,N_14711);
or UO_772 (O_772,N_14067,N_14043);
nand UO_773 (O_773,N_14389,N_14814);
nand UO_774 (O_774,N_14424,N_14765);
and UO_775 (O_775,N_14327,N_14686);
or UO_776 (O_776,N_14434,N_14642);
nor UO_777 (O_777,N_14192,N_14700);
nand UO_778 (O_778,N_14109,N_14434);
nand UO_779 (O_779,N_14123,N_14624);
nand UO_780 (O_780,N_14246,N_14925);
xor UO_781 (O_781,N_14803,N_14174);
nand UO_782 (O_782,N_14942,N_14231);
nor UO_783 (O_783,N_14823,N_14898);
xnor UO_784 (O_784,N_14515,N_14745);
and UO_785 (O_785,N_14344,N_14863);
or UO_786 (O_786,N_14688,N_14107);
nor UO_787 (O_787,N_14275,N_14180);
nand UO_788 (O_788,N_14654,N_14040);
and UO_789 (O_789,N_14002,N_14114);
or UO_790 (O_790,N_14156,N_14965);
or UO_791 (O_791,N_14279,N_14228);
nand UO_792 (O_792,N_14344,N_14925);
nand UO_793 (O_793,N_14344,N_14023);
xor UO_794 (O_794,N_14899,N_14716);
or UO_795 (O_795,N_14598,N_14712);
or UO_796 (O_796,N_14041,N_14485);
nand UO_797 (O_797,N_14039,N_14909);
xor UO_798 (O_798,N_14713,N_14560);
or UO_799 (O_799,N_14247,N_14197);
and UO_800 (O_800,N_14271,N_14804);
or UO_801 (O_801,N_14966,N_14092);
or UO_802 (O_802,N_14440,N_14248);
nand UO_803 (O_803,N_14925,N_14659);
or UO_804 (O_804,N_14968,N_14306);
or UO_805 (O_805,N_14450,N_14423);
xor UO_806 (O_806,N_14149,N_14900);
nor UO_807 (O_807,N_14460,N_14387);
nor UO_808 (O_808,N_14120,N_14253);
and UO_809 (O_809,N_14389,N_14686);
nand UO_810 (O_810,N_14951,N_14751);
and UO_811 (O_811,N_14380,N_14379);
or UO_812 (O_812,N_14212,N_14789);
or UO_813 (O_813,N_14953,N_14965);
xor UO_814 (O_814,N_14843,N_14460);
or UO_815 (O_815,N_14815,N_14256);
and UO_816 (O_816,N_14022,N_14224);
or UO_817 (O_817,N_14018,N_14249);
xor UO_818 (O_818,N_14525,N_14559);
and UO_819 (O_819,N_14925,N_14366);
and UO_820 (O_820,N_14771,N_14686);
nor UO_821 (O_821,N_14235,N_14312);
or UO_822 (O_822,N_14093,N_14513);
nand UO_823 (O_823,N_14834,N_14582);
and UO_824 (O_824,N_14640,N_14663);
xnor UO_825 (O_825,N_14872,N_14506);
nor UO_826 (O_826,N_14146,N_14661);
xnor UO_827 (O_827,N_14449,N_14202);
nand UO_828 (O_828,N_14727,N_14480);
nor UO_829 (O_829,N_14619,N_14043);
xnor UO_830 (O_830,N_14991,N_14456);
nand UO_831 (O_831,N_14675,N_14233);
or UO_832 (O_832,N_14768,N_14281);
xor UO_833 (O_833,N_14360,N_14704);
and UO_834 (O_834,N_14193,N_14903);
nor UO_835 (O_835,N_14079,N_14006);
nand UO_836 (O_836,N_14998,N_14841);
and UO_837 (O_837,N_14995,N_14084);
nor UO_838 (O_838,N_14159,N_14247);
nand UO_839 (O_839,N_14767,N_14935);
xnor UO_840 (O_840,N_14096,N_14123);
nand UO_841 (O_841,N_14345,N_14552);
or UO_842 (O_842,N_14556,N_14906);
xnor UO_843 (O_843,N_14437,N_14961);
xor UO_844 (O_844,N_14337,N_14591);
nand UO_845 (O_845,N_14361,N_14904);
xor UO_846 (O_846,N_14840,N_14386);
and UO_847 (O_847,N_14346,N_14909);
nand UO_848 (O_848,N_14623,N_14434);
xnor UO_849 (O_849,N_14969,N_14543);
or UO_850 (O_850,N_14685,N_14073);
and UO_851 (O_851,N_14868,N_14216);
nor UO_852 (O_852,N_14203,N_14688);
nor UO_853 (O_853,N_14449,N_14511);
xnor UO_854 (O_854,N_14173,N_14439);
or UO_855 (O_855,N_14438,N_14088);
nor UO_856 (O_856,N_14856,N_14961);
and UO_857 (O_857,N_14836,N_14080);
nor UO_858 (O_858,N_14578,N_14416);
nand UO_859 (O_859,N_14461,N_14043);
nand UO_860 (O_860,N_14165,N_14178);
nor UO_861 (O_861,N_14646,N_14938);
xor UO_862 (O_862,N_14609,N_14788);
and UO_863 (O_863,N_14215,N_14028);
nor UO_864 (O_864,N_14148,N_14576);
or UO_865 (O_865,N_14506,N_14813);
and UO_866 (O_866,N_14027,N_14922);
nand UO_867 (O_867,N_14016,N_14419);
nand UO_868 (O_868,N_14924,N_14934);
nor UO_869 (O_869,N_14491,N_14177);
and UO_870 (O_870,N_14416,N_14561);
and UO_871 (O_871,N_14177,N_14605);
and UO_872 (O_872,N_14826,N_14284);
xnor UO_873 (O_873,N_14090,N_14092);
nand UO_874 (O_874,N_14533,N_14535);
nor UO_875 (O_875,N_14993,N_14918);
or UO_876 (O_876,N_14552,N_14678);
xnor UO_877 (O_877,N_14369,N_14172);
or UO_878 (O_878,N_14761,N_14179);
nand UO_879 (O_879,N_14954,N_14652);
and UO_880 (O_880,N_14132,N_14136);
or UO_881 (O_881,N_14405,N_14039);
and UO_882 (O_882,N_14982,N_14728);
xor UO_883 (O_883,N_14509,N_14845);
and UO_884 (O_884,N_14017,N_14297);
nand UO_885 (O_885,N_14237,N_14636);
nor UO_886 (O_886,N_14917,N_14751);
nand UO_887 (O_887,N_14407,N_14981);
nand UO_888 (O_888,N_14213,N_14890);
nor UO_889 (O_889,N_14726,N_14210);
and UO_890 (O_890,N_14821,N_14249);
or UO_891 (O_891,N_14358,N_14829);
nand UO_892 (O_892,N_14037,N_14141);
or UO_893 (O_893,N_14047,N_14941);
and UO_894 (O_894,N_14424,N_14660);
xor UO_895 (O_895,N_14453,N_14381);
nor UO_896 (O_896,N_14458,N_14110);
nand UO_897 (O_897,N_14187,N_14049);
xor UO_898 (O_898,N_14135,N_14115);
xor UO_899 (O_899,N_14362,N_14890);
and UO_900 (O_900,N_14364,N_14740);
xnor UO_901 (O_901,N_14459,N_14421);
and UO_902 (O_902,N_14636,N_14700);
and UO_903 (O_903,N_14655,N_14620);
or UO_904 (O_904,N_14723,N_14373);
and UO_905 (O_905,N_14936,N_14694);
or UO_906 (O_906,N_14022,N_14972);
nor UO_907 (O_907,N_14357,N_14050);
and UO_908 (O_908,N_14183,N_14232);
nor UO_909 (O_909,N_14329,N_14171);
nor UO_910 (O_910,N_14453,N_14709);
or UO_911 (O_911,N_14319,N_14457);
or UO_912 (O_912,N_14851,N_14053);
nor UO_913 (O_913,N_14374,N_14918);
or UO_914 (O_914,N_14687,N_14669);
or UO_915 (O_915,N_14449,N_14049);
nor UO_916 (O_916,N_14828,N_14142);
xor UO_917 (O_917,N_14075,N_14727);
or UO_918 (O_918,N_14789,N_14724);
or UO_919 (O_919,N_14436,N_14859);
and UO_920 (O_920,N_14617,N_14856);
nand UO_921 (O_921,N_14208,N_14095);
nor UO_922 (O_922,N_14617,N_14342);
xnor UO_923 (O_923,N_14847,N_14115);
nand UO_924 (O_924,N_14622,N_14599);
nor UO_925 (O_925,N_14442,N_14356);
and UO_926 (O_926,N_14548,N_14920);
and UO_927 (O_927,N_14553,N_14140);
nand UO_928 (O_928,N_14471,N_14389);
nor UO_929 (O_929,N_14116,N_14267);
or UO_930 (O_930,N_14012,N_14518);
or UO_931 (O_931,N_14547,N_14319);
nor UO_932 (O_932,N_14330,N_14955);
nand UO_933 (O_933,N_14139,N_14548);
or UO_934 (O_934,N_14101,N_14288);
nand UO_935 (O_935,N_14637,N_14253);
or UO_936 (O_936,N_14628,N_14848);
xnor UO_937 (O_937,N_14917,N_14389);
and UO_938 (O_938,N_14874,N_14056);
nor UO_939 (O_939,N_14584,N_14711);
or UO_940 (O_940,N_14054,N_14486);
xor UO_941 (O_941,N_14626,N_14916);
or UO_942 (O_942,N_14606,N_14632);
xnor UO_943 (O_943,N_14657,N_14929);
or UO_944 (O_944,N_14537,N_14001);
xor UO_945 (O_945,N_14195,N_14076);
xnor UO_946 (O_946,N_14528,N_14844);
xor UO_947 (O_947,N_14264,N_14175);
nor UO_948 (O_948,N_14357,N_14421);
nand UO_949 (O_949,N_14772,N_14671);
or UO_950 (O_950,N_14480,N_14484);
and UO_951 (O_951,N_14694,N_14551);
and UO_952 (O_952,N_14569,N_14137);
or UO_953 (O_953,N_14401,N_14249);
nand UO_954 (O_954,N_14045,N_14916);
nand UO_955 (O_955,N_14954,N_14818);
and UO_956 (O_956,N_14308,N_14521);
xor UO_957 (O_957,N_14315,N_14593);
or UO_958 (O_958,N_14303,N_14567);
nor UO_959 (O_959,N_14089,N_14287);
or UO_960 (O_960,N_14497,N_14442);
or UO_961 (O_961,N_14785,N_14412);
nand UO_962 (O_962,N_14693,N_14636);
or UO_963 (O_963,N_14366,N_14822);
nand UO_964 (O_964,N_14676,N_14408);
and UO_965 (O_965,N_14844,N_14986);
and UO_966 (O_966,N_14430,N_14257);
nand UO_967 (O_967,N_14147,N_14154);
nand UO_968 (O_968,N_14814,N_14486);
and UO_969 (O_969,N_14202,N_14385);
nor UO_970 (O_970,N_14525,N_14618);
and UO_971 (O_971,N_14418,N_14944);
xnor UO_972 (O_972,N_14548,N_14338);
or UO_973 (O_973,N_14429,N_14196);
or UO_974 (O_974,N_14415,N_14555);
or UO_975 (O_975,N_14552,N_14180);
nor UO_976 (O_976,N_14926,N_14134);
xnor UO_977 (O_977,N_14543,N_14322);
or UO_978 (O_978,N_14629,N_14143);
or UO_979 (O_979,N_14997,N_14185);
or UO_980 (O_980,N_14438,N_14993);
nand UO_981 (O_981,N_14629,N_14334);
xnor UO_982 (O_982,N_14895,N_14339);
nor UO_983 (O_983,N_14839,N_14788);
nor UO_984 (O_984,N_14194,N_14516);
nor UO_985 (O_985,N_14586,N_14834);
or UO_986 (O_986,N_14163,N_14720);
nand UO_987 (O_987,N_14014,N_14513);
xor UO_988 (O_988,N_14503,N_14590);
xor UO_989 (O_989,N_14946,N_14049);
and UO_990 (O_990,N_14341,N_14122);
nand UO_991 (O_991,N_14414,N_14115);
nor UO_992 (O_992,N_14276,N_14073);
xnor UO_993 (O_993,N_14593,N_14926);
nor UO_994 (O_994,N_14607,N_14546);
nand UO_995 (O_995,N_14969,N_14353);
and UO_996 (O_996,N_14987,N_14420);
and UO_997 (O_997,N_14778,N_14299);
and UO_998 (O_998,N_14275,N_14671);
and UO_999 (O_999,N_14899,N_14100);
nand UO_1000 (O_1000,N_14005,N_14845);
nand UO_1001 (O_1001,N_14385,N_14554);
and UO_1002 (O_1002,N_14043,N_14197);
and UO_1003 (O_1003,N_14866,N_14791);
and UO_1004 (O_1004,N_14273,N_14830);
xor UO_1005 (O_1005,N_14254,N_14837);
nand UO_1006 (O_1006,N_14809,N_14981);
nor UO_1007 (O_1007,N_14321,N_14592);
or UO_1008 (O_1008,N_14625,N_14147);
nor UO_1009 (O_1009,N_14522,N_14376);
nor UO_1010 (O_1010,N_14063,N_14160);
and UO_1011 (O_1011,N_14102,N_14911);
and UO_1012 (O_1012,N_14847,N_14705);
nand UO_1013 (O_1013,N_14539,N_14649);
and UO_1014 (O_1014,N_14468,N_14434);
xnor UO_1015 (O_1015,N_14897,N_14756);
nor UO_1016 (O_1016,N_14536,N_14791);
nor UO_1017 (O_1017,N_14957,N_14085);
nor UO_1018 (O_1018,N_14041,N_14773);
nor UO_1019 (O_1019,N_14878,N_14702);
nor UO_1020 (O_1020,N_14827,N_14167);
or UO_1021 (O_1021,N_14250,N_14285);
nand UO_1022 (O_1022,N_14275,N_14814);
nand UO_1023 (O_1023,N_14512,N_14454);
nand UO_1024 (O_1024,N_14699,N_14628);
and UO_1025 (O_1025,N_14073,N_14693);
xnor UO_1026 (O_1026,N_14056,N_14128);
nand UO_1027 (O_1027,N_14425,N_14205);
and UO_1028 (O_1028,N_14356,N_14647);
xnor UO_1029 (O_1029,N_14253,N_14492);
xnor UO_1030 (O_1030,N_14707,N_14010);
xor UO_1031 (O_1031,N_14776,N_14779);
xnor UO_1032 (O_1032,N_14706,N_14642);
xor UO_1033 (O_1033,N_14580,N_14256);
nand UO_1034 (O_1034,N_14781,N_14488);
or UO_1035 (O_1035,N_14503,N_14561);
and UO_1036 (O_1036,N_14433,N_14330);
nand UO_1037 (O_1037,N_14420,N_14603);
or UO_1038 (O_1038,N_14816,N_14615);
nand UO_1039 (O_1039,N_14392,N_14295);
or UO_1040 (O_1040,N_14682,N_14175);
xnor UO_1041 (O_1041,N_14099,N_14582);
or UO_1042 (O_1042,N_14457,N_14206);
and UO_1043 (O_1043,N_14061,N_14607);
and UO_1044 (O_1044,N_14225,N_14294);
nand UO_1045 (O_1045,N_14146,N_14851);
xor UO_1046 (O_1046,N_14999,N_14013);
nor UO_1047 (O_1047,N_14255,N_14006);
or UO_1048 (O_1048,N_14250,N_14549);
nand UO_1049 (O_1049,N_14511,N_14859);
or UO_1050 (O_1050,N_14669,N_14400);
nor UO_1051 (O_1051,N_14260,N_14840);
nand UO_1052 (O_1052,N_14941,N_14874);
xnor UO_1053 (O_1053,N_14435,N_14958);
xor UO_1054 (O_1054,N_14387,N_14177);
nor UO_1055 (O_1055,N_14597,N_14565);
and UO_1056 (O_1056,N_14930,N_14749);
nor UO_1057 (O_1057,N_14325,N_14945);
and UO_1058 (O_1058,N_14073,N_14151);
or UO_1059 (O_1059,N_14974,N_14767);
nor UO_1060 (O_1060,N_14143,N_14369);
or UO_1061 (O_1061,N_14060,N_14203);
or UO_1062 (O_1062,N_14968,N_14194);
nor UO_1063 (O_1063,N_14974,N_14391);
nor UO_1064 (O_1064,N_14094,N_14394);
nor UO_1065 (O_1065,N_14994,N_14203);
nand UO_1066 (O_1066,N_14819,N_14771);
nor UO_1067 (O_1067,N_14238,N_14241);
or UO_1068 (O_1068,N_14793,N_14621);
nor UO_1069 (O_1069,N_14393,N_14267);
xor UO_1070 (O_1070,N_14793,N_14720);
or UO_1071 (O_1071,N_14318,N_14749);
or UO_1072 (O_1072,N_14846,N_14849);
nor UO_1073 (O_1073,N_14506,N_14891);
nor UO_1074 (O_1074,N_14680,N_14031);
or UO_1075 (O_1075,N_14670,N_14313);
and UO_1076 (O_1076,N_14791,N_14629);
nand UO_1077 (O_1077,N_14689,N_14369);
nand UO_1078 (O_1078,N_14423,N_14498);
or UO_1079 (O_1079,N_14924,N_14200);
nand UO_1080 (O_1080,N_14041,N_14696);
nand UO_1081 (O_1081,N_14550,N_14132);
xnor UO_1082 (O_1082,N_14060,N_14813);
nor UO_1083 (O_1083,N_14569,N_14500);
xnor UO_1084 (O_1084,N_14967,N_14704);
and UO_1085 (O_1085,N_14706,N_14678);
and UO_1086 (O_1086,N_14937,N_14045);
xnor UO_1087 (O_1087,N_14225,N_14020);
nor UO_1088 (O_1088,N_14304,N_14171);
xor UO_1089 (O_1089,N_14433,N_14909);
and UO_1090 (O_1090,N_14166,N_14462);
and UO_1091 (O_1091,N_14808,N_14385);
nand UO_1092 (O_1092,N_14902,N_14598);
xor UO_1093 (O_1093,N_14326,N_14435);
nor UO_1094 (O_1094,N_14162,N_14818);
nand UO_1095 (O_1095,N_14023,N_14088);
xnor UO_1096 (O_1096,N_14038,N_14911);
nor UO_1097 (O_1097,N_14157,N_14016);
and UO_1098 (O_1098,N_14511,N_14790);
nand UO_1099 (O_1099,N_14062,N_14178);
xor UO_1100 (O_1100,N_14441,N_14032);
nand UO_1101 (O_1101,N_14481,N_14859);
or UO_1102 (O_1102,N_14549,N_14107);
xnor UO_1103 (O_1103,N_14410,N_14766);
xor UO_1104 (O_1104,N_14478,N_14150);
and UO_1105 (O_1105,N_14989,N_14053);
or UO_1106 (O_1106,N_14690,N_14442);
or UO_1107 (O_1107,N_14632,N_14161);
and UO_1108 (O_1108,N_14455,N_14378);
nand UO_1109 (O_1109,N_14370,N_14389);
xor UO_1110 (O_1110,N_14081,N_14164);
and UO_1111 (O_1111,N_14339,N_14814);
and UO_1112 (O_1112,N_14301,N_14791);
and UO_1113 (O_1113,N_14961,N_14130);
nor UO_1114 (O_1114,N_14931,N_14466);
nor UO_1115 (O_1115,N_14727,N_14219);
nor UO_1116 (O_1116,N_14004,N_14241);
or UO_1117 (O_1117,N_14931,N_14190);
xor UO_1118 (O_1118,N_14924,N_14719);
nand UO_1119 (O_1119,N_14156,N_14248);
or UO_1120 (O_1120,N_14363,N_14290);
or UO_1121 (O_1121,N_14093,N_14564);
nor UO_1122 (O_1122,N_14407,N_14992);
or UO_1123 (O_1123,N_14087,N_14686);
xor UO_1124 (O_1124,N_14052,N_14317);
xnor UO_1125 (O_1125,N_14722,N_14823);
and UO_1126 (O_1126,N_14719,N_14625);
xor UO_1127 (O_1127,N_14286,N_14586);
nand UO_1128 (O_1128,N_14647,N_14951);
nor UO_1129 (O_1129,N_14984,N_14659);
nor UO_1130 (O_1130,N_14812,N_14344);
xor UO_1131 (O_1131,N_14501,N_14452);
nor UO_1132 (O_1132,N_14238,N_14532);
xnor UO_1133 (O_1133,N_14167,N_14475);
nor UO_1134 (O_1134,N_14951,N_14277);
xor UO_1135 (O_1135,N_14905,N_14935);
nor UO_1136 (O_1136,N_14852,N_14638);
and UO_1137 (O_1137,N_14250,N_14767);
or UO_1138 (O_1138,N_14483,N_14213);
or UO_1139 (O_1139,N_14224,N_14479);
nand UO_1140 (O_1140,N_14787,N_14045);
nand UO_1141 (O_1141,N_14560,N_14786);
nor UO_1142 (O_1142,N_14162,N_14667);
xor UO_1143 (O_1143,N_14993,N_14220);
nor UO_1144 (O_1144,N_14703,N_14242);
nand UO_1145 (O_1145,N_14166,N_14387);
nor UO_1146 (O_1146,N_14875,N_14183);
and UO_1147 (O_1147,N_14874,N_14772);
nor UO_1148 (O_1148,N_14361,N_14080);
or UO_1149 (O_1149,N_14661,N_14751);
and UO_1150 (O_1150,N_14123,N_14084);
and UO_1151 (O_1151,N_14877,N_14475);
and UO_1152 (O_1152,N_14324,N_14060);
and UO_1153 (O_1153,N_14804,N_14690);
xor UO_1154 (O_1154,N_14162,N_14842);
and UO_1155 (O_1155,N_14535,N_14548);
or UO_1156 (O_1156,N_14965,N_14872);
nor UO_1157 (O_1157,N_14850,N_14319);
xor UO_1158 (O_1158,N_14260,N_14647);
or UO_1159 (O_1159,N_14940,N_14113);
or UO_1160 (O_1160,N_14058,N_14391);
nand UO_1161 (O_1161,N_14861,N_14758);
xor UO_1162 (O_1162,N_14045,N_14991);
nor UO_1163 (O_1163,N_14523,N_14305);
nand UO_1164 (O_1164,N_14248,N_14973);
and UO_1165 (O_1165,N_14021,N_14335);
or UO_1166 (O_1166,N_14476,N_14542);
nor UO_1167 (O_1167,N_14852,N_14315);
and UO_1168 (O_1168,N_14002,N_14107);
and UO_1169 (O_1169,N_14897,N_14206);
and UO_1170 (O_1170,N_14020,N_14678);
or UO_1171 (O_1171,N_14837,N_14621);
or UO_1172 (O_1172,N_14685,N_14950);
xnor UO_1173 (O_1173,N_14673,N_14364);
xnor UO_1174 (O_1174,N_14606,N_14351);
nor UO_1175 (O_1175,N_14900,N_14131);
or UO_1176 (O_1176,N_14039,N_14851);
and UO_1177 (O_1177,N_14507,N_14362);
nor UO_1178 (O_1178,N_14487,N_14248);
xnor UO_1179 (O_1179,N_14719,N_14801);
and UO_1180 (O_1180,N_14389,N_14417);
xnor UO_1181 (O_1181,N_14577,N_14213);
xnor UO_1182 (O_1182,N_14348,N_14498);
or UO_1183 (O_1183,N_14566,N_14903);
or UO_1184 (O_1184,N_14621,N_14438);
and UO_1185 (O_1185,N_14035,N_14821);
or UO_1186 (O_1186,N_14256,N_14701);
nor UO_1187 (O_1187,N_14877,N_14360);
and UO_1188 (O_1188,N_14769,N_14685);
xor UO_1189 (O_1189,N_14863,N_14182);
and UO_1190 (O_1190,N_14520,N_14494);
nor UO_1191 (O_1191,N_14159,N_14919);
nor UO_1192 (O_1192,N_14095,N_14674);
nor UO_1193 (O_1193,N_14571,N_14789);
xor UO_1194 (O_1194,N_14978,N_14925);
nor UO_1195 (O_1195,N_14339,N_14161);
or UO_1196 (O_1196,N_14894,N_14446);
and UO_1197 (O_1197,N_14753,N_14840);
or UO_1198 (O_1198,N_14014,N_14239);
or UO_1199 (O_1199,N_14638,N_14591);
or UO_1200 (O_1200,N_14796,N_14519);
or UO_1201 (O_1201,N_14153,N_14301);
or UO_1202 (O_1202,N_14678,N_14350);
xnor UO_1203 (O_1203,N_14163,N_14571);
nor UO_1204 (O_1204,N_14711,N_14165);
nor UO_1205 (O_1205,N_14262,N_14356);
and UO_1206 (O_1206,N_14691,N_14942);
nand UO_1207 (O_1207,N_14127,N_14027);
nand UO_1208 (O_1208,N_14658,N_14015);
or UO_1209 (O_1209,N_14921,N_14053);
or UO_1210 (O_1210,N_14271,N_14365);
nor UO_1211 (O_1211,N_14457,N_14518);
nand UO_1212 (O_1212,N_14364,N_14572);
nand UO_1213 (O_1213,N_14107,N_14273);
and UO_1214 (O_1214,N_14668,N_14879);
nand UO_1215 (O_1215,N_14873,N_14491);
or UO_1216 (O_1216,N_14852,N_14241);
and UO_1217 (O_1217,N_14604,N_14676);
xor UO_1218 (O_1218,N_14639,N_14499);
nand UO_1219 (O_1219,N_14641,N_14616);
xor UO_1220 (O_1220,N_14782,N_14425);
xor UO_1221 (O_1221,N_14144,N_14272);
nand UO_1222 (O_1222,N_14173,N_14154);
nor UO_1223 (O_1223,N_14252,N_14654);
nand UO_1224 (O_1224,N_14396,N_14430);
and UO_1225 (O_1225,N_14204,N_14306);
nor UO_1226 (O_1226,N_14461,N_14545);
xor UO_1227 (O_1227,N_14716,N_14049);
xor UO_1228 (O_1228,N_14257,N_14711);
nand UO_1229 (O_1229,N_14452,N_14915);
and UO_1230 (O_1230,N_14343,N_14819);
and UO_1231 (O_1231,N_14911,N_14226);
nand UO_1232 (O_1232,N_14199,N_14455);
and UO_1233 (O_1233,N_14644,N_14812);
xnor UO_1234 (O_1234,N_14652,N_14481);
xnor UO_1235 (O_1235,N_14656,N_14613);
nor UO_1236 (O_1236,N_14686,N_14183);
nor UO_1237 (O_1237,N_14771,N_14517);
nand UO_1238 (O_1238,N_14996,N_14457);
or UO_1239 (O_1239,N_14999,N_14816);
nor UO_1240 (O_1240,N_14956,N_14953);
or UO_1241 (O_1241,N_14278,N_14495);
or UO_1242 (O_1242,N_14510,N_14493);
or UO_1243 (O_1243,N_14289,N_14939);
nand UO_1244 (O_1244,N_14130,N_14618);
nand UO_1245 (O_1245,N_14066,N_14497);
xnor UO_1246 (O_1246,N_14979,N_14813);
nor UO_1247 (O_1247,N_14550,N_14668);
and UO_1248 (O_1248,N_14428,N_14469);
xnor UO_1249 (O_1249,N_14148,N_14816);
xor UO_1250 (O_1250,N_14624,N_14933);
and UO_1251 (O_1251,N_14981,N_14446);
xor UO_1252 (O_1252,N_14730,N_14853);
or UO_1253 (O_1253,N_14027,N_14909);
and UO_1254 (O_1254,N_14170,N_14725);
xor UO_1255 (O_1255,N_14140,N_14697);
nor UO_1256 (O_1256,N_14099,N_14132);
nor UO_1257 (O_1257,N_14413,N_14244);
and UO_1258 (O_1258,N_14658,N_14363);
nor UO_1259 (O_1259,N_14075,N_14553);
xor UO_1260 (O_1260,N_14175,N_14655);
and UO_1261 (O_1261,N_14669,N_14986);
and UO_1262 (O_1262,N_14718,N_14324);
or UO_1263 (O_1263,N_14857,N_14084);
xnor UO_1264 (O_1264,N_14361,N_14231);
nand UO_1265 (O_1265,N_14484,N_14737);
and UO_1266 (O_1266,N_14973,N_14836);
nor UO_1267 (O_1267,N_14024,N_14370);
and UO_1268 (O_1268,N_14119,N_14762);
or UO_1269 (O_1269,N_14862,N_14059);
nand UO_1270 (O_1270,N_14303,N_14122);
xor UO_1271 (O_1271,N_14539,N_14484);
nor UO_1272 (O_1272,N_14282,N_14227);
nand UO_1273 (O_1273,N_14684,N_14542);
xnor UO_1274 (O_1274,N_14299,N_14055);
xnor UO_1275 (O_1275,N_14904,N_14795);
nand UO_1276 (O_1276,N_14607,N_14063);
nand UO_1277 (O_1277,N_14408,N_14659);
xnor UO_1278 (O_1278,N_14088,N_14419);
nor UO_1279 (O_1279,N_14358,N_14151);
nand UO_1280 (O_1280,N_14434,N_14310);
xnor UO_1281 (O_1281,N_14471,N_14319);
and UO_1282 (O_1282,N_14178,N_14988);
and UO_1283 (O_1283,N_14969,N_14653);
or UO_1284 (O_1284,N_14538,N_14181);
or UO_1285 (O_1285,N_14602,N_14910);
and UO_1286 (O_1286,N_14020,N_14202);
xnor UO_1287 (O_1287,N_14149,N_14742);
and UO_1288 (O_1288,N_14255,N_14187);
and UO_1289 (O_1289,N_14634,N_14942);
and UO_1290 (O_1290,N_14073,N_14721);
nor UO_1291 (O_1291,N_14907,N_14780);
and UO_1292 (O_1292,N_14553,N_14262);
xor UO_1293 (O_1293,N_14982,N_14977);
xor UO_1294 (O_1294,N_14738,N_14983);
nor UO_1295 (O_1295,N_14604,N_14394);
nor UO_1296 (O_1296,N_14868,N_14685);
nand UO_1297 (O_1297,N_14454,N_14062);
xor UO_1298 (O_1298,N_14815,N_14805);
nand UO_1299 (O_1299,N_14643,N_14963);
or UO_1300 (O_1300,N_14741,N_14704);
or UO_1301 (O_1301,N_14476,N_14381);
nand UO_1302 (O_1302,N_14926,N_14324);
nand UO_1303 (O_1303,N_14433,N_14384);
or UO_1304 (O_1304,N_14270,N_14631);
nor UO_1305 (O_1305,N_14746,N_14832);
and UO_1306 (O_1306,N_14754,N_14059);
or UO_1307 (O_1307,N_14778,N_14345);
and UO_1308 (O_1308,N_14942,N_14965);
nor UO_1309 (O_1309,N_14889,N_14370);
and UO_1310 (O_1310,N_14747,N_14392);
xnor UO_1311 (O_1311,N_14655,N_14276);
and UO_1312 (O_1312,N_14766,N_14348);
xor UO_1313 (O_1313,N_14787,N_14641);
and UO_1314 (O_1314,N_14448,N_14414);
nor UO_1315 (O_1315,N_14040,N_14258);
nor UO_1316 (O_1316,N_14120,N_14495);
or UO_1317 (O_1317,N_14334,N_14678);
and UO_1318 (O_1318,N_14636,N_14748);
xnor UO_1319 (O_1319,N_14709,N_14845);
xor UO_1320 (O_1320,N_14654,N_14509);
xnor UO_1321 (O_1321,N_14763,N_14317);
and UO_1322 (O_1322,N_14339,N_14088);
xor UO_1323 (O_1323,N_14574,N_14255);
and UO_1324 (O_1324,N_14665,N_14699);
or UO_1325 (O_1325,N_14835,N_14869);
or UO_1326 (O_1326,N_14058,N_14118);
xnor UO_1327 (O_1327,N_14946,N_14655);
nand UO_1328 (O_1328,N_14356,N_14962);
xnor UO_1329 (O_1329,N_14874,N_14394);
or UO_1330 (O_1330,N_14483,N_14050);
xor UO_1331 (O_1331,N_14974,N_14017);
xnor UO_1332 (O_1332,N_14585,N_14179);
or UO_1333 (O_1333,N_14336,N_14177);
nor UO_1334 (O_1334,N_14072,N_14194);
xor UO_1335 (O_1335,N_14566,N_14410);
xnor UO_1336 (O_1336,N_14961,N_14160);
xor UO_1337 (O_1337,N_14656,N_14849);
nand UO_1338 (O_1338,N_14147,N_14999);
nand UO_1339 (O_1339,N_14625,N_14924);
nor UO_1340 (O_1340,N_14386,N_14011);
or UO_1341 (O_1341,N_14863,N_14948);
xnor UO_1342 (O_1342,N_14520,N_14193);
nor UO_1343 (O_1343,N_14295,N_14762);
xor UO_1344 (O_1344,N_14385,N_14447);
xor UO_1345 (O_1345,N_14746,N_14353);
and UO_1346 (O_1346,N_14822,N_14732);
nor UO_1347 (O_1347,N_14457,N_14202);
xnor UO_1348 (O_1348,N_14300,N_14405);
nand UO_1349 (O_1349,N_14933,N_14163);
nor UO_1350 (O_1350,N_14475,N_14600);
nand UO_1351 (O_1351,N_14841,N_14407);
or UO_1352 (O_1352,N_14662,N_14738);
and UO_1353 (O_1353,N_14623,N_14729);
and UO_1354 (O_1354,N_14405,N_14072);
and UO_1355 (O_1355,N_14877,N_14411);
nor UO_1356 (O_1356,N_14795,N_14238);
xor UO_1357 (O_1357,N_14757,N_14747);
or UO_1358 (O_1358,N_14959,N_14238);
and UO_1359 (O_1359,N_14966,N_14181);
and UO_1360 (O_1360,N_14541,N_14267);
or UO_1361 (O_1361,N_14320,N_14259);
nor UO_1362 (O_1362,N_14990,N_14767);
and UO_1363 (O_1363,N_14960,N_14766);
and UO_1364 (O_1364,N_14324,N_14000);
or UO_1365 (O_1365,N_14423,N_14012);
xnor UO_1366 (O_1366,N_14906,N_14605);
and UO_1367 (O_1367,N_14645,N_14760);
nor UO_1368 (O_1368,N_14434,N_14257);
nor UO_1369 (O_1369,N_14844,N_14950);
xnor UO_1370 (O_1370,N_14255,N_14694);
nand UO_1371 (O_1371,N_14479,N_14370);
nand UO_1372 (O_1372,N_14166,N_14291);
xnor UO_1373 (O_1373,N_14752,N_14753);
nor UO_1374 (O_1374,N_14179,N_14651);
xnor UO_1375 (O_1375,N_14939,N_14507);
nand UO_1376 (O_1376,N_14972,N_14045);
nor UO_1377 (O_1377,N_14132,N_14332);
or UO_1378 (O_1378,N_14358,N_14061);
xnor UO_1379 (O_1379,N_14112,N_14988);
or UO_1380 (O_1380,N_14461,N_14669);
and UO_1381 (O_1381,N_14707,N_14911);
xnor UO_1382 (O_1382,N_14144,N_14295);
or UO_1383 (O_1383,N_14023,N_14961);
nand UO_1384 (O_1384,N_14607,N_14552);
and UO_1385 (O_1385,N_14861,N_14458);
and UO_1386 (O_1386,N_14218,N_14383);
and UO_1387 (O_1387,N_14897,N_14158);
and UO_1388 (O_1388,N_14604,N_14476);
nor UO_1389 (O_1389,N_14385,N_14942);
xnor UO_1390 (O_1390,N_14505,N_14817);
nand UO_1391 (O_1391,N_14964,N_14490);
nand UO_1392 (O_1392,N_14500,N_14606);
xor UO_1393 (O_1393,N_14949,N_14589);
or UO_1394 (O_1394,N_14338,N_14279);
nor UO_1395 (O_1395,N_14297,N_14374);
nor UO_1396 (O_1396,N_14945,N_14998);
xor UO_1397 (O_1397,N_14922,N_14936);
or UO_1398 (O_1398,N_14624,N_14287);
or UO_1399 (O_1399,N_14526,N_14686);
nand UO_1400 (O_1400,N_14512,N_14837);
xnor UO_1401 (O_1401,N_14987,N_14135);
xor UO_1402 (O_1402,N_14550,N_14883);
xor UO_1403 (O_1403,N_14157,N_14591);
nand UO_1404 (O_1404,N_14477,N_14534);
xnor UO_1405 (O_1405,N_14495,N_14151);
and UO_1406 (O_1406,N_14969,N_14878);
nand UO_1407 (O_1407,N_14748,N_14189);
xor UO_1408 (O_1408,N_14745,N_14335);
nand UO_1409 (O_1409,N_14220,N_14840);
nand UO_1410 (O_1410,N_14041,N_14934);
xnor UO_1411 (O_1411,N_14915,N_14234);
or UO_1412 (O_1412,N_14448,N_14249);
nand UO_1413 (O_1413,N_14573,N_14511);
xnor UO_1414 (O_1414,N_14049,N_14394);
xor UO_1415 (O_1415,N_14727,N_14169);
and UO_1416 (O_1416,N_14370,N_14707);
xor UO_1417 (O_1417,N_14473,N_14727);
nand UO_1418 (O_1418,N_14372,N_14577);
nor UO_1419 (O_1419,N_14241,N_14054);
and UO_1420 (O_1420,N_14395,N_14486);
nor UO_1421 (O_1421,N_14851,N_14860);
nor UO_1422 (O_1422,N_14188,N_14850);
nand UO_1423 (O_1423,N_14313,N_14650);
xor UO_1424 (O_1424,N_14110,N_14788);
nor UO_1425 (O_1425,N_14949,N_14756);
nor UO_1426 (O_1426,N_14877,N_14586);
xnor UO_1427 (O_1427,N_14847,N_14609);
xnor UO_1428 (O_1428,N_14402,N_14548);
xor UO_1429 (O_1429,N_14358,N_14117);
or UO_1430 (O_1430,N_14981,N_14039);
and UO_1431 (O_1431,N_14517,N_14329);
nand UO_1432 (O_1432,N_14951,N_14518);
and UO_1433 (O_1433,N_14339,N_14326);
nand UO_1434 (O_1434,N_14074,N_14485);
nor UO_1435 (O_1435,N_14546,N_14682);
nand UO_1436 (O_1436,N_14821,N_14676);
nand UO_1437 (O_1437,N_14217,N_14547);
nand UO_1438 (O_1438,N_14656,N_14674);
and UO_1439 (O_1439,N_14657,N_14529);
and UO_1440 (O_1440,N_14158,N_14076);
nand UO_1441 (O_1441,N_14940,N_14364);
nand UO_1442 (O_1442,N_14953,N_14929);
nor UO_1443 (O_1443,N_14799,N_14084);
or UO_1444 (O_1444,N_14454,N_14972);
or UO_1445 (O_1445,N_14701,N_14387);
nand UO_1446 (O_1446,N_14935,N_14404);
nor UO_1447 (O_1447,N_14031,N_14354);
or UO_1448 (O_1448,N_14383,N_14148);
nor UO_1449 (O_1449,N_14230,N_14400);
nand UO_1450 (O_1450,N_14333,N_14736);
nor UO_1451 (O_1451,N_14361,N_14690);
or UO_1452 (O_1452,N_14741,N_14808);
or UO_1453 (O_1453,N_14400,N_14273);
and UO_1454 (O_1454,N_14441,N_14157);
nand UO_1455 (O_1455,N_14688,N_14404);
and UO_1456 (O_1456,N_14775,N_14313);
nor UO_1457 (O_1457,N_14562,N_14820);
or UO_1458 (O_1458,N_14696,N_14595);
nand UO_1459 (O_1459,N_14116,N_14640);
nor UO_1460 (O_1460,N_14899,N_14951);
xor UO_1461 (O_1461,N_14139,N_14161);
nand UO_1462 (O_1462,N_14422,N_14569);
xor UO_1463 (O_1463,N_14078,N_14088);
xnor UO_1464 (O_1464,N_14830,N_14044);
nor UO_1465 (O_1465,N_14406,N_14798);
xor UO_1466 (O_1466,N_14539,N_14865);
xnor UO_1467 (O_1467,N_14597,N_14241);
xnor UO_1468 (O_1468,N_14995,N_14298);
nor UO_1469 (O_1469,N_14144,N_14816);
and UO_1470 (O_1470,N_14350,N_14230);
and UO_1471 (O_1471,N_14715,N_14691);
and UO_1472 (O_1472,N_14928,N_14840);
and UO_1473 (O_1473,N_14794,N_14392);
or UO_1474 (O_1474,N_14427,N_14665);
xor UO_1475 (O_1475,N_14839,N_14658);
nand UO_1476 (O_1476,N_14786,N_14088);
or UO_1477 (O_1477,N_14694,N_14195);
xnor UO_1478 (O_1478,N_14832,N_14555);
or UO_1479 (O_1479,N_14347,N_14992);
or UO_1480 (O_1480,N_14205,N_14276);
nand UO_1481 (O_1481,N_14169,N_14490);
and UO_1482 (O_1482,N_14717,N_14762);
nor UO_1483 (O_1483,N_14923,N_14434);
or UO_1484 (O_1484,N_14377,N_14363);
nand UO_1485 (O_1485,N_14818,N_14110);
nor UO_1486 (O_1486,N_14517,N_14845);
nor UO_1487 (O_1487,N_14245,N_14092);
and UO_1488 (O_1488,N_14644,N_14660);
or UO_1489 (O_1489,N_14423,N_14902);
and UO_1490 (O_1490,N_14706,N_14454);
or UO_1491 (O_1491,N_14900,N_14306);
and UO_1492 (O_1492,N_14567,N_14850);
nand UO_1493 (O_1493,N_14543,N_14814);
nor UO_1494 (O_1494,N_14271,N_14774);
and UO_1495 (O_1495,N_14755,N_14233);
nand UO_1496 (O_1496,N_14378,N_14627);
xnor UO_1497 (O_1497,N_14866,N_14724);
xnor UO_1498 (O_1498,N_14290,N_14643);
and UO_1499 (O_1499,N_14004,N_14437);
or UO_1500 (O_1500,N_14519,N_14209);
nand UO_1501 (O_1501,N_14379,N_14523);
xor UO_1502 (O_1502,N_14202,N_14989);
xnor UO_1503 (O_1503,N_14188,N_14052);
nand UO_1504 (O_1504,N_14382,N_14127);
or UO_1505 (O_1505,N_14770,N_14283);
nand UO_1506 (O_1506,N_14585,N_14110);
or UO_1507 (O_1507,N_14632,N_14800);
nand UO_1508 (O_1508,N_14509,N_14773);
nand UO_1509 (O_1509,N_14678,N_14028);
xnor UO_1510 (O_1510,N_14659,N_14594);
nor UO_1511 (O_1511,N_14632,N_14287);
nand UO_1512 (O_1512,N_14873,N_14272);
nand UO_1513 (O_1513,N_14553,N_14589);
nor UO_1514 (O_1514,N_14993,N_14667);
or UO_1515 (O_1515,N_14447,N_14705);
nor UO_1516 (O_1516,N_14009,N_14411);
nor UO_1517 (O_1517,N_14037,N_14573);
or UO_1518 (O_1518,N_14119,N_14198);
nor UO_1519 (O_1519,N_14714,N_14069);
or UO_1520 (O_1520,N_14117,N_14928);
nor UO_1521 (O_1521,N_14734,N_14752);
nand UO_1522 (O_1522,N_14977,N_14163);
and UO_1523 (O_1523,N_14231,N_14932);
xor UO_1524 (O_1524,N_14584,N_14109);
or UO_1525 (O_1525,N_14484,N_14788);
and UO_1526 (O_1526,N_14761,N_14559);
xor UO_1527 (O_1527,N_14981,N_14622);
nor UO_1528 (O_1528,N_14602,N_14202);
nand UO_1529 (O_1529,N_14484,N_14194);
xor UO_1530 (O_1530,N_14134,N_14011);
and UO_1531 (O_1531,N_14602,N_14880);
nor UO_1532 (O_1532,N_14919,N_14509);
or UO_1533 (O_1533,N_14044,N_14862);
or UO_1534 (O_1534,N_14037,N_14281);
and UO_1535 (O_1535,N_14517,N_14813);
nor UO_1536 (O_1536,N_14939,N_14026);
or UO_1537 (O_1537,N_14546,N_14936);
nand UO_1538 (O_1538,N_14183,N_14997);
xnor UO_1539 (O_1539,N_14476,N_14680);
and UO_1540 (O_1540,N_14538,N_14696);
nor UO_1541 (O_1541,N_14897,N_14301);
nor UO_1542 (O_1542,N_14320,N_14210);
nand UO_1543 (O_1543,N_14997,N_14041);
nor UO_1544 (O_1544,N_14853,N_14092);
or UO_1545 (O_1545,N_14879,N_14349);
nand UO_1546 (O_1546,N_14127,N_14471);
nand UO_1547 (O_1547,N_14499,N_14865);
xor UO_1548 (O_1548,N_14703,N_14597);
and UO_1549 (O_1549,N_14532,N_14089);
xor UO_1550 (O_1550,N_14504,N_14399);
and UO_1551 (O_1551,N_14150,N_14569);
xnor UO_1552 (O_1552,N_14219,N_14754);
nand UO_1553 (O_1553,N_14376,N_14832);
and UO_1554 (O_1554,N_14903,N_14646);
nor UO_1555 (O_1555,N_14221,N_14717);
nand UO_1556 (O_1556,N_14179,N_14120);
or UO_1557 (O_1557,N_14424,N_14494);
nand UO_1558 (O_1558,N_14993,N_14604);
nor UO_1559 (O_1559,N_14236,N_14652);
or UO_1560 (O_1560,N_14196,N_14056);
and UO_1561 (O_1561,N_14631,N_14356);
xor UO_1562 (O_1562,N_14882,N_14787);
xor UO_1563 (O_1563,N_14552,N_14002);
and UO_1564 (O_1564,N_14865,N_14834);
or UO_1565 (O_1565,N_14061,N_14093);
or UO_1566 (O_1566,N_14970,N_14724);
xnor UO_1567 (O_1567,N_14080,N_14593);
or UO_1568 (O_1568,N_14980,N_14697);
xnor UO_1569 (O_1569,N_14537,N_14912);
nor UO_1570 (O_1570,N_14240,N_14313);
nor UO_1571 (O_1571,N_14502,N_14593);
nand UO_1572 (O_1572,N_14115,N_14273);
and UO_1573 (O_1573,N_14195,N_14767);
nor UO_1574 (O_1574,N_14080,N_14708);
and UO_1575 (O_1575,N_14265,N_14652);
nor UO_1576 (O_1576,N_14669,N_14835);
or UO_1577 (O_1577,N_14666,N_14573);
nor UO_1578 (O_1578,N_14749,N_14585);
and UO_1579 (O_1579,N_14622,N_14760);
or UO_1580 (O_1580,N_14785,N_14245);
nand UO_1581 (O_1581,N_14326,N_14597);
nand UO_1582 (O_1582,N_14582,N_14883);
nand UO_1583 (O_1583,N_14397,N_14004);
nand UO_1584 (O_1584,N_14153,N_14697);
nand UO_1585 (O_1585,N_14877,N_14659);
nand UO_1586 (O_1586,N_14943,N_14227);
nand UO_1587 (O_1587,N_14601,N_14501);
and UO_1588 (O_1588,N_14212,N_14886);
nor UO_1589 (O_1589,N_14688,N_14871);
nor UO_1590 (O_1590,N_14815,N_14004);
xnor UO_1591 (O_1591,N_14264,N_14216);
nand UO_1592 (O_1592,N_14905,N_14878);
nor UO_1593 (O_1593,N_14787,N_14770);
nand UO_1594 (O_1594,N_14055,N_14593);
xor UO_1595 (O_1595,N_14494,N_14993);
nor UO_1596 (O_1596,N_14084,N_14686);
or UO_1597 (O_1597,N_14332,N_14466);
nor UO_1598 (O_1598,N_14616,N_14166);
xnor UO_1599 (O_1599,N_14390,N_14339);
or UO_1600 (O_1600,N_14454,N_14043);
or UO_1601 (O_1601,N_14854,N_14425);
nand UO_1602 (O_1602,N_14685,N_14915);
or UO_1603 (O_1603,N_14865,N_14615);
or UO_1604 (O_1604,N_14460,N_14537);
nand UO_1605 (O_1605,N_14668,N_14623);
or UO_1606 (O_1606,N_14371,N_14902);
or UO_1607 (O_1607,N_14912,N_14210);
xor UO_1608 (O_1608,N_14358,N_14759);
nand UO_1609 (O_1609,N_14557,N_14195);
nor UO_1610 (O_1610,N_14264,N_14755);
nor UO_1611 (O_1611,N_14593,N_14855);
or UO_1612 (O_1612,N_14870,N_14391);
nand UO_1613 (O_1613,N_14700,N_14054);
and UO_1614 (O_1614,N_14437,N_14914);
nand UO_1615 (O_1615,N_14644,N_14816);
and UO_1616 (O_1616,N_14615,N_14167);
nand UO_1617 (O_1617,N_14575,N_14517);
or UO_1618 (O_1618,N_14129,N_14984);
nor UO_1619 (O_1619,N_14681,N_14769);
xnor UO_1620 (O_1620,N_14717,N_14198);
or UO_1621 (O_1621,N_14823,N_14581);
xor UO_1622 (O_1622,N_14883,N_14413);
nand UO_1623 (O_1623,N_14833,N_14587);
nand UO_1624 (O_1624,N_14304,N_14461);
xor UO_1625 (O_1625,N_14796,N_14680);
or UO_1626 (O_1626,N_14844,N_14732);
or UO_1627 (O_1627,N_14898,N_14924);
nor UO_1628 (O_1628,N_14850,N_14307);
nor UO_1629 (O_1629,N_14661,N_14654);
nor UO_1630 (O_1630,N_14047,N_14064);
xor UO_1631 (O_1631,N_14115,N_14942);
nand UO_1632 (O_1632,N_14733,N_14813);
and UO_1633 (O_1633,N_14395,N_14035);
xnor UO_1634 (O_1634,N_14981,N_14523);
nand UO_1635 (O_1635,N_14011,N_14423);
and UO_1636 (O_1636,N_14925,N_14307);
nand UO_1637 (O_1637,N_14682,N_14247);
nand UO_1638 (O_1638,N_14417,N_14643);
or UO_1639 (O_1639,N_14691,N_14103);
nand UO_1640 (O_1640,N_14039,N_14305);
nand UO_1641 (O_1641,N_14319,N_14734);
and UO_1642 (O_1642,N_14882,N_14497);
and UO_1643 (O_1643,N_14137,N_14232);
and UO_1644 (O_1644,N_14542,N_14122);
nand UO_1645 (O_1645,N_14623,N_14971);
nor UO_1646 (O_1646,N_14788,N_14835);
nor UO_1647 (O_1647,N_14622,N_14909);
xor UO_1648 (O_1648,N_14785,N_14276);
xnor UO_1649 (O_1649,N_14614,N_14610);
nand UO_1650 (O_1650,N_14143,N_14714);
or UO_1651 (O_1651,N_14051,N_14174);
or UO_1652 (O_1652,N_14854,N_14752);
or UO_1653 (O_1653,N_14640,N_14982);
or UO_1654 (O_1654,N_14536,N_14805);
and UO_1655 (O_1655,N_14616,N_14170);
nor UO_1656 (O_1656,N_14007,N_14308);
nand UO_1657 (O_1657,N_14207,N_14216);
nor UO_1658 (O_1658,N_14261,N_14563);
nand UO_1659 (O_1659,N_14540,N_14447);
and UO_1660 (O_1660,N_14348,N_14723);
xnor UO_1661 (O_1661,N_14142,N_14093);
nor UO_1662 (O_1662,N_14406,N_14493);
nor UO_1663 (O_1663,N_14965,N_14519);
nor UO_1664 (O_1664,N_14807,N_14747);
nor UO_1665 (O_1665,N_14329,N_14166);
or UO_1666 (O_1666,N_14979,N_14239);
nand UO_1667 (O_1667,N_14555,N_14474);
or UO_1668 (O_1668,N_14835,N_14411);
or UO_1669 (O_1669,N_14670,N_14299);
or UO_1670 (O_1670,N_14185,N_14902);
and UO_1671 (O_1671,N_14417,N_14275);
or UO_1672 (O_1672,N_14820,N_14864);
nand UO_1673 (O_1673,N_14928,N_14650);
or UO_1674 (O_1674,N_14409,N_14581);
nor UO_1675 (O_1675,N_14189,N_14446);
or UO_1676 (O_1676,N_14671,N_14087);
nor UO_1677 (O_1677,N_14024,N_14299);
or UO_1678 (O_1678,N_14550,N_14313);
nor UO_1679 (O_1679,N_14726,N_14391);
and UO_1680 (O_1680,N_14139,N_14768);
nor UO_1681 (O_1681,N_14398,N_14687);
nand UO_1682 (O_1682,N_14510,N_14087);
nor UO_1683 (O_1683,N_14219,N_14645);
nor UO_1684 (O_1684,N_14626,N_14573);
nor UO_1685 (O_1685,N_14273,N_14408);
nor UO_1686 (O_1686,N_14710,N_14781);
nor UO_1687 (O_1687,N_14377,N_14915);
nand UO_1688 (O_1688,N_14921,N_14725);
xnor UO_1689 (O_1689,N_14982,N_14399);
nand UO_1690 (O_1690,N_14484,N_14927);
and UO_1691 (O_1691,N_14231,N_14404);
xor UO_1692 (O_1692,N_14922,N_14270);
nor UO_1693 (O_1693,N_14921,N_14782);
or UO_1694 (O_1694,N_14877,N_14613);
xor UO_1695 (O_1695,N_14261,N_14840);
nor UO_1696 (O_1696,N_14568,N_14619);
or UO_1697 (O_1697,N_14928,N_14212);
nand UO_1698 (O_1698,N_14507,N_14948);
nand UO_1699 (O_1699,N_14826,N_14396);
nor UO_1700 (O_1700,N_14367,N_14809);
and UO_1701 (O_1701,N_14404,N_14550);
nand UO_1702 (O_1702,N_14867,N_14248);
and UO_1703 (O_1703,N_14724,N_14067);
or UO_1704 (O_1704,N_14908,N_14035);
and UO_1705 (O_1705,N_14680,N_14910);
and UO_1706 (O_1706,N_14889,N_14423);
xnor UO_1707 (O_1707,N_14348,N_14460);
or UO_1708 (O_1708,N_14002,N_14184);
xnor UO_1709 (O_1709,N_14704,N_14572);
xor UO_1710 (O_1710,N_14220,N_14837);
nor UO_1711 (O_1711,N_14965,N_14185);
or UO_1712 (O_1712,N_14431,N_14706);
nand UO_1713 (O_1713,N_14196,N_14972);
nand UO_1714 (O_1714,N_14803,N_14977);
nor UO_1715 (O_1715,N_14951,N_14964);
nand UO_1716 (O_1716,N_14844,N_14771);
xnor UO_1717 (O_1717,N_14158,N_14979);
xor UO_1718 (O_1718,N_14906,N_14260);
or UO_1719 (O_1719,N_14392,N_14525);
xnor UO_1720 (O_1720,N_14750,N_14445);
and UO_1721 (O_1721,N_14453,N_14332);
nor UO_1722 (O_1722,N_14099,N_14268);
xor UO_1723 (O_1723,N_14640,N_14267);
or UO_1724 (O_1724,N_14701,N_14928);
nand UO_1725 (O_1725,N_14601,N_14872);
and UO_1726 (O_1726,N_14839,N_14031);
xor UO_1727 (O_1727,N_14234,N_14874);
nor UO_1728 (O_1728,N_14071,N_14081);
nor UO_1729 (O_1729,N_14961,N_14086);
xor UO_1730 (O_1730,N_14032,N_14779);
and UO_1731 (O_1731,N_14789,N_14628);
or UO_1732 (O_1732,N_14338,N_14100);
or UO_1733 (O_1733,N_14735,N_14289);
xor UO_1734 (O_1734,N_14719,N_14186);
or UO_1735 (O_1735,N_14315,N_14567);
nor UO_1736 (O_1736,N_14454,N_14340);
or UO_1737 (O_1737,N_14026,N_14263);
nor UO_1738 (O_1738,N_14747,N_14494);
nand UO_1739 (O_1739,N_14359,N_14894);
nor UO_1740 (O_1740,N_14354,N_14116);
or UO_1741 (O_1741,N_14278,N_14071);
xor UO_1742 (O_1742,N_14480,N_14748);
or UO_1743 (O_1743,N_14131,N_14762);
or UO_1744 (O_1744,N_14474,N_14106);
or UO_1745 (O_1745,N_14231,N_14828);
nor UO_1746 (O_1746,N_14517,N_14105);
xor UO_1747 (O_1747,N_14111,N_14675);
xnor UO_1748 (O_1748,N_14514,N_14895);
or UO_1749 (O_1749,N_14126,N_14243);
or UO_1750 (O_1750,N_14365,N_14611);
nor UO_1751 (O_1751,N_14087,N_14733);
xor UO_1752 (O_1752,N_14180,N_14060);
nand UO_1753 (O_1753,N_14094,N_14578);
xnor UO_1754 (O_1754,N_14437,N_14030);
nand UO_1755 (O_1755,N_14344,N_14851);
nor UO_1756 (O_1756,N_14710,N_14828);
or UO_1757 (O_1757,N_14518,N_14273);
nand UO_1758 (O_1758,N_14545,N_14833);
or UO_1759 (O_1759,N_14240,N_14756);
or UO_1760 (O_1760,N_14862,N_14505);
nand UO_1761 (O_1761,N_14592,N_14559);
nor UO_1762 (O_1762,N_14571,N_14225);
nand UO_1763 (O_1763,N_14689,N_14357);
and UO_1764 (O_1764,N_14616,N_14053);
and UO_1765 (O_1765,N_14091,N_14422);
nand UO_1766 (O_1766,N_14567,N_14652);
nand UO_1767 (O_1767,N_14294,N_14759);
nand UO_1768 (O_1768,N_14154,N_14756);
or UO_1769 (O_1769,N_14133,N_14425);
nor UO_1770 (O_1770,N_14716,N_14607);
and UO_1771 (O_1771,N_14026,N_14592);
nand UO_1772 (O_1772,N_14636,N_14498);
nor UO_1773 (O_1773,N_14248,N_14067);
and UO_1774 (O_1774,N_14085,N_14864);
nand UO_1775 (O_1775,N_14723,N_14038);
or UO_1776 (O_1776,N_14791,N_14630);
and UO_1777 (O_1777,N_14408,N_14773);
nor UO_1778 (O_1778,N_14965,N_14462);
nand UO_1779 (O_1779,N_14699,N_14238);
or UO_1780 (O_1780,N_14292,N_14986);
nor UO_1781 (O_1781,N_14444,N_14068);
nand UO_1782 (O_1782,N_14167,N_14084);
and UO_1783 (O_1783,N_14400,N_14820);
nor UO_1784 (O_1784,N_14559,N_14879);
or UO_1785 (O_1785,N_14460,N_14946);
xnor UO_1786 (O_1786,N_14574,N_14917);
or UO_1787 (O_1787,N_14560,N_14581);
nor UO_1788 (O_1788,N_14910,N_14811);
xor UO_1789 (O_1789,N_14233,N_14052);
and UO_1790 (O_1790,N_14368,N_14479);
xnor UO_1791 (O_1791,N_14318,N_14585);
or UO_1792 (O_1792,N_14028,N_14236);
or UO_1793 (O_1793,N_14254,N_14226);
nor UO_1794 (O_1794,N_14934,N_14325);
nor UO_1795 (O_1795,N_14461,N_14487);
and UO_1796 (O_1796,N_14390,N_14538);
or UO_1797 (O_1797,N_14585,N_14162);
or UO_1798 (O_1798,N_14053,N_14471);
or UO_1799 (O_1799,N_14433,N_14741);
xor UO_1800 (O_1800,N_14866,N_14705);
xnor UO_1801 (O_1801,N_14314,N_14848);
nor UO_1802 (O_1802,N_14841,N_14825);
or UO_1803 (O_1803,N_14717,N_14769);
and UO_1804 (O_1804,N_14820,N_14285);
nor UO_1805 (O_1805,N_14520,N_14518);
nand UO_1806 (O_1806,N_14208,N_14850);
or UO_1807 (O_1807,N_14408,N_14709);
or UO_1808 (O_1808,N_14532,N_14805);
xor UO_1809 (O_1809,N_14109,N_14291);
xor UO_1810 (O_1810,N_14884,N_14649);
xor UO_1811 (O_1811,N_14167,N_14270);
xor UO_1812 (O_1812,N_14375,N_14057);
and UO_1813 (O_1813,N_14323,N_14654);
and UO_1814 (O_1814,N_14701,N_14685);
and UO_1815 (O_1815,N_14980,N_14196);
xnor UO_1816 (O_1816,N_14877,N_14804);
nand UO_1817 (O_1817,N_14662,N_14068);
nand UO_1818 (O_1818,N_14362,N_14696);
and UO_1819 (O_1819,N_14335,N_14118);
nor UO_1820 (O_1820,N_14791,N_14725);
or UO_1821 (O_1821,N_14255,N_14599);
xnor UO_1822 (O_1822,N_14642,N_14832);
nand UO_1823 (O_1823,N_14849,N_14142);
and UO_1824 (O_1824,N_14748,N_14209);
or UO_1825 (O_1825,N_14404,N_14325);
or UO_1826 (O_1826,N_14393,N_14050);
xor UO_1827 (O_1827,N_14701,N_14342);
nand UO_1828 (O_1828,N_14901,N_14599);
xnor UO_1829 (O_1829,N_14947,N_14324);
nand UO_1830 (O_1830,N_14858,N_14469);
and UO_1831 (O_1831,N_14900,N_14901);
nand UO_1832 (O_1832,N_14133,N_14867);
xor UO_1833 (O_1833,N_14758,N_14403);
or UO_1834 (O_1834,N_14414,N_14343);
or UO_1835 (O_1835,N_14909,N_14679);
xnor UO_1836 (O_1836,N_14696,N_14495);
and UO_1837 (O_1837,N_14064,N_14298);
and UO_1838 (O_1838,N_14417,N_14266);
xnor UO_1839 (O_1839,N_14501,N_14489);
nand UO_1840 (O_1840,N_14140,N_14258);
nand UO_1841 (O_1841,N_14522,N_14260);
xor UO_1842 (O_1842,N_14908,N_14045);
xor UO_1843 (O_1843,N_14157,N_14527);
and UO_1844 (O_1844,N_14781,N_14033);
or UO_1845 (O_1845,N_14879,N_14352);
xor UO_1846 (O_1846,N_14980,N_14575);
nor UO_1847 (O_1847,N_14586,N_14042);
xor UO_1848 (O_1848,N_14445,N_14143);
xor UO_1849 (O_1849,N_14206,N_14382);
nor UO_1850 (O_1850,N_14165,N_14819);
or UO_1851 (O_1851,N_14037,N_14305);
xnor UO_1852 (O_1852,N_14383,N_14087);
nor UO_1853 (O_1853,N_14560,N_14228);
xor UO_1854 (O_1854,N_14605,N_14501);
or UO_1855 (O_1855,N_14907,N_14934);
or UO_1856 (O_1856,N_14021,N_14893);
xnor UO_1857 (O_1857,N_14620,N_14049);
nand UO_1858 (O_1858,N_14950,N_14084);
nand UO_1859 (O_1859,N_14875,N_14730);
nor UO_1860 (O_1860,N_14807,N_14050);
and UO_1861 (O_1861,N_14219,N_14518);
xnor UO_1862 (O_1862,N_14644,N_14811);
nor UO_1863 (O_1863,N_14956,N_14163);
and UO_1864 (O_1864,N_14393,N_14696);
xor UO_1865 (O_1865,N_14788,N_14773);
nor UO_1866 (O_1866,N_14886,N_14418);
nand UO_1867 (O_1867,N_14620,N_14897);
nor UO_1868 (O_1868,N_14068,N_14634);
nand UO_1869 (O_1869,N_14355,N_14240);
nor UO_1870 (O_1870,N_14137,N_14625);
xor UO_1871 (O_1871,N_14979,N_14830);
nand UO_1872 (O_1872,N_14658,N_14775);
xor UO_1873 (O_1873,N_14593,N_14312);
and UO_1874 (O_1874,N_14405,N_14915);
and UO_1875 (O_1875,N_14184,N_14349);
or UO_1876 (O_1876,N_14651,N_14523);
nand UO_1877 (O_1877,N_14122,N_14682);
xnor UO_1878 (O_1878,N_14266,N_14332);
nand UO_1879 (O_1879,N_14013,N_14369);
or UO_1880 (O_1880,N_14152,N_14368);
or UO_1881 (O_1881,N_14880,N_14782);
or UO_1882 (O_1882,N_14924,N_14622);
xor UO_1883 (O_1883,N_14838,N_14675);
nor UO_1884 (O_1884,N_14183,N_14203);
nand UO_1885 (O_1885,N_14472,N_14336);
and UO_1886 (O_1886,N_14286,N_14816);
or UO_1887 (O_1887,N_14484,N_14029);
nor UO_1888 (O_1888,N_14272,N_14997);
nand UO_1889 (O_1889,N_14496,N_14765);
and UO_1890 (O_1890,N_14553,N_14970);
and UO_1891 (O_1891,N_14351,N_14406);
and UO_1892 (O_1892,N_14345,N_14474);
nand UO_1893 (O_1893,N_14550,N_14743);
or UO_1894 (O_1894,N_14917,N_14107);
nor UO_1895 (O_1895,N_14692,N_14606);
and UO_1896 (O_1896,N_14796,N_14101);
xnor UO_1897 (O_1897,N_14545,N_14859);
nand UO_1898 (O_1898,N_14395,N_14948);
and UO_1899 (O_1899,N_14265,N_14441);
xor UO_1900 (O_1900,N_14812,N_14327);
and UO_1901 (O_1901,N_14415,N_14161);
or UO_1902 (O_1902,N_14375,N_14402);
or UO_1903 (O_1903,N_14256,N_14321);
xor UO_1904 (O_1904,N_14395,N_14802);
nor UO_1905 (O_1905,N_14581,N_14347);
nand UO_1906 (O_1906,N_14978,N_14969);
and UO_1907 (O_1907,N_14488,N_14213);
and UO_1908 (O_1908,N_14032,N_14996);
or UO_1909 (O_1909,N_14963,N_14748);
xnor UO_1910 (O_1910,N_14376,N_14099);
nor UO_1911 (O_1911,N_14859,N_14022);
or UO_1912 (O_1912,N_14176,N_14293);
nor UO_1913 (O_1913,N_14992,N_14965);
and UO_1914 (O_1914,N_14519,N_14067);
nor UO_1915 (O_1915,N_14032,N_14681);
or UO_1916 (O_1916,N_14368,N_14494);
nand UO_1917 (O_1917,N_14655,N_14110);
xor UO_1918 (O_1918,N_14277,N_14901);
nor UO_1919 (O_1919,N_14876,N_14566);
or UO_1920 (O_1920,N_14176,N_14406);
or UO_1921 (O_1921,N_14200,N_14779);
nor UO_1922 (O_1922,N_14558,N_14135);
xnor UO_1923 (O_1923,N_14493,N_14322);
and UO_1924 (O_1924,N_14319,N_14529);
nand UO_1925 (O_1925,N_14779,N_14917);
and UO_1926 (O_1926,N_14974,N_14955);
xnor UO_1927 (O_1927,N_14231,N_14115);
nand UO_1928 (O_1928,N_14553,N_14348);
or UO_1929 (O_1929,N_14403,N_14344);
xor UO_1930 (O_1930,N_14222,N_14442);
xor UO_1931 (O_1931,N_14733,N_14959);
or UO_1932 (O_1932,N_14745,N_14463);
and UO_1933 (O_1933,N_14460,N_14359);
xnor UO_1934 (O_1934,N_14570,N_14070);
nor UO_1935 (O_1935,N_14269,N_14729);
or UO_1936 (O_1936,N_14556,N_14856);
nor UO_1937 (O_1937,N_14121,N_14426);
nor UO_1938 (O_1938,N_14762,N_14243);
and UO_1939 (O_1939,N_14331,N_14718);
xor UO_1940 (O_1940,N_14510,N_14461);
xor UO_1941 (O_1941,N_14465,N_14598);
xnor UO_1942 (O_1942,N_14359,N_14010);
and UO_1943 (O_1943,N_14588,N_14652);
and UO_1944 (O_1944,N_14550,N_14050);
or UO_1945 (O_1945,N_14382,N_14835);
nand UO_1946 (O_1946,N_14691,N_14820);
xnor UO_1947 (O_1947,N_14841,N_14072);
nor UO_1948 (O_1948,N_14274,N_14128);
xor UO_1949 (O_1949,N_14779,N_14819);
and UO_1950 (O_1950,N_14481,N_14365);
xnor UO_1951 (O_1951,N_14213,N_14952);
or UO_1952 (O_1952,N_14675,N_14378);
and UO_1953 (O_1953,N_14632,N_14902);
and UO_1954 (O_1954,N_14008,N_14711);
xor UO_1955 (O_1955,N_14366,N_14365);
and UO_1956 (O_1956,N_14958,N_14320);
and UO_1957 (O_1957,N_14751,N_14580);
or UO_1958 (O_1958,N_14272,N_14445);
or UO_1959 (O_1959,N_14442,N_14915);
nor UO_1960 (O_1960,N_14844,N_14547);
nor UO_1961 (O_1961,N_14537,N_14660);
or UO_1962 (O_1962,N_14700,N_14812);
nand UO_1963 (O_1963,N_14647,N_14473);
nand UO_1964 (O_1964,N_14104,N_14875);
nor UO_1965 (O_1965,N_14304,N_14006);
xor UO_1966 (O_1966,N_14158,N_14385);
and UO_1967 (O_1967,N_14888,N_14395);
xor UO_1968 (O_1968,N_14950,N_14382);
and UO_1969 (O_1969,N_14942,N_14176);
or UO_1970 (O_1970,N_14454,N_14586);
nor UO_1971 (O_1971,N_14451,N_14419);
nor UO_1972 (O_1972,N_14802,N_14599);
and UO_1973 (O_1973,N_14831,N_14485);
xor UO_1974 (O_1974,N_14571,N_14411);
nand UO_1975 (O_1975,N_14583,N_14899);
and UO_1976 (O_1976,N_14774,N_14412);
and UO_1977 (O_1977,N_14420,N_14965);
nor UO_1978 (O_1978,N_14027,N_14661);
or UO_1979 (O_1979,N_14044,N_14189);
xor UO_1980 (O_1980,N_14043,N_14593);
nand UO_1981 (O_1981,N_14415,N_14376);
or UO_1982 (O_1982,N_14585,N_14963);
and UO_1983 (O_1983,N_14115,N_14589);
and UO_1984 (O_1984,N_14998,N_14593);
xor UO_1985 (O_1985,N_14542,N_14469);
xnor UO_1986 (O_1986,N_14434,N_14024);
nand UO_1987 (O_1987,N_14827,N_14384);
nor UO_1988 (O_1988,N_14864,N_14977);
nand UO_1989 (O_1989,N_14191,N_14646);
nand UO_1990 (O_1990,N_14806,N_14681);
xnor UO_1991 (O_1991,N_14703,N_14116);
or UO_1992 (O_1992,N_14970,N_14995);
nand UO_1993 (O_1993,N_14264,N_14039);
nor UO_1994 (O_1994,N_14560,N_14756);
nor UO_1995 (O_1995,N_14473,N_14401);
nand UO_1996 (O_1996,N_14208,N_14115);
nor UO_1997 (O_1997,N_14925,N_14314);
nand UO_1998 (O_1998,N_14948,N_14508);
xnor UO_1999 (O_1999,N_14891,N_14649);
endmodule