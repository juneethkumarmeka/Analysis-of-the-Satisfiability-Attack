module basic_1000_10000_1500_4_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_368,In_465);
and U1 (N_1,In_313,In_376);
or U2 (N_2,In_576,In_998);
nand U3 (N_3,In_686,In_370);
or U4 (N_4,In_191,In_121);
nand U5 (N_5,In_603,In_25);
nor U6 (N_6,In_402,In_839);
nor U7 (N_7,In_367,In_705);
or U8 (N_8,In_981,In_428);
or U9 (N_9,In_305,In_371);
nand U10 (N_10,In_444,In_909);
xnor U11 (N_11,In_729,In_627);
and U12 (N_12,In_299,In_386);
nand U13 (N_13,In_393,In_12);
nor U14 (N_14,In_319,In_252);
xnor U15 (N_15,In_961,In_820);
and U16 (N_16,In_274,In_82);
nor U17 (N_17,In_118,In_328);
nand U18 (N_18,In_90,In_674);
and U19 (N_19,In_356,In_267);
or U20 (N_20,In_427,In_993);
and U21 (N_21,In_460,In_492);
nor U22 (N_22,In_680,In_872);
or U23 (N_23,In_781,In_303);
or U24 (N_24,In_439,In_149);
xnor U25 (N_25,In_726,In_631);
nor U26 (N_26,In_525,In_296);
nand U27 (N_27,In_780,In_792);
xnor U28 (N_28,In_553,In_81);
nor U29 (N_29,In_84,In_656);
nor U30 (N_30,In_456,In_441);
and U31 (N_31,In_298,In_33);
or U32 (N_32,In_752,In_203);
or U33 (N_33,In_127,In_128);
xor U34 (N_34,In_806,In_504);
or U35 (N_35,In_589,In_2);
and U36 (N_36,In_103,In_355);
nand U37 (N_37,In_605,In_32);
nand U38 (N_38,In_5,In_623);
or U39 (N_39,In_440,In_655);
nand U40 (N_40,In_206,In_881);
nor U41 (N_41,In_60,In_707);
nor U42 (N_42,In_99,In_249);
nand U43 (N_43,In_162,In_31);
xor U44 (N_44,In_884,In_721);
nor U45 (N_45,In_475,In_934);
or U46 (N_46,In_258,In_119);
nor U47 (N_47,In_192,In_116);
nand U48 (N_48,In_836,In_843);
or U49 (N_49,In_777,In_636);
and U50 (N_50,In_422,In_442);
xnor U51 (N_51,In_600,In_970);
xor U52 (N_52,In_858,In_318);
and U53 (N_53,In_459,In_415);
and U54 (N_54,In_113,In_885);
nor U55 (N_55,In_886,In_853);
and U56 (N_56,In_26,In_276);
nand U57 (N_57,In_96,In_50);
or U58 (N_58,In_754,In_129);
nor U59 (N_59,In_642,In_698);
and U60 (N_60,In_41,In_932);
nand U61 (N_61,In_30,In_659);
and U62 (N_62,In_351,In_247);
or U63 (N_63,In_257,In_300);
and U64 (N_64,In_408,In_384);
xnor U65 (N_65,In_547,In_329);
xnor U66 (N_66,In_95,In_180);
nor U67 (N_67,In_530,In_581);
or U68 (N_68,In_542,In_816);
or U69 (N_69,In_235,In_764);
or U70 (N_70,In_864,In_464);
nor U71 (N_71,In_549,In_529);
xnor U72 (N_72,In_317,In_683);
nor U73 (N_73,In_785,In_900);
and U74 (N_74,In_652,In_874);
nor U75 (N_75,In_394,In_353);
nor U76 (N_76,In_234,In_463);
nand U77 (N_77,In_702,In_972);
or U78 (N_78,In_811,In_828);
nand U79 (N_79,In_759,In_722);
nand U80 (N_80,In_499,In_633);
nand U81 (N_81,In_143,In_124);
and U82 (N_82,In_221,In_878);
or U83 (N_83,In_832,In_115);
or U84 (N_84,In_395,In_724);
nand U85 (N_85,In_995,In_323);
xor U86 (N_86,In_20,In_924);
nand U87 (N_87,In_526,In_834);
nor U88 (N_88,In_967,In_689);
xor U89 (N_89,In_228,In_174);
or U90 (N_90,In_937,In_434);
nand U91 (N_91,In_810,In_331);
xnor U92 (N_92,In_582,In_840);
xor U93 (N_93,In_406,In_639);
nor U94 (N_94,In_264,In_378);
nand U95 (N_95,In_420,In_342);
or U96 (N_96,In_75,In_193);
xnor U97 (N_97,In_933,In_256);
nand U98 (N_98,In_560,In_915);
nor U99 (N_99,In_634,In_23);
or U100 (N_100,In_541,In_69);
and U101 (N_101,In_546,In_288);
nor U102 (N_102,In_346,In_158);
xor U103 (N_103,In_963,In_18);
nor U104 (N_104,In_848,In_992);
nand U105 (N_105,In_169,In_518);
nand U106 (N_106,In_808,In_941);
xor U107 (N_107,In_629,In_154);
or U108 (N_108,In_105,In_663);
nor U109 (N_109,In_22,In_246);
nor U110 (N_110,In_573,In_562);
and U111 (N_111,In_958,In_760);
or U112 (N_112,In_965,In_311);
or U113 (N_113,In_374,In_259);
xor U114 (N_114,In_215,In_350);
nor U115 (N_115,In_236,In_521);
xor U116 (N_116,In_163,In_423);
or U117 (N_117,In_142,In_513);
nand U118 (N_118,In_641,In_845);
xor U119 (N_119,In_438,In_93);
nor U120 (N_120,In_635,In_97);
nor U121 (N_121,In_467,In_731);
xor U122 (N_122,In_92,In_385);
xor U123 (N_123,In_742,In_260);
xor U124 (N_124,In_672,In_536);
nor U125 (N_125,In_263,In_833);
nor U126 (N_126,In_57,In_111);
nand U127 (N_127,In_502,In_640);
or U128 (N_128,In_988,In_156);
nor U129 (N_129,In_59,In_114);
and U130 (N_130,In_925,In_52);
nand U131 (N_131,In_125,In_667);
nand U132 (N_132,In_574,In_102);
nand U133 (N_133,In_744,In_265);
and U134 (N_134,In_857,In_272);
nor U135 (N_135,In_47,In_891);
or U136 (N_136,In_682,In_852);
nand U137 (N_137,In_533,In_939);
nor U138 (N_138,In_185,In_743);
and U139 (N_139,In_150,In_822);
xnor U140 (N_140,In_363,In_910);
nor U141 (N_141,In_799,In_851);
or U142 (N_142,In_120,In_849);
xor U143 (N_143,In_737,In_804);
or U144 (N_144,In_710,In_271);
and U145 (N_145,In_280,In_45);
nor U146 (N_146,In_658,In_622);
or U147 (N_147,In_916,In_575);
nand U148 (N_148,In_68,In_40);
nand U149 (N_149,In_468,In_784);
and U150 (N_150,In_486,In_903);
or U151 (N_151,In_39,In_196);
and U152 (N_152,In_229,In_644);
and U153 (N_153,In_951,In_74);
nor U154 (N_154,In_699,In_889);
or U155 (N_155,In_137,In_223);
and U156 (N_156,In_283,In_865);
nand U157 (N_157,In_83,In_746);
nand U158 (N_158,In_362,In_58);
nor U159 (N_159,In_245,In_380);
nand U160 (N_160,In_94,In_918);
and U161 (N_161,In_159,In_835);
and U162 (N_162,In_692,In_66);
and U163 (N_163,In_268,In_70);
nor U164 (N_164,In_955,In_358);
nand U165 (N_165,In_190,In_253);
and U166 (N_166,In_330,In_776);
or U167 (N_167,In_231,In_36);
nand U168 (N_168,In_333,In_433);
xnor U169 (N_169,In_572,In_999);
or U170 (N_170,In_819,In_21);
xor U171 (N_171,In_867,In_711);
nor U172 (N_172,In_585,In_130);
nand U173 (N_173,In_237,In_117);
xnor U174 (N_174,In_275,In_315);
or U175 (N_175,In_500,In_261);
xnor U176 (N_176,In_814,In_568);
nor U177 (N_177,In_487,In_497);
nor U178 (N_178,In_586,In_902);
nand U179 (N_179,In_557,In_210);
and U180 (N_180,In_239,In_179);
nor U181 (N_181,In_314,In_134);
and U182 (N_182,In_449,In_519);
or U183 (N_183,In_751,In_919);
xnor U184 (N_184,In_873,In_322);
or U185 (N_185,In_991,In_3);
and U186 (N_186,In_681,In_278);
xnor U187 (N_187,In_688,In_653);
nor U188 (N_188,In_501,In_11);
nor U189 (N_189,In_930,In_396);
nor U190 (N_190,In_602,In_607);
or U191 (N_191,In_827,In_167);
and U192 (N_192,In_880,In_701);
nand U193 (N_193,In_517,In_352);
and U194 (N_194,In_15,In_953);
and U195 (N_195,In_282,In_982);
and U196 (N_196,In_212,In_462);
nand U197 (N_197,In_997,In_977);
and U198 (N_198,In_301,In_382);
xnor U199 (N_199,In_205,In_986);
and U200 (N_200,In_709,In_676);
nor U201 (N_201,In_757,In_430);
and U202 (N_202,In_860,In_42);
nand U203 (N_203,In_620,In_431);
xnor U204 (N_204,In_304,In_898);
nor U205 (N_205,In_775,In_78);
or U206 (N_206,In_1,In_454);
or U207 (N_207,In_364,In_535);
nand U208 (N_208,In_8,In_537);
nor U209 (N_209,In_911,In_369);
nor U210 (N_210,In_250,In_291);
or U211 (N_211,In_720,In_324);
nand U212 (N_212,In_238,In_690);
and U213 (N_213,In_522,In_453);
and U214 (N_214,In_146,In_509);
nand U215 (N_215,In_326,In_387);
nor U216 (N_216,In_591,In_877);
or U217 (N_217,In_532,In_110);
nor U218 (N_218,In_98,In_336);
nor U219 (N_219,In_490,In_85);
or U220 (N_220,In_214,In_365);
or U221 (N_221,In_426,In_470);
nand U222 (N_222,In_178,In_728);
nor U223 (N_223,In_354,In_649);
nor U224 (N_224,In_974,In_771);
nor U225 (N_225,In_375,In_181);
and U226 (N_226,In_863,In_233);
nand U227 (N_227,In_875,In_461);
or U228 (N_228,In_748,In_538);
or U229 (N_229,In_978,In_989);
or U230 (N_230,In_379,In_971);
or U231 (N_231,In_347,In_604);
or U232 (N_232,In_917,In_184);
xor U233 (N_233,In_739,In_209);
nor U234 (N_234,In_309,In_53);
nor U235 (N_235,In_778,In_44);
and U236 (N_236,In_914,In_7);
nor U237 (N_237,In_100,In_71);
or U238 (N_238,In_392,In_928);
and U239 (N_239,In_929,In_197);
nand U240 (N_240,In_964,In_716);
and U241 (N_241,In_213,In_446);
and U242 (N_242,In_227,In_173);
or U243 (N_243,In_388,In_225);
xnor U244 (N_244,In_801,In_0);
xnor U245 (N_245,In_219,In_452);
nor U246 (N_246,In_199,In_651);
nand U247 (N_247,In_766,In_590);
xnor U248 (N_248,In_165,In_505);
and U249 (N_249,In_908,In_222);
and U250 (N_250,In_132,In_139);
or U251 (N_251,In_477,In_638);
xnor U252 (N_252,In_170,In_548);
nor U253 (N_253,In_65,In_512);
nand U254 (N_254,In_944,In_782);
and U255 (N_255,In_554,In_940);
and U256 (N_256,In_664,In_335);
or U257 (N_257,In_14,In_484);
nand U258 (N_258,In_745,In_412);
nor U259 (N_259,In_401,In_284);
xor U260 (N_260,In_935,In_64);
nor U261 (N_261,In_482,In_841);
nand U262 (N_262,In_515,In_520);
and U263 (N_263,In_725,In_344);
and U264 (N_264,In_949,In_9);
xnor U265 (N_265,In_957,In_826);
and U266 (N_266,In_51,In_62);
or U267 (N_267,In_77,In_232);
nand U268 (N_268,In_896,In_437);
xor U269 (N_269,In_545,In_262);
nor U270 (N_270,In_244,In_443);
nor U271 (N_271,In_740,In_703);
and U272 (N_272,In_24,In_708);
or U273 (N_273,In_567,In_63);
nor U274 (N_274,In_421,In_101);
and U275 (N_275,In_947,In_779);
nor U276 (N_276,In_34,In_540);
nand U277 (N_277,In_104,In_691);
or U278 (N_278,In_770,In_618);
and U279 (N_279,In_593,In_194);
or U280 (N_280,In_558,In_145);
and U281 (N_281,In_416,In_962);
xor U282 (N_282,In_140,In_73);
and U283 (N_283,In_838,In_306);
nand U284 (N_284,In_469,In_802);
nor U285 (N_285,In_450,In_800);
nor U286 (N_286,In_601,In_447);
xor U287 (N_287,In_458,In_398);
or U288 (N_288,In_417,In_534);
nand U289 (N_289,In_507,In_543);
or U290 (N_290,In_606,In_292);
nor U291 (N_291,In_187,In_905);
xnor U292 (N_292,In_56,In_678);
nand U293 (N_293,In_281,In_868);
nand U294 (N_294,In_55,In_768);
nor U295 (N_295,In_783,In_657);
xnor U296 (N_296,In_931,In_866);
nor U297 (N_297,In_208,In_666);
xor U298 (N_298,In_155,In_88);
or U299 (N_299,In_609,In_308);
nor U300 (N_300,In_307,In_43);
and U301 (N_301,In_825,In_736);
and U302 (N_302,In_735,In_767);
nor U303 (N_303,In_481,In_798);
nand U304 (N_304,In_859,In_337);
nand U305 (N_305,In_942,In_508);
or U306 (N_306,In_587,In_619);
or U307 (N_307,In_334,In_566);
xor U308 (N_308,In_144,In_87);
nand U309 (N_309,In_290,In_630);
and U310 (N_310,In_645,In_493);
or U311 (N_311,In_687,In_455);
nor U312 (N_312,In_815,In_220);
xnor U313 (N_313,In_890,In_407);
or U314 (N_314,In_183,In_425);
and U315 (N_315,In_797,In_432);
nor U316 (N_316,In_157,In_943);
nor U317 (N_317,In_251,In_13);
xnor U318 (N_318,In_539,In_413);
and U319 (N_319,In_37,In_954);
xnor U320 (N_320,In_54,In_202);
and U321 (N_321,In_550,In_528);
nand U322 (N_322,In_38,In_706);
xnor U323 (N_323,In_171,In_847);
and U324 (N_324,In_624,In_429);
nand U325 (N_325,In_803,In_632);
xnor U326 (N_326,In_795,In_791);
or U327 (N_327,In_531,In_474);
xor U328 (N_328,In_109,In_414);
or U329 (N_329,In_503,In_926);
nor U330 (N_330,In_479,In_790);
or U331 (N_331,In_491,In_559);
nor U332 (N_332,In_599,In_489);
nor U333 (N_333,In_749,In_793);
nor U334 (N_334,In_359,In_189);
or U335 (N_335,In_817,In_200);
xnor U336 (N_336,In_694,In_86);
and U337 (N_337,In_17,In_769);
nor U338 (N_338,In_869,In_389);
nor U339 (N_339,In_610,In_277);
or U340 (N_340,In_883,In_854);
xnor U341 (N_341,In_823,In_621);
nand U342 (N_342,In_987,In_399);
and U343 (N_343,In_168,In_611);
and U344 (N_344,In_661,In_108);
nor U345 (N_345,In_765,In_787);
nor U346 (N_346,In_968,In_671);
and U347 (N_347,In_693,In_391);
nor U348 (N_348,In_812,In_161);
nor U349 (N_349,In_166,In_138);
and U350 (N_350,In_985,In_913);
and U351 (N_351,In_871,In_718);
xnor U352 (N_352,In_662,In_218);
or U353 (N_353,In_626,In_552);
nor U354 (N_354,In_584,In_608);
nor U355 (N_355,In_279,In_879);
nand U356 (N_356,In_16,In_106);
and U357 (N_357,In_856,In_4);
or U358 (N_358,In_451,In_295);
nor U359 (N_359,In_485,In_48);
xnor U360 (N_360,In_435,In_654);
nand U361 (N_361,In_152,In_466);
and U362 (N_362,In_471,In_758);
nor U363 (N_363,In_842,In_660);
and U364 (N_364,In_28,In_400);
nor U365 (N_365,In_445,In_887);
xor U366 (N_366,In_677,In_506);
xor U367 (N_367,In_579,In_756);
nand U368 (N_368,In_571,In_325);
xor U369 (N_369,In_946,In_457);
nand U370 (N_370,In_405,In_418);
and U371 (N_371,In_616,In_224);
and U372 (N_372,In_226,In_945);
or U373 (N_373,In_561,In_821);
and U374 (N_374,In_950,In_478);
or U375 (N_375,In_670,In_556);
and U376 (N_376,In_516,In_696);
nand U377 (N_377,In_569,In_809);
nand U378 (N_378,In_813,In_927);
nand U379 (N_379,In_788,In_46);
nor U380 (N_380,In_870,In_357);
and U381 (N_381,In_348,In_147);
xor U382 (N_382,In_983,In_476);
xor U383 (N_383,In_523,In_888);
and U384 (N_384,In_302,In_80);
or U385 (N_385,In_175,In_270);
nor U386 (N_386,In_480,In_498);
and U387 (N_387,In_381,In_254);
or U388 (N_388,In_555,In_794);
nand U389 (N_389,In_126,In_207);
nor U390 (N_390,In_29,In_973);
and U391 (N_391,In_483,In_789);
nor U392 (N_392,In_133,In_597);
nor U393 (N_393,In_327,In_565);
xor U394 (N_394,In_390,In_772);
xor U395 (N_395,In_818,In_240);
or U396 (N_396,In_959,In_182);
and U397 (N_397,In_894,In_614);
nor U398 (N_398,In_920,In_637);
xnor U399 (N_399,In_19,In_293);
and U400 (N_400,In_360,In_366);
xnor U401 (N_401,In_730,In_738);
xor U402 (N_402,In_266,In_665);
nor U403 (N_403,In_831,In_316);
and U404 (N_404,In_979,In_829);
xnor U405 (N_405,In_527,In_976);
and U406 (N_406,In_89,In_172);
and U407 (N_407,In_321,In_122);
and U408 (N_408,In_844,In_10);
or U409 (N_409,In_289,In_273);
and U410 (N_410,In_901,In_343);
or U411 (N_411,In_613,In_732);
nor U412 (N_412,In_862,In_612);
or U413 (N_413,In_141,In_876);
and U414 (N_414,In_176,In_773);
nor U415 (N_415,In_948,In_669);
or U416 (N_416,In_938,In_980);
and U417 (N_417,In_824,In_424);
xnor U418 (N_418,In_960,In_753);
xor U419 (N_419,In_216,In_675);
or U420 (N_420,In_6,In_700);
xnor U421 (N_421,In_830,In_312);
nand U422 (N_422,In_338,In_419);
xnor U423 (N_423,In_846,In_715);
nor U424 (N_424,In_341,In_345);
nand U425 (N_425,In_695,In_112);
nand U426 (N_426,In_592,In_761);
and U427 (N_427,In_741,In_211);
xnor U428 (N_428,In_135,In_294);
or U429 (N_429,In_598,In_164);
nor U430 (N_430,In_511,In_595);
xor U431 (N_431,In_248,In_61);
and U432 (N_432,In_850,In_403);
or U433 (N_433,In_747,In_763);
or U434 (N_434,In_975,In_855);
and U435 (N_435,In_123,In_628);
nor U436 (N_436,In_241,In_996);
and U437 (N_437,In_892,In_966);
and U438 (N_438,In_310,In_684);
or U439 (N_439,In_733,In_936);
or U440 (N_440,In_410,In_243);
nor U441 (N_441,In_339,In_242);
or U442 (N_442,In_712,In_151);
nand U443 (N_443,In_837,In_679);
nand U444 (N_444,In_899,In_136);
and U445 (N_445,In_160,In_195);
or U446 (N_446,In_922,In_588);
xnor U447 (N_447,In_177,In_969);
or U448 (N_448,In_990,In_727);
xor U449 (N_449,In_495,In_786);
xnor U450 (N_450,In_580,In_131);
and U451 (N_451,In_79,In_72);
and U452 (N_452,In_332,In_564);
nor U453 (N_453,In_397,In_668);
xnor U454 (N_454,In_340,In_255);
or U455 (N_455,In_488,In_956);
or U456 (N_456,In_188,In_646);
nor U457 (N_457,In_372,In_912);
xor U458 (N_458,In_615,In_409);
nand U459 (N_459,In_49,In_895);
or U460 (N_460,In_230,In_551);
nand U461 (N_461,In_186,In_750);
nand U462 (N_462,In_472,In_411);
xor U463 (N_463,In_320,In_383);
or U464 (N_464,In_906,In_882);
nor U465 (N_465,In_719,In_201);
and U466 (N_466,In_27,In_373);
and U467 (N_467,In_448,In_377);
nand U468 (N_468,In_704,In_286);
xor U469 (N_469,In_578,In_514);
or U470 (N_470,In_76,In_685);
and U471 (N_471,In_861,In_650);
nand U472 (N_472,In_594,In_897);
xnor U473 (N_473,In_807,In_904);
xor U474 (N_474,In_723,In_805);
nor U475 (N_475,In_625,In_734);
xor U476 (N_476,In_287,In_148);
xor U477 (N_477,In_697,In_510);
and U478 (N_478,In_217,In_893);
and U479 (N_479,In_577,In_907);
and U480 (N_480,In_643,In_494);
xnor U481 (N_481,In_361,In_713);
nand U482 (N_482,In_755,In_570);
nor U483 (N_483,In_35,In_269);
and U484 (N_484,In_544,In_297);
nand U485 (N_485,In_107,In_921);
nand U486 (N_486,In_563,In_617);
or U487 (N_487,In_774,In_648);
or U488 (N_488,In_762,In_994);
nor U489 (N_489,In_198,In_404);
nand U490 (N_490,In_349,In_473);
nand U491 (N_491,In_524,In_952);
nor U492 (N_492,In_714,In_673);
nand U493 (N_493,In_436,In_67);
nor U494 (N_494,In_984,In_204);
nor U495 (N_495,In_717,In_583);
nor U496 (N_496,In_153,In_285);
nor U497 (N_497,In_923,In_647);
nor U498 (N_498,In_91,In_796);
or U499 (N_499,In_496,In_596);
and U500 (N_500,In_488,In_146);
nor U501 (N_501,In_501,In_110);
xnor U502 (N_502,In_527,In_922);
and U503 (N_503,In_698,In_261);
and U504 (N_504,In_70,In_198);
and U505 (N_505,In_636,In_467);
nand U506 (N_506,In_793,In_361);
xor U507 (N_507,In_300,In_265);
nor U508 (N_508,In_818,In_225);
nand U509 (N_509,In_874,In_18);
and U510 (N_510,In_706,In_718);
or U511 (N_511,In_867,In_494);
and U512 (N_512,In_65,In_229);
or U513 (N_513,In_139,In_679);
and U514 (N_514,In_357,In_84);
nand U515 (N_515,In_913,In_635);
nand U516 (N_516,In_36,In_980);
nor U517 (N_517,In_704,In_380);
nand U518 (N_518,In_85,In_672);
nand U519 (N_519,In_119,In_611);
or U520 (N_520,In_394,In_466);
or U521 (N_521,In_854,In_769);
and U522 (N_522,In_607,In_836);
and U523 (N_523,In_413,In_130);
or U524 (N_524,In_46,In_66);
nand U525 (N_525,In_925,In_162);
and U526 (N_526,In_559,In_211);
or U527 (N_527,In_936,In_17);
or U528 (N_528,In_665,In_204);
nand U529 (N_529,In_139,In_763);
or U530 (N_530,In_860,In_755);
or U531 (N_531,In_326,In_304);
nor U532 (N_532,In_351,In_495);
xor U533 (N_533,In_664,In_202);
nor U534 (N_534,In_901,In_980);
xnor U535 (N_535,In_662,In_865);
xor U536 (N_536,In_365,In_742);
and U537 (N_537,In_806,In_610);
and U538 (N_538,In_996,In_564);
nand U539 (N_539,In_824,In_813);
xnor U540 (N_540,In_787,In_658);
xor U541 (N_541,In_773,In_198);
nand U542 (N_542,In_254,In_397);
nand U543 (N_543,In_529,In_339);
nor U544 (N_544,In_563,In_0);
nand U545 (N_545,In_686,In_907);
and U546 (N_546,In_874,In_165);
and U547 (N_547,In_861,In_113);
or U548 (N_548,In_582,In_822);
or U549 (N_549,In_642,In_726);
and U550 (N_550,In_755,In_714);
xnor U551 (N_551,In_708,In_304);
or U552 (N_552,In_383,In_761);
nor U553 (N_553,In_375,In_499);
and U554 (N_554,In_98,In_356);
xor U555 (N_555,In_21,In_476);
or U556 (N_556,In_843,In_214);
nand U557 (N_557,In_844,In_462);
nand U558 (N_558,In_895,In_465);
and U559 (N_559,In_398,In_254);
nor U560 (N_560,In_172,In_528);
or U561 (N_561,In_500,In_763);
xnor U562 (N_562,In_962,In_534);
xor U563 (N_563,In_372,In_466);
nand U564 (N_564,In_570,In_378);
and U565 (N_565,In_841,In_229);
nand U566 (N_566,In_487,In_509);
and U567 (N_567,In_148,In_59);
and U568 (N_568,In_524,In_722);
nand U569 (N_569,In_367,In_543);
or U570 (N_570,In_366,In_284);
nand U571 (N_571,In_928,In_555);
nand U572 (N_572,In_763,In_134);
nor U573 (N_573,In_664,In_474);
and U574 (N_574,In_653,In_112);
nor U575 (N_575,In_529,In_635);
nand U576 (N_576,In_569,In_226);
and U577 (N_577,In_710,In_550);
xnor U578 (N_578,In_386,In_739);
nor U579 (N_579,In_951,In_48);
nor U580 (N_580,In_330,In_950);
nor U581 (N_581,In_913,In_385);
nand U582 (N_582,In_327,In_113);
and U583 (N_583,In_803,In_982);
nor U584 (N_584,In_670,In_660);
nand U585 (N_585,In_692,In_211);
or U586 (N_586,In_732,In_921);
nor U587 (N_587,In_773,In_183);
nand U588 (N_588,In_289,In_378);
nor U589 (N_589,In_466,In_449);
and U590 (N_590,In_70,In_803);
xor U591 (N_591,In_663,In_808);
nor U592 (N_592,In_899,In_115);
and U593 (N_593,In_818,In_348);
xor U594 (N_594,In_833,In_858);
or U595 (N_595,In_496,In_82);
nor U596 (N_596,In_124,In_531);
nand U597 (N_597,In_163,In_45);
nand U598 (N_598,In_88,In_433);
nor U599 (N_599,In_260,In_797);
and U600 (N_600,In_918,In_847);
and U601 (N_601,In_220,In_571);
xnor U602 (N_602,In_297,In_859);
xor U603 (N_603,In_661,In_172);
nand U604 (N_604,In_461,In_196);
and U605 (N_605,In_697,In_475);
or U606 (N_606,In_782,In_679);
nor U607 (N_607,In_109,In_752);
or U608 (N_608,In_820,In_468);
nand U609 (N_609,In_943,In_186);
xnor U610 (N_610,In_100,In_2);
xor U611 (N_611,In_922,In_786);
nor U612 (N_612,In_598,In_346);
xnor U613 (N_613,In_214,In_341);
or U614 (N_614,In_713,In_661);
and U615 (N_615,In_91,In_942);
nand U616 (N_616,In_197,In_389);
nand U617 (N_617,In_709,In_786);
or U618 (N_618,In_951,In_755);
or U619 (N_619,In_161,In_57);
nand U620 (N_620,In_918,In_655);
and U621 (N_621,In_409,In_988);
xor U622 (N_622,In_411,In_833);
or U623 (N_623,In_40,In_902);
and U624 (N_624,In_268,In_443);
xnor U625 (N_625,In_663,In_631);
nor U626 (N_626,In_667,In_463);
and U627 (N_627,In_285,In_203);
xnor U628 (N_628,In_763,In_510);
and U629 (N_629,In_537,In_45);
nor U630 (N_630,In_897,In_24);
nand U631 (N_631,In_350,In_999);
xnor U632 (N_632,In_745,In_135);
nor U633 (N_633,In_710,In_263);
nand U634 (N_634,In_393,In_109);
or U635 (N_635,In_287,In_370);
xor U636 (N_636,In_871,In_222);
or U637 (N_637,In_226,In_646);
or U638 (N_638,In_436,In_157);
and U639 (N_639,In_540,In_111);
nand U640 (N_640,In_553,In_413);
xor U641 (N_641,In_354,In_416);
and U642 (N_642,In_342,In_974);
xor U643 (N_643,In_7,In_620);
xor U644 (N_644,In_189,In_517);
or U645 (N_645,In_930,In_313);
nand U646 (N_646,In_380,In_135);
and U647 (N_647,In_449,In_163);
nand U648 (N_648,In_633,In_628);
nand U649 (N_649,In_564,In_703);
nand U650 (N_650,In_24,In_445);
xor U651 (N_651,In_571,In_161);
or U652 (N_652,In_247,In_379);
nand U653 (N_653,In_335,In_734);
nand U654 (N_654,In_809,In_284);
nand U655 (N_655,In_812,In_958);
nand U656 (N_656,In_446,In_979);
xor U657 (N_657,In_458,In_234);
and U658 (N_658,In_423,In_776);
and U659 (N_659,In_738,In_104);
nand U660 (N_660,In_450,In_821);
nor U661 (N_661,In_356,In_508);
or U662 (N_662,In_267,In_825);
xor U663 (N_663,In_656,In_350);
xnor U664 (N_664,In_28,In_680);
nand U665 (N_665,In_4,In_294);
nor U666 (N_666,In_419,In_639);
xnor U667 (N_667,In_333,In_844);
xnor U668 (N_668,In_227,In_883);
xnor U669 (N_669,In_285,In_44);
or U670 (N_670,In_89,In_936);
nor U671 (N_671,In_509,In_147);
and U672 (N_672,In_644,In_602);
nand U673 (N_673,In_481,In_690);
xnor U674 (N_674,In_830,In_1);
nor U675 (N_675,In_958,In_841);
and U676 (N_676,In_172,In_351);
or U677 (N_677,In_914,In_848);
xor U678 (N_678,In_639,In_897);
nor U679 (N_679,In_723,In_758);
xor U680 (N_680,In_449,In_505);
or U681 (N_681,In_819,In_686);
and U682 (N_682,In_881,In_364);
nand U683 (N_683,In_690,In_585);
nand U684 (N_684,In_594,In_347);
nand U685 (N_685,In_85,In_728);
or U686 (N_686,In_621,In_115);
or U687 (N_687,In_261,In_613);
nor U688 (N_688,In_60,In_518);
and U689 (N_689,In_9,In_510);
nor U690 (N_690,In_264,In_676);
and U691 (N_691,In_430,In_475);
xnor U692 (N_692,In_323,In_28);
nor U693 (N_693,In_476,In_44);
nor U694 (N_694,In_110,In_548);
or U695 (N_695,In_746,In_846);
nand U696 (N_696,In_582,In_959);
and U697 (N_697,In_596,In_791);
and U698 (N_698,In_828,In_63);
and U699 (N_699,In_963,In_248);
or U700 (N_700,In_604,In_99);
xnor U701 (N_701,In_112,In_305);
nor U702 (N_702,In_524,In_454);
nor U703 (N_703,In_754,In_802);
and U704 (N_704,In_409,In_477);
or U705 (N_705,In_641,In_586);
and U706 (N_706,In_755,In_596);
xnor U707 (N_707,In_30,In_257);
and U708 (N_708,In_10,In_913);
nor U709 (N_709,In_617,In_263);
xor U710 (N_710,In_410,In_739);
nand U711 (N_711,In_161,In_326);
nor U712 (N_712,In_486,In_992);
xor U713 (N_713,In_425,In_88);
and U714 (N_714,In_929,In_137);
and U715 (N_715,In_817,In_373);
or U716 (N_716,In_146,In_956);
or U717 (N_717,In_689,In_719);
nor U718 (N_718,In_755,In_204);
nor U719 (N_719,In_90,In_651);
nor U720 (N_720,In_576,In_242);
or U721 (N_721,In_17,In_894);
or U722 (N_722,In_828,In_964);
and U723 (N_723,In_235,In_872);
or U724 (N_724,In_478,In_414);
nand U725 (N_725,In_537,In_774);
or U726 (N_726,In_384,In_471);
xnor U727 (N_727,In_982,In_824);
or U728 (N_728,In_140,In_106);
and U729 (N_729,In_687,In_795);
nand U730 (N_730,In_382,In_802);
xnor U731 (N_731,In_72,In_83);
and U732 (N_732,In_180,In_751);
nand U733 (N_733,In_97,In_731);
nand U734 (N_734,In_735,In_333);
xor U735 (N_735,In_851,In_766);
nor U736 (N_736,In_856,In_738);
nand U737 (N_737,In_550,In_86);
and U738 (N_738,In_357,In_830);
nand U739 (N_739,In_59,In_925);
xnor U740 (N_740,In_393,In_529);
nand U741 (N_741,In_116,In_119);
and U742 (N_742,In_947,In_281);
and U743 (N_743,In_947,In_56);
and U744 (N_744,In_486,In_117);
xnor U745 (N_745,In_949,In_92);
nand U746 (N_746,In_28,In_892);
xnor U747 (N_747,In_447,In_68);
xor U748 (N_748,In_531,In_728);
xor U749 (N_749,In_686,In_509);
xor U750 (N_750,In_265,In_4);
nand U751 (N_751,In_266,In_227);
nand U752 (N_752,In_405,In_300);
nor U753 (N_753,In_309,In_723);
or U754 (N_754,In_982,In_132);
xnor U755 (N_755,In_480,In_288);
nor U756 (N_756,In_944,In_616);
or U757 (N_757,In_803,In_905);
and U758 (N_758,In_174,In_408);
or U759 (N_759,In_228,In_229);
and U760 (N_760,In_122,In_897);
nor U761 (N_761,In_19,In_520);
xor U762 (N_762,In_211,In_778);
xnor U763 (N_763,In_419,In_520);
nor U764 (N_764,In_296,In_95);
and U765 (N_765,In_588,In_484);
nor U766 (N_766,In_220,In_338);
and U767 (N_767,In_816,In_291);
or U768 (N_768,In_595,In_105);
xnor U769 (N_769,In_396,In_20);
xor U770 (N_770,In_646,In_973);
xnor U771 (N_771,In_590,In_195);
nand U772 (N_772,In_657,In_560);
or U773 (N_773,In_413,In_732);
xnor U774 (N_774,In_406,In_189);
or U775 (N_775,In_795,In_432);
nor U776 (N_776,In_729,In_439);
or U777 (N_777,In_862,In_758);
nand U778 (N_778,In_414,In_871);
and U779 (N_779,In_332,In_68);
nand U780 (N_780,In_958,In_154);
nand U781 (N_781,In_288,In_236);
and U782 (N_782,In_896,In_701);
nand U783 (N_783,In_808,In_912);
xor U784 (N_784,In_104,In_125);
nor U785 (N_785,In_938,In_87);
or U786 (N_786,In_411,In_707);
nand U787 (N_787,In_959,In_447);
or U788 (N_788,In_388,In_807);
or U789 (N_789,In_662,In_10);
xor U790 (N_790,In_541,In_401);
and U791 (N_791,In_256,In_675);
and U792 (N_792,In_145,In_829);
and U793 (N_793,In_831,In_874);
nand U794 (N_794,In_449,In_654);
nand U795 (N_795,In_572,In_844);
nor U796 (N_796,In_109,In_134);
nand U797 (N_797,In_158,In_960);
nand U798 (N_798,In_783,In_506);
nand U799 (N_799,In_197,In_7);
xor U800 (N_800,In_437,In_272);
nand U801 (N_801,In_141,In_891);
nor U802 (N_802,In_80,In_655);
and U803 (N_803,In_377,In_950);
and U804 (N_804,In_339,In_198);
and U805 (N_805,In_589,In_535);
xor U806 (N_806,In_146,In_799);
xor U807 (N_807,In_952,In_22);
nand U808 (N_808,In_390,In_361);
and U809 (N_809,In_612,In_784);
xor U810 (N_810,In_381,In_29);
or U811 (N_811,In_740,In_142);
or U812 (N_812,In_754,In_223);
nand U813 (N_813,In_771,In_520);
xor U814 (N_814,In_62,In_528);
nor U815 (N_815,In_441,In_814);
nor U816 (N_816,In_861,In_294);
nand U817 (N_817,In_105,In_841);
nand U818 (N_818,In_532,In_162);
or U819 (N_819,In_867,In_265);
and U820 (N_820,In_20,In_686);
or U821 (N_821,In_884,In_562);
xor U822 (N_822,In_870,In_258);
xnor U823 (N_823,In_862,In_467);
or U824 (N_824,In_516,In_679);
nand U825 (N_825,In_122,In_358);
and U826 (N_826,In_657,In_8);
and U827 (N_827,In_657,In_728);
xor U828 (N_828,In_998,In_780);
and U829 (N_829,In_446,In_429);
xnor U830 (N_830,In_637,In_745);
or U831 (N_831,In_762,In_498);
nor U832 (N_832,In_574,In_522);
nand U833 (N_833,In_9,In_815);
and U834 (N_834,In_629,In_414);
nand U835 (N_835,In_664,In_268);
nor U836 (N_836,In_614,In_132);
or U837 (N_837,In_753,In_381);
and U838 (N_838,In_829,In_446);
nor U839 (N_839,In_734,In_839);
or U840 (N_840,In_676,In_621);
and U841 (N_841,In_338,In_140);
nor U842 (N_842,In_58,In_17);
nand U843 (N_843,In_796,In_54);
nand U844 (N_844,In_698,In_438);
or U845 (N_845,In_537,In_522);
nor U846 (N_846,In_395,In_887);
nand U847 (N_847,In_345,In_425);
nand U848 (N_848,In_186,In_909);
nor U849 (N_849,In_418,In_818);
nand U850 (N_850,In_359,In_323);
nand U851 (N_851,In_71,In_796);
nand U852 (N_852,In_227,In_488);
and U853 (N_853,In_592,In_795);
nand U854 (N_854,In_490,In_949);
nand U855 (N_855,In_765,In_214);
nor U856 (N_856,In_505,In_884);
xnor U857 (N_857,In_912,In_784);
and U858 (N_858,In_824,In_882);
nor U859 (N_859,In_305,In_887);
nor U860 (N_860,In_891,In_46);
xnor U861 (N_861,In_546,In_648);
nor U862 (N_862,In_829,In_582);
and U863 (N_863,In_522,In_485);
and U864 (N_864,In_501,In_930);
nor U865 (N_865,In_203,In_347);
xnor U866 (N_866,In_99,In_112);
nor U867 (N_867,In_954,In_852);
nand U868 (N_868,In_182,In_658);
xor U869 (N_869,In_282,In_555);
and U870 (N_870,In_210,In_856);
nand U871 (N_871,In_958,In_32);
and U872 (N_872,In_569,In_57);
nor U873 (N_873,In_151,In_23);
nor U874 (N_874,In_997,In_188);
xnor U875 (N_875,In_533,In_508);
nand U876 (N_876,In_588,In_100);
and U877 (N_877,In_193,In_545);
nor U878 (N_878,In_752,In_928);
nand U879 (N_879,In_194,In_351);
or U880 (N_880,In_311,In_849);
or U881 (N_881,In_531,In_840);
xor U882 (N_882,In_753,In_323);
nand U883 (N_883,In_504,In_689);
xnor U884 (N_884,In_653,In_709);
nor U885 (N_885,In_603,In_819);
or U886 (N_886,In_204,In_773);
nand U887 (N_887,In_453,In_699);
nor U888 (N_888,In_865,In_540);
or U889 (N_889,In_912,In_149);
nand U890 (N_890,In_87,In_478);
nor U891 (N_891,In_141,In_154);
xnor U892 (N_892,In_100,In_142);
and U893 (N_893,In_923,In_94);
nor U894 (N_894,In_664,In_831);
and U895 (N_895,In_232,In_616);
xor U896 (N_896,In_343,In_792);
nand U897 (N_897,In_982,In_919);
and U898 (N_898,In_945,In_910);
nor U899 (N_899,In_905,In_658);
xor U900 (N_900,In_520,In_229);
nand U901 (N_901,In_73,In_651);
nor U902 (N_902,In_241,In_605);
nor U903 (N_903,In_135,In_273);
nor U904 (N_904,In_995,In_821);
nor U905 (N_905,In_498,In_130);
xor U906 (N_906,In_270,In_781);
and U907 (N_907,In_576,In_219);
nand U908 (N_908,In_731,In_32);
or U909 (N_909,In_224,In_72);
or U910 (N_910,In_715,In_255);
or U911 (N_911,In_94,In_975);
or U912 (N_912,In_246,In_644);
xnor U913 (N_913,In_183,In_589);
xnor U914 (N_914,In_70,In_255);
and U915 (N_915,In_936,In_138);
nand U916 (N_916,In_210,In_358);
xor U917 (N_917,In_973,In_929);
xnor U918 (N_918,In_914,In_474);
nor U919 (N_919,In_13,In_306);
nand U920 (N_920,In_862,In_123);
and U921 (N_921,In_83,In_130);
nand U922 (N_922,In_349,In_403);
or U923 (N_923,In_833,In_116);
xor U924 (N_924,In_453,In_216);
and U925 (N_925,In_5,In_758);
xor U926 (N_926,In_712,In_305);
or U927 (N_927,In_348,In_956);
or U928 (N_928,In_818,In_398);
nor U929 (N_929,In_46,In_251);
nand U930 (N_930,In_154,In_81);
xor U931 (N_931,In_263,In_278);
xnor U932 (N_932,In_709,In_104);
nand U933 (N_933,In_63,In_821);
nand U934 (N_934,In_36,In_4);
nand U935 (N_935,In_801,In_802);
nor U936 (N_936,In_74,In_339);
and U937 (N_937,In_32,In_59);
nand U938 (N_938,In_603,In_879);
xor U939 (N_939,In_625,In_643);
and U940 (N_940,In_173,In_554);
and U941 (N_941,In_482,In_673);
nor U942 (N_942,In_66,In_152);
xor U943 (N_943,In_55,In_659);
or U944 (N_944,In_858,In_97);
nor U945 (N_945,In_78,In_640);
nand U946 (N_946,In_639,In_955);
nor U947 (N_947,In_307,In_775);
or U948 (N_948,In_607,In_412);
nor U949 (N_949,In_881,In_584);
nor U950 (N_950,In_724,In_432);
nand U951 (N_951,In_64,In_621);
nand U952 (N_952,In_634,In_852);
or U953 (N_953,In_996,In_358);
and U954 (N_954,In_786,In_145);
and U955 (N_955,In_175,In_411);
xnor U956 (N_956,In_506,In_139);
nor U957 (N_957,In_38,In_903);
xnor U958 (N_958,In_873,In_924);
xnor U959 (N_959,In_375,In_587);
and U960 (N_960,In_795,In_164);
nand U961 (N_961,In_651,In_579);
nand U962 (N_962,In_227,In_143);
and U963 (N_963,In_696,In_9);
and U964 (N_964,In_360,In_525);
xnor U965 (N_965,In_953,In_468);
xnor U966 (N_966,In_645,In_150);
xnor U967 (N_967,In_593,In_563);
and U968 (N_968,In_87,In_197);
or U969 (N_969,In_984,In_293);
nor U970 (N_970,In_858,In_723);
xor U971 (N_971,In_279,In_338);
and U972 (N_972,In_906,In_478);
nor U973 (N_973,In_283,In_410);
nand U974 (N_974,In_267,In_583);
nor U975 (N_975,In_61,In_69);
nand U976 (N_976,In_456,In_220);
nor U977 (N_977,In_276,In_724);
and U978 (N_978,In_495,In_832);
or U979 (N_979,In_516,In_676);
and U980 (N_980,In_293,In_314);
nor U981 (N_981,In_429,In_824);
and U982 (N_982,In_678,In_92);
xor U983 (N_983,In_541,In_99);
nor U984 (N_984,In_702,In_294);
xnor U985 (N_985,In_489,In_341);
nand U986 (N_986,In_31,In_823);
and U987 (N_987,In_230,In_488);
nor U988 (N_988,In_536,In_36);
nand U989 (N_989,In_160,In_461);
nor U990 (N_990,In_121,In_284);
xnor U991 (N_991,In_502,In_557);
and U992 (N_992,In_893,In_776);
nor U993 (N_993,In_861,In_719);
nand U994 (N_994,In_613,In_313);
or U995 (N_995,In_37,In_790);
nor U996 (N_996,In_750,In_794);
xnor U997 (N_997,In_861,In_886);
and U998 (N_998,In_459,In_344);
and U999 (N_999,In_131,In_754);
nor U1000 (N_1000,In_809,In_400);
nor U1001 (N_1001,In_531,In_632);
xor U1002 (N_1002,In_63,In_216);
nand U1003 (N_1003,In_213,In_952);
nand U1004 (N_1004,In_981,In_589);
or U1005 (N_1005,In_798,In_506);
or U1006 (N_1006,In_936,In_157);
xnor U1007 (N_1007,In_257,In_675);
and U1008 (N_1008,In_99,In_33);
nor U1009 (N_1009,In_809,In_435);
and U1010 (N_1010,In_575,In_345);
or U1011 (N_1011,In_463,In_579);
or U1012 (N_1012,In_752,In_16);
xnor U1013 (N_1013,In_11,In_854);
or U1014 (N_1014,In_109,In_814);
nor U1015 (N_1015,In_879,In_324);
nor U1016 (N_1016,In_564,In_384);
or U1017 (N_1017,In_134,In_202);
xor U1018 (N_1018,In_62,In_424);
nand U1019 (N_1019,In_679,In_241);
nand U1020 (N_1020,In_791,In_583);
and U1021 (N_1021,In_991,In_937);
nand U1022 (N_1022,In_34,In_509);
nand U1023 (N_1023,In_516,In_152);
xor U1024 (N_1024,In_3,In_911);
xor U1025 (N_1025,In_36,In_468);
nor U1026 (N_1026,In_422,In_303);
xnor U1027 (N_1027,In_731,In_447);
or U1028 (N_1028,In_342,In_288);
xnor U1029 (N_1029,In_11,In_396);
and U1030 (N_1030,In_912,In_540);
or U1031 (N_1031,In_648,In_535);
or U1032 (N_1032,In_84,In_530);
and U1033 (N_1033,In_116,In_663);
xnor U1034 (N_1034,In_577,In_444);
xnor U1035 (N_1035,In_206,In_806);
nor U1036 (N_1036,In_584,In_605);
xnor U1037 (N_1037,In_57,In_669);
and U1038 (N_1038,In_409,In_368);
or U1039 (N_1039,In_357,In_349);
nor U1040 (N_1040,In_803,In_910);
xor U1041 (N_1041,In_24,In_223);
nor U1042 (N_1042,In_546,In_620);
nor U1043 (N_1043,In_13,In_634);
and U1044 (N_1044,In_447,In_735);
or U1045 (N_1045,In_223,In_1);
xnor U1046 (N_1046,In_801,In_260);
or U1047 (N_1047,In_583,In_119);
xor U1048 (N_1048,In_725,In_399);
xnor U1049 (N_1049,In_31,In_370);
and U1050 (N_1050,In_975,In_143);
and U1051 (N_1051,In_243,In_779);
nand U1052 (N_1052,In_57,In_884);
or U1053 (N_1053,In_385,In_152);
or U1054 (N_1054,In_443,In_987);
nand U1055 (N_1055,In_751,In_814);
nand U1056 (N_1056,In_116,In_731);
nor U1057 (N_1057,In_33,In_655);
nor U1058 (N_1058,In_156,In_807);
and U1059 (N_1059,In_315,In_942);
and U1060 (N_1060,In_276,In_801);
xnor U1061 (N_1061,In_273,In_701);
or U1062 (N_1062,In_645,In_844);
nand U1063 (N_1063,In_98,In_348);
or U1064 (N_1064,In_716,In_709);
and U1065 (N_1065,In_785,In_458);
or U1066 (N_1066,In_901,In_730);
nor U1067 (N_1067,In_497,In_648);
or U1068 (N_1068,In_302,In_17);
xor U1069 (N_1069,In_191,In_11);
or U1070 (N_1070,In_570,In_181);
xor U1071 (N_1071,In_8,In_831);
or U1072 (N_1072,In_518,In_824);
nand U1073 (N_1073,In_95,In_776);
or U1074 (N_1074,In_17,In_590);
nor U1075 (N_1075,In_460,In_370);
and U1076 (N_1076,In_641,In_614);
xnor U1077 (N_1077,In_820,In_825);
or U1078 (N_1078,In_82,In_39);
xnor U1079 (N_1079,In_907,In_874);
or U1080 (N_1080,In_751,In_817);
nor U1081 (N_1081,In_178,In_585);
nor U1082 (N_1082,In_727,In_916);
xnor U1083 (N_1083,In_41,In_363);
nor U1084 (N_1084,In_885,In_575);
and U1085 (N_1085,In_53,In_599);
or U1086 (N_1086,In_640,In_109);
xnor U1087 (N_1087,In_663,In_942);
and U1088 (N_1088,In_649,In_917);
and U1089 (N_1089,In_619,In_845);
or U1090 (N_1090,In_750,In_771);
or U1091 (N_1091,In_39,In_739);
nand U1092 (N_1092,In_95,In_33);
xor U1093 (N_1093,In_552,In_959);
xnor U1094 (N_1094,In_26,In_892);
xor U1095 (N_1095,In_625,In_541);
nand U1096 (N_1096,In_305,In_198);
nand U1097 (N_1097,In_436,In_348);
xor U1098 (N_1098,In_315,In_156);
and U1099 (N_1099,In_693,In_745);
nor U1100 (N_1100,In_274,In_197);
and U1101 (N_1101,In_572,In_898);
nor U1102 (N_1102,In_911,In_838);
nor U1103 (N_1103,In_26,In_159);
or U1104 (N_1104,In_304,In_186);
and U1105 (N_1105,In_861,In_658);
nand U1106 (N_1106,In_638,In_38);
or U1107 (N_1107,In_71,In_336);
nor U1108 (N_1108,In_78,In_585);
and U1109 (N_1109,In_927,In_828);
nor U1110 (N_1110,In_780,In_499);
xor U1111 (N_1111,In_827,In_337);
nor U1112 (N_1112,In_489,In_318);
nand U1113 (N_1113,In_406,In_732);
xor U1114 (N_1114,In_786,In_550);
and U1115 (N_1115,In_106,In_534);
and U1116 (N_1116,In_723,In_426);
nor U1117 (N_1117,In_856,In_637);
or U1118 (N_1118,In_697,In_201);
nor U1119 (N_1119,In_92,In_236);
or U1120 (N_1120,In_613,In_175);
nor U1121 (N_1121,In_32,In_281);
nor U1122 (N_1122,In_25,In_287);
nor U1123 (N_1123,In_785,In_407);
nor U1124 (N_1124,In_521,In_31);
xnor U1125 (N_1125,In_161,In_602);
nand U1126 (N_1126,In_56,In_548);
nand U1127 (N_1127,In_924,In_711);
or U1128 (N_1128,In_558,In_476);
or U1129 (N_1129,In_460,In_58);
or U1130 (N_1130,In_457,In_287);
nand U1131 (N_1131,In_34,In_30);
nor U1132 (N_1132,In_432,In_354);
nand U1133 (N_1133,In_847,In_830);
and U1134 (N_1134,In_718,In_976);
xnor U1135 (N_1135,In_268,In_543);
xnor U1136 (N_1136,In_989,In_95);
nor U1137 (N_1137,In_912,In_816);
and U1138 (N_1138,In_894,In_302);
or U1139 (N_1139,In_6,In_712);
or U1140 (N_1140,In_881,In_506);
xnor U1141 (N_1141,In_765,In_259);
nand U1142 (N_1142,In_0,In_362);
and U1143 (N_1143,In_882,In_149);
or U1144 (N_1144,In_519,In_903);
nand U1145 (N_1145,In_600,In_509);
and U1146 (N_1146,In_377,In_306);
and U1147 (N_1147,In_662,In_797);
nor U1148 (N_1148,In_607,In_49);
nor U1149 (N_1149,In_304,In_550);
nand U1150 (N_1150,In_800,In_56);
and U1151 (N_1151,In_298,In_181);
and U1152 (N_1152,In_613,In_836);
xnor U1153 (N_1153,In_269,In_92);
xor U1154 (N_1154,In_328,In_964);
nor U1155 (N_1155,In_75,In_618);
nor U1156 (N_1156,In_940,In_67);
xor U1157 (N_1157,In_383,In_609);
and U1158 (N_1158,In_455,In_717);
and U1159 (N_1159,In_438,In_168);
and U1160 (N_1160,In_892,In_792);
and U1161 (N_1161,In_145,In_260);
xnor U1162 (N_1162,In_821,In_97);
nor U1163 (N_1163,In_213,In_409);
nor U1164 (N_1164,In_856,In_235);
xor U1165 (N_1165,In_470,In_28);
nor U1166 (N_1166,In_256,In_200);
nand U1167 (N_1167,In_442,In_677);
and U1168 (N_1168,In_238,In_555);
and U1169 (N_1169,In_649,In_138);
nand U1170 (N_1170,In_738,In_952);
nand U1171 (N_1171,In_425,In_485);
and U1172 (N_1172,In_996,In_545);
and U1173 (N_1173,In_101,In_877);
and U1174 (N_1174,In_64,In_90);
or U1175 (N_1175,In_678,In_176);
xnor U1176 (N_1176,In_790,In_84);
nand U1177 (N_1177,In_381,In_329);
xnor U1178 (N_1178,In_925,In_83);
nor U1179 (N_1179,In_570,In_846);
xnor U1180 (N_1180,In_139,In_371);
nand U1181 (N_1181,In_455,In_976);
nand U1182 (N_1182,In_894,In_661);
and U1183 (N_1183,In_58,In_953);
nor U1184 (N_1184,In_198,In_224);
or U1185 (N_1185,In_56,In_216);
nor U1186 (N_1186,In_655,In_969);
or U1187 (N_1187,In_107,In_580);
and U1188 (N_1188,In_396,In_971);
nor U1189 (N_1189,In_921,In_806);
xor U1190 (N_1190,In_670,In_542);
nor U1191 (N_1191,In_604,In_464);
and U1192 (N_1192,In_477,In_968);
nor U1193 (N_1193,In_456,In_904);
nand U1194 (N_1194,In_861,In_396);
and U1195 (N_1195,In_460,In_455);
nand U1196 (N_1196,In_558,In_707);
xor U1197 (N_1197,In_892,In_772);
and U1198 (N_1198,In_193,In_639);
or U1199 (N_1199,In_262,In_368);
nand U1200 (N_1200,In_356,In_494);
and U1201 (N_1201,In_504,In_490);
xor U1202 (N_1202,In_220,In_177);
xnor U1203 (N_1203,In_392,In_884);
and U1204 (N_1204,In_148,In_236);
or U1205 (N_1205,In_62,In_297);
nor U1206 (N_1206,In_831,In_778);
xor U1207 (N_1207,In_729,In_259);
or U1208 (N_1208,In_160,In_966);
xor U1209 (N_1209,In_773,In_661);
nand U1210 (N_1210,In_416,In_861);
or U1211 (N_1211,In_120,In_358);
and U1212 (N_1212,In_917,In_290);
and U1213 (N_1213,In_599,In_20);
or U1214 (N_1214,In_190,In_688);
xnor U1215 (N_1215,In_659,In_69);
xnor U1216 (N_1216,In_180,In_474);
xor U1217 (N_1217,In_370,In_983);
nand U1218 (N_1218,In_49,In_528);
xnor U1219 (N_1219,In_961,In_360);
xnor U1220 (N_1220,In_952,In_634);
nand U1221 (N_1221,In_775,In_793);
nand U1222 (N_1222,In_929,In_19);
nor U1223 (N_1223,In_793,In_952);
and U1224 (N_1224,In_247,In_854);
xor U1225 (N_1225,In_839,In_421);
nand U1226 (N_1226,In_943,In_273);
and U1227 (N_1227,In_898,In_306);
nand U1228 (N_1228,In_892,In_71);
nor U1229 (N_1229,In_722,In_458);
nor U1230 (N_1230,In_696,In_590);
nand U1231 (N_1231,In_65,In_237);
xnor U1232 (N_1232,In_159,In_413);
or U1233 (N_1233,In_473,In_772);
nand U1234 (N_1234,In_440,In_986);
or U1235 (N_1235,In_826,In_576);
nand U1236 (N_1236,In_602,In_370);
nand U1237 (N_1237,In_111,In_469);
nand U1238 (N_1238,In_623,In_525);
nor U1239 (N_1239,In_111,In_141);
and U1240 (N_1240,In_965,In_559);
nand U1241 (N_1241,In_408,In_491);
and U1242 (N_1242,In_278,In_361);
nor U1243 (N_1243,In_819,In_959);
nor U1244 (N_1244,In_213,In_202);
xnor U1245 (N_1245,In_307,In_370);
xor U1246 (N_1246,In_679,In_817);
nor U1247 (N_1247,In_0,In_433);
xor U1248 (N_1248,In_440,In_447);
nand U1249 (N_1249,In_975,In_279);
xor U1250 (N_1250,In_274,In_629);
and U1251 (N_1251,In_176,In_8);
or U1252 (N_1252,In_466,In_159);
nand U1253 (N_1253,In_767,In_837);
and U1254 (N_1254,In_595,In_982);
nor U1255 (N_1255,In_627,In_599);
nand U1256 (N_1256,In_348,In_301);
nor U1257 (N_1257,In_218,In_577);
or U1258 (N_1258,In_652,In_237);
nand U1259 (N_1259,In_23,In_755);
nor U1260 (N_1260,In_324,In_2);
and U1261 (N_1261,In_356,In_257);
and U1262 (N_1262,In_494,In_79);
or U1263 (N_1263,In_756,In_175);
nand U1264 (N_1264,In_524,In_817);
nor U1265 (N_1265,In_211,In_657);
nor U1266 (N_1266,In_79,In_699);
or U1267 (N_1267,In_795,In_187);
xor U1268 (N_1268,In_450,In_660);
nor U1269 (N_1269,In_549,In_129);
nor U1270 (N_1270,In_334,In_901);
nor U1271 (N_1271,In_575,In_948);
nor U1272 (N_1272,In_75,In_213);
and U1273 (N_1273,In_323,In_954);
and U1274 (N_1274,In_780,In_284);
or U1275 (N_1275,In_834,In_628);
nor U1276 (N_1276,In_229,In_270);
or U1277 (N_1277,In_573,In_405);
and U1278 (N_1278,In_445,In_698);
nor U1279 (N_1279,In_771,In_506);
nor U1280 (N_1280,In_583,In_934);
nand U1281 (N_1281,In_874,In_152);
or U1282 (N_1282,In_443,In_975);
and U1283 (N_1283,In_52,In_903);
nand U1284 (N_1284,In_509,In_128);
or U1285 (N_1285,In_815,In_255);
or U1286 (N_1286,In_228,In_181);
xor U1287 (N_1287,In_454,In_549);
nand U1288 (N_1288,In_712,In_998);
and U1289 (N_1289,In_925,In_793);
nor U1290 (N_1290,In_158,In_463);
nor U1291 (N_1291,In_599,In_670);
nand U1292 (N_1292,In_773,In_814);
or U1293 (N_1293,In_43,In_997);
and U1294 (N_1294,In_778,In_517);
and U1295 (N_1295,In_700,In_239);
nor U1296 (N_1296,In_417,In_478);
xnor U1297 (N_1297,In_695,In_913);
or U1298 (N_1298,In_799,In_645);
nand U1299 (N_1299,In_653,In_931);
nand U1300 (N_1300,In_916,In_919);
and U1301 (N_1301,In_623,In_719);
xnor U1302 (N_1302,In_343,In_119);
xnor U1303 (N_1303,In_508,In_758);
xor U1304 (N_1304,In_194,In_881);
or U1305 (N_1305,In_713,In_698);
nor U1306 (N_1306,In_998,In_316);
nor U1307 (N_1307,In_814,In_375);
and U1308 (N_1308,In_420,In_74);
and U1309 (N_1309,In_598,In_790);
xnor U1310 (N_1310,In_318,In_538);
nand U1311 (N_1311,In_108,In_980);
or U1312 (N_1312,In_353,In_667);
and U1313 (N_1313,In_705,In_19);
and U1314 (N_1314,In_172,In_851);
or U1315 (N_1315,In_39,In_675);
xor U1316 (N_1316,In_784,In_84);
xor U1317 (N_1317,In_613,In_634);
and U1318 (N_1318,In_176,In_82);
or U1319 (N_1319,In_238,In_672);
xnor U1320 (N_1320,In_8,In_129);
xnor U1321 (N_1321,In_389,In_376);
nor U1322 (N_1322,In_472,In_223);
nor U1323 (N_1323,In_880,In_130);
and U1324 (N_1324,In_376,In_944);
and U1325 (N_1325,In_423,In_817);
nor U1326 (N_1326,In_32,In_504);
nor U1327 (N_1327,In_472,In_106);
nor U1328 (N_1328,In_256,In_942);
nor U1329 (N_1329,In_686,In_149);
nand U1330 (N_1330,In_503,In_246);
and U1331 (N_1331,In_933,In_95);
nand U1332 (N_1332,In_441,In_830);
xnor U1333 (N_1333,In_114,In_57);
or U1334 (N_1334,In_815,In_819);
and U1335 (N_1335,In_35,In_887);
and U1336 (N_1336,In_56,In_606);
nand U1337 (N_1337,In_796,In_506);
xor U1338 (N_1338,In_39,In_98);
or U1339 (N_1339,In_937,In_782);
nor U1340 (N_1340,In_905,In_922);
or U1341 (N_1341,In_620,In_690);
or U1342 (N_1342,In_972,In_947);
and U1343 (N_1343,In_304,In_242);
nand U1344 (N_1344,In_21,In_87);
xnor U1345 (N_1345,In_878,In_731);
or U1346 (N_1346,In_745,In_113);
nor U1347 (N_1347,In_852,In_744);
and U1348 (N_1348,In_392,In_57);
xor U1349 (N_1349,In_501,In_687);
nor U1350 (N_1350,In_563,In_453);
and U1351 (N_1351,In_984,In_796);
and U1352 (N_1352,In_722,In_916);
or U1353 (N_1353,In_484,In_143);
or U1354 (N_1354,In_884,In_330);
nor U1355 (N_1355,In_562,In_347);
and U1356 (N_1356,In_156,In_223);
and U1357 (N_1357,In_608,In_832);
and U1358 (N_1358,In_544,In_73);
xnor U1359 (N_1359,In_114,In_416);
nor U1360 (N_1360,In_75,In_973);
and U1361 (N_1361,In_865,In_523);
nand U1362 (N_1362,In_510,In_747);
nand U1363 (N_1363,In_33,In_46);
xnor U1364 (N_1364,In_668,In_328);
nand U1365 (N_1365,In_62,In_933);
nor U1366 (N_1366,In_899,In_322);
nand U1367 (N_1367,In_273,In_104);
nand U1368 (N_1368,In_16,In_301);
and U1369 (N_1369,In_89,In_981);
and U1370 (N_1370,In_633,In_350);
or U1371 (N_1371,In_912,In_579);
and U1372 (N_1372,In_32,In_741);
or U1373 (N_1373,In_298,In_494);
nand U1374 (N_1374,In_739,In_131);
xor U1375 (N_1375,In_527,In_233);
nand U1376 (N_1376,In_969,In_676);
nor U1377 (N_1377,In_747,In_429);
and U1378 (N_1378,In_958,In_93);
or U1379 (N_1379,In_66,In_839);
xor U1380 (N_1380,In_543,In_664);
or U1381 (N_1381,In_220,In_830);
or U1382 (N_1382,In_236,In_484);
nand U1383 (N_1383,In_169,In_784);
xnor U1384 (N_1384,In_480,In_368);
nand U1385 (N_1385,In_416,In_153);
and U1386 (N_1386,In_508,In_869);
or U1387 (N_1387,In_750,In_438);
nor U1388 (N_1388,In_401,In_746);
nand U1389 (N_1389,In_366,In_957);
and U1390 (N_1390,In_62,In_373);
and U1391 (N_1391,In_728,In_500);
and U1392 (N_1392,In_280,In_293);
and U1393 (N_1393,In_135,In_727);
xor U1394 (N_1394,In_814,In_258);
and U1395 (N_1395,In_226,In_113);
or U1396 (N_1396,In_832,In_989);
nor U1397 (N_1397,In_316,In_489);
or U1398 (N_1398,In_210,In_420);
xor U1399 (N_1399,In_583,In_970);
xor U1400 (N_1400,In_64,In_242);
nand U1401 (N_1401,In_839,In_996);
nor U1402 (N_1402,In_474,In_586);
xnor U1403 (N_1403,In_796,In_982);
or U1404 (N_1404,In_614,In_405);
or U1405 (N_1405,In_521,In_144);
nor U1406 (N_1406,In_632,In_237);
nand U1407 (N_1407,In_49,In_989);
and U1408 (N_1408,In_137,In_790);
nor U1409 (N_1409,In_130,In_934);
or U1410 (N_1410,In_428,In_838);
xnor U1411 (N_1411,In_56,In_646);
nand U1412 (N_1412,In_182,In_566);
nor U1413 (N_1413,In_13,In_715);
and U1414 (N_1414,In_33,In_442);
or U1415 (N_1415,In_266,In_796);
nand U1416 (N_1416,In_951,In_605);
nor U1417 (N_1417,In_403,In_97);
and U1418 (N_1418,In_519,In_495);
nor U1419 (N_1419,In_228,In_11);
or U1420 (N_1420,In_795,In_591);
or U1421 (N_1421,In_343,In_582);
nand U1422 (N_1422,In_161,In_428);
xnor U1423 (N_1423,In_68,In_184);
nor U1424 (N_1424,In_706,In_376);
or U1425 (N_1425,In_719,In_563);
xnor U1426 (N_1426,In_746,In_22);
xnor U1427 (N_1427,In_768,In_342);
nand U1428 (N_1428,In_472,In_234);
xor U1429 (N_1429,In_904,In_120);
or U1430 (N_1430,In_171,In_316);
or U1431 (N_1431,In_940,In_922);
nor U1432 (N_1432,In_402,In_433);
nor U1433 (N_1433,In_822,In_110);
nor U1434 (N_1434,In_212,In_755);
nor U1435 (N_1435,In_534,In_412);
and U1436 (N_1436,In_436,In_132);
and U1437 (N_1437,In_728,In_732);
nand U1438 (N_1438,In_229,In_41);
nand U1439 (N_1439,In_630,In_682);
xor U1440 (N_1440,In_64,In_58);
or U1441 (N_1441,In_47,In_319);
xnor U1442 (N_1442,In_618,In_136);
and U1443 (N_1443,In_280,In_655);
xor U1444 (N_1444,In_933,In_420);
xor U1445 (N_1445,In_171,In_709);
or U1446 (N_1446,In_639,In_907);
nand U1447 (N_1447,In_401,In_86);
or U1448 (N_1448,In_804,In_448);
and U1449 (N_1449,In_749,In_744);
or U1450 (N_1450,In_557,In_29);
or U1451 (N_1451,In_209,In_914);
nand U1452 (N_1452,In_967,In_335);
or U1453 (N_1453,In_943,In_225);
nand U1454 (N_1454,In_280,In_343);
or U1455 (N_1455,In_766,In_49);
or U1456 (N_1456,In_429,In_779);
and U1457 (N_1457,In_100,In_846);
xnor U1458 (N_1458,In_636,In_97);
xor U1459 (N_1459,In_863,In_326);
nand U1460 (N_1460,In_443,In_584);
nand U1461 (N_1461,In_730,In_991);
or U1462 (N_1462,In_115,In_710);
xor U1463 (N_1463,In_726,In_396);
nor U1464 (N_1464,In_664,In_418);
nand U1465 (N_1465,In_187,In_678);
and U1466 (N_1466,In_931,In_832);
and U1467 (N_1467,In_162,In_763);
nand U1468 (N_1468,In_498,In_607);
xor U1469 (N_1469,In_120,In_934);
nand U1470 (N_1470,In_494,In_613);
and U1471 (N_1471,In_201,In_379);
nand U1472 (N_1472,In_175,In_453);
and U1473 (N_1473,In_620,In_990);
nor U1474 (N_1474,In_381,In_80);
nor U1475 (N_1475,In_531,In_688);
nor U1476 (N_1476,In_933,In_626);
nor U1477 (N_1477,In_522,In_868);
nand U1478 (N_1478,In_883,In_829);
nand U1479 (N_1479,In_21,In_557);
xnor U1480 (N_1480,In_399,In_656);
xnor U1481 (N_1481,In_374,In_850);
nand U1482 (N_1482,In_186,In_157);
or U1483 (N_1483,In_604,In_945);
and U1484 (N_1484,In_817,In_205);
and U1485 (N_1485,In_963,In_613);
xor U1486 (N_1486,In_983,In_500);
nor U1487 (N_1487,In_94,In_995);
and U1488 (N_1488,In_726,In_458);
nor U1489 (N_1489,In_695,In_613);
or U1490 (N_1490,In_802,In_11);
nand U1491 (N_1491,In_7,In_331);
nand U1492 (N_1492,In_736,In_531);
nand U1493 (N_1493,In_872,In_23);
nand U1494 (N_1494,In_168,In_345);
nor U1495 (N_1495,In_590,In_38);
and U1496 (N_1496,In_37,In_886);
nor U1497 (N_1497,In_401,In_741);
and U1498 (N_1498,In_7,In_803);
xor U1499 (N_1499,In_962,In_985);
nand U1500 (N_1500,In_303,In_130);
xnor U1501 (N_1501,In_98,In_539);
nand U1502 (N_1502,In_735,In_585);
nand U1503 (N_1503,In_427,In_621);
nand U1504 (N_1504,In_158,In_584);
or U1505 (N_1505,In_133,In_420);
xor U1506 (N_1506,In_806,In_892);
nor U1507 (N_1507,In_420,In_633);
or U1508 (N_1508,In_443,In_444);
nand U1509 (N_1509,In_933,In_211);
nor U1510 (N_1510,In_364,In_74);
nand U1511 (N_1511,In_664,In_504);
or U1512 (N_1512,In_940,In_468);
nor U1513 (N_1513,In_938,In_174);
or U1514 (N_1514,In_962,In_859);
nand U1515 (N_1515,In_551,In_40);
xor U1516 (N_1516,In_67,In_328);
or U1517 (N_1517,In_178,In_349);
nand U1518 (N_1518,In_946,In_756);
xnor U1519 (N_1519,In_122,In_783);
xor U1520 (N_1520,In_489,In_333);
or U1521 (N_1521,In_269,In_406);
nor U1522 (N_1522,In_872,In_985);
and U1523 (N_1523,In_101,In_972);
nand U1524 (N_1524,In_302,In_857);
or U1525 (N_1525,In_387,In_495);
xnor U1526 (N_1526,In_472,In_898);
or U1527 (N_1527,In_770,In_587);
and U1528 (N_1528,In_173,In_65);
and U1529 (N_1529,In_855,In_794);
or U1530 (N_1530,In_23,In_89);
xnor U1531 (N_1531,In_566,In_707);
nand U1532 (N_1532,In_757,In_621);
nand U1533 (N_1533,In_733,In_130);
or U1534 (N_1534,In_88,In_599);
or U1535 (N_1535,In_906,In_711);
or U1536 (N_1536,In_314,In_254);
or U1537 (N_1537,In_319,In_558);
and U1538 (N_1538,In_471,In_151);
nor U1539 (N_1539,In_958,In_339);
and U1540 (N_1540,In_518,In_181);
nand U1541 (N_1541,In_119,In_168);
nor U1542 (N_1542,In_318,In_601);
nand U1543 (N_1543,In_207,In_37);
nor U1544 (N_1544,In_5,In_285);
or U1545 (N_1545,In_424,In_236);
nor U1546 (N_1546,In_631,In_405);
nand U1547 (N_1547,In_841,In_936);
xor U1548 (N_1548,In_873,In_951);
nor U1549 (N_1549,In_152,In_75);
xnor U1550 (N_1550,In_159,In_0);
xor U1551 (N_1551,In_6,In_678);
nand U1552 (N_1552,In_275,In_505);
nor U1553 (N_1553,In_539,In_52);
nor U1554 (N_1554,In_648,In_852);
and U1555 (N_1555,In_693,In_349);
nand U1556 (N_1556,In_908,In_929);
xnor U1557 (N_1557,In_126,In_192);
or U1558 (N_1558,In_707,In_212);
nand U1559 (N_1559,In_694,In_392);
nand U1560 (N_1560,In_753,In_417);
nor U1561 (N_1561,In_735,In_496);
and U1562 (N_1562,In_5,In_443);
nor U1563 (N_1563,In_668,In_274);
or U1564 (N_1564,In_636,In_682);
nor U1565 (N_1565,In_689,In_941);
xor U1566 (N_1566,In_197,In_568);
or U1567 (N_1567,In_386,In_322);
or U1568 (N_1568,In_119,In_34);
and U1569 (N_1569,In_828,In_237);
nor U1570 (N_1570,In_229,In_733);
nand U1571 (N_1571,In_615,In_590);
nor U1572 (N_1572,In_168,In_103);
nor U1573 (N_1573,In_347,In_983);
and U1574 (N_1574,In_208,In_543);
xor U1575 (N_1575,In_984,In_527);
or U1576 (N_1576,In_637,In_851);
xor U1577 (N_1577,In_497,In_397);
nor U1578 (N_1578,In_125,In_16);
xnor U1579 (N_1579,In_600,In_323);
xnor U1580 (N_1580,In_34,In_668);
xnor U1581 (N_1581,In_73,In_302);
and U1582 (N_1582,In_749,In_359);
xor U1583 (N_1583,In_490,In_723);
xor U1584 (N_1584,In_461,In_876);
nand U1585 (N_1585,In_522,In_132);
or U1586 (N_1586,In_338,In_403);
xnor U1587 (N_1587,In_187,In_846);
and U1588 (N_1588,In_369,In_707);
nor U1589 (N_1589,In_985,In_981);
nand U1590 (N_1590,In_330,In_584);
xor U1591 (N_1591,In_403,In_447);
and U1592 (N_1592,In_9,In_408);
nand U1593 (N_1593,In_349,In_3);
nand U1594 (N_1594,In_199,In_478);
nor U1595 (N_1595,In_353,In_6);
nand U1596 (N_1596,In_279,In_219);
or U1597 (N_1597,In_197,In_253);
or U1598 (N_1598,In_560,In_603);
xor U1599 (N_1599,In_32,In_288);
or U1600 (N_1600,In_985,In_820);
nor U1601 (N_1601,In_282,In_397);
nor U1602 (N_1602,In_928,In_55);
and U1603 (N_1603,In_547,In_715);
or U1604 (N_1604,In_132,In_729);
nand U1605 (N_1605,In_346,In_626);
nand U1606 (N_1606,In_476,In_832);
nand U1607 (N_1607,In_720,In_66);
nor U1608 (N_1608,In_359,In_781);
and U1609 (N_1609,In_609,In_283);
or U1610 (N_1610,In_807,In_836);
or U1611 (N_1611,In_664,In_641);
nand U1612 (N_1612,In_904,In_289);
and U1613 (N_1613,In_359,In_28);
nor U1614 (N_1614,In_284,In_649);
nor U1615 (N_1615,In_94,In_465);
nor U1616 (N_1616,In_490,In_755);
or U1617 (N_1617,In_220,In_968);
and U1618 (N_1618,In_723,In_108);
or U1619 (N_1619,In_996,In_18);
or U1620 (N_1620,In_573,In_959);
nand U1621 (N_1621,In_461,In_637);
and U1622 (N_1622,In_359,In_751);
xor U1623 (N_1623,In_885,In_201);
and U1624 (N_1624,In_561,In_118);
and U1625 (N_1625,In_996,In_385);
and U1626 (N_1626,In_457,In_841);
or U1627 (N_1627,In_835,In_746);
nor U1628 (N_1628,In_994,In_25);
and U1629 (N_1629,In_585,In_441);
nor U1630 (N_1630,In_538,In_616);
nor U1631 (N_1631,In_82,In_430);
nor U1632 (N_1632,In_339,In_870);
or U1633 (N_1633,In_367,In_51);
nor U1634 (N_1634,In_865,In_590);
xor U1635 (N_1635,In_588,In_711);
xnor U1636 (N_1636,In_937,In_545);
or U1637 (N_1637,In_195,In_395);
and U1638 (N_1638,In_715,In_53);
nor U1639 (N_1639,In_938,In_531);
xnor U1640 (N_1640,In_793,In_800);
and U1641 (N_1641,In_322,In_458);
or U1642 (N_1642,In_282,In_561);
nand U1643 (N_1643,In_571,In_354);
nand U1644 (N_1644,In_278,In_863);
and U1645 (N_1645,In_397,In_628);
nand U1646 (N_1646,In_239,In_153);
nor U1647 (N_1647,In_66,In_408);
xnor U1648 (N_1648,In_0,In_31);
nor U1649 (N_1649,In_726,In_169);
xor U1650 (N_1650,In_567,In_879);
and U1651 (N_1651,In_188,In_793);
or U1652 (N_1652,In_344,In_242);
or U1653 (N_1653,In_110,In_40);
nand U1654 (N_1654,In_256,In_46);
or U1655 (N_1655,In_714,In_977);
xor U1656 (N_1656,In_759,In_293);
nor U1657 (N_1657,In_929,In_16);
nand U1658 (N_1658,In_587,In_455);
nor U1659 (N_1659,In_795,In_330);
and U1660 (N_1660,In_362,In_507);
nor U1661 (N_1661,In_985,In_564);
nor U1662 (N_1662,In_436,In_553);
or U1663 (N_1663,In_639,In_659);
and U1664 (N_1664,In_120,In_235);
nor U1665 (N_1665,In_601,In_817);
nand U1666 (N_1666,In_967,In_612);
and U1667 (N_1667,In_96,In_61);
or U1668 (N_1668,In_599,In_28);
or U1669 (N_1669,In_712,In_173);
nand U1670 (N_1670,In_647,In_433);
and U1671 (N_1671,In_432,In_114);
xnor U1672 (N_1672,In_260,In_403);
nand U1673 (N_1673,In_725,In_560);
nand U1674 (N_1674,In_91,In_853);
nand U1675 (N_1675,In_374,In_187);
xor U1676 (N_1676,In_363,In_629);
or U1677 (N_1677,In_154,In_484);
or U1678 (N_1678,In_387,In_428);
and U1679 (N_1679,In_6,In_578);
or U1680 (N_1680,In_732,In_750);
nor U1681 (N_1681,In_495,In_148);
nor U1682 (N_1682,In_416,In_753);
nand U1683 (N_1683,In_876,In_974);
or U1684 (N_1684,In_788,In_371);
xor U1685 (N_1685,In_163,In_207);
nand U1686 (N_1686,In_614,In_897);
and U1687 (N_1687,In_514,In_40);
or U1688 (N_1688,In_238,In_588);
or U1689 (N_1689,In_85,In_835);
and U1690 (N_1690,In_748,In_418);
nand U1691 (N_1691,In_997,In_570);
xor U1692 (N_1692,In_686,In_70);
and U1693 (N_1693,In_477,In_445);
nand U1694 (N_1694,In_425,In_65);
and U1695 (N_1695,In_476,In_309);
xnor U1696 (N_1696,In_107,In_811);
and U1697 (N_1697,In_739,In_99);
nor U1698 (N_1698,In_573,In_785);
xor U1699 (N_1699,In_93,In_905);
xor U1700 (N_1700,In_491,In_808);
nor U1701 (N_1701,In_140,In_684);
nand U1702 (N_1702,In_549,In_113);
nand U1703 (N_1703,In_901,In_947);
nor U1704 (N_1704,In_297,In_957);
or U1705 (N_1705,In_921,In_589);
nor U1706 (N_1706,In_961,In_108);
xor U1707 (N_1707,In_656,In_815);
or U1708 (N_1708,In_61,In_600);
nor U1709 (N_1709,In_236,In_907);
nand U1710 (N_1710,In_81,In_780);
and U1711 (N_1711,In_656,In_765);
nand U1712 (N_1712,In_762,In_564);
xnor U1713 (N_1713,In_427,In_848);
nand U1714 (N_1714,In_654,In_252);
nor U1715 (N_1715,In_272,In_123);
or U1716 (N_1716,In_202,In_319);
nand U1717 (N_1717,In_326,In_969);
or U1718 (N_1718,In_113,In_311);
xor U1719 (N_1719,In_787,In_640);
and U1720 (N_1720,In_501,In_593);
xnor U1721 (N_1721,In_434,In_697);
xor U1722 (N_1722,In_42,In_569);
xnor U1723 (N_1723,In_762,In_507);
xor U1724 (N_1724,In_515,In_841);
xnor U1725 (N_1725,In_407,In_62);
or U1726 (N_1726,In_66,In_813);
nor U1727 (N_1727,In_987,In_408);
nor U1728 (N_1728,In_533,In_320);
nor U1729 (N_1729,In_556,In_743);
and U1730 (N_1730,In_942,In_50);
and U1731 (N_1731,In_657,In_707);
and U1732 (N_1732,In_461,In_415);
xor U1733 (N_1733,In_349,In_290);
and U1734 (N_1734,In_136,In_600);
and U1735 (N_1735,In_446,In_79);
xor U1736 (N_1736,In_375,In_448);
or U1737 (N_1737,In_994,In_621);
xor U1738 (N_1738,In_335,In_769);
and U1739 (N_1739,In_923,In_839);
and U1740 (N_1740,In_215,In_171);
nand U1741 (N_1741,In_169,In_706);
nor U1742 (N_1742,In_122,In_327);
nand U1743 (N_1743,In_440,In_563);
nand U1744 (N_1744,In_825,In_668);
nand U1745 (N_1745,In_685,In_968);
nor U1746 (N_1746,In_941,In_243);
nor U1747 (N_1747,In_87,In_210);
and U1748 (N_1748,In_73,In_667);
and U1749 (N_1749,In_650,In_696);
or U1750 (N_1750,In_879,In_158);
nand U1751 (N_1751,In_569,In_471);
or U1752 (N_1752,In_610,In_978);
nand U1753 (N_1753,In_765,In_238);
nor U1754 (N_1754,In_189,In_970);
or U1755 (N_1755,In_349,In_303);
or U1756 (N_1756,In_195,In_385);
nand U1757 (N_1757,In_171,In_636);
nand U1758 (N_1758,In_871,In_983);
and U1759 (N_1759,In_950,In_852);
nor U1760 (N_1760,In_550,In_898);
xor U1761 (N_1761,In_890,In_719);
xnor U1762 (N_1762,In_771,In_947);
and U1763 (N_1763,In_622,In_196);
nor U1764 (N_1764,In_136,In_893);
xor U1765 (N_1765,In_597,In_569);
nand U1766 (N_1766,In_324,In_564);
nand U1767 (N_1767,In_203,In_700);
or U1768 (N_1768,In_201,In_681);
or U1769 (N_1769,In_623,In_189);
and U1770 (N_1770,In_640,In_146);
nor U1771 (N_1771,In_927,In_516);
nand U1772 (N_1772,In_371,In_752);
and U1773 (N_1773,In_502,In_96);
nor U1774 (N_1774,In_495,In_502);
xor U1775 (N_1775,In_777,In_177);
nand U1776 (N_1776,In_352,In_324);
xor U1777 (N_1777,In_735,In_261);
nand U1778 (N_1778,In_419,In_948);
or U1779 (N_1779,In_210,In_647);
nand U1780 (N_1780,In_758,In_206);
and U1781 (N_1781,In_514,In_651);
nor U1782 (N_1782,In_339,In_686);
xnor U1783 (N_1783,In_695,In_904);
or U1784 (N_1784,In_258,In_52);
nand U1785 (N_1785,In_342,In_729);
xor U1786 (N_1786,In_596,In_462);
nor U1787 (N_1787,In_662,In_815);
or U1788 (N_1788,In_226,In_110);
xor U1789 (N_1789,In_936,In_443);
nor U1790 (N_1790,In_277,In_693);
xnor U1791 (N_1791,In_890,In_359);
or U1792 (N_1792,In_149,In_327);
nor U1793 (N_1793,In_598,In_880);
nand U1794 (N_1794,In_626,In_613);
nand U1795 (N_1795,In_301,In_654);
nand U1796 (N_1796,In_178,In_950);
or U1797 (N_1797,In_503,In_324);
nor U1798 (N_1798,In_159,In_344);
nor U1799 (N_1799,In_722,In_17);
xnor U1800 (N_1800,In_418,In_9);
nand U1801 (N_1801,In_974,In_692);
xor U1802 (N_1802,In_849,In_62);
xnor U1803 (N_1803,In_472,In_257);
and U1804 (N_1804,In_34,In_406);
or U1805 (N_1805,In_189,In_71);
xor U1806 (N_1806,In_143,In_938);
xnor U1807 (N_1807,In_899,In_148);
and U1808 (N_1808,In_456,In_478);
nand U1809 (N_1809,In_310,In_583);
or U1810 (N_1810,In_246,In_873);
nor U1811 (N_1811,In_685,In_790);
or U1812 (N_1812,In_92,In_158);
or U1813 (N_1813,In_500,In_3);
or U1814 (N_1814,In_343,In_181);
or U1815 (N_1815,In_341,In_702);
and U1816 (N_1816,In_668,In_234);
and U1817 (N_1817,In_579,In_134);
nand U1818 (N_1818,In_604,In_344);
and U1819 (N_1819,In_243,In_167);
nand U1820 (N_1820,In_566,In_989);
and U1821 (N_1821,In_453,In_621);
nand U1822 (N_1822,In_249,In_930);
nand U1823 (N_1823,In_910,In_283);
nand U1824 (N_1824,In_708,In_445);
and U1825 (N_1825,In_972,In_47);
xnor U1826 (N_1826,In_151,In_812);
nor U1827 (N_1827,In_381,In_179);
nand U1828 (N_1828,In_991,In_235);
or U1829 (N_1829,In_918,In_350);
or U1830 (N_1830,In_208,In_868);
xnor U1831 (N_1831,In_774,In_62);
or U1832 (N_1832,In_208,In_639);
nand U1833 (N_1833,In_736,In_633);
xor U1834 (N_1834,In_904,In_468);
and U1835 (N_1835,In_157,In_995);
or U1836 (N_1836,In_801,In_923);
nor U1837 (N_1837,In_321,In_868);
nor U1838 (N_1838,In_834,In_699);
nor U1839 (N_1839,In_237,In_617);
nor U1840 (N_1840,In_911,In_540);
xnor U1841 (N_1841,In_359,In_853);
or U1842 (N_1842,In_226,In_777);
nand U1843 (N_1843,In_287,In_32);
nor U1844 (N_1844,In_727,In_777);
xnor U1845 (N_1845,In_199,In_193);
or U1846 (N_1846,In_423,In_395);
or U1847 (N_1847,In_974,In_965);
nand U1848 (N_1848,In_586,In_69);
and U1849 (N_1849,In_934,In_265);
or U1850 (N_1850,In_313,In_132);
xnor U1851 (N_1851,In_122,In_633);
nand U1852 (N_1852,In_872,In_785);
xnor U1853 (N_1853,In_449,In_379);
nand U1854 (N_1854,In_882,In_700);
xnor U1855 (N_1855,In_947,In_978);
and U1856 (N_1856,In_905,In_26);
xnor U1857 (N_1857,In_854,In_675);
or U1858 (N_1858,In_784,In_649);
or U1859 (N_1859,In_278,In_552);
xor U1860 (N_1860,In_143,In_457);
and U1861 (N_1861,In_429,In_603);
and U1862 (N_1862,In_936,In_124);
or U1863 (N_1863,In_386,In_661);
xnor U1864 (N_1864,In_714,In_318);
or U1865 (N_1865,In_178,In_478);
xor U1866 (N_1866,In_496,In_589);
or U1867 (N_1867,In_846,In_838);
or U1868 (N_1868,In_627,In_640);
nand U1869 (N_1869,In_682,In_522);
and U1870 (N_1870,In_996,In_625);
nand U1871 (N_1871,In_590,In_562);
or U1872 (N_1872,In_773,In_442);
nor U1873 (N_1873,In_550,In_465);
and U1874 (N_1874,In_211,In_892);
or U1875 (N_1875,In_113,In_379);
xnor U1876 (N_1876,In_821,In_586);
nor U1877 (N_1877,In_562,In_301);
nand U1878 (N_1878,In_920,In_690);
nor U1879 (N_1879,In_582,In_223);
nor U1880 (N_1880,In_510,In_4);
or U1881 (N_1881,In_837,In_877);
and U1882 (N_1882,In_431,In_885);
nor U1883 (N_1883,In_909,In_168);
xnor U1884 (N_1884,In_419,In_296);
nor U1885 (N_1885,In_113,In_880);
and U1886 (N_1886,In_762,In_429);
nor U1887 (N_1887,In_823,In_998);
or U1888 (N_1888,In_225,In_573);
and U1889 (N_1889,In_777,In_81);
nand U1890 (N_1890,In_650,In_305);
or U1891 (N_1891,In_389,In_991);
xor U1892 (N_1892,In_412,In_834);
xnor U1893 (N_1893,In_594,In_986);
nor U1894 (N_1894,In_985,In_75);
and U1895 (N_1895,In_723,In_836);
xor U1896 (N_1896,In_853,In_745);
nor U1897 (N_1897,In_644,In_724);
xnor U1898 (N_1898,In_769,In_489);
or U1899 (N_1899,In_657,In_711);
or U1900 (N_1900,In_69,In_959);
and U1901 (N_1901,In_337,In_534);
xnor U1902 (N_1902,In_307,In_375);
nand U1903 (N_1903,In_815,In_479);
nor U1904 (N_1904,In_3,In_913);
nor U1905 (N_1905,In_994,In_325);
nand U1906 (N_1906,In_879,In_656);
or U1907 (N_1907,In_125,In_763);
or U1908 (N_1908,In_161,In_294);
xnor U1909 (N_1909,In_915,In_260);
nor U1910 (N_1910,In_337,In_475);
and U1911 (N_1911,In_724,In_95);
nor U1912 (N_1912,In_117,In_826);
nor U1913 (N_1913,In_438,In_902);
and U1914 (N_1914,In_503,In_290);
nor U1915 (N_1915,In_347,In_453);
nand U1916 (N_1916,In_918,In_570);
or U1917 (N_1917,In_350,In_638);
nand U1918 (N_1918,In_537,In_790);
or U1919 (N_1919,In_120,In_593);
or U1920 (N_1920,In_628,In_365);
or U1921 (N_1921,In_364,In_311);
xor U1922 (N_1922,In_698,In_166);
nor U1923 (N_1923,In_324,In_183);
and U1924 (N_1924,In_151,In_941);
xor U1925 (N_1925,In_883,In_106);
or U1926 (N_1926,In_327,In_59);
nand U1927 (N_1927,In_410,In_131);
nand U1928 (N_1928,In_464,In_725);
or U1929 (N_1929,In_624,In_111);
nor U1930 (N_1930,In_873,In_853);
nand U1931 (N_1931,In_185,In_424);
nand U1932 (N_1932,In_699,In_632);
nand U1933 (N_1933,In_733,In_832);
or U1934 (N_1934,In_719,In_464);
nand U1935 (N_1935,In_310,In_487);
nand U1936 (N_1936,In_107,In_599);
or U1937 (N_1937,In_641,In_850);
xnor U1938 (N_1938,In_14,In_578);
or U1939 (N_1939,In_885,In_182);
xor U1940 (N_1940,In_453,In_300);
nand U1941 (N_1941,In_908,In_296);
nand U1942 (N_1942,In_196,In_546);
nor U1943 (N_1943,In_879,In_757);
nor U1944 (N_1944,In_884,In_890);
xor U1945 (N_1945,In_80,In_76);
or U1946 (N_1946,In_411,In_726);
xnor U1947 (N_1947,In_634,In_625);
or U1948 (N_1948,In_467,In_545);
xor U1949 (N_1949,In_35,In_856);
nor U1950 (N_1950,In_358,In_487);
nand U1951 (N_1951,In_40,In_337);
nand U1952 (N_1952,In_553,In_401);
or U1953 (N_1953,In_52,In_295);
or U1954 (N_1954,In_930,In_628);
nor U1955 (N_1955,In_846,In_244);
nor U1956 (N_1956,In_495,In_220);
nor U1957 (N_1957,In_60,In_50);
nor U1958 (N_1958,In_56,In_550);
xor U1959 (N_1959,In_946,In_736);
xnor U1960 (N_1960,In_696,In_475);
xnor U1961 (N_1961,In_823,In_294);
or U1962 (N_1962,In_32,In_197);
nand U1963 (N_1963,In_806,In_856);
nand U1964 (N_1964,In_173,In_930);
or U1965 (N_1965,In_862,In_672);
and U1966 (N_1966,In_426,In_631);
nor U1967 (N_1967,In_684,In_606);
xor U1968 (N_1968,In_194,In_9);
nor U1969 (N_1969,In_717,In_232);
xor U1970 (N_1970,In_996,In_159);
xor U1971 (N_1971,In_22,In_493);
or U1972 (N_1972,In_174,In_794);
xnor U1973 (N_1973,In_924,In_951);
and U1974 (N_1974,In_733,In_824);
nand U1975 (N_1975,In_192,In_673);
nand U1976 (N_1976,In_800,In_768);
nor U1977 (N_1977,In_810,In_369);
xor U1978 (N_1978,In_798,In_263);
and U1979 (N_1979,In_443,In_279);
nand U1980 (N_1980,In_884,In_954);
and U1981 (N_1981,In_714,In_170);
nor U1982 (N_1982,In_808,In_416);
and U1983 (N_1983,In_725,In_217);
or U1984 (N_1984,In_347,In_445);
and U1985 (N_1985,In_750,In_170);
nor U1986 (N_1986,In_308,In_921);
nand U1987 (N_1987,In_520,In_175);
nor U1988 (N_1988,In_810,In_69);
xor U1989 (N_1989,In_594,In_978);
nor U1990 (N_1990,In_284,In_737);
nand U1991 (N_1991,In_642,In_838);
nor U1992 (N_1992,In_312,In_641);
nand U1993 (N_1993,In_489,In_809);
nor U1994 (N_1994,In_876,In_467);
nand U1995 (N_1995,In_805,In_694);
or U1996 (N_1996,In_300,In_627);
or U1997 (N_1997,In_142,In_901);
nor U1998 (N_1998,In_173,In_975);
nor U1999 (N_1999,In_106,In_379);
and U2000 (N_2000,In_291,In_679);
nand U2001 (N_2001,In_398,In_931);
nor U2002 (N_2002,In_285,In_806);
nor U2003 (N_2003,In_567,In_978);
nor U2004 (N_2004,In_672,In_250);
or U2005 (N_2005,In_681,In_422);
xor U2006 (N_2006,In_846,In_858);
and U2007 (N_2007,In_172,In_167);
or U2008 (N_2008,In_623,In_601);
nor U2009 (N_2009,In_336,In_643);
nand U2010 (N_2010,In_986,In_558);
or U2011 (N_2011,In_305,In_467);
nor U2012 (N_2012,In_900,In_419);
nand U2013 (N_2013,In_252,In_118);
nor U2014 (N_2014,In_555,In_672);
and U2015 (N_2015,In_198,In_392);
or U2016 (N_2016,In_37,In_122);
or U2017 (N_2017,In_236,In_394);
xnor U2018 (N_2018,In_621,In_260);
nand U2019 (N_2019,In_876,In_494);
nand U2020 (N_2020,In_974,In_891);
xnor U2021 (N_2021,In_976,In_624);
or U2022 (N_2022,In_302,In_250);
nor U2023 (N_2023,In_192,In_605);
xor U2024 (N_2024,In_506,In_156);
xor U2025 (N_2025,In_426,In_19);
nand U2026 (N_2026,In_163,In_246);
or U2027 (N_2027,In_95,In_544);
or U2028 (N_2028,In_905,In_818);
nor U2029 (N_2029,In_442,In_192);
and U2030 (N_2030,In_222,In_104);
or U2031 (N_2031,In_293,In_481);
xnor U2032 (N_2032,In_497,In_994);
nand U2033 (N_2033,In_957,In_862);
nand U2034 (N_2034,In_818,In_753);
and U2035 (N_2035,In_187,In_361);
nor U2036 (N_2036,In_429,In_115);
nand U2037 (N_2037,In_630,In_247);
nand U2038 (N_2038,In_759,In_986);
xor U2039 (N_2039,In_43,In_682);
xor U2040 (N_2040,In_895,In_709);
nor U2041 (N_2041,In_994,In_962);
nor U2042 (N_2042,In_575,In_485);
nand U2043 (N_2043,In_447,In_944);
nor U2044 (N_2044,In_376,In_50);
nor U2045 (N_2045,In_474,In_493);
xnor U2046 (N_2046,In_86,In_270);
or U2047 (N_2047,In_647,In_608);
and U2048 (N_2048,In_88,In_457);
nand U2049 (N_2049,In_31,In_527);
xor U2050 (N_2050,In_123,In_759);
nor U2051 (N_2051,In_655,In_926);
and U2052 (N_2052,In_525,In_451);
nand U2053 (N_2053,In_848,In_162);
nand U2054 (N_2054,In_534,In_254);
nor U2055 (N_2055,In_866,In_738);
nor U2056 (N_2056,In_686,In_188);
xnor U2057 (N_2057,In_555,In_779);
or U2058 (N_2058,In_479,In_767);
xnor U2059 (N_2059,In_188,In_214);
and U2060 (N_2060,In_785,In_353);
or U2061 (N_2061,In_159,In_347);
and U2062 (N_2062,In_281,In_680);
nand U2063 (N_2063,In_836,In_862);
nand U2064 (N_2064,In_101,In_238);
nand U2065 (N_2065,In_581,In_478);
and U2066 (N_2066,In_908,In_447);
xnor U2067 (N_2067,In_187,In_570);
nand U2068 (N_2068,In_902,In_137);
nor U2069 (N_2069,In_146,In_368);
nor U2070 (N_2070,In_707,In_808);
or U2071 (N_2071,In_116,In_753);
and U2072 (N_2072,In_88,In_808);
xor U2073 (N_2073,In_331,In_524);
xnor U2074 (N_2074,In_935,In_497);
nor U2075 (N_2075,In_186,In_977);
nand U2076 (N_2076,In_755,In_381);
nand U2077 (N_2077,In_883,In_810);
or U2078 (N_2078,In_499,In_960);
and U2079 (N_2079,In_950,In_510);
and U2080 (N_2080,In_989,In_761);
xor U2081 (N_2081,In_936,In_444);
nand U2082 (N_2082,In_957,In_489);
nor U2083 (N_2083,In_890,In_211);
or U2084 (N_2084,In_19,In_496);
nand U2085 (N_2085,In_716,In_538);
xnor U2086 (N_2086,In_724,In_259);
or U2087 (N_2087,In_631,In_361);
nand U2088 (N_2088,In_317,In_856);
nand U2089 (N_2089,In_336,In_404);
nor U2090 (N_2090,In_968,In_892);
nor U2091 (N_2091,In_385,In_119);
or U2092 (N_2092,In_706,In_957);
or U2093 (N_2093,In_148,In_450);
or U2094 (N_2094,In_801,In_523);
or U2095 (N_2095,In_167,In_959);
or U2096 (N_2096,In_298,In_198);
and U2097 (N_2097,In_136,In_898);
nor U2098 (N_2098,In_221,In_369);
xnor U2099 (N_2099,In_328,In_965);
nor U2100 (N_2100,In_621,In_868);
nand U2101 (N_2101,In_246,In_448);
or U2102 (N_2102,In_259,In_407);
nand U2103 (N_2103,In_313,In_1);
and U2104 (N_2104,In_785,In_957);
nor U2105 (N_2105,In_803,In_924);
xnor U2106 (N_2106,In_323,In_381);
xnor U2107 (N_2107,In_26,In_156);
nand U2108 (N_2108,In_780,In_506);
and U2109 (N_2109,In_44,In_921);
nor U2110 (N_2110,In_827,In_304);
or U2111 (N_2111,In_498,In_645);
xor U2112 (N_2112,In_749,In_672);
or U2113 (N_2113,In_354,In_559);
or U2114 (N_2114,In_673,In_439);
nor U2115 (N_2115,In_899,In_218);
nand U2116 (N_2116,In_681,In_654);
nand U2117 (N_2117,In_676,In_743);
xnor U2118 (N_2118,In_73,In_182);
and U2119 (N_2119,In_717,In_330);
nand U2120 (N_2120,In_164,In_959);
nor U2121 (N_2121,In_678,In_932);
and U2122 (N_2122,In_16,In_668);
or U2123 (N_2123,In_606,In_545);
xor U2124 (N_2124,In_664,In_331);
or U2125 (N_2125,In_909,In_158);
nor U2126 (N_2126,In_734,In_280);
or U2127 (N_2127,In_821,In_474);
xor U2128 (N_2128,In_946,In_431);
nand U2129 (N_2129,In_287,In_154);
nor U2130 (N_2130,In_682,In_492);
nor U2131 (N_2131,In_749,In_474);
xor U2132 (N_2132,In_883,In_129);
nor U2133 (N_2133,In_759,In_42);
nand U2134 (N_2134,In_587,In_712);
xnor U2135 (N_2135,In_356,In_370);
or U2136 (N_2136,In_142,In_761);
and U2137 (N_2137,In_861,In_155);
nand U2138 (N_2138,In_340,In_951);
xor U2139 (N_2139,In_131,In_233);
nand U2140 (N_2140,In_273,In_155);
and U2141 (N_2141,In_898,In_189);
xnor U2142 (N_2142,In_382,In_623);
nand U2143 (N_2143,In_793,In_904);
and U2144 (N_2144,In_869,In_560);
or U2145 (N_2145,In_854,In_334);
nand U2146 (N_2146,In_77,In_905);
nor U2147 (N_2147,In_911,In_818);
and U2148 (N_2148,In_589,In_92);
nor U2149 (N_2149,In_285,In_763);
xor U2150 (N_2150,In_200,In_57);
or U2151 (N_2151,In_895,In_766);
nand U2152 (N_2152,In_578,In_816);
nor U2153 (N_2153,In_594,In_829);
and U2154 (N_2154,In_991,In_342);
and U2155 (N_2155,In_643,In_415);
nand U2156 (N_2156,In_957,In_53);
or U2157 (N_2157,In_499,In_609);
xor U2158 (N_2158,In_992,In_835);
nor U2159 (N_2159,In_410,In_843);
nor U2160 (N_2160,In_661,In_302);
or U2161 (N_2161,In_957,In_248);
xnor U2162 (N_2162,In_998,In_171);
nor U2163 (N_2163,In_268,In_817);
or U2164 (N_2164,In_496,In_191);
or U2165 (N_2165,In_669,In_641);
nor U2166 (N_2166,In_412,In_857);
and U2167 (N_2167,In_964,In_474);
xnor U2168 (N_2168,In_354,In_710);
xor U2169 (N_2169,In_706,In_625);
nor U2170 (N_2170,In_148,In_342);
nand U2171 (N_2171,In_370,In_321);
xor U2172 (N_2172,In_899,In_578);
or U2173 (N_2173,In_15,In_88);
or U2174 (N_2174,In_843,In_408);
xor U2175 (N_2175,In_758,In_374);
nand U2176 (N_2176,In_73,In_392);
and U2177 (N_2177,In_496,In_894);
nor U2178 (N_2178,In_867,In_386);
and U2179 (N_2179,In_924,In_742);
nor U2180 (N_2180,In_201,In_133);
and U2181 (N_2181,In_815,In_992);
nor U2182 (N_2182,In_759,In_187);
nor U2183 (N_2183,In_553,In_106);
nor U2184 (N_2184,In_944,In_332);
nand U2185 (N_2185,In_107,In_467);
xor U2186 (N_2186,In_794,In_155);
xor U2187 (N_2187,In_835,In_326);
or U2188 (N_2188,In_510,In_142);
nand U2189 (N_2189,In_575,In_708);
and U2190 (N_2190,In_384,In_751);
nand U2191 (N_2191,In_886,In_652);
nand U2192 (N_2192,In_756,In_105);
and U2193 (N_2193,In_188,In_308);
or U2194 (N_2194,In_378,In_830);
and U2195 (N_2195,In_350,In_938);
nor U2196 (N_2196,In_45,In_150);
nor U2197 (N_2197,In_668,In_522);
or U2198 (N_2198,In_129,In_541);
nand U2199 (N_2199,In_352,In_170);
xor U2200 (N_2200,In_513,In_32);
and U2201 (N_2201,In_197,In_319);
and U2202 (N_2202,In_246,In_684);
nand U2203 (N_2203,In_346,In_293);
nand U2204 (N_2204,In_480,In_874);
nand U2205 (N_2205,In_880,In_102);
or U2206 (N_2206,In_995,In_22);
xnor U2207 (N_2207,In_420,In_901);
or U2208 (N_2208,In_261,In_916);
nand U2209 (N_2209,In_543,In_982);
xnor U2210 (N_2210,In_606,In_818);
nand U2211 (N_2211,In_232,In_356);
and U2212 (N_2212,In_26,In_222);
and U2213 (N_2213,In_377,In_804);
nand U2214 (N_2214,In_984,In_721);
xor U2215 (N_2215,In_434,In_911);
nor U2216 (N_2216,In_407,In_811);
xor U2217 (N_2217,In_253,In_102);
and U2218 (N_2218,In_693,In_237);
or U2219 (N_2219,In_510,In_520);
and U2220 (N_2220,In_330,In_137);
nand U2221 (N_2221,In_594,In_27);
or U2222 (N_2222,In_320,In_30);
or U2223 (N_2223,In_429,In_441);
nand U2224 (N_2224,In_307,In_454);
xor U2225 (N_2225,In_139,In_993);
nand U2226 (N_2226,In_985,In_632);
and U2227 (N_2227,In_488,In_10);
nor U2228 (N_2228,In_20,In_240);
xor U2229 (N_2229,In_926,In_794);
and U2230 (N_2230,In_491,In_501);
nand U2231 (N_2231,In_193,In_9);
nand U2232 (N_2232,In_548,In_352);
xnor U2233 (N_2233,In_159,In_753);
or U2234 (N_2234,In_316,In_289);
nand U2235 (N_2235,In_549,In_54);
nand U2236 (N_2236,In_806,In_864);
xor U2237 (N_2237,In_781,In_226);
and U2238 (N_2238,In_630,In_839);
and U2239 (N_2239,In_540,In_765);
or U2240 (N_2240,In_46,In_948);
and U2241 (N_2241,In_870,In_984);
nor U2242 (N_2242,In_466,In_793);
nor U2243 (N_2243,In_564,In_196);
or U2244 (N_2244,In_740,In_374);
nor U2245 (N_2245,In_950,In_833);
and U2246 (N_2246,In_149,In_747);
nor U2247 (N_2247,In_71,In_12);
xnor U2248 (N_2248,In_687,In_388);
xnor U2249 (N_2249,In_592,In_499);
nand U2250 (N_2250,In_745,In_751);
and U2251 (N_2251,In_865,In_457);
nor U2252 (N_2252,In_238,In_356);
or U2253 (N_2253,In_994,In_838);
and U2254 (N_2254,In_412,In_139);
xor U2255 (N_2255,In_58,In_294);
and U2256 (N_2256,In_502,In_592);
nand U2257 (N_2257,In_353,In_551);
and U2258 (N_2258,In_605,In_965);
nor U2259 (N_2259,In_887,In_450);
nand U2260 (N_2260,In_500,In_696);
and U2261 (N_2261,In_315,In_245);
and U2262 (N_2262,In_893,In_257);
and U2263 (N_2263,In_612,In_632);
or U2264 (N_2264,In_292,In_360);
and U2265 (N_2265,In_183,In_428);
and U2266 (N_2266,In_750,In_216);
xor U2267 (N_2267,In_126,In_889);
xor U2268 (N_2268,In_167,In_197);
or U2269 (N_2269,In_651,In_386);
nor U2270 (N_2270,In_192,In_90);
or U2271 (N_2271,In_706,In_727);
xnor U2272 (N_2272,In_495,In_392);
xnor U2273 (N_2273,In_114,In_25);
nand U2274 (N_2274,In_907,In_322);
xor U2275 (N_2275,In_439,In_281);
nor U2276 (N_2276,In_532,In_758);
and U2277 (N_2277,In_131,In_590);
nor U2278 (N_2278,In_346,In_383);
or U2279 (N_2279,In_867,In_457);
xnor U2280 (N_2280,In_554,In_901);
and U2281 (N_2281,In_823,In_305);
nor U2282 (N_2282,In_235,In_269);
nor U2283 (N_2283,In_700,In_739);
nand U2284 (N_2284,In_158,In_772);
nor U2285 (N_2285,In_369,In_815);
or U2286 (N_2286,In_278,In_141);
nor U2287 (N_2287,In_183,In_540);
xor U2288 (N_2288,In_821,In_119);
nor U2289 (N_2289,In_432,In_663);
and U2290 (N_2290,In_973,In_818);
xnor U2291 (N_2291,In_20,In_954);
xor U2292 (N_2292,In_918,In_11);
xor U2293 (N_2293,In_461,In_488);
nor U2294 (N_2294,In_751,In_898);
nor U2295 (N_2295,In_530,In_140);
and U2296 (N_2296,In_448,In_939);
xnor U2297 (N_2297,In_844,In_151);
and U2298 (N_2298,In_719,In_281);
nor U2299 (N_2299,In_46,In_642);
xor U2300 (N_2300,In_118,In_168);
and U2301 (N_2301,In_179,In_762);
nor U2302 (N_2302,In_507,In_222);
nand U2303 (N_2303,In_859,In_22);
xor U2304 (N_2304,In_76,In_23);
and U2305 (N_2305,In_525,In_482);
or U2306 (N_2306,In_191,In_710);
nand U2307 (N_2307,In_343,In_90);
nand U2308 (N_2308,In_770,In_925);
or U2309 (N_2309,In_903,In_624);
xnor U2310 (N_2310,In_195,In_411);
nand U2311 (N_2311,In_867,In_689);
and U2312 (N_2312,In_850,In_57);
or U2313 (N_2313,In_146,In_948);
nor U2314 (N_2314,In_372,In_170);
nand U2315 (N_2315,In_904,In_119);
and U2316 (N_2316,In_651,In_467);
and U2317 (N_2317,In_212,In_422);
nor U2318 (N_2318,In_394,In_322);
and U2319 (N_2319,In_353,In_813);
or U2320 (N_2320,In_212,In_913);
or U2321 (N_2321,In_948,In_987);
nor U2322 (N_2322,In_369,In_75);
or U2323 (N_2323,In_760,In_853);
nor U2324 (N_2324,In_125,In_837);
nand U2325 (N_2325,In_47,In_327);
nand U2326 (N_2326,In_687,In_627);
nand U2327 (N_2327,In_162,In_726);
nor U2328 (N_2328,In_211,In_101);
and U2329 (N_2329,In_376,In_409);
xor U2330 (N_2330,In_625,In_243);
or U2331 (N_2331,In_220,In_693);
nand U2332 (N_2332,In_227,In_415);
nor U2333 (N_2333,In_336,In_938);
nand U2334 (N_2334,In_37,In_917);
nand U2335 (N_2335,In_524,In_188);
or U2336 (N_2336,In_423,In_162);
nor U2337 (N_2337,In_371,In_666);
xor U2338 (N_2338,In_676,In_299);
and U2339 (N_2339,In_623,In_61);
nand U2340 (N_2340,In_861,In_630);
and U2341 (N_2341,In_741,In_607);
nor U2342 (N_2342,In_847,In_915);
or U2343 (N_2343,In_511,In_565);
nor U2344 (N_2344,In_246,In_799);
nand U2345 (N_2345,In_43,In_269);
or U2346 (N_2346,In_454,In_898);
nand U2347 (N_2347,In_128,In_178);
xor U2348 (N_2348,In_538,In_350);
and U2349 (N_2349,In_594,In_896);
nor U2350 (N_2350,In_232,In_110);
nor U2351 (N_2351,In_501,In_291);
or U2352 (N_2352,In_9,In_905);
nand U2353 (N_2353,In_978,In_209);
or U2354 (N_2354,In_714,In_715);
or U2355 (N_2355,In_821,In_315);
xnor U2356 (N_2356,In_358,In_91);
nand U2357 (N_2357,In_726,In_673);
and U2358 (N_2358,In_691,In_775);
xnor U2359 (N_2359,In_105,In_798);
xnor U2360 (N_2360,In_853,In_250);
nand U2361 (N_2361,In_529,In_284);
nand U2362 (N_2362,In_552,In_243);
nor U2363 (N_2363,In_68,In_410);
nor U2364 (N_2364,In_903,In_239);
or U2365 (N_2365,In_260,In_846);
or U2366 (N_2366,In_732,In_379);
nor U2367 (N_2367,In_573,In_678);
nand U2368 (N_2368,In_841,In_949);
or U2369 (N_2369,In_567,In_339);
nor U2370 (N_2370,In_710,In_198);
or U2371 (N_2371,In_744,In_237);
and U2372 (N_2372,In_980,In_350);
nor U2373 (N_2373,In_634,In_732);
nor U2374 (N_2374,In_733,In_50);
and U2375 (N_2375,In_957,In_133);
nor U2376 (N_2376,In_953,In_692);
and U2377 (N_2377,In_194,In_941);
nor U2378 (N_2378,In_590,In_974);
nand U2379 (N_2379,In_616,In_177);
xnor U2380 (N_2380,In_401,In_105);
and U2381 (N_2381,In_733,In_232);
or U2382 (N_2382,In_881,In_49);
or U2383 (N_2383,In_149,In_624);
xor U2384 (N_2384,In_106,In_723);
and U2385 (N_2385,In_309,In_294);
and U2386 (N_2386,In_740,In_667);
nor U2387 (N_2387,In_925,In_745);
xor U2388 (N_2388,In_660,In_910);
nand U2389 (N_2389,In_990,In_548);
and U2390 (N_2390,In_876,In_401);
xor U2391 (N_2391,In_399,In_215);
nand U2392 (N_2392,In_271,In_472);
xor U2393 (N_2393,In_892,In_729);
nand U2394 (N_2394,In_161,In_14);
xnor U2395 (N_2395,In_987,In_405);
xnor U2396 (N_2396,In_872,In_432);
or U2397 (N_2397,In_282,In_976);
nand U2398 (N_2398,In_489,In_421);
and U2399 (N_2399,In_988,In_870);
nor U2400 (N_2400,In_761,In_660);
or U2401 (N_2401,In_748,In_179);
and U2402 (N_2402,In_768,In_764);
xnor U2403 (N_2403,In_27,In_104);
nand U2404 (N_2404,In_234,In_170);
nor U2405 (N_2405,In_664,In_890);
nor U2406 (N_2406,In_513,In_951);
nor U2407 (N_2407,In_454,In_849);
nor U2408 (N_2408,In_311,In_765);
xor U2409 (N_2409,In_482,In_273);
nand U2410 (N_2410,In_252,In_710);
nor U2411 (N_2411,In_568,In_247);
or U2412 (N_2412,In_29,In_976);
or U2413 (N_2413,In_757,In_790);
nand U2414 (N_2414,In_548,In_544);
nand U2415 (N_2415,In_998,In_801);
xnor U2416 (N_2416,In_361,In_235);
nor U2417 (N_2417,In_843,In_420);
and U2418 (N_2418,In_533,In_525);
or U2419 (N_2419,In_902,In_107);
or U2420 (N_2420,In_165,In_162);
nor U2421 (N_2421,In_168,In_907);
nand U2422 (N_2422,In_330,In_349);
nor U2423 (N_2423,In_321,In_0);
nand U2424 (N_2424,In_830,In_735);
and U2425 (N_2425,In_93,In_975);
and U2426 (N_2426,In_967,In_254);
nand U2427 (N_2427,In_237,In_963);
nand U2428 (N_2428,In_39,In_58);
and U2429 (N_2429,In_206,In_538);
or U2430 (N_2430,In_588,In_751);
nor U2431 (N_2431,In_821,In_229);
or U2432 (N_2432,In_227,In_501);
or U2433 (N_2433,In_981,In_749);
xnor U2434 (N_2434,In_271,In_408);
or U2435 (N_2435,In_835,In_784);
xor U2436 (N_2436,In_477,In_449);
nor U2437 (N_2437,In_69,In_32);
xnor U2438 (N_2438,In_622,In_9);
nor U2439 (N_2439,In_905,In_809);
or U2440 (N_2440,In_292,In_438);
nand U2441 (N_2441,In_798,In_546);
nor U2442 (N_2442,In_643,In_430);
or U2443 (N_2443,In_975,In_536);
xor U2444 (N_2444,In_562,In_607);
xnor U2445 (N_2445,In_842,In_183);
nand U2446 (N_2446,In_332,In_70);
or U2447 (N_2447,In_121,In_422);
and U2448 (N_2448,In_708,In_341);
and U2449 (N_2449,In_259,In_366);
nand U2450 (N_2450,In_65,In_176);
xnor U2451 (N_2451,In_168,In_261);
and U2452 (N_2452,In_131,In_42);
and U2453 (N_2453,In_905,In_685);
nor U2454 (N_2454,In_495,In_870);
and U2455 (N_2455,In_12,In_952);
and U2456 (N_2456,In_560,In_924);
and U2457 (N_2457,In_482,In_328);
nor U2458 (N_2458,In_290,In_598);
nand U2459 (N_2459,In_570,In_1);
nor U2460 (N_2460,In_937,In_202);
or U2461 (N_2461,In_524,In_128);
nand U2462 (N_2462,In_558,In_869);
and U2463 (N_2463,In_108,In_654);
or U2464 (N_2464,In_376,In_395);
or U2465 (N_2465,In_756,In_165);
nand U2466 (N_2466,In_298,In_636);
xor U2467 (N_2467,In_455,In_782);
xnor U2468 (N_2468,In_709,In_998);
or U2469 (N_2469,In_347,In_375);
or U2470 (N_2470,In_882,In_643);
xnor U2471 (N_2471,In_551,In_949);
xnor U2472 (N_2472,In_621,In_272);
or U2473 (N_2473,In_289,In_649);
or U2474 (N_2474,In_83,In_189);
nor U2475 (N_2475,In_23,In_777);
or U2476 (N_2476,In_739,In_282);
or U2477 (N_2477,In_206,In_780);
xnor U2478 (N_2478,In_685,In_736);
and U2479 (N_2479,In_811,In_376);
xor U2480 (N_2480,In_846,In_834);
xnor U2481 (N_2481,In_571,In_654);
nand U2482 (N_2482,In_615,In_943);
and U2483 (N_2483,In_705,In_650);
nor U2484 (N_2484,In_301,In_770);
xnor U2485 (N_2485,In_69,In_230);
and U2486 (N_2486,In_815,In_183);
and U2487 (N_2487,In_583,In_972);
and U2488 (N_2488,In_622,In_214);
or U2489 (N_2489,In_736,In_20);
nand U2490 (N_2490,In_758,In_109);
nand U2491 (N_2491,In_539,In_827);
nor U2492 (N_2492,In_582,In_233);
xnor U2493 (N_2493,In_424,In_967);
or U2494 (N_2494,In_844,In_502);
xnor U2495 (N_2495,In_581,In_838);
xnor U2496 (N_2496,In_556,In_890);
or U2497 (N_2497,In_532,In_805);
nand U2498 (N_2498,In_611,In_752);
or U2499 (N_2499,In_958,In_821);
nor U2500 (N_2500,N_1095,N_1412);
or U2501 (N_2501,N_1367,N_1971);
nor U2502 (N_2502,N_1697,N_780);
nor U2503 (N_2503,N_265,N_96);
or U2504 (N_2504,N_1411,N_601);
xnor U2505 (N_2505,N_118,N_366);
or U2506 (N_2506,N_881,N_758);
nand U2507 (N_2507,N_193,N_1829);
or U2508 (N_2508,N_2361,N_1600);
nand U2509 (N_2509,N_1693,N_1135);
and U2510 (N_2510,N_2493,N_2403);
or U2511 (N_2511,N_2191,N_888);
nor U2512 (N_2512,N_213,N_1319);
or U2513 (N_2513,N_389,N_1247);
or U2514 (N_2514,N_2266,N_1884);
nand U2515 (N_2515,N_1796,N_1136);
nor U2516 (N_2516,N_1432,N_2458);
nor U2517 (N_2517,N_1063,N_1535);
nand U2518 (N_2518,N_1107,N_2042);
or U2519 (N_2519,N_1056,N_198);
nor U2520 (N_2520,N_678,N_1210);
nor U2521 (N_2521,N_1325,N_830);
xor U2522 (N_2522,N_561,N_2419);
or U2523 (N_2523,N_2321,N_2429);
xnor U2524 (N_2524,N_2330,N_897);
nor U2525 (N_2525,N_651,N_1397);
xnor U2526 (N_2526,N_2380,N_1916);
and U2527 (N_2527,N_1553,N_622);
and U2528 (N_2528,N_1880,N_794);
or U2529 (N_2529,N_2464,N_548);
nand U2530 (N_2530,N_946,N_924);
nand U2531 (N_2531,N_14,N_104);
xor U2532 (N_2532,N_1155,N_330);
and U2533 (N_2533,N_2444,N_2479);
and U2534 (N_2534,N_869,N_1595);
and U2535 (N_2535,N_2433,N_683);
xnor U2536 (N_2536,N_2317,N_537);
nand U2537 (N_2537,N_1741,N_55);
xor U2538 (N_2538,N_1685,N_1018);
or U2539 (N_2539,N_880,N_1439);
and U2540 (N_2540,N_2267,N_2214);
nor U2541 (N_2541,N_1800,N_696);
nand U2542 (N_2542,N_287,N_783);
or U2543 (N_2543,N_1583,N_655);
nor U2544 (N_2544,N_268,N_2074);
nor U2545 (N_2545,N_2408,N_370);
and U2546 (N_2546,N_1363,N_1249);
or U2547 (N_2547,N_2168,N_484);
and U2548 (N_2548,N_1536,N_1642);
and U2549 (N_2549,N_1573,N_522);
xnor U2550 (N_2550,N_412,N_1031);
xor U2551 (N_2551,N_2044,N_1586);
xnor U2552 (N_2552,N_738,N_1818);
nand U2553 (N_2553,N_1620,N_2348);
or U2554 (N_2554,N_378,N_511);
nor U2555 (N_2555,N_823,N_525);
and U2556 (N_2556,N_886,N_441);
xnor U2557 (N_2557,N_75,N_1477);
xnor U2558 (N_2558,N_1719,N_917);
nand U2559 (N_2559,N_306,N_832);
or U2560 (N_2560,N_1455,N_2067);
xor U2561 (N_2561,N_1372,N_1323);
or U2562 (N_2562,N_1767,N_2095);
and U2563 (N_2563,N_439,N_178);
xor U2564 (N_2564,N_1085,N_1705);
and U2565 (N_2565,N_227,N_938);
nor U2566 (N_2566,N_175,N_2017);
nand U2567 (N_2567,N_2309,N_1909);
or U2568 (N_2568,N_637,N_600);
nor U2569 (N_2569,N_160,N_2012);
xor U2570 (N_2570,N_221,N_440);
nor U2571 (N_2571,N_803,N_183);
nand U2572 (N_2572,N_1288,N_1799);
and U2573 (N_2573,N_1327,N_593);
xnor U2574 (N_2574,N_1656,N_2430);
and U2575 (N_2575,N_2307,N_592);
xor U2576 (N_2576,N_515,N_2313);
xor U2577 (N_2577,N_1175,N_871);
nor U2578 (N_2578,N_1366,N_292);
xnor U2579 (N_2579,N_1330,N_2206);
nor U2580 (N_2580,N_1383,N_266);
nand U2581 (N_2581,N_2421,N_1130);
and U2582 (N_2582,N_1087,N_2287);
or U2583 (N_2583,N_749,N_1520);
nand U2584 (N_2584,N_752,N_58);
xnor U2585 (N_2585,N_902,N_1471);
nor U2586 (N_2586,N_1089,N_1368);
xnor U2587 (N_2587,N_813,N_1446);
or U2588 (N_2588,N_156,N_2473);
nor U2589 (N_2589,N_1613,N_144);
nand U2590 (N_2590,N_485,N_1710);
nand U2591 (N_2591,N_1202,N_801);
xor U2592 (N_2592,N_2412,N_1540);
or U2593 (N_2593,N_2056,N_984);
nand U2594 (N_2594,N_2132,N_1351);
xnor U2595 (N_2595,N_1533,N_429);
and U2596 (N_2596,N_455,N_559);
xor U2597 (N_2597,N_1352,N_730);
xor U2598 (N_2598,N_682,N_1810);
nor U2599 (N_2599,N_239,N_1606);
and U2600 (N_2600,N_1804,N_1762);
and U2601 (N_2601,N_2085,N_861);
or U2602 (N_2602,N_2183,N_566);
or U2603 (N_2603,N_69,N_1547);
xor U2604 (N_2604,N_1371,N_2410);
nor U2605 (N_2605,N_2450,N_1433);
nand U2606 (N_2606,N_1273,N_2062);
nor U2607 (N_2607,N_2010,N_164);
xor U2608 (N_2608,N_27,N_6);
and U2609 (N_2609,N_101,N_1773);
xor U2610 (N_2610,N_754,N_2050);
xnor U2611 (N_2611,N_840,N_1088);
nor U2612 (N_2612,N_1222,N_771);
xor U2613 (N_2613,N_2089,N_1476);
or U2614 (N_2614,N_271,N_1612);
nor U2615 (N_2615,N_661,N_1322);
nor U2616 (N_2616,N_1567,N_531);
nand U2617 (N_2617,N_1895,N_1725);
nor U2618 (N_2618,N_473,N_17);
and U2619 (N_2619,N_461,N_2277);
xor U2620 (N_2620,N_550,N_417);
xor U2621 (N_2621,N_1442,N_2388);
and U2622 (N_2622,N_1472,N_2019);
and U2623 (N_2623,N_2396,N_1918);
nor U2624 (N_2624,N_248,N_594);
nand U2625 (N_2625,N_505,N_1309);
nor U2626 (N_2626,N_2188,N_2407);
xor U2627 (N_2627,N_908,N_544);
xor U2628 (N_2628,N_1184,N_1188);
nor U2629 (N_2629,N_1931,N_2013);
nor U2630 (N_2630,N_2286,N_1444);
nor U2631 (N_2631,N_368,N_401);
and U2632 (N_2632,N_1126,N_1294);
xnor U2633 (N_2633,N_2457,N_769);
or U2634 (N_2634,N_1146,N_1002);
xor U2635 (N_2635,N_380,N_873);
nand U2636 (N_2636,N_512,N_1234);
or U2637 (N_2637,N_1060,N_2071);
or U2638 (N_2638,N_705,N_2283);
and U2639 (N_2639,N_1374,N_735);
xor U2640 (N_2640,N_451,N_2490);
xnor U2641 (N_2641,N_2375,N_2364);
nor U2642 (N_2642,N_1326,N_643);
and U2643 (N_2643,N_1317,N_2166);
xnor U2644 (N_2644,N_2088,N_1912);
xnor U2645 (N_2645,N_307,N_1496);
nand U2646 (N_2646,N_1039,N_234);
or U2647 (N_2647,N_639,N_1751);
and U2648 (N_2648,N_740,N_1350);
nand U2649 (N_2649,N_1101,N_2463);
nand U2650 (N_2650,N_961,N_932);
xor U2651 (N_2651,N_940,N_2365);
nand U2652 (N_2652,N_398,N_2440);
and U2653 (N_2653,N_2125,N_766);
nand U2654 (N_2654,N_2108,N_2338);
and U2655 (N_2655,N_1394,N_2387);
and U2656 (N_2656,N_2483,N_991);
nor U2657 (N_2657,N_952,N_1935);
or U2658 (N_2658,N_1193,N_145);
nor U2659 (N_2659,N_1008,N_1292);
nor U2660 (N_2660,N_2289,N_1783);
xor U2661 (N_2661,N_1297,N_706);
nand U2662 (N_2662,N_1438,N_1836);
nand U2663 (N_2663,N_720,N_2308);
nand U2664 (N_2664,N_1587,N_312);
or U2665 (N_2665,N_2343,N_1965);
nand U2666 (N_2666,N_826,N_1923);
or U2667 (N_2667,N_1563,N_475);
nand U2668 (N_2668,N_1359,N_1760);
nand U2669 (N_2669,N_1788,N_2219);
and U2670 (N_2670,N_2259,N_2316);
xnor U2671 (N_2671,N_1584,N_867);
or U2672 (N_2672,N_1118,N_1001);
nor U2673 (N_2673,N_648,N_588);
xnor U2674 (N_2674,N_1639,N_751);
or U2675 (N_2675,N_545,N_1734);
or U2676 (N_2676,N_2098,N_1548);
xnor U2677 (N_2677,N_1354,N_1930);
or U2678 (N_2678,N_486,N_778);
and U2679 (N_2679,N_2237,N_1495);
nor U2680 (N_2680,N_2101,N_2109);
or U2681 (N_2681,N_2350,N_963);
xnor U2682 (N_2682,N_1917,N_89);
nor U2683 (N_2683,N_857,N_650);
or U2684 (N_2684,N_1744,N_1956);
nor U2685 (N_2685,N_405,N_1882);
nor U2686 (N_2686,N_1399,N_246);
and U2687 (N_2687,N_1423,N_1950);
nor U2688 (N_2688,N_2366,N_1947);
xor U2689 (N_2689,N_1792,N_452);
or U2690 (N_2690,N_689,N_1979);
and U2691 (N_2691,N_806,N_1034);
nor U2692 (N_2692,N_2402,N_1329);
and U2693 (N_2693,N_2282,N_1516);
and U2694 (N_2694,N_553,N_812);
or U2695 (N_2695,N_1459,N_1772);
or U2696 (N_2696,N_1050,N_2244);
or U2697 (N_2697,N_1414,N_504);
nand U2698 (N_2698,N_976,N_2138);
and U2699 (N_2699,N_1901,N_1231);
nor U2700 (N_2700,N_1219,N_113);
xnor U2701 (N_2701,N_877,N_1190);
nand U2702 (N_2702,N_1504,N_797);
xnor U2703 (N_2703,N_304,N_1173);
xor U2704 (N_2704,N_2293,N_858);
or U2705 (N_2705,N_2498,N_937);
or U2706 (N_2706,N_189,N_392);
xor U2707 (N_2707,N_767,N_2294);
nand U2708 (N_2708,N_742,N_2137);
and U2709 (N_2709,N_1360,N_1550);
nand U2710 (N_2710,N_365,N_1942);
and U2711 (N_2711,N_158,N_2064);
or U2712 (N_2712,N_447,N_2130);
nor U2713 (N_2713,N_1373,N_2149);
and U2714 (N_2714,N_1825,N_586);
xor U2715 (N_2715,N_1742,N_19);
xor U2716 (N_2716,N_1053,N_1035);
xnor U2717 (N_2717,N_281,N_1384);
nor U2718 (N_2718,N_1278,N_1166);
or U2719 (N_2719,N_68,N_2382);
and U2720 (N_2720,N_1183,N_1740);
and U2721 (N_2721,N_2275,N_2416);
xnor U2722 (N_2722,N_1978,N_807);
xnor U2723 (N_2723,N_1889,N_1284);
nor U2724 (N_2724,N_980,N_2154);
nor U2725 (N_2725,N_1749,N_1280);
nand U2726 (N_2726,N_332,N_362);
or U2727 (N_2727,N_88,N_1057);
or U2728 (N_2728,N_2379,N_351);
xor U2729 (N_2729,N_2385,N_558);
nor U2730 (N_2730,N_646,N_149);
and U2731 (N_2731,N_381,N_1353);
or U2732 (N_2732,N_290,N_1843);
nand U2733 (N_2733,N_2371,N_151);
nor U2734 (N_2734,N_2049,N_264);
and U2735 (N_2735,N_1811,N_1678);
and U2736 (N_2736,N_2469,N_492);
and U2737 (N_2737,N_1827,N_192);
xor U2738 (N_2738,N_1908,N_1892);
or U2739 (N_2739,N_263,N_1768);
nand U2740 (N_2740,N_2273,N_1470);
xnor U2741 (N_2741,N_1750,N_50);
nand U2742 (N_2742,N_107,N_2424);
nor U2743 (N_2743,N_916,N_532);
xnor U2744 (N_2744,N_2492,N_1921);
or U2745 (N_2745,N_2376,N_1874);
xor U2746 (N_2746,N_513,N_1541);
or U2747 (N_2747,N_1066,N_1185);
xnor U2748 (N_2748,N_2081,N_1551);
or U2749 (N_2749,N_635,N_568);
nand U2750 (N_2750,N_49,N_1515);
nor U2751 (N_2751,N_2092,N_579);
nand U2752 (N_2752,N_1561,N_1481);
or U2753 (N_2753,N_708,N_37);
nand U2754 (N_2754,N_929,N_1664);
nand U2755 (N_2755,N_326,N_15);
or U2756 (N_2756,N_2008,N_1953);
or U2757 (N_2757,N_636,N_1969);
nor U2758 (N_2758,N_619,N_1047);
xor U2759 (N_2759,N_411,N_2076);
nor U2760 (N_2760,N_499,N_139);
or U2761 (N_2761,N_1659,N_704);
or U2762 (N_2762,N_575,N_785);
or U2763 (N_2763,N_895,N_1336);
and U2764 (N_2764,N_1011,N_2038);
nand U2765 (N_2765,N_2423,N_542);
or U2766 (N_2766,N_324,N_2115);
or U2767 (N_2767,N_2060,N_2271);
nand U2768 (N_2768,N_1159,N_1485);
or U2769 (N_2769,N_737,N_1033);
nor U2770 (N_2770,N_1267,N_755);
xnor U2771 (N_2771,N_1526,N_2459);
xnor U2772 (N_2772,N_1770,N_1487);
and U2773 (N_2773,N_339,N_1029);
nor U2774 (N_2774,N_2482,N_46);
nand U2775 (N_2775,N_2193,N_224);
nor U2776 (N_2776,N_2370,N_2028);
nand U2777 (N_2777,N_1915,N_746);
and U2778 (N_2778,N_465,N_186);
and U2779 (N_2779,N_2190,N_2180);
nor U2780 (N_2780,N_853,N_2356);
nor U2781 (N_2781,N_1385,N_2362);
and U2782 (N_2782,N_388,N_1198);
xnor U2783 (N_2783,N_2200,N_1262);
nand U2784 (N_2784,N_955,N_111);
nor U2785 (N_2785,N_2055,N_106);
and U2786 (N_2786,N_1165,N_2497);
xnor U2787 (N_2787,N_998,N_1502);
and U2788 (N_2788,N_317,N_623);
xnor U2789 (N_2789,N_663,N_1492);
nand U2790 (N_2790,N_358,N_1051);
xnor U2791 (N_2791,N_1524,N_1622);
and U2792 (N_2792,N_1009,N_2300);
nor U2793 (N_2793,N_349,N_702);
or U2794 (N_2794,N_2021,N_626);
nand U2795 (N_2795,N_933,N_1797);
and U2796 (N_2796,N_1562,N_1410);
and U2797 (N_2797,N_316,N_200);
or U2798 (N_2798,N_2318,N_296);
or U2799 (N_2799,N_483,N_2030);
xor U2800 (N_2800,N_1939,N_195);
xor U2801 (N_2801,N_1665,N_61);
or U2802 (N_2802,N_1589,N_1236);
nor U2803 (N_2803,N_1180,N_1940);
nand U2804 (N_2804,N_1084,N_1871);
or U2805 (N_2805,N_157,N_846);
and U2806 (N_2806,N_2220,N_115);
or U2807 (N_2807,N_1531,N_819);
nand U2808 (N_2808,N_2155,N_1679);
and U2809 (N_2809,N_141,N_2036);
and U2810 (N_2810,N_387,N_988);
nor U2811 (N_2811,N_2032,N_1582);
and U2812 (N_2812,N_876,N_1929);
or U2813 (N_2813,N_2007,N_864);
nand U2814 (N_2814,N_620,N_293);
and U2815 (N_2815,N_1069,N_957);
nand U2816 (N_2816,N_87,N_130);
or U2817 (N_2817,N_233,N_1452);
nand U2818 (N_2818,N_2290,N_2488);
xor U2819 (N_2819,N_294,N_1856);
nand U2820 (N_2820,N_43,N_533);
and U2821 (N_2821,N_1704,N_2360);
nor U2822 (N_2822,N_1689,N_2196);
nor U2823 (N_2823,N_887,N_1872);
nand U2824 (N_2824,N_1957,N_347);
xor U2825 (N_2825,N_267,N_97);
or U2826 (N_2826,N_904,N_2305);
nor U2827 (N_2827,N_1900,N_2248);
or U2828 (N_2828,N_1290,N_2175);
and U2829 (N_2829,N_1793,N_38);
xnor U2830 (N_2830,N_1698,N_674);
nor U2831 (N_2831,N_1149,N_1835);
xor U2832 (N_2832,N_975,N_1640);
xnor U2833 (N_2833,N_1102,N_1743);
nor U2834 (N_2834,N_1806,N_1464);
nor U2835 (N_2835,N_489,N_2009);
nor U2836 (N_2836,N_1898,N_1615);
nor U2837 (N_2837,N_1182,N_299);
xor U2838 (N_2838,N_1154,N_8);
or U2839 (N_2839,N_1143,N_1370);
and U2840 (N_2840,N_1728,N_2198);
xor U2841 (N_2841,N_2094,N_2186);
xor U2842 (N_2842,N_928,N_1150);
and U2843 (N_2843,N_926,N_1708);
or U2844 (N_2844,N_2241,N_1883);
nor U2845 (N_2845,N_12,N_2034);
and U2846 (N_2846,N_578,N_1514);
nand U2847 (N_2847,N_2112,N_2058);
nor U2848 (N_2848,N_2406,N_1733);
or U2849 (N_2849,N_260,N_194);
and U2850 (N_2850,N_76,N_1724);
and U2851 (N_2851,N_507,N_110);
xor U2852 (N_2852,N_434,N_1295);
and U2853 (N_2853,N_1120,N_182);
or U2854 (N_2854,N_1241,N_1272);
nand U2855 (N_2855,N_217,N_694);
and U2856 (N_2856,N_628,N_2075);
nand U2857 (N_2857,N_1924,N_787);
xnor U2858 (N_2858,N_2003,N_279);
nor U2859 (N_2859,N_1736,N_1707);
nand U2860 (N_2860,N_1824,N_1555);
nand U2861 (N_2861,N_2254,N_236);
or U2862 (N_2862,N_1177,N_2389);
nand U2863 (N_2863,N_53,N_1113);
xor U2864 (N_2864,N_2068,N_44);
and U2865 (N_2865,N_384,N_743);
or U2866 (N_2866,N_1505,N_1075);
xnor U2867 (N_2867,N_261,N_1259);
or U2868 (N_2868,N_1672,N_59);
and U2869 (N_2869,N_2472,N_2024);
nor U2870 (N_2870,N_2359,N_1137);
nor U2871 (N_2871,N_1176,N_1546);
nor U2872 (N_2872,N_1730,N_922);
nor U2873 (N_2873,N_1807,N_92);
xnor U2874 (N_2874,N_1129,N_1687);
nand U2875 (N_2875,N_2462,N_280);
or U2876 (N_2876,N_1049,N_199);
nor U2877 (N_2877,N_245,N_1192);
or U2878 (N_2878,N_1233,N_2461);
nand U2879 (N_2879,N_1349,N_1127);
nor U2880 (N_2880,N_1142,N_2331);
xor U2881 (N_2881,N_1320,N_135);
xnor U2882 (N_2882,N_1287,N_2182);
or U2883 (N_2883,N_218,N_1568);
or U2884 (N_2884,N_133,N_2026);
nor U2885 (N_2885,N_1922,N_257);
or U2886 (N_2886,N_659,N_1839);
nor U2887 (N_2887,N_1346,N_176);
xnor U2888 (N_2888,N_1885,N_2079);
or U2889 (N_2889,N_1948,N_1162);
nor U2890 (N_2890,N_894,N_2199);
and U2891 (N_2891,N_810,N_2097);
nand U2892 (N_2892,N_642,N_555);
or U2893 (N_2893,N_2128,N_1105);
nand U2894 (N_2894,N_1324,N_1347);
or U2895 (N_2895,N_796,N_2415);
xor U2896 (N_2896,N_1043,N_1691);
or U2897 (N_2897,N_2442,N_856);
xnor U2898 (N_2898,N_563,N_2054);
xnor U2899 (N_2899,N_2127,N_1610);
nand U2900 (N_2900,N_2288,N_1868);
nor U2901 (N_2901,N_1103,N_1906);
or U2902 (N_2902,N_855,N_374);
and U2903 (N_2903,N_1226,N_1987);
xor U2904 (N_2904,N_1172,N_1430);
xnor U2905 (N_2905,N_2306,N_1096);
and U2906 (N_2906,N_2373,N_445);
nor U2907 (N_2907,N_722,N_841);
nor U2908 (N_2908,N_2118,N_1756);
or U2909 (N_2909,N_1409,N_1614);
nand U2910 (N_2910,N_2184,N_1275);
or U2911 (N_2911,N_1914,N_725);
and U2912 (N_2912,N_656,N_212);
and U2913 (N_2913,N_1318,N_822);
nand U2914 (N_2914,N_424,N_571);
xnor U2915 (N_2915,N_1869,N_353);
nor U2916 (N_2916,N_1519,N_879);
and U2917 (N_2917,N_1626,N_2392);
nor U2918 (N_2918,N_1920,N_331);
nand U2919 (N_2919,N_1787,N_2156);
and U2920 (N_2920,N_1440,N_2414);
nand U2921 (N_2921,N_828,N_2411);
and U2922 (N_2922,N_1712,N_2192);
or U2923 (N_2923,N_1377,N_1201);
nor U2924 (N_2924,N_2471,N_123);
and U2925 (N_2925,N_632,N_786);
nor U2926 (N_2926,N_1237,N_476);
or U2927 (N_2927,N_1598,N_231);
xnor U2928 (N_2928,N_800,N_510);
nor U2929 (N_2929,N_993,N_2351);
xnor U2930 (N_2930,N_2453,N_30);
nor U2931 (N_2931,N_729,N_480);
nand U2932 (N_2932,N_1450,N_662);
and U2933 (N_2933,N_56,N_383);
and U2934 (N_2934,N_2016,N_216);
nor U2935 (N_2935,N_1308,N_1534);
xor U2936 (N_2936,N_891,N_762);
and U2937 (N_2937,N_538,N_1132);
xnor U2938 (N_2938,N_1268,N_2185);
nand U2939 (N_2939,N_1955,N_369);
and U2940 (N_2940,N_953,N_314);
and U2941 (N_2941,N_905,N_1167);
nand U2942 (N_2942,N_631,N_354);
nor U2943 (N_2943,N_676,N_1304);
xnor U2944 (N_2944,N_337,N_1988);
nand U2945 (N_2945,N_671,N_1170);
and U2946 (N_2946,N_313,N_892);
xor U2947 (N_2947,N_495,N_1688);
and U2948 (N_2948,N_1858,N_74);
nor U2949 (N_2949,N_413,N_2393);
or U2950 (N_2950,N_1980,N_1048);
nand U2951 (N_2951,N_1484,N_1161);
nand U2952 (N_2952,N_1617,N_1990);
nand U2953 (N_2953,N_284,N_1842);
xnor U2954 (N_2954,N_2436,N_634);
or U2955 (N_2955,N_968,N_1422);
or U2956 (N_2956,N_2466,N_1195);
and U2957 (N_2957,N_2377,N_1023);
nor U2958 (N_2958,N_969,N_909);
nand U2959 (N_2959,N_576,N_372);
nor U2960 (N_2960,N_1673,N_912);
xnor U2961 (N_2961,N_93,N_493);
or U2962 (N_2962,N_1572,N_1966);
and U2963 (N_2963,N_1337,N_2230);
nor U2964 (N_2964,N_1343,N_1151);
nand U2965 (N_2965,N_2123,N_143);
nor U2966 (N_2966,N_2104,N_1599);
or U2967 (N_2967,N_885,N_1960);
nand U2968 (N_2968,N_2255,N_535);
and U2969 (N_2969,N_1164,N_361);
xor U2970 (N_2970,N_971,N_1702);
nand U2971 (N_2971,N_1257,N_2195);
and U2972 (N_2972,N_2443,N_309);
nor U2973 (N_2973,N_836,N_272);
and U2974 (N_2974,N_835,N_915);
nand U2975 (N_2975,N_502,N_1396);
or U2976 (N_2976,N_2489,N_432);
or U2977 (N_2977,N_2435,N_1427);
and U2978 (N_2978,N_948,N_2209);
nand U2979 (N_2979,N_589,N_1527);
nand U2980 (N_2980,N_1671,N_477);
or U2981 (N_2981,N_181,N_1059);
and U2982 (N_2982,N_1191,N_1071);
nand U2983 (N_2983,N_709,N_1067);
nor U2984 (N_2984,N_2023,N_1072);
nor U2985 (N_2985,N_1755,N_630);
nor U2986 (N_2986,N_1356,N_2001);
or U2987 (N_2987,N_42,N_686);
nand U2988 (N_2988,N_1932,N_2378);
nand U2989 (N_2989,N_757,N_2027);
or U2990 (N_2990,N_1925,N_1348);
nor U2991 (N_2991,N_1566,N_2173);
xnor U2992 (N_2992,N_1285,N_2404);
nand U2993 (N_2993,N_668,N_277);
xnor U2994 (N_2994,N_845,N_2301);
nor U2995 (N_2995,N_1111,N_346);
nand U2996 (N_2996,N_1194,N_1601);
nor U2997 (N_2997,N_478,N_1879);
or U2998 (N_2998,N_155,N_2124);
xor U2999 (N_2999,N_1602,N_204);
xnor U3000 (N_3000,N_196,N_1860);
nor U3001 (N_3001,N_519,N_1577);
or U3002 (N_3002,N_1823,N_298);
nor U3003 (N_3003,N_591,N_1624);
nand U3004 (N_3004,N_863,N_1058);
nand U3005 (N_3005,N_638,N_2153);
xor U3006 (N_3006,N_1229,N_1675);
nor U3007 (N_3007,N_125,N_1692);
xor U3008 (N_3008,N_2323,N_1419);
and U3009 (N_3009,N_1670,N_1016);
or U3010 (N_3010,N_1260,N_1511);
and U3011 (N_3011,N_913,N_1303);
nand U3012 (N_3012,N_994,N_1019);
and U3013 (N_3013,N_291,N_1890);
or U3014 (N_3014,N_344,N_1886);
nand U3015 (N_3015,N_660,N_711);
and U3016 (N_3016,N_983,N_1493);
xnor U3017 (N_3017,N_718,N_1809);
and U3018 (N_3018,N_1144,N_1716);
nand U3019 (N_3019,N_142,N_2122);
or U3020 (N_3020,N_1061,N_464);
and U3021 (N_3021,N_2131,N_1145);
nor U3022 (N_3022,N_1400,N_1498);
nand U3023 (N_3023,N_816,N_1936);
xnor U3024 (N_3024,N_174,N_2272);
xnor U3025 (N_3025,N_2087,N_310);
and U3026 (N_3026,N_1635,N_450);
nor U3027 (N_3027,N_645,N_54);
xor U3028 (N_3028,N_159,N_1240);
nand U3029 (N_3029,N_860,N_136);
and U3030 (N_3030,N_893,N_1896);
or U3031 (N_3031,N_102,N_1156);
nand U3032 (N_3032,N_252,N_35);
nor U3033 (N_3033,N_1334,N_649);
nor U3034 (N_3034,N_2181,N_1134);
and U3035 (N_3035,N_396,N_792);
nor U3036 (N_3036,N_397,N_2033);
nor U3037 (N_3037,N_2400,N_1604);
or U3038 (N_3038,N_446,N_2434);
nand U3039 (N_3039,N_528,N_112);
xnor U3040 (N_3040,N_1482,N_691);
nor U3041 (N_3041,N_1510,N_1565);
nor U3042 (N_3042,N_105,N_2386);
nor U3043 (N_3043,N_1913,N_2136);
nand U3044 (N_3044,N_1388,N_616);
nand U3045 (N_3045,N_2349,N_2213);
xor U3046 (N_3046,N_1831,N_516);
and U3047 (N_3047,N_73,N_700);
nor U3048 (N_3048,N_851,N_2358);
nor U3049 (N_3049,N_884,N_852);
or U3050 (N_3050,N_163,N_2203);
nand U3051 (N_3051,N_1596,N_1844);
and U3052 (N_3052,N_972,N_1832);
and U3053 (N_3053,N_2102,N_540);
xor U3054 (N_3054,N_153,N_1274);
and U3055 (N_3055,N_2086,N_936);
nor U3056 (N_3056,N_2481,N_1949);
nor U3057 (N_3057,N_2228,N_1790);
and U3058 (N_3058,N_415,N_166);
or U3059 (N_3059,N_1657,N_1299);
nand U3060 (N_3060,N_1116,N_1616);
nand U3061 (N_3061,N_48,N_608);
nor U3062 (N_3062,N_169,N_1952);
xor U3063 (N_3063,N_422,N_318);
or U3064 (N_3064,N_918,N_79);
and U3065 (N_3065,N_1379,N_1000);
nor U3066 (N_3066,N_802,N_250);
nand U3067 (N_3067,N_629,N_2263);
nor U3068 (N_3068,N_1757,N_1888);
xor U3069 (N_3069,N_697,N_615);
and U3070 (N_3070,N_1305,N_1147);
and U3071 (N_3071,N_2151,N_1628);
nand U3072 (N_3072,N_315,N_744);
xnor U3073 (N_3073,N_1068,N_167);
nor U3074 (N_3074,N_1774,N_501);
and U3075 (N_3075,N_470,N_1878);
nor U3076 (N_3076,N_2212,N_1253);
nand U3077 (N_3077,N_1648,N_825);
nand U3078 (N_3078,N_161,N_1431);
or U3079 (N_3079,N_573,N_914);
and U3080 (N_3080,N_554,N_2096);
and U3081 (N_3081,N_214,N_1441);
xor U3082 (N_3082,N_494,N_99);
nor U3083 (N_3083,N_2035,N_419);
nand U3084 (N_3084,N_1927,N_1951);
nand U3085 (N_3085,N_2363,N_1763);
nand U3086 (N_3086,N_1121,N_1104);
nand U3087 (N_3087,N_1281,N_1243);
and U3088 (N_3088,N_225,N_2211);
nor U3089 (N_3089,N_1814,N_81);
or U3090 (N_3090,N_1518,N_596);
xnor U3091 (N_3091,N_1752,N_541);
or U3092 (N_3092,N_1458,N_844);
xnor U3093 (N_3093,N_2120,N_1296);
and U3094 (N_3094,N_753,N_1479);
nor U3095 (N_3095,N_18,N_459);
nor U3096 (N_3096,N_360,N_1578);
nor U3097 (N_3097,N_2157,N_180);
xnor U3098 (N_3098,N_944,N_1228);
or U3099 (N_3099,N_16,N_1390);
nand U3100 (N_3100,N_1298,N_2484);
nor U3101 (N_3101,N_1208,N_1808);
or U3102 (N_3102,N_109,N_1361);
or U3103 (N_3103,N_1417,N_866);
nand U3104 (N_3104,N_2070,N_2452);
or U3105 (N_3105,N_1517,N_530);
nor U3106 (N_3106,N_1769,N_1425);
and U3107 (N_3107,N_2409,N_1434);
and U3108 (N_3108,N_1037,N_1475);
or U3109 (N_3109,N_1025,N_1168);
and U3110 (N_3110,N_1682,N_1300);
and U3111 (N_3111,N_2384,N_2091);
or U3112 (N_3112,N_824,N_1532);
nor U3113 (N_3113,N_2161,N_262);
xor U3114 (N_3114,N_1786,N_259);
xnor U3115 (N_3115,N_698,N_2170);
xor U3116 (N_3116,N_1010,N_336);
nand U3117 (N_3117,N_40,N_1503);
nand U3118 (N_3118,N_1585,N_973);
or U3119 (N_3119,N_154,N_179);
nand U3120 (N_3120,N_831,N_2000);
xor U3121 (N_3121,N_52,N_2390);
xor U3122 (N_3122,N_1250,N_2);
or U3123 (N_3123,N_1854,N_2221);
nand U3124 (N_3124,N_1701,N_1497);
nor U3125 (N_3125,N_2210,N_2004);
nor U3126 (N_3126,N_673,N_818);
nor U3127 (N_3127,N_376,N_2285);
nand U3128 (N_3128,N_2395,N_2105);
nand U3129 (N_3129,N_2320,N_633);
xor U3130 (N_3130,N_232,N_60);
and U3131 (N_3131,N_2073,N_2047);
and U3132 (N_3132,N_308,N_41);
nand U3133 (N_3133,N_1469,N_872);
and U3134 (N_3134,N_29,N_784);
and U3135 (N_3135,N_128,N_1220);
nor U3136 (N_3136,N_1603,N_170);
xnor U3137 (N_3137,N_1451,N_235);
nand U3138 (N_3138,N_2456,N_274);
or U3139 (N_3139,N_203,N_1777);
or U3140 (N_3140,N_2218,N_2340);
and U3141 (N_3141,N_2332,N_719);
xor U3142 (N_3142,N_311,N_606);
nor U3143 (N_3143,N_1928,N_959);
nand U3144 (N_3144,N_408,N_300);
xor U3145 (N_3145,N_875,N_282);
nand U3146 (N_3146,N_1402,N_1958);
and U3147 (N_3147,N_1785,N_1509);
nor U3148 (N_3148,N_2401,N_1429);
and U3149 (N_3149,N_2239,N_1065);
xor U3150 (N_3150,N_241,N_1114);
nor U3151 (N_3151,N_574,N_865);
nand U3152 (N_3152,N_707,N_188);
or U3153 (N_3153,N_251,N_2278);
nand U3154 (N_3154,N_211,N_1209);
nor U3155 (N_3155,N_1386,N_114);
nor U3156 (N_3156,N_1128,N_1082);
or U3157 (N_3157,N_1643,N_564);
nor U3158 (N_3158,N_433,N_1408);
or U3159 (N_3159,N_2325,N_171);
xnor U3160 (N_3160,N_1711,N_13);
xor U3161 (N_3161,N_1086,N_805);
xnor U3162 (N_3162,N_958,N_1158);
xnor U3163 (N_3163,N_2291,N_527);
nor U3164 (N_3164,N_1232,N_24);
nand U3165 (N_3165,N_1982,N_609);
nand U3166 (N_3166,N_581,N_1647);
or U3167 (N_3167,N_927,N_1339);
nor U3168 (N_3168,N_423,N_1462);
nand U3169 (N_3169,N_243,N_2279);
xor U3170 (N_3170,N_2417,N_254);
nor U3171 (N_3171,N_2246,N_2225);
and U3172 (N_3172,N_1403,N_364);
and U3173 (N_3173,N_1761,N_301);
and U3174 (N_3174,N_333,N_1062);
nor U3175 (N_3175,N_140,N_456);
and U3176 (N_3176,N_652,N_1694);
xor U3177 (N_3177,N_2253,N_1283);
nand U3178 (N_3178,N_1560,N_1539);
nand U3179 (N_3179,N_2270,N_1798);
nand U3180 (N_3180,N_966,N_931);
nor U3181 (N_3181,N_1301,N_2355);
nand U3182 (N_3182,N_4,N_1124);
or U3183 (N_3183,N_1235,N_624);
xor U3184 (N_3184,N_1748,N_1052);
xnor U3185 (N_3185,N_701,N_741);
or U3186 (N_3186,N_1859,N_9);
xnor U3187 (N_3187,N_562,N_1621);
and U3188 (N_3188,N_1212,N_1508);
xnor U3189 (N_3189,N_47,N_1506);
xor U3190 (N_3190,N_585,N_416);
or U3191 (N_3191,N_1491,N_1406);
xor U3192 (N_3192,N_1112,N_1131);
nand U3193 (N_3193,N_1244,N_500);
nand U3194 (N_3194,N_614,N_95);
or U3195 (N_3195,N_848,N_1893);
nor U3196 (N_3196,N_2418,N_750);
nand U3197 (N_3197,N_1448,N_1381);
or U3198 (N_3198,N_1530,N_1703);
and U3199 (N_3199,N_1905,N_610);
or U3200 (N_3200,N_605,N_479);
nor U3201 (N_3201,N_1378,N_275);
xnor U3202 (N_3202,N_960,N_2468);
or U3203 (N_3203,N_1211,N_2235);
nand U3204 (N_3204,N_409,N_64);
nor U3205 (N_3205,N_1251,N_1254);
nand U3206 (N_3206,N_509,N_165);
xnor U3207 (N_3207,N_1611,N_2141);
nand U3208 (N_3208,N_2425,N_1090);
or U3209 (N_3209,N_1863,N_205);
and U3210 (N_3210,N_920,N_1331);
or U3211 (N_3211,N_2140,N_2159);
xnor U3212 (N_3212,N_138,N_2150);
nand U3213 (N_3213,N_1415,N_2252);
or U3214 (N_3214,N_1311,N_1593);
xnor U3215 (N_3215,N_2441,N_177);
nand U3216 (N_3216,N_517,N_2158);
and U3217 (N_3217,N_2245,N_103);
nor U3218 (N_3218,N_1847,N_1405);
and U3219 (N_3219,N_288,N_1046);
nand U3220 (N_3220,N_1269,N_2327);
and U3221 (N_3221,N_1108,N_728);
and U3222 (N_3222,N_1332,N_748);
xor U3223 (N_3223,N_172,N_685);
or U3224 (N_3224,N_2116,N_393);
xor U3225 (N_3225,N_989,N_453);
nand U3226 (N_3226,N_837,N_657);
nand U3227 (N_3227,N_108,N_799);
xor U3228 (N_3228,N_173,N_1674);
or U3229 (N_3229,N_1588,N_1099);
nand U3230 (N_3230,N_297,N_400);
nor U3231 (N_3231,N_703,N_1812);
xnor U3232 (N_3232,N_463,N_2480);
nor U3233 (N_3233,N_1115,N_2179);
xor U3234 (N_3234,N_1467,N_1307);
or U3235 (N_3235,N_1775,N_448);
nor U3236 (N_3236,N_1865,N_2238);
and U3237 (N_3237,N_1306,N_1213);
or U3238 (N_3238,N_1791,N_1457);
nand U3239 (N_3239,N_190,N_436);
or U3240 (N_3240,N_418,N_1934);
nor U3241 (N_3241,N_62,N_2224);
and U3242 (N_3242,N_1594,N_1737);
and U3243 (N_3243,N_2465,N_1853);
or U3244 (N_3244,N_1246,N_1499);
and U3245 (N_3245,N_1521,N_2052);
nor U3246 (N_3246,N_772,N_850);
or U3247 (N_3247,N_2448,N_1091);
xor U3248 (N_3248,N_1970,N_641);
and U3249 (N_3249,N_57,N_1501);
xor U3250 (N_3250,N_1849,N_2276);
xnor U3251 (N_3251,N_1005,N_1816);
nor U3252 (N_3252,N_1653,N_2121);
xor U3253 (N_3253,N_675,N_1081);
and U3254 (N_3254,N_1522,N_1215);
or U3255 (N_3255,N_739,N_595);
xor U3256 (N_3256,N_1972,N_2041);
nor U3257 (N_3257,N_759,N_1677);
nand U3258 (N_3258,N_1828,N_2084);
and U3259 (N_3259,N_230,N_134);
xor U3260 (N_3260,N_1255,N_839);
nor U3261 (N_3261,N_911,N_654);
nand U3262 (N_3262,N_467,N_2051);
xor U3263 (N_3263,N_2176,N_1026);
or U3264 (N_3264,N_1666,N_687);
nand U3265 (N_3265,N_2217,N_1223);
nor U3266 (N_3266,N_1852,N_402);
and U3267 (N_3267,N_1413,N_2284);
and U3268 (N_3268,N_1478,N_1512);
or U3269 (N_3269,N_1681,N_1999);
nor U3270 (N_3270,N_520,N_352);
or U3271 (N_3271,N_191,N_2455);
nor U3272 (N_3272,N_543,N_2326);
nand U3273 (N_3273,N_677,N_1894);
nor U3274 (N_3274,N_951,N_974);
xnor U3275 (N_3275,N_1608,N_1207);
xnor U3276 (N_3276,N_714,N_1735);
or U3277 (N_3277,N_699,N_1);
and U3278 (N_3278,N_63,N_947);
and U3279 (N_3279,N_693,N_1876);
or U3280 (N_3280,N_2142,N_2165);
xor U3281 (N_3281,N_1391,N_66);
or U3282 (N_3282,N_2207,N_420);
nor U3283 (N_3283,N_1851,N_1315);
and U3284 (N_3284,N_1739,N_1174);
nor U3285 (N_3285,N_1041,N_1358);
xnor U3286 (N_3286,N_1765,N_430);
or U3287 (N_3287,N_695,N_26);
nand U3288 (N_3288,N_1552,N_1080);
nand U3289 (N_3289,N_1899,N_1109);
or U3290 (N_3290,N_119,N_1821);
nor U3291 (N_3291,N_613,N_2240);
and U3292 (N_3292,N_255,N_1313);
nor U3293 (N_3293,N_583,N_90);
and U3294 (N_3294,N_777,N_1977);
xor U3295 (N_3295,N_1022,N_2432);
xor U3296 (N_3296,N_612,N_1850);
nor U3297 (N_3297,N_244,N_1286);
or U3298 (N_3298,N_2113,N_647);
xor U3299 (N_3299,N_1661,N_658);
nand U3300 (N_3300,N_1178,N_1110);
nand U3301 (N_3301,N_1845,N_406);
and U3302 (N_3302,N_286,N_25);
nor U3303 (N_3303,N_466,N_1658);
or U3304 (N_3304,N_2189,N_2059);
and U3305 (N_3305,N_1911,N_2256);
xnor U3306 (N_3306,N_1731,N_2445);
and U3307 (N_3307,N_1570,N_906);
nand U3308 (N_3308,N_2303,N_1722);
nor U3309 (N_3309,N_1224,N_1024);
or U3310 (N_3310,N_428,N_1962);
nor U3311 (N_3311,N_2110,N_2268);
and U3312 (N_3312,N_2446,N_1013);
xor U3313 (N_3313,N_356,N_1864);
and U3314 (N_3314,N_209,N_1727);
nand U3315 (N_3315,N_375,N_1314);
or U3316 (N_3316,N_2187,N_1686);
xor U3317 (N_3317,N_1345,N_2339);
and U3318 (N_3318,N_2460,N_228);
and U3319 (N_3319,N_363,N_549);
xor U3320 (N_3320,N_391,N_2139);
and U3321 (N_3321,N_442,N_1579);
nor U3322 (N_3322,N_1746,N_223);
xor U3323 (N_3323,N_2439,N_518);
nand U3324 (N_3324,N_1830,N_2477);
and U3325 (N_3325,N_2280,N_404);
nor U3326 (N_3326,N_427,N_1139);
or U3327 (N_3327,N_2106,N_2226);
nand U3328 (N_3328,N_2274,N_970);
nand U3329 (N_3329,N_2449,N_31);
xor U3330 (N_3330,N_1242,N_2144);
xnor U3331 (N_3331,N_2045,N_854);
and U3332 (N_3332,N_1776,N_1203);
nor U3333 (N_3333,N_2496,N_72);
xor U3334 (N_3334,N_1407,N_2258);
nand U3335 (N_3335,N_129,N_1891);
nor U3336 (N_3336,N_978,N_2133);
nor U3337 (N_3337,N_900,N_2039);
and U3338 (N_3338,N_1395,N_798);
nor U3339 (N_3339,N_421,N_890);
or U3340 (N_3340,N_1834,N_23);
xnor U3341 (N_3341,N_2428,N_506);
or U3342 (N_3342,N_1416,N_1239);
nor U3343 (N_3343,N_2099,N_1862);
nor U3344 (N_3344,N_2397,N_2447);
nand U3345 (N_3345,N_1160,N_552);
nor U3346 (N_3346,N_1044,N_491);
and U3347 (N_3347,N_2312,N_21);
nor U3348 (N_3348,N_2302,N_2269);
xor U3349 (N_3349,N_1684,N_1632);
nor U3350 (N_3350,N_723,N_116);
nand U3351 (N_3351,N_2061,N_1967);
or U3352 (N_3352,N_386,N_390);
xor U3353 (N_3353,N_664,N_982);
or U3354 (N_3354,N_1263,N_1592);
and U3355 (N_3355,N_2345,N_775);
or U3356 (N_3356,N_222,N_1873);
or U3357 (N_3357,N_1848,N_1456);
nand U3358 (N_3358,N_1754,N_2262);
nand U3359 (N_3359,N_577,N_2494);
nor U3360 (N_3360,N_3,N_127);
xor U3361 (N_3361,N_2357,N_1238);
and U3362 (N_3362,N_514,N_1357);
nor U3363 (N_3363,N_1073,N_1074);
nor U3364 (N_3364,N_793,N_1460);
and U3365 (N_3365,N_438,N_1994);
or U3366 (N_3366,N_907,N_237);
and U3367 (N_3367,N_458,N_2374);
nand U3368 (N_3368,N_882,N_2103);
nand U3369 (N_3369,N_2249,N_148);
or U3370 (N_3370,N_811,N_1045);
xnor U3371 (N_3371,N_1523,N_1070);
xnor U3372 (N_3372,N_295,N_2216);
and U3373 (N_3373,N_791,N_941);
xnor U3374 (N_3374,N_2474,N_1780);
nand U3375 (N_3375,N_903,N_2148);
nor U3376 (N_3376,N_1020,N_1214);
xnor U3377 (N_3377,N_747,N_2117);
xor U3378 (N_3378,N_469,N_327);
and U3379 (N_3379,N_1186,N_1597);
or U3380 (N_3380,N_379,N_1903);
and U3381 (N_3381,N_1718,N_1076);
xor U3382 (N_3382,N_584,N_348);
xor U3383 (N_3383,N_1758,N_2486);
or U3384 (N_3384,N_534,N_2369);
xnor U3385 (N_3385,N_2243,N_385);
or U3386 (N_3386,N_868,N_665);
nand U3387 (N_3387,N_329,N_1466);
nor U3388 (N_3388,N_2080,N_2025);
and U3389 (N_3389,N_2295,N_2005);
nand U3390 (N_3390,N_621,N_1837);
nand U3391 (N_3391,N_950,N_2162);
nor U3392 (N_3392,N_910,N_435);
xnor U3393 (N_3393,N_956,N_152);
nand U3394 (N_3394,N_1012,N_91);
nand U3395 (N_3395,N_1729,N_734);
xor U3396 (N_3396,N_1206,N_2352);
or U3397 (N_3397,N_618,N_782);
nor U3398 (N_3398,N_921,N_80);
nor U3399 (N_3399,N_1513,N_644);
and U3400 (N_3400,N_1205,N_2328);
and U3401 (N_3401,N_2476,N_779);
and U3402 (N_3402,N_833,N_33);
nor U3403 (N_3403,N_1445,N_2082);
and U3404 (N_3404,N_2065,N_2146);
and U3405 (N_3405,N_1720,N_488);
or U3406 (N_3406,N_45,N_1083);
xnor U3407 (N_3407,N_2354,N_611);
nor U3408 (N_3408,N_220,N_1557);
nor U3409 (N_3409,N_2311,N_487);
or U3410 (N_3410,N_2223,N_367);
or U3411 (N_3411,N_670,N_1453);
nand U3412 (N_3412,N_896,N_1655);
nand U3413 (N_3413,N_1549,N_2383);
and U3414 (N_3414,N_1803,N_1680);
or U3415 (N_3415,N_874,N_1463);
or U3416 (N_3416,N_472,N_849);
nor U3417 (N_3417,N_1380,N_399);
and U3418 (N_3418,N_2093,N_2090);
or U3419 (N_3419,N_1813,N_1996);
xnor U3420 (N_3420,N_1625,N_981);
and U3421 (N_3421,N_1974,N_2197);
or U3422 (N_3422,N_1537,N_817);
xor U3423 (N_3423,N_712,N_2431);
nand U3424 (N_3424,N_444,N_1590);
xor U3425 (N_3425,N_1265,N_862);
and U3426 (N_3426,N_1276,N_2368);
or U3427 (N_3427,N_736,N_1078);
nand U3428 (N_3428,N_2031,N_1338);
and U3429 (N_3429,N_1820,N_2399);
or U3430 (N_3430,N_1556,N_2367);
xor U3431 (N_3431,N_82,N_2002);
or U3432 (N_3432,N_350,N_1486);
or U3433 (N_3433,N_1870,N_1857);
nand U3434 (N_3434,N_1375,N_901);
nand U3435 (N_3435,N_2329,N_1230);
nor U3436 (N_3436,N_1645,N_1291);
nand U3437 (N_3437,N_667,N_1042);
nand U3438 (N_3438,N_1634,N_1545);
nor U3439 (N_3439,N_870,N_1805);
nor U3440 (N_3440,N_1525,N_790);
nand U3441 (N_3441,N_1569,N_343);
nand U3442 (N_3442,N_2126,N_2134);
and U3443 (N_3443,N_1316,N_1310);
or U3444 (N_3444,N_1745,N_2057);
xnor U3445 (N_3445,N_1003,N_1261);
nand U3446 (N_3446,N_1778,N_289);
nand U3447 (N_3447,N_2143,N_1875);
and U3448 (N_3448,N_2167,N_2053);
and U3449 (N_3449,N_137,N_1855);
xor U3450 (N_3450,N_774,N_834);
or U3451 (N_3451,N_580,N_1529);
nand U3452 (N_3452,N_878,N_1125);
nor U3453 (N_3453,N_2236,N_1248);
and U3454 (N_3454,N_1293,N_2135);
or U3455 (N_3455,N_1507,N_1877);
nor U3456 (N_3456,N_2420,N_1976);
xnor U3457 (N_3457,N_2495,N_2454);
xnor U3458 (N_3458,N_1961,N_320);
nand U3459 (N_3459,N_1264,N_2171);
and U3460 (N_3460,N_842,N_1437);
nor U3461 (N_3461,N_1833,N_1328);
nand U3462 (N_3462,N_1954,N_1822);
nand U3463 (N_3463,N_551,N_529);
or U3464 (N_3464,N_1169,N_508);
or U3465 (N_3465,N_319,N_1218);
or U3466 (N_3466,N_1838,N_1092);
and U3467 (N_3467,N_1897,N_1654);
xor U3468 (N_3468,N_999,N_185);
or U3469 (N_3469,N_1544,N_2438);
or U3470 (N_3470,N_2297,N_1271);
and U3471 (N_3471,N_2072,N_377);
xnor U3472 (N_3472,N_604,N_2398);
and U3473 (N_3473,N_51,N_1941);
and U3474 (N_3474,N_724,N_503);
or U3475 (N_3475,N_1717,N_765);
nand U3476 (N_3476,N_809,N_2296);
or U3477 (N_3477,N_1993,N_124);
nand U3478 (N_3478,N_1335,N_949);
nor U3479 (N_3479,N_1006,N_2422);
xnor U3480 (N_3480,N_2314,N_1344);
xnor U3481 (N_3481,N_2202,N_208);
or U3482 (N_3482,N_763,N_727);
nor U3483 (N_3483,N_602,N_2251);
xor U3484 (N_3484,N_2215,N_1795);
nand U3485 (N_3485,N_2169,N_126);
and U3486 (N_3486,N_617,N_1683);
nor U3487 (N_3487,N_342,N_2178);
nor U3488 (N_3488,N_283,N_1919);
nand U3489 (N_3489,N_640,N_1991);
xnor U3490 (N_3490,N_1782,N_2310);
nor U3491 (N_3491,N_1100,N_215);
and U3492 (N_3492,N_2029,N_395);
and U3493 (N_3493,N_546,N_919);
nor U3494 (N_3494,N_1968,N_431);
xor U3495 (N_3495,N_679,N_1538);
and U3496 (N_3496,N_1985,N_954);
nor U3497 (N_3497,N_1926,N_276);
and U3498 (N_3498,N_247,N_2381);
or U3499 (N_3499,N_2391,N_1392);
xnor U3500 (N_3500,N_672,N_1881);
and U3501 (N_3501,N_1571,N_1989);
nand U3502 (N_3502,N_70,N_2231);
xnor U3503 (N_3503,N_425,N_795);
nor U3504 (N_3504,N_745,N_1424);
or U3505 (N_3505,N_1696,N_1644);
xor U3506 (N_3506,N_147,N_2470);
and U3507 (N_3507,N_925,N_1771);
and U3508 (N_3508,N_990,N_407);
xnor U3509 (N_3509,N_1983,N_229);
or U3510 (N_3510,N_2205,N_403);
xor U3511 (N_3511,N_1910,N_2487);
and U3512 (N_3512,N_690,N_2485);
or U3513 (N_3513,N_1138,N_2324);
xnor U3514 (N_3514,N_2234,N_1591);
or U3515 (N_3515,N_979,N_1866);
nor U3516 (N_3516,N_1488,N_788);
xnor U3517 (N_3517,N_1428,N_2346);
and U3518 (N_3518,N_1054,N_1633);
nand U3519 (N_3519,N_1706,N_1017);
xnor U3520 (N_3520,N_899,N_1163);
xor U3521 (N_3521,N_1279,N_603);
nor U3522 (N_3522,N_2069,N_773);
nor U3523 (N_3523,N_1064,N_201);
nand U3524 (N_3524,N_582,N_1197);
and U3525 (N_3525,N_1365,N_207);
or U3526 (N_3526,N_84,N_680);
xor U3527 (N_3527,N_1418,N_526);
or U3528 (N_3528,N_1867,N_131);
or U3529 (N_3529,N_242,N_1270);
nor U3530 (N_3530,N_1699,N_2451);
and U3531 (N_3531,N_36,N_569);
nand U3532 (N_3532,N_1543,N_460);
xnor U3533 (N_3533,N_1646,N_721);
nor U3534 (N_3534,N_627,N_2174);
nor U3535 (N_3535,N_1559,N_847);
xnor U3536 (N_3536,N_1153,N_2242);
or U3537 (N_3537,N_2164,N_2043);
and U3538 (N_3538,N_71,N_1436);
or U3539 (N_3539,N_1030,N_1963);
nand U3540 (N_3540,N_768,N_1468);
nor U3541 (N_3541,N_820,N_1490);
xnor U3542 (N_3542,N_83,N_28);
or U3543 (N_3543,N_437,N_1618);
nor U3544 (N_3544,N_838,N_789);
nor U3545 (N_3545,N_557,N_1738);
nand U3546 (N_3546,N_1216,N_1630);
and U3547 (N_3547,N_821,N_1097);
xnor U3548 (N_3548,N_1055,N_2018);
xor U3549 (N_3549,N_1122,N_539);
xnor U3550 (N_3550,N_2077,N_1027);
nand U3551 (N_3551,N_964,N_713);
nand U3552 (N_3552,N_1171,N_468);
and U3553 (N_3553,N_2405,N_1542);
nor U3554 (N_3554,N_1494,N_1401);
or U3555 (N_3555,N_1605,N_0);
xnor U3556 (N_3556,N_1937,N_1997);
xor U3557 (N_3557,N_65,N_2322);
nand U3558 (N_3558,N_1489,N_2233);
nand U3559 (N_3559,N_1225,N_2194);
and U3560 (N_3560,N_607,N_2040);
nand U3561 (N_3561,N_2078,N_498);
or U3562 (N_3562,N_1021,N_1846);
xnor U3563 (N_3563,N_32,N_2037);
xnor U3564 (N_3564,N_341,N_2344);
and U3565 (N_3565,N_1117,N_939);
and U3566 (N_3566,N_1959,N_565);
nand U3567 (N_3567,N_22,N_132);
xor U3568 (N_3568,N_394,N_78);
and U3569 (N_3569,N_942,N_462);
nor U3570 (N_3570,N_883,N_967);
xnor U3571 (N_3571,N_1528,N_1732);
xor U3572 (N_3572,N_1904,N_776);
nor U3573 (N_3573,N_1981,N_1123);
and U3574 (N_3574,N_1652,N_1179);
xnor U3575 (N_3575,N_117,N_2372);
nor U3576 (N_3576,N_625,N_1028);
nand U3577 (N_3577,N_1461,N_1181);
or U3578 (N_3578,N_570,N_781);
or U3579 (N_3579,N_2083,N_2264);
or U3580 (N_3580,N_1077,N_1651);
xor U3581 (N_3581,N_1333,N_1801);
xor U3582 (N_3582,N_2163,N_669);
and U3583 (N_3583,N_325,N_815);
nand U3584 (N_3584,N_410,N_210);
nand U3585 (N_3585,N_567,N_1641);
nor U3586 (N_3586,N_1500,N_2353);
and U3587 (N_3587,N_1945,N_1695);
and U3588 (N_3588,N_1943,N_77);
xor U3589 (N_3589,N_1721,N_1764);
or U3590 (N_3590,N_497,N_808);
or U3591 (N_3591,N_1341,N_2046);
xor U3592 (N_3592,N_987,N_1637);
xnor U3593 (N_3593,N_340,N_731);
and U3594 (N_3594,N_2119,N_1714);
and U3595 (N_3595,N_2499,N_1669);
or U3596 (N_3596,N_1662,N_184);
nor U3597 (N_3597,N_2160,N_688);
nand U3598 (N_3598,N_1340,N_1631);
or U3599 (N_3599,N_1938,N_1819);
and U3600 (N_3600,N_1690,N_524);
nand U3601 (N_3601,N_345,N_1887);
or U3602 (N_3602,N_39,N_2250);
nor U3603 (N_3603,N_1474,N_162);
xor U3604 (N_3604,N_590,N_965);
or U3605 (N_3605,N_2426,N_1382);
or U3606 (N_3606,N_338,N_2201);
xor U3607 (N_3607,N_2304,N_2342);
xnor U3608 (N_3608,N_426,N_1040);
or U3609 (N_3609,N_373,N_1093);
or U3610 (N_3610,N_1404,N_187);
and U3611 (N_3611,N_1266,N_2152);
or U3612 (N_3612,N_1364,N_572);
or U3613 (N_3613,N_1036,N_1389);
nand U3614 (N_3614,N_1668,N_253);
or U3615 (N_3615,N_726,N_997);
nand U3616 (N_3616,N_355,N_2020);
or U3617 (N_3617,N_85,N_2114);
and U3618 (N_3618,N_1362,N_1933);
xnor U3619 (N_3619,N_2129,N_1355);
xor U3620 (N_3620,N_1342,N_547);
nor U3621 (N_3621,N_449,N_1014);
and U3622 (N_3622,N_985,N_86);
nor U3623 (N_3623,N_587,N_1700);
nor U3624 (N_3624,N_482,N_2022);
or U3625 (N_3625,N_328,N_1826);
nand U3626 (N_3626,N_710,N_1676);
xnor U3627 (N_3627,N_934,N_1709);
xor U3628 (N_3628,N_1581,N_206);
nand U3629 (N_3629,N_285,N_1079);
and U3630 (N_3630,N_303,N_1815);
nor U3631 (N_3631,N_2204,N_930);
nor U3632 (N_3632,N_7,N_760);
or U3633 (N_3633,N_2427,N_1221);
xnor U3634 (N_3634,N_2467,N_2394);
and U3635 (N_3635,N_556,N_1447);
nor U3636 (N_3636,N_2298,N_321);
nor U3637 (N_3637,N_1794,N_219);
xnor U3638 (N_3638,N_827,N_1321);
xor U3639 (N_3639,N_2107,N_2100);
or U3640 (N_3640,N_1964,N_273);
or U3641 (N_3641,N_1148,N_2147);
nor U3642 (N_3642,N_1106,N_1607);
nor U3643 (N_3643,N_335,N_2177);
nor U3644 (N_3644,N_943,N_1766);
or U3645 (N_3645,N_1227,N_1840);
and U3646 (N_3646,N_5,N_2478);
nor U3647 (N_3647,N_2063,N_1376);
xnor U3648 (N_3648,N_1907,N_1119);
nor U3649 (N_3649,N_1619,N_717);
xnor U3650 (N_3650,N_1667,N_1638);
or U3651 (N_3651,N_1189,N_322);
nand U3652 (N_3652,N_1973,N_1558);
nor U3653 (N_3653,N_1861,N_1726);
nand U3654 (N_3654,N_2145,N_1944);
nor U3655 (N_3655,N_121,N_1574);
xnor U3656 (N_3656,N_1609,N_1984);
nand U3657 (N_3657,N_2319,N_226);
or U3658 (N_3658,N_2475,N_1289);
nor U3659 (N_3659,N_443,N_1258);
or U3660 (N_3660,N_2066,N_1454);
or U3661 (N_3661,N_10,N_202);
and U3662 (N_3662,N_2315,N_716);
nand U3663 (N_3663,N_599,N_2335);
and U3664 (N_3664,N_414,N_681);
and U3665 (N_3665,N_2292,N_1480);
xor U3666 (N_3666,N_490,N_1660);
or U3667 (N_3667,N_715,N_2299);
nor U3668 (N_3668,N_1152,N_1623);
or U3669 (N_3669,N_34,N_2227);
nand U3670 (N_3670,N_1098,N_1252);
or U3671 (N_3671,N_1200,N_1196);
or U3672 (N_3672,N_2413,N_1449);
xor U3673 (N_3673,N_1369,N_457);
nor U3674 (N_3674,N_2172,N_598);
nand U3675 (N_3675,N_1443,N_122);
nor U3676 (N_3676,N_371,N_357);
nand U3677 (N_3677,N_2208,N_382);
xor U3678 (N_3678,N_1629,N_2232);
or U3679 (N_3679,N_684,N_120);
nor U3680 (N_3680,N_2006,N_258);
nand U3681 (N_3681,N_843,N_1784);
xor U3682 (N_3682,N_1627,N_1554);
or U3683 (N_3683,N_2048,N_1986);
and U3684 (N_3684,N_764,N_1998);
xor U3685 (N_3685,N_756,N_1421);
nor U3686 (N_3686,N_1841,N_1465);
nand U3687 (N_3687,N_1992,N_814);
or U3688 (N_3688,N_597,N_2334);
xnor U3689 (N_3689,N_692,N_761);
xnor U3690 (N_3690,N_1580,N_474);
or U3691 (N_3691,N_302,N_1781);
nand U3692 (N_3692,N_945,N_521);
nor U3693 (N_3693,N_2261,N_249);
xor U3694 (N_3694,N_1282,N_1398);
and U3695 (N_3695,N_278,N_1157);
xnor U3696 (N_3696,N_197,N_996);
nand U3697 (N_3697,N_2260,N_150);
xnor U3698 (N_3698,N_1564,N_2247);
xor U3699 (N_3699,N_1312,N_496);
nor U3700 (N_3700,N_240,N_2265);
nand U3701 (N_3701,N_67,N_923);
and U3702 (N_3702,N_334,N_1140);
nor U3703 (N_3703,N_359,N_1217);
xor U3704 (N_3704,N_94,N_1245);
xor U3705 (N_3705,N_1483,N_269);
and U3706 (N_3706,N_1789,N_732);
xor U3707 (N_3707,N_2333,N_1256);
nor U3708 (N_3708,N_889,N_1004);
nor U3709 (N_3709,N_20,N_2111);
xor U3710 (N_3710,N_962,N_1038);
and U3711 (N_3711,N_1420,N_1779);
or U3712 (N_3712,N_1649,N_100);
nand U3713 (N_3713,N_305,N_995);
nor U3714 (N_3714,N_146,N_256);
or U3715 (N_3715,N_98,N_1650);
or U3716 (N_3716,N_1713,N_1902);
and U3717 (N_3717,N_1723,N_1302);
xnor U3718 (N_3718,N_2011,N_481);
xor U3719 (N_3719,N_1817,N_1473);
nor U3720 (N_3720,N_2281,N_1015);
and U3721 (N_3721,N_977,N_1187);
nor U3722 (N_3722,N_829,N_1133);
and U3723 (N_3723,N_2222,N_1435);
nor U3724 (N_3724,N_2229,N_666);
or U3725 (N_3725,N_1277,N_454);
xor U3726 (N_3726,N_1199,N_898);
nand U3727 (N_3727,N_1032,N_1636);
and U3728 (N_3728,N_2014,N_770);
nand U3729 (N_3729,N_1426,N_992);
xnor U3730 (N_3730,N_536,N_1204);
nand U3731 (N_3731,N_804,N_323);
nand U3732 (N_3732,N_1576,N_1802);
xor U3733 (N_3733,N_1759,N_2437);
nor U3734 (N_3734,N_2347,N_1663);
nand U3735 (N_3735,N_238,N_986);
and U3736 (N_3736,N_1393,N_653);
nand U3737 (N_3737,N_2257,N_2341);
or U3738 (N_3738,N_1007,N_935);
nand U3739 (N_3739,N_2491,N_1094);
xor U3740 (N_3740,N_2337,N_859);
and U3741 (N_3741,N_2015,N_1995);
nand U3742 (N_3742,N_471,N_1575);
xnor U3743 (N_3743,N_2336,N_1753);
nor U3744 (N_3744,N_523,N_1715);
and U3745 (N_3745,N_270,N_1975);
xor U3746 (N_3746,N_1387,N_11);
or U3747 (N_3747,N_1141,N_560);
and U3748 (N_3748,N_1946,N_1747);
nand U3749 (N_3749,N_733,N_168);
nor U3750 (N_3750,N_2264,N_2080);
xnor U3751 (N_3751,N_1451,N_2414);
nor U3752 (N_3752,N_1831,N_2035);
and U3753 (N_3753,N_117,N_1704);
or U3754 (N_3754,N_1338,N_1915);
nor U3755 (N_3755,N_861,N_1594);
and U3756 (N_3756,N_1665,N_710);
or U3757 (N_3757,N_779,N_1632);
nand U3758 (N_3758,N_899,N_1201);
and U3759 (N_3759,N_2196,N_2435);
or U3760 (N_3760,N_418,N_2106);
nand U3761 (N_3761,N_488,N_349);
nand U3762 (N_3762,N_2087,N_2140);
nor U3763 (N_3763,N_1212,N_137);
nand U3764 (N_3764,N_596,N_1015);
and U3765 (N_3765,N_1743,N_1877);
nor U3766 (N_3766,N_1151,N_1693);
xor U3767 (N_3767,N_1748,N_2113);
nor U3768 (N_3768,N_1940,N_135);
and U3769 (N_3769,N_1920,N_515);
and U3770 (N_3770,N_580,N_777);
and U3771 (N_3771,N_1788,N_2120);
or U3772 (N_3772,N_2454,N_546);
or U3773 (N_3773,N_903,N_1880);
and U3774 (N_3774,N_2222,N_1371);
and U3775 (N_3775,N_965,N_2369);
xor U3776 (N_3776,N_299,N_185);
and U3777 (N_3777,N_351,N_167);
nand U3778 (N_3778,N_506,N_1855);
or U3779 (N_3779,N_224,N_1099);
nand U3780 (N_3780,N_1648,N_347);
nand U3781 (N_3781,N_1194,N_1007);
nand U3782 (N_3782,N_2156,N_2270);
nor U3783 (N_3783,N_476,N_1982);
nand U3784 (N_3784,N_488,N_1054);
nand U3785 (N_3785,N_1877,N_1958);
xnor U3786 (N_3786,N_2311,N_206);
or U3787 (N_3787,N_1623,N_1075);
nor U3788 (N_3788,N_143,N_1990);
xor U3789 (N_3789,N_1716,N_1196);
nand U3790 (N_3790,N_359,N_993);
nor U3791 (N_3791,N_1469,N_783);
nand U3792 (N_3792,N_750,N_385);
nor U3793 (N_3793,N_1077,N_1901);
or U3794 (N_3794,N_2030,N_1940);
nor U3795 (N_3795,N_242,N_2004);
and U3796 (N_3796,N_2343,N_2351);
nor U3797 (N_3797,N_1552,N_1707);
nand U3798 (N_3798,N_454,N_2018);
nor U3799 (N_3799,N_817,N_2416);
nand U3800 (N_3800,N_1045,N_1488);
and U3801 (N_3801,N_1505,N_443);
and U3802 (N_3802,N_559,N_233);
xnor U3803 (N_3803,N_1536,N_2012);
nand U3804 (N_3804,N_817,N_2092);
xnor U3805 (N_3805,N_42,N_501);
nand U3806 (N_3806,N_1203,N_1235);
and U3807 (N_3807,N_1328,N_901);
and U3808 (N_3808,N_1928,N_1585);
or U3809 (N_3809,N_2076,N_587);
xnor U3810 (N_3810,N_2190,N_2321);
nand U3811 (N_3811,N_2106,N_2351);
xor U3812 (N_3812,N_1679,N_676);
xor U3813 (N_3813,N_1172,N_1566);
nand U3814 (N_3814,N_964,N_153);
xor U3815 (N_3815,N_1855,N_219);
nor U3816 (N_3816,N_2161,N_1269);
nand U3817 (N_3817,N_738,N_544);
and U3818 (N_3818,N_114,N_165);
or U3819 (N_3819,N_1458,N_878);
nand U3820 (N_3820,N_1917,N_1347);
nor U3821 (N_3821,N_1497,N_1072);
nand U3822 (N_3822,N_660,N_1486);
nand U3823 (N_3823,N_1091,N_1710);
xor U3824 (N_3824,N_2068,N_216);
xor U3825 (N_3825,N_9,N_952);
or U3826 (N_3826,N_1938,N_1532);
nor U3827 (N_3827,N_630,N_202);
and U3828 (N_3828,N_1142,N_1856);
and U3829 (N_3829,N_1778,N_513);
xnor U3830 (N_3830,N_1574,N_2318);
or U3831 (N_3831,N_1549,N_188);
or U3832 (N_3832,N_2277,N_322);
xnor U3833 (N_3833,N_2399,N_2362);
and U3834 (N_3834,N_1137,N_371);
or U3835 (N_3835,N_1533,N_1439);
xor U3836 (N_3836,N_2049,N_2296);
nand U3837 (N_3837,N_1477,N_1461);
or U3838 (N_3838,N_290,N_1730);
nor U3839 (N_3839,N_784,N_148);
or U3840 (N_3840,N_1296,N_44);
xnor U3841 (N_3841,N_64,N_2400);
or U3842 (N_3842,N_2465,N_989);
nor U3843 (N_3843,N_1134,N_1795);
and U3844 (N_3844,N_206,N_669);
and U3845 (N_3845,N_118,N_57);
or U3846 (N_3846,N_1544,N_2484);
and U3847 (N_3847,N_2214,N_329);
nand U3848 (N_3848,N_1689,N_548);
nand U3849 (N_3849,N_1538,N_2005);
xnor U3850 (N_3850,N_104,N_1303);
or U3851 (N_3851,N_2452,N_2119);
and U3852 (N_3852,N_2434,N_2371);
and U3853 (N_3853,N_1176,N_818);
xor U3854 (N_3854,N_495,N_1903);
xor U3855 (N_3855,N_2008,N_219);
or U3856 (N_3856,N_1769,N_48);
xor U3857 (N_3857,N_1769,N_2197);
or U3858 (N_3858,N_1041,N_1047);
and U3859 (N_3859,N_33,N_2381);
or U3860 (N_3860,N_963,N_2481);
nor U3861 (N_3861,N_1195,N_2495);
or U3862 (N_3862,N_2084,N_1731);
xnor U3863 (N_3863,N_425,N_383);
or U3864 (N_3864,N_685,N_916);
or U3865 (N_3865,N_2177,N_694);
xor U3866 (N_3866,N_1334,N_199);
nor U3867 (N_3867,N_2066,N_1315);
or U3868 (N_3868,N_631,N_1787);
and U3869 (N_3869,N_415,N_1474);
and U3870 (N_3870,N_639,N_1052);
nor U3871 (N_3871,N_1668,N_1855);
and U3872 (N_3872,N_50,N_1668);
nand U3873 (N_3873,N_2278,N_955);
nand U3874 (N_3874,N_1694,N_1882);
or U3875 (N_3875,N_743,N_14);
or U3876 (N_3876,N_1498,N_904);
xnor U3877 (N_3877,N_2319,N_1084);
and U3878 (N_3878,N_1758,N_2227);
nand U3879 (N_3879,N_2225,N_1969);
and U3880 (N_3880,N_1561,N_994);
or U3881 (N_3881,N_1636,N_475);
xnor U3882 (N_3882,N_1236,N_1730);
nor U3883 (N_3883,N_1599,N_441);
nor U3884 (N_3884,N_463,N_1309);
or U3885 (N_3885,N_1416,N_2363);
nor U3886 (N_3886,N_219,N_680);
and U3887 (N_3887,N_2184,N_77);
and U3888 (N_3888,N_2025,N_914);
or U3889 (N_3889,N_1574,N_198);
nor U3890 (N_3890,N_657,N_148);
or U3891 (N_3891,N_1765,N_914);
nand U3892 (N_3892,N_1529,N_1498);
nand U3893 (N_3893,N_2056,N_1839);
or U3894 (N_3894,N_926,N_194);
and U3895 (N_3895,N_2205,N_351);
or U3896 (N_3896,N_1430,N_653);
nor U3897 (N_3897,N_1133,N_71);
or U3898 (N_3898,N_1875,N_2368);
nor U3899 (N_3899,N_1747,N_544);
or U3900 (N_3900,N_1988,N_441);
xor U3901 (N_3901,N_435,N_2201);
nand U3902 (N_3902,N_1948,N_1300);
or U3903 (N_3903,N_2006,N_1418);
nand U3904 (N_3904,N_194,N_1006);
xnor U3905 (N_3905,N_1509,N_2197);
and U3906 (N_3906,N_415,N_754);
nand U3907 (N_3907,N_2304,N_77);
nor U3908 (N_3908,N_942,N_1325);
nor U3909 (N_3909,N_973,N_2248);
nor U3910 (N_3910,N_1761,N_546);
and U3911 (N_3911,N_377,N_1771);
xor U3912 (N_3912,N_2494,N_1524);
and U3913 (N_3913,N_1076,N_1917);
or U3914 (N_3914,N_867,N_1118);
nand U3915 (N_3915,N_806,N_2095);
or U3916 (N_3916,N_1276,N_2014);
nand U3917 (N_3917,N_2152,N_736);
nand U3918 (N_3918,N_256,N_2366);
xor U3919 (N_3919,N_70,N_1536);
nand U3920 (N_3920,N_2460,N_1205);
nand U3921 (N_3921,N_627,N_2128);
nand U3922 (N_3922,N_1424,N_331);
nand U3923 (N_3923,N_632,N_567);
and U3924 (N_3924,N_1549,N_1868);
xor U3925 (N_3925,N_337,N_1900);
nand U3926 (N_3926,N_631,N_2302);
or U3927 (N_3927,N_2011,N_1542);
nor U3928 (N_3928,N_996,N_1669);
xnor U3929 (N_3929,N_1199,N_970);
nand U3930 (N_3930,N_796,N_1258);
and U3931 (N_3931,N_1287,N_1770);
xnor U3932 (N_3932,N_1756,N_373);
or U3933 (N_3933,N_1987,N_1012);
xnor U3934 (N_3934,N_719,N_1963);
nor U3935 (N_3935,N_2423,N_796);
and U3936 (N_3936,N_193,N_1544);
xnor U3937 (N_3937,N_1447,N_1261);
and U3938 (N_3938,N_2408,N_2492);
nor U3939 (N_3939,N_1741,N_1483);
nand U3940 (N_3940,N_662,N_94);
or U3941 (N_3941,N_1989,N_1733);
and U3942 (N_3942,N_1321,N_812);
nor U3943 (N_3943,N_303,N_1305);
or U3944 (N_3944,N_1982,N_1268);
and U3945 (N_3945,N_69,N_1900);
nand U3946 (N_3946,N_510,N_873);
and U3947 (N_3947,N_499,N_730);
nand U3948 (N_3948,N_30,N_964);
and U3949 (N_3949,N_1855,N_526);
nor U3950 (N_3950,N_266,N_1577);
or U3951 (N_3951,N_581,N_1211);
or U3952 (N_3952,N_206,N_1871);
and U3953 (N_3953,N_782,N_2107);
and U3954 (N_3954,N_1153,N_2393);
xor U3955 (N_3955,N_531,N_1904);
nor U3956 (N_3956,N_2330,N_1694);
or U3957 (N_3957,N_835,N_976);
or U3958 (N_3958,N_2268,N_1625);
and U3959 (N_3959,N_1445,N_1852);
nor U3960 (N_3960,N_737,N_2487);
xor U3961 (N_3961,N_1012,N_2202);
nand U3962 (N_3962,N_949,N_738);
and U3963 (N_3963,N_155,N_596);
nand U3964 (N_3964,N_939,N_197);
and U3965 (N_3965,N_734,N_30);
and U3966 (N_3966,N_1588,N_1439);
nor U3967 (N_3967,N_1031,N_710);
or U3968 (N_3968,N_547,N_58);
or U3969 (N_3969,N_715,N_418);
xor U3970 (N_3970,N_442,N_982);
xor U3971 (N_3971,N_1312,N_1545);
and U3972 (N_3972,N_1331,N_343);
and U3973 (N_3973,N_1297,N_1571);
nor U3974 (N_3974,N_1887,N_1838);
and U3975 (N_3975,N_2220,N_539);
or U3976 (N_3976,N_1412,N_1612);
or U3977 (N_3977,N_2423,N_301);
and U3978 (N_3978,N_2072,N_1308);
nand U3979 (N_3979,N_395,N_1022);
nor U3980 (N_3980,N_742,N_769);
xor U3981 (N_3981,N_1640,N_882);
nand U3982 (N_3982,N_273,N_2387);
nor U3983 (N_3983,N_113,N_725);
nand U3984 (N_3984,N_1513,N_1935);
or U3985 (N_3985,N_1027,N_506);
nor U3986 (N_3986,N_1271,N_2428);
xnor U3987 (N_3987,N_2280,N_2406);
nand U3988 (N_3988,N_466,N_1693);
nand U3989 (N_3989,N_457,N_1794);
or U3990 (N_3990,N_270,N_2034);
nand U3991 (N_3991,N_2495,N_1935);
xor U3992 (N_3992,N_2329,N_854);
nand U3993 (N_3993,N_2014,N_222);
and U3994 (N_3994,N_236,N_1071);
or U3995 (N_3995,N_2193,N_2062);
and U3996 (N_3996,N_276,N_2430);
or U3997 (N_3997,N_2418,N_1153);
and U3998 (N_3998,N_911,N_78);
or U3999 (N_3999,N_2030,N_1627);
nand U4000 (N_4000,N_165,N_1755);
and U4001 (N_4001,N_1912,N_911);
and U4002 (N_4002,N_916,N_175);
nand U4003 (N_4003,N_1665,N_1115);
nor U4004 (N_4004,N_2158,N_154);
nor U4005 (N_4005,N_2083,N_1064);
or U4006 (N_4006,N_1116,N_877);
nor U4007 (N_4007,N_89,N_1940);
nor U4008 (N_4008,N_293,N_2420);
nand U4009 (N_4009,N_1865,N_1463);
and U4010 (N_4010,N_1442,N_790);
or U4011 (N_4011,N_680,N_2369);
nor U4012 (N_4012,N_1140,N_1953);
xnor U4013 (N_4013,N_1075,N_466);
nand U4014 (N_4014,N_2188,N_2316);
or U4015 (N_4015,N_617,N_248);
nor U4016 (N_4016,N_637,N_2073);
or U4017 (N_4017,N_95,N_855);
or U4018 (N_4018,N_2292,N_1831);
and U4019 (N_4019,N_1253,N_635);
and U4020 (N_4020,N_2111,N_1855);
nor U4021 (N_4021,N_1742,N_2284);
nand U4022 (N_4022,N_862,N_561);
and U4023 (N_4023,N_2069,N_1387);
and U4024 (N_4024,N_2226,N_1679);
nand U4025 (N_4025,N_1791,N_80);
nor U4026 (N_4026,N_2362,N_1595);
nor U4027 (N_4027,N_551,N_937);
nor U4028 (N_4028,N_599,N_67);
and U4029 (N_4029,N_2493,N_2343);
nand U4030 (N_4030,N_2452,N_2496);
nand U4031 (N_4031,N_1465,N_1154);
or U4032 (N_4032,N_1098,N_1615);
nor U4033 (N_4033,N_913,N_1719);
nand U4034 (N_4034,N_1161,N_18);
nand U4035 (N_4035,N_1968,N_1192);
xor U4036 (N_4036,N_416,N_389);
nand U4037 (N_4037,N_1898,N_82);
xnor U4038 (N_4038,N_1815,N_585);
xnor U4039 (N_4039,N_1883,N_2134);
xor U4040 (N_4040,N_397,N_2212);
nand U4041 (N_4041,N_1860,N_706);
or U4042 (N_4042,N_2038,N_461);
or U4043 (N_4043,N_1625,N_1434);
xor U4044 (N_4044,N_2244,N_1594);
and U4045 (N_4045,N_2271,N_439);
nor U4046 (N_4046,N_843,N_1081);
nor U4047 (N_4047,N_707,N_1321);
xor U4048 (N_4048,N_419,N_2325);
xor U4049 (N_4049,N_1831,N_707);
or U4050 (N_4050,N_1249,N_2359);
xor U4051 (N_4051,N_1811,N_534);
or U4052 (N_4052,N_2347,N_2127);
and U4053 (N_4053,N_1101,N_2377);
nand U4054 (N_4054,N_1033,N_1613);
and U4055 (N_4055,N_1733,N_1029);
nand U4056 (N_4056,N_326,N_977);
xor U4057 (N_4057,N_2037,N_837);
and U4058 (N_4058,N_117,N_1539);
and U4059 (N_4059,N_1035,N_1940);
nor U4060 (N_4060,N_1098,N_461);
nor U4061 (N_4061,N_2004,N_206);
nand U4062 (N_4062,N_1069,N_1930);
and U4063 (N_4063,N_2283,N_595);
nor U4064 (N_4064,N_1419,N_643);
nand U4065 (N_4065,N_1162,N_2066);
nand U4066 (N_4066,N_1735,N_2377);
nand U4067 (N_4067,N_1291,N_492);
nand U4068 (N_4068,N_2156,N_511);
or U4069 (N_4069,N_896,N_2156);
nor U4070 (N_4070,N_1186,N_773);
and U4071 (N_4071,N_261,N_798);
nor U4072 (N_4072,N_906,N_931);
nor U4073 (N_4073,N_1856,N_2346);
nor U4074 (N_4074,N_305,N_2273);
nor U4075 (N_4075,N_2258,N_956);
nor U4076 (N_4076,N_1027,N_746);
nand U4077 (N_4077,N_2069,N_1136);
and U4078 (N_4078,N_385,N_595);
nor U4079 (N_4079,N_1567,N_1331);
xor U4080 (N_4080,N_343,N_1743);
xnor U4081 (N_4081,N_1864,N_2371);
nand U4082 (N_4082,N_442,N_1863);
xor U4083 (N_4083,N_123,N_1935);
and U4084 (N_4084,N_1060,N_2289);
xor U4085 (N_4085,N_1992,N_301);
nor U4086 (N_4086,N_2178,N_1641);
and U4087 (N_4087,N_1463,N_1473);
xor U4088 (N_4088,N_154,N_1379);
or U4089 (N_4089,N_2210,N_2092);
and U4090 (N_4090,N_1288,N_1972);
xnor U4091 (N_4091,N_131,N_1647);
and U4092 (N_4092,N_1189,N_368);
and U4093 (N_4093,N_1990,N_1054);
and U4094 (N_4094,N_120,N_173);
and U4095 (N_4095,N_1995,N_1649);
or U4096 (N_4096,N_360,N_56);
nand U4097 (N_4097,N_70,N_2209);
xnor U4098 (N_4098,N_1112,N_1631);
xor U4099 (N_4099,N_568,N_1067);
or U4100 (N_4100,N_731,N_1440);
xor U4101 (N_4101,N_1094,N_215);
nor U4102 (N_4102,N_1956,N_161);
nand U4103 (N_4103,N_996,N_1821);
and U4104 (N_4104,N_121,N_993);
nor U4105 (N_4105,N_2142,N_1446);
and U4106 (N_4106,N_1123,N_502);
nor U4107 (N_4107,N_2339,N_1857);
and U4108 (N_4108,N_966,N_1485);
or U4109 (N_4109,N_746,N_1828);
or U4110 (N_4110,N_2374,N_1514);
xor U4111 (N_4111,N_965,N_1402);
nor U4112 (N_4112,N_515,N_2395);
xnor U4113 (N_4113,N_2414,N_2341);
and U4114 (N_4114,N_1202,N_1453);
nand U4115 (N_4115,N_1087,N_1131);
nand U4116 (N_4116,N_2199,N_1579);
and U4117 (N_4117,N_2087,N_1310);
or U4118 (N_4118,N_562,N_2407);
nand U4119 (N_4119,N_40,N_1852);
nor U4120 (N_4120,N_1661,N_2159);
xor U4121 (N_4121,N_87,N_285);
nor U4122 (N_4122,N_1007,N_1078);
nand U4123 (N_4123,N_674,N_253);
or U4124 (N_4124,N_1570,N_795);
and U4125 (N_4125,N_1143,N_1856);
nand U4126 (N_4126,N_2462,N_21);
nor U4127 (N_4127,N_2105,N_121);
and U4128 (N_4128,N_2291,N_2391);
or U4129 (N_4129,N_667,N_1517);
nand U4130 (N_4130,N_1817,N_154);
or U4131 (N_4131,N_540,N_6);
xnor U4132 (N_4132,N_1600,N_1402);
nor U4133 (N_4133,N_523,N_1748);
nor U4134 (N_4134,N_582,N_723);
or U4135 (N_4135,N_365,N_66);
xnor U4136 (N_4136,N_906,N_2377);
nand U4137 (N_4137,N_1071,N_540);
and U4138 (N_4138,N_714,N_2295);
and U4139 (N_4139,N_983,N_194);
nand U4140 (N_4140,N_419,N_1768);
xor U4141 (N_4141,N_2300,N_186);
nand U4142 (N_4142,N_778,N_2454);
xnor U4143 (N_4143,N_680,N_769);
or U4144 (N_4144,N_1507,N_2369);
xor U4145 (N_4145,N_968,N_2166);
xnor U4146 (N_4146,N_1506,N_2358);
nand U4147 (N_4147,N_1325,N_1025);
or U4148 (N_4148,N_1016,N_1493);
and U4149 (N_4149,N_2440,N_2450);
nor U4150 (N_4150,N_1230,N_2001);
nor U4151 (N_4151,N_1148,N_1195);
nor U4152 (N_4152,N_819,N_2471);
or U4153 (N_4153,N_1320,N_1086);
xnor U4154 (N_4154,N_460,N_1963);
nor U4155 (N_4155,N_1644,N_1807);
or U4156 (N_4156,N_101,N_124);
nor U4157 (N_4157,N_747,N_496);
nor U4158 (N_4158,N_2274,N_782);
and U4159 (N_4159,N_1564,N_33);
or U4160 (N_4160,N_1552,N_1227);
and U4161 (N_4161,N_873,N_963);
xnor U4162 (N_4162,N_1853,N_1811);
nand U4163 (N_4163,N_1707,N_1131);
xnor U4164 (N_4164,N_159,N_275);
nand U4165 (N_4165,N_1991,N_1207);
or U4166 (N_4166,N_551,N_2454);
nand U4167 (N_4167,N_1451,N_27);
nand U4168 (N_4168,N_435,N_804);
and U4169 (N_4169,N_1772,N_2474);
nor U4170 (N_4170,N_2335,N_541);
nand U4171 (N_4171,N_1376,N_2137);
nor U4172 (N_4172,N_2137,N_1131);
nand U4173 (N_4173,N_2421,N_632);
or U4174 (N_4174,N_2496,N_1363);
nand U4175 (N_4175,N_2476,N_1866);
nand U4176 (N_4176,N_51,N_1878);
xor U4177 (N_4177,N_346,N_328);
or U4178 (N_4178,N_269,N_365);
xor U4179 (N_4179,N_1467,N_633);
nand U4180 (N_4180,N_1262,N_1943);
or U4181 (N_4181,N_1517,N_1032);
or U4182 (N_4182,N_1400,N_527);
or U4183 (N_4183,N_1509,N_1444);
and U4184 (N_4184,N_514,N_1577);
xnor U4185 (N_4185,N_1034,N_633);
nand U4186 (N_4186,N_616,N_640);
or U4187 (N_4187,N_1025,N_2138);
nor U4188 (N_4188,N_1847,N_2381);
nand U4189 (N_4189,N_1490,N_1780);
xnor U4190 (N_4190,N_432,N_516);
nand U4191 (N_4191,N_679,N_2119);
nor U4192 (N_4192,N_1075,N_1629);
and U4193 (N_4193,N_597,N_234);
nand U4194 (N_4194,N_2181,N_1020);
or U4195 (N_4195,N_1543,N_2066);
xnor U4196 (N_4196,N_376,N_862);
or U4197 (N_4197,N_1100,N_1506);
and U4198 (N_4198,N_192,N_903);
nand U4199 (N_4199,N_2325,N_2337);
and U4200 (N_4200,N_1033,N_2294);
and U4201 (N_4201,N_221,N_1765);
and U4202 (N_4202,N_2,N_991);
and U4203 (N_4203,N_2344,N_338);
nor U4204 (N_4204,N_1469,N_2409);
nand U4205 (N_4205,N_955,N_715);
xnor U4206 (N_4206,N_1999,N_1912);
nand U4207 (N_4207,N_2168,N_2484);
nand U4208 (N_4208,N_331,N_489);
and U4209 (N_4209,N_560,N_663);
nand U4210 (N_4210,N_2199,N_524);
nand U4211 (N_4211,N_791,N_2140);
nand U4212 (N_4212,N_1288,N_487);
nor U4213 (N_4213,N_152,N_630);
nor U4214 (N_4214,N_720,N_2108);
and U4215 (N_4215,N_1874,N_2414);
nor U4216 (N_4216,N_1689,N_416);
nand U4217 (N_4217,N_2288,N_1423);
xor U4218 (N_4218,N_1724,N_442);
xnor U4219 (N_4219,N_519,N_1220);
xor U4220 (N_4220,N_714,N_1573);
nand U4221 (N_4221,N_2325,N_1704);
and U4222 (N_4222,N_2344,N_96);
or U4223 (N_4223,N_1225,N_1761);
xor U4224 (N_4224,N_341,N_1173);
xnor U4225 (N_4225,N_1378,N_1089);
nand U4226 (N_4226,N_665,N_24);
nand U4227 (N_4227,N_37,N_1076);
nand U4228 (N_4228,N_1389,N_2059);
or U4229 (N_4229,N_1558,N_149);
and U4230 (N_4230,N_1204,N_1511);
nor U4231 (N_4231,N_1444,N_1896);
or U4232 (N_4232,N_1914,N_668);
nor U4233 (N_4233,N_227,N_2132);
and U4234 (N_4234,N_679,N_193);
and U4235 (N_4235,N_470,N_1904);
and U4236 (N_4236,N_281,N_2023);
nand U4237 (N_4237,N_1897,N_321);
nand U4238 (N_4238,N_1495,N_2067);
xor U4239 (N_4239,N_2177,N_1515);
xnor U4240 (N_4240,N_139,N_2365);
nor U4241 (N_4241,N_954,N_1766);
xor U4242 (N_4242,N_860,N_157);
or U4243 (N_4243,N_71,N_17);
or U4244 (N_4244,N_808,N_2451);
or U4245 (N_4245,N_2290,N_1625);
or U4246 (N_4246,N_730,N_305);
or U4247 (N_4247,N_293,N_827);
xnor U4248 (N_4248,N_1338,N_377);
and U4249 (N_4249,N_2000,N_135);
xnor U4250 (N_4250,N_1756,N_1592);
nand U4251 (N_4251,N_1416,N_1146);
or U4252 (N_4252,N_568,N_1550);
nand U4253 (N_4253,N_1171,N_1882);
nor U4254 (N_4254,N_142,N_1121);
or U4255 (N_4255,N_2426,N_651);
and U4256 (N_4256,N_1755,N_2407);
and U4257 (N_4257,N_134,N_1768);
or U4258 (N_4258,N_1734,N_1389);
xor U4259 (N_4259,N_850,N_1354);
and U4260 (N_4260,N_2218,N_322);
nor U4261 (N_4261,N_383,N_507);
and U4262 (N_4262,N_955,N_845);
and U4263 (N_4263,N_795,N_1761);
xor U4264 (N_4264,N_1928,N_1712);
nand U4265 (N_4265,N_66,N_906);
nor U4266 (N_4266,N_1247,N_1836);
and U4267 (N_4267,N_408,N_899);
or U4268 (N_4268,N_1931,N_2420);
or U4269 (N_4269,N_2322,N_2210);
nor U4270 (N_4270,N_2319,N_1150);
nand U4271 (N_4271,N_249,N_1485);
or U4272 (N_4272,N_1425,N_1078);
nor U4273 (N_4273,N_412,N_2361);
xnor U4274 (N_4274,N_8,N_1944);
or U4275 (N_4275,N_53,N_2362);
nor U4276 (N_4276,N_1863,N_950);
nand U4277 (N_4277,N_2354,N_1931);
nand U4278 (N_4278,N_97,N_1829);
nor U4279 (N_4279,N_273,N_643);
nor U4280 (N_4280,N_1260,N_380);
and U4281 (N_4281,N_1284,N_1727);
xnor U4282 (N_4282,N_719,N_1900);
and U4283 (N_4283,N_378,N_572);
nand U4284 (N_4284,N_1681,N_1177);
and U4285 (N_4285,N_195,N_1955);
nand U4286 (N_4286,N_195,N_1287);
nor U4287 (N_4287,N_743,N_1446);
or U4288 (N_4288,N_204,N_1684);
or U4289 (N_4289,N_1899,N_1584);
or U4290 (N_4290,N_82,N_1498);
and U4291 (N_4291,N_2152,N_656);
xnor U4292 (N_4292,N_129,N_847);
and U4293 (N_4293,N_1738,N_32);
or U4294 (N_4294,N_144,N_350);
and U4295 (N_4295,N_1348,N_282);
xor U4296 (N_4296,N_1339,N_662);
nand U4297 (N_4297,N_2452,N_1381);
or U4298 (N_4298,N_370,N_1044);
xor U4299 (N_4299,N_322,N_2188);
xor U4300 (N_4300,N_1659,N_491);
or U4301 (N_4301,N_659,N_476);
or U4302 (N_4302,N_582,N_832);
nor U4303 (N_4303,N_231,N_545);
nor U4304 (N_4304,N_136,N_284);
and U4305 (N_4305,N_523,N_3);
and U4306 (N_4306,N_1116,N_1956);
and U4307 (N_4307,N_579,N_1562);
or U4308 (N_4308,N_1253,N_2109);
and U4309 (N_4309,N_1081,N_70);
nor U4310 (N_4310,N_243,N_1032);
nor U4311 (N_4311,N_1461,N_88);
nand U4312 (N_4312,N_785,N_2198);
nor U4313 (N_4313,N_1480,N_847);
nor U4314 (N_4314,N_839,N_1878);
and U4315 (N_4315,N_1831,N_1148);
or U4316 (N_4316,N_769,N_390);
nand U4317 (N_4317,N_67,N_2345);
nor U4318 (N_4318,N_2071,N_316);
and U4319 (N_4319,N_861,N_791);
and U4320 (N_4320,N_635,N_2282);
or U4321 (N_4321,N_1257,N_1001);
or U4322 (N_4322,N_1593,N_364);
or U4323 (N_4323,N_1911,N_1752);
nor U4324 (N_4324,N_1147,N_267);
nor U4325 (N_4325,N_766,N_1350);
or U4326 (N_4326,N_1905,N_2038);
xnor U4327 (N_4327,N_1060,N_715);
xnor U4328 (N_4328,N_1903,N_1383);
nor U4329 (N_4329,N_996,N_1854);
or U4330 (N_4330,N_1873,N_1583);
and U4331 (N_4331,N_385,N_432);
and U4332 (N_4332,N_1913,N_90);
and U4333 (N_4333,N_930,N_429);
nor U4334 (N_4334,N_2165,N_1485);
nor U4335 (N_4335,N_1856,N_2453);
or U4336 (N_4336,N_2153,N_838);
or U4337 (N_4337,N_1755,N_1733);
nor U4338 (N_4338,N_196,N_1234);
and U4339 (N_4339,N_72,N_1801);
nand U4340 (N_4340,N_1206,N_2274);
nand U4341 (N_4341,N_992,N_1256);
and U4342 (N_4342,N_2078,N_1439);
nor U4343 (N_4343,N_763,N_1747);
or U4344 (N_4344,N_769,N_2360);
nor U4345 (N_4345,N_1324,N_2288);
nor U4346 (N_4346,N_641,N_620);
and U4347 (N_4347,N_562,N_2205);
nand U4348 (N_4348,N_313,N_1860);
and U4349 (N_4349,N_702,N_1450);
and U4350 (N_4350,N_851,N_1157);
and U4351 (N_4351,N_214,N_1757);
nor U4352 (N_4352,N_2251,N_944);
and U4353 (N_4353,N_1577,N_1415);
nand U4354 (N_4354,N_1059,N_552);
xor U4355 (N_4355,N_806,N_2270);
or U4356 (N_4356,N_739,N_386);
and U4357 (N_4357,N_2367,N_939);
and U4358 (N_4358,N_2007,N_2425);
and U4359 (N_4359,N_2336,N_1447);
nor U4360 (N_4360,N_1105,N_828);
nand U4361 (N_4361,N_2452,N_265);
xor U4362 (N_4362,N_2482,N_1981);
or U4363 (N_4363,N_346,N_1989);
and U4364 (N_4364,N_500,N_2106);
nand U4365 (N_4365,N_1752,N_529);
or U4366 (N_4366,N_1114,N_111);
and U4367 (N_4367,N_2129,N_487);
xor U4368 (N_4368,N_643,N_2155);
xor U4369 (N_4369,N_865,N_886);
and U4370 (N_4370,N_981,N_1361);
nand U4371 (N_4371,N_170,N_1213);
nor U4372 (N_4372,N_2106,N_2387);
or U4373 (N_4373,N_396,N_965);
nor U4374 (N_4374,N_1879,N_358);
nor U4375 (N_4375,N_261,N_431);
nand U4376 (N_4376,N_2219,N_415);
and U4377 (N_4377,N_1565,N_1248);
or U4378 (N_4378,N_2078,N_1569);
nand U4379 (N_4379,N_1134,N_1407);
nor U4380 (N_4380,N_1921,N_627);
xor U4381 (N_4381,N_2417,N_7);
xor U4382 (N_4382,N_60,N_1121);
nor U4383 (N_4383,N_2273,N_2176);
xnor U4384 (N_4384,N_908,N_1818);
and U4385 (N_4385,N_2422,N_2436);
xor U4386 (N_4386,N_2226,N_2111);
or U4387 (N_4387,N_751,N_808);
nor U4388 (N_4388,N_579,N_1073);
xor U4389 (N_4389,N_1688,N_411);
xor U4390 (N_4390,N_2494,N_296);
and U4391 (N_4391,N_1264,N_105);
or U4392 (N_4392,N_585,N_129);
or U4393 (N_4393,N_287,N_551);
nor U4394 (N_4394,N_1615,N_2137);
and U4395 (N_4395,N_1136,N_397);
and U4396 (N_4396,N_482,N_191);
nor U4397 (N_4397,N_1856,N_1913);
and U4398 (N_4398,N_679,N_1908);
nand U4399 (N_4399,N_1354,N_1936);
nor U4400 (N_4400,N_1405,N_2329);
xor U4401 (N_4401,N_1919,N_1949);
nor U4402 (N_4402,N_156,N_1603);
nor U4403 (N_4403,N_1236,N_933);
nor U4404 (N_4404,N_2481,N_103);
or U4405 (N_4405,N_1868,N_1787);
nor U4406 (N_4406,N_1089,N_2258);
nand U4407 (N_4407,N_1557,N_2348);
nor U4408 (N_4408,N_2428,N_2094);
xor U4409 (N_4409,N_1792,N_52);
or U4410 (N_4410,N_247,N_1198);
nor U4411 (N_4411,N_1620,N_1);
xor U4412 (N_4412,N_1040,N_817);
and U4413 (N_4413,N_1659,N_1596);
or U4414 (N_4414,N_415,N_2180);
nor U4415 (N_4415,N_2344,N_753);
xor U4416 (N_4416,N_652,N_349);
xor U4417 (N_4417,N_79,N_204);
nand U4418 (N_4418,N_673,N_1953);
and U4419 (N_4419,N_2484,N_2009);
nand U4420 (N_4420,N_1486,N_1330);
and U4421 (N_4421,N_101,N_472);
and U4422 (N_4422,N_1430,N_1516);
nand U4423 (N_4423,N_1089,N_2354);
nand U4424 (N_4424,N_1918,N_501);
xnor U4425 (N_4425,N_328,N_911);
xnor U4426 (N_4426,N_2388,N_736);
xor U4427 (N_4427,N_981,N_1822);
or U4428 (N_4428,N_1007,N_1403);
nand U4429 (N_4429,N_1182,N_1109);
or U4430 (N_4430,N_699,N_362);
nor U4431 (N_4431,N_867,N_898);
xnor U4432 (N_4432,N_886,N_2064);
nand U4433 (N_4433,N_86,N_849);
xnor U4434 (N_4434,N_1391,N_2373);
nand U4435 (N_4435,N_1823,N_680);
and U4436 (N_4436,N_1252,N_1520);
nand U4437 (N_4437,N_1676,N_1981);
nand U4438 (N_4438,N_502,N_1667);
or U4439 (N_4439,N_1668,N_2073);
xnor U4440 (N_4440,N_719,N_585);
and U4441 (N_4441,N_680,N_1716);
and U4442 (N_4442,N_798,N_306);
nand U4443 (N_4443,N_1765,N_1639);
xor U4444 (N_4444,N_2374,N_1340);
nor U4445 (N_4445,N_1392,N_340);
and U4446 (N_4446,N_2126,N_904);
and U4447 (N_4447,N_899,N_448);
and U4448 (N_4448,N_2109,N_1450);
or U4449 (N_4449,N_1052,N_1212);
xnor U4450 (N_4450,N_2048,N_1823);
xnor U4451 (N_4451,N_648,N_1119);
and U4452 (N_4452,N_2376,N_1034);
xnor U4453 (N_4453,N_981,N_2392);
nand U4454 (N_4454,N_378,N_12);
or U4455 (N_4455,N_2447,N_1119);
xor U4456 (N_4456,N_1097,N_1784);
and U4457 (N_4457,N_1928,N_405);
or U4458 (N_4458,N_1665,N_2063);
nor U4459 (N_4459,N_321,N_2);
nor U4460 (N_4460,N_2181,N_1936);
nor U4461 (N_4461,N_1325,N_2005);
and U4462 (N_4462,N_585,N_909);
xnor U4463 (N_4463,N_992,N_2029);
nand U4464 (N_4464,N_2456,N_2194);
xor U4465 (N_4465,N_2477,N_22);
xnor U4466 (N_4466,N_2482,N_1924);
nor U4467 (N_4467,N_1653,N_2257);
or U4468 (N_4468,N_842,N_1317);
nand U4469 (N_4469,N_747,N_2344);
or U4470 (N_4470,N_838,N_2221);
nor U4471 (N_4471,N_23,N_173);
or U4472 (N_4472,N_2100,N_502);
nand U4473 (N_4473,N_983,N_1348);
and U4474 (N_4474,N_1742,N_626);
or U4475 (N_4475,N_2487,N_299);
nor U4476 (N_4476,N_1409,N_1516);
xnor U4477 (N_4477,N_2002,N_404);
xor U4478 (N_4478,N_2450,N_230);
or U4479 (N_4479,N_760,N_437);
nor U4480 (N_4480,N_1391,N_1700);
nor U4481 (N_4481,N_1280,N_240);
nor U4482 (N_4482,N_979,N_626);
and U4483 (N_4483,N_1795,N_676);
or U4484 (N_4484,N_2289,N_1577);
xor U4485 (N_4485,N_850,N_377);
nand U4486 (N_4486,N_117,N_1090);
and U4487 (N_4487,N_1227,N_2053);
nor U4488 (N_4488,N_1389,N_1288);
or U4489 (N_4489,N_1267,N_744);
or U4490 (N_4490,N_2466,N_897);
xor U4491 (N_4491,N_2094,N_2036);
nand U4492 (N_4492,N_1969,N_1618);
xor U4493 (N_4493,N_743,N_1363);
or U4494 (N_4494,N_430,N_1987);
and U4495 (N_4495,N_1844,N_471);
nand U4496 (N_4496,N_2176,N_845);
nand U4497 (N_4497,N_1425,N_1208);
xnor U4498 (N_4498,N_2215,N_1459);
nor U4499 (N_4499,N_2487,N_1145);
xor U4500 (N_4500,N_503,N_1925);
xnor U4501 (N_4501,N_293,N_1982);
nand U4502 (N_4502,N_908,N_2352);
xor U4503 (N_4503,N_1498,N_1071);
or U4504 (N_4504,N_590,N_1923);
nor U4505 (N_4505,N_2010,N_1608);
nor U4506 (N_4506,N_31,N_132);
or U4507 (N_4507,N_407,N_2455);
xor U4508 (N_4508,N_695,N_125);
nand U4509 (N_4509,N_1614,N_358);
xnor U4510 (N_4510,N_1919,N_2442);
nand U4511 (N_4511,N_144,N_1546);
or U4512 (N_4512,N_332,N_125);
nand U4513 (N_4513,N_1176,N_1414);
xnor U4514 (N_4514,N_1803,N_1711);
nor U4515 (N_4515,N_26,N_437);
nand U4516 (N_4516,N_1064,N_2229);
nand U4517 (N_4517,N_782,N_1122);
or U4518 (N_4518,N_1193,N_2089);
and U4519 (N_4519,N_548,N_619);
nand U4520 (N_4520,N_1714,N_1899);
or U4521 (N_4521,N_549,N_669);
nand U4522 (N_4522,N_2341,N_2024);
nor U4523 (N_4523,N_1022,N_1771);
nand U4524 (N_4524,N_1904,N_2189);
and U4525 (N_4525,N_514,N_394);
and U4526 (N_4526,N_703,N_931);
and U4527 (N_4527,N_372,N_27);
nor U4528 (N_4528,N_2254,N_1276);
and U4529 (N_4529,N_587,N_2355);
nand U4530 (N_4530,N_680,N_579);
and U4531 (N_4531,N_1147,N_283);
nand U4532 (N_4532,N_949,N_82);
nor U4533 (N_4533,N_670,N_1295);
or U4534 (N_4534,N_2472,N_2122);
xor U4535 (N_4535,N_2073,N_947);
nand U4536 (N_4536,N_1765,N_2349);
or U4537 (N_4537,N_215,N_377);
or U4538 (N_4538,N_1094,N_47);
xor U4539 (N_4539,N_1666,N_974);
nor U4540 (N_4540,N_2459,N_428);
nor U4541 (N_4541,N_1011,N_814);
nor U4542 (N_4542,N_121,N_867);
nand U4543 (N_4543,N_2248,N_376);
or U4544 (N_4544,N_2383,N_354);
or U4545 (N_4545,N_2485,N_312);
nand U4546 (N_4546,N_384,N_2170);
nor U4547 (N_4547,N_2439,N_2042);
or U4548 (N_4548,N_1345,N_2192);
and U4549 (N_4549,N_1012,N_536);
nand U4550 (N_4550,N_1393,N_1904);
nand U4551 (N_4551,N_885,N_1532);
and U4552 (N_4552,N_1405,N_1588);
nand U4553 (N_4553,N_817,N_1495);
xor U4554 (N_4554,N_351,N_127);
xor U4555 (N_4555,N_338,N_2439);
nor U4556 (N_4556,N_992,N_637);
nor U4557 (N_4557,N_1232,N_1797);
or U4558 (N_4558,N_231,N_2136);
nand U4559 (N_4559,N_350,N_1300);
and U4560 (N_4560,N_1939,N_376);
or U4561 (N_4561,N_2278,N_821);
nor U4562 (N_4562,N_286,N_1818);
or U4563 (N_4563,N_1528,N_2495);
and U4564 (N_4564,N_385,N_500);
and U4565 (N_4565,N_2178,N_1995);
nand U4566 (N_4566,N_1360,N_2499);
and U4567 (N_4567,N_1452,N_840);
nand U4568 (N_4568,N_304,N_566);
or U4569 (N_4569,N_1836,N_2455);
or U4570 (N_4570,N_504,N_41);
nand U4571 (N_4571,N_659,N_2240);
xnor U4572 (N_4572,N_2235,N_2257);
nor U4573 (N_4573,N_1669,N_417);
nand U4574 (N_4574,N_1053,N_918);
nor U4575 (N_4575,N_1352,N_1338);
and U4576 (N_4576,N_1666,N_506);
or U4577 (N_4577,N_1818,N_739);
nand U4578 (N_4578,N_266,N_1648);
nor U4579 (N_4579,N_2422,N_1622);
xor U4580 (N_4580,N_1449,N_1786);
xor U4581 (N_4581,N_170,N_1030);
xnor U4582 (N_4582,N_492,N_924);
xnor U4583 (N_4583,N_1572,N_674);
and U4584 (N_4584,N_39,N_2151);
xnor U4585 (N_4585,N_1315,N_1805);
and U4586 (N_4586,N_857,N_1722);
and U4587 (N_4587,N_1870,N_1319);
nor U4588 (N_4588,N_204,N_1750);
nand U4589 (N_4589,N_2313,N_1484);
nand U4590 (N_4590,N_2005,N_1237);
and U4591 (N_4591,N_1969,N_218);
xor U4592 (N_4592,N_294,N_327);
xor U4593 (N_4593,N_1173,N_2359);
and U4594 (N_4594,N_485,N_881);
xor U4595 (N_4595,N_446,N_673);
and U4596 (N_4596,N_1849,N_776);
and U4597 (N_4597,N_1247,N_1675);
nand U4598 (N_4598,N_1845,N_2182);
xnor U4599 (N_4599,N_366,N_1983);
nand U4600 (N_4600,N_1763,N_77);
nor U4601 (N_4601,N_1472,N_1458);
nand U4602 (N_4602,N_1729,N_1502);
nand U4603 (N_4603,N_424,N_864);
and U4604 (N_4604,N_1643,N_2205);
nor U4605 (N_4605,N_2457,N_2184);
nor U4606 (N_4606,N_508,N_892);
or U4607 (N_4607,N_2107,N_1970);
nor U4608 (N_4608,N_741,N_2192);
nor U4609 (N_4609,N_545,N_1544);
nand U4610 (N_4610,N_783,N_1946);
or U4611 (N_4611,N_243,N_2098);
xnor U4612 (N_4612,N_1091,N_1242);
nand U4613 (N_4613,N_2381,N_1605);
nor U4614 (N_4614,N_664,N_1507);
and U4615 (N_4615,N_2067,N_2339);
xnor U4616 (N_4616,N_457,N_1279);
xor U4617 (N_4617,N_693,N_2020);
xnor U4618 (N_4618,N_2135,N_1875);
or U4619 (N_4619,N_3,N_111);
or U4620 (N_4620,N_667,N_115);
nor U4621 (N_4621,N_615,N_591);
nor U4622 (N_4622,N_542,N_1938);
nand U4623 (N_4623,N_159,N_560);
nand U4624 (N_4624,N_2188,N_1131);
nor U4625 (N_4625,N_1682,N_383);
and U4626 (N_4626,N_1370,N_1745);
nand U4627 (N_4627,N_1504,N_1539);
or U4628 (N_4628,N_2088,N_2185);
or U4629 (N_4629,N_366,N_1369);
and U4630 (N_4630,N_1044,N_2095);
or U4631 (N_4631,N_823,N_2044);
or U4632 (N_4632,N_2072,N_2150);
xnor U4633 (N_4633,N_1028,N_2058);
nor U4634 (N_4634,N_2307,N_669);
nand U4635 (N_4635,N_2048,N_1592);
or U4636 (N_4636,N_1437,N_2421);
xor U4637 (N_4637,N_1532,N_1346);
nand U4638 (N_4638,N_2202,N_209);
nor U4639 (N_4639,N_407,N_4);
or U4640 (N_4640,N_1792,N_2494);
nand U4641 (N_4641,N_1888,N_1653);
xnor U4642 (N_4642,N_2074,N_1104);
and U4643 (N_4643,N_1699,N_493);
or U4644 (N_4644,N_947,N_297);
nand U4645 (N_4645,N_1655,N_687);
nand U4646 (N_4646,N_2156,N_945);
or U4647 (N_4647,N_2139,N_929);
xor U4648 (N_4648,N_2409,N_436);
and U4649 (N_4649,N_883,N_127);
or U4650 (N_4650,N_1745,N_1055);
nand U4651 (N_4651,N_1298,N_2364);
and U4652 (N_4652,N_1426,N_1158);
or U4653 (N_4653,N_227,N_2477);
or U4654 (N_4654,N_1376,N_1129);
or U4655 (N_4655,N_356,N_255);
and U4656 (N_4656,N_1205,N_2397);
xor U4657 (N_4657,N_269,N_201);
nor U4658 (N_4658,N_77,N_225);
or U4659 (N_4659,N_678,N_1710);
nand U4660 (N_4660,N_2430,N_1418);
nor U4661 (N_4661,N_1130,N_954);
xnor U4662 (N_4662,N_92,N_796);
xor U4663 (N_4663,N_1272,N_1402);
nand U4664 (N_4664,N_577,N_1497);
xor U4665 (N_4665,N_1818,N_1677);
xor U4666 (N_4666,N_1499,N_186);
and U4667 (N_4667,N_2214,N_1643);
xor U4668 (N_4668,N_2084,N_471);
or U4669 (N_4669,N_78,N_2485);
and U4670 (N_4670,N_1908,N_1654);
or U4671 (N_4671,N_928,N_205);
xor U4672 (N_4672,N_1805,N_540);
or U4673 (N_4673,N_652,N_1512);
and U4674 (N_4674,N_1599,N_659);
nor U4675 (N_4675,N_82,N_427);
nand U4676 (N_4676,N_1377,N_49);
or U4677 (N_4677,N_1151,N_1171);
xor U4678 (N_4678,N_1720,N_521);
nand U4679 (N_4679,N_2372,N_759);
nor U4680 (N_4680,N_1847,N_1264);
or U4681 (N_4681,N_1248,N_2132);
xor U4682 (N_4682,N_276,N_4);
xor U4683 (N_4683,N_1047,N_127);
or U4684 (N_4684,N_294,N_389);
nor U4685 (N_4685,N_34,N_1080);
or U4686 (N_4686,N_704,N_1448);
xnor U4687 (N_4687,N_969,N_2435);
nand U4688 (N_4688,N_1253,N_80);
or U4689 (N_4689,N_1504,N_2408);
nand U4690 (N_4690,N_774,N_767);
xnor U4691 (N_4691,N_1787,N_2297);
nor U4692 (N_4692,N_1775,N_50);
and U4693 (N_4693,N_935,N_1654);
xnor U4694 (N_4694,N_577,N_941);
xnor U4695 (N_4695,N_503,N_2331);
or U4696 (N_4696,N_1854,N_2040);
xnor U4697 (N_4697,N_145,N_290);
or U4698 (N_4698,N_1438,N_361);
nor U4699 (N_4699,N_2072,N_1039);
or U4700 (N_4700,N_833,N_1645);
xor U4701 (N_4701,N_363,N_1211);
nor U4702 (N_4702,N_855,N_1472);
or U4703 (N_4703,N_652,N_1417);
nand U4704 (N_4704,N_2022,N_132);
and U4705 (N_4705,N_285,N_1247);
and U4706 (N_4706,N_2344,N_1143);
xnor U4707 (N_4707,N_442,N_1044);
nor U4708 (N_4708,N_2230,N_557);
nor U4709 (N_4709,N_19,N_1446);
and U4710 (N_4710,N_168,N_51);
xor U4711 (N_4711,N_2143,N_534);
nand U4712 (N_4712,N_1162,N_137);
or U4713 (N_4713,N_925,N_431);
or U4714 (N_4714,N_1144,N_102);
or U4715 (N_4715,N_599,N_229);
nand U4716 (N_4716,N_686,N_2442);
nor U4717 (N_4717,N_486,N_938);
and U4718 (N_4718,N_2013,N_2286);
nand U4719 (N_4719,N_464,N_694);
nor U4720 (N_4720,N_245,N_367);
nor U4721 (N_4721,N_2270,N_1569);
nand U4722 (N_4722,N_1940,N_2352);
nand U4723 (N_4723,N_1783,N_1826);
or U4724 (N_4724,N_271,N_1039);
or U4725 (N_4725,N_2436,N_2409);
nand U4726 (N_4726,N_2020,N_257);
or U4727 (N_4727,N_736,N_2144);
xor U4728 (N_4728,N_1308,N_1296);
nand U4729 (N_4729,N_1416,N_1982);
or U4730 (N_4730,N_1378,N_244);
nor U4731 (N_4731,N_2029,N_2326);
nand U4732 (N_4732,N_2134,N_152);
xor U4733 (N_4733,N_876,N_1731);
or U4734 (N_4734,N_1307,N_2005);
or U4735 (N_4735,N_2462,N_1174);
nand U4736 (N_4736,N_1090,N_1848);
nand U4737 (N_4737,N_1263,N_1058);
xor U4738 (N_4738,N_383,N_862);
nor U4739 (N_4739,N_475,N_1951);
nor U4740 (N_4740,N_1914,N_302);
xnor U4741 (N_4741,N_1844,N_698);
nor U4742 (N_4742,N_1732,N_1649);
or U4743 (N_4743,N_195,N_395);
nand U4744 (N_4744,N_1191,N_202);
xnor U4745 (N_4745,N_1898,N_2392);
or U4746 (N_4746,N_971,N_161);
and U4747 (N_4747,N_1564,N_1279);
nor U4748 (N_4748,N_1344,N_325);
nor U4749 (N_4749,N_1197,N_2165);
nor U4750 (N_4750,N_1538,N_1026);
or U4751 (N_4751,N_1004,N_118);
or U4752 (N_4752,N_919,N_816);
or U4753 (N_4753,N_1892,N_2370);
and U4754 (N_4754,N_747,N_659);
xnor U4755 (N_4755,N_1210,N_1996);
and U4756 (N_4756,N_407,N_1429);
xnor U4757 (N_4757,N_446,N_1787);
nand U4758 (N_4758,N_344,N_1122);
xor U4759 (N_4759,N_972,N_630);
xnor U4760 (N_4760,N_626,N_935);
nand U4761 (N_4761,N_1937,N_1855);
nand U4762 (N_4762,N_2092,N_1602);
or U4763 (N_4763,N_1033,N_436);
xnor U4764 (N_4764,N_1666,N_1577);
or U4765 (N_4765,N_1745,N_920);
nor U4766 (N_4766,N_1713,N_1681);
and U4767 (N_4767,N_1218,N_1452);
or U4768 (N_4768,N_1855,N_462);
xor U4769 (N_4769,N_112,N_1401);
nor U4770 (N_4770,N_595,N_1067);
nand U4771 (N_4771,N_180,N_67);
nor U4772 (N_4772,N_1749,N_1227);
nand U4773 (N_4773,N_1095,N_792);
xor U4774 (N_4774,N_1154,N_1622);
and U4775 (N_4775,N_288,N_1121);
nand U4776 (N_4776,N_1466,N_546);
and U4777 (N_4777,N_1424,N_1989);
nor U4778 (N_4778,N_1208,N_1063);
nand U4779 (N_4779,N_1883,N_530);
and U4780 (N_4780,N_335,N_1273);
nand U4781 (N_4781,N_2245,N_0);
or U4782 (N_4782,N_204,N_2365);
xnor U4783 (N_4783,N_2403,N_1075);
or U4784 (N_4784,N_1180,N_848);
or U4785 (N_4785,N_221,N_964);
nor U4786 (N_4786,N_1461,N_1386);
nand U4787 (N_4787,N_1079,N_2152);
or U4788 (N_4788,N_1696,N_373);
nand U4789 (N_4789,N_2127,N_24);
nor U4790 (N_4790,N_2177,N_78);
and U4791 (N_4791,N_1455,N_397);
and U4792 (N_4792,N_972,N_241);
xor U4793 (N_4793,N_1320,N_2019);
and U4794 (N_4794,N_1814,N_1870);
nand U4795 (N_4795,N_396,N_1213);
nand U4796 (N_4796,N_2224,N_266);
nand U4797 (N_4797,N_2197,N_1664);
or U4798 (N_4798,N_514,N_1759);
nand U4799 (N_4799,N_802,N_361);
nor U4800 (N_4800,N_347,N_1221);
or U4801 (N_4801,N_1644,N_864);
nor U4802 (N_4802,N_2495,N_1499);
nor U4803 (N_4803,N_273,N_289);
nand U4804 (N_4804,N_1881,N_1286);
or U4805 (N_4805,N_645,N_542);
xnor U4806 (N_4806,N_294,N_966);
nor U4807 (N_4807,N_1071,N_222);
nand U4808 (N_4808,N_1135,N_1262);
or U4809 (N_4809,N_551,N_697);
nor U4810 (N_4810,N_1159,N_2134);
or U4811 (N_4811,N_1535,N_1798);
nor U4812 (N_4812,N_1867,N_1887);
or U4813 (N_4813,N_475,N_678);
nor U4814 (N_4814,N_2215,N_1339);
and U4815 (N_4815,N_1640,N_142);
or U4816 (N_4816,N_965,N_282);
nand U4817 (N_4817,N_2112,N_1292);
and U4818 (N_4818,N_10,N_369);
or U4819 (N_4819,N_1996,N_1357);
nor U4820 (N_4820,N_1513,N_1598);
or U4821 (N_4821,N_1730,N_1466);
and U4822 (N_4822,N_175,N_1419);
or U4823 (N_4823,N_1885,N_1353);
and U4824 (N_4824,N_723,N_369);
and U4825 (N_4825,N_1633,N_1243);
nand U4826 (N_4826,N_1352,N_2301);
and U4827 (N_4827,N_56,N_2239);
and U4828 (N_4828,N_872,N_1244);
and U4829 (N_4829,N_2255,N_1876);
and U4830 (N_4830,N_1353,N_2466);
xor U4831 (N_4831,N_44,N_2024);
nor U4832 (N_4832,N_1359,N_63);
nand U4833 (N_4833,N_370,N_2086);
or U4834 (N_4834,N_777,N_361);
and U4835 (N_4835,N_722,N_2145);
or U4836 (N_4836,N_1101,N_2077);
nand U4837 (N_4837,N_784,N_1207);
nor U4838 (N_4838,N_555,N_1394);
nor U4839 (N_4839,N_2375,N_52);
and U4840 (N_4840,N_2270,N_1519);
or U4841 (N_4841,N_944,N_780);
or U4842 (N_4842,N_2486,N_2109);
nor U4843 (N_4843,N_2217,N_2058);
xnor U4844 (N_4844,N_300,N_1709);
nor U4845 (N_4845,N_1883,N_2230);
or U4846 (N_4846,N_577,N_2239);
nand U4847 (N_4847,N_1864,N_1204);
nand U4848 (N_4848,N_2322,N_2074);
or U4849 (N_4849,N_960,N_1940);
nor U4850 (N_4850,N_2405,N_1086);
xor U4851 (N_4851,N_2267,N_1341);
xnor U4852 (N_4852,N_2280,N_62);
and U4853 (N_4853,N_1262,N_668);
nand U4854 (N_4854,N_923,N_1266);
and U4855 (N_4855,N_2411,N_1518);
and U4856 (N_4856,N_2154,N_160);
and U4857 (N_4857,N_768,N_1310);
nand U4858 (N_4858,N_1736,N_2360);
nor U4859 (N_4859,N_1837,N_275);
and U4860 (N_4860,N_2466,N_1680);
xor U4861 (N_4861,N_717,N_264);
nor U4862 (N_4862,N_522,N_1745);
and U4863 (N_4863,N_1260,N_102);
nor U4864 (N_4864,N_1971,N_312);
or U4865 (N_4865,N_8,N_1806);
nor U4866 (N_4866,N_2244,N_1327);
xnor U4867 (N_4867,N_89,N_789);
and U4868 (N_4868,N_1766,N_2139);
xnor U4869 (N_4869,N_999,N_835);
nor U4870 (N_4870,N_463,N_484);
xnor U4871 (N_4871,N_1504,N_586);
nor U4872 (N_4872,N_1899,N_1778);
or U4873 (N_4873,N_985,N_903);
or U4874 (N_4874,N_1508,N_2427);
nand U4875 (N_4875,N_598,N_1471);
nand U4876 (N_4876,N_1134,N_2032);
nand U4877 (N_4877,N_1657,N_837);
and U4878 (N_4878,N_258,N_1587);
nor U4879 (N_4879,N_1199,N_804);
or U4880 (N_4880,N_1126,N_1989);
nand U4881 (N_4881,N_756,N_1911);
and U4882 (N_4882,N_835,N_502);
or U4883 (N_4883,N_295,N_166);
and U4884 (N_4884,N_300,N_1052);
xnor U4885 (N_4885,N_1573,N_1930);
or U4886 (N_4886,N_316,N_486);
nor U4887 (N_4887,N_491,N_2120);
nor U4888 (N_4888,N_2064,N_2381);
xnor U4889 (N_4889,N_2259,N_1101);
and U4890 (N_4890,N_130,N_1529);
nand U4891 (N_4891,N_51,N_613);
nor U4892 (N_4892,N_2289,N_636);
nor U4893 (N_4893,N_406,N_1790);
xnor U4894 (N_4894,N_1707,N_2016);
or U4895 (N_4895,N_868,N_113);
nand U4896 (N_4896,N_2071,N_337);
nand U4897 (N_4897,N_1567,N_1160);
xor U4898 (N_4898,N_862,N_1006);
nor U4899 (N_4899,N_1351,N_834);
or U4900 (N_4900,N_1798,N_1165);
and U4901 (N_4901,N_1839,N_1312);
nand U4902 (N_4902,N_380,N_1548);
nand U4903 (N_4903,N_1035,N_2088);
nand U4904 (N_4904,N_1733,N_986);
and U4905 (N_4905,N_1696,N_2289);
nand U4906 (N_4906,N_2489,N_194);
or U4907 (N_4907,N_1011,N_359);
xor U4908 (N_4908,N_108,N_2133);
and U4909 (N_4909,N_496,N_364);
or U4910 (N_4910,N_2217,N_484);
and U4911 (N_4911,N_976,N_151);
nor U4912 (N_4912,N_2038,N_446);
nor U4913 (N_4913,N_1624,N_529);
or U4914 (N_4914,N_143,N_2260);
xnor U4915 (N_4915,N_851,N_464);
nor U4916 (N_4916,N_2008,N_1541);
and U4917 (N_4917,N_555,N_795);
and U4918 (N_4918,N_1651,N_2168);
nand U4919 (N_4919,N_690,N_1040);
or U4920 (N_4920,N_1195,N_24);
xor U4921 (N_4921,N_2349,N_400);
xnor U4922 (N_4922,N_2409,N_2451);
nand U4923 (N_4923,N_1516,N_664);
xnor U4924 (N_4924,N_1575,N_424);
xor U4925 (N_4925,N_1590,N_2007);
nand U4926 (N_4926,N_1588,N_2199);
nor U4927 (N_4927,N_2249,N_1912);
or U4928 (N_4928,N_1968,N_1495);
or U4929 (N_4929,N_1478,N_360);
and U4930 (N_4930,N_1474,N_2188);
nor U4931 (N_4931,N_2024,N_2418);
nand U4932 (N_4932,N_1740,N_1474);
xor U4933 (N_4933,N_995,N_635);
or U4934 (N_4934,N_1095,N_1139);
xor U4935 (N_4935,N_1858,N_793);
and U4936 (N_4936,N_2423,N_1583);
or U4937 (N_4937,N_2373,N_536);
and U4938 (N_4938,N_1189,N_429);
nand U4939 (N_4939,N_1442,N_2271);
or U4940 (N_4940,N_1479,N_1854);
xor U4941 (N_4941,N_110,N_1396);
and U4942 (N_4942,N_464,N_2355);
nand U4943 (N_4943,N_2020,N_1653);
xnor U4944 (N_4944,N_1390,N_2035);
and U4945 (N_4945,N_1910,N_1056);
or U4946 (N_4946,N_590,N_1688);
xnor U4947 (N_4947,N_2473,N_150);
and U4948 (N_4948,N_1209,N_2061);
and U4949 (N_4949,N_842,N_1179);
nor U4950 (N_4950,N_1194,N_1440);
nor U4951 (N_4951,N_1064,N_1865);
xor U4952 (N_4952,N_2213,N_1154);
nand U4953 (N_4953,N_1017,N_1090);
and U4954 (N_4954,N_1568,N_2300);
xor U4955 (N_4955,N_706,N_533);
xnor U4956 (N_4956,N_210,N_1825);
xor U4957 (N_4957,N_2191,N_754);
and U4958 (N_4958,N_1675,N_1264);
nor U4959 (N_4959,N_140,N_689);
nand U4960 (N_4960,N_833,N_1802);
nor U4961 (N_4961,N_220,N_1589);
and U4962 (N_4962,N_2165,N_1650);
or U4963 (N_4963,N_2447,N_262);
or U4964 (N_4964,N_337,N_423);
xnor U4965 (N_4965,N_1030,N_503);
nand U4966 (N_4966,N_1287,N_1029);
and U4967 (N_4967,N_1118,N_1032);
nor U4968 (N_4968,N_131,N_1906);
nand U4969 (N_4969,N_1703,N_2453);
or U4970 (N_4970,N_2200,N_1999);
nor U4971 (N_4971,N_2346,N_1995);
and U4972 (N_4972,N_1429,N_1027);
nor U4973 (N_4973,N_1770,N_1483);
nand U4974 (N_4974,N_1332,N_1553);
or U4975 (N_4975,N_111,N_1883);
or U4976 (N_4976,N_2110,N_1659);
or U4977 (N_4977,N_2242,N_407);
nand U4978 (N_4978,N_173,N_2226);
and U4979 (N_4979,N_1925,N_1056);
nor U4980 (N_4980,N_954,N_1962);
xnor U4981 (N_4981,N_863,N_1874);
nor U4982 (N_4982,N_2116,N_2485);
xnor U4983 (N_4983,N_2333,N_429);
xnor U4984 (N_4984,N_433,N_769);
nand U4985 (N_4985,N_2424,N_767);
nand U4986 (N_4986,N_318,N_1663);
or U4987 (N_4987,N_1324,N_1296);
or U4988 (N_4988,N_1253,N_1260);
or U4989 (N_4989,N_290,N_975);
and U4990 (N_4990,N_1525,N_43);
nand U4991 (N_4991,N_211,N_2284);
nor U4992 (N_4992,N_1918,N_810);
nor U4993 (N_4993,N_2474,N_1642);
nand U4994 (N_4994,N_1899,N_949);
nor U4995 (N_4995,N_1539,N_671);
xor U4996 (N_4996,N_135,N_1774);
xnor U4997 (N_4997,N_2486,N_551);
or U4998 (N_4998,N_1585,N_746);
nor U4999 (N_4999,N_1933,N_2237);
nor U5000 (N_5000,N_3457,N_4375);
or U5001 (N_5001,N_4535,N_4866);
or U5002 (N_5002,N_3496,N_3207);
nand U5003 (N_5003,N_3978,N_3368);
and U5004 (N_5004,N_2992,N_4622);
or U5005 (N_5005,N_3498,N_3410);
nor U5006 (N_5006,N_3754,N_3329);
nor U5007 (N_5007,N_3305,N_4021);
xnor U5008 (N_5008,N_3282,N_3309);
or U5009 (N_5009,N_4997,N_3490);
nand U5010 (N_5010,N_3701,N_4121);
nand U5011 (N_5011,N_2519,N_2870);
nand U5012 (N_5012,N_3009,N_4367);
and U5013 (N_5013,N_4448,N_2949);
and U5014 (N_5014,N_4054,N_3893);
nand U5015 (N_5015,N_3447,N_3458);
nor U5016 (N_5016,N_4165,N_3685);
xnor U5017 (N_5017,N_3507,N_3155);
xnor U5018 (N_5018,N_4899,N_4842);
xnor U5019 (N_5019,N_4976,N_2551);
xor U5020 (N_5020,N_4679,N_4699);
or U5021 (N_5021,N_3828,N_2877);
or U5022 (N_5022,N_2871,N_4939);
and U5023 (N_5023,N_4212,N_4916);
nor U5024 (N_5024,N_4896,N_3246);
or U5025 (N_5025,N_2858,N_3208);
nand U5026 (N_5026,N_4494,N_2698);
nor U5027 (N_5027,N_4194,N_4401);
xor U5028 (N_5028,N_4973,N_4484);
xor U5029 (N_5029,N_3688,N_4928);
xnor U5030 (N_5030,N_4168,N_4096);
or U5031 (N_5031,N_4368,N_3802);
nor U5032 (N_5032,N_2863,N_4336);
or U5033 (N_5033,N_4644,N_4733);
or U5034 (N_5034,N_2711,N_4028);
nand U5035 (N_5035,N_2503,N_4618);
and U5036 (N_5036,N_3232,N_2534);
xor U5037 (N_5037,N_2866,N_2608);
xnor U5038 (N_5038,N_4822,N_2731);
or U5039 (N_5039,N_4462,N_3431);
and U5040 (N_5040,N_3593,N_4291);
nand U5041 (N_5041,N_4849,N_3074);
nor U5042 (N_5042,N_3965,N_3137);
and U5043 (N_5043,N_3994,N_3381);
nor U5044 (N_5044,N_4205,N_3929);
nand U5045 (N_5045,N_3642,N_2543);
nand U5046 (N_5046,N_4949,N_3669);
xor U5047 (N_5047,N_4171,N_2744);
nor U5048 (N_5048,N_3915,N_4583);
xnor U5049 (N_5049,N_3653,N_4472);
and U5050 (N_5050,N_2854,N_4693);
nand U5051 (N_5051,N_4027,N_2962);
nand U5052 (N_5052,N_3409,N_3334);
nand U5053 (N_5053,N_4546,N_3079);
or U5054 (N_5054,N_4247,N_4923);
or U5055 (N_5055,N_3575,N_3338);
nor U5056 (N_5056,N_4774,N_4049);
and U5057 (N_5057,N_4469,N_3779);
nor U5058 (N_5058,N_2690,N_4736);
nor U5059 (N_5059,N_3933,N_2624);
nand U5060 (N_5060,N_4875,N_3146);
xnor U5061 (N_5061,N_3563,N_4681);
xnor U5062 (N_5062,N_4598,N_2825);
nand U5063 (N_5063,N_3408,N_2823);
nor U5064 (N_5064,N_3818,N_4754);
and U5065 (N_5065,N_3921,N_2599);
xnor U5066 (N_5066,N_3151,N_2838);
and U5067 (N_5067,N_4688,N_4035);
xnor U5068 (N_5068,N_3036,N_3860);
xor U5069 (N_5069,N_3216,N_4773);
nor U5070 (N_5070,N_4238,N_3161);
and U5071 (N_5071,N_4600,N_4978);
and U5072 (N_5072,N_4189,N_2940);
xnor U5073 (N_5073,N_2953,N_4652);
or U5074 (N_5074,N_4541,N_3252);
nand U5075 (N_5075,N_3227,N_4363);
nand U5076 (N_5076,N_2650,N_3681);
and U5077 (N_5077,N_3240,N_3995);
xor U5078 (N_5078,N_4783,N_2548);
nand U5079 (N_5079,N_4180,N_4629);
or U5080 (N_5080,N_4468,N_2814);
xor U5081 (N_5081,N_4789,N_4422);
nor U5082 (N_5082,N_3570,N_3533);
or U5083 (N_5083,N_4214,N_3784);
or U5084 (N_5084,N_4474,N_2564);
xor U5085 (N_5085,N_4145,N_2558);
and U5086 (N_5086,N_4383,N_2905);
xnor U5087 (N_5087,N_3322,N_4139);
nand U5088 (N_5088,N_3082,N_4686);
nor U5089 (N_5089,N_2756,N_4534);
xnor U5090 (N_5090,N_3778,N_3595);
xnor U5091 (N_5091,N_3157,N_3165);
and U5092 (N_5092,N_2724,N_3990);
and U5093 (N_5093,N_3220,N_2970);
and U5094 (N_5094,N_4560,N_4898);
and U5095 (N_5095,N_4345,N_2899);
nor U5096 (N_5096,N_4843,N_3594);
and U5097 (N_5097,N_4625,N_2634);
or U5098 (N_5098,N_4073,N_3635);
nor U5099 (N_5099,N_3640,N_3848);
or U5100 (N_5100,N_4612,N_2582);
nor U5101 (N_5101,N_4955,N_4564);
xnor U5102 (N_5102,N_4846,N_3485);
and U5103 (N_5103,N_3486,N_3274);
and U5104 (N_5104,N_4132,N_3659);
or U5105 (N_5105,N_4926,N_3942);
nor U5106 (N_5106,N_2964,N_3327);
or U5107 (N_5107,N_3858,N_4816);
nor U5108 (N_5108,N_4911,N_4539);
or U5109 (N_5109,N_3621,N_3065);
nand U5110 (N_5110,N_4596,N_4196);
nand U5111 (N_5111,N_3158,N_4431);
nand U5112 (N_5112,N_3150,N_3697);
xnor U5113 (N_5113,N_4497,N_2879);
or U5114 (N_5114,N_3526,N_2986);
nor U5115 (N_5115,N_4714,N_3364);
and U5116 (N_5116,N_4316,N_3733);
nand U5117 (N_5117,N_3819,N_4201);
and U5118 (N_5118,N_4133,N_2555);
xnor U5119 (N_5119,N_2750,N_4830);
and U5120 (N_5120,N_3977,N_3646);
xnor U5121 (N_5121,N_3928,N_4356);
xor U5122 (N_5122,N_3992,N_3123);
nand U5123 (N_5123,N_3029,N_4909);
and U5124 (N_5124,N_4515,N_2827);
xnor U5125 (N_5125,N_4473,N_3047);
xnor U5126 (N_5126,N_4162,N_4533);
or U5127 (N_5127,N_3285,N_4210);
xnor U5128 (N_5128,N_2583,N_4251);
nand U5129 (N_5129,N_2754,N_4695);
and U5130 (N_5130,N_2795,N_4586);
or U5131 (N_5131,N_4292,N_4660);
xor U5132 (N_5132,N_2820,N_3537);
nand U5133 (N_5133,N_3665,N_4112);
nor U5134 (N_5134,N_4776,N_4461);
or U5135 (N_5135,N_2628,N_2762);
xor U5136 (N_5136,N_3742,N_3390);
nor U5137 (N_5137,N_4682,N_4325);
or U5138 (N_5138,N_3461,N_3766);
xor U5139 (N_5139,N_3710,N_4404);
nand U5140 (N_5140,N_2613,N_4507);
nor U5141 (N_5141,N_4421,N_4200);
or U5142 (N_5142,N_4000,N_4985);
and U5143 (N_5143,N_4913,N_4304);
nor U5144 (N_5144,N_4946,N_4319);
or U5145 (N_5145,N_3395,N_3234);
xnor U5146 (N_5146,N_3935,N_4272);
nand U5147 (N_5147,N_3986,N_4847);
or U5148 (N_5148,N_4364,N_3948);
nand U5149 (N_5149,N_4142,N_4762);
or U5150 (N_5150,N_2873,N_4701);
or U5151 (N_5151,N_3156,N_2654);
xor U5152 (N_5152,N_3926,N_4640);
or U5153 (N_5153,N_3293,N_3188);
or U5154 (N_5154,N_3820,N_4175);
nor U5155 (N_5155,N_4256,N_4127);
and U5156 (N_5156,N_3435,N_3266);
or U5157 (N_5157,N_4153,N_3326);
xnor U5158 (N_5158,N_2719,N_4123);
or U5159 (N_5159,N_3470,N_3023);
nand U5160 (N_5160,N_3854,N_4055);
xnor U5161 (N_5161,N_3297,N_4280);
xnor U5162 (N_5162,N_4837,N_4927);
nor U5163 (N_5163,N_4149,N_2995);
nand U5164 (N_5164,N_3342,N_2614);
nor U5165 (N_5165,N_2641,N_3280);
nor U5166 (N_5166,N_4502,N_3522);
xnor U5167 (N_5167,N_3940,N_4906);
or U5168 (N_5168,N_3463,N_3983);
xnor U5169 (N_5169,N_3981,N_3196);
or U5170 (N_5170,N_2955,N_4530);
nand U5171 (N_5171,N_4078,N_3476);
nand U5172 (N_5172,N_4820,N_2510);
xor U5173 (N_5173,N_2511,N_3279);
or U5174 (N_5174,N_2669,N_3159);
or U5175 (N_5175,N_4258,N_2813);
nor U5176 (N_5176,N_3959,N_4721);
and U5177 (N_5177,N_3693,N_4910);
xor U5178 (N_5178,N_4342,N_3260);
nand U5179 (N_5179,N_3465,N_2770);
nand U5180 (N_5180,N_3696,N_3233);
xnor U5181 (N_5181,N_2596,N_4388);
nand U5182 (N_5182,N_4097,N_3442);
nand U5183 (N_5183,N_4881,N_2906);
and U5184 (N_5184,N_3626,N_4282);
or U5185 (N_5185,N_3063,N_2980);
xor U5186 (N_5186,N_3172,N_3675);
or U5187 (N_5187,N_3468,N_3907);
nor U5188 (N_5188,N_4440,N_2531);
nand U5189 (N_5189,N_4182,N_4329);
and U5190 (N_5190,N_4536,N_3270);
and U5191 (N_5191,N_3980,N_2586);
nand U5192 (N_5192,N_2876,N_4449);
nand U5193 (N_5193,N_3816,N_3174);
nand U5194 (N_5194,N_4992,N_4274);
nor U5195 (N_5195,N_3712,N_4796);
nand U5196 (N_5196,N_4912,N_3292);
nand U5197 (N_5197,N_3734,N_3231);
or U5198 (N_5198,N_4435,N_3973);
xor U5199 (N_5199,N_2942,N_2612);
nor U5200 (N_5200,N_3198,N_3142);
nand U5201 (N_5201,N_2723,N_2682);
and U5202 (N_5202,N_4397,N_2990);
and U5203 (N_5203,N_4943,N_3949);
nor U5204 (N_5204,N_3616,N_3866);
or U5205 (N_5205,N_4755,N_4349);
and U5206 (N_5206,N_3918,N_2733);
or U5207 (N_5207,N_4861,N_4752);
and U5208 (N_5208,N_4917,N_2956);
or U5209 (N_5209,N_2793,N_3441);
xnor U5210 (N_5210,N_2755,N_2891);
nor U5211 (N_5211,N_2946,N_4979);
or U5212 (N_5212,N_2729,N_3643);
xnor U5213 (N_5213,N_3492,N_3005);
and U5214 (N_5214,N_4181,N_4931);
or U5215 (N_5215,N_3107,N_2853);
nand U5216 (N_5216,N_3695,N_3308);
or U5217 (N_5217,N_2715,N_2670);
and U5218 (N_5218,N_2716,N_3702);
nand U5219 (N_5219,N_4457,N_3917);
nor U5220 (N_5220,N_4977,N_3055);
xor U5221 (N_5221,N_3826,N_3609);
xnor U5222 (N_5222,N_2959,N_3124);
nand U5223 (N_5223,N_3467,N_3691);
nand U5224 (N_5224,N_4170,N_4608);
nor U5225 (N_5225,N_3275,N_3713);
and U5226 (N_5226,N_3972,N_2785);
or U5227 (N_5227,N_3169,N_3876);
nor U5228 (N_5228,N_4084,N_3104);
xor U5229 (N_5229,N_2842,N_3737);
or U5230 (N_5230,N_3755,N_4982);
or U5231 (N_5231,N_2622,N_3077);
nor U5232 (N_5232,N_2645,N_3251);
nand U5233 (N_5233,N_4657,N_4414);
nor U5234 (N_5234,N_2725,N_3262);
or U5235 (N_5235,N_4744,N_3128);
nand U5236 (N_5236,N_2666,N_4022);
and U5237 (N_5237,N_3328,N_3956);
nor U5238 (N_5238,N_3413,N_4989);
nand U5239 (N_5239,N_4108,N_2774);
nor U5240 (N_5240,N_4047,N_3690);
and U5241 (N_5241,N_3641,N_4290);
nor U5242 (N_5242,N_3186,N_3898);
nand U5243 (N_5243,N_2796,N_3471);
and U5244 (N_5244,N_2741,N_3098);
xor U5245 (N_5245,N_3599,N_3885);
and U5246 (N_5246,N_3925,N_3011);
nand U5247 (N_5247,N_2517,N_4335);
and U5248 (N_5248,N_4443,N_2701);
xor U5249 (N_5249,N_4211,N_4423);
xor U5250 (N_5250,N_4516,N_2562);
or U5251 (N_5251,N_2790,N_3117);
and U5252 (N_5252,N_3684,N_4808);
and U5253 (N_5253,N_4738,N_4174);
nor U5254 (N_5254,N_4878,N_3615);
xor U5255 (N_5255,N_3515,N_2544);
nor U5256 (N_5256,N_4405,N_4244);
nand U5257 (N_5257,N_4353,N_4557);
xor U5258 (N_5258,N_4555,N_4760);
and U5259 (N_5259,N_3394,N_4630);
xor U5260 (N_5260,N_4880,N_4716);
and U5261 (N_5261,N_2506,N_2742);
nor U5262 (N_5262,N_4591,N_4601);
nor U5263 (N_5263,N_3379,N_3518);
nor U5264 (N_5264,N_4587,N_2661);
nor U5265 (N_5265,N_2563,N_4452);
and U5266 (N_5266,N_4865,N_3529);
nand U5267 (N_5267,N_2800,N_3756);
nor U5268 (N_5268,N_4039,N_4260);
nand U5269 (N_5269,N_2933,N_4963);
nor U5270 (N_5270,N_3844,N_2789);
and U5271 (N_5271,N_3878,N_4143);
nor U5272 (N_5272,N_3096,N_3969);
xor U5273 (N_5273,N_4677,N_3738);
or U5274 (N_5274,N_3213,N_3139);
or U5275 (N_5275,N_4966,N_3066);
and U5276 (N_5276,N_3000,N_3206);
nor U5277 (N_5277,N_3782,N_3789);
nand U5278 (N_5278,N_4347,N_3562);
or U5279 (N_5279,N_2928,N_3423);
nand U5280 (N_5280,N_4848,N_3606);
nor U5281 (N_5281,N_4611,N_2592);
or U5282 (N_5282,N_3554,N_3068);
xnor U5283 (N_5283,N_4167,N_4713);
nand U5284 (N_5284,N_3323,N_2904);
nand U5285 (N_5285,N_4144,N_4542);
and U5286 (N_5286,N_4859,N_3312);
nand U5287 (N_5287,N_3436,N_4011);
and U5288 (N_5288,N_4751,N_3824);
nor U5289 (N_5289,N_3794,N_3548);
and U5290 (N_5290,N_3731,N_4960);
nor U5291 (N_5291,N_3783,N_3375);
xnor U5292 (N_5292,N_3369,N_2625);
nand U5293 (N_5293,N_3791,N_3460);
nand U5294 (N_5294,N_3145,N_2894);
xor U5295 (N_5295,N_4753,N_3194);
xnor U5296 (N_5296,N_3887,N_4044);
and U5297 (N_5297,N_4565,N_3572);
nor U5298 (N_5298,N_3135,N_4633);
or U5299 (N_5299,N_2809,N_3610);
nand U5300 (N_5300,N_3010,N_4801);
nand U5301 (N_5301,N_4777,N_3088);
or U5302 (N_5302,N_3052,N_4505);
and U5303 (N_5303,N_3429,N_2610);
or U5304 (N_5304,N_4434,N_3163);
or U5305 (N_5305,N_3474,N_4302);
nand U5306 (N_5306,N_3633,N_2950);
or U5307 (N_5307,N_4506,N_4825);
and U5308 (N_5308,N_4259,N_3420);
or U5309 (N_5309,N_4176,N_3686);
or U5310 (N_5310,N_3244,N_3725);
nor U5311 (N_5311,N_2501,N_4286);
and U5312 (N_5312,N_4178,N_3914);
xor U5313 (N_5313,N_4905,N_4020);
and U5314 (N_5314,N_4571,N_3936);
nor U5315 (N_5315,N_2938,N_3757);
or U5316 (N_5316,N_3941,N_2937);
xnor U5317 (N_5317,N_3298,N_3719);
and U5318 (N_5318,N_4191,N_3099);
nand U5319 (N_5319,N_4263,N_2673);
or U5320 (N_5320,N_3625,N_3013);
and U5321 (N_5321,N_3661,N_4081);
and U5322 (N_5322,N_3865,N_3551);
xor U5323 (N_5323,N_3834,N_3149);
and U5324 (N_5324,N_2726,N_4856);
nand U5325 (N_5325,N_3489,N_4902);
nor U5326 (N_5326,N_2978,N_4990);
and U5327 (N_5327,N_4420,N_4278);
nand U5328 (N_5328,N_4467,N_4897);
or U5329 (N_5329,N_4340,N_3604);
nand U5330 (N_5330,N_3114,N_3565);
or U5331 (N_5331,N_3552,N_4791);
nor U5332 (N_5332,N_4236,N_4412);
nand U5333 (N_5333,N_3475,N_4545);
nor U5334 (N_5334,N_4662,N_4346);
nor U5335 (N_5335,N_3836,N_4962);
or U5336 (N_5336,N_4293,N_4582);
and U5337 (N_5337,N_4159,N_4231);
and U5338 (N_5338,N_4602,N_4550);
nor U5339 (N_5339,N_4839,N_4815);
nor U5340 (N_5340,N_4115,N_2536);
and U5341 (N_5341,N_3030,N_3437);
or U5342 (N_5342,N_4155,N_4454);
xnor U5343 (N_5343,N_4128,N_4694);
nand U5344 (N_5344,N_4313,N_3739);
nand U5345 (N_5345,N_4066,N_4046);
xnor U5346 (N_5346,N_3652,N_4122);
xnor U5347 (N_5347,N_3888,N_4137);
xor U5348 (N_5348,N_3049,N_2588);
xnor U5349 (N_5349,N_4409,N_2893);
and U5350 (N_5350,N_4350,N_2507);
and U5351 (N_5351,N_3201,N_3937);
nand U5352 (N_5352,N_4790,N_4935);
nor U5353 (N_5353,N_3358,N_3225);
and U5354 (N_5354,N_3272,N_2761);
and U5355 (N_5355,N_4988,N_3830);
and U5356 (N_5356,N_2930,N_3401);
xnor U5357 (N_5357,N_2554,N_2901);
xor U5358 (N_5358,N_4664,N_3190);
or U5359 (N_5359,N_3164,N_2925);
and U5360 (N_5360,N_4481,N_3530);
nand U5361 (N_5361,N_3982,N_3454);
nand U5362 (N_5362,N_4882,N_4965);
or U5363 (N_5363,N_4958,N_3979);
nand U5364 (N_5364,N_4800,N_3373);
xor U5365 (N_5365,N_3303,N_2663);
or U5366 (N_5366,N_3953,N_3176);
or U5367 (N_5367,N_4719,N_4396);
nand U5368 (N_5368,N_4206,N_4951);
or U5369 (N_5369,N_3415,N_4863);
xnor U5370 (N_5370,N_3863,N_4737);
and U5371 (N_5371,N_3171,N_4584);
nor U5372 (N_5372,N_4821,N_2892);
nand U5373 (N_5373,N_3185,N_4741);
nand U5374 (N_5374,N_3359,N_4438);
or U5375 (N_5375,N_4001,N_3152);
or U5376 (N_5376,N_3060,N_3456);
nor U5377 (N_5377,N_2607,N_3264);
nor U5378 (N_5378,N_4482,N_3452);
and U5379 (N_5379,N_4855,N_4219);
and U5380 (N_5380,N_4378,N_4567);
and U5381 (N_5381,N_3545,N_3775);
nor U5382 (N_5382,N_3497,N_4471);
nand U5383 (N_5383,N_3908,N_4854);
xnor U5384 (N_5384,N_4059,N_2571);
or U5385 (N_5385,N_4092,N_3307);
nor U5386 (N_5386,N_4797,N_3763);
xor U5387 (N_5387,N_4580,N_4980);
or U5388 (N_5388,N_3187,N_4068);
or U5389 (N_5389,N_3668,N_4060);
nand U5390 (N_5390,N_2584,N_4413);
xnor U5391 (N_5391,N_3944,N_4261);
xor U5392 (N_5392,N_4314,N_2749);
xnor U5393 (N_5393,N_4298,N_4945);
and U5394 (N_5394,N_3101,N_2890);
nor U5395 (N_5395,N_2515,N_3842);
xnor U5396 (N_5396,N_4944,N_3683);
and U5397 (N_5397,N_4594,N_3481);
and U5398 (N_5398,N_4130,N_3058);
xor U5399 (N_5399,N_3038,N_2627);
nor U5400 (N_5400,N_2695,N_3771);
nand U5401 (N_5401,N_3070,N_3923);
nand U5402 (N_5402,N_4496,N_2851);
nand U5403 (N_5403,N_4747,N_3897);
and U5404 (N_5404,N_3179,N_3277);
and U5405 (N_5405,N_3875,N_2822);
nor U5406 (N_5406,N_4495,N_4391);
nor U5407 (N_5407,N_3955,N_4860);
and U5408 (N_5408,N_3504,N_4470);
nand U5409 (N_5409,N_3817,N_4332);
and U5410 (N_5410,N_3541,N_3366);
and U5411 (N_5411,N_2739,N_4673);
nor U5412 (N_5412,N_3720,N_4013);
or U5413 (N_5413,N_4003,N_3374);
or U5414 (N_5414,N_4903,N_3085);
or U5415 (N_5415,N_4779,N_3823);
or U5416 (N_5416,N_3516,N_4488);
nand U5417 (N_5417,N_2685,N_3717);
nand U5418 (N_5418,N_2769,N_3472);
nand U5419 (N_5419,N_3112,N_3735);
and U5420 (N_5420,N_2537,N_4592);
nor U5421 (N_5421,N_4643,N_4498);
or U5422 (N_5422,N_3574,N_3178);
or U5423 (N_5423,N_3662,N_2948);
or U5424 (N_5424,N_3017,N_3879);
or U5425 (N_5425,N_2764,N_4240);
or U5426 (N_5426,N_3881,N_4551);
or U5427 (N_5427,N_4163,N_4070);
or U5428 (N_5428,N_3718,N_2617);
nand U5429 (N_5429,N_3257,N_4793);
xnor U5430 (N_5430,N_3118,N_4840);
or U5431 (N_5431,N_4327,N_2700);
nor U5432 (N_5432,N_3512,N_4953);
nand U5433 (N_5433,N_4374,N_4532);
or U5434 (N_5434,N_4617,N_3283);
nor U5435 (N_5435,N_3748,N_2806);
xor U5436 (N_5436,N_2887,N_4769);
or U5437 (N_5437,N_3352,N_3709);
xor U5438 (N_5438,N_2856,N_4025);
xnor U5439 (N_5439,N_4704,N_4510);
xor U5440 (N_5440,N_2604,N_4748);
nor U5441 (N_5441,N_3350,N_4154);
and U5442 (N_5442,N_3378,N_4079);
xnor U5443 (N_5443,N_4879,N_3193);
and U5444 (N_5444,N_3245,N_3601);
xnor U5445 (N_5445,N_2572,N_3539);
nor U5446 (N_5446,N_4606,N_3051);
nor U5447 (N_5447,N_2874,N_2801);
and U5448 (N_5448,N_3509,N_4938);
or U5449 (N_5449,N_2797,N_4919);
nor U5450 (N_5450,N_4463,N_4465);
nand U5451 (N_5451,N_2678,N_3964);
nand U5452 (N_5452,N_3989,N_2912);
nor U5453 (N_5453,N_4718,N_2969);
nor U5454 (N_5454,N_4080,N_4004);
nor U5455 (N_5455,N_4008,N_2589);
nand U5456 (N_5456,N_4692,N_2975);
xor U5457 (N_5457,N_3673,N_2915);
nand U5458 (N_5458,N_4101,N_4503);
or U5459 (N_5459,N_3692,N_3938);
and U5460 (N_5460,N_2603,N_3287);
xnor U5461 (N_5461,N_2713,N_3611);
nand U5462 (N_5462,N_4573,N_2821);
and U5463 (N_5463,N_4563,N_3294);
or U5464 (N_5464,N_4745,N_2691);
or U5465 (N_5465,N_3667,N_3167);
xnor U5466 (N_5466,N_3024,N_4424);
xor U5467 (N_5467,N_4500,N_3622);
and U5468 (N_5468,N_3744,N_3841);
or U5469 (N_5469,N_4276,N_3416);
nor U5470 (N_5470,N_4117,N_3090);
nand U5471 (N_5471,N_4684,N_2699);
nand U5472 (N_5472,N_3064,N_3527);
nand U5473 (N_5473,N_2524,N_3803);
nand U5474 (N_5474,N_2803,N_3950);
and U5475 (N_5475,N_4243,N_3008);
xnor U5476 (N_5476,N_3805,N_4088);
xnor U5477 (N_5477,N_3125,N_2606);
nand U5478 (N_5478,N_4894,N_2845);
xor U5479 (N_5479,N_3785,N_4283);
nor U5480 (N_5480,N_3920,N_4838);
or U5481 (N_5481,N_4017,N_3110);
xor U5482 (N_5482,N_4845,N_3822);
nor U5483 (N_5483,N_4869,N_2815);
nor U5484 (N_5484,N_3962,N_3567);
xor U5485 (N_5485,N_3493,N_3448);
nand U5486 (N_5486,N_4520,N_4828);
nand U5487 (N_5487,N_3511,N_4224);
or U5488 (N_5488,N_4941,N_3016);
nor U5489 (N_5489,N_4217,N_3067);
and U5490 (N_5490,N_2730,N_4607);
nand U5491 (N_5491,N_3462,N_4930);
nand U5492 (N_5492,N_4914,N_2734);
and U5493 (N_5493,N_4058,N_4746);
xnor U5494 (N_5494,N_4802,N_3411);
xnor U5495 (N_5495,N_4169,N_4250);
nor U5496 (N_5496,N_4442,N_4957);
xor U5497 (N_5497,N_3434,N_4307);
xor U5498 (N_5498,N_4296,N_3414);
nand U5499 (N_5499,N_4784,N_4086);
xnor U5500 (N_5500,N_3650,N_2587);
and U5501 (N_5501,N_2881,N_3957);
or U5502 (N_5502,N_4844,N_4810);
or U5503 (N_5503,N_3175,N_3761);
or U5504 (N_5504,N_4277,N_2565);
xnor U5505 (N_5505,N_3954,N_4402);
nor U5506 (N_5506,N_3976,N_3549);
xnor U5507 (N_5507,N_2985,N_2917);
nand U5508 (N_5508,N_3094,N_3741);
xor U5509 (N_5509,N_3081,N_2798);
xnor U5510 (N_5510,N_3310,N_2527);
or U5511 (N_5511,N_4991,N_2861);
or U5512 (N_5512,N_4411,N_4289);
xor U5513 (N_5513,N_4799,N_4116);
xnor U5514 (N_5514,N_4104,N_2740);
or U5515 (N_5515,N_4483,N_3634);
and U5516 (N_5516,N_3397,N_3422);
or U5517 (N_5517,N_3578,N_3376);
nor U5518 (N_5518,N_4439,N_2696);
and U5519 (N_5519,N_4295,N_3687);
and U5520 (N_5520,N_3573,N_4156);
or U5521 (N_5521,N_4841,N_4357);
xnor U5522 (N_5522,N_4014,N_3093);
nand U5523 (N_5523,N_3506,N_2520);
nand U5524 (N_5524,N_4249,N_2834);
nor U5525 (N_5525,N_3586,N_3655);
nand U5526 (N_5526,N_4576,N_4823);
xnor U5527 (N_5527,N_2500,N_2530);
nand U5528 (N_5528,N_3459,N_3613);
nor U5529 (N_5529,N_3086,N_4665);
nor U5530 (N_5530,N_3271,N_3916);
and U5531 (N_5531,N_2570,N_3212);
or U5532 (N_5532,N_4729,N_2528);
nand U5533 (N_5533,N_3555,N_4197);
and U5534 (N_5534,N_2602,N_3400);
and U5535 (N_5535,N_3349,N_3396);
xor U5536 (N_5536,N_3619,N_4009);
xnor U5537 (N_5537,N_4893,N_2872);
xnor U5538 (N_5538,N_4778,N_3727);
nand U5539 (N_5539,N_3729,N_4148);
xor U5540 (N_5540,N_3988,N_4297);
nor U5541 (N_5541,N_4676,N_4659);
or U5542 (N_5542,N_4445,N_2652);
xnor U5543 (N_5543,N_2843,N_4226);
nor U5544 (N_5544,N_2704,N_3795);
or U5545 (N_5545,N_2545,N_2960);
or U5546 (N_5546,N_3591,N_3343);
and U5547 (N_5547,N_3335,N_3367);
nand U5548 (N_5548,N_2738,N_2810);
and U5549 (N_5549,N_3707,N_3597);
or U5550 (N_5550,N_3815,N_3018);
xor U5551 (N_5551,N_3069,N_2643);
and U5552 (N_5552,N_4177,N_4354);
xor U5553 (N_5553,N_3451,N_3630);
nor U5554 (N_5554,N_4106,N_4102);
and U5555 (N_5555,N_4675,N_2846);
nand U5556 (N_5556,N_3050,N_2763);
or U5557 (N_5557,N_4871,N_3056);
xor U5558 (N_5558,N_4392,N_4524);
xor U5559 (N_5559,N_3774,N_3600);
and U5560 (N_5560,N_3062,N_3810);
xnor U5561 (N_5561,N_3523,N_3821);
or U5562 (N_5562,N_3540,N_3446);
nor U5563 (N_5563,N_3189,N_3106);
nor U5564 (N_5564,N_4339,N_4750);
nor U5565 (N_5565,N_4759,N_4786);
nor U5566 (N_5566,N_2816,N_2683);
and U5567 (N_5567,N_3542,N_4782);
and U5568 (N_5568,N_4886,N_4616);
or U5569 (N_5569,N_4868,N_2841);
or U5570 (N_5570,N_4715,N_2971);
or U5571 (N_5571,N_2888,N_3300);
nand U5572 (N_5572,N_4103,N_3825);
nor U5573 (N_5573,N_4408,N_4418);
nand U5574 (N_5574,N_3347,N_3910);
and U5575 (N_5575,N_3153,N_3804);
xnor U5576 (N_5576,N_4273,N_2623);
nor U5577 (N_5577,N_2760,N_2923);
or U5578 (N_5578,N_3180,N_4956);
nor U5579 (N_5579,N_4002,N_3874);
or U5580 (N_5580,N_4034,N_4831);
or U5581 (N_5581,N_3318,N_4430);
and U5582 (N_5582,N_3556,N_4650);
nand U5583 (N_5583,N_4399,N_3404);
and U5584 (N_5584,N_3872,N_2573);
nand U5585 (N_5585,N_4253,N_4062);
nand U5586 (N_5586,N_3239,N_3215);
and U5587 (N_5587,N_4372,N_2883);
or U5588 (N_5588,N_3331,N_4974);
or U5589 (N_5589,N_4727,N_4284);
nor U5590 (N_5590,N_4382,N_3632);
nor U5591 (N_5591,N_3663,N_2694);
and U5592 (N_5592,N_3028,N_2772);
nand U5593 (N_5593,N_3867,N_4235);
xor U5594 (N_5594,N_3838,N_3746);
nor U5595 (N_5595,N_2830,N_2556);
nor U5596 (N_5596,N_4222,N_4940);
xor U5597 (N_5597,N_4232,N_4813);
or U5598 (N_5598,N_3528,N_2646);
or U5599 (N_5599,N_4126,N_4365);
xor U5600 (N_5600,N_4362,N_3182);
nand U5601 (N_5601,N_2984,N_3571);
and U5602 (N_5602,N_4671,N_3631);
nand U5603 (N_5603,N_4647,N_4666);
nor U5604 (N_5604,N_4519,N_2736);
nand U5605 (N_5605,N_4242,N_4087);
nand U5606 (N_5606,N_3249,N_2514);
and U5607 (N_5607,N_3048,N_3205);
or U5608 (N_5608,N_4766,N_3544);
nor U5609 (N_5609,N_4892,N_4269);
or U5610 (N_5610,N_2708,N_3608);
nand U5611 (N_5611,N_2751,N_2848);
nor U5612 (N_5612,N_3267,N_2999);
xor U5613 (N_5613,N_2943,N_3391);
nand U5614 (N_5614,N_3596,N_3807);
xor U5615 (N_5615,N_4901,N_3419);
xnor U5616 (N_5616,N_2997,N_3314);
or U5617 (N_5617,N_3403,N_3660);
xnor U5618 (N_5618,N_2941,N_2550);
and U5619 (N_5619,N_2522,N_3348);
nor U5620 (N_5620,N_4763,N_2581);
nand U5621 (N_5621,N_3053,N_3627);
or U5622 (N_5622,N_4575,N_3083);
or U5623 (N_5623,N_4239,N_4877);
xnor U5624 (N_5624,N_2835,N_2637);
xnor U5625 (N_5625,N_4486,N_4604);
nand U5626 (N_5626,N_2907,N_4136);
or U5627 (N_5627,N_2567,N_3387);
nor U5628 (N_5628,N_4628,N_2811);
nand U5629 (N_5629,N_4798,N_3852);
xnor U5630 (N_5630,N_3412,N_3333);
nand U5631 (N_5631,N_3568,N_3793);
nand U5632 (N_5632,N_3525,N_3590);
nand U5633 (N_5633,N_4700,N_2847);
nand U5634 (N_5634,N_2653,N_3877);
xnor U5635 (N_5635,N_3671,N_3857);
and U5636 (N_5636,N_4639,N_4056);
xor U5637 (N_5637,N_2918,N_4433);
and U5638 (N_5638,N_3813,N_4348);
or U5639 (N_5639,N_4947,N_2927);
or U5640 (N_5640,N_4147,N_3091);
and U5641 (N_5641,N_3261,N_2868);
nor U5642 (N_5642,N_2512,N_4215);
xor U5643 (N_5643,N_4164,N_3945);
xor U5644 (N_5644,N_4544,N_4385);
and U5645 (N_5645,N_4152,N_4994);
or U5646 (N_5646,N_2513,N_4562);
or U5647 (N_5647,N_4403,N_4306);
nor U5648 (N_5648,N_3587,N_4605);
or U5649 (N_5649,N_4883,N_2590);
or U5650 (N_5650,N_3799,N_3780);
nand U5651 (N_5651,N_3508,N_2712);
nand U5652 (N_5652,N_2780,N_2860);
and U5653 (N_5653,N_2597,N_4466);
nor U5654 (N_5654,N_4585,N_4780);
or U5655 (N_5655,N_3203,N_2737);
nand U5656 (N_5656,N_2629,N_4221);
nor U5657 (N_5657,N_4105,N_2791);
and U5658 (N_5658,N_3007,N_4959);
nand U5659 (N_5659,N_4379,N_3535);
or U5660 (N_5660,N_3195,N_3421);
nand U5661 (N_5661,N_3398,N_2542);
xor U5662 (N_5662,N_3097,N_2585);
nor U5663 (N_5663,N_3426,N_3177);
nand U5664 (N_5664,N_3122,N_2605);
or U5665 (N_5665,N_3214,N_2799);
and U5666 (N_5666,N_3624,N_4588);
or U5667 (N_5667,N_2919,N_3044);
or U5668 (N_5668,N_2649,N_4265);
nand U5669 (N_5669,N_4380,N_3495);
nor U5670 (N_5670,N_3576,N_4743);
xnor U5671 (N_5671,N_3095,N_4687);
nor U5672 (N_5672,N_4225,N_3943);
or U5673 (N_5673,N_2676,N_2687);
nand U5674 (N_5674,N_4521,N_3361);
nand U5675 (N_5675,N_2508,N_4888);
or U5676 (N_5676,N_4918,N_4477);
and U5677 (N_5677,N_3357,N_3952);
and U5678 (N_5678,N_3311,N_2884);
or U5679 (N_5679,N_3281,N_3612);
nor U5680 (N_5680,N_4040,N_4389);
nor U5681 (N_5681,N_4566,N_3843);
and U5682 (N_5682,N_4255,N_3002);
nand U5683 (N_5683,N_2837,N_4832);
and U5684 (N_5684,N_4884,N_4853);
nor U5685 (N_5685,N_3217,N_4161);
nand U5686 (N_5686,N_4303,N_2595);
nand U5687 (N_5687,N_3682,N_3080);
xor U5688 (N_5688,N_4241,N_2703);
nand U5689 (N_5689,N_2748,N_4333);
nand U5690 (N_5690,N_4873,N_3930);
nand U5691 (N_5691,N_2559,N_3483);
nand U5692 (N_5692,N_4835,N_2983);
nand U5693 (N_5693,N_2771,N_4954);
nor U5694 (N_5694,N_4330,N_4908);
and U5695 (N_5695,N_3730,N_3740);
and U5696 (N_5696,N_2908,N_3870);
or U5697 (N_5697,N_3134,N_3100);
xnor U5698 (N_5698,N_4485,N_4281);
or U5699 (N_5699,N_4436,N_3985);
xor U5700 (N_5700,N_2611,N_3019);
and U5701 (N_5701,N_2601,N_4809);
xor U5702 (N_5702,N_4981,N_4045);
xor U5703 (N_5703,N_2709,N_4570);
nand U5704 (N_5704,N_2996,N_4775);
nand U5705 (N_5705,N_2776,N_2720);
or U5706 (N_5706,N_3753,N_2552);
or U5707 (N_5707,N_4971,N_4792);
nor U5708 (N_5708,N_4384,N_4455);
xnor U5709 (N_5709,N_3399,N_3168);
nor U5710 (N_5710,N_4220,N_2523);
or U5711 (N_5711,N_3229,N_3623);
or U5712 (N_5712,N_3773,N_4287);
xnor U5713 (N_5713,N_4740,N_4033);
xnor U5714 (N_5714,N_2898,N_3290);
and U5715 (N_5715,N_3677,N_2509);
nor U5716 (N_5716,N_3278,N_2805);
nor U5717 (N_5717,N_2541,N_3202);
or U5718 (N_5718,N_3603,N_3859);
and U5719 (N_5719,N_3315,N_4537);
or U5720 (N_5720,N_2878,N_2674);
or U5721 (N_5721,N_4098,N_4538);
xnor U5722 (N_5722,N_3389,N_4862);
and U5723 (N_5723,N_3120,N_4310);
nand U5724 (N_5724,N_4305,N_3380);
and U5725 (N_5725,N_4326,N_2794);
nand U5726 (N_5726,N_4031,N_2664);
nand U5727 (N_5727,N_3041,N_3583);
nor U5728 (N_5728,N_3302,N_4728);
or U5729 (N_5729,N_4109,N_4514);
and U5730 (N_5730,N_3012,N_2561);
nor U5731 (N_5731,N_4726,N_3140);
or U5732 (N_5732,N_4048,N_3678);
nand U5733 (N_5733,N_2538,N_3078);
or U5734 (N_5734,N_4450,N_4301);
or U5735 (N_5735,N_3054,N_4999);
or U5736 (N_5736,N_4275,N_4857);
and U5737 (N_5737,N_4361,N_4267);
nor U5738 (N_5738,N_2991,N_3382);
nor U5739 (N_5739,N_3644,N_4120);
or U5740 (N_5740,N_3071,N_4512);
nor U5741 (N_5741,N_3919,N_3230);
nand U5742 (N_5742,N_2880,N_3765);
nand U5743 (N_5743,N_2945,N_2518);
nand U5744 (N_5744,N_4437,N_4885);
or U5745 (N_5745,N_4019,N_2504);
and U5746 (N_5746,N_3582,N_3851);
nor U5747 (N_5747,N_2546,N_3473);
nand U5748 (N_5748,N_4805,N_4271);
nand U5749 (N_5749,N_4936,N_4257);
or U5750 (N_5750,N_4065,N_3255);
and U5751 (N_5751,N_4720,N_2705);
or U5752 (N_5752,N_2658,N_3968);
nand U5753 (N_5753,N_4441,N_4285);
nor U5754 (N_5754,N_4623,N_4007);
and U5755 (N_5755,N_2746,N_3762);
nand U5756 (N_5756,N_3108,N_4279);
nor U5757 (N_5757,N_4826,N_4501);
or U5758 (N_5758,N_3922,N_4620);
nand U5759 (N_5759,N_2849,N_4311);
nand U5760 (N_5760,N_4195,N_4366);
or U5761 (N_5761,N_3491,N_2886);
or U5762 (N_5762,N_3443,N_3751);
nor U5763 (N_5763,N_4589,N_3557);
nor U5764 (N_5764,N_3076,N_2633);
xor U5765 (N_5765,N_4561,N_3371);
and U5766 (N_5766,N_3598,N_3647);
or U5767 (N_5767,N_3464,N_3383);
or U5768 (N_5768,N_4322,N_2900);
xnor U5769 (N_5769,N_3405,N_2783);
nand U5770 (N_5770,N_2897,N_4937);
nand U5771 (N_5771,N_4669,N_3478);
xnor U5772 (N_5772,N_4053,N_3034);
nor U5773 (N_5773,N_4493,N_4107);
nand U5774 (N_5774,N_3487,N_3336);
nand U5775 (N_5775,N_2957,N_3645);
nand U5776 (N_5776,N_4315,N_2920);
nand U5777 (N_5777,N_3021,N_4141);
xor U5778 (N_5778,N_3449,N_3250);
nand U5779 (N_5779,N_2639,N_2875);
xor U5780 (N_5780,N_4621,N_4491);
xor U5781 (N_5781,N_4270,N_2707);
and U5782 (N_5782,N_3704,N_3500);
or U5783 (N_5783,N_3042,N_3265);
xnor U5784 (N_5784,N_4426,N_4234);
nand U5785 (N_5785,N_2882,N_4969);
nor U5786 (N_5786,N_3708,N_2965);
or U5787 (N_5787,N_3466,N_2655);
nand U5788 (N_5788,N_3705,N_4248);
xor U5789 (N_5789,N_3564,N_3247);
nor U5790 (N_5790,N_4987,N_4158);
xnor U5791 (N_5791,N_4245,N_3868);
nand U5792 (N_5792,N_4138,N_4627);
xnor U5793 (N_5793,N_4785,N_2560);
xor U5794 (N_5794,N_4406,N_3679);
and U5795 (N_5795,N_3126,N_2672);
or U5796 (N_5796,N_3003,N_3767);
nand U5797 (N_5797,N_3801,N_4795);
nand U5798 (N_5798,N_4230,N_2636);
nand U5799 (N_5799,N_4328,N_2626);
xnor U5800 (N_5800,N_4344,N_4183);
or U5801 (N_5801,N_4061,N_4052);
or U5802 (N_5802,N_2914,N_3832);
or U5803 (N_5803,N_3951,N_3228);
or U5804 (N_5804,N_3806,N_4824);
and U5805 (N_5805,N_2895,N_3853);
or U5806 (N_5806,N_2916,N_4113);
and U5807 (N_5807,N_2569,N_4803);
xor U5808 (N_5808,N_4649,N_3132);
xnor U5809 (N_5809,N_4114,N_3934);
nand U5810 (N_5810,N_4597,N_3649);
nand U5811 (N_5811,N_2743,N_2525);
nand U5812 (N_5812,N_4995,N_2757);
or U5813 (N_5813,N_3809,N_4707);
nand U5814 (N_5814,N_3750,N_4950);
nor U5815 (N_5815,N_2934,N_3984);
nor U5816 (N_5816,N_3325,N_4895);
xnor U5817 (N_5817,N_4864,N_4513);
and U5818 (N_5818,N_3316,N_4499);
nand U5819 (N_5819,N_2766,N_3129);
nor U5820 (N_5820,N_4645,N_2577);
nand U5821 (N_5821,N_2721,N_2580);
and U5822 (N_5822,N_2665,N_3337);
and U5823 (N_5823,N_3520,N_3694);
and U5824 (N_5824,N_3269,N_4717);
or U5825 (N_5825,N_4479,N_3306);
nor U5826 (N_5826,N_4920,N_2832);
and U5827 (N_5827,N_4609,N_3602);
nand U5828 (N_5828,N_2994,N_2977);
and U5829 (N_5829,N_3840,N_4578);
and U5830 (N_5830,N_3637,N_3344);
and U5831 (N_5831,N_4858,N_4579);
nor U5832 (N_5832,N_4460,N_2574);
and U5833 (N_5833,N_4288,N_3883);
nor U5834 (N_5834,N_3676,N_3911);
nand U5835 (N_5835,N_4228,N_2885);
xor U5836 (N_5836,N_4308,N_3903);
or U5837 (N_5837,N_3392,N_3480);
xor U5838 (N_5838,N_3061,N_4262);
or U5839 (N_5839,N_2779,N_3769);
nor U5840 (N_5840,N_3706,N_2889);
nand U5841 (N_5841,N_3654,N_2855);
xor U5842 (N_5842,N_3510,N_4377);
and U5843 (N_5843,N_2535,N_4553);
xnor U5844 (N_5844,N_4904,N_4151);
xnor U5845 (N_5845,N_3424,N_3797);
nor U5846 (N_5846,N_3927,N_3835);
or U5847 (N_5847,N_4626,N_3931);
nor U5848 (N_5848,N_3736,N_4077);
and U5849 (N_5849,N_3726,N_3006);
nor U5850 (N_5850,N_4634,N_4967);
nand U5851 (N_5851,N_4207,N_4509);
or U5852 (N_5852,N_3295,N_4184);
nor U5853 (N_5853,N_4756,N_4648);
or U5854 (N_5854,N_3538,N_2981);
nand U5855 (N_5855,N_3289,N_4690);
or U5856 (N_5856,N_3996,N_2759);
and U5857 (N_5857,N_3469,N_2647);
and U5858 (N_5858,N_4321,N_3722);
or U5859 (N_5859,N_2516,N_3363);
or U5860 (N_5860,N_3909,N_4651);
nor U5861 (N_5861,N_2638,N_3882);
nand U5862 (N_5862,N_2502,N_3211);
xor U5863 (N_5863,N_2656,N_3524);
or U5864 (N_5864,N_3505,N_4697);
and U5865 (N_5865,N_4531,N_3324);
xor U5866 (N_5866,N_2993,N_4160);
nand U5867 (N_5867,N_4089,N_3004);
nor U5868 (N_5868,N_3913,N_4026);
or U5869 (N_5869,N_3276,N_4487);
nand U5870 (N_5870,N_3732,N_4093);
nor U5871 (N_5871,N_4661,N_2781);
and U5872 (N_5872,N_3248,N_3788);
nor U5873 (N_5873,N_3698,N_4173);
nor U5874 (N_5874,N_4199,N_2747);
or U5875 (N_5875,N_3284,N_3902);
nor U5876 (N_5876,N_2910,N_4731);
nor U5877 (N_5877,N_3192,N_4934);
and U5878 (N_5878,N_4432,N_3362);
or U5879 (N_5879,N_3402,N_4540);
nand U5880 (N_5880,N_3072,N_3113);
and U5881 (N_5881,N_4552,N_3022);
or U5882 (N_5882,N_3618,N_2692);
nor U5883 (N_5883,N_3222,N_3869);
xor U5884 (N_5884,N_3658,N_2828);
nand U5885 (N_5885,N_3884,N_2896);
and U5886 (N_5886,N_3263,N_4549);
xor U5887 (N_5887,N_4814,N_3224);
or U5888 (N_5888,N_3714,N_3974);
and U5889 (N_5889,N_3758,N_3427);
and U5890 (N_5890,N_4998,N_3235);
xnor U5891 (N_5891,N_3313,N_3519);
xor U5892 (N_5892,N_4386,N_2566);
nand U5893 (N_5893,N_4668,N_3116);
nand U5894 (N_5894,N_4095,N_4124);
nor U5895 (N_5895,N_4119,N_3880);
or U5896 (N_5896,N_4459,N_4525);
nand U5897 (N_5897,N_3059,N_4480);
xnor U5898 (N_5898,N_2775,N_3559);
xnor U5899 (N_5899,N_3291,N_3546);
and U5900 (N_5900,N_2786,N_2850);
xor U5901 (N_5901,N_4360,N_3341);
or U5902 (N_5902,N_2911,N_3716);
nor U5903 (N_5903,N_4577,N_3027);
and U5904 (N_5904,N_4915,N_4674);
nand U5905 (N_5905,N_2630,N_4593);
or U5906 (N_5906,N_2998,N_4932);
or U5907 (N_5907,N_4203,N_2961);
nor U5908 (N_5908,N_4975,N_3620);
or U5909 (N_5909,N_4654,N_4429);
xnor U5910 (N_5910,N_3455,N_2732);
nand U5911 (N_5911,N_3040,N_3184);
and U5912 (N_5912,N_3450,N_2728);
or U5913 (N_5913,N_4925,N_4029);
and U5914 (N_5914,N_4118,N_3745);
xnor U5915 (N_5915,N_4458,N_4416);
and U5916 (N_5916,N_4369,N_3484);
and U5917 (N_5917,N_4511,N_2579);
nor U5918 (N_5918,N_4051,N_2718);
xnor U5919 (N_5919,N_3340,N_4190);
nor U5920 (N_5920,N_4338,N_4807);
nand U5921 (N_5921,N_4683,N_3259);
xor U5922 (N_5922,N_2807,N_4787);
and U5923 (N_5923,N_3115,N_2951);
nor U5924 (N_5924,N_4610,N_4192);
or U5925 (N_5925,N_4638,N_3242);
xnor U5926 (N_5926,N_3724,N_3998);
xnor U5927 (N_5927,N_4834,N_2792);
nand U5928 (N_5928,N_4768,N_4179);
or U5929 (N_5929,N_3856,N_4724);
or U5930 (N_5930,N_2802,N_4264);
nor U5931 (N_5931,N_4523,N_2974);
or U5932 (N_5932,N_3657,N_4015);
or U5933 (N_5933,N_3723,N_3670);
nor U5934 (N_5934,N_4900,N_2782);
or U5935 (N_5935,N_4016,N_4772);
nor U5936 (N_5936,N_2667,N_3092);
nor U5937 (N_5937,N_3617,N_2921);
nor U5938 (N_5938,N_3811,N_4185);
nor U5939 (N_5939,N_2932,N_4739);
and U5940 (N_5940,N_2867,N_4111);
nor U5941 (N_5941,N_2529,N_2680);
nor U5942 (N_5942,N_3440,N_3651);
and U5943 (N_5943,N_3543,N_3345);
and U5944 (N_5944,N_3760,N_2540);
nor U5945 (N_5945,N_4504,N_3223);
or U5946 (N_5946,N_2903,N_4172);
and U5947 (N_5947,N_2804,N_4407);
xor U5948 (N_5948,N_4723,N_3946);
or U5949 (N_5949,N_4984,N_4094);
nand U5950 (N_5950,N_4233,N_4646);
nand U5951 (N_5951,N_2758,N_2521);
nor U5952 (N_5952,N_3162,N_3895);
nand U5953 (N_5953,N_4030,N_2677);
xor U5954 (N_5954,N_4085,N_3254);
nor U5955 (N_5955,N_3243,N_3963);
xor U5956 (N_5956,N_3033,N_4558);
nand U5957 (N_5957,N_2862,N_2635);
nor U5958 (N_5958,N_3967,N_2826);
nor U5959 (N_5959,N_3700,N_4615);
nand U5960 (N_5960,N_3210,N_4952);
nor U5961 (N_5961,N_3947,N_4672);
or U5962 (N_5962,N_2657,N_3721);
nor U5963 (N_5963,N_2591,N_2735);
nand U5964 (N_5964,N_4996,N_3614);
nor U5965 (N_5965,N_4572,N_2958);
or U5966 (N_5966,N_4964,N_4667);
nor U5967 (N_5967,N_2697,N_3433);
nor U5968 (N_5968,N_2578,N_4198);
xnor U5969 (N_5969,N_2929,N_4732);
nand U5970 (N_5970,N_4656,N_4010);
nand U5971 (N_5971,N_3997,N_2593);
nor U5972 (N_5972,N_4870,N_2935);
nor U5973 (N_5973,N_2829,N_3531);
nor U5974 (N_5974,N_2533,N_4761);
and U5975 (N_5975,N_3939,N_3892);
or U5976 (N_5976,N_3273,N_2926);
and U5977 (N_5977,N_3075,N_3517);
xnor U5978 (N_5978,N_3131,N_4351);
or U5979 (N_5979,N_4492,N_3046);
nand U5980 (N_5980,N_4475,N_4157);
and U5981 (N_5981,N_4266,N_3605);
nand U5982 (N_5982,N_3147,N_3296);
or U5983 (N_5983,N_4722,N_3130);
nand U5984 (N_5984,N_3393,N_2594);
and U5985 (N_5985,N_3861,N_3589);
nand U5986 (N_5986,N_3200,N_4370);
or U5987 (N_5987,N_3320,N_3536);
nor U5988 (N_5988,N_3864,N_4268);
and U5989 (N_5989,N_3747,N_4050);
xor U5990 (N_5990,N_3901,N_2788);
xnor U5991 (N_5991,N_3237,N_3577);
nor U5992 (N_5992,N_4711,N_3638);
or U5993 (N_5993,N_4341,N_3428);
xor U5994 (N_5994,N_3971,N_3204);
and U5995 (N_5995,N_4670,N_4922);
and U5996 (N_5996,N_3584,N_4569);
xor U5997 (N_5997,N_4359,N_2632);
nand U5998 (N_5998,N_2688,N_2944);
xnor U5999 (N_5999,N_4057,N_3932);
xnor U6000 (N_6000,N_4129,N_2681);
xnor U6001 (N_6001,N_4696,N_3790);
or U6002 (N_6002,N_3432,N_2864);
or U6003 (N_6003,N_3896,N_2784);
and U6004 (N_6004,N_2640,N_4091);
or U6005 (N_6005,N_4705,N_4036);
or U6006 (N_6006,N_3674,N_4131);
xnor U6007 (N_6007,N_2526,N_4734);
or U6008 (N_6008,N_2702,N_3043);
or U6009 (N_6009,N_3579,N_3585);
or U6010 (N_6010,N_3166,N_3384);
nand U6011 (N_6011,N_4574,N_3768);
nand U6012 (N_6012,N_4827,N_4619);
and U6013 (N_6013,N_2924,N_2982);
xor U6014 (N_6014,N_4812,N_4208);
nand U6015 (N_6015,N_2777,N_4986);
and U6016 (N_6016,N_3301,N_4698);
xor U6017 (N_6017,N_4890,N_4135);
nand U6018 (N_6018,N_3664,N_4395);
or U6019 (N_6019,N_3772,N_4794);
nand U6020 (N_6020,N_2967,N_3479);
nor U6021 (N_6021,N_4850,N_4508);
nand U6022 (N_6022,N_2819,N_4082);
xnor U6023 (N_6023,N_2824,N_3031);
xor U6024 (N_6024,N_3588,N_4804);
and U6025 (N_6025,N_4038,N_3906);
nand U6026 (N_6026,N_4323,N_4685);
or U6027 (N_6027,N_3236,N_4653);
nor U6028 (N_6028,N_3812,N_2987);
nor U6029 (N_6029,N_4358,N_3087);
or U6030 (N_6030,N_3299,N_3105);
nor U6031 (N_6031,N_3639,N_2773);
and U6032 (N_6032,N_2913,N_2808);
and U6033 (N_6033,N_3871,N_3849);
xnor U6034 (N_6034,N_2840,N_3960);
nand U6035 (N_6035,N_4320,N_4818);
nor U6036 (N_6036,N_4317,N_4075);
or U6037 (N_6037,N_4490,N_3924);
or U6038 (N_6038,N_3847,N_4188);
xor U6039 (N_6039,N_4309,N_3386);
nor U6040 (N_6040,N_3966,N_4706);
xnor U6041 (N_6041,N_3777,N_4876);
xnor U6042 (N_6042,N_3958,N_4100);
nor U6043 (N_6043,N_2745,N_3351);
xnor U6044 (N_6044,N_3102,N_3814);
nand U6045 (N_6045,N_4451,N_2765);
or U6046 (N_6046,N_2839,N_4559);
and U6047 (N_6047,N_3499,N_4146);
nand U6048 (N_6048,N_3057,N_3592);
and U6049 (N_6049,N_3181,N_3786);
nor U6050 (N_6050,N_3330,N_3197);
nor U6051 (N_6051,N_4972,N_3561);
nand U6052 (N_6052,N_2549,N_3482);
nor U6053 (N_6053,N_3226,N_4543);
nor U6054 (N_6054,N_4453,N_3109);
and U6055 (N_6055,N_3961,N_4658);
nand U6056 (N_6056,N_4970,N_2539);
nand U6057 (N_6057,N_4186,N_3987);
or U6058 (N_6058,N_3417,N_3569);
nor U6059 (N_6059,N_2642,N_4603);
nand U6060 (N_6060,N_4213,N_3749);
and U6061 (N_6061,N_3221,N_4632);
nor U6062 (N_6062,N_4229,N_3304);
or U6063 (N_6063,N_2671,N_4125);
nor U6064 (N_6064,N_3138,N_4218);
xnor U6065 (N_6065,N_3581,N_3711);
xor U6066 (N_6066,N_4836,N_4961);
xnor U6067 (N_6067,N_4770,N_2976);
xor U6068 (N_6068,N_3689,N_4829);
nor U6069 (N_6069,N_3899,N_3026);
or U6070 (N_6070,N_4806,N_2869);
nand U6071 (N_6071,N_3846,N_4252);
nand U6072 (N_6072,N_4355,N_2989);
nor U6073 (N_6073,N_3770,N_4294);
nand U6074 (N_6074,N_4874,N_4613);
nor U6075 (N_6075,N_4948,N_4334);
nand U6076 (N_6076,N_3680,N_2660);
xor U6077 (N_6077,N_2616,N_4547);
or U6078 (N_6078,N_3258,N_4771);
or U6079 (N_6079,N_3905,N_4993);
and U6080 (N_6080,N_3365,N_2778);
and U6081 (N_6081,N_4464,N_4522);
or U6082 (N_6082,N_3502,N_2576);
or U6083 (N_6083,N_4083,N_4635);
and U6084 (N_6084,N_4312,N_2722);
and U6085 (N_6085,N_2865,N_2644);
and U6086 (N_6086,N_4400,N_3045);
nand U6087 (N_6087,N_2857,N_3385);
xnor U6088 (N_6088,N_3547,N_2631);
nor U6089 (N_6089,N_3521,N_4764);
xnor U6090 (N_6090,N_3356,N_4702);
or U6091 (N_6091,N_4064,N_2902);
or U6092 (N_6092,N_3648,N_3219);
or U6093 (N_6093,N_4254,N_3438);
nand U6094 (N_6094,N_4387,N_4376);
and U6095 (N_6095,N_4708,N_4852);
nor U6096 (N_6096,N_4393,N_3133);
nor U6097 (N_6097,N_3607,N_2651);
xor U6098 (N_6098,N_3513,N_2659);
or U6099 (N_6099,N_3672,N_3103);
nor U6100 (N_6100,N_4758,N_4891);
xnor U6101 (N_6101,N_2817,N_4765);
and U6102 (N_6102,N_3514,N_3288);
and U6103 (N_6103,N_3894,N_4556);
or U6104 (N_6104,N_2752,N_3975);
nand U6105 (N_6105,N_3388,N_3141);
nand U6106 (N_6106,N_4921,N_4417);
nand U6107 (N_6107,N_4352,N_4590);
nand U6108 (N_6108,N_3032,N_3143);
nor U6109 (N_6109,N_4624,N_3354);
and U6110 (N_6110,N_3360,N_3355);
nor U6111 (N_6111,N_4517,N_4554);
nor U6112 (N_6112,N_4410,N_3798);
xor U6113 (N_6113,N_4209,N_4447);
nand U6114 (N_6114,N_2963,N_2620);
and U6115 (N_6115,N_3477,N_4641);
xnor U6116 (N_6116,N_3183,N_3553);
and U6117 (N_6117,N_4398,N_4595);
nand U6118 (N_6118,N_3862,N_4907);
nand U6119 (N_6119,N_4223,N_3993);
nor U6120 (N_6120,N_4709,N_3001);
nor U6121 (N_6121,N_4749,N_2553);
nor U6122 (N_6122,N_3488,N_4663);
and U6123 (N_6123,N_4599,N_3430);
xnor U6124 (N_6124,N_3286,N_3445);
and U6125 (N_6125,N_3039,N_3873);
and U6126 (N_6126,N_3035,N_2689);
and U6127 (N_6127,N_3119,N_4811);
and U6128 (N_6128,N_2988,N_4069);
or U6129 (N_6129,N_3136,N_4872);
xnor U6130 (N_6130,N_3241,N_4614);
or U6131 (N_6131,N_3890,N_3558);
or U6132 (N_6132,N_3776,N_4216);
nand U6133 (N_6133,N_4518,N_2727);
or U6134 (N_6134,N_4725,N_2547);
xor U6135 (N_6135,N_4134,N_4851);
nand U6136 (N_6136,N_3370,N_4187);
xnor U6137 (N_6137,N_4024,N_4023);
xnor U6138 (N_6138,N_4110,N_2833);
or U6139 (N_6139,N_2568,N_2922);
and U6140 (N_6140,N_3728,N_4043);
xor U6141 (N_6141,N_3317,N_2648);
and U6142 (N_6142,N_3501,N_3015);
xnor U6143 (N_6143,N_3014,N_3912);
nor U6144 (N_6144,N_2575,N_3991);
nor U6145 (N_6145,N_4371,N_2615);
or U6146 (N_6146,N_3453,N_3566);
and U6147 (N_6147,N_4005,N_4767);
xnor U6148 (N_6148,N_3319,N_2710);
and U6149 (N_6149,N_4655,N_2686);
nand U6150 (N_6150,N_3256,N_4887);
and U6151 (N_6151,N_2968,N_2836);
nor U6152 (N_6152,N_4425,N_2973);
nor U6153 (N_6153,N_3891,N_2859);
and U6154 (N_6154,N_4394,N_4331);
xnor U6155 (N_6155,N_2717,N_3199);
nor U6156 (N_6156,N_3037,N_4781);
nand U6157 (N_6157,N_2668,N_4444);
nor U6158 (N_6158,N_4476,N_4788);
xnor U6159 (N_6159,N_3332,N_4428);
and U6160 (N_6160,N_4071,N_4090);
or U6161 (N_6161,N_4193,N_2966);
and U6162 (N_6162,N_2936,N_4933);
and U6163 (N_6163,N_3831,N_3407);
nand U6164 (N_6164,N_4166,N_3781);
xor U6165 (N_6165,N_3020,N_3084);
nor U6166 (N_6166,N_3218,N_4037);
or U6167 (N_6167,N_3764,N_3850);
or U6168 (N_6168,N_3444,N_4526);
xor U6169 (N_6169,N_2767,N_2621);
or U6170 (N_6170,N_4427,N_2532);
nor U6171 (N_6171,N_3808,N_3377);
or U6172 (N_6172,N_3580,N_4150);
nor U6173 (N_6173,N_4637,N_3173);
or U6174 (N_6174,N_3268,N_3111);
nand U6175 (N_6175,N_2952,N_4929);
or U6176 (N_6176,N_4390,N_3827);
nand U6177 (N_6177,N_4456,N_2939);
and U6178 (N_6178,N_3845,N_2818);
nor U6179 (N_6179,N_2609,N_4527);
nand U6180 (N_6180,N_3550,N_4074);
nand U6181 (N_6181,N_3886,N_3148);
xnor U6182 (N_6182,N_2600,N_4678);
or U6183 (N_6183,N_4730,N_3406);
or U6184 (N_6184,N_4867,N_2947);
xor U6185 (N_6185,N_4710,N_3503);
nor U6186 (N_6186,N_4833,N_3346);
and U6187 (N_6187,N_4006,N_4742);
xor U6188 (N_6188,N_3796,N_2787);
xor U6189 (N_6189,N_2954,N_2684);
xor U6190 (N_6190,N_3353,N_4324);
nand U6191 (N_6191,N_2557,N_4735);
xnor U6192 (N_6192,N_4032,N_2768);
xnor U6193 (N_6193,N_3629,N_4381);
nand U6194 (N_6194,N_4072,N_3800);
nor U6195 (N_6195,N_2852,N_3253);
nand U6196 (N_6196,N_4489,N_4703);
xor U6197 (N_6197,N_4042,N_2972);
or U6198 (N_6198,N_4076,N_2662);
nand U6199 (N_6199,N_4012,N_4041);
or U6200 (N_6200,N_3792,N_2675);
nor U6201 (N_6201,N_4478,N_4689);
nand U6202 (N_6202,N_3170,N_3127);
and U6203 (N_6203,N_4415,N_3839);
and U6204 (N_6204,N_2931,N_3339);
xor U6205 (N_6205,N_2693,N_3889);
nand U6206 (N_6206,N_4227,N_2598);
or U6207 (N_6207,N_3154,N_4529);
nand U6208 (N_6208,N_3636,N_2909);
or U6209 (N_6209,N_2679,N_4373);
nand U6210 (N_6210,N_2714,N_4446);
nor U6211 (N_6211,N_3787,N_3191);
nand U6212 (N_6212,N_2753,N_2844);
and U6213 (N_6213,N_4817,N_3703);
and U6214 (N_6214,N_3425,N_3418);
or U6215 (N_6215,N_4636,N_4548);
nor U6216 (N_6216,N_4140,N_4528);
and U6217 (N_6217,N_3121,N_4642);
and U6218 (N_6218,N_2831,N_4568);
or U6219 (N_6219,N_3089,N_3532);
or U6220 (N_6220,N_3855,N_4924);
and U6221 (N_6221,N_3656,N_3534);
nand U6222 (N_6222,N_2706,N_3209);
nor U6223 (N_6223,N_3560,N_2619);
and U6224 (N_6224,N_3900,N_4202);
and U6225 (N_6225,N_4983,N_2812);
nor U6226 (N_6226,N_4099,N_4419);
or U6227 (N_6227,N_3073,N_4680);
and U6228 (N_6228,N_4712,N_4343);
nand U6229 (N_6229,N_4067,N_3144);
or U6230 (N_6230,N_3160,N_4237);
xor U6231 (N_6231,N_3833,N_3321);
and U6232 (N_6232,N_3752,N_3494);
nor U6233 (N_6233,N_3743,N_4063);
nor U6234 (N_6234,N_4889,N_4204);
xor U6235 (N_6235,N_4018,N_3999);
xnor U6236 (N_6236,N_3759,N_3666);
nand U6237 (N_6237,N_3628,N_4691);
and U6238 (N_6238,N_3829,N_4337);
or U6239 (N_6239,N_3904,N_3372);
nand U6240 (N_6240,N_3715,N_4631);
or U6241 (N_6241,N_4246,N_3699);
nor U6242 (N_6242,N_4757,N_3238);
xnor U6243 (N_6243,N_3025,N_4299);
nor U6244 (N_6244,N_3439,N_2618);
and U6245 (N_6245,N_4318,N_2505);
and U6246 (N_6246,N_4819,N_4300);
or U6247 (N_6247,N_2979,N_4968);
nand U6248 (N_6248,N_4942,N_4581);
nand U6249 (N_6249,N_3837,N_3970);
or U6250 (N_6250,N_3219,N_4085);
and U6251 (N_6251,N_4859,N_3948);
and U6252 (N_6252,N_3992,N_4250);
or U6253 (N_6253,N_2963,N_2538);
nor U6254 (N_6254,N_4697,N_4853);
and U6255 (N_6255,N_4246,N_3643);
xnor U6256 (N_6256,N_4712,N_2531);
and U6257 (N_6257,N_4496,N_2805);
nand U6258 (N_6258,N_4664,N_2715);
nand U6259 (N_6259,N_2759,N_3518);
nor U6260 (N_6260,N_4397,N_2612);
and U6261 (N_6261,N_2948,N_3985);
xnor U6262 (N_6262,N_4485,N_3712);
nor U6263 (N_6263,N_3090,N_3955);
nand U6264 (N_6264,N_4062,N_3501);
and U6265 (N_6265,N_2713,N_2732);
nand U6266 (N_6266,N_3822,N_4214);
nand U6267 (N_6267,N_3330,N_3151);
xor U6268 (N_6268,N_3754,N_4361);
nor U6269 (N_6269,N_3373,N_3206);
nor U6270 (N_6270,N_4734,N_2854);
nor U6271 (N_6271,N_4841,N_3683);
and U6272 (N_6272,N_3001,N_4722);
and U6273 (N_6273,N_3157,N_2513);
or U6274 (N_6274,N_4134,N_3235);
or U6275 (N_6275,N_4907,N_2538);
nor U6276 (N_6276,N_3205,N_4902);
nor U6277 (N_6277,N_2706,N_3034);
nor U6278 (N_6278,N_4421,N_3176);
xor U6279 (N_6279,N_4211,N_3958);
nand U6280 (N_6280,N_4824,N_3271);
or U6281 (N_6281,N_3153,N_4173);
xnor U6282 (N_6282,N_2863,N_4700);
nand U6283 (N_6283,N_3087,N_4451);
nand U6284 (N_6284,N_2715,N_3827);
or U6285 (N_6285,N_4353,N_3287);
or U6286 (N_6286,N_3055,N_3261);
and U6287 (N_6287,N_3586,N_3624);
or U6288 (N_6288,N_2835,N_3380);
and U6289 (N_6289,N_3097,N_3697);
and U6290 (N_6290,N_2889,N_4600);
nor U6291 (N_6291,N_3370,N_4113);
or U6292 (N_6292,N_3752,N_2879);
nand U6293 (N_6293,N_2531,N_3919);
nand U6294 (N_6294,N_2798,N_2970);
or U6295 (N_6295,N_3413,N_3012);
and U6296 (N_6296,N_4694,N_3756);
and U6297 (N_6297,N_3074,N_3286);
or U6298 (N_6298,N_4045,N_2764);
xor U6299 (N_6299,N_4261,N_4018);
nor U6300 (N_6300,N_3472,N_2691);
nand U6301 (N_6301,N_4147,N_3599);
nand U6302 (N_6302,N_3171,N_3368);
and U6303 (N_6303,N_4016,N_4797);
or U6304 (N_6304,N_3819,N_3723);
nand U6305 (N_6305,N_4642,N_3397);
nand U6306 (N_6306,N_3324,N_2586);
xor U6307 (N_6307,N_4190,N_3504);
xor U6308 (N_6308,N_4216,N_4775);
and U6309 (N_6309,N_4751,N_3462);
or U6310 (N_6310,N_4728,N_3095);
and U6311 (N_6311,N_2885,N_4647);
or U6312 (N_6312,N_4474,N_3228);
nor U6313 (N_6313,N_4921,N_2873);
xnor U6314 (N_6314,N_4167,N_3192);
xor U6315 (N_6315,N_4664,N_3563);
or U6316 (N_6316,N_4767,N_4330);
and U6317 (N_6317,N_4795,N_4628);
and U6318 (N_6318,N_3946,N_3035);
nand U6319 (N_6319,N_3436,N_3432);
or U6320 (N_6320,N_3446,N_2799);
xnor U6321 (N_6321,N_4649,N_3502);
nand U6322 (N_6322,N_3882,N_3007);
xor U6323 (N_6323,N_3967,N_4445);
nor U6324 (N_6324,N_4627,N_4843);
nor U6325 (N_6325,N_3476,N_2590);
or U6326 (N_6326,N_4352,N_2636);
xor U6327 (N_6327,N_3303,N_2747);
xnor U6328 (N_6328,N_3818,N_3682);
nand U6329 (N_6329,N_3993,N_3312);
nand U6330 (N_6330,N_4856,N_3010);
nand U6331 (N_6331,N_2546,N_4193);
or U6332 (N_6332,N_3737,N_3622);
or U6333 (N_6333,N_3776,N_2602);
nand U6334 (N_6334,N_3660,N_3664);
xnor U6335 (N_6335,N_3910,N_3601);
or U6336 (N_6336,N_4065,N_3166);
and U6337 (N_6337,N_2817,N_3436);
nor U6338 (N_6338,N_4462,N_4723);
nor U6339 (N_6339,N_2775,N_3602);
and U6340 (N_6340,N_3219,N_2604);
nand U6341 (N_6341,N_4467,N_4634);
nand U6342 (N_6342,N_2916,N_4712);
xor U6343 (N_6343,N_3692,N_3369);
xor U6344 (N_6344,N_3950,N_2996);
and U6345 (N_6345,N_2644,N_3062);
nand U6346 (N_6346,N_3813,N_2755);
xor U6347 (N_6347,N_3488,N_4561);
nand U6348 (N_6348,N_4793,N_2552);
nand U6349 (N_6349,N_3576,N_3207);
nand U6350 (N_6350,N_2716,N_3816);
nand U6351 (N_6351,N_4137,N_4661);
nand U6352 (N_6352,N_4455,N_2903);
and U6353 (N_6353,N_3263,N_2784);
nor U6354 (N_6354,N_3837,N_4786);
nand U6355 (N_6355,N_2858,N_4265);
nand U6356 (N_6356,N_2776,N_2564);
xnor U6357 (N_6357,N_2705,N_4723);
nor U6358 (N_6358,N_4430,N_2871);
or U6359 (N_6359,N_2975,N_2911);
or U6360 (N_6360,N_4166,N_3569);
xor U6361 (N_6361,N_3166,N_3242);
xnor U6362 (N_6362,N_3539,N_3968);
nor U6363 (N_6363,N_3270,N_3871);
xnor U6364 (N_6364,N_3452,N_2737);
nor U6365 (N_6365,N_2661,N_2973);
or U6366 (N_6366,N_3822,N_2755);
and U6367 (N_6367,N_3804,N_4227);
xnor U6368 (N_6368,N_4861,N_2541);
xnor U6369 (N_6369,N_4575,N_4851);
nor U6370 (N_6370,N_2965,N_4555);
or U6371 (N_6371,N_4379,N_4386);
xnor U6372 (N_6372,N_3380,N_3169);
nand U6373 (N_6373,N_2652,N_4784);
or U6374 (N_6374,N_4249,N_4122);
nand U6375 (N_6375,N_4343,N_2872);
nand U6376 (N_6376,N_2893,N_4850);
or U6377 (N_6377,N_3006,N_2896);
nand U6378 (N_6378,N_2608,N_2729);
nor U6379 (N_6379,N_3693,N_3657);
nor U6380 (N_6380,N_3010,N_4241);
nor U6381 (N_6381,N_3600,N_4909);
nor U6382 (N_6382,N_2639,N_4958);
nand U6383 (N_6383,N_4294,N_4561);
xor U6384 (N_6384,N_2818,N_3679);
nand U6385 (N_6385,N_4382,N_2661);
nor U6386 (N_6386,N_4859,N_3888);
nand U6387 (N_6387,N_3440,N_4207);
nor U6388 (N_6388,N_3808,N_3869);
xor U6389 (N_6389,N_3305,N_2608);
nor U6390 (N_6390,N_2857,N_4996);
nor U6391 (N_6391,N_2742,N_4370);
or U6392 (N_6392,N_4502,N_3935);
xor U6393 (N_6393,N_4926,N_4109);
or U6394 (N_6394,N_4546,N_3501);
nand U6395 (N_6395,N_4240,N_3531);
or U6396 (N_6396,N_3415,N_3527);
nor U6397 (N_6397,N_3204,N_4473);
nor U6398 (N_6398,N_3908,N_3607);
xnor U6399 (N_6399,N_4553,N_3267);
xor U6400 (N_6400,N_3932,N_3885);
or U6401 (N_6401,N_4231,N_2589);
and U6402 (N_6402,N_2650,N_4921);
or U6403 (N_6403,N_3638,N_4135);
and U6404 (N_6404,N_2614,N_4813);
and U6405 (N_6405,N_4205,N_2547);
and U6406 (N_6406,N_3894,N_4940);
xor U6407 (N_6407,N_4668,N_3214);
nand U6408 (N_6408,N_3443,N_2760);
or U6409 (N_6409,N_3044,N_4472);
xor U6410 (N_6410,N_4704,N_4151);
xor U6411 (N_6411,N_4627,N_4932);
nor U6412 (N_6412,N_4585,N_3050);
nand U6413 (N_6413,N_3666,N_2902);
and U6414 (N_6414,N_2596,N_3890);
or U6415 (N_6415,N_3120,N_4753);
nand U6416 (N_6416,N_4414,N_3609);
nand U6417 (N_6417,N_2768,N_3531);
or U6418 (N_6418,N_2771,N_2557);
or U6419 (N_6419,N_4260,N_4831);
or U6420 (N_6420,N_2858,N_3068);
nand U6421 (N_6421,N_3159,N_3172);
xor U6422 (N_6422,N_4313,N_2756);
xor U6423 (N_6423,N_4898,N_4156);
or U6424 (N_6424,N_4464,N_2750);
or U6425 (N_6425,N_4751,N_4308);
nand U6426 (N_6426,N_4911,N_4217);
nor U6427 (N_6427,N_3879,N_4248);
xnor U6428 (N_6428,N_3816,N_3932);
nand U6429 (N_6429,N_4808,N_4689);
nor U6430 (N_6430,N_2633,N_3340);
xor U6431 (N_6431,N_3767,N_3525);
or U6432 (N_6432,N_4086,N_4130);
nor U6433 (N_6433,N_3794,N_3194);
xor U6434 (N_6434,N_4419,N_2984);
nand U6435 (N_6435,N_4195,N_4422);
or U6436 (N_6436,N_2850,N_3685);
nand U6437 (N_6437,N_4351,N_4781);
or U6438 (N_6438,N_2851,N_4127);
nor U6439 (N_6439,N_3341,N_4666);
and U6440 (N_6440,N_3328,N_4406);
and U6441 (N_6441,N_4536,N_2766);
nor U6442 (N_6442,N_3393,N_2778);
and U6443 (N_6443,N_2880,N_3873);
or U6444 (N_6444,N_3020,N_4898);
nand U6445 (N_6445,N_4255,N_3565);
nand U6446 (N_6446,N_4810,N_2909);
nand U6447 (N_6447,N_3122,N_4323);
or U6448 (N_6448,N_3323,N_3520);
and U6449 (N_6449,N_3620,N_3826);
or U6450 (N_6450,N_4180,N_3581);
nand U6451 (N_6451,N_4654,N_4281);
nor U6452 (N_6452,N_3911,N_2564);
xor U6453 (N_6453,N_4218,N_3388);
and U6454 (N_6454,N_2825,N_4653);
nand U6455 (N_6455,N_4127,N_4789);
nor U6456 (N_6456,N_4766,N_4527);
and U6457 (N_6457,N_4393,N_3852);
xor U6458 (N_6458,N_2908,N_3500);
xor U6459 (N_6459,N_4364,N_2543);
xor U6460 (N_6460,N_3301,N_2672);
xor U6461 (N_6461,N_4152,N_3538);
or U6462 (N_6462,N_3164,N_2536);
and U6463 (N_6463,N_4102,N_3703);
nand U6464 (N_6464,N_4754,N_4300);
nor U6465 (N_6465,N_4635,N_4193);
and U6466 (N_6466,N_3527,N_3641);
xor U6467 (N_6467,N_3723,N_4535);
or U6468 (N_6468,N_3665,N_2787);
and U6469 (N_6469,N_3050,N_4122);
or U6470 (N_6470,N_3314,N_4988);
or U6471 (N_6471,N_3203,N_3466);
nand U6472 (N_6472,N_4453,N_4307);
xnor U6473 (N_6473,N_3373,N_4966);
and U6474 (N_6474,N_4791,N_4414);
or U6475 (N_6475,N_3703,N_3378);
xnor U6476 (N_6476,N_4251,N_3078);
and U6477 (N_6477,N_4977,N_3028);
nor U6478 (N_6478,N_3111,N_2639);
xnor U6479 (N_6479,N_2901,N_3053);
and U6480 (N_6480,N_4584,N_2594);
nor U6481 (N_6481,N_4192,N_4144);
and U6482 (N_6482,N_4729,N_2625);
nor U6483 (N_6483,N_2583,N_3487);
nor U6484 (N_6484,N_4095,N_2959);
and U6485 (N_6485,N_3061,N_3397);
and U6486 (N_6486,N_3077,N_3072);
and U6487 (N_6487,N_2794,N_4943);
and U6488 (N_6488,N_2680,N_3985);
or U6489 (N_6489,N_4774,N_4093);
or U6490 (N_6490,N_3257,N_4023);
nor U6491 (N_6491,N_2843,N_3017);
nand U6492 (N_6492,N_3814,N_2566);
nand U6493 (N_6493,N_3174,N_4225);
xor U6494 (N_6494,N_4310,N_3535);
or U6495 (N_6495,N_2661,N_4015);
nand U6496 (N_6496,N_4917,N_4130);
and U6497 (N_6497,N_4454,N_4603);
or U6498 (N_6498,N_3485,N_2840);
nor U6499 (N_6499,N_4568,N_3919);
xor U6500 (N_6500,N_4437,N_3163);
xnor U6501 (N_6501,N_4421,N_2875);
and U6502 (N_6502,N_3748,N_2547);
nor U6503 (N_6503,N_2907,N_4087);
xnor U6504 (N_6504,N_3394,N_4764);
nor U6505 (N_6505,N_4898,N_4311);
nor U6506 (N_6506,N_2959,N_3938);
nor U6507 (N_6507,N_2506,N_4846);
nor U6508 (N_6508,N_2560,N_3445);
xnor U6509 (N_6509,N_3125,N_3963);
nand U6510 (N_6510,N_3706,N_2683);
nor U6511 (N_6511,N_2715,N_4384);
and U6512 (N_6512,N_2692,N_4305);
nand U6513 (N_6513,N_3018,N_3251);
nand U6514 (N_6514,N_2867,N_2805);
xnor U6515 (N_6515,N_4783,N_4791);
and U6516 (N_6516,N_2511,N_2966);
xor U6517 (N_6517,N_4905,N_4706);
nand U6518 (N_6518,N_4289,N_3649);
and U6519 (N_6519,N_3164,N_3582);
and U6520 (N_6520,N_4353,N_4424);
xor U6521 (N_6521,N_4150,N_3632);
nor U6522 (N_6522,N_3453,N_2963);
nand U6523 (N_6523,N_2658,N_4537);
and U6524 (N_6524,N_3384,N_3726);
xor U6525 (N_6525,N_4947,N_2788);
nor U6526 (N_6526,N_3769,N_3309);
xnor U6527 (N_6527,N_4116,N_4857);
nand U6528 (N_6528,N_4457,N_3832);
nand U6529 (N_6529,N_2875,N_4551);
nor U6530 (N_6530,N_4454,N_3137);
or U6531 (N_6531,N_4003,N_3533);
and U6532 (N_6532,N_3135,N_4585);
and U6533 (N_6533,N_4601,N_3441);
or U6534 (N_6534,N_3236,N_2909);
xor U6535 (N_6535,N_3867,N_2782);
xor U6536 (N_6536,N_3248,N_4059);
xor U6537 (N_6537,N_4023,N_3282);
xnor U6538 (N_6538,N_2753,N_4462);
nor U6539 (N_6539,N_4162,N_3393);
xor U6540 (N_6540,N_4691,N_3727);
nor U6541 (N_6541,N_3846,N_3639);
xnor U6542 (N_6542,N_4577,N_3118);
or U6543 (N_6543,N_4629,N_3651);
or U6544 (N_6544,N_2701,N_2691);
and U6545 (N_6545,N_4736,N_4302);
nand U6546 (N_6546,N_4906,N_3920);
nand U6547 (N_6547,N_4178,N_3233);
or U6548 (N_6548,N_3142,N_4076);
nor U6549 (N_6549,N_4390,N_2936);
and U6550 (N_6550,N_2972,N_3674);
xor U6551 (N_6551,N_3811,N_3477);
xnor U6552 (N_6552,N_3051,N_2883);
and U6553 (N_6553,N_4322,N_3383);
nor U6554 (N_6554,N_4193,N_4636);
nand U6555 (N_6555,N_3026,N_3381);
nand U6556 (N_6556,N_4124,N_3300);
and U6557 (N_6557,N_4915,N_3937);
or U6558 (N_6558,N_4853,N_4319);
nand U6559 (N_6559,N_4218,N_4868);
and U6560 (N_6560,N_3314,N_4419);
xor U6561 (N_6561,N_3329,N_4716);
nor U6562 (N_6562,N_3110,N_3074);
nor U6563 (N_6563,N_2602,N_3551);
xor U6564 (N_6564,N_3732,N_3816);
nand U6565 (N_6565,N_3663,N_3299);
or U6566 (N_6566,N_2826,N_2827);
xor U6567 (N_6567,N_4164,N_4193);
or U6568 (N_6568,N_3388,N_2590);
and U6569 (N_6569,N_3242,N_3750);
or U6570 (N_6570,N_3091,N_3226);
and U6571 (N_6571,N_4727,N_3885);
and U6572 (N_6572,N_2990,N_3213);
and U6573 (N_6573,N_4879,N_3177);
and U6574 (N_6574,N_3260,N_3338);
xor U6575 (N_6575,N_3177,N_3251);
and U6576 (N_6576,N_4892,N_4434);
and U6577 (N_6577,N_3649,N_4766);
or U6578 (N_6578,N_4796,N_4329);
xor U6579 (N_6579,N_4925,N_4517);
nor U6580 (N_6580,N_4686,N_3099);
nand U6581 (N_6581,N_4917,N_4670);
or U6582 (N_6582,N_3839,N_2699);
and U6583 (N_6583,N_2958,N_2999);
nor U6584 (N_6584,N_2813,N_2694);
and U6585 (N_6585,N_2815,N_4878);
nor U6586 (N_6586,N_4687,N_2984);
nor U6587 (N_6587,N_2782,N_3462);
nor U6588 (N_6588,N_4990,N_4180);
xor U6589 (N_6589,N_2624,N_2540);
xor U6590 (N_6590,N_2702,N_4225);
nand U6591 (N_6591,N_3125,N_3224);
and U6592 (N_6592,N_3785,N_3069);
and U6593 (N_6593,N_3727,N_3079);
or U6594 (N_6594,N_4508,N_4204);
and U6595 (N_6595,N_4718,N_2626);
nand U6596 (N_6596,N_3296,N_2603);
nor U6597 (N_6597,N_3179,N_3585);
nor U6598 (N_6598,N_4656,N_3950);
nor U6599 (N_6599,N_4663,N_4289);
nand U6600 (N_6600,N_4833,N_4479);
and U6601 (N_6601,N_3507,N_2892);
nand U6602 (N_6602,N_4957,N_4928);
nor U6603 (N_6603,N_3287,N_3800);
xor U6604 (N_6604,N_2980,N_3743);
and U6605 (N_6605,N_2965,N_4703);
and U6606 (N_6606,N_2920,N_3108);
nand U6607 (N_6607,N_3924,N_3491);
nand U6608 (N_6608,N_3537,N_4878);
or U6609 (N_6609,N_4873,N_2978);
xnor U6610 (N_6610,N_2503,N_4813);
or U6611 (N_6611,N_4078,N_2860);
and U6612 (N_6612,N_2866,N_3238);
xnor U6613 (N_6613,N_3473,N_2682);
and U6614 (N_6614,N_4365,N_4478);
and U6615 (N_6615,N_2794,N_3210);
or U6616 (N_6616,N_4802,N_4282);
and U6617 (N_6617,N_2842,N_3003);
and U6618 (N_6618,N_3392,N_4583);
xnor U6619 (N_6619,N_3890,N_3591);
nand U6620 (N_6620,N_3535,N_3927);
and U6621 (N_6621,N_3874,N_4140);
xor U6622 (N_6622,N_3970,N_3909);
nand U6623 (N_6623,N_3956,N_4564);
nor U6624 (N_6624,N_3054,N_4443);
xnor U6625 (N_6625,N_4299,N_2909);
or U6626 (N_6626,N_2559,N_3986);
xor U6627 (N_6627,N_3273,N_3768);
nor U6628 (N_6628,N_3425,N_3440);
or U6629 (N_6629,N_2626,N_4092);
nor U6630 (N_6630,N_3937,N_3169);
nand U6631 (N_6631,N_3105,N_3543);
nor U6632 (N_6632,N_2589,N_4506);
nand U6633 (N_6633,N_2658,N_4477);
nor U6634 (N_6634,N_4666,N_2772);
nand U6635 (N_6635,N_2874,N_4543);
or U6636 (N_6636,N_4444,N_4253);
nor U6637 (N_6637,N_3588,N_4829);
and U6638 (N_6638,N_4259,N_3835);
nor U6639 (N_6639,N_3988,N_4745);
xnor U6640 (N_6640,N_4050,N_4612);
or U6641 (N_6641,N_3288,N_4351);
xor U6642 (N_6642,N_4901,N_2978);
xor U6643 (N_6643,N_4952,N_3723);
xor U6644 (N_6644,N_2618,N_4490);
and U6645 (N_6645,N_3351,N_4959);
nand U6646 (N_6646,N_3507,N_2627);
xnor U6647 (N_6647,N_4326,N_4374);
or U6648 (N_6648,N_3029,N_3063);
or U6649 (N_6649,N_4090,N_2563);
and U6650 (N_6650,N_3269,N_3201);
nor U6651 (N_6651,N_2613,N_4810);
or U6652 (N_6652,N_3519,N_2641);
nand U6653 (N_6653,N_2663,N_3368);
nand U6654 (N_6654,N_2726,N_4365);
nand U6655 (N_6655,N_4165,N_3408);
nand U6656 (N_6656,N_3027,N_2677);
and U6657 (N_6657,N_2842,N_4290);
and U6658 (N_6658,N_3307,N_3339);
xor U6659 (N_6659,N_3643,N_4016);
xor U6660 (N_6660,N_3709,N_4559);
or U6661 (N_6661,N_4380,N_4821);
xnor U6662 (N_6662,N_4439,N_2673);
nand U6663 (N_6663,N_3618,N_3534);
or U6664 (N_6664,N_3530,N_4068);
nor U6665 (N_6665,N_3913,N_3369);
nor U6666 (N_6666,N_3219,N_3071);
and U6667 (N_6667,N_4834,N_2793);
or U6668 (N_6668,N_3360,N_2777);
nor U6669 (N_6669,N_4229,N_4149);
nand U6670 (N_6670,N_4993,N_2942);
nor U6671 (N_6671,N_2956,N_2997);
or U6672 (N_6672,N_4667,N_4806);
or U6673 (N_6673,N_3093,N_4344);
nor U6674 (N_6674,N_3020,N_3506);
xnor U6675 (N_6675,N_3983,N_4997);
and U6676 (N_6676,N_4118,N_4468);
xor U6677 (N_6677,N_3417,N_4024);
xnor U6678 (N_6678,N_4734,N_4544);
and U6679 (N_6679,N_3756,N_3783);
xnor U6680 (N_6680,N_3414,N_4566);
nor U6681 (N_6681,N_4463,N_4838);
xor U6682 (N_6682,N_3088,N_3397);
xor U6683 (N_6683,N_3655,N_4999);
nand U6684 (N_6684,N_4141,N_3073);
and U6685 (N_6685,N_4160,N_3119);
nor U6686 (N_6686,N_3635,N_3108);
xor U6687 (N_6687,N_4767,N_3090);
nor U6688 (N_6688,N_3440,N_3190);
nand U6689 (N_6689,N_2934,N_4699);
or U6690 (N_6690,N_4369,N_3035);
or U6691 (N_6691,N_3994,N_4798);
nor U6692 (N_6692,N_3203,N_2920);
nand U6693 (N_6693,N_3644,N_2985);
or U6694 (N_6694,N_4231,N_3978);
and U6695 (N_6695,N_4842,N_3432);
nand U6696 (N_6696,N_4131,N_3233);
nor U6697 (N_6697,N_2919,N_3327);
and U6698 (N_6698,N_4978,N_4788);
or U6699 (N_6699,N_3406,N_3341);
nor U6700 (N_6700,N_3396,N_2930);
and U6701 (N_6701,N_3777,N_2863);
or U6702 (N_6702,N_2783,N_3273);
nand U6703 (N_6703,N_2949,N_4700);
and U6704 (N_6704,N_3253,N_3406);
nand U6705 (N_6705,N_4557,N_3786);
or U6706 (N_6706,N_4135,N_4825);
nor U6707 (N_6707,N_4327,N_2890);
xor U6708 (N_6708,N_4033,N_3887);
or U6709 (N_6709,N_3545,N_3013);
nand U6710 (N_6710,N_4640,N_3288);
and U6711 (N_6711,N_3126,N_2642);
nand U6712 (N_6712,N_3035,N_4972);
and U6713 (N_6713,N_4645,N_4850);
or U6714 (N_6714,N_3839,N_4785);
or U6715 (N_6715,N_2871,N_4193);
and U6716 (N_6716,N_2865,N_3939);
nand U6717 (N_6717,N_3774,N_4118);
xnor U6718 (N_6718,N_4794,N_2683);
or U6719 (N_6719,N_3970,N_2922);
and U6720 (N_6720,N_4151,N_3713);
and U6721 (N_6721,N_4618,N_4284);
or U6722 (N_6722,N_3659,N_2603);
xnor U6723 (N_6723,N_3753,N_4351);
nor U6724 (N_6724,N_3171,N_4188);
nor U6725 (N_6725,N_3673,N_3289);
or U6726 (N_6726,N_4065,N_4989);
xor U6727 (N_6727,N_3195,N_4170);
xor U6728 (N_6728,N_4708,N_2582);
nor U6729 (N_6729,N_4406,N_4646);
or U6730 (N_6730,N_3863,N_2558);
xor U6731 (N_6731,N_4900,N_4156);
nand U6732 (N_6732,N_2742,N_4100);
xor U6733 (N_6733,N_4239,N_4307);
nand U6734 (N_6734,N_2634,N_3632);
or U6735 (N_6735,N_4082,N_4843);
or U6736 (N_6736,N_2543,N_4047);
nor U6737 (N_6737,N_4616,N_4922);
nand U6738 (N_6738,N_2713,N_4734);
or U6739 (N_6739,N_3089,N_4205);
and U6740 (N_6740,N_3025,N_3286);
or U6741 (N_6741,N_4399,N_4341);
and U6742 (N_6742,N_4076,N_2937);
and U6743 (N_6743,N_2915,N_2986);
and U6744 (N_6744,N_2918,N_2774);
xor U6745 (N_6745,N_4582,N_3373);
nor U6746 (N_6746,N_3380,N_2862);
xor U6747 (N_6747,N_3832,N_3303);
or U6748 (N_6748,N_2961,N_4130);
nand U6749 (N_6749,N_4835,N_4089);
or U6750 (N_6750,N_4703,N_4872);
or U6751 (N_6751,N_4622,N_2862);
and U6752 (N_6752,N_4381,N_4179);
or U6753 (N_6753,N_3330,N_2724);
nor U6754 (N_6754,N_3426,N_2568);
nand U6755 (N_6755,N_3098,N_3495);
nand U6756 (N_6756,N_2525,N_4258);
and U6757 (N_6757,N_4765,N_4305);
nor U6758 (N_6758,N_3689,N_3837);
nand U6759 (N_6759,N_4334,N_3127);
and U6760 (N_6760,N_3626,N_4788);
xnor U6761 (N_6761,N_2595,N_4415);
nor U6762 (N_6762,N_4692,N_3035);
or U6763 (N_6763,N_3477,N_3723);
nor U6764 (N_6764,N_3753,N_4142);
and U6765 (N_6765,N_3178,N_3489);
nor U6766 (N_6766,N_3464,N_3024);
and U6767 (N_6767,N_4623,N_4091);
xnor U6768 (N_6768,N_4759,N_4737);
and U6769 (N_6769,N_4350,N_2595);
nor U6770 (N_6770,N_3348,N_2932);
and U6771 (N_6771,N_4051,N_4766);
and U6772 (N_6772,N_3731,N_4124);
and U6773 (N_6773,N_4755,N_2817);
xor U6774 (N_6774,N_3026,N_4989);
or U6775 (N_6775,N_2905,N_3453);
nand U6776 (N_6776,N_2605,N_4412);
nand U6777 (N_6777,N_3702,N_2647);
nor U6778 (N_6778,N_4493,N_4161);
nand U6779 (N_6779,N_3170,N_3593);
xor U6780 (N_6780,N_2681,N_4923);
nor U6781 (N_6781,N_4700,N_3883);
or U6782 (N_6782,N_4513,N_3838);
and U6783 (N_6783,N_3613,N_3195);
and U6784 (N_6784,N_4624,N_4940);
xor U6785 (N_6785,N_3390,N_4851);
or U6786 (N_6786,N_3699,N_3924);
xnor U6787 (N_6787,N_4187,N_4562);
nand U6788 (N_6788,N_4294,N_3329);
xor U6789 (N_6789,N_2802,N_2865);
xor U6790 (N_6790,N_3395,N_3669);
xnor U6791 (N_6791,N_4393,N_3655);
nor U6792 (N_6792,N_2660,N_4612);
and U6793 (N_6793,N_3411,N_4047);
or U6794 (N_6794,N_2798,N_3311);
nor U6795 (N_6795,N_4439,N_4009);
or U6796 (N_6796,N_4913,N_4292);
and U6797 (N_6797,N_3629,N_4034);
xnor U6798 (N_6798,N_3875,N_2597);
nand U6799 (N_6799,N_4734,N_2978);
and U6800 (N_6800,N_3440,N_2633);
and U6801 (N_6801,N_3742,N_4831);
and U6802 (N_6802,N_4064,N_3221);
and U6803 (N_6803,N_2795,N_4159);
or U6804 (N_6804,N_2972,N_3009);
and U6805 (N_6805,N_3170,N_2621);
and U6806 (N_6806,N_4937,N_3183);
xnor U6807 (N_6807,N_4243,N_2943);
nor U6808 (N_6808,N_4518,N_3774);
xor U6809 (N_6809,N_2907,N_3433);
or U6810 (N_6810,N_4867,N_2927);
nor U6811 (N_6811,N_2604,N_3562);
nand U6812 (N_6812,N_3279,N_3329);
nor U6813 (N_6813,N_3198,N_3747);
nand U6814 (N_6814,N_3448,N_3247);
or U6815 (N_6815,N_4891,N_4974);
and U6816 (N_6816,N_3360,N_3549);
xor U6817 (N_6817,N_3365,N_4170);
xor U6818 (N_6818,N_4794,N_3730);
xnor U6819 (N_6819,N_3845,N_4123);
and U6820 (N_6820,N_2611,N_4696);
and U6821 (N_6821,N_4595,N_3015);
and U6822 (N_6822,N_2702,N_3034);
xnor U6823 (N_6823,N_3556,N_3386);
nand U6824 (N_6824,N_3591,N_3022);
nor U6825 (N_6825,N_3578,N_4044);
nand U6826 (N_6826,N_4768,N_4670);
or U6827 (N_6827,N_2726,N_2645);
nand U6828 (N_6828,N_3266,N_4783);
or U6829 (N_6829,N_3080,N_3888);
or U6830 (N_6830,N_2856,N_3929);
nor U6831 (N_6831,N_4309,N_2551);
nor U6832 (N_6832,N_3499,N_3801);
xor U6833 (N_6833,N_3682,N_2633);
or U6834 (N_6834,N_3599,N_4312);
nand U6835 (N_6835,N_4658,N_4108);
nor U6836 (N_6836,N_3809,N_4520);
xor U6837 (N_6837,N_4149,N_4886);
nor U6838 (N_6838,N_3665,N_4300);
or U6839 (N_6839,N_4899,N_4462);
and U6840 (N_6840,N_3560,N_3004);
and U6841 (N_6841,N_3620,N_2731);
xnor U6842 (N_6842,N_3498,N_2944);
nand U6843 (N_6843,N_2832,N_2761);
nor U6844 (N_6844,N_3448,N_4255);
and U6845 (N_6845,N_3970,N_4472);
xor U6846 (N_6846,N_4409,N_3867);
nor U6847 (N_6847,N_4402,N_4048);
xnor U6848 (N_6848,N_2725,N_3099);
nor U6849 (N_6849,N_2776,N_3942);
nor U6850 (N_6850,N_4376,N_3908);
and U6851 (N_6851,N_4246,N_4634);
xnor U6852 (N_6852,N_2824,N_4734);
nand U6853 (N_6853,N_3543,N_3712);
xor U6854 (N_6854,N_4078,N_3901);
xor U6855 (N_6855,N_4247,N_4596);
and U6856 (N_6856,N_4977,N_2712);
and U6857 (N_6857,N_3585,N_2857);
xor U6858 (N_6858,N_3976,N_2565);
nor U6859 (N_6859,N_2767,N_4199);
nor U6860 (N_6860,N_4055,N_4061);
nor U6861 (N_6861,N_3736,N_4902);
nor U6862 (N_6862,N_4794,N_2807);
or U6863 (N_6863,N_3442,N_4636);
xor U6864 (N_6864,N_2638,N_2907);
nor U6865 (N_6865,N_2625,N_4167);
xnor U6866 (N_6866,N_4198,N_4407);
nor U6867 (N_6867,N_4289,N_3396);
or U6868 (N_6868,N_4047,N_4793);
xor U6869 (N_6869,N_4343,N_4588);
or U6870 (N_6870,N_3483,N_3774);
nand U6871 (N_6871,N_2569,N_4977);
nand U6872 (N_6872,N_3343,N_4197);
and U6873 (N_6873,N_2812,N_4649);
nand U6874 (N_6874,N_4492,N_4531);
nor U6875 (N_6875,N_4944,N_4341);
or U6876 (N_6876,N_3715,N_3227);
nor U6877 (N_6877,N_4383,N_4832);
nor U6878 (N_6878,N_3611,N_4904);
nor U6879 (N_6879,N_3853,N_3248);
nand U6880 (N_6880,N_3804,N_3491);
nand U6881 (N_6881,N_4772,N_4775);
and U6882 (N_6882,N_2834,N_3617);
nor U6883 (N_6883,N_4734,N_3835);
xnor U6884 (N_6884,N_3985,N_3601);
nand U6885 (N_6885,N_4219,N_4026);
xor U6886 (N_6886,N_4988,N_4330);
nand U6887 (N_6887,N_3979,N_4811);
xnor U6888 (N_6888,N_4974,N_4561);
nand U6889 (N_6889,N_3670,N_4219);
nor U6890 (N_6890,N_4301,N_4956);
and U6891 (N_6891,N_3134,N_4743);
xnor U6892 (N_6892,N_3646,N_3261);
nand U6893 (N_6893,N_3096,N_2869);
nand U6894 (N_6894,N_2653,N_3077);
nor U6895 (N_6895,N_4791,N_4959);
and U6896 (N_6896,N_4703,N_3529);
nand U6897 (N_6897,N_3946,N_2971);
or U6898 (N_6898,N_2838,N_2743);
nand U6899 (N_6899,N_4348,N_3991);
xnor U6900 (N_6900,N_4534,N_3227);
xnor U6901 (N_6901,N_3020,N_4164);
nand U6902 (N_6902,N_4634,N_3660);
and U6903 (N_6903,N_3395,N_4415);
nand U6904 (N_6904,N_2881,N_3905);
nand U6905 (N_6905,N_2998,N_3329);
and U6906 (N_6906,N_3569,N_4260);
or U6907 (N_6907,N_2673,N_3916);
or U6908 (N_6908,N_3068,N_3779);
nand U6909 (N_6909,N_4295,N_4831);
xnor U6910 (N_6910,N_3616,N_4305);
and U6911 (N_6911,N_2536,N_4503);
xnor U6912 (N_6912,N_2951,N_4632);
and U6913 (N_6913,N_3034,N_4625);
nor U6914 (N_6914,N_4696,N_3304);
xnor U6915 (N_6915,N_3667,N_4474);
and U6916 (N_6916,N_2635,N_3528);
or U6917 (N_6917,N_4518,N_3996);
nor U6918 (N_6918,N_4304,N_2815);
or U6919 (N_6919,N_4561,N_3320);
xor U6920 (N_6920,N_2992,N_4914);
and U6921 (N_6921,N_2520,N_4712);
nand U6922 (N_6922,N_4692,N_4726);
and U6923 (N_6923,N_3172,N_4260);
or U6924 (N_6924,N_2901,N_3391);
and U6925 (N_6925,N_4968,N_3608);
and U6926 (N_6926,N_4367,N_4909);
nand U6927 (N_6927,N_2603,N_2975);
xor U6928 (N_6928,N_4424,N_4156);
and U6929 (N_6929,N_3600,N_4798);
and U6930 (N_6930,N_3216,N_2680);
nand U6931 (N_6931,N_3049,N_4945);
or U6932 (N_6932,N_2889,N_4178);
xnor U6933 (N_6933,N_2593,N_3976);
and U6934 (N_6934,N_3464,N_4196);
nor U6935 (N_6935,N_3791,N_4945);
and U6936 (N_6936,N_4486,N_4614);
nor U6937 (N_6937,N_3862,N_2649);
and U6938 (N_6938,N_4838,N_2878);
nand U6939 (N_6939,N_2926,N_2829);
nor U6940 (N_6940,N_3557,N_3830);
nand U6941 (N_6941,N_2644,N_3014);
or U6942 (N_6942,N_4891,N_3183);
and U6943 (N_6943,N_3273,N_3816);
nor U6944 (N_6944,N_3059,N_3506);
or U6945 (N_6945,N_3266,N_3877);
xnor U6946 (N_6946,N_2639,N_4265);
and U6947 (N_6947,N_4091,N_2523);
or U6948 (N_6948,N_4049,N_3283);
and U6949 (N_6949,N_3505,N_4900);
nor U6950 (N_6950,N_3536,N_2940);
nor U6951 (N_6951,N_4715,N_2993);
nor U6952 (N_6952,N_3270,N_3879);
or U6953 (N_6953,N_4079,N_4187);
nand U6954 (N_6954,N_2893,N_4201);
nor U6955 (N_6955,N_4553,N_3246);
or U6956 (N_6956,N_4455,N_4901);
and U6957 (N_6957,N_4513,N_2688);
nor U6958 (N_6958,N_2510,N_3906);
nand U6959 (N_6959,N_2728,N_2836);
and U6960 (N_6960,N_2872,N_4502);
nand U6961 (N_6961,N_4131,N_2675);
nand U6962 (N_6962,N_3545,N_4025);
nand U6963 (N_6963,N_3652,N_4424);
and U6964 (N_6964,N_4335,N_2888);
nand U6965 (N_6965,N_3588,N_3501);
nor U6966 (N_6966,N_4083,N_4136);
nand U6967 (N_6967,N_2753,N_3558);
or U6968 (N_6968,N_3591,N_4857);
or U6969 (N_6969,N_3933,N_3965);
xor U6970 (N_6970,N_3756,N_3105);
and U6971 (N_6971,N_3706,N_3182);
nand U6972 (N_6972,N_4908,N_3490);
xor U6973 (N_6973,N_4710,N_2639);
and U6974 (N_6974,N_4356,N_3597);
xnor U6975 (N_6975,N_3021,N_4623);
and U6976 (N_6976,N_4243,N_2765);
xor U6977 (N_6977,N_3731,N_2640);
xor U6978 (N_6978,N_4043,N_4501);
xor U6979 (N_6979,N_3105,N_4734);
and U6980 (N_6980,N_4476,N_3508);
nand U6981 (N_6981,N_4345,N_3503);
or U6982 (N_6982,N_2873,N_3217);
and U6983 (N_6983,N_3267,N_2858);
nor U6984 (N_6984,N_2572,N_2840);
and U6985 (N_6985,N_3713,N_3583);
and U6986 (N_6986,N_4539,N_4080);
nor U6987 (N_6987,N_3642,N_4141);
nor U6988 (N_6988,N_2712,N_2648);
xnor U6989 (N_6989,N_4473,N_4053);
nor U6990 (N_6990,N_4390,N_3033);
nor U6991 (N_6991,N_2861,N_2526);
or U6992 (N_6992,N_2603,N_2596);
or U6993 (N_6993,N_3200,N_2700);
or U6994 (N_6994,N_4827,N_3477);
xnor U6995 (N_6995,N_4657,N_2537);
nand U6996 (N_6996,N_3951,N_4312);
nand U6997 (N_6997,N_4803,N_4684);
nor U6998 (N_6998,N_3502,N_3595);
nand U6999 (N_6999,N_4490,N_2721);
nor U7000 (N_7000,N_4356,N_3555);
xor U7001 (N_7001,N_4151,N_2530);
nand U7002 (N_7002,N_3162,N_3664);
nor U7003 (N_7003,N_3792,N_3993);
and U7004 (N_7004,N_4183,N_3600);
nor U7005 (N_7005,N_4263,N_2925);
nand U7006 (N_7006,N_3240,N_3734);
nor U7007 (N_7007,N_3240,N_3453);
xnor U7008 (N_7008,N_3606,N_4749);
nor U7009 (N_7009,N_4004,N_2829);
nand U7010 (N_7010,N_4606,N_3685);
and U7011 (N_7011,N_3234,N_2663);
nor U7012 (N_7012,N_3023,N_3669);
xor U7013 (N_7013,N_4311,N_4267);
and U7014 (N_7014,N_3181,N_2942);
nand U7015 (N_7015,N_2840,N_3328);
xor U7016 (N_7016,N_3978,N_3543);
and U7017 (N_7017,N_3756,N_4918);
and U7018 (N_7018,N_2722,N_2951);
nand U7019 (N_7019,N_2742,N_3995);
nand U7020 (N_7020,N_4959,N_3898);
xnor U7021 (N_7021,N_3751,N_3497);
or U7022 (N_7022,N_2753,N_3098);
or U7023 (N_7023,N_2881,N_4381);
nor U7024 (N_7024,N_4710,N_4039);
nor U7025 (N_7025,N_3868,N_3627);
or U7026 (N_7026,N_2840,N_3194);
nor U7027 (N_7027,N_2564,N_4941);
nor U7028 (N_7028,N_2522,N_2779);
and U7029 (N_7029,N_3058,N_4510);
xnor U7030 (N_7030,N_4761,N_4804);
and U7031 (N_7031,N_4578,N_3263);
and U7032 (N_7032,N_3154,N_3741);
or U7033 (N_7033,N_2794,N_2538);
nand U7034 (N_7034,N_2893,N_3197);
nand U7035 (N_7035,N_4777,N_4958);
nor U7036 (N_7036,N_4642,N_2518);
and U7037 (N_7037,N_4445,N_3218);
or U7038 (N_7038,N_3879,N_3030);
nor U7039 (N_7039,N_4677,N_4738);
or U7040 (N_7040,N_2741,N_4622);
nand U7041 (N_7041,N_4099,N_4226);
nor U7042 (N_7042,N_3114,N_4564);
xnor U7043 (N_7043,N_3151,N_3284);
nand U7044 (N_7044,N_3872,N_3720);
nor U7045 (N_7045,N_3896,N_3903);
nor U7046 (N_7046,N_3181,N_2960);
nand U7047 (N_7047,N_3363,N_4649);
xnor U7048 (N_7048,N_4246,N_2721);
nand U7049 (N_7049,N_4064,N_2700);
and U7050 (N_7050,N_3957,N_4797);
nor U7051 (N_7051,N_3382,N_4900);
xnor U7052 (N_7052,N_4741,N_4342);
and U7053 (N_7053,N_2607,N_4568);
nand U7054 (N_7054,N_3214,N_3064);
nand U7055 (N_7055,N_2721,N_3767);
or U7056 (N_7056,N_4190,N_3312);
and U7057 (N_7057,N_3629,N_3023);
and U7058 (N_7058,N_3044,N_4486);
xnor U7059 (N_7059,N_4546,N_4583);
nor U7060 (N_7060,N_4920,N_3009);
nor U7061 (N_7061,N_2614,N_4915);
or U7062 (N_7062,N_3616,N_4599);
and U7063 (N_7063,N_2579,N_3579);
or U7064 (N_7064,N_2921,N_2876);
nor U7065 (N_7065,N_4220,N_3422);
and U7066 (N_7066,N_2761,N_4769);
and U7067 (N_7067,N_2596,N_4939);
nor U7068 (N_7068,N_2767,N_4598);
nor U7069 (N_7069,N_3743,N_4207);
nor U7070 (N_7070,N_4491,N_3308);
nor U7071 (N_7071,N_3194,N_3373);
nand U7072 (N_7072,N_3974,N_3771);
and U7073 (N_7073,N_4562,N_2720);
xor U7074 (N_7074,N_4272,N_2858);
or U7075 (N_7075,N_3614,N_2899);
nor U7076 (N_7076,N_3434,N_2510);
nor U7077 (N_7077,N_4182,N_3016);
xnor U7078 (N_7078,N_3140,N_4829);
nor U7079 (N_7079,N_3450,N_4712);
xor U7080 (N_7080,N_4982,N_4181);
and U7081 (N_7081,N_3592,N_3006);
nor U7082 (N_7082,N_2596,N_4532);
nor U7083 (N_7083,N_3670,N_2621);
or U7084 (N_7084,N_4903,N_4281);
or U7085 (N_7085,N_3816,N_2618);
nand U7086 (N_7086,N_3131,N_4437);
xnor U7087 (N_7087,N_2866,N_4202);
nor U7088 (N_7088,N_3480,N_2834);
or U7089 (N_7089,N_3450,N_4843);
nand U7090 (N_7090,N_4058,N_2792);
and U7091 (N_7091,N_3937,N_3157);
xnor U7092 (N_7092,N_3777,N_4136);
nand U7093 (N_7093,N_3967,N_3105);
and U7094 (N_7094,N_2873,N_2524);
xor U7095 (N_7095,N_4338,N_4111);
nand U7096 (N_7096,N_4386,N_4088);
nor U7097 (N_7097,N_4385,N_3045);
or U7098 (N_7098,N_3146,N_3224);
nor U7099 (N_7099,N_4558,N_3584);
or U7100 (N_7100,N_2919,N_2567);
nand U7101 (N_7101,N_4066,N_2707);
nand U7102 (N_7102,N_4467,N_4191);
xnor U7103 (N_7103,N_2677,N_4118);
nand U7104 (N_7104,N_3473,N_2813);
xnor U7105 (N_7105,N_3567,N_4781);
nand U7106 (N_7106,N_2993,N_3695);
nor U7107 (N_7107,N_4902,N_2775);
or U7108 (N_7108,N_2956,N_2814);
or U7109 (N_7109,N_4173,N_3049);
nand U7110 (N_7110,N_4626,N_4273);
and U7111 (N_7111,N_2880,N_2676);
nand U7112 (N_7112,N_4555,N_2693);
nand U7113 (N_7113,N_4431,N_3726);
xor U7114 (N_7114,N_4806,N_2825);
xor U7115 (N_7115,N_2907,N_2868);
nand U7116 (N_7116,N_2885,N_2767);
or U7117 (N_7117,N_4287,N_3923);
nor U7118 (N_7118,N_3221,N_3306);
or U7119 (N_7119,N_4454,N_4642);
nor U7120 (N_7120,N_2973,N_3244);
and U7121 (N_7121,N_2771,N_2514);
xor U7122 (N_7122,N_4993,N_4992);
nor U7123 (N_7123,N_4777,N_4811);
or U7124 (N_7124,N_3987,N_2843);
xnor U7125 (N_7125,N_4962,N_3698);
or U7126 (N_7126,N_3763,N_3507);
and U7127 (N_7127,N_4679,N_4502);
xnor U7128 (N_7128,N_3667,N_3290);
nor U7129 (N_7129,N_4516,N_4843);
nor U7130 (N_7130,N_4147,N_4855);
and U7131 (N_7131,N_2798,N_4019);
xnor U7132 (N_7132,N_4043,N_4254);
or U7133 (N_7133,N_3655,N_4508);
or U7134 (N_7134,N_4907,N_3604);
nand U7135 (N_7135,N_3279,N_3947);
or U7136 (N_7136,N_2803,N_4288);
or U7137 (N_7137,N_4168,N_2967);
nor U7138 (N_7138,N_3006,N_2741);
nor U7139 (N_7139,N_4058,N_3285);
xnor U7140 (N_7140,N_4643,N_4239);
or U7141 (N_7141,N_4969,N_4276);
xnor U7142 (N_7142,N_4637,N_4620);
nand U7143 (N_7143,N_2617,N_2965);
xnor U7144 (N_7144,N_3946,N_3998);
xnor U7145 (N_7145,N_4574,N_3370);
nand U7146 (N_7146,N_4079,N_3345);
nand U7147 (N_7147,N_3894,N_2708);
nor U7148 (N_7148,N_3000,N_3270);
nand U7149 (N_7149,N_2631,N_4364);
and U7150 (N_7150,N_4557,N_4271);
and U7151 (N_7151,N_3759,N_3559);
nand U7152 (N_7152,N_3084,N_4463);
nand U7153 (N_7153,N_4134,N_4800);
and U7154 (N_7154,N_3411,N_3196);
nand U7155 (N_7155,N_2536,N_4927);
or U7156 (N_7156,N_2796,N_4547);
xnor U7157 (N_7157,N_3580,N_3785);
or U7158 (N_7158,N_3563,N_4704);
nor U7159 (N_7159,N_4920,N_2537);
nor U7160 (N_7160,N_3621,N_3446);
and U7161 (N_7161,N_4391,N_3277);
nand U7162 (N_7162,N_4454,N_3125);
nor U7163 (N_7163,N_3814,N_4126);
nor U7164 (N_7164,N_2722,N_3071);
xnor U7165 (N_7165,N_4180,N_2511);
or U7166 (N_7166,N_4144,N_3146);
or U7167 (N_7167,N_3888,N_3576);
and U7168 (N_7168,N_3334,N_3318);
nor U7169 (N_7169,N_3442,N_4794);
and U7170 (N_7170,N_3984,N_3280);
nand U7171 (N_7171,N_3575,N_4223);
nor U7172 (N_7172,N_4327,N_2608);
or U7173 (N_7173,N_3366,N_2861);
xor U7174 (N_7174,N_3342,N_3402);
nor U7175 (N_7175,N_3685,N_4409);
nand U7176 (N_7176,N_2995,N_3150);
or U7177 (N_7177,N_4231,N_4926);
nor U7178 (N_7178,N_2756,N_3830);
and U7179 (N_7179,N_4269,N_4973);
or U7180 (N_7180,N_3359,N_4515);
or U7181 (N_7181,N_4227,N_2603);
nand U7182 (N_7182,N_4833,N_3360);
nor U7183 (N_7183,N_3121,N_2658);
xnor U7184 (N_7184,N_2649,N_3741);
or U7185 (N_7185,N_3244,N_3039);
and U7186 (N_7186,N_4258,N_2781);
nand U7187 (N_7187,N_3831,N_4708);
nor U7188 (N_7188,N_3848,N_3054);
or U7189 (N_7189,N_4212,N_4317);
xnor U7190 (N_7190,N_4646,N_2520);
nor U7191 (N_7191,N_4399,N_4402);
nand U7192 (N_7192,N_2840,N_4467);
nand U7193 (N_7193,N_2979,N_4342);
nand U7194 (N_7194,N_4581,N_4333);
nor U7195 (N_7195,N_4714,N_4812);
xnor U7196 (N_7196,N_3328,N_2730);
xnor U7197 (N_7197,N_3672,N_2809);
and U7198 (N_7198,N_3893,N_3014);
xnor U7199 (N_7199,N_4526,N_3692);
nand U7200 (N_7200,N_2635,N_3884);
nand U7201 (N_7201,N_4776,N_4101);
and U7202 (N_7202,N_4917,N_3115);
xor U7203 (N_7203,N_4686,N_4986);
nor U7204 (N_7204,N_3106,N_4810);
or U7205 (N_7205,N_3574,N_3979);
xnor U7206 (N_7206,N_3354,N_3941);
nor U7207 (N_7207,N_4166,N_4332);
nand U7208 (N_7208,N_4613,N_4224);
nor U7209 (N_7209,N_3615,N_4277);
nand U7210 (N_7210,N_2985,N_2737);
xnor U7211 (N_7211,N_3175,N_3824);
nand U7212 (N_7212,N_3578,N_4622);
or U7213 (N_7213,N_4777,N_3480);
nand U7214 (N_7214,N_4992,N_4002);
nor U7215 (N_7215,N_2552,N_2820);
nor U7216 (N_7216,N_2843,N_4860);
nor U7217 (N_7217,N_4015,N_3708);
and U7218 (N_7218,N_4070,N_4322);
nor U7219 (N_7219,N_4227,N_3317);
nand U7220 (N_7220,N_3361,N_2931);
and U7221 (N_7221,N_4622,N_4161);
xnor U7222 (N_7222,N_2802,N_3226);
nand U7223 (N_7223,N_4131,N_4717);
xnor U7224 (N_7224,N_3319,N_3698);
nand U7225 (N_7225,N_3186,N_3665);
nor U7226 (N_7226,N_3831,N_4339);
xor U7227 (N_7227,N_3359,N_3144);
xnor U7228 (N_7228,N_4912,N_3112);
xor U7229 (N_7229,N_3619,N_4949);
xor U7230 (N_7230,N_4352,N_4620);
and U7231 (N_7231,N_4116,N_2971);
and U7232 (N_7232,N_3460,N_3462);
nor U7233 (N_7233,N_4563,N_4741);
or U7234 (N_7234,N_3477,N_4663);
nor U7235 (N_7235,N_4548,N_4023);
or U7236 (N_7236,N_3960,N_3514);
xnor U7237 (N_7237,N_3626,N_4167);
or U7238 (N_7238,N_2799,N_3442);
or U7239 (N_7239,N_4079,N_2934);
nor U7240 (N_7240,N_4446,N_3925);
xnor U7241 (N_7241,N_3235,N_4306);
xnor U7242 (N_7242,N_3357,N_3314);
nand U7243 (N_7243,N_4753,N_3369);
xnor U7244 (N_7244,N_4173,N_2752);
nor U7245 (N_7245,N_3606,N_3633);
or U7246 (N_7246,N_4609,N_3576);
nand U7247 (N_7247,N_4850,N_3894);
nor U7248 (N_7248,N_3301,N_3876);
and U7249 (N_7249,N_3161,N_3339);
nor U7250 (N_7250,N_3782,N_4390);
nand U7251 (N_7251,N_4051,N_2820);
or U7252 (N_7252,N_3874,N_4179);
xor U7253 (N_7253,N_4110,N_4841);
nor U7254 (N_7254,N_2793,N_3597);
xnor U7255 (N_7255,N_4321,N_4835);
or U7256 (N_7256,N_3988,N_3195);
xnor U7257 (N_7257,N_2752,N_3558);
and U7258 (N_7258,N_4812,N_2674);
nor U7259 (N_7259,N_3094,N_4755);
xnor U7260 (N_7260,N_3824,N_3051);
xor U7261 (N_7261,N_3438,N_3432);
and U7262 (N_7262,N_2714,N_3545);
nor U7263 (N_7263,N_3084,N_4160);
nand U7264 (N_7264,N_4094,N_3687);
xnor U7265 (N_7265,N_2852,N_4566);
xor U7266 (N_7266,N_3741,N_3642);
and U7267 (N_7267,N_2778,N_3569);
xor U7268 (N_7268,N_3971,N_4749);
nand U7269 (N_7269,N_4353,N_3109);
nor U7270 (N_7270,N_2977,N_2794);
nand U7271 (N_7271,N_4238,N_3153);
nand U7272 (N_7272,N_2530,N_3672);
nand U7273 (N_7273,N_2906,N_4303);
xor U7274 (N_7274,N_4213,N_2961);
or U7275 (N_7275,N_4112,N_2745);
xnor U7276 (N_7276,N_2626,N_4590);
nand U7277 (N_7277,N_4517,N_3139);
or U7278 (N_7278,N_2990,N_4146);
nor U7279 (N_7279,N_3305,N_4476);
nand U7280 (N_7280,N_3128,N_3462);
nand U7281 (N_7281,N_3294,N_3835);
and U7282 (N_7282,N_4906,N_3945);
nor U7283 (N_7283,N_2633,N_3212);
nor U7284 (N_7284,N_4743,N_4117);
nor U7285 (N_7285,N_4970,N_3254);
or U7286 (N_7286,N_4312,N_3130);
or U7287 (N_7287,N_3338,N_3599);
xor U7288 (N_7288,N_3596,N_3218);
nand U7289 (N_7289,N_4579,N_3918);
nor U7290 (N_7290,N_2878,N_2795);
xor U7291 (N_7291,N_2983,N_3671);
xor U7292 (N_7292,N_2819,N_3873);
and U7293 (N_7293,N_2857,N_3780);
nor U7294 (N_7294,N_4310,N_4596);
xnor U7295 (N_7295,N_3305,N_2977);
or U7296 (N_7296,N_3450,N_3058);
xnor U7297 (N_7297,N_4820,N_4301);
xnor U7298 (N_7298,N_3013,N_3591);
xnor U7299 (N_7299,N_4787,N_3993);
nand U7300 (N_7300,N_3348,N_3679);
nand U7301 (N_7301,N_4496,N_4881);
and U7302 (N_7302,N_2584,N_4609);
xnor U7303 (N_7303,N_3847,N_4738);
or U7304 (N_7304,N_3066,N_3931);
and U7305 (N_7305,N_3636,N_3919);
or U7306 (N_7306,N_2881,N_3943);
xnor U7307 (N_7307,N_4529,N_4548);
nand U7308 (N_7308,N_3646,N_4130);
or U7309 (N_7309,N_3327,N_3684);
or U7310 (N_7310,N_2867,N_4173);
nor U7311 (N_7311,N_4031,N_2708);
and U7312 (N_7312,N_4496,N_4806);
and U7313 (N_7313,N_4383,N_2520);
xnor U7314 (N_7314,N_4970,N_4490);
nand U7315 (N_7315,N_4415,N_3279);
nand U7316 (N_7316,N_3389,N_4570);
nor U7317 (N_7317,N_3905,N_3426);
nor U7318 (N_7318,N_3634,N_3658);
or U7319 (N_7319,N_2658,N_3032);
nor U7320 (N_7320,N_2771,N_3399);
xor U7321 (N_7321,N_2778,N_4943);
nor U7322 (N_7322,N_3093,N_2578);
nand U7323 (N_7323,N_4638,N_2879);
or U7324 (N_7324,N_3992,N_4153);
nor U7325 (N_7325,N_4289,N_4632);
nand U7326 (N_7326,N_4047,N_4717);
and U7327 (N_7327,N_4754,N_3203);
or U7328 (N_7328,N_3463,N_4673);
xnor U7329 (N_7329,N_4864,N_4170);
or U7330 (N_7330,N_3287,N_4823);
xnor U7331 (N_7331,N_3105,N_3740);
or U7332 (N_7332,N_2670,N_4955);
nand U7333 (N_7333,N_3496,N_4198);
nor U7334 (N_7334,N_2968,N_3136);
or U7335 (N_7335,N_4791,N_2980);
and U7336 (N_7336,N_4959,N_3688);
xor U7337 (N_7337,N_4623,N_3586);
nor U7338 (N_7338,N_3382,N_2660);
nand U7339 (N_7339,N_2667,N_3509);
nand U7340 (N_7340,N_3868,N_4139);
or U7341 (N_7341,N_4292,N_4842);
or U7342 (N_7342,N_2722,N_2731);
nor U7343 (N_7343,N_4067,N_3460);
xor U7344 (N_7344,N_2804,N_3134);
nor U7345 (N_7345,N_3218,N_2717);
nor U7346 (N_7346,N_4997,N_3705);
nand U7347 (N_7347,N_2910,N_3657);
xnor U7348 (N_7348,N_4928,N_3871);
nor U7349 (N_7349,N_4044,N_3339);
nor U7350 (N_7350,N_3148,N_4714);
nor U7351 (N_7351,N_2572,N_3994);
or U7352 (N_7352,N_3549,N_3362);
and U7353 (N_7353,N_4820,N_4780);
nor U7354 (N_7354,N_3134,N_4223);
or U7355 (N_7355,N_2859,N_3853);
nand U7356 (N_7356,N_4369,N_3289);
nand U7357 (N_7357,N_4946,N_2647);
or U7358 (N_7358,N_2847,N_3218);
xnor U7359 (N_7359,N_3375,N_4464);
or U7360 (N_7360,N_3491,N_3291);
nand U7361 (N_7361,N_3581,N_3199);
nand U7362 (N_7362,N_2742,N_2919);
nor U7363 (N_7363,N_4006,N_2874);
xnor U7364 (N_7364,N_4374,N_4981);
and U7365 (N_7365,N_3681,N_3378);
or U7366 (N_7366,N_4811,N_3514);
xor U7367 (N_7367,N_3042,N_4122);
or U7368 (N_7368,N_4361,N_4570);
xor U7369 (N_7369,N_3591,N_4252);
xnor U7370 (N_7370,N_3731,N_4847);
xnor U7371 (N_7371,N_3325,N_4795);
nand U7372 (N_7372,N_4036,N_4355);
nor U7373 (N_7373,N_4182,N_3702);
and U7374 (N_7374,N_4773,N_3622);
nand U7375 (N_7375,N_4659,N_4857);
or U7376 (N_7376,N_3605,N_4308);
and U7377 (N_7377,N_3504,N_2762);
xnor U7378 (N_7378,N_3463,N_3237);
nor U7379 (N_7379,N_2642,N_3932);
nor U7380 (N_7380,N_2626,N_4431);
or U7381 (N_7381,N_4504,N_4713);
nor U7382 (N_7382,N_4313,N_4538);
xor U7383 (N_7383,N_4733,N_3682);
and U7384 (N_7384,N_3172,N_4793);
nor U7385 (N_7385,N_4401,N_4753);
nand U7386 (N_7386,N_2740,N_2832);
nor U7387 (N_7387,N_3669,N_2546);
nor U7388 (N_7388,N_2919,N_3033);
xor U7389 (N_7389,N_2811,N_2954);
or U7390 (N_7390,N_2775,N_4517);
and U7391 (N_7391,N_3812,N_4293);
xnor U7392 (N_7392,N_2713,N_2856);
nand U7393 (N_7393,N_3144,N_2713);
nand U7394 (N_7394,N_3153,N_2501);
nor U7395 (N_7395,N_2707,N_3236);
and U7396 (N_7396,N_2679,N_3369);
nor U7397 (N_7397,N_3094,N_3555);
nor U7398 (N_7398,N_3060,N_4448);
nor U7399 (N_7399,N_3067,N_4849);
and U7400 (N_7400,N_3833,N_3002);
nor U7401 (N_7401,N_3882,N_2878);
nand U7402 (N_7402,N_2850,N_3914);
nor U7403 (N_7403,N_4137,N_3507);
or U7404 (N_7404,N_4362,N_3791);
nor U7405 (N_7405,N_4425,N_3394);
nand U7406 (N_7406,N_2930,N_2697);
nand U7407 (N_7407,N_3908,N_4226);
nor U7408 (N_7408,N_4509,N_4120);
and U7409 (N_7409,N_4310,N_3867);
and U7410 (N_7410,N_3092,N_2712);
nand U7411 (N_7411,N_3232,N_3034);
nor U7412 (N_7412,N_4001,N_2771);
or U7413 (N_7413,N_4647,N_3833);
nand U7414 (N_7414,N_4682,N_3957);
or U7415 (N_7415,N_3989,N_3933);
nand U7416 (N_7416,N_4193,N_3513);
nand U7417 (N_7417,N_4060,N_4764);
xor U7418 (N_7418,N_4713,N_4478);
xor U7419 (N_7419,N_4455,N_4356);
xor U7420 (N_7420,N_3398,N_4936);
xnor U7421 (N_7421,N_4916,N_4407);
and U7422 (N_7422,N_4186,N_3051);
xor U7423 (N_7423,N_3777,N_3369);
xor U7424 (N_7424,N_4889,N_4094);
and U7425 (N_7425,N_2796,N_2634);
nor U7426 (N_7426,N_2749,N_4547);
or U7427 (N_7427,N_3895,N_2526);
and U7428 (N_7428,N_3715,N_3473);
xnor U7429 (N_7429,N_3467,N_4971);
and U7430 (N_7430,N_3404,N_2787);
nand U7431 (N_7431,N_3383,N_3977);
xnor U7432 (N_7432,N_3659,N_2972);
xor U7433 (N_7433,N_4599,N_2996);
and U7434 (N_7434,N_3818,N_4498);
and U7435 (N_7435,N_4222,N_3682);
xor U7436 (N_7436,N_3265,N_2511);
xor U7437 (N_7437,N_4848,N_3925);
nor U7438 (N_7438,N_4318,N_4345);
nor U7439 (N_7439,N_4612,N_2760);
xor U7440 (N_7440,N_4921,N_3105);
nand U7441 (N_7441,N_4811,N_2981);
nor U7442 (N_7442,N_4416,N_2674);
nand U7443 (N_7443,N_3032,N_2995);
nand U7444 (N_7444,N_4705,N_3031);
nand U7445 (N_7445,N_3741,N_4803);
nor U7446 (N_7446,N_2705,N_4201);
nor U7447 (N_7447,N_3342,N_4535);
nand U7448 (N_7448,N_3251,N_4021);
nor U7449 (N_7449,N_4623,N_4923);
nand U7450 (N_7450,N_3309,N_3346);
nor U7451 (N_7451,N_2753,N_3953);
and U7452 (N_7452,N_4838,N_4700);
or U7453 (N_7453,N_3876,N_2970);
nor U7454 (N_7454,N_3837,N_4354);
or U7455 (N_7455,N_3896,N_3446);
or U7456 (N_7456,N_4136,N_4952);
nor U7457 (N_7457,N_3461,N_4625);
or U7458 (N_7458,N_2686,N_4088);
and U7459 (N_7459,N_3583,N_3172);
and U7460 (N_7460,N_3309,N_3959);
xor U7461 (N_7461,N_2730,N_3144);
and U7462 (N_7462,N_2927,N_4456);
and U7463 (N_7463,N_4666,N_2818);
xnor U7464 (N_7464,N_4157,N_3028);
nand U7465 (N_7465,N_3740,N_2632);
nor U7466 (N_7466,N_3208,N_4959);
xnor U7467 (N_7467,N_3974,N_4387);
or U7468 (N_7468,N_3080,N_2578);
and U7469 (N_7469,N_3817,N_3969);
xnor U7470 (N_7470,N_3736,N_4493);
and U7471 (N_7471,N_4835,N_4481);
nor U7472 (N_7472,N_4108,N_3492);
nand U7473 (N_7473,N_4750,N_2654);
xor U7474 (N_7474,N_4533,N_4864);
xor U7475 (N_7475,N_2731,N_3642);
xor U7476 (N_7476,N_4343,N_2785);
nand U7477 (N_7477,N_2796,N_2719);
or U7478 (N_7478,N_3358,N_4250);
or U7479 (N_7479,N_2945,N_2758);
nand U7480 (N_7480,N_3381,N_2579);
nor U7481 (N_7481,N_3886,N_2565);
nand U7482 (N_7482,N_3265,N_4362);
and U7483 (N_7483,N_3214,N_2798);
nor U7484 (N_7484,N_4303,N_4147);
nand U7485 (N_7485,N_2622,N_2907);
or U7486 (N_7486,N_4076,N_4668);
or U7487 (N_7487,N_4372,N_3009);
and U7488 (N_7488,N_3811,N_4135);
and U7489 (N_7489,N_4029,N_3897);
xnor U7490 (N_7490,N_3106,N_3280);
nor U7491 (N_7491,N_4509,N_4855);
xor U7492 (N_7492,N_4720,N_3947);
nor U7493 (N_7493,N_4541,N_4414);
nand U7494 (N_7494,N_3489,N_4315);
and U7495 (N_7495,N_4397,N_4378);
nand U7496 (N_7496,N_4248,N_3025);
nand U7497 (N_7497,N_3716,N_3482);
or U7498 (N_7498,N_3831,N_4181);
or U7499 (N_7499,N_3147,N_3482);
nor U7500 (N_7500,N_6940,N_6678);
or U7501 (N_7501,N_7000,N_6786);
nor U7502 (N_7502,N_6714,N_5919);
xor U7503 (N_7503,N_6433,N_6145);
nand U7504 (N_7504,N_5416,N_6115);
and U7505 (N_7505,N_5210,N_6595);
nor U7506 (N_7506,N_6090,N_6460);
nor U7507 (N_7507,N_6455,N_5658);
nand U7508 (N_7508,N_7035,N_6651);
or U7509 (N_7509,N_7498,N_7420);
and U7510 (N_7510,N_6841,N_5630);
xor U7511 (N_7511,N_6180,N_7412);
nand U7512 (N_7512,N_6753,N_6482);
nor U7513 (N_7513,N_6472,N_6950);
nand U7514 (N_7514,N_6134,N_7195);
nor U7515 (N_7515,N_6930,N_5415);
and U7516 (N_7516,N_5321,N_5284);
xor U7517 (N_7517,N_7271,N_5510);
nor U7518 (N_7518,N_5074,N_6812);
nand U7519 (N_7519,N_6619,N_6633);
xor U7520 (N_7520,N_6888,N_6994);
or U7521 (N_7521,N_5958,N_6889);
nand U7522 (N_7522,N_5078,N_7041);
or U7523 (N_7523,N_5069,N_5299);
xnor U7524 (N_7524,N_5914,N_5361);
nor U7525 (N_7525,N_6341,N_5347);
and U7526 (N_7526,N_7369,N_6388);
or U7527 (N_7527,N_6095,N_6112);
or U7528 (N_7528,N_6993,N_6294);
and U7529 (N_7529,N_5500,N_6347);
and U7530 (N_7530,N_6526,N_6811);
nand U7531 (N_7531,N_7255,N_6567);
nand U7532 (N_7532,N_7269,N_5833);
xnor U7533 (N_7533,N_7134,N_5103);
xor U7534 (N_7534,N_5834,N_6211);
and U7535 (N_7535,N_6334,N_6412);
xor U7536 (N_7536,N_6259,N_7266);
nor U7537 (N_7537,N_6017,N_6673);
nand U7538 (N_7538,N_5434,N_7380);
xor U7539 (N_7539,N_5750,N_5997);
nand U7540 (N_7540,N_7361,N_6260);
xor U7541 (N_7541,N_7175,N_5012);
xor U7542 (N_7542,N_6667,N_5717);
and U7543 (N_7543,N_7217,N_6537);
nor U7544 (N_7544,N_6337,N_5785);
xor U7545 (N_7545,N_6688,N_7357);
or U7546 (N_7546,N_5720,N_6013);
or U7547 (N_7547,N_7497,N_5405);
nor U7548 (N_7548,N_7477,N_7478);
nand U7549 (N_7549,N_6147,N_7423);
and U7550 (N_7550,N_5723,N_7199);
or U7551 (N_7551,N_5026,N_5377);
xnor U7552 (N_7552,N_6458,N_5033);
nor U7553 (N_7553,N_7260,N_6784);
and U7554 (N_7554,N_6317,N_7076);
and U7555 (N_7555,N_6061,N_7065);
or U7556 (N_7556,N_5503,N_7379);
or U7557 (N_7557,N_5089,N_6133);
or U7558 (N_7558,N_5136,N_5946);
nor U7559 (N_7559,N_5056,N_5135);
and U7560 (N_7560,N_6923,N_7499);
nor U7561 (N_7561,N_5517,N_6252);
nor U7562 (N_7562,N_5961,N_6826);
and U7563 (N_7563,N_5877,N_6542);
and U7564 (N_7564,N_6071,N_5665);
xor U7565 (N_7565,N_7452,N_5110);
nor U7566 (N_7566,N_5054,N_6282);
and U7567 (N_7567,N_7064,N_6223);
xor U7568 (N_7568,N_5220,N_6383);
nand U7569 (N_7569,N_6646,N_6301);
nand U7570 (N_7570,N_7228,N_5280);
xnor U7571 (N_7571,N_7216,N_6903);
and U7572 (N_7572,N_5037,N_6033);
or U7573 (N_7573,N_6418,N_5697);
xor U7574 (N_7574,N_5085,N_6516);
nand U7575 (N_7575,N_6424,N_6397);
nor U7576 (N_7576,N_5302,N_5443);
nand U7577 (N_7577,N_7408,N_5094);
xor U7578 (N_7578,N_6363,N_6591);
xor U7579 (N_7579,N_7012,N_5937);
nor U7580 (N_7580,N_6517,N_5605);
nor U7581 (N_7581,N_5813,N_6988);
and U7582 (N_7582,N_5974,N_6932);
or U7583 (N_7583,N_7395,N_5516);
xnor U7584 (N_7584,N_6298,N_6519);
or U7585 (N_7585,N_5985,N_5562);
nor U7586 (N_7586,N_5841,N_7085);
xor U7587 (N_7587,N_6879,N_5338);
or U7588 (N_7588,N_6356,N_5366);
nand U7589 (N_7589,N_5447,N_7278);
nand U7590 (N_7590,N_5451,N_6401);
and U7591 (N_7591,N_6375,N_6783);
xnor U7592 (N_7592,N_5777,N_7356);
and U7593 (N_7593,N_6419,N_5050);
nand U7594 (N_7594,N_5906,N_5827);
or U7595 (N_7595,N_6330,N_6638);
nor U7596 (N_7596,N_6159,N_5905);
or U7597 (N_7597,N_6428,N_7120);
xor U7598 (N_7598,N_6348,N_6410);
and U7599 (N_7599,N_5943,N_6142);
and U7600 (N_7600,N_7407,N_5980);
and U7601 (N_7601,N_5794,N_5725);
nor U7602 (N_7602,N_7440,N_7323);
nor U7603 (N_7603,N_6055,N_6637);
nor U7604 (N_7604,N_6524,N_6630);
nand U7605 (N_7605,N_5560,N_7386);
xnor U7606 (N_7606,N_6871,N_5496);
nor U7607 (N_7607,N_6528,N_5076);
nand U7608 (N_7608,N_7224,N_5628);
or U7609 (N_7609,N_6631,N_7203);
nor U7610 (N_7610,N_6878,N_6427);
and U7611 (N_7611,N_6649,N_6832);
or U7612 (N_7612,N_6978,N_6436);
or U7613 (N_7613,N_5741,N_6350);
nor U7614 (N_7614,N_6746,N_6407);
or U7615 (N_7615,N_5912,N_7054);
xor U7616 (N_7616,N_6729,N_5365);
nor U7617 (N_7617,N_7005,N_5409);
nor U7618 (N_7618,N_6741,N_6261);
and U7619 (N_7619,N_5576,N_5801);
nand U7620 (N_7620,N_6722,N_5079);
nor U7621 (N_7621,N_5825,N_7157);
nand U7622 (N_7622,N_5820,N_5335);
or U7623 (N_7623,N_5013,N_6882);
nand U7624 (N_7624,N_7250,N_6610);
nand U7625 (N_7625,N_5549,N_6942);
and U7626 (N_7626,N_7354,N_7337);
nor U7627 (N_7627,N_5818,N_5786);
xor U7628 (N_7628,N_5298,N_6668);
nand U7629 (N_7629,N_5408,N_6676);
nand U7630 (N_7630,N_6721,N_5792);
xor U7631 (N_7631,N_5838,N_5346);
nor U7632 (N_7632,N_7114,N_5533);
or U7633 (N_7633,N_7472,N_5350);
xnor U7634 (N_7634,N_5973,N_6331);
xor U7635 (N_7635,N_6558,N_5198);
and U7636 (N_7636,N_7342,N_5247);
xnor U7637 (N_7637,N_7291,N_6273);
xor U7638 (N_7638,N_5970,N_6205);
nor U7639 (N_7639,N_6484,N_7460);
and U7640 (N_7640,N_6225,N_5543);
xnor U7641 (N_7641,N_6338,N_5940);
nand U7642 (N_7642,N_5169,N_5018);
xnor U7643 (N_7643,N_5459,N_7463);
xnor U7644 (N_7644,N_7014,N_6265);
or U7645 (N_7645,N_5354,N_7074);
nand U7646 (N_7646,N_7394,N_5715);
and U7647 (N_7647,N_6662,N_6488);
nor U7648 (N_7648,N_6439,N_5622);
xnor U7649 (N_7649,N_5633,N_6025);
nor U7650 (N_7650,N_7042,N_7002);
and U7651 (N_7651,N_5646,N_5647);
xor U7652 (N_7652,N_5716,N_6696);
and U7653 (N_7653,N_7070,N_6322);
nand U7654 (N_7654,N_6764,N_6659);
or U7655 (N_7655,N_5222,N_5066);
or U7656 (N_7656,N_5507,N_6757);
nand U7657 (N_7657,N_5132,N_7084);
xnor U7658 (N_7658,N_5735,N_5472);
nand U7659 (N_7659,N_7450,N_5291);
or U7660 (N_7660,N_7075,N_6078);
or U7661 (N_7661,N_6563,N_5602);
nor U7662 (N_7662,N_5143,N_6155);
or U7663 (N_7663,N_6157,N_5843);
nor U7664 (N_7664,N_6733,N_7221);
xnor U7665 (N_7665,N_6110,N_6480);
and U7666 (N_7666,N_5608,N_5372);
or U7667 (N_7667,N_7311,N_7262);
xor U7668 (N_7668,N_6283,N_5036);
nand U7669 (N_7669,N_7371,N_6052);
nand U7670 (N_7670,N_6303,N_6049);
xor U7671 (N_7671,N_5855,N_5326);
or U7672 (N_7672,N_7147,N_7392);
nor U7673 (N_7673,N_6496,N_5854);
nand U7674 (N_7674,N_5096,N_6343);
nand U7675 (N_7675,N_7404,N_7229);
or U7676 (N_7676,N_6816,N_7415);
nand U7677 (N_7677,N_5739,N_7086);
xnor U7678 (N_7678,N_5755,N_5252);
and U7679 (N_7679,N_7048,N_7272);
nand U7680 (N_7680,N_7313,N_6309);
xor U7681 (N_7681,N_7170,N_6856);
nand U7682 (N_7682,N_6704,N_7491);
or U7683 (N_7683,N_7326,N_5520);
and U7684 (N_7684,N_6750,N_6953);
xnor U7685 (N_7685,N_6467,N_5241);
xnor U7686 (N_7686,N_5484,N_5534);
xnor U7687 (N_7687,N_5362,N_6596);
and U7688 (N_7688,N_7190,N_5891);
xnor U7689 (N_7689,N_6626,N_6902);
or U7690 (N_7690,N_7124,N_5556);
xor U7691 (N_7691,N_5042,N_7487);
and U7692 (N_7692,N_5444,N_5677);
and U7693 (N_7693,N_5676,N_7368);
xor U7694 (N_7694,N_5882,N_6057);
or U7695 (N_7695,N_7339,N_7061);
nor U7696 (N_7696,N_5221,N_6996);
and U7697 (N_7697,N_7307,N_7052);
xor U7698 (N_7698,N_5123,N_6779);
and U7699 (N_7699,N_5816,N_6569);
xnor U7700 (N_7700,N_5315,N_6904);
or U7701 (N_7701,N_5866,N_7430);
xnor U7702 (N_7702,N_5903,N_6872);
nand U7703 (N_7703,N_7492,N_6192);
nand U7704 (N_7704,N_5967,N_7039);
nor U7705 (N_7705,N_5823,N_6380);
xor U7706 (N_7706,N_7340,N_5144);
or U7707 (N_7707,N_6821,N_7429);
or U7708 (N_7708,N_6046,N_5743);
nand U7709 (N_7709,N_5863,N_7155);
and U7710 (N_7710,N_6394,N_5343);
or U7711 (N_7711,N_6937,N_7287);
xnor U7712 (N_7712,N_6587,N_5203);
and U7713 (N_7713,N_6617,N_6128);
nand U7714 (N_7714,N_7471,N_7367);
nor U7715 (N_7715,N_6374,N_6794);
and U7716 (N_7716,N_5711,N_5617);
nand U7717 (N_7717,N_6890,N_6756);
nor U7718 (N_7718,N_5563,N_6158);
and U7719 (N_7719,N_5407,N_6098);
nor U7720 (N_7720,N_5614,N_6847);
nor U7721 (N_7721,N_5043,N_7439);
or U7722 (N_7722,N_7008,N_6060);
or U7723 (N_7723,N_7037,N_6429);
and U7724 (N_7724,N_5975,N_7372);
nor U7725 (N_7725,N_6984,N_6468);
xnor U7726 (N_7726,N_5933,N_6612);
nand U7727 (N_7727,N_5681,N_5703);
or U7728 (N_7728,N_6384,N_5462);
nand U7729 (N_7729,N_6747,N_6765);
nor U7730 (N_7730,N_6464,N_6728);
and U7731 (N_7731,N_7459,N_5045);
nor U7732 (N_7732,N_7210,N_5800);
nor U7733 (N_7733,N_5088,N_7118);
nand U7734 (N_7734,N_5190,N_7001);
and U7735 (N_7735,N_5402,N_5944);
nand U7736 (N_7736,N_5511,N_6402);
nor U7737 (N_7737,N_6613,N_5293);
nor U7738 (N_7738,N_6062,N_7265);
or U7739 (N_7739,N_5464,N_6312);
and U7740 (N_7740,N_7159,N_6555);
nor U7741 (N_7741,N_7276,N_6578);
or U7742 (N_7742,N_6197,N_5615);
and U7743 (N_7743,N_5260,N_6672);
and U7744 (N_7744,N_6691,N_5766);
nand U7745 (N_7745,N_5683,N_6475);
xor U7746 (N_7746,N_6190,N_7348);
nand U7747 (N_7747,N_6014,N_5465);
and U7748 (N_7748,N_6236,N_5945);
xor U7749 (N_7749,N_7149,N_6852);
nand U7750 (N_7750,N_7239,N_7322);
xnor U7751 (N_7751,N_7243,N_5979);
nor U7752 (N_7752,N_5494,N_5957);
and U7753 (N_7753,N_5240,N_6835);
xor U7754 (N_7754,N_7174,N_7451);
and U7755 (N_7755,N_6342,N_7316);
nand U7756 (N_7756,N_5784,N_6103);
xor U7757 (N_7757,N_7066,N_5490);
nor U7758 (N_7758,N_6502,N_7122);
xor U7759 (N_7759,N_5585,N_5861);
nand U7760 (N_7760,N_6102,N_7106);
or U7761 (N_7761,N_7033,N_5577);
or U7762 (N_7762,N_5911,N_6615);
xnor U7763 (N_7763,N_6124,N_7082);
nor U7764 (N_7764,N_5883,N_6800);
nand U7765 (N_7765,N_6024,N_6562);
and U7766 (N_7766,N_7081,N_6997);
nor U7767 (N_7767,N_6719,N_6680);
nor U7768 (N_7768,N_6725,N_6803);
xor U7769 (N_7769,N_5003,N_7441);
nand U7770 (N_7770,N_6226,N_6834);
nor U7771 (N_7771,N_5782,N_7484);
or U7772 (N_7772,N_7464,N_6361);
nor U7773 (N_7773,N_7044,N_5173);
nor U7774 (N_7774,N_6791,N_5776);
nand U7775 (N_7775,N_6830,N_6952);
and U7776 (N_7776,N_5899,N_5192);
nor U7777 (N_7777,N_7290,N_5994);
or U7778 (N_7778,N_6644,N_6174);
and U7779 (N_7779,N_7251,N_5704);
or U7780 (N_7780,N_5215,N_6987);
xnor U7781 (N_7781,N_5020,N_6804);
or U7782 (N_7782,N_7140,N_7335);
xnor U7783 (N_7783,N_5783,N_6168);
and U7784 (N_7784,N_5699,N_7467);
or U7785 (N_7785,N_6699,N_5673);
and U7786 (N_7786,N_5461,N_5938);
nand U7787 (N_7787,N_7456,N_6598);
and U7788 (N_7788,N_5152,N_5236);
or U7789 (N_7789,N_5864,N_5381);
nand U7790 (N_7790,N_6951,N_5038);
or U7791 (N_7791,N_5852,N_6810);
nand U7792 (N_7792,N_7179,N_5039);
xor U7793 (N_7793,N_5186,N_5194);
and U7794 (N_7794,N_6556,N_6495);
nand U7795 (N_7795,N_6525,N_5672);
xnor U7796 (N_7796,N_5448,N_6479);
and U7797 (N_7797,N_5521,N_5445);
nor U7798 (N_7798,N_5356,N_6059);
nor U7799 (N_7799,N_5106,N_5319);
or U7800 (N_7800,N_5401,N_5330);
and U7801 (N_7801,N_5080,N_6588);
xnor U7802 (N_7802,N_5223,N_5047);
or U7803 (N_7803,N_5548,N_5529);
nor U7804 (N_7804,N_6200,N_5273);
and U7805 (N_7805,N_7454,N_5688);
nand U7806 (N_7806,N_5770,N_5803);
nand U7807 (N_7807,N_7355,N_5292);
xor U7808 (N_7808,N_5340,N_5865);
xnor U7809 (N_7809,N_5331,N_5489);
and U7810 (N_7810,N_5467,N_5892);
and U7811 (N_7811,N_5027,N_7034);
or U7812 (N_7812,N_5508,N_6916);
nand U7813 (N_7813,N_6539,N_7049);
nor U7814 (N_7814,N_6070,N_5468);
nor U7815 (N_7815,N_7150,N_6447);
nor U7816 (N_7816,N_7030,N_5706);
nand U7817 (N_7817,N_5540,N_6970);
nand U7818 (N_7818,N_6353,N_6827);
nand U7819 (N_7819,N_5607,N_6685);
nand U7820 (N_7820,N_5601,N_6144);
and U7821 (N_7821,N_5010,N_6789);
or U7822 (N_7822,N_6431,N_6831);
or U7823 (N_7823,N_5286,N_5239);
xor U7824 (N_7824,N_6692,N_7448);
and U7825 (N_7825,N_7209,N_6257);
nor U7826 (N_7826,N_5493,N_5421);
nor U7827 (N_7827,N_6445,N_6976);
or U7828 (N_7828,N_5460,N_6828);
and U7829 (N_7829,N_7067,N_6648);
nor U7830 (N_7830,N_7309,N_5237);
or U7831 (N_7831,N_5126,N_7164);
nand U7832 (N_7832,N_7489,N_7235);
nor U7833 (N_7833,N_7344,N_7305);
xnor U7834 (N_7834,N_6677,N_6026);
xnor U7835 (N_7835,N_5138,N_7178);
or U7836 (N_7836,N_7100,N_5684);
xor U7837 (N_7837,N_5624,N_6481);
nand U7838 (N_7838,N_5971,N_5998);
nor U7839 (N_7839,N_6231,N_5413);
nor U7840 (N_7840,N_5713,N_7088);
nor U7841 (N_7841,N_6998,N_7453);
xnor U7842 (N_7842,N_5774,N_6371);
xor U7843 (N_7843,N_6915,N_5141);
nand U7844 (N_7844,N_6358,N_6173);
and U7845 (N_7845,N_6570,N_6576);
xnor U7846 (N_7846,N_6408,N_5650);
nor U7847 (N_7847,N_6802,N_5155);
xor U7848 (N_7848,N_5364,N_5748);
nand U7849 (N_7849,N_5555,N_5707);
or U7850 (N_7850,N_6221,N_7176);
xor U7851 (N_7851,N_5234,N_6286);
nand U7852 (N_7852,N_5118,N_7314);
nand U7853 (N_7853,N_5368,N_5049);
or U7854 (N_7854,N_6671,N_5426);
nor U7855 (N_7855,N_5456,N_5011);
xnor U7856 (N_7856,N_6565,N_7197);
nor U7857 (N_7857,N_6921,N_5644);
or U7858 (N_7858,N_5370,N_7447);
or U7859 (N_7859,N_6561,N_5154);
nor U7860 (N_7860,N_5246,N_6191);
xor U7861 (N_7861,N_5499,N_6087);
and U7862 (N_7862,N_7069,N_7194);
or U7863 (N_7863,N_5875,N_6302);
xor U7864 (N_7864,N_6601,N_6875);
or U7865 (N_7865,N_6707,N_7156);
xor U7866 (N_7866,N_5856,N_5351);
nor U7867 (N_7867,N_6584,N_5317);
nor U7868 (N_7868,N_5098,N_5634);
nand U7869 (N_7869,N_5400,N_7173);
nor U7870 (N_7870,N_5603,N_7053);
nor U7871 (N_7871,N_5272,N_6602);
xnor U7872 (N_7872,N_7162,N_6774);
or U7873 (N_7873,N_7377,N_5469);
nor U7874 (N_7874,N_6136,N_5251);
xor U7875 (N_7875,N_6378,N_5059);
or U7876 (N_7876,N_6417,N_7360);
xor U7877 (N_7877,N_5081,N_6104);
or U7878 (N_7878,N_7101,N_6344);
and U7879 (N_7879,N_5373,N_6179);
nor U7880 (N_7880,N_5787,N_7027);
nor U7881 (N_7881,N_6399,N_7144);
and U7882 (N_7882,N_5289,N_6256);
xor U7883 (N_7883,N_7189,N_7182);
nand U7884 (N_7884,N_5120,N_7324);
xor U7885 (N_7885,N_5454,N_5918);
or U7886 (N_7886,N_6980,N_6043);
nand U7887 (N_7887,N_5573,N_6700);
and U7888 (N_7888,N_5148,N_5837);
nand U7889 (N_7889,N_6697,N_5431);
nand U7890 (N_7890,N_5959,N_7284);
or U7891 (N_7891,N_7116,N_7365);
and U7892 (N_7892,N_5184,N_7396);
nand U7893 (N_7893,N_6137,N_7298);
or U7894 (N_7894,N_6518,N_7438);
xor U7895 (N_7895,N_7185,N_5742);
nor U7896 (N_7896,N_6961,N_6497);
xor U7897 (N_7897,N_6165,N_7214);
nor U7898 (N_7898,N_6778,N_7241);
xor U7899 (N_7899,N_5759,N_6958);
xnor U7900 (N_7900,N_6067,N_6076);
and U7901 (N_7901,N_6928,N_7071);
or U7902 (N_7902,N_7056,N_5333);
nor U7903 (N_7903,N_6867,N_6805);
xnor U7904 (N_7904,N_5474,N_6981);
nor U7905 (N_7905,N_6123,N_5449);
nand U7906 (N_7906,N_6547,N_7043);
and U7907 (N_7907,N_7138,N_6829);
or U7908 (N_7908,N_5336,N_5031);
xnor U7909 (N_7909,N_5982,N_5276);
nand U7910 (N_7910,N_5840,N_5566);
and U7911 (N_7911,N_6606,N_7462);
or U7912 (N_7912,N_6193,N_5383);
nand U7913 (N_7913,N_5737,N_6400);
nor U7914 (N_7914,N_5926,N_6772);
xnor U7915 (N_7915,N_6270,N_6850);
nand U7916 (N_7916,N_5802,N_7388);
xnor U7917 (N_7917,N_5515,N_6097);
xor U7918 (N_7918,N_6652,N_5609);
nand U7919 (N_7919,N_7201,N_5376);
and U7920 (N_7920,N_6532,N_5032);
nand U7921 (N_7921,N_6434,N_5807);
nor U7922 (N_7922,N_6459,N_6895);
nand U7923 (N_7923,N_7105,N_6105);
xor U7924 (N_7924,N_5492,N_5436);
xor U7925 (N_7925,N_7400,N_5073);
and U7926 (N_7926,N_6645,N_6823);
nor U7927 (N_7927,N_5285,N_6476);
nand U7928 (N_7928,N_7200,N_7091);
nor U7929 (N_7929,N_6354,N_6487);
or U7930 (N_7930,N_7133,N_6316);
nor U7931 (N_7931,N_5015,N_7399);
or U7932 (N_7932,N_6385,N_6332);
nor U7933 (N_7933,N_6553,N_5789);
xnor U7934 (N_7934,N_5977,N_5966);
or U7935 (N_7935,N_5679,N_6790);
nor U7936 (N_7936,N_5191,N_7072);
nand U7937 (N_7937,N_6290,N_5878);
nand U7938 (N_7938,N_5592,N_6204);
nand U7939 (N_7939,N_6642,N_5927);
and U7940 (N_7940,N_6416,N_6058);
and U7941 (N_7941,N_5374,N_5301);
nand U7942 (N_7942,N_6771,N_6040);
xnor U7943 (N_7943,N_6001,N_7329);
and U7944 (N_7944,N_5654,N_7320);
xnor U7945 (N_7945,N_7032,N_6106);
and U7946 (N_7946,N_6176,N_5068);
or U7947 (N_7947,N_5900,N_5583);
nand U7948 (N_7948,N_6263,N_5916);
xnor U7949 (N_7949,N_5146,N_5637);
xor U7950 (N_7950,N_6392,N_5232);
nand U7951 (N_7951,N_6611,N_6213);
or U7952 (N_7952,N_6366,N_6127);
or U7953 (N_7953,N_6409,N_5831);
nor U7954 (N_7954,N_5310,N_6508);
or U7955 (N_7955,N_7475,N_5125);
and U7956 (N_7956,N_7424,N_5675);
or U7957 (N_7957,N_5425,N_5153);
xor U7958 (N_7958,N_6411,N_5157);
and U7959 (N_7959,N_5908,N_7004);
xor U7960 (N_7960,N_6536,N_6369);
or U7961 (N_7961,N_6228,N_5450);
nor U7962 (N_7962,N_6511,N_5128);
nand U7963 (N_7963,N_6308,N_5754);
or U7964 (N_7964,N_5969,N_5483);
and U7965 (N_7965,N_5606,N_6592);
xor U7966 (N_7966,N_5275,N_5839);
xor U7967 (N_7967,N_6574,N_6664);
nor U7968 (N_7968,N_6470,N_6579);
nand U7969 (N_7969,N_6089,N_6491);
nor U7970 (N_7970,N_7097,N_5962);
or U7971 (N_7971,N_5751,N_7023);
xor U7972 (N_7972,N_6838,N_6003);
nand U7973 (N_7973,N_5862,N_5504);
nand U7974 (N_7974,N_5822,N_6974);
and U7975 (N_7975,N_6899,N_6207);
nor U7976 (N_7976,N_6845,N_6364);
xor U7977 (N_7977,N_6109,N_7443);
or U7978 (N_7978,N_5653,N_7129);
and U7979 (N_7979,N_6297,N_6766);
nor U7980 (N_7980,N_5224,N_5851);
nor U7981 (N_7981,N_6299,N_6842);
nand U7982 (N_7982,N_5631,N_7083);
nor U7983 (N_7983,N_5257,N_7073);
or U7984 (N_7984,N_6111,N_7103);
xor U7985 (N_7985,N_7319,N_7449);
xor U7986 (N_7986,N_5430,N_7347);
or U7987 (N_7987,N_5501,N_5261);
and U7988 (N_7988,N_6448,N_6202);
and U7989 (N_7989,N_6126,N_6622);
and U7990 (N_7990,N_6809,N_6501);
and U7991 (N_7991,N_5404,N_6403);
or U7992 (N_7992,N_5968,N_6189);
and U7993 (N_7993,N_5001,N_5663);
xor U7994 (N_7994,N_6351,N_5989);
and U7995 (N_7995,N_5890,N_6275);
and U7996 (N_7996,N_6698,N_5314);
and U7997 (N_7997,N_6277,N_7213);
nor U7998 (N_7998,N_5561,N_6718);
or U7999 (N_7999,N_6734,N_5196);
or U8000 (N_8000,N_6934,N_5424);
and U8001 (N_8001,N_6372,N_5214);
xnor U8002 (N_8002,N_6245,N_5283);
xor U8003 (N_8003,N_7013,N_5728);
or U8004 (N_8004,N_7442,N_6284);
xor U8005 (N_8005,N_6887,N_6959);
or U8006 (N_8006,N_6510,N_5440);
xor U8007 (N_8007,N_6689,N_7141);
nand U8008 (N_8008,N_6203,N_5178);
xor U8009 (N_8009,N_6768,N_6359);
and U8010 (N_8010,N_5296,N_5611);
nor U8011 (N_8011,N_5535,N_6170);
and U8012 (N_8012,N_6920,N_6912);
nand U8013 (N_8013,N_7495,N_7142);
nor U8014 (N_8014,N_5395,N_6435);
xnor U8015 (N_8015,N_6665,N_6088);
or U8016 (N_8016,N_6593,N_7154);
nor U8017 (N_8017,N_6381,N_5850);
nand U8018 (N_8018,N_6064,N_7096);
or U8019 (N_8019,N_5745,N_6292);
nor U8020 (N_8020,N_6583,N_7426);
and U8021 (N_8021,N_6545,N_6466);
and U8022 (N_8022,N_6084,N_5009);
nand U8023 (N_8023,N_5312,N_7432);
or U8024 (N_8024,N_7406,N_6745);
xnor U8025 (N_8025,N_6865,N_5258);
nor U8026 (N_8026,N_5553,N_6761);
nand U8027 (N_8027,N_7482,N_6007);
and U8028 (N_8028,N_7051,N_6995);
xnor U8029 (N_8029,N_5625,N_5419);
nand U8030 (N_8030,N_6075,N_6880);
or U8031 (N_8031,N_6184,N_6314);
and U8032 (N_8032,N_5696,N_5768);
nor U8033 (N_8033,N_7373,N_6770);
or U8034 (N_8034,N_6627,N_5396);
nand U8035 (N_8035,N_5846,N_7268);
nand U8036 (N_8036,N_5303,N_5359);
and U8037 (N_8037,N_5034,N_6325);
nand U8038 (N_8038,N_7363,N_5572);
nand U8039 (N_8039,N_6011,N_6319);
nor U8040 (N_8040,N_6727,N_5528);
nand U8041 (N_8041,N_7480,N_5264);
nand U8042 (N_8042,N_6239,N_6474);
nor U8043 (N_8043,N_5116,N_5379);
and U8044 (N_8044,N_5996,N_5880);
or U8045 (N_8045,N_7425,N_6846);
xor U8046 (N_8046,N_6340,N_5052);
and U8047 (N_8047,N_7172,N_7183);
or U8048 (N_8048,N_5709,N_5568);
or U8049 (N_8049,N_7028,N_6224);
nor U8050 (N_8050,N_7437,N_5002);
xnor U8051 (N_8051,N_6732,N_6990);
and U8052 (N_8052,N_5243,N_6621);
xnor U8053 (N_8053,N_6955,N_5597);
xor U8054 (N_8054,N_6541,N_7233);
nor U8055 (N_8055,N_5932,N_6512);
and U8056 (N_8056,N_5130,N_7446);
nand U8057 (N_8057,N_5021,N_5661);
and U8058 (N_8058,N_6012,N_5799);
nand U8059 (N_8059,N_5435,N_6035);
nand U8060 (N_8060,N_7128,N_6876);
nand U8061 (N_8061,N_5718,N_5772);
or U8062 (N_8062,N_7029,N_6679);
and U8063 (N_8063,N_7328,N_6045);
and U8064 (N_8064,N_7204,N_7295);
nand U8065 (N_8065,N_5951,N_6478);
or U8066 (N_8066,N_5922,N_6682);
and U8067 (N_8067,N_5557,N_7115);
xnor U8068 (N_8068,N_5271,N_5064);
and U8069 (N_8069,N_5177,N_5921);
xor U8070 (N_8070,N_5527,N_6599);
nand U8071 (N_8071,N_5902,N_6492);
or U8072 (N_8072,N_6254,N_7249);
nor U8073 (N_8073,N_6819,N_6234);
xor U8074 (N_8074,N_5762,N_7226);
xor U8075 (N_8075,N_7024,N_7181);
nor U8076 (N_8076,N_5904,N_5086);
and U8077 (N_8077,N_6504,N_6908);
xnor U8078 (N_8078,N_5168,N_6370);
or U8079 (N_8079,N_6019,N_6367);
nand U8080 (N_8080,N_7009,N_5995);
xnor U8081 (N_8081,N_7285,N_6047);
and U8082 (N_8082,N_6861,N_5438);
and U8083 (N_8083,N_6268,N_6398);
and U8084 (N_8084,N_6129,N_5005);
or U8085 (N_8085,N_5337,N_5526);
nor U8086 (N_8086,N_6486,N_7237);
and U8087 (N_8087,N_6559,N_7031);
xnor U8088 (N_8088,N_6730,N_6485);
nand U8089 (N_8089,N_6605,N_5060);
or U8090 (N_8090,N_6860,N_6675);
xnor U8091 (N_8091,N_6452,N_7109);
nor U8092 (N_8092,N_6632,N_5756);
xor U8093 (N_8093,N_7455,N_6198);
xnor U8094 (N_8094,N_5847,N_5389);
or U8095 (N_8095,N_5250,N_5197);
xor U8096 (N_8096,N_6177,N_7434);
and U8097 (N_8097,N_5212,N_5790);
and U8098 (N_8098,N_5948,N_6883);
xnor U8099 (N_8099,N_7288,N_7483);
xor U8100 (N_8100,N_5269,N_6796);
nand U8101 (N_8101,N_7018,N_7378);
xor U8102 (N_8102,N_6949,N_6266);
nor U8103 (N_8103,N_6395,N_5671);
and U8104 (N_8104,N_5667,N_7332);
xor U8105 (N_8105,N_6969,N_7089);
nor U8106 (N_8106,N_6215,N_5277);
or U8107 (N_8107,N_7301,N_7304);
xor U8108 (N_8108,N_6822,N_5410);
nor U8109 (N_8109,N_6405,N_5327);
xnor U8110 (N_8110,N_5344,N_5869);
or U8111 (N_8111,N_5781,N_6328);
nand U8112 (N_8112,N_5439,N_5131);
and U8113 (N_8113,N_6146,N_6320);
xor U8114 (N_8114,N_6313,N_6653);
xor U8115 (N_8115,N_6140,N_5329);
nor U8116 (N_8116,N_6181,N_6941);
and U8117 (N_8117,N_6853,N_6715);
nor U8118 (N_8118,N_5433,N_6919);
nand U8119 (N_8119,N_5669,N_6138);
xnor U8120 (N_8120,N_7325,N_6851);
nand U8121 (N_8121,N_6125,N_6623);
nand U8122 (N_8122,N_6507,N_6752);
nand U8123 (N_8123,N_6513,N_6130);
or U8124 (N_8124,N_6131,N_6139);
xor U8125 (N_8125,N_5999,N_7366);
or U8126 (N_8126,N_5769,N_6787);
nand U8127 (N_8127,N_5988,N_6580);
xnor U8128 (N_8128,N_7299,N_6963);
and U8129 (N_8129,N_7161,N_7253);
nor U8130 (N_8130,N_6844,N_7110);
and U8131 (N_8131,N_7349,N_7006);
or U8132 (N_8132,N_6527,N_5167);
or U8133 (N_8133,N_6982,N_5701);
or U8134 (N_8134,N_5101,N_7206);
or U8135 (N_8135,N_6849,N_6708);
and U8136 (N_8136,N_6540,N_5205);
xnor U8137 (N_8137,N_6654,N_6641);
nor U8138 (N_8138,N_5541,N_5149);
xnor U8139 (N_8139,N_5714,N_6329);
nor U8140 (N_8140,N_5092,N_6833);
nor U8141 (N_8141,N_6603,N_5466);
nand U8142 (N_8142,N_6233,N_5710);
nand U8143 (N_8143,N_5339,N_6051);
xnor U8144 (N_8144,N_6016,N_6767);
nand U8145 (N_8145,N_7193,N_5599);
and U8146 (N_8146,N_7321,N_6118);
nor U8147 (N_8147,N_6933,N_6683);
nor U8148 (N_8148,N_7261,N_7211);
or U8149 (N_8149,N_6333,N_7330);
and U8150 (N_8150,N_6581,N_7263);
nor U8151 (N_8151,N_6742,N_6135);
and U8152 (N_8152,N_6163,N_6042);
and U8153 (N_8153,N_5532,N_5963);
nand U8154 (N_8154,N_5917,N_6443);
nor U8155 (N_8155,N_6247,N_5266);
xor U8156 (N_8156,N_6989,N_6008);
and U8157 (N_8157,N_6777,N_6628);
and U8158 (N_8158,N_7315,N_5140);
or U8159 (N_8159,N_6454,N_7188);
and U8160 (N_8160,N_6336,N_5227);
nand U8161 (N_8161,N_5981,N_7135);
or U8162 (N_8162,N_6490,N_6175);
and U8163 (N_8163,N_6237,N_6551);
xnor U8164 (N_8164,N_6289,N_5091);
nand U8165 (N_8165,N_6954,N_5910);
nand U8166 (N_8166,N_6701,N_5305);
and U8167 (N_8167,N_5964,N_6391);
and U8168 (N_8168,N_6446,N_6469);
nand U8169 (N_8169,N_7234,N_5845);
nor U8170 (N_8170,N_6195,N_6743);
xor U8171 (N_8171,N_6149,N_6438);
nand U8172 (N_8172,N_6305,N_6607);
xnor U8173 (N_8173,N_7095,N_5987);
and U8174 (N_8174,N_5061,N_7391);
nand U8175 (N_8175,N_5552,N_5235);
nand U8176 (N_8176,N_5112,N_6922);
and U8177 (N_8177,N_6549,N_5505);
or U8178 (N_8178,N_6999,N_5537);
xnor U8179 (N_8179,N_6781,N_6992);
and U8180 (N_8180,N_5730,N_6534);
xnor U8181 (N_8181,N_5095,N_7187);
nor U8182 (N_8182,N_5023,N_6453);
and U8183 (N_8183,N_5209,N_5947);
or U8184 (N_8184,N_5244,N_5418);
nor U8185 (N_8185,N_5295,N_6575);
nand U8186 (N_8186,N_7177,N_7153);
and U8187 (N_8187,N_6597,N_7059);
or U8188 (N_8188,N_5513,N_5897);
nor U8189 (N_8189,N_7108,N_6094);
xor U8190 (N_8190,N_5000,N_7063);
or U8191 (N_8191,N_5477,N_5216);
and U8192 (N_8192,N_5287,N_6280);
and U8193 (N_8193,N_7016,N_6877);
nor U8194 (N_8194,N_6709,N_7111);
or U8195 (N_8195,N_5065,N_7419);
and U8196 (N_8196,N_7422,N_6421);
or U8197 (N_8197,N_6246,N_6624);
nand U8198 (N_8198,N_6212,N_5328);
or U8199 (N_8199,N_5281,N_7436);
xnor U8200 (N_8200,N_5342,N_5797);
nor U8201 (N_8201,N_6209,N_6711);
nand U8202 (N_8202,N_6080,N_6738);
nor U8203 (N_8203,N_6931,N_6107);
xnor U8204 (N_8204,N_5334,N_6010);
and U8205 (N_8205,N_6194,N_6620);
and U8206 (N_8206,N_6379,N_6893);
xor U8207 (N_8207,N_7435,N_6218);
and U8208 (N_8208,N_7252,N_5930);
nand U8209 (N_8209,N_6586,N_5779);
xor U8210 (N_8210,N_5114,N_6712);
xor U8211 (N_8211,N_6160,N_6188);
and U8212 (N_8212,N_5238,N_6975);
and U8213 (N_8213,N_7236,N_5811);
xnor U8214 (N_8214,N_6346,N_5524);
nor U8215 (N_8215,N_6083,N_6171);
and U8216 (N_8216,N_6749,N_6020);
or U8217 (N_8217,N_5693,N_6857);
nand U8218 (N_8218,N_5884,N_7151);
nor U8219 (N_8219,N_7026,N_5752);
nand U8220 (N_8220,N_7117,N_6658);
nand U8221 (N_8221,N_6201,N_5437);
nand U8222 (N_8222,N_5618,N_5249);
and U8223 (N_8223,N_7417,N_7145);
xor U8224 (N_8224,N_7264,N_7242);
nor U8225 (N_8225,N_7405,N_7123);
nand U8226 (N_8226,N_7160,N_6530);
nor U8227 (N_8227,N_7046,N_5369);
or U8228 (N_8228,N_7302,N_6151);
xnor U8229 (N_8229,N_6178,N_5547);
xnor U8230 (N_8230,N_6608,N_6039);
nand U8231 (N_8231,N_5690,N_6006);
nor U8232 (N_8232,N_5488,N_5753);
or U8233 (N_8233,N_5832,N_6706);
xnor U8234 (N_8234,N_7341,N_6296);
nor U8235 (N_8235,N_7445,N_5668);
nor U8236 (N_8236,N_5388,N_6120);
and U8237 (N_8237,N_6962,N_7476);
nor U8238 (N_8238,N_6731,N_7409);
and U8239 (N_8239,N_5780,N_7254);
nor U8240 (N_8240,N_6858,N_6977);
or U8241 (N_8241,N_5480,N_5984);
nor U8242 (N_8242,N_5719,N_5041);
nor U8243 (N_8243,N_5200,N_7077);
nor U8244 (N_8244,N_6377,N_6086);
xnor U8245 (N_8245,N_7343,N_7334);
nor U8246 (N_8246,N_5954,N_6897);
or U8247 (N_8247,N_5458,N_6339);
nand U8248 (N_8248,N_5849,N_5726);
xnor U8249 (N_8249,N_6550,N_5145);
xor U8250 (N_8250,N_7444,N_7238);
nand U8251 (N_8251,N_5007,N_6387);
or U8252 (N_8252,N_7007,N_6947);
and U8253 (N_8253,N_7468,N_6230);
nor U8254 (N_8254,N_5629,N_6894);
and U8255 (N_8255,N_6015,N_5992);
xnor U8256 (N_8256,N_6892,N_6068);
nor U8257 (N_8257,N_5639,N_5872);
or U8258 (N_8258,N_5478,N_7421);
nor U8259 (N_8259,N_7205,N_5360);
xor U8260 (N_8260,N_6072,N_7384);
nand U8261 (N_8261,N_6966,N_7219);
and U8262 (N_8262,N_5868,N_6153);
nand U8263 (N_8263,N_6925,N_7202);
nand U8264 (N_8264,N_7220,N_6287);
xor U8265 (N_8265,N_5102,N_7163);
nand U8266 (N_8266,N_6911,N_5187);
nor U8267 (N_8267,N_5531,N_7112);
or U8268 (N_8268,N_6293,N_5022);
and U8269 (N_8269,N_6240,N_6735);
xor U8270 (N_8270,N_5757,N_7146);
or U8271 (N_8271,N_5546,N_5931);
xnor U8272 (N_8272,N_6660,N_7017);
nor U8273 (N_8273,N_6169,N_7186);
or U8274 (N_8274,N_5161,N_5025);
nand U8275 (N_8275,N_5255,N_7474);
or U8276 (N_8276,N_7136,N_5055);
and U8277 (N_8277,N_5898,N_5795);
nor U8278 (N_8278,N_5313,N_6393);
nand U8279 (N_8279,N_5767,N_5530);
nor U8280 (N_8280,N_5687,N_7382);
nor U8281 (N_8281,N_6748,N_5219);
or U8282 (N_8282,N_5765,N_7093);
and U8283 (N_8283,N_7336,N_5485);
nand U8284 (N_8284,N_6028,N_5763);
and U8285 (N_8285,N_6462,N_6241);
and U8286 (N_8286,N_7376,N_5812);
nor U8287 (N_8287,N_6032,N_6817);
xnor U8288 (N_8288,N_6639,N_6069);
nor U8289 (N_8289,N_5942,N_5357);
nor U8290 (N_8290,N_5457,N_6538);
xor U8291 (N_8291,N_7256,N_6244);
xnor U8292 (N_8292,N_5016,N_5844);
nand U8293 (N_8293,N_5051,N_6253);
nor U8294 (N_8294,N_6864,N_6352);
or U8295 (N_8295,N_6506,N_5949);
nor U8296 (N_8296,N_7050,N_5363);
or U8297 (N_8297,N_6187,N_5189);
nand U8298 (N_8298,N_6414,N_6636);
and U8299 (N_8299,N_5712,N_6820);
or U8300 (N_8300,N_5406,N_6441);
or U8301 (N_8301,N_7413,N_7414);
or U8302 (N_8302,N_7130,N_5808);
xnor U8303 (N_8303,N_5708,N_5506);
or U8304 (N_8304,N_5124,N_6185);
and U8305 (N_8305,N_5965,N_6690);
xnor U8306 (N_8306,N_6985,N_6030);
nand U8307 (N_8307,N_5030,N_6927);
or U8308 (N_8308,N_5817,N_5638);
and U8309 (N_8309,N_5188,N_7060);
nor U8310 (N_8310,N_5689,N_6795);
nand U8311 (N_8311,N_6004,N_5048);
nor U8312 (N_8312,N_5934,N_6917);
xnor U8313 (N_8313,N_5659,N_7139);
and U8314 (N_8314,N_6235,N_5040);
and U8315 (N_8315,N_5482,N_5746);
xnor U8316 (N_8316,N_6248,N_7486);
or U8317 (N_8317,N_6432,N_5107);
nor U8318 (N_8318,N_6262,N_6449);
xnor U8319 (N_8319,N_5225,N_5657);
xnor U8320 (N_8320,N_6323,N_5441);
and U8321 (N_8321,N_5035,N_6498);
nor U8322 (N_8322,N_5087,N_7496);
nand U8323 (N_8323,N_7098,N_7240);
and U8324 (N_8324,N_5432,N_5819);
and U8325 (N_8325,N_6220,N_7078);
or U8326 (N_8326,N_7351,N_5893);
nor U8327 (N_8327,N_6196,N_5788);
and U8328 (N_8328,N_7296,N_5183);
or U8329 (N_8329,N_5382,N_6206);
nor U8330 (N_8330,N_6091,N_6081);
nand U8331 (N_8331,N_6824,N_5509);
xor U8332 (N_8332,N_5635,N_5939);
xor U8333 (N_8333,N_5545,N_5263);
xor U8334 (N_8334,N_5874,N_5166);
nand U8335 (N_8335,N_5691,N_5195);
nor U8336 (N_8336,N_5348,N_6898);
or U8337 (N_8337,N_6686,N_5479);
or U8338 (N_8338,N_7466,N_6214);
xnor U8339 (N_8339,N_5185,N_5129);
nor U8340 (N_8340,N_7165,N_5670);
nand U8341 (N_8341,N_6531,N_7308);
nor U8342 (N_8342,N_6148,N_5297);
and U8343 (N_8343,N_6891,N_6957);
xnor U8344 (N_8344,N_6544,N_6515);
or U8345 (N_8345,N_6413,N_5217);
and U8346 (N_8346,N_6848,N_6430);
or U8347 (N_8347,N_5384,N_7047);
and U8348 (N_8348,N_6884,N_5452);
xor U8349 (N_8349,N_6493,N_5544);
nand U8350 (N_8350,N_5632,N_6855);
nand U8351 (N_8351,N_6814,N_6041);
or U8352 (N_8352,N_5270,N_6382);
nand U8353 (N_8353,N_5353,N_7458);
or U8354 (N_8354,N_7318,N_6840);
nand U8355 (N_8355,N_6021,N_6295);
nor U8356 (N_8356,N_5978,N_6780);
nand U8357 (N_8357,N_6762,N_7055);
nand U8358 (N_8358,N_7196,N_6625);
xnor U8359 (N_8359,N_7180,N_5610);
xor U8360 (N_8360,N_5824,N_5621);
or U8361 (N_8361,N_5705,N_5262);
and U8362 (N_8362,N_6907,N_6389);
xor U8363 (N_8363,N_6788,N_7246);
xnor U8364 (N_8364,N_5427,N_5386);
or U8365 (N_8365,N_5796,N_6368);
and U8366 (N_8366,N_6546,N_7364);
nand U8367 (N_8367,N_5349,N_5093);
and U8368 (N_8368,N_5620,N_6590);
nand U8369 (N_8369,N_5685,N_7232);
and U8370 (N_8370,N_5798,N_5233);
xnor U8371 (N_8371,N_5702,N_6815);
nor U8372 (N_8372,N_5151,N_6227);
or U8373 (N_8373,N_5993,N_5744);
or U8374 (N_8374,N_7244,N_6113);
or U8375 (N_8375,N_5108,N_5859);
nand U8376 (N_8376,N_7277,N_7087);
nor U8377 (N_8377,N_6250,N_6943);
nand U8378 (N_8378,N_6494,N_5598);
or U8379 (N_8379,N_5495,N_5156);
and U8380 (N_8380,N_5213,N_6415);
nand U8381 (N_8381,N_6863,N_5324);
or U8382 (N_8382,N_6503,N_6634);
or U8383 (N_8383,N_6744,N_7020);
and U8384 (N_8384,N_7353,N_6085);
or U8385 (N_8385,N_5174,N_5476);
xor U8386 (N_8386,N_6900,N_5316);
xnor U8387 (N_8387,N_5695,N_6635);
nand U8388 (N_8388,N_5972,N_6423);
nand U8389 (N_8389,N_7143,N_5542);
or U8390 (N_8390,N_6573,N_5641);
nor U8391 (N_8391,N_7428,N_6687);
nor U8392 (N_8392,N_6050,N_7215);
and U8393 (N_8393,N_7286,N_6684);
nor U8394 (N_8394,N_5636,N_6885);
and U8395 (N_8395,N_5267,N_6710);
or U8396 (N_8396,N_6114,N_5991);
or U8397 (N_8397,N_5692,N_6758);
nand U8398 (N_8398,N_7350,N_7402);
and U8399 (N_8399,N_5896,N_7469);
or U8400 (N_8400,N_7171,N_5550);
xor U8401 (N_8401,N_5160,N_6210);
xor U8402 (N_8402,N_5895,N_5867);
nand U8403 (N_8403,N_6948,N_6514);
nor U8404 (N_8404,N_7281,N_7062);
xor U8405 (N_8405,N_5952,N_6594);
xor U8406 (N_8406,N_7119,N_5953);
xnor U8407 (N_8407,N_7258,N_5071);
xor U8408 (N_8408,N_5829,N_5062);
and U8409 (N_8409,N_7148,N_6278);
or U8410 (N_8410,N_7282,N_7218);
nor U8411 (N_8411,N_5888,N_6005);
or U8412 (N_8412,N_5570,N_6096);
and U8413 (N_8413,N_7275,N_5805);
nand U8414 (N_8414,N_6154,N_6755);
and U8415 (N_8415,N_5179,N_5810);
and U8416 (N_8416,N_5612,N_5518);
nor U8417 (N_8417,N_7104,N_6529);
xor U8418 (N_8418,N_6208,N_5853);
or U8419 (N_8419,N_6500,N_5871);
nor U8420 (N_8420,N_5165,N_7389);
xor U8421 (N_8421,N_6264,N_6886);
or U8422 (N_8422,N_6905,N_7390);
nand U8423 (N_8423,N_5738,N_6219);
and U8424 (N_8424,N_6967,N_7393);
and U8425 (N_8425,N_5385,N_5539);
xnor U8426 (N_8426,N_7025,N_6009);
or U8427 (N_8427,N_7015,N_5941);
and U8428 (N_8428,N_5278,N_6944);
nor U8429 (N_8429,N_6018,N_5873);
or U8430 (N_8430,N_5595,N_5886);
and U8431 (N_8431,N_5133,N_5590);
xor U8432 (N_8432,N_7208,N_6807);
or U8433 (N_8433,N_5809,N_6866);
nor U8434 (N_8434,N_5355,N_6801);
xor U8435 (N_8435,N_5821,N_6079);
nand U8436 (N_8436,N_5180,N_5181);
or U8437 (N_8437,N_5594,N_7121);
or U8438 (N_8438,N_7212,N_7137);
or U8439 (N_8439,N_6054,N_5127);
and U8440 (N_8440,N_7019,N_6420);
nor U8441 (N_8441,N_7125,N_6666);
xor U8442 (N_8442,N_5075,N_6798);
or U8443 (N_8443,N_5375,N_5428);
or U8444 (N_8444,N_5306,N_5057);
nand U8445 (N_8445,N_7245,N_5523);
or U8446 (N_8446,N_5986,N_7168);
nor U8447 (N_8447,N_6983,N_5736);
and U8448 (N_8448,N_5920,N_6360);
or U8449 (N_8449,N_6870,N_5522);
nor U8450 (N_8450,N_7166,N_5643);
nor U8451 (N_8451,N_7280,N_5345);
or U8452 (N_8452,N_5894,N_6335);
and U8453 (N_8453,N_5498,N_5204);
xnor U8454 (N_8454,N_7068,N_6036);
or U8455 (N_8455,N_5084,N_5613);
xor U8456 (N_8456,N_6152,N_7131);
or U8457 (N_8457,N_6461,N_5446);
nand U8458 (N_8458,N_7222,N_6695);
or U8459 (N_8459,N_6473,N_7207);
or U8460 (N_8460,N_7292,N_5793);
nor U8461 (N_8461,N_6285,N_6979);
or U8462 (N_8462,N_5245,N_6238);
or U8463 (N_8463,N_6669,N_7397);
and U8464 (N_8464,N_6782,N_6968);
nand U8465 (N_8465,N_5567,N_6451);
nand U8466 (N_8466,N_6813,N_5950);
xor U8467 (N_8467,N_6038,N_5558);
xor U8468 (N_8468,N_6543,N_7198);
nor U8469 (N_8469,N_6914,N_5090);
or U8470 (N_8470,N_6609,N_5619);
nor U8471 (N_8471,N_5536,N_6792);
xor U8472 (N_8472,N_5105,N_5682);
xnor U8473 (N_8473,N_5815,N_5870);
nor U8474 (N_8474,N_6463,N_5656);
nand U8475 (N_8475,N_7317,N_5976);
or U8476 (N_8476,N_6065,N_5230);
xnor U8477 (N_8477,N_6945,N_7338);
or U8478 (N_8478,N_5473,N_6557);
nand U8479 (N_8479,N_7375,N_6315);
nand U8480 (N_8480,N_5077,N_5578);
xor U8481 (N_8481,N_5925,N_7470);
nor U8482 (N_8482,N_7127,N_7398);
nor U8483 (N_8483,N_6099,N_6074);
nor U8484 (N_8484,N_5733,N_5028);
xor U8485 (N_8485,N_7132,N_5860);
nor U8486 (N_8486,N_7092,N_6535);
nand U8487 (N_8487,N_5308,N_5889);
nor U8488 (N_8488,N_7312,N_5700);
nor U8489 (N_8489,N_6396,N_6799);
or U8490 (N_8490,N_6656,N_7036);
nor U8491 (N_8491,N_5318,N_6156);
or U8492 (N_8492,N_7045,N_6837);
or U8493 (N_8493,N_6763,N_6465);
nand U8494 (N_8494,N_5722,N_6505);
nand U8495 (N_8495,N_6906,N_5423);
and U8496 (N_8496,N_6604,N_5698);
and U8497 (N_8497,N_6705,N_7223);
xor U8498 (N_8498,N_6376,N_6773);
or U8499 (N_8499,N_5304,N_6349);
nand U8500 (N_8500,N_5193,N_5928);
and U8501 (N_8501,N_6918,N_5662);
xor U8502 (N_8502,N_6913,N_5724);
nand U8503 (N_8503,N_7410,N_6568);
nor U8504 (N_8504,N_7248,N_5274);
xor U8505 (N_8505,N_5371,N_5442);
or U8506 (N_8506,N_5387,N_5290);
xnor U8507 (N_8507,N_6121,N_7273);
or U8508 (N_8508,N_5175,N_5024);
and U8509 (N_8509,N_6063,N_5731);
and U8510 (N_8510,N_7300,N_6751);
xnor U8511 (N_8511,N_7370,N_7303);
nor U8512 (N_8512,N_5575,N_6267);
xor U8513 (N_8513,N_5403,N_6618);
or U8514 (N_8514,N_6232,N_6477);
or U8515 (N_8515,N_6279,N_7169);
nand U8516 (N_8516,N_5554,N_5616);
or U8517 (N_8517,N_6406,N_6172);
or U8518 (N_8518,N_6161,N_6029);
nand U8519 (N_8519,N_5139,N_5836);
nand U8520 (N_8520,N_6141,N_6037);
nor U8521 (N_8521,N_5771,N_6670);
nand U8522 (N_8522,N_5758,N_6362);
nor U8523 (N_8523,N_7003,N_6548);
nand U8524 (N_8524,N_5778,N_5414);
xor U8525 (N_8525,N_5211,N_6723);
and U8526 (N_8526,N_7473,N_6564);
xnor U8527 (N_8527,N_7358,N_5242);
xor U8528 (N_8528,N_7080,N_7010);
nand U8529 (N_8529,N_5029,N_5881);
xor U8530 (N_8530,N_7167,N_5749);
xnor U8531 (N_8531,N_5857,N_5773);
or U8532 (N_8532,N_6442,N_5288);
or U8533 (N_8533,N_5150,N_6661);
nand U8534 (N_8534,N_6216,N_5655);
and U8535 (N_8535,N_5814,N_5311);
nand U8536 (N_8536,N_5909,N_5806);
or U8537 (N_8537,N_5649,N_6736);
or U8538 (N_8538,N_5367,N_6199);
or U8539 (N_8539,N_5248,N_5104);
nand U8540 (N_8540,N_6910,N_6345);
and U8541 (N_8541,N_6276,N_6357);
xnor U8542 (N_8542,N_5341,N_7279);
xor U8543 (N_8543,N_7385,N_5502);
or U8544 (N_8544,N_6629,N_7331);
and U8545 (N_8545,N_6056,N_6939);
nor U8546 (N_8546,N_7107,N_5046);
nand U8547 (N_8547,N_5067,N_5412);
xnor U8548 (N_8548,N_6450,N_7099);
or U8549 (N_8549,N_5591,N_5323);
nand U8550 (N_8550,N_5887,N_6306);
or U8551 (N_8551,N_6909,N_6986);
xor U8552 (N_8552,N_5006,N_6122);
nand U8553 (N_8553,N_6724,N_6924);
nor U8554 (N_8554,N_7457,N_5470);
and U8555 (N_8555,N_5332,N_5514);
nand U8556 (N_8556,N_7427,N_5058);
nor U8557 (N_8557,N_5924,N_5471);
and U8558 (N_8558,N_6217,N_5119);
xor U8559 (N_8559,N_5206,N_6258);
or U8560 (N_8560,N_5497,N_6935);
or U8561 (N_8561,N_5147,N_6186);
and U8562 (N_8562,N_7152,N_5564);
or U8563 (N_8563,N_5923,N_7113);
nor U8564 (N_8564,N_5579,N_5913);
nor U8565 (N_8565,N_5642,N_6640);
or U8566 (N_8566,N_6971,N_6108);
and U8567 (N_8567,N_6053,N_5378);
nand U8568 (N_8568,N_5587,N_7381);
xor U8569 (N_8569,N_5960,N_5764);
nor U8570 (N_8570,N_7040,N_6582);
nand U8571 (N_8571,N_5588,N_5019);
and U8572 (N_8572,N_5835,N_6255);
nand U8573 (N_8573,N_5380,N_5014);
xor U8574 (N_8574,N_6717,N_5256);
and U8575 (N_8575,N_5008,N_6274);
and U8576 (N_8576,N_6288,N_6600);
nand U8577 (N_8577,N_5455,N_7079);
or U8578 (N_8578,N_5727,N_5229);
xnor U8579 (N_8579,N_7479,N_6093);
nor U8580 (N_8580,N_6327,N_5645);
nor U8581 (N_8581,N_5162,N_5475);
nand U8582 (N_8582,N_6713,N_6566);
nor U8583 (N_8583,N_5411,N_5142);
nand U8584 (N_8584,N_5593,N_6521);
xor U8585 (N_8585,N_6936,N_5660);
nor U8586 (N_8586,N_5172,N_6291);
or U8587 (N_8587,N_7488,N_5115);
nor U8588 (N_8588,N_6874,N_7327);
nand U8589 (N_8589,N_6271,N_6117);
nand U8590 (N_8590,N_6390,N_5393);
nand U8591 (N_8591,N_5551,N_6614);
nand U8592 (N_8592,N_6101,N_6242);
nor U8593 (N_8593,N_6166,N_6854);
nand U8594 (N_8594,N_5201,N_6162);
or U8595 (N_8595,N_5254,N_7494);
xor U8596 (N_8596,N_5651,N_6457);
and U8597 (N_8597,N_6694,N_7310);
and U8598 (N_8598,N_5487,N_7283);
and U8599 (N_8599,N_7011,N_7247);
or U8600 (N_8600,N_5117,N_6044);
xor U8601 (N_8601,N_5486,N_5182);
or U8602 (N_8602,N_6077,N_5664);
nand U8603 (N_8603,N_6737,N_5582);
nor U8604 (N_8604,N_6754,N_7411);
and U8605 (N_8605,N_7401,N_5137);
or U8606 (N_8606,N_5747,N_6249);
nor U8607 (N_8607,N_5109,N_6843);
nand U8608 (N_8608,N_6896,N_5322);
nand U8609 (N_8609,N_7191,N_5652);
xnor U8610 (N_8610,N_6881,N_6150);
nor U8611 (N_8611,N_5231,N_5163);
and U8612 (N_8612,N_7270,N_6440);
nor U8613 (N_8613,N_5732,N_6681);
nand U8614 (N_8614,N_5053,N_6355);
nor U8615 (N_8615,N_5218,N_5761);
xnor U8616 (N_8616,N_5171,N_6929);
or U8617 (N_8617,N_7293,N_5828);
and U8618 (N_8618,N_5390,N_5265);
and U8619 (N_8619,N_6404,N_6002);
or U8620 (N_8620,N_6938,N_5804);
nor U8621 (N_8621,N_6716,N_5399);
nor U8622 (N_8622,N_5307,N_5491);
or U8623 (N_8623,N_6825,N_6785);
and U8624 (N_8624,N_6926,N_6818);
nor U8625 (N_8625,N_5352,N_7485);
xnor U8626 (N_8626,N_7416,N_5848);
nor U8627 (N_8627,N_5729,N_6143);
or U8628 (N_8628,N_6183,N_5565);
nor U8629 (N_8629,N_6321,N_7102);
nor U8630 (N_8630,N_6386,N_6793);
and U8631 (N_8631,N_7465,N_5678);
xnor U8632 (N_8632,N_6326,N_5596);
xnor U8633 (N_8633,N_5325,N_5320);
xor U8634 (N_8634,N_6499,N_7230);
xnor U8635 (N_8635,N_6533,N_7192);
nor U8636 (N_8636,N_7094,N_5627);
xor U8637 (N_8637,N_5300,N_6776);
and U8638 (N_8638,N_5983,N_6167);
or U8639 (N_8639,N_5907,N_5004);
or U8640 (N_8640,N_6243,N_6965);
and U8641 (N_8641,N_5394,N_5207);
and U8642 (N_8642,N_5600,N_5397);
nand U8643 (N_8643,N_7225,N_5044);
nand U8644 (N_8644,N_5279,N_5392);
nor U8645 (N_8645,N_5775,N_7257);
nor U8646 (N_8646,N_7352,N_5070);
xor U8647 (N_8647,N_6307,N_6946);
nand U8648 (N_8648,N_5929,N_5259);
nand U8649 (N_8649,N_5580,N_5694);
nor U8650 (N_8650,N_6571,N_6655);
and U8651 (N_8651,N_5422,N_6119);
and U8652 (N_8652,N_5512,N_6520);
nor U8653 (N_8653,N_6522,N_5569);
or U8654 (N_8654,N_6132,N_6643);
and U8655 (N_8655,N_6972,N_6616);
xor U8656 (N_8656,N_7383,N_7022);
or U8657 (N_8657,N_5791,N_5111);
xnor U8658 (N_8658,N_5122,N_6100);
or U8659 (N_8659,N_6222,N_5623);
xnor U8660 (N_8660,N_5268,N_7294);
or U8661 (N_8661,N_6862,N_6693);
nand U8662 (N_8662,N_6775,N_6873);
or U8663 (N_8663,N_5604,N_6740);
and U8664 (N_8664,N_5100,N_6073);
or U8665 (N_8665,N_6960,N_6956);
nand U8666 (N_8666,N_5734,N_6471);
or U8667 (N_8667,N_5228,N_5648);
and U8668 (N_8668,N_6229,N_6048);
or U8669 (N_8669,N_6552,N_6726);
and U8670 (N_8670,N_7057,N_5226);
nor U8671 (N_8671,N_7431,N_5901);
xnor U8672 (N_8672,N_6589,N_6066);
or U8673 (N_8673,N_6444,N_5072);
and U8674 (N_8674,N_6901,N_5170);
nand U8675 (N_8675,N_6836,N_5581);
and U8676 (N_8676,N_5429,N_5159);
xor U8677 (N_8677,N_5398,N_5879);
or U8678 (N_8678,N_5586,N_5559);
or U8679 (N_8679,N_5674,N_6031);
or U8680 (N_8680,N_5538,N_6868);
nand U8681 (N_8681,N_5990,N_6964);
or U8682 (N_8682,N_5017,N_5956);
and U8683 (N_8683,N_6769,N_7126);
xnor U8684 (N_8684,N_6577,N_7184);
nand U8685 (N_8685,N_6034,N_6523);
or U8686 (N_8686,N_5915,N_6674);
and U8687 (N_8687,N_5885,N_6182);
or U8688 (N_8688,N_7387,N_5113);
and U8689 (N_8689,N_6304,N_5294);
nor U8690 (N_8690,N_5680,N_5309);
nor U8691 (N_8691,N_5760,N_6720);
nor U8692 (N_8692,N_5584,N_6869);
or U8693 (N_8693,N_5525,N_5199);
nand U8694 (N_8694,N_7345,N_7021);
xor U8695 (N_8695,N_7374,N_6426);
xnor U8696 (N_8696,N_6269,N_6797);
or U8697 (N_8697,N_5176,N_6324);
xor U8698 (N_8698,N_5097,N_6859);
or U8699 (N_8699,N_7090,N_5391);
and U8700 (N_8700,N_5686,N_6647);
or U8701 (N_8701,N_6703,N_5858);
nand U8702 (N_8702,N_5830,N_6272);
nor U8703 (N_8703,N_5208,N_5453);
and U8704 (N_8704,N_6554,N_6311);
and U8705 (N_8705,N_7231,N_5063);
nor U8706 (N_8706,N_5626,N_5666);
or U8707 (N_8707,N_6437,N_5574);
nor U8708 (N_8708,N_7158,N_5481);
nand U8709 (N_8709,N_5571,N_7297);
and U8710 (N_8710,N_7333,N_5589);
xor U8711 (N_8711,N_7490,N_5164);
or U8712 (N_8712,N_6483,N_7403);
nand U8713 (N_8713,N_6739,N_6509);
nand U8714 (N_8714,N_6991,N_6839);
nand U8715 (N_8715,N_6425,N_5134);
nor U8716 (N_8716,N_7306,N_7274);
and U8717 (N_8717,N_6663,N_5640);
or U8718 (N_8718,N_5876,N_7058);
and U8719 (N_8719,N_6000,N_6759);
or U8720 (N_8720,N_6251,N_6585);
nand U8721 (N_8721,N_6281,N_5519);
and U8722 (N_8722,N_7461,N_6760);
xnor U8723 (N_8723,N_5121,N_7362);
xor U8724 (N_8724,N_6022,N_7433);
and U8725 (N_8725,N_7359,N_5420);
nand U8726 (N_8726,N_6027,N_5099);
nand U8727 (N_8727,N_7267,N_6082);
xnor U8728 (N_8728,N_5082,N_6365);
nor U8729 (N_8729,N_7259,N_6456);
nand U8730 (N_8730,N_7227,N_5936);
xor U8731 (N_8731,N_6657,N_6422);
or U8732 (N_8732,N_6023,N_6973);
or U8733 (N_8733,N_6164,N_6310);
and U8734 (N_8734,N_7418,N_5826);
or U8735 (N_8735,N_5842,N_7346);
xnor U8736 (N_8736,N_6489,N_6092);
xor U8737 (N_8737,N_5158,N_5358);
or U8738 (N_8738,N_6806,N_5083);
nor U8739 (N_8739,N_5955,N_5740);
xor U8740 (N_8740,N_6572,N_6300);
nor U8741 (N_8741,N_5463,N_7481);
and U8742 (N_8742,N_5253,N_7493);
nand U8743 (N_8743,N_5935,N_5202);
and U8744 (N_8744,N_7038,N_6318);
xor U8745 (N_8745,N_7289,N_6650);
or U8746 (N_8746,N_5282,N_6808);
xnor U8747 (N_8747,N_6116,N_5721);
or U8748 (N_8748,N_6702,N_5417);
xnor U8749 (N_8749,N_6373,N_6560);
nor U8750 (N_8750,N_6469,N_5568);
xnor U8751 (N_8751,N_7188,N_6319);
nand U8752 (N_8752,N_7041,N_5727);
nand U8753 (N_8753,N_6188,N_5166);
or U8754 (N_8754,N_6621,N_6649);
xor U8755 (N_8755,N_6533,N_5435);
xor U8756 (N_8756,N_6144,N_5955);
nor U8757 (N_8757,N_7085,N_6087);
nor U8758 (N_8758,N_5555,N_6500);
or U8759 (N_8759,N_7014,N_5151);
or U8760 (N_8760,N_5943,N_6965);
and U8761 (N_8761,N_5998,N_5217);
or U8762 (N_8762,N_5134,N_7369);
and U8763 (N_8763,N_6248,N_5187);
nand U8764 (N_8764,N_7361,N_5956);
and U8765 (N_8765,N_5759,N_6932);
xor U8766 (N_8766,N_6807,N_5500);
or U8767 (N_8767,N_5092,N_5867);
and U8768 (N_8768,N_6126,N_6961);
xor U8769 (N_8769,N_5237,N_5354);
nand U8770 (N_8770,N_7492,N_5938);
and U8771 (N_8771,N_5319,N_6890);
or U8772 (N_8772,N_5310,N_7111);
or U8773 (N_8773,N_6724,N_6375);
or U8774 (N_8774,N_5467,N_5437);
or U8775 (N_8775,N_5700,N_5965);
nor U8776 (N_8776,N_5042,N_5624);
nor U8777 (N_8777,N_5607,N_7257);
xor U8778 (N_8778,N_6271,N_6886);
and U8779 (N_8779,N_7179,N_6739);
and U8780 (N_8780,N_6373,N_5595);
nor U8781 (N_8781,N_7450,N_6632);
and U8782 (N_8782,N_5302,N_5099);
and U8783 (N_8783,N_6498,N_5936);
or U8784 (N_8784,N_5094,N_7288);
nand U8785 (N_8785,N_5710,N_5275);
xor U8786 (N_8786,N_6748,N_6779);
nor U8787 (N_8787,N_6020,N_5385);
xnor U8788 (N_8788,N_5883,N_6006);
nor U8789 (N_8789,N_6673,N_6996);
nor U8790 (N_8790,N_6693,N_6965);
and U8791 (N_8791,N_5346,N_6250);
or U8792 (N_8792,N_7099,N_7398);
xnor U8793 (N_8793,N_6914,N_6812);
or U8794 (N_8794,N_6565,N_5217);
and U8795 (N_8795,N_6126,N_5535);
or U8796 (N_8796,N_6070,N_5968);
nor U8797 (N_8797,N_6307,N_5464);
xnor U8798 (N_8798,N_6418,N_6124);
xor U8799 (N_8799,N_5910,N_5082);
nand U8800 (N_8800,N_6067,N_6083);
nor U8801 (N_8801,N_7427,N_5271);
nor U8802 (N_8802,N_7032,N_5290);
nand U8803 (N_8803,N_6920,N_6000);
nand U8804 (N_8804,N_7425,N_7217);
and U8805 (N_8805,N_5275,N_7440);
nor U8806 (N_8806,N_5584,N_7494);
and U8807 (N_8807,N_5567,N_6292);
and U8808 (N_8808,N_5758,N_6383);
and U8809 (N_8809,N_6931,N_5053);
and U8810 (N_8810,N_5909,N_5255);
xor U8811 (N_8811,N_6296,N_6932);
xnor U8812 (N_8812,N_6873,N_5078);
nand U8813 (N_8813,N_6903,N_7454);
xor U8814 (N_8814,N_5407,N_5917);
and U8815 (N_8815,N_7005,N_5630);
xor U8816 (N_8816,N_5795,N_5729);
nand U8817 (N_8817,N_5103,N_7357);
xnor U8818 (N_8818,N_6227,N_6298);
nand U8819 (N_8819,N_5599,N_6203);
nor U8820 (N_8820,N_5912,N_5253);
nand U8821 (N_8821,N_6269,N_7427);
or U8822 (N_8822,N_6871,N_5375);
and U8823 (N_8823,N_7436,N_6068);
or U8824 (N_8824,N_7189,N_5223);
xor U8825 (N_8825,N_5998,N_7497);
nand U8826 (N_8826,N_5360,N_6031);
or U8827 (N_8827,N_5398,N_6292);
nand U8828 (N_8828,N_6856,N_6396);
nor U8829 (N_8829,N_5240,N_6397);
xnor U8830 (N_8830,N_5078,N_7492);
or U8831 (N_8831,N_5101,N_6247);
xnor U8832 (N_8832,N_7109,N_7143);
or U8833 (N_8833,N_6377,N_7165);
or U8834 (N_8834,N_6575,N_6027);
and U8835 (N_8835,N_6988,N_6618);
nand U8836 (N_8836,N_5281,N_6981);
or U8837 (N_8837,N_6719,N_5649);
xor U8838 (N_8838,N_6710,N_6774);
nand U8839 (N_8839,N_5975,N_7232);
and U8840 (N_8840,N_5195,N_5876);
xor U8841 (N_8841,N_5408,N_7389);
xor U8842 (N_8842,N_6318,N_5560);
nor U8843 (N_8843,N_6324,N_6237);
or U8844 (N_8844,N_7357,N_5504);
nand U8845 (N_8845,N_6327,N_7133);
xnor U8846 (N_8846,N_6905,N_6522);
and U8847 (N_8847,N_6863,N_6060);
and U8848 (N_8848,N_7077,N_5584);
or U8849 (N_8849,N_6777,N_6900);
nand U8850 (N_8850,N_5958,N_6011);
xnor U8851 (N_8851,N_7268,N_6205);
nand U8852 (N_8852,N_5224,N_5282);
and U8853 (N_8853,N_6765,N_5484);
xor U8854 (N_8854,N_5212,N_6370);
and U8855 (N_8855,N_5642,N_7446);
or U8856 (N_8856,N_5264,N_6615);
and U8857 (N_8857,N_6384,N_7456);
xnor U8858 (N_8858,N_5968,N_6934);
nand U8859 (N_8859,N_6108,N_7338);
nor U8860 (N_8860,N_5163,N_5239);
xor U8861 (N_8861,N_5933,N_5338);
nand U8862 (N_8862,N_6178,N_6175);
xnor U8863 (N_8863,N_7242,N_5176);
xnor U8864 (N_8864,N_7065,N_7280);
nand U8865 (N_8865,N_5786,N_6119);
and U8866 (N_8866,N_6969,N_6475);
or U8867 (N_8867,N_6882,N_6658);
nor U8868 (N_8868,N_6357,N_7147);
and U8869 (N_8869,N_6660,N_6734);
and U8870 (N_8870,N_5878,N_7120);
or U8871 (N_8871,N_5880,N_5148);
nand U8872 (N_8872,N_5950,N_6358);
nand U8873 (N_8873,N_7289,N_5372);
xnor U8874 (N_8874,N_5051,N_7036);
nor U8875 (N_8875,N_5702,N_6230);
and U8876 (N_8876,N_5483,N_7099);
nand U8877 (N_8877,N_6285,N_6089);
or U8878 (N_8878,N_7473,N_6274);
nor U8879 (N_8879,N_5814,N_5141);
xnor U8880 (N_8880,N_5742,N_6529);
or U8881 (N_8881,N_7039,N_6034);
xnor U8882 (N_8882,N_5802,N_6691);
xnor U8883 (N_8883,N_6422,N_6337);
or U8884 (N_8884,N_6858,N_6751);
xor U8885 (N_8885,N_6975,N_7414);
xnor U8886 (N_8886,N_5955,N_5382);
and U8887 (N_8887,N_5490,N_5771);
nand U8888 (N_8888,N_6665,N_6009);
xor U8889 (N_8889,N_6125,N_7480);
nand U8890 (N_8890,N_5761,N_7437);
xnor U8891 (N_8891,N_5961,N_7263);
or U8892 (N_8892,N_5772,N_6984);
nand U8893 (N_8893,N_7023,N_5538);
xor U8894 (N_8894,N_5070,N_7017);
xnor U8895 (N_8895,N_5688,N_5229);
xor U8896 (N_8896,N_5667,N_5794);
nand U8897 (N_8897,N_5394,N_6817);
nor U8898 (N_8898,N_5745,N_5689);
nand U8899 (N_8899,N_5171,N_6736);
xnor U8900 (N_8900,N_7220,N_5735);
xor U8901 (N_8901,N_6829,N_7474);
and U8902 (N_8902,N_6565,N_5417);
and U8903 (N_8903,N_5499,N_7223);
or U8904 (N_8904,N_7001,N_6516);
xor U8905 (N_8905,N_7092,N_6259);
xnor U8906 (N_8906,N_6543,N_6013);
xor U8907 (N_8907,N_7158,N_6401);
nand U8908 (N_8908,N_5512,N_7411);
xnor U8909 (N_8909,N_5952,N_6710);
or U8910 (N_8910,N_6624,N_6036);
nor U8911 (N_8911,N_6029,N_7360);
nand U8912 (N_8912,N_6315,N_5280);
nand U8913 (N_8913,N_6773,N_6246);
and U8914 (N_8914,N_5375,N_5113);
xor U8915 (N_8915,N_5127,N_5095);
and U8916 (N_8916,N_6862,N_5017);
nor U8917 (N_8917,N_5276,N_5845);
or U8918 (N_8918,N_5931,N_5900);
nor U8919 (N_8919,N_5520,N_6646);
nor U8920 (N_8920,N_6796,N_7078);
xnor U8921 (N_8921,N_5664,N_6010);
or U8922 (N_8922,N_5087,N_5556);
xor U8923 (N_8923,N_6166,N_5314);
nor U8924 (N_8924,N_5724,N_6431);
or U8925 (N_8925,N_5839,N_7416);
xor U8926 (N_8926,N_5521,N_5622);
or U8927 (N_8927,N_6331,N_6769);
and U8928 (N_8928,N_5580,N_5404);
nor U8929 (N_8929,N_6291,N_5376);
nand U8930 (N_8930,N_6160,N_7401);
nand U8931 (N_8931,N_6377,N_6070);
xnor U8932 (N_8932,N_6752,N_6588);
and U8933 (N_8933,N_5160,N_5824);
xnor U8934 (N_8934,N_7034,N_7094);
or U8935 (N_8935,N_6240,N_6708);
xor U8936 (N_8936,N_6407,N_5013);
and U8937 (N_8937,N_5106,N_7024);
or U8938 (N_8938,N_6251,N_7001);
or U8939 (N_8939,N_5099,N_5939);
xnor U8940 (N_8940,N_5966,N_6609);
nand U8941 (N_8941,N_7002,N_7236);
and U8942 (N_8942,N_7455,N_7121);
xnor U8943 (N_8943,N_6128,N_6180);
and U8944 (N_8944,N_5978,N_7215);
or U8945 (N_8945,N_5585,N_6349);
or U8946 (N_8946,N_5479,N_5507);
or U8947 (N_8947,N_7203,N_5246);
nand U8948 (N_8948,N_7134,N_6259);
nor U8949 (N_8949,N_6484,N_6706);
and U8950 (N_8950,N_5995,N_5765);
nand U8951 (N_8951,N_7425,N_5065);
or U8952 (N_8952,N_6242,N_5094);
or U8953 (N_8953,N_6994,N_5703);
nor U8954 (N_8954,N_5488,N_6286);
nand U8955 (N_8955,N_5770,N_5554);
and U8956 (N_8956,N_6581,N_5811);
xor U8957 (N_8957,N_7352,N_7003);
or U8958 (N_8958,N_6240,N_6037);
and U8959 (N_8959,N_5303,N_5097);
nor U8960 (N_8960,N_6115,N_7319);
nor U8961 (N_8961,N_5022,N_6522);
nor U8962 (N_8962,N_7175,N_6337);
nor U8963 (N_8963,N_7016,N_5730);
and U8964 (N_8964,N_5396,N_6005);
or U8965 (N_8965,N_7133,N_7015);
and U8966 (N_8966,N_5901,N_7247);
and U8967 (N_8967,N_5032,N_6136);
xnor U8968 (N_8968,N_6433,N_6583);
nand U8969 (N_8969,N_5256,N_7275);
xor U8970 (N_8970,N_6976,N_6594);
or U8971 (N_8971,N_7325,N_6185);
nor U8972 (N_8972,N_6334,N_6403);
xnor U8973 (N_8973,N_6543,N_5587);
nor U8974 (N_8974,N_7033,N_7391);
xor U8975 (N_8975,N_5256,N_5229);
and U8976 (N_8976,N_7197,N_5561);
or U8977 (N_8977,N_5603,N_7253);
nand U8978 (N_8978,N_7456,N_6171);
and U8979 (N_8979,N_7184,N_7410);
and U8980 (N_8980,N_6451,N_6013);
nand U8981 (N_8981,N_5316,N_6467);
and U8982 (N_8982,N_5888,N_6680);
nor U8983 (N_8983,N_5230,N_6197);
and U8984 (N_8984,N_7115,N_5417);
and U8985 (N_8985,N_5873,N_6489);
nand U8986 (N_8986,N_7359,N_6364);
or U8987 (N_8987,N_5858,N_5570);
nand U8988 (N_8988,N_7105,N_7346);
nand U8989 (N_8989,N_5763,N_5941);
or U8990 (N_8990,N_7260,N_5057);
nor U8991 (N_8991,N_6255,N_5894);
and U8992 (N_8992,N_5681,N_5231);
or U8993 (N_8993,N_6810,N_5586);
nor U8994 (N_8994,N_6937,N_6471);
nor U8995 (N_8995,N_6921,N_7022);
and U8996 (N_8996,N_7249,N_6665);
nand U8997 (N_8997,N_5118,N_6689);
or U8998 (N_8998,N_7404,N_7161);
and U8999 (N_8999,N_6814,N_6480);
nand U9000 (N_9000,N_6132,N_6033);
or U9001 (N_9001,N_5173,N_5370);
nand U9002 (N_9002,N_7467,N_5155);
nor U9003 (N_9003,N_7149,N_7342);
nor U9004 (N_9004,N_6059,N_6434);
nand U9005 (N_9005,N_6835,N_7350);
or U9006 (N_9006,N_5989,N_5610);
nor U9007 (N_9007,N_7232,N_5414);
nor U9008 (N_9008,N_5665,N_5208);
and U9009 (N_9009,N_6250,N_5954);
nor U9010 (N_9010,N_5614,N_6894);
xnor U9011 (N_9011,N_6805,N_6041);
and U9012 (N_9012,N_5014,N_6990);
or U9013 (N_9013,N_5716,N_7023);
or U9014 (N_9014,N_6644,N_7295);
nor U9015 (N_9015,N_5419,N_6856);
xnor U9016 (N_9016,N_7219,N_6413);
nor U9017 (N_9017,N_5729,N_5244);
and U9018 (N_9018,N_6865,N_5213);
and U9019 (N_9019,N_5389,N_6782);
nand U9020 (N_9020,N_7091,N_7163);
nand U9021 (N_9021,N_5122,N_6561);
nor U9022 (N_9022,N_6995,N_6315);
nand U9023 (N_9023,N_6700,N_5560);
or U9024 (N_9024,N_6770,N_6942);
or U9025 (N_9025,N_5594,N_7257);
and U9026 (N_9026,N_6508,N_7232);
xor U9027 (N_9027,N_5890,N_6207);
nand U9028 (N_9028,N_6933,N_7331);
xnor U9029 (N_9029,N_5747,N_5665);
or U9030 (N_9030,N_6441,N_6904);
or U9031 (N_9031,N_6261,N_6937);
or U9032 (N_9032,N_6381,N_5013);
or U9033 (N_9033,N_6635,N_5289);
and U9034 (N_9034,N_5190,N_6977);
xor U9035 (N_9035,N_7241,N_5724);
or U9036 (N_9036,N_5627,N_6729);
nand U9037 (N_9037,N_5682,N_6975);
nor U9038 (N_9038,N_5775,N_7279);
xnor U9039 (N_9039,N_6177,N_6673);
nor U9040 (N_9040,N_5035,N_5209);
and U9041 (N_9041,N_6368,N_5742);
or U9042 (N_9042,N_6292,N_6956);
or U9043 (N_9043,N_6959,N_5221);
and U9044 (N_9044,N_6900,N_6862);
nor U9045 (N_9045,N_6371,N_7399);
and U9046 (N_9046,N_6261,N_5675);
xnor U9047 (N_9047,N_6763,N_5771);
and U9048 (N_9048,N_5994,N_5425);
nor U9049 (N_9049,N_5263,N_6108);
nor U9050 (N_9050,N_6168,N_7393);
xnor U9051 (N_9051,N_6482,N_7119);
xor U9052 (N_9052,N_5811,N_5795);
and U9053 (N_9053,N_5587,N_7402);
or U9054 (N_9054,N_7216,N_6140);
or U9055 (N_9055,N_6682,N_6999);
and U9056 (N_9056,N_6934,N_5441);
and U9057 (N_9057,N_5215,N_6171);
or U9058 (N_9058,N_5002,N_6248);
and U9059 (N_9059,N_6022,N_5677);
and U9060 (N_9060,N_7304,N_6378);
nor U9061 (N_9061,N_5971,N_7230);
and U9062 (N_9062,N_7295,N_5499);
nand U9063 (N_9063,N_6444,N_5064);
nor U9064 (N_9064,N_5841,N_7082);
nor U9065 (N_9065,N_7138,N_5559);
and U9066 (N_9066,N_5858,N_5089);
nand U9067 (N_9067,N_5975,N_5416);
or U9068 (N_9068,N_6520,N_6769);
and U9069 (N_9069,N_6666,N_6203);
xor U9070 (N_9070,N_5437,N_5341);
or U9071 (N_9071,N_6968,N_5551);
and U9072 (N_9072,N_6087,N_5541);
nand U9073 (N_9073,N_6861,N_5621);
xnor U9074 (N_9074,N_5195,N_6066);
xor U9075 (N_9075,N_6032,N_6203);
xnor U9076 (N_9076,N_6127,N_6819);
and U9077 (N_9077,N_5803,N_5592);
and U9078 (N_9078,N_5637,N_5792);
xnor U9079 (N_9079,N_6854,N_5832);
xor U9080 (N_9080,N_5125,N_5858);
nor U9081 (N_9081,N_6620,N_7097);
nor U9082 (N_9082,N_6426,N_5701);
and U9083 (N_9083,N_6922,N_7312);
nor U9084 (N_9084,N_7357,N_5084);
xnor U9085 (N_9085,N_5599,N_5122);
nand U9086 (N_9086,N_5048,N_6071);
xnor U9087 (N_9087,N_6002,N_5248);
nor U9088 (N_9088,N_5800,N_6523);
and U9089 (N_9089,N_6444,N_6453);
and U9090 (N_9090,N_5239,N_5445);
and U9091 (N_9091,N_5159,N_5735);
nor U9092 (N_9092,N_5005,N_6311);
xnor U9093 (N_9093,N_5916,N_6663);
and U9094 (N_9094,N_6702,N_6856);
and U9095 (N_9095,N_7186,N_5874);
xor U9096 (N_9096,N_6463,N_6751);
nor U9097 (N_9097,N_6538,N_7001);
nor U9098 (N_9098,N_6248,N_5267);
xor U9099 (N_9099,N_5898,N_5199);
or U9100 (N_9100,N_6295,N_6091);
and U9101 (N_9101,N_5757,N_6113);
nand U9102 (N_9102,N_7230,N_6539);
xnor U9103 (N_9103,N_7463,N_6849);
nor U9104 (N_9104,N_6642,N_5478);
xnor U9105 (N_9105,N_7121,N_5526);
nor U9106 (N_9106,N_5329,N_5059);
xor U9107 (N_9107,N_7008,N_6788);
and U9108 (N_9108,N_6343,N_6842);
xor U9109 (N_9109,N_5362,N_7330);
nor U9110 (N_9110,N_6380,N_5408);
nand U9111 (N_9111,N_5453,N_7456);
nor U9112 (N_9112,N_6905,N_5017);
xnor U9113 (N_9113,N_5016,N_6634);
nor U9114 (N_9114,N_5124,N_5067);
or U9115 (N_9115,N_5404,N_7094);
and U9116 (N_9116,N_6106,N_5233);
or U9117 (N_9117,N_6831,N_5788);
xnor U9118 (N_9118,N_7411,N_5650);
nor U9119 (N_9119,N_6126,N_6342);
xor U9120 (N_9120,N_5200,N_7163);
xnor U9121 (N_9121,N_5823,N_5314);
nor U9122 (N_9122,N_6077,N_6739);
nand U9123 (N_9123,N_7007,N_6614);
or U9124 (N_9124,N_6108,N_5112);
or U9125 (N_9125,N_5193,N_5403);
nor U9126 (N_9126,N_5490,N_7209);
or U9127 (N_9127,N_6404,N_6564);
nor U9128 (N_9128,N_5449,N_7140);
xor U9129 (N_9129,N_6956,N_6116);
or U9130 (N_9130,N_5368,N_7022);
and U9131 (N_9131,N_6031,N_6444);
nand U9132 (N_9132,N_5535,N_5224);
and U9133 (N_9133,N_7309,N_6572);
or U9134 (N_9134,N_7473,N_7141);
and U9135 (N_9135,N_6776,N_6657);
nor U9136 (N_9136,N_5064,N_5195);
nor U9137 (N_9137,N_7490,N_5449);
xor U9138 (N_9138,N_5189,N_7068);
nor U9139 (N_9139,N_5786,N_6574);
nor U9140 (N_9140,N_6158,N_5945);
or U9141 (N_9141,N_5528,N_5267);
or U9142 (N_9142,N_6683,N_5240);
or U9143 (N_9143,N_5054,N_5186);
nor U9144 (N_9144,N_5470,N_6820);
nor U9145 (N_9145,N_7097,N_7157);
nor U9146 (N_9146,N_5610,N_7069);
nor U9147 (N_9147,N_5989,N_6998);
and U9148 (N_9148,N_5009,N_7194);
or U9149 (N_9149,N_7005,N_5711);
nor U9150 (N_9150,N_6152,N_6396);
xor U9151 (N_9151,N_5695,N_6410);
or U9152 (N_9152,N_6094,N_5266);
xor U9153 (N_9153,N_5492,N_5637);
or U9154 (N_9154,N_6933,N_6758);
nor U9155 (N_9155,N_5073,N_6138);
or U9156 (N_9156,N_6821,N_6764);
or U9157 (N_9157,N_7234,N_6867);
or U9158 (N_9158,N_5563,N_6707);
nand U9159 (N_9159,N_5517,N_6701);
nor U9160 (N_9160,N_5220,N_5065);
or U9161 (N_9161,N_5901,N_5860);
nand U9162 (N_9162,N_7140,N_6206);
xor U9163 (N_9163,N_5930,N_7206);
nand U9164 (N_9164,N_5308,N_7021);
and U9165 (N_9165,N_5049,N_6648);
or U9166 (N_9166,N_5309,N_5821);
or U9167 (N_9167,N_5048,N_5156);
or U9168 (N_9168,N_5451,N_5275);
or U9169 (N_9169,N_6216,N_5447);
and U9170 (N_9170,N_7234,N_5263);
or U9171 (N_9171,N_6541,N_7397);
xnor U9172 (N_9172,N_5753,N_5358);
or U9173 (N_9173,N_7428,N_5230);
xnor U9174 (N_9174,N_6898,N_5124);
nor U9175 (N_9175,N_6169,N_5612);
or U9176 (N_9176,N_6177,N_5131);
nor U9177 (N_9177,N_6338,N_7045);
or U9178 (N_9178,N_5636,N_6591);
nor U9179 (N_9179,N_5934,N_5189);
and U9180 (N_9180,N_5776,N_5925);
nand U9181 (N_9181,N_6915,N_6024);
or U9182 (N_9182,N_5708,N_7238);
nand U9183 (N_9183,N_6466,N_7092);
nor U9184 (N_9184,N_5335,N_5476);
nor U9185 (N_9185,N_5823,N_6858);
or U9186 (N_9186,N_7006,N_6084);
xor U9187 (N_9187,N_5503,N_6974);
and U9188 (N_9188,N_5416,N_6785);
nand U9189 (N_9189,N_6084,N_5120);
nand U9190 (N_9190,N_5894,N_5696);
xnor U9191 (N_9191,N_5287,N_7310);
or U9192 (N_9192,N_5483,N_7296);
and U9193 (N_9193,N_6294,N_7212);
nand U9194 (N_9194,N_7206,N_7009);
nand U9195 (N_9195,N_5102,N_6276);
or U9196 (N_9196,N_6611,N_5729);
nor U9197 (N_9197,N_6271,N_5189);
nor U9198 (N_9198,N_7076,N_7099);
xnor U9199 (N_9199,N_6421,N_6717);
and U9200 (N_9200,N_7310,N_5812);
and U9201 (N_9201,N_5506,N_5353);
and U9202 (N_9202,N_7199,N_6899);
nand U9203 (N_9203,N_6879,N_5092);
nand U9204 (N_9204,N_7265,N_7337);
nand U9205 (N_9205,N_7019,N_5970);
nand U9206 (N_9206,N_6825,N_6412);
xor U9207 (N_9207,N_6117,N_6880);
or U9208 (N_9208,N_6458,N_6052);
and U9209 (N_9209,N_7061,N_6937);
nand U9210 (N_9210,N_6058,N_7415);
and U9211 (N_9211,N_6178,N_7384);
and U9212 (N_9212,N_5033,N_5314);
nor U9213 (N_9213,N_5956,N_5411);
nor U9214 (N_9214,N_6384,N_5951);
xnor U9215 (N_9215,N_6565,N_6874);
xnor U9216 (N_9216,N_5174,N_5758);
xnor U9217 (N_9217,N_5084,N_7402);
and U9218 (N_9218,N_6063,N_7165);
xor U9219 (N_9219,N_7209,N_5417);
nor U9220 (N_9220,N_7468,N_5937);
xor U9221 (N_9221,N_5711,N_6104);
nand U9222 (N_9222,N_6314,N_7090);
or U9223 (N_9223,N_6944,N_7285);
xnor U9224 (N_9224,N_5789,N_5192);
or U9225 (N_9225,N_6851,N_5903);
nor U9226 (N_9226,N_7416,N_5812);
xor U9227 (N_9227,N_7001,N_6115);
xnor U9228 (N_9228,N_5139,N_5143);
and U9229 (N_9229,N_5739,N_6827);
nand U9230 (N_9230,N_5307,N_5308);
nand U9231 (N_9231,N_6400,N_5084);
and U9232 (N_9232,N_6163,N_6449);
or U9233 (N_9233,N_7478,N_7159);
and U9234 (N_9234,N_6534,N_5330);
xor U9235 (N_9235,N_7053,N_6841);
nand U9236 (N_9236,N_5372,N_7112);
nor U9237 (N_9237,N_6144,N_5739);
xor U9238 (N_9238,N_7461,N_7271);
or U9239 (N_9239,N_7361,N_5389);
or U9240 (N_9240,N_6926,N_6551);
nor U9241 (N_9241,N_6993,N_6489);
and U9242 (N_9242,N_5424,N_6653);
nor U9243 (N_9243,N_7065,N_5400);
nor U9244 (N_9244,N_5189,N_7176);
nor U9245 (N_9245,N_6565,N_5377);
nor U9246 (N_9246,N_6282,N_5517);
xor U9247 (N_9247,N_5989,N_6302);
and U9248 (N_9248,N_5431,N_5209);
nand U9249 (N_9249,N_6212,N_5917);
nand U9250 (N_9250,N_6710,N_5081);
xor U9251 (N_9251,N_7118,N_5149);
or U9252 (N_9252,N_6683,N_6503);
or U9253 (N_9253,N_5076,N_5469);
xnor U9254 (N_9254,N_6416,N_7465);
xnor U9255 (N_9255,N_7226,N_5965);
nor U9256 (N_9256,N_7346,N_7373);
or U9257 (N_9257,N_5803,N_5330);
and U9258 (N_9258,N_6951,N_6301);
or U9259 (N_9259,N_5542,N_7089);
xor U9260 (N_9260,N_6582,N_5149);
nor U9261 (N_9261,N_6808,N_5830);
or U9262 (N_9262,N_6319,N_6320);
xor U9263 (N_9263,N_7158,N_6569);
nand U9264 (N_9264,N_7286,N_7129);
nand U9265 (N_9265,N_5679,N_6160);
nand U9266 (N_9266,N_6702,N_5722);
or U9267 (N_9267,N_5692,N_6993);
nor U9268 (N_9268,N_7272,N_6822);
nor U9269 (N_9269,N_5709,N_5672);
xnor U9270 (N_9270,N_6996,N_7231);
xnor U9271 (N_9271,N_6701,N_7077);
or U9272 (N_9272,N_7437,N_7084);
and U9273 (N_9273,N_6431,N_6637);
xnor U9274 (N_9274,N_6381,N_5114);
and U9275 (N_9275,N_6271,N_7480);
nor U9276 (N_9276,N_5551,N_5850);
nor U9277 (N_9277,N_6197,N_6668);
nor U9278 (N_9278,N_6758,N_7220);
nand U9279 (N_9279,N_6423,N_5303);
and U9280 (N_9280,N_6001,N_5953);
xnor U9281 (N_9281,N_6597,N_7002);
nor U9282 (N_9282,N_5043,N_5052);
xor U9283 (N_9283,N_7394,N_5555);
and U9284 (N_9284,N_7316,N_5561);
xor U9285 (N_9285,N_6108,N_5968);
or U9286 (N_9286,N_6309,N_7195);
xnor U9287 (N_9287,N_5923,N_7013);
or U9288 (N_9288,N_5998,N_7399);
and U9289 (N_9289,N_5180,N_6254);
nand U9290 (N_9290,N_6795,N_5226);
nor U9291 (N_9291,N_7308,N_7159);
or U9292 (N_9292,N_5158,N_6913);
xnor U9293 (N_9293,N_5031,N_5561);
or U9294 (N_9294,N_5353,N_7068);
or U9295 (N_9295,N_5253,N_6992);
and U9296 (N_9296,N_5321,N_5762);
or U9297 (N_9297,N_6133,N_5290);
xnor U9298 (N_9298,N_5380,N_6207);
nor U9299 (N_9299,N_6760,N_6608);
or U9300 (N_9300,N_5865,N_7173);
nor U9301 (N_9301,N_7299,N_5350);
or U9302 (N_9302,N_5789,N_6057);
xnor U9303 (N_9303,N_5299,N_6918);
nor U9304 (N_9304,N_6194,N_5157);
or U9305 (N_9305,N_7047,N_5740);
xnor U9306 (N_9306,N_6825,N_6056);
and U9307 (N_9307,N_6015,N_7134);
or U9308 (N_9308,N_6179,N_5774);
and U9309 (N_9309,N_7064,N_5948);
and U9310 (N_9310,N_6648,N_6022);
nand U9311 (N_9311,N_6055,N_6441);
xnor U9312 (N_9312,N_7238,N_7219);
xnor U9313 (N_9313,N_7370,N_5273);
or U9314 (N_9314,N_5044,N_5851);
xnor U9315 (N_9315,N_6160,N_7163);
nand U9316 (N_9316,N_6611,N_6880);
or U9317 (N_9317,N_5639,N_5916);
nand U9318 (N_9318,N_7136,N_5682);
xnor U9319 (N_9319,N_6643,N_5434);
or U9320 (N_9320,N_6033,N_6104);
nor U9321 (N_9321,N_6237,N_6146);
nor U9322 (N_9322,N_6663,N_5498);
nand U9323 (N_9323,N_6934,N_7156);
xor U9324 (N_9324,N_5875,N_6114);
nor U9325 (N_9325,N_5132,N_5991);
nand U9326 (N_9326,N_6279,N_6264);
or U9327 (N_9327,N_5660,N_5045);
nand U9328 (N_9328,N_5397,N_5279);
and U9329 (N_9329,N_7491,N_5523);
nor U9330 (N_9330,N_7495,N_6718);
xnor U9331 (N_9331,N_6953,N_6720);
and U9332 (N_9332,N_6600,N_5466);
or U9333 (N_9333,N_5940,N_7002);
nand U9334 (N_9334,N_5585,N_6351);
nand U9335 (N_9335,N_5273,N_7182);
or U9336 (N_9336,N_7378,N_5312);
and U9337 (N_9337,N_5147,N_5411);
or U9338 (N_9338,N_5769,N_7226);
or U9339 (N_9339,N_6200,N_6415);
or U9340 (N_9340,N_6349,N_5922);
xor U9341 (N_9341,N_6744,N_6516);
and U9342 (N_9342,N_6921,N_7426);
and U9343 (N_9343,N_6021,N_5537);
or U9344 (N_9344,N_5776,N_6394);
xor U9345 (N_9345,N_5977,N_6319);
nand U9346 (N_9346,N_6253,N_5537);
nor U9347 (N_9347,N_6183,N_6071);
and U9348 (N_9348,N_7011,N_6227);
or U9349 (N_9349,N_7451,N_5313);
or U9350 (N_9350,N_7418,N_6240);
or U9351 (N_9351,N_5272,N_7192);
xor U9352 (N_9352,N_6438,N_6854);
or U9353 (N_9353,N_5279,N_6699);
xnor U9354 (N_9354,N_5921,N_6553);
xnor U9355 (N_9355,N_6262,N_6348);
nor U9356 (N_9356,N_7372,N_5638);
xor U9357 (N_9357,N_6474,N_6831);
nand U9358 (N_9358,N_5372,N_5743);
nor U9359 (N_9359,N_5447,N_5363);
nand U9360 (N_9360,N_5039,N_6897);
or U9361 (N_9361,N_6820,N_5118);
nand U9362 (N_9362,N_5075,N_6971);
nor U9363 (N_9363,N_6469,N_5693);
xnor U9364 (N_9364,N_5650,N_7210);
or U9365 (N_9365,N_6871,N_5619);
or U9366 (N_9366,N_6270,N_6878);
xor U9367 (N_9367,N_7196,N_6569);
xor U9368 (N_9368,N_7323,N_5581);
and U9369 (N_9369,N_7255,N_7239);
nor U9370 (N_9370,N_6701,N_7078);
nor U9371 (N_9371,N_5692,N_6382);
nand U9372 (N_9372,N_5126,N_6024);
and U9373 (N_9373,N_5361,N_6721);
or U9374 (N_9374,N_5633,N_6890);
or U9375 (N_9375,N_6072,N_6655);
and U9376 (N_9376,N_6931,N_5629);
or U9377 (N_9377,N_6821,N_5954);
nor U9378 (N_9378,N_6395,N_5839);
nand U9379 (N_9379,N_5359,N_5177);
nor U9380 (N_9380,N_6357,N_6557);
xnor U9381 (N_9381,N_6746,N_6787);
nor U9382 (N_9382,N_6009,N_7215);
or U9383 (N_9383,N_7040,N_6285);
xnor U9384 (N_9384,N_6348,N_5614);
or U9385 (N_9385,N_5477,N_5382);
xor U9386 (N_9386,N_5326,N_6631);
nand U9387 (N_9387,N_5984,N_6878);
and U9388 (N_9388,N_7458,N_6426);
nor U9389 (N_9389,N_5509,N_6326);
nor U9390 (N_9390,N_5457,N_5987);
nor U9391 (N_9391,N_5124,N_6752);
nor U9392 (N_9392,N_6295,N_6894);
nor U9393 (N_9393,N_6323,N_6893);
xor U9394 (N_9394,N_7095,N_7022);
and U9395 (N_9395,N_5808,N_5434);
or U9396 (N_9396,N_7461,N_6579);
or U9397 (N_9397,N_6967,N_6553);
xor U9398 (N_9398,N_6527,N_5776);
or U9399 (N_9399,N_5153,N_6955);
xnor U9400 (N_9400,N_6580,N_5510);
nor U9401 (N_9401,N_7233,N_5180);
and U9402 (N_9402,N_5924,N_6827);
and U9403 (N_9403,N_6324,N_5430);
nand U9404 (N_9404,N_5273,N_5030);
xor U9405 (N_9405,N_6351,N_5980);
xnor U9406 (N_9406,N_5358,N_7319);
xnor U9407 (N_9407,N_6285,N_5159);
and U9408 (N_9408,N_7151,N_6491);
or U9409 (N_9409,N_5286,N_5064);
nor U9410 (N_9410,N_5119,N_7431);
and U9411 (N_9411,N_5369,N_7496);
nor U9412 (N_9412,N_5602,N_5622);
or U9413 (N_9413,N_6312,N_5396);
xnor U9414 (N_9414,N_7190,N_6041);
nor U9415 (N_9415,N_7217,N_5331);
nor U9416 (N_9416,N_5283,N_6738);
nor U9417 (N_9417,N_5904,N_5579);
nand U9418 (N_9418,N_5702,N_5893);
xor U9419 (N_9419,N_5057,N_7202);
or U9420 (N_9420,N_6960,N_6209);
nand U9421 (N_9421,N_5115,N_6009);
xnor U9422 (N_9422,N_6352,N_7025);
xor U9423 (N_9423,N_6219,N_7476);
and U9424 (N_9424,N_6304,N_6490);
nor U9425 (N_9425,N_7339,N_7252);
xnor U9426 (N_9426,N_6246,N_7193);
nor U9427 (N_9427,N_5630,N_6557);
or U9428 (N_9428,N_5678,N_6550);
and U9429 (N_9429,N_6183,N_6399);
or U9430 (N_9430,N_7413,N_5151);
and U9431 (N_9431,N_5746,N_5447);
or U9432 (N_9432,N_7182,N_6407);
or U9433 (N_9433,N_6210,N_5969);
nand U9434 (N_9434,N_5350,N_5311);
nor U9435 (N_9435,N_7078,N_6859);
and U9436 (N_9436,N_7005,N_5969);
nand U9437 (N_9437,N_5320,N_6075);
nor U9438 (N_9438,N_6897,N_5600);
and U9439 (N_9439,N_5698,N_5031);
or U9440 (N_9440,N_6955,N_6051);
and U9441 (N_9441,N_5452,N_5036);
or U9442 (N_9442,N_6113,N_6593);
nor U9443 (N_9443,N_7251,N_5048);
and U9444 (N_9444,N_7173,N_6284);
nor U9445 (N_9445,N_6749,N_6569);
and U9446 (N_9446,N_6934,N_5115);
or U9447 (N_9447,N_6218,N_5778);
and U9448 (N_9448,N_6924,N_7149);
and U9449 (N_9449,N_5239,N_6069);
xnor U9450 (N_9450,N_6466,N_6076);
or U9451 (N_9451,N_6337,N_6999);
nand U9452 (N_9452,N_7012,N_6867);
and U9453 (N_9453,N_6687,N_5743);
or U9454 (N_9454,N_6756,N_5391);
nand U9455 (N_9455,N_6858,N_5357);
xnor U9456 (N_9456,N_5613,N_6249);
nor U9457 (N_9457,N_6886,N_7198);
nand U9458 (N_9458,N_7358,N_7448);
and U9459 (N_9459,N_5824,N_6681);
nand U9460 (N_9460,N_5747,N_5090);
nor U9461 (N_9461,N_5690,N_5045);
nor U9462 (N_9462,N_7174,N_7094);
nand U9463 (N_9463,N_5922,N_6710);
and U9464 (N_9464,N_6538,N_7314);
or U9465 (N_9465,N_6090,N_6776);
and U9466 (N_9466,N_5600,N_6457);
nor U9467 (N_9467,N_6626,N_5239);
or U9468 (N_9468,N_6405,N_6933);
or U9469 (N_9469,N_6047,N_5507);
or U9470 (N_9470,N_6883,N_7176);
nor U9471 (N_9471,N_5675,N_5700);
xnor U9472 (N_9472,N_5705,N_5865);
and U9473 (N_9473,N_5557,N_6014);
or U9474 (N_9474,N_6419,N_7121);
and U9475 (N_9475,N_7208,N_5267);
xor U9476 (N_9476,N_6570,N_5140);
xnor U9477 (N_9477,N_5432,N_6075);
or U9478 (N_9478,N_5828,N_5979);
nand U9479 (N_9479,N_5881,N_6517);
xnor U9480 (N_9480,N_6203,N_7279);
or U9481 (N_9481,N_6511,N_6286);
and U9482 (N_9482,N_5129,N_6400);
or U9483 (N_9483,N_6478,N_6916);
and U9484 (N_9484,N_7011,N_5739);
nor U9485 (N_9485,N_6522,N_5870);
xor U9486 (N_9486,N_7288,N_6965);
xnor U9487 (N_9487,N_6538,N_5155);
nand U9488 (N_9488,N_6016,N_7212);
nand U9489 (N_9489,N_6752,N_6464);
and U9490 (N_9490,N_5662,N_7300);
nor U9491 (N_9491,N_6495,N_6740);
nor U9492 (N_9492,N_5120,N_6386);
or U9493 (N_9493,N_7224,N_6387);
or U9494 (N_9494,N_5939,N_6059);
and U9495 (N_9495,N_5479,N_6870);
nand U9496 (N_9496,N_7408,N_6551);
xnor U9497 (N_9497,N_6671,N_7220);
or U9498 (N_9498,N_5606,N_6539);
or U9499 (N_9499,N_5251,N_7169);
nand U9500 (N_9500,N_5891,N_6891);
nor U9501 (N_9501,N_5691,N_6246);
xnor U9502 (N_9502,N_6753,N_6686);
nand U9503 (N_9503,N_6303,N_7317);
nor U9504 (N_9504,N_5445,N_7219);
and U9505 (N_9505,N_5582,N_5881);
xnor U9506 (N_9506,N_6771,N_5690);
and U9507 (N_9507,N_6708,N_6144);
or U9508 (N_9508,N_7490,N_6652);
and U9509 (N_9509,N_5584,N_6894);
nand U9510 (N_9510,N_6594,N_5107);
nand U9511 (N_9511,N_5729,N_6700);
and U9512 (N_9512,N_7250,N_7144);
and U9513 (N_9513,N_6159,N_6333);
nand U9514 (N_9514,N_6914,N_5681);
nor U9515 (N_9515,N_5049,N_5636);
nor U9516 (N_9516,N_5414,N_5901);
xnor U9517 (N_9517,N_6735,N_6400);
and U9518 (N_9518,N_5082,N_6612);
or U9519 (N_9519,N_5810,N_7332);
or U9520 (N_9520,N_6927,N_7209);
nand U9521 (N_9521,N_6218,N_5531);
and U9522 (N_9522,N_7083,N_7200);
nor U9523 (N_9523,N_7411,N_6266);
or U9524 (N_9524,N_5822,N_7165);
or U9525 (N_9525,N_7356,N_6753);
nand U9526 (N_9526,N_6913,N_5229);
or U9527 (N_9527,N_6660,N_7166);
nand U9528 (N_9528,N_5918,N_5891);
nor U9529 (N_9529,N_5228,N_7202);
xnor U9530 (N_9530,N_5635,N_5845);
and U9531 (N_9531,N_6058,N_5130);
and U9532 (N_9532,N_7109,N_5804);
nor U9533 (N_9533,N_7037,N_6896);
or U9534 (N_9534,N_6320,N_5130);
nor U9535 (N_9535,N_6250,N_6283);
nor U9536 (N_9536,N_5582,N_5923);
xnor U9537 (N_9537,N_7280,N_5965);
nand U9538 (N_9538,N_6647,N_6897);
nand U9539 (N_9539,N_6018,N_5087);
nand U9540 (N_9540,N_7160,N_5757);
or U9541 (N_9541,N_6358,N_5222);
or U9542 (N_9542,N_6268,N_5356);
or U9543 (N_9543,N_5241,N_6319);
nand U9544 (N_9544,N_5982,N_5191);
or U9545 (N_9545,N_6113,N_5091);
or U9546 (N_9546,N_6380,N_7363);
xnor U9547 (N_9547,N_6808,N_6946);
or U9548 (N_9548,N_7397,N_7355);
and U9549 (N_9549,N_6561,N_6369);
nand U9550 (N_9550,N_5820,N_5362);
xnor U9551 (N_9551,N_7150,N_6368);
nor U9552 (N_9552,N_5889,N_6087);
nand U9553 (N_9553,N_6739,N_7343);
and U9554 (N_9554,N_6073,N_5799);
or U9555 (N_9555,N_6678,N_5181);
or U9556 (N_9556,N_6635,N_6803);
or U9557 (N_9557,N_5672,N_7163);
nor U9558 (N_9558,N_5726,N_5449);
nand U9559 (N_9559,N_7484,N_6573);
and U9560 (N_9560,N_5003,N_6240);
and U9561 (N_9561,N_6683,N_5992);
xor U9562 (N_9562,N_6805,N_5483);
and U9563 (N_9563,N_5902,N_5605);
nand U9564 (N_9564,N_5972,N_6621);
or U9565 (N_9565,N_6269,N_7171);
nor U9566 (N_9566,N_5780,N_6565);
nor U9567 (N_9567,N_7452,N_7347);
or U9568 (N_9568,N_6851,N_5905);
or U9569 (N_9569,N_6423,N_5708);
and U9570 (N_9570,N_7110,N_6731);
nor U9571 (N_9571,N_5725,N_7056);
or U9572 (N_9572,N_7446,N_6550);
and U9573 (N_9573,N_6220,N_5509);
nand U9574 (N_9574,N_6955,N_5213);
xor U9575 (N_9575,N_6360,N_5424);
nor U9576 (N_9576,N_5057,N_6029);
nand U9577 (N_9577,N_7265,N_5909);
xnor U9578 (N_9578,N_5733,N_6453);
or U9579 (N_9579,N_5071,N_5562);
and U9580 (N_9580,N_7319,N_6703);
and U9581 (N_9581,N_5020,N_6303);
nand U9582 (N_9582,N_6734,N_6203);
xnor U9583 (N_9583,N_7456,N_6414);
nor U9584 (N_9584,N_7328,N_5967);
nor U9585 (N_9585,N_5180,N_6931);
xnor U9586 (N_9586,N_6632,N_5434);
and U9587 (N_9587,N_5624,N_6146);
nand U9588 (N_9588,N_6664,N_6628);
nand U9589 (N_9589,N_6894,N_6663);
or U9590 (N_9590,N_6205,N_6290);
nand U9591 (N_9591,N_5037,N_6986);
nand U9592 (N_9592,N_7415,N_7243);
nand U9593 (N_9593,N_5981,N_6244);
nand U9594 (N_9594,N_6291,N_6477);
xor U9595 (N_9595,N_5662,N_5177);
nand U9596 (N_9596,N_7488,N_5164);
nand U9597 (N_9597,N_5103,N_5853);
or U9598 (N_9598,N_6746,N_6847);
nor U9599 (N_9599,N_5955,N_6930);
nor U9600 (N_9600,N_5014,N_5226);
or U9601 (N_9601,N_6226,N_5634);
and U9602 (N_9602,N_6052,N_5494);
nor U9603 (N_9603,N_7028,N_7103);
or U9604 (N_9604,N_6041,N_6681);
xor U9605 (N_9605,N_5246,N_6469);
xnor U9606 (N_9606,N_7329,N_7409);
or U9607 (N_9607,N_7039,N_5740);
and U9608 (N_9608,N_6318,N_6422);
and U9609 (N_9609,N_6055,N_5434);
and U9610 (N_9610,N_6725,N_5606);
and U9611 (N_9611,N_5641,N_7195);
xnor U9612 (N_9612,N_7082,N_5959);
xnor U9613 (N_9613,N_5886,N_5357);
xor U9614 (N_9614,N_7344,N_6686);
and U9615 (N_9615,N_5948,N_6032);
nor U9616 (N_9616,N_5120,N_5678);
or U9617 (N_9617,N_7112,N_5938);
xnor U9618 (N_9618,N_5013,N_6818);
and U9619 (N_9619,N_6380,N_6578);
and U9620 (N_9620,N_6114,N_6523);
and U9621 (N_9621,N_5833,N_5974);
and U9622 (N_9622,N_5826,N_6018);
or U9623 (N_9623,N_5765,N_6549);
xnor U9624 (N_9624,N_6413,N_6411);
xnor U9625 (N_9625,N_6508,N_7269);
nand U9626 (N_9626,N_5187,N_5592);
or U9627 (N_9627,N_5609,N_5220);
xor U9628 (N_9628,N_6411,N_5891);
nor U9629 (N_9629,N_5866,N_5857);
or U9630 (N_9630,N_5902,N_5223);
nor U9631 (N_9631,N_5810,N_5045);
or U9632 (N_9632,N_7342,N_6664);
xnor U9633 (N_9633,N_6806,N_6988);
or U9634 (N_9634,N_7475,N_6960);
or U9635 (N_9635,N_6047,N_5922);
xor U9636 (N_9636,N_6745,N_5267);
and U9637 (N_9637,N_5615,N_6921);
and U9638 (N_9638,N_6291,N_6842);
nor U9639 (N_9639,N_5601,N_5626);
nor U9640 (N_9640,N_5710,N_5828);
xor U9641 (N_9641,N_6401,N_5093);
nor U9642 (N_9642,N_6605,N_5153);
and U9643 (N_9643,N_5188,N_6755);
nand U9644 (N_9644,N_5919,N_7291);
xnor U9645 (N_9645,N_7277,N_6931);
and U9646 (N_9646,N_5393,N_7324);
nor U9647 (N_9647,N_6551,N_7440);
and U9648 (N_9648,N_7490,N_6702);
nand U9649 (N_9649,N_7003,N_6078);
nor U9650 (N_9650,N_7367,N_7107);
and U9651 (N_9651,N_7117,N_6119);
nor U9652 (N_9652,N_6844,N_6430);
or U9653 (N_9653,N_5588,N_7465);
or U9654 (N_9654,N_5156,N_6329);
xnor U9655 (N_9655,N_5768,N_6404);
or U9656 (N_9656,N_5752,N_7270);
or U9657 (N_9657,N_5157,N_6484);
or U9658 (N_9658,N_5936,N_7465);
nand U9659 (N_9659,N_6378,N_5166);
and U9660 (N_9660,N_6261,N_5414);
nor U9661 (N_9661,N_6302,N_5050);
nor U9662 (N_9662,N_5727,N_6318);
xor U9663 (N_9663,N_5941,N_5747);
or U9664 (N_9664,N_6400,N_5462);
xnor U9665 (N_9665,N_5937,N_5022);
nor U9666 (N_9666,N_6851,N_5241);
and U9667 (N_9667,N_7088,N_7224);
xor U9668 (N_9668,N_6025,N_5137);
and U9669 (N_9669,N_6122,N_6753);
nand U9670 (N_9670,N_7131,N_6276);
or U9671 (N_9671,N_7205,N_7062);
nor U9672 (N_9672,N_6774,N_6848);
nand U9673 (N_9673,N_7038,N_6576);
or U9674 (N_9674,N_5077,N_7379);
nor U9675 (N_9675,N_5763,N_6011);
nor U9676 (N_9676,N_6594,N_7144);
xnor U9677 (N_9677,N_6744,N_5336);
xor U9678 (N_9678,N_7265,N_5814);
nor U9679 (N_9679,N_5049,N_5418);
or U9680 (N_9680,N_6701,N_6938);
nor U9681 (N_9681,N_5868,N_5499);
xor U9682 (N_9682,N_6139,N_5870);
nand U9683 (N_9683,N_6653,N_5102);
nand U9684 (N_9684,N_7019,N_6983);
and U9685 (N_9685,N_7170,N_6473);
and U9686 (N_9686,N_5458,N_6610);
xor U9687 (N_9687,N_7435,N_5027);
nand U9688 (N_9688,N_6632,N_7094);
nor U9689 (N_9689,N_7494,N_6846);
nor U9690 (N_9690,N_6843,N_7479);
or U9691 (N_9691,N_6381,N_5491);
or U9692 (N_9692,N_7022,N_6268);
xor U9693 (N_9693,N_6347,N_5888);
xor U9694 (N_9694,N_5869,N_5241);
nor U9695 (N_9695,N_6375,N_5586);
or U9696 (N_9696,N_5099,N_5337);
nor U9697 (N_9697,N_6377,N_6071);
nand U9698 (N_9698,N_7397,N_6481);
nor U9699 (N_9699,N_6457,N_5893);
or U9700 (N_9700,N_7015,N_5278);
or U9701 (N_9701,N_6791,N_6100);
nand U9702 (N_9702,N_6487,N_5112);
nand U9703 (N_9703,N_7130,N_5747);
or U9704 (N_9704,N_7248,N_5958);
xor U9705 (N_9705,N_6861,N_7196);
nand U9706 (N_9706,N_6201,N_6667);
or U9707 (N_9707,N_5974,N_7020);
nor U9708 (N_9708,N_5400,N_5682);
nor U9709 (N_9709,N_5527,N_6392);
nand U9710 (N_9710,N_7210,N_6291);
nand U9711 (N_9711,N_6529,N_6227);
and U9712 (N_9712,N_7465,N_6252);
nor U9713 (N_9713,N_5318,N_5498);
nand U9714 (N_9714,N_7398,N_5628);
or U9715 (N_9715,N_6221,N_5654);
nor U9716 (N_9716,N_5640,N_7102);
and U9717 (N_9717,N_7499,N_5501);
and U9718 (N_9718,N_5888,N_5000);
or U9719 (N_9719,N_7415,N_5762);
xnor U9720 (N_9720,N_6124,N_6838);
or U9721 (N_9721,N_6366,N_6860);
nand U9722 (N_9722,N_7226,N_6549);
nand U9723 (N_9723,N_5340,N_5709);
and U9724 (N_9724,N_5132,N_5369);
nand U9725 (N_9725,N_7032,N_5854);
or U9726 (N_9726,N_6676,N_5173);
and U9727 (N_9727,N_5068,N_6623);
nand U9728 (N_9728,N_7493,N_6231);
nor U9729 (N_9729,N_5284,N_6827);
xor U9730 (N_9730,N_5361,N_6858);
and U9731 (N_9731,N_5032,N_5820);
or U9732 (N_9732,N_6200,N_5935);
xor U9733 (N_9733,N_7053,N_6933);
or U9734 (N_9734,N_7301,N_6436);
nor U9735 (N_9735,N_5999,N_5556);
nor U9736 (N_9736,N_5801,N_5359);
and U9737 (N_9737,N_5888,N_6385);
nand U9738 (N_9738,N_5609,N_5307);
or U9739 (N_9739,N_7390,N_5790);
nand U9740 (N_9740,N_6205,N_7419);
xor U9741 (N_9741,N_6164,N_5995);
nor U9742 (N_9742,N_7255,N_7198);
or U9743 (N_9743,N_6288,N_6687);
nand U9744 (N_9744,N_5802,N_7464);
xor U9745 (N_9745,N_6229,N_5658);
or U9746 (N_9746,N_7482,N_6100);
and U9747 (N_9747,N_6105,N_6623);
nor U9748 (N_9748,N_7361,N_6658);
or U9749 (N_9749,N_6312,N_6962);
or U9750 (N_9750,N_6581,N_5672);
nor U9751 (N_9751,N_7194,N_5798);
nor U9752 (N_9752,N_5276,N_5480);
or U9753 (N_9753,N_6953,N_6913);
or U9754 (N_9754,N_5214,N_7025);
nor U9755 (N_9755,N_5625,N_7081);
xor U9756 (N_9756,N_5165,N_7282);
and U9757 (N_9757,N_6071,N_6422);
nand U9758 (N_9758,N_6902,N_6806);
nor U9759 (N_9759,N_5369,N_6992);
or U9760 (N_9760,N_7108,N_6833);
xnor U9761 (N_9761,N_5735,N_7250);
nor U9762 (N_9762,N_6274,N_6947);
and U9763 (N_9763,N_5486,N_6715);
or U9764 (N_9764,N_5507,N_6420);
xnor U9765 (N_9765,N_5303,N_5107);
xnor U9766 (N_9766,N_5748,N_6456);
xnor U9767 (N_9767,N_6842,N_5573);
and U9768 (N_9768,N_5650,N_5353);
nor U9769 (N_9769,N_6649,N_6503);
xor U9770 (N_9770,N_5914,N_5514);
nand U9771 (N_9771,N_5710,N_6987);
xnor U9772 (N_9772,N_5194,N_5572);
xor U9773 (N_9773,N_5973,N_7404);
or U9774 (N_9774,N_5170,N_5065);
nor U9775 (N_9775,N_6638,N_7087);
nand U9776 (N_9776,N_6101,N_5830);
nand U9777 (N_9777,N_5989,N_5005);
nand U9778 (N_9778,N_7139,N_5837);
nand U9779 (N_9779,N_5447,N_6066);
and U9780 (N_9780,N_5286,N_5226);
or U9781 (N_9781,N_6608,N_5764);
nor U9782 (N_9782,N_7025,N_6184);
xnor U9783 (N_9783,N_6248,N_5798);
nor U9784 (N_9784,N_6835,N_5702);
or U9785 (N_9785,N_7127,N_6267);
or U9786 (N_9786,N_5994,N_6875);
nand U9787 (N_9787,N_5458,N_6135);
xnor U9788 (N_9788,N_6153,N_7331);
nand U9789 (N_9789,N_7198,N_5867);
xnor U9790 (N_9790,N_5995,N_7075);
and U9791 (N_9791,N_7393,N_5098);
xor U9792 (N_9792,N_5657,N_6774);
or U9793 (N_9793,N_5509,N_6781);
nand U9794 (N_9794,N_6427,N_6204);
nor U9795 (N_9795,N_5580,N_5239);
nor U9796 (N_9796,N_5332,N_6592);
nand U9797 (N_9797,N_5092,N_5367);
or U9798 (N_9798,N_6189,N_7298);
or U9799 (N_9799,N_7168,N_5832);
and U9800 (N_9800,N_6698,N_6745);
and U9801 (N_9801,N_5675,N_5349);
or U9802 (N_9802,N_5079,N_6856);
or U9803 (N_9803,N_5283,N_5203);
xnor U9804 (N_9804,N_5168,N_6034);
nor U9805 (N_9805,N_6493,N_5856);
nor U9806 (N_9806,N_7220,N_6113);
nor U9807 (N_9807,N_5873,N_6864);
nor U9808 (N_9808,N_5415,N_5144);
xnor U9809 (N_9809,N_6566,N_6256);
and U9810 (N_9810,N_5646,N_5335);
xor U9811 (N_9811,N_7128,N_6233);
and U9812 (N_9812,N_5925,N_6607);
or U9813 (N_9813,N_5461,N_6891);
and U9814 (N_9814,N_6460,N_7041);
xor U9815 (N_9815,N_5700,N_6387);
and U9816 (N_9816,N_7277,N_5167);
or U9817 (N_9817,N_6242,N_5039);
xnor U9818 (N_9818,N_6192,N_6816);
and U9819 (N_9819,N_6719,N_7498);
and U9820 (N_9820,N_5349,N_7156);
and U9821 (N_9821,N_6013,N_5883);
xor U9822 (N_9822,N_5970,N_6781);
nand U9823 (N_9823,N_5656,N_5869);
xor U9824 (N_9824,N_5137,N_6090);
nand U9825 (N_9825,N_5417,N_5765);
nand U9826 (N_9826,N_5443,N_6298);
nand U9827 (N_9827,N_7196,N_6690);
and U9828 (N_9828,N_7039,N_5843);
or U9829 (N_9829,N_6243,N_7070);
or U9830 (N_9830,N_5065,N_5002);
and U9831 (N_9831,N_7099,N_5996);
nand U9832 (N_9832,N_7473,N_6389);
nor U9833 (N_9833,N_6815,N_6378);
and U9834 (N_9834,N_5310,N_6263);
or U9835 (N_9835,N_5042,N_7058);
or U9836 (N_9836,N_6385,N_6068);
and U9837 (N_9837,N_6327,N_6894);
and U9838 (N_9838,N_6041,N_5402);
nand U9839 (N_9839,N_7077,N_6647);
or U9840 (N_9840,N_6953,N_5351);
or U9841 (N_9841,N_6620,N_5686);
nand U9842 (N_9842,N_7274,N_5061);
nand U9843 (N_9843,N_5273,N_5025);
nor U9844 (N_9844,N_5036,N_7225);
and U9845 (N_9845,N_6745,N_5220);
nand U9846 (N_9846,N_5142,N_6483);
nand U9847 (N_9847,N_5289,N_5688);
nor U9848 (N_9848,N_5390,N_6001);
or U9849 (N_9849,N_7132,N_5820);
xor U9850 (N_9850,N_5861,N_6363);
or U9851 (N_9851,N_5388,N_6790);
nand U9852 (N_9852,N_7151,N_6801);
or U9853 (N_9853,N_7359,N_5352);
xnor U9854 (N_9854,N_5802,N_5361);
and U9855 (N_9855,N_5984,N_5056);
xnor U9856 (N_9856,N_6950,N_5773);
or U9857 (N_9857,N_7012,N_5848);
and U9858 (N_9858,N_6333,N_5150);
and U9859 (N_9859,N_6533,N_6459);
xnor U9860 (N_9860,N_6982,N_5622);
nand U9861 (N_9861,N_7143,N_7172);
nor U9862 (N_9862,N_6242,N_5713);
nor U9863 (N_9863,N_6111,N_6666);
or U9864 (N_9864,N_6160,N_5062);
or U9865 (N_9865,N_7493,N_5688);
or U9866 (N_9866,N_6506,N_5390);
nor U9867 (N_9867,N_7373,N_5804);
nand U9868 (N_9868,N_7270,N_5234);
or U9869 (N_9869,N_5732,N_6955);
nor U9870 (N_9870,N_6353,N_6304);
and U9871 (N_9871,N_6926,N_6557);
nor U9872 (N_9872,N_6554,N_5193);
or U9873 (N_9873,N_5608,N_5023);
nor U9874 (N_9874,N_5108,N_7225);
or U9875 (N_9875,N_7290,N_5738);
or U9876 (N_9876,N_5385,N_7262);
and U9877 (N_9877,N_6762,N_5531);
nand U9878 (N_9878,N_5321,N_5033);
nand U9879 (N_9879,N_7270,N_6444);
and U9880 (N_9880,N_5229,N_6825);
or U9881 (N_9881,N_5842,N_7381);
xor U9882 (N_9882,N_6778,N_6956);
xnor U9883 (N_9883,N_7224,N_6686);
xnor U9884 (N_9884,N_5755,N_7393);
nor U9885 (N_9885,N_5240,N_5128);
nand U9886 (N_9886,N_6903,N_5335);
xor U9887 (N_9887,N_6138,N_6588);
or U9888 (N_9888,N_5965,N_5263);
xnor U9889 (N_9889,N_6770,N_5371);
nand U9890 (N_9890,N_5195,N_5112);
nand U9891 (N_9891,N_5824,N_6702);
and U9892 (N_9892,N_5167,N_5551);
or U9893 (N_9893,N_7465,N_5397);
xor U9894 (N_9894,N_5023,N_6779);
nor U9895 (N_9895,N_5690,N_6376);
or U9896 (N_9896,N_5801,N_5744);
and U9897 (N_9897,N_7327,N_6663);
xnor U9898 (N_9898,N_5361,N_6368);
xnor U9899 (N_9899,N_6506,N_5459);
or U9900 (N_9900,N_7309,N_6416);
nor U9901 (N_9901,N_6889,N_7238);
xor U9902 (N_9902,N_7057,N_5886);
nor U9903 (N_9903,N_6273,N_6589);
and U9904 (N_9904,N_5102,N_5492);
nor U9905 (N_9905,N_5213,N_5161);
and U9906 (N_9906,N_7260,N_7026);
nor U9907 (N_9907,N_7466,N_5812);
xor U9908 (N_9908,N_5268,N_5536);
or U9909 (N_9909,N_5629,N_6315);
nor U9910 (N_9910,N_5958,N_7384);
nand U9911 (N_9911,N_7128,N_5390);
nor U9912 (N_9912,N_7219,N_6561);
xnor U9913 (N_9913,N_6812,N_5280);
nor U9914 (N_9914,N_7191,N_6925);
nor U9915 (N_9915,N_6037,N_6236);
nand U9916 (N_9916,N_7380,N_5975);
or U9917 (N_9917,N_7357,N_6731);
and U9918 (N_9918,N_5943,N_5766);
nor U9919 (N_9919,N_6414,N_7309);
nand U9920 (N_9920,N_6723,N_7274);
or U9921 (N_9921,N_7457,N_5389);
or U9922 (N_9922,N_5137,N_5452);
and U9923 (N_9923,N_6924,N_6321);
xor U9924 (N_9924,N_5558,N_5872);
and U9925 (N_9925,N_6461,N_6033);
or U9926 (N_9926,N_6788,N_5001);
nand U9927 (N_9927,N_6372,N_5545);
nand U9928 (N_9928,N_6756,N_5452);
nand U9929 (N_9929,N_6964,N_6879);
or U9930 (N_9930,N_6995,N_6073);
xor U9931 (N_9931,N_6958,N_5564);
xor U9932 (N_9932,N_6521,N_5233);
or U9933 (N_9933,N_7345,N_6486);
or U9934 (N_9934,N_5799,N_5101);
and U9935 (N_9935,N_5364,N_5986);
nand U9936 (N_9936,N_5886,N_7107);
nand U9937 (N_9937,N_7417,N_5558);
xnor U9938 (N_9938,N_6517,N_5643);
nor U9939 (N_9939,N_6760,N_5727);
or U9940 (N_9940,N_5622,N_6062);
nand U9941 (N_9941,N_5642,N_6502);
or U9942 (N_9942,N_6280,N_5007);
and U9943 (N_9943,N_6654,N_7126);
and U9944 (N_9944,N_5182,N_5893);
or U9945 (N_9945,N_6638,N_7485);
nor U9946 (N_9946,N_5586,N_6000);
nor U9947 (N_9947,N_6596,N_6209);
nand U9948 (N_9948,N_5297,N_5598);
and U9949 (N_9949,N_6054,N_7206);
xnor U9950 (N_9950,N_6584,N_6177);
xor U9951 (N_9951,N_6411,N_5332);
and U9952 (N_9952,N_7126,N_6587);
nor U9953 (N_9953,N_5243,N_6772);
or U9954 (N_9954,N_6634,N_7480);
xnor U9955 (N_9955,N_6228,N_5876);
nand U9956 (N_9956,N_6256,N_7345);
nor U9957 (N_9957,N_7236,N_7026);
nand U9958 (N_9958,N_5018,N_5354);
nor U9959 (N_9959,N_5330,N_5725);
and U9960 (N_9960,N_5627,N_5595);
or U9961 (N_9961,N_5050,N_6650);
nor U9962 (N_9962,N_5675,N_7225);
xor U9963 (N_9963,N_6612,N_5268);
nor U9964 (N_9964,N_6518,N_5915);
or U9965 (N_9965,N_5135,N_7033);
nor U9966 (N_9966,N_5711,N_5501);
xor U9967 (N_9967,N_7371,N_6566);
nand U9968 (N_9968,N_6590,N_5112);
and U9969 (N_9969,N_5423,N_7127);
nor U9970 (N_9970,N_5894,N_5091);
or U9971 (N_9971,N_5762,N_5004);
or U9972 (N_9972,N_6866,N_5234);
or U9973 (N_9973,N_5370,N_6895);
or U9974 (N_9974,N_6667,N_5616);
nor U9975 (N_9975,N_5254,N_6018);
nor U9976 (N_9976,N_5237,N_6088);
xor U9977 (N_9977,N_6641,N_6717);
and U9978 (N_9978,N_6376,N_6889);
or U9979 (N_9979,N_6886,N_7437);
or U9980 (N_9980,N_5640,N_6004);
xor U9981 (N_9981,N_5655,N_5190);
nand U9982 (N_9982,N_5815,N_5960);
nor U9983 (N_9983,N_5745,N_5187);
xnor U9984 (N_9984,N_5570,N_6538);
or U9985 (N_9985,N_5361,N_6201);
nand U9986 (N_9986,N_6585,N_6213);
or U9987 (N_9987,N_6644,N_5359);
xor U9988 (N_9988,N_5511,N_6166);
or U9989 (N_9989,N_6119,N_6330);
xor U9990 (N_9990,N_7054,N_6122);
and U9991 (N_9991,N_7142,N_5475);
nand U9992 (N_9992,N_5572,N_5573);
and U9993 (N_9993,N_7138,N_6269);
and U9994 (N_9994,N_7376,N_7472);
and U9995 (N_9995,N_5178,N_5652);
nand U9996 (N_9996,N_7378,N_7163);
nand U9997 (N_9997,N_5483,N_6067);
or U9998 (N_9998,N_7301,N_6742);
and U9999 (N_9999,N_7416,N_6850);
nor UO_0 (O_0,N_7531,N_8410);
nor UO_1 (O_1,N_9600,N_8532);
nor UO_2 (O_2,N_8567,N_9057);
and UO_3 (O_3,N_8165,N_7807);
or UO_4 (O_4,N_8407,N_8266);
and UO_5 (O_5,N_9851,N_7950);
and UO_6 (O_6,N_9116,N_9718);
nor UO_7 (O_7,N_8578,N_8894);
and UO_8 (O_8,N_7551,N_8088);
nand UO_9 (O_9,N_8649,N_8505);
nand UO_10 (O_10,N_9836,N_8246);
nor UO_11 (O_11,N_9816,N_8178);
xnor UO_12 (O_12,N_9393,N_9170);
and UO_13 (O_13,N_8226,N_7841);
xor UO_14 (O_14,N_8106,N_8613);
nand UO_15 (O_15,N_8022,N_9192);
or UO_16 (O_16,N_8768,N_9987);
and UO_17 (O_17,N_8187,N_7568);
nand UO_18 (O_18,N_7720,N_8946);
nor UO_19 (O_19,N_7595,N_8597);
xnor UO_20 (O_20,N_7715,N_9276);
nor UO_21 (O_21,N_7828,N_9713);
nor UO_22 (O_22,N_8412,N_9859);
nand UO_23 (O_23,N_9082,N_7819);
nand UO_24 (O_24,N_9607,N_9847);
nor UO_25 (O_25,N_9819,N_7849);
xnor UO_26 (O_26,N_7528,N_7578);
or UO_27 (O_27,N_7876,N_9824);
or UO_28 (O_28,N_9783,N_9461);
xor UO_29 (O_29,N_9845,N_9390);
nor UO_30 (O_30,N_8205,N_9140);
nor UO_31 (O_31,N_9232,N_7729);
and UO_32 (O_32,N_8150,N_8896);
and UO_33 (O_33,N_7795,N_7530);
nand UO_34 (O_34,N_8814,N_9242);
nor UO_35 (O_35,N_7652,N_9490);
nand UO_36 (O_36,N_9411,N_7862);
xnor UO_37 (O_37,N_8213,N_8858);
xor UO_38 (O_38,N_8760,N_8541);
nand UO_39 (O_39,N_9483,N_9946);
nand UO_40 (O_40,N_8061,N_8604);
nand UO_41 (O_41,N_9820,N_7920);
nand UO_42 (O_42,N_9583,N_8902);
xnor UO_43 (O_43,N_8476,N_7627);
nand UO_44 (O_44,N_8718,N_9281);
xnor UO_45 (O_45,N_9703,N_8575);
nand UO_46 (O_46,N_8228,N_9065);
or UO_47 (O_47,N_8565,N_9273);
xor UO_48 (O_48,N_7509,N_8382);
nor UO_49 (O_49,N_8588,N_9993);
xnor UO_50 (O_50,N_8610,N_8669);
nand UO_51 (O_51,N_9710,N_8563);
xor UO_52 (O_52,N_8183,N_9727);
or UO_53 (O_53,N_7544,N_8711);
and UO_54 (O_54,N_8630,N_7585);
and UO_55 (O_55,N_9387,N_8839);
xor UO_56 (O_56,N_8821,N_9911);
or UO_57 (O_57,N_8800,N_9794);
nand UO_58 (O_58,N_8646,N_8314);
xor UO_59 (O_59,N_8693,N_8857);
and UO_60 (O_60,N_9489,N_8548);
nor UO_61 (O_61,N_8687,N_9077);
and UO_62 (O_62,N_9969,N_9491);
nand UO_63 (O_63,N_9428,N_8999);
and UO_64 (O_64,N_8891,N_8851);
nand UO_65 (O_65,N_9218,N_8437);
or UO_66 (O_66,N_9750,N_8348);
or UO_67 (O_67,N_8642,N_8663);
or UO_68 (O_68,N_9303,N_9451);
or UO_69 (O_69,N_9740,N_9267);
and UO_70 (O_70,N_9823,N_8932);
or UO_71 (O_71,N_9195,N_8392);
or UO_72 (O_72,N_8385,N_9472);
nor UO_73 (O_73,N_9834,N_9511);
or UO_74 (O_74,N_9257,N_7688);
and UO_75 (O_75,N_8511,N_7955);
or UO_76 (O_76,N_7889,N_8250);
nand UO_77 (O_77,N_9027,N_8121);
or UO_78 (O_78,N_7780,N_9655);
xnor UO_79 (O_79,N_8453,N_7655);
or UO_80 (O_80,N_8915,N_7882);
nor UO_81 (O_81,N_8301,N_9021);
and UO_82 (O_82,N_9869,N_8979);
xor UO_83 (O_83,N_8355,N_8728);
nor UO_84 (O_84,N_8370,N_8546);
and UO_85 (O_85,N_7691,N_7890);
nand UO_86 (O_86,N_7789,N_9348);
or UO_87 (O_87,N_8904,N_8601);
xor UO_88 (O_88,N_8201,N_7887);
and UO_89 (O_89,N_9403,N_8318);
nand UO_90 (O_90,N_8306,N_8787);
and UO_91 (O_91,N_8569,N_8340);
and UO_92 (O_92,N_7880,N_9376);
or UO_93 (O_93,N_8551,N_9687);
nor UO_94 (O_94,N_8115,N_8050);
and UO_95 (O_95,N_9357,N_9111);
or UO_96 (O_96,N_9646,N_9271);
nand UO_97 (O_97,N_7933,N_9494);
and UO_98 (O_98,N_9106,N_9593);
nor UO_99 (O_99,N_8162,N_9962);
nor UO_100 (O_100,N_9720,N_7705);
and UO_101 (O_101,N_7963,N_8184);
nand UO_102 (O_102,N_8124,N_7784);
nand UO_103 (O_103,N_8449,N_8985);
nor UO_104 (O_104,N_8369,N_8923);
nand UO_105 (O_105,N_9689,N_9066);
and UO_106 (O_106,N_8105,N_8239);
or UO_107 (O_107,N_8953,N_7860);
xor UO_108 (O_108,N_9323,N_8095);
nand UO_109 (O_109,N_9202,N_9531);
and UO_110 (O_110,N_8917,N_9807);
nand UO_111 (O_111,N_8867,N_9688);
nand UO_112 (O_112,N_7896,N_9258);
or UO_113 (O_113,N_9768,N_7523);
nand UO_114 (O_114,N_9180,N_8652);
nand UO_115 (O_115,N_7596,N_9322);
nor UO_116 (O_116,N_8496,N_8877);
nor UO_117 (O_117,N_8014,N_8018);
nand UO_118 (O_118,N_9132,N_7782);
nor UO_119 (O_119,N_8712,N_9282);
and UO_120 (O_120,N_8155,N_9592);
nor UO_121 (O_121,N_9810,N_8102);
nor UO_122 (O_122,N_9166,N_7559);
and UO_123 (O_123,N_9255,N_8114);
xnor UO_124 (O_124,N_9204,N_7952);
or UO_125 (O_125,N_9647,N_8905);
or UO_126 (O_126,N_9153,N_7805);
nor UO_127 (O_127,N_9216,N_8886);
xor UO_128 (O_128,N_8016,N_8174);
nor UO_129 (O_129,N_9105,N_9844);
or UO_130 (O_130,N_7659,N_7878);
or UO_131 (O_131,N_9006,N_8729);
and UO_132 (O_132,N_9838,N_8884);
and UO_133 (O_133,N_8328,N_7993);
xor UO_134 (O_134,N_9199,N_7796);
nand UO_135 (O_135,N_9039,N_8265);
nor UO_136 (O_136,N_9488,N_9527);
or UO_137 (O_137,N_8179,N_7811);
xor UO_138 (O_138,N_8745,N_8364);
and UO_139 (O_139,N_9220,N_8947);
and UO_140 (O_140,N_8817,N_7845);
or UO_141 (O_141,N_7972,N_9857);
nor UO_142 (O_142,N_8397,N_9389);
or UO_143 (O_143,N_9415,N_9030);
xor UO_144 (O_144,N_7614,N_9040);
xnor UO_145 (O_145,N_9585,N_7566);
nor UO_146 (O_146,N_8142,N_9353);
and UO_147 (O_147,N_7975,N_9943);
xor UO_148 (O_148,N_9044,N_8376);
nand UO_149 (O_149,N_9072,N_9509);
xnor UO_150 (O_150,N_9139,N_9289);
or UO_151 (O_151,N_8519,N_7689);
nand UO_152 (O_152,N_9564,N_9977);
or UO_153 (O_153,N_8697,N_7518);
nand UO_154 (O_154,N_8998,N_8277);
xor UO_155 (O_155,N_7765,N_7747);
and UO_156 (O_156,N_8076,N_9501);
nor UO_157 (O_157,N_8833,N_8607);
nand UO_158 (O_158,N_8835,N_9552);
or UO_159 (O_159,N_9539,N_9230);
or UO_160 (O_160,N_8522,N_9885);
xor UO_161 (O_161,N_8020,N_7730);
and UO_162 (O_162,N_8084,N_9274);
or UO_163 (O_163,N_9799,N_9115);
or UO_164 (O_164,N_7851,N_9961);
xor UO_165 (O_165,N_7554,N_9396);
nor UO_166 (O_166,N_8801,N_9723);
nor UO_167 (O_167,N_9528,N_9701);
and UO_168 (O_168,N_9705,N_9979);
xnor UO_169 (O_169,N_9645,N_8761);
and UO_170 (O_170,N_7776,N_9171);
and UO_171 (O_171,N_9515,N_9888);
nand UO_172 (O_172,N_8864,N_8900);
and UO_173 (O_173,N_9830,N_7918);
nor UO_174 (O_174,N_8918,N_8557);
xor UO_175 (O_175,N_7542,N_9413);
and UO_176 (O_176,N_8104,N_7623);
and UO_177 (O_177,N_8866,N_7884);
nand UO_178 (O_178,N_8276,N_8230);
xnor UO_179 (O_179,N_8543,N_9912);
and UO_180 (O_180,N_8815,N_9486);
nand UO_181 (O_181,N_8278,N_8117);
or UO_182 (O_182,N_8462,N_9404);
and UO_183 (O_183,N_7602,N_9938);
and UO_184 (O_184,N_8722,N_7501);
nor UO_185 (O_185,N_9133,N_8012);
or UO_186 (O_186,N_8176,N_8307);
nand UO_187 (O_187,N_9431,N_9638);
xor UO_188 (O_188,N_8868,N_7939);
or UO_189 (O_189,N_8000,N_9444);
or UO_190 (O_190,N_8427,N_7982);
nor UO_191 (O_191,N_9878,N_8171);
xnor UO_192 (O_192,N_8158,N_9758);
or UO_193 (O_193,N_9658,N_9037);
xor UO_194 (O_194,N_7822,N_9523);
and UO_195 (O_195,N_7543,N_9164);
nor UO_196 (O_196,N_8730,N_9866);
and UO_197 (O_197,N_9023,N_8691);
nor UO_198 (O_198,N_7583,N_9302);
xnor UO_199 (O_199,N_9317,N_8464);
nor UO_200 (O_200,N_9229,N_9391);
nor UO_201 (O_201,N_9529,N_8068);
nand UO_202 (O_202,N_8818,N_9328);
or UO_203 (O_203,N_7867,N_9695);
nand UO_204 (O_204,N_9620,N_9124);
nand UO_205 (O_205,N_7942,N_7500);
or UO_206 (O_206,N_9201,N_9679);
nor UO_207 (O_207,N_8043,N_9746);
nor UO_208 (O_208,N_9252,N_8190);
or UO_209 (O_209,N_8714,N_7708);
nor UO_210 (O_210,N_8680,N_8304);
xor UO_211 (O_211,N_9992,N_9045);
nor UO_212 (O_212,N_7970,N_8200);
xor UO_213 (O_213,N_8120,N_9575);
or UO_214 (O_214,N_8589,N_9112);
nand UO_215 (O_215,N_7863,N_8622);
xor UO_216 (O_216,N_8836,N_9015);
nor UO_217 (O_217,N_9541,N_7683);
nor UO_218 (O_218,N_9660,N_8220);
xor UO_219 (O_219,N_9898,N_8925);
or UO_220 (O_220,N_9612,N_9340);
nand UO_221 (O_221,N_7616,N_9475);
nor UO_222 (O_222,N_7662,N_8756);
nor UO_223 (O_223,N_8389,N_8152);
nor UO_224 (O_224,N_9492,N_8770);
and UO_225 (O_225,N_9563,N_9073);
and UO_226 (O_226,N_9706,N_8128);
and UO_227 (O_227,N_7928,N_8843);
or UO_228 (O_228,N_9361,N_8032);
nor UO_229 (O_229,N_9239,N_8353);
or UO_230 (O_230,N_9188,N_9137);
nor UO_231 (O_231,N_8963,N_9788);
nor UO_232 (O_232,N_7755,N_9381);
nor UO_233 (O_233,N_9756,N_7908);
and UO_234 (O_234,N_7599,N_9757);
or UO_235 (O_235,N_8677,N_9096);
xnor UO_236 (O_236,N_7612,N_8173);
or UO_237 (O_237,N_8252,N_8931);
nand UO_238 (O_238,N_7941,N_9359);
nand UO_239 (O_239,N_9837,N_9923);
nor UO_240 (O_240,N_8292,N_8309);
xnor UO_241 (O_241,N_8363,N_8500);
and UO_242 (O_242,N_8240,N_9372);
nor UO_243 (O_243,N_7816,N_9731);
and UO_244 (O_244,N_9903,N_7524);
nor UO_245 (O_245,N_9884,N_8447);
nand UO_246 (O_246,N_9558,N_7693);
or UO_247 (O_247,N_8542,N_7598);
and UO_248 (O_248,N_7858,N_9277);
xor UO_249 (O_249,N_9835,N_7638);
xnor UO_250 (O_250,N_8809,N_9010);
nor UO_251 (O_251,N_8899,N_8494);
or UO_252 (O_252,N_9925,N_9599);
xnor UO_253 (O_253,N_9036,N_9767);
nand UO_254 (O_254,N_9861,N_8862);
nor UO_255 (O_255,N_9468,N_8263);
nor UO_256 (O_256,N_9743,N_9297);
nor UO_257 (O_257,N_8566,N_7676);
nor UO_258 (O_258,N_8454,N_9875);
or UO_259 (O_259,N_7752,N_8317);
nand UO_260 (O_260,N_9392,N_8927);
xor UO_261 (O_261,N_9554,N_9333);
or UO_262 (O_262,N_8063,N_8041);
nand UO_263 (O_263,N_7737,N_7671);
nor UO_264 (O_264,N_9846,N_9628);
xnor UO_265 (O_265,N_8164,N_8731);
nand UO_266 (O_266,N_8323,N_9292);
or UO_267 (O_267,N_8244,N_8666);
nand UO_268 (O_268,N_9167,N_8248);
or UO_269 (O_269,N_7865,N_9084);
or UO_270 (O_270,N_7685,N_9092);
xnor UO_271 (O_271,N_8111,N_9457);
or UO_272 (O_272,N_8049,N_9315);
or UO_273 (O_273,N_9046,N_8638);
nand UO_274 (O_274,N_8737,N_8118);
xor UO_275 (O_275,N_9284,N_9121);
and UO_276 (O_276,N_8572,N_9832);
nand UO_277 (O_277,N_8094,N_9193);
nand UO_278 (O_278,N_7525,N_9806);
and UO_279 (O_279,N_8206,N_7549);
and UO_280 (O_280,N_8571,N_8508);
nor UO_281 (O_281,N_7600,N_8335);
and UO_282 (O_282,N_8879,N_8218);
xor UO_283 (O_283,N_9398,N_9769);
nand UO_284 (O_284,N_8941,N_8643);
or UO_285 (O_285,N_9508,N_8856);
or UO_286 (O_286,N_8161,N_9998);
nor UO_287 (O_287,N_7775,N_8208);
and UO_288 (O_288,N_7753,N_8038);
xor UO_289 (O_289,N_8876,N_9991);
nor UO_290 (O_290,N_7597,N_8198);
xor UO_291 (O_291,N_8002,N_8327);
and UO_292 (O_292,N_8460,N_8763);
or UO_293 (O_293,N_8186,N_9543);
nor UO_294 (O_294,N_9680,N_9334);
and UO_295 (O_295,N_9410,N_7745);
xor UO_296 (O_296,N_8689,N_8299);
and UO_297 (O_297,N_9981,N_9187);
or UO_298 (O_298,N_9748,N_9012);
nor UO_299 (O_299,N_9573,N_8368);
or UO_300 (O_300,N_8129,N_7726);
xor UO_301 (O_301,N_9568,N_9432);
or UO_302 (O_302,N_8315,N_8144);
xor UO_303 (O_303,N_9726,N_9858);
nor UO_304 (O_304,N_7793,N_7813);
or UO_305 (O_305,N_9248,N_9352);
xor UO_306 (O_306,N_7579,N_7658);
or UO_307 (O_307,N_8893,N_8160);
nand UO_308 (O_308,N_8577,N_8311);
nand UO_309 (O_309,N_8977,N_8650);
and UO_310 (O_310,N_7569,N_8655);
nor UO_311 (O_311,N_7757,N_7962);
and UO_312 (O_312,N_8432,N_9548);
or UO_313 (O_313,N_9293,N_7879);
nand UO_314 (O_314,N_8702,N_9296);
xor UO_315 (O_315,N_8873,N_9555);
nor UO_316 (O_316,N_9692,N_9329);
nor UO_317 (O_317,N_8721,N_7728);
nor UO_318 (O_318,N_8074,N_9463);
xor UO_319 (O_319,N_8882,N_9957);
and UO_320 (O_320,N_8668,N_8690);
nand UO_321 (O_321,N_9742,N_8455);
or UO_322 (O_322,N_9177,N_9759);
nor UO_323 (O_323,N_8243,N_8196);
or UO_324 (O_324,N_8796,N_9143);
or UO_325 (O_325,N_8602,N_7703);
nand UO_326 (O_326,N_8320,N_9452);
or UO_327 (O_327,N_8598,N_9175);
and UO_328 (O_328,N_9278,N_8040);
xnor UO_329 (O_329,N_8209,N_9433);
and UO_330 (O_330,N_8769,N_8970);
or UO_331 (O_331,N_8849,N_7938);
or UO_332 (O_332,N_9939,N_8520);
nand UO_333 (O_333,N_9028,N_9691);
nand UO_334 (O_334,N_9661,N_7800);
nand UO_335 (O_335,N_9590,N_9146);
or UO_336 (O_336,N_7820,N_9536);
and UO_337 (O_337,N_9775,N_9753);
xnor UO_338 (O_338,N_9454,N_8847);
and UO_339 (O_339,N_7607,N_7631);
xor UO_340 (O_340,N_9930,N_7700);
nor UO_341 (O_341,N_9205,N_8350);
nor UO_342 (O_342,N_8280,N_7736);
and UO_343 (O_343,N_8986,N_8929);
and UO_344 (O_344,N_9147,N_9250);
and UO_345 (O_345,N_7644,N_9920);
or UO_346 (O_346,N_7673,N_8285);
and UO_347 (O_347,N_8659,N_8959);
and UO_348 (O_348,N_8223,N_9308);
and UO_349 (O_349,N_9182,N_9363);
nor UO_350 (O_350,N_9470,N_8224);
xnor UO_351 (O_351,N_9752,N_7810);
or UO_352 (O_352,N_9260,N_8470);
and UO_353 (O_353,N_9609,N_7682);
nor UO_354 (O_354,N_8268,N_9450);
xor UO_355 (O_355,N_8426,N_7885);
xnor UO_356 (O_356,N_8440,N_8834);
and UO_357 (O_357,N_9813,N_7520);
nor UO_358 (O_358,N_9110,N_9963);
nor UO_359 (O_359,N_8291,N_9342);
and UO_360 (O_360,N_8980,N_8402);
nor UO_361 (O_361,N_8221,N_8048);
nand UO_362 (O_362,N_8725,N_8694);
and UO_363 (O_363,N_7951,N_9471);
or UO_364 (O_364,N_7572,N_7762);
or UO_365 (O_365,N_9784,N_8726);
and UO_366 (O_366,N_8069,N_9053);
xor UO_367 (O_367,N_8077,N_8034);
and UO_368 (O_368,N_8359,N_7617);
and UO_369 (O_369,N_9643,N_9673);
nand UO_370 (O_370,N_9190,N_7791);
nand UO_371 (O_371,N_9225,N_9123);
xor UO_372 (O_372,N_9029,N_8294);
nor UO_373 (O_373,N_8555,N_8310);
nand UO_374 (O_374,N_9200,N_7985);
nand UO_375 (O_375,N_8481,N_8249);
or UO_376 (O_376,N_9294,N_9702);
nand UO_377 (O_377,N_8717,N_8343);
nand UO_378 (O_378,N_8089,N_8850);
xnor UO_379 (O_379,N_7995,N_8633);
nor UO_380 (O_380,N_7738,N_9364);
or UO_381 (O_381,N_9196,N_7959);
nand UO_382 (O_382,N_8791,N_8443);
nor UO_383 (O_383,N_7586,N_8568);
or UO_384 (O_384,N_8639,N_7949);
nor UO_385 (O_385,N_8550,N_9712);
xor UO_386 (O_386,N_9034,N_8428);
nand UO_387 (O_387,N_8180,N_8295);
and UO_388 (O_388,N_9151,N_8991);
and UO_389 (O_389,N_9427,N_7749);
nor UO_390 (O_390,N_9227,N_9429);
and UO_391 (O_391,N_7786,N_8067);
nor UO_392 (O_392,N_8695,N_9644);
nor UO_393 (O_393,N_8776,N_9498);
and UO_394 (O_394,N_9553,N_9533);
nor UO_395 (O_395,N_8260,N_8047);
or UO_396 (O_396,N_8234,N_8583);
nor UO_397 (O_397,N_8326,N_9306);
and UO_398 (O_398,N_7536,N_8608);
or UO_399 (O_399,N_7628,N_9394);
nor UO_400 (O_400,N_7923,N_9426);
nand UO_401 (O_401,N_8938,N_8499);
or UO_402 (O_402,N_9311,N_8145);
nor UO_403 (O_403,N_9780,N_8138);
and UO_404 (O_404,N_8685,N_8869);
xnor UO_405 (O_405,N_8143,N_8006);
nand UO_406 (O_406,N_7893,N_9360);
xor UO_407 (O_407,N_8674,N_8514);
nor UO_408 (O_408,N_8997,N_8881);
and UO_409 (O_409,N_8346,N_9997);
xnor UO_410 (O_410,N_7721,N_9493);
nor UO_411 (O_411,N_8510,N_8972);
and UO_412 (O_412,N_9244,N_7792);
nor UO_413 (O_413,N_8219,N_9954);
nor UO_414 (O_414,N_9074,N_8182);
nor UO_415 (O_415,N_9677,N_9056);
nor UO_416 (O_416,N_8241,N_9236);
or UO_417 (O_417,N_9633,N_8888);
xor UO_418 (O_418,N_7582,N_8284);
and UO_419 (O_419,N_9521,N_7934);
nor UO_420 (O_420,N_9319,N_8842);
and UO_421 (O_421,N_7677,N_8880);
and UO_422 (O_422,N_8556,N_9212);
and UO_423 (O_423,N_9545,N_9478);
nand UO_424 (O_424,N_9058,N_8672);
xor UO_425 (O_425,N_8387,N_8042);
nand UO_426 (O_426,N_8484,N_8487);
nor UO_427 (O_427,N_7667,N_9722);
or UO_428 (O_428,N_9988,N_9174);
and UO_429 (O_429,N_9291,N_8781);
nor UO_430 (O_430,N_8540,N_9574);
and UO_431 (O_431,N_7668,N_8420);
nor UO_432 (O_432,N_7944,N_7680);
xnor UO_433 (O_433,N_7678,N_9902);
or UO_434 (O_434,N_7725,N_7636);
xnor UO_435 (O_435,N_9312,N_7648);
xor UO_436 (O_436,N_9815,N_9785);
xor UO_437 (O_437,N_8175,N_9373);
or UO_438 (O_438,N_9362,N_7684);
and UO_439 (O_439,N_9540,N_7548);
nor UO_440 (O_440,N_8459,N_9886);
or UO_441 (O_441,N_8081,N_8762);
and UO_442 (O_442,N_7779,N_8709);
and UO_443 (O_443,N_9439,N_8586);
nand UO_444 (O_444,N_9399,N_8055);
nand UO_445 (O_445,N_9386,N_9922);
nor UO_446 (O_446,N_7718,N_8808);
and UO_447 (O_447,N_8199,N_9455);
and UO_448 (O_448,N_9777,N_8181);
and UO_449 (O_449,N_8059,N_7892);
nor UO_450 (O_450,N_9653,N_9458);
xnor UO_451 (O_451,N_8878,N_8995);
and UO_452 (O_452,N_7584,N_8778);
nor UO_453 (O_453,N_8134,N_9916);
and UO_454 (O_454,N_8914,N_7912);
or UO_455 (O_455,N_9222,N_8937);
or UO_456 (O_456,N_9502,N_7641);
nor UO_457 (O_457,N_8676,N_8490);
xnor UO_458 (O_458,N_8793,N_8297);
nor UO_459 (O_459,N_9755,N_9141);
or UO_460 (O_460,N_8498,N_7783);
nand UO_461 (O_461,N_8751,N_9559);
nand UO_462 (O_462,N_9063,N_8706);
xor UO_463 (O_463,N_8231,N_8573);
xor UO_464 (O_464,N_9899,N_7850);
xor UO_465 (O_465,N_8251,N_8823);
or UO_466 (O_466,N_9960,N_7588);
nor UO_467 (O_467,N_9109,N_8748);
and UO_468 (O_468,N_8361,N_9052);
xor UO_469 (O_469,N_7533,N_7534);
nand UO_470 (O_470,N_7553,N_7560);
and UO_471 (O_471,N_7681,N_8909);
or UO_472 (O_472,N_8513,N_9246);
and UO_473 (O_473,N_9717,N_9941);
or UO_474 (O_474,N_9640,N_7741);
nand UO_475 (O_475,N_8988,N_8395);
or UO_476 (O_476,N_7802,N_7989);
nand UO_477 (O_477,N_9605,N_8101);
or UO_478 (O_478,N_7927,N_9589);
nand UO_479 (O_479,N_7756,N_9013);
and UO_480 (O_480,N_7592,N_9270);
xnor UO_481 (O_481,N_9233,N_9667);
and UO_482 (O_482,N_8859,N_7695);
xor UO_483 (O_483,N_7570,N_9374);
or UO_484 (O_484,N_9649,N_7855);
or UO_485 (O_485,N_8993,N_8810);
and UO_486 (O_486,N_7519,N_7564);
or UO_487 (O_487,N_7917,N_7545);
or UO_488 (O_488,N_9272,N_7732);
nand UO_489 (O_489,N_9546,N_9161);
xor UO_490 (O_490,N_8347,N_7540);
nand UO_491 (O_491,N_7587,N_9125);
xor UO_492 (O_492,N_8419,N_9578);
and UO_493 (O_493,N_9290,N_8113);
and UO_494 (O_494,N_8509,N_8456);
nand UO_495 (O_495,N_7826,N_9840);
or UO_496 (O_496,N_9324,N_9516);
xor UO_497 (O_497,N_8269,N_9382);
or UO_498 (O_498,N_9388,N_9976);
xor UO_499 (O_499,N_8848,N_9108);
nand UO_500 (O_500,N_8400,N_8388);
and UO_501 (O_501,N_8298,N_8708);
nor UO_502 (O_502,N_7690,N_9127);
or UO_503 (O_503,N_8125,N_8281);
or UO_504 (O_504,N_7926,N_8156);
nor UO_505 (O_505,N_9917,N_7646);
nand UO_506 (O_506,N_8619,N_9208);
or UO_507 (O_507,N_9926,N_9479);
or UO_508 (O_508,N_9179,N_8013);
xor UO_509 (O_509,N_8092,N_7639);
or UO_510 (O_510,N_9318,N_7526);
nor UO_511 (O_511,N_8789,N_9480);
or UO_512 (O_512,N_7630,N_8536);
or UO_513 (O_513,N_7861,N_9622);
and UO_514 (O_514,N_8788,N_9335);
xor UO_515 (O_515,N_7911,N_9796);
nor UO_516 (O_516,N_9668,N_8952);
nand UO_517 (O_517,N_8906,N_9771);
or UO_518 (O_518,N_7935,N_8830);
nand UO_519 (O_519,N_9513,N_8448);
xor UO_520 (O_520,N_8657,N_8625);
or UO_521 (O_521,N_8242,N_7897);
nor UO_522 (O_522,N_9214,N_8194);
or UO_523 (O_523,N_7704,N_8469);
xnor UO_524 (O_524,N_9715,N_7637);
xnor UO_525 (O_525,N_9978,N_9579);
or UO_526 (O_526,N_9809,N_9662);
and UO_527 (O_527,N_9751,N_8008);
and UO_528 (O_528,N_9581,N_8795);
nor UO_529 (O_529,N_9944,N_8060);
nor UO_530 (O_530,N_9049,N_7854);
nand UO_531 (O_531,N_9253,N_9664);
nand UO_532 (O_532,N_9079,N_7620);
nand UO_533 (O_533,N_8892,N_8273);
nand UO_534 (O_534,N_7870,N_8517);
and UO_535 (O_535,N_7521,N_7769);
or UO_536 (O_536,N_9422,N_9280);
or UO_537 (O_537,N_9826,N_9093);
and UO_538 (O_538,N_9269,N_9737);
nor UO_539 (O_539,N_8110,N_9665);
nor UO_540 (O_540,N_9500,N_7669);
and UO_541 (O_541,N_9226,N_9224);
nand UO_542 (O_542,N_8300,N_8961);
or UO_543 (O_543,N_8558,N_7983);
nor UO_544 (O_544,N_9972,N_9685);
nor UO_545 (O_545,N_8724,N_8215);
nor UO_546 (O_546,N_8667,N_9055);
and UO_547 (O_547,N_9595,N_8141);
nor UO_548 (O_548,N_9300,N_9584);
or UO_549 (O_549,N_9889,N_7723);
nand UO_550 (O_550,N_9154,N_8495);
or UO_551 (O_551,N_7555,N_8338);
and UO_552 (O_552,N_7750,N_7625);
or UO_553 (O_553,N_8579,N_9973);
xor UO_554 (O_554,N_9183,N_8112);
nand UO_555 (O_555,N_8930,N_9909);
or UO_556 (O_556,N_9142,N_7710);
nand UO_557 (O_557,N_9395,N_9409);
xnor UO_558 (O_558,N_8135,N_8261);
nor UO_559 (O_559,N_8660,N_9839);
nand UO_560 (O_560,N_8978,N_9418);
nor UO_561 (O_561,N_8530,N_7785);
nor UO_562 (O_562,N_9378,N_8584);
nor UO_563 (O_563,N_9670,N_9526);
nor UO_564 (O_564,N_8853,N_8011);
and UO_565 (O_565,N_8009,N_8895);
or UO_566 (O_566,N_7575,N_8803);
nand UO_567 (O_567,N_8418,N_7808);
xnor UO_568 (O_568,N_8560,N_7877);
and UO_569 (O_569,N_8005,N_9934);
xor UO_570 (O_570,N_8393,N_8855);
nand UO_571 (O_571,N_9828,N_9591);
xor UO_572 (O_572,N_7976,N_8766);
nand UO_573 (O_573,N_7891,N_7840);
or UO_574 (O_574,N_7594,N_9327);
nand UO_575 (O_575,N_8169,N_8130);
xnor UO_576 (O_576,N_8096,N_8637);
and UO_577 (O_577,N_9022,N_9356);
nor UO_578 (O_578,N_9304,N_9031);
xnor UO_579 (O_579,N_8401,N_8107);
or UO_580 (O_580,N_8564,N_8151);
or UO_581 (O_581,N_8794,N_7714);
xnor UO_582 (O_582,N_9614,N_7895);
and UO_583 (O_583,N_8373,N_8203);
xnor UO_584 (O_584,N_8606,N_9243);
nand UO_585 (O_585,N_9950,N_9275);
nand UO_586 (O_586,N_8620,N_7727);
and UO_587 (O_587,N_9896,N_9014);
or UO_588 (O_588,N_8651,N_9562);
or UO_589 (O_589,N_9719,N_9524);
nor UO_590 (O_590,N_8958,N_8245);
and UO_591 (O_591,N_8384,N_9764);
nor UO_592 (O_592,N_8330,N_8482);
xor UO_593 (O_593,N_8197,N_9874);
nor UO_594 (O_594,N_9514,N_7731);
nand UO_595 (O_595,N_7832,N_8480);
nand UO_596 (O_596,N_8802,N_8434);
and UO_597 (O_597,N_9295,N_8716);
nand UO_598 (O_598,N_8545,N_8837);
xor UO_599 (O_599,N_8679,N_8202);
nand UO_600 (O_600,N_8422,N_8331);
and UO_601 (O_601,N_7823,N_8705);
nand UO_602 (O_602,N_7556,N_9038);
or UO_603 (O_603,N_9402,N_8525);
nand UO_604 (O_604,N_8475,N_9245);
nand UO_605 (O_605,N_9790,N_7799);
xnor UO_606 (O_606,N_7716,N_8439);
or UO_607 (O_607,N_9495,N_8819);
xnor UO_608 (O_608,N_8085,N_7839);
xor UO_609 (O_609,N_9380,N_9129);
nor UO_610 (O_610,N_8272,N_9940);
nand UO_611 (O_611,N_9577,N_8216);
nand UO_612 (O_612,N_8897,N_9408);
nand UO_613 (O_613,N_8492,N_8468);
xor UO_614 (O_614,N_9877,N_8365);
nand UO_615 (O_615,N_7932,N_8574);
nor UO_616 (O_616,N_8631,N_8624);
nor UO_617 (O_617,N_7653,N_9496);
nor UO_618 (O_618,N_7674,N_7567);
nor UO_619 (O_619,N_8673,N_9765);
and UO_620 (O_620,N_8287,N_9003);
and UO_621 (O_621,N_8149,N_8362);
nor UO_622 (O_622,N_9598,N_9157);
nor UO_623 (O_623,N_7605,N_8430);
nand UO_624 (O_624,N_7990,N_7954);
nand UO_625 (O_625,N_8783,N_8099);
or UO_626 (O_626,N_8671,N_9017);
xor UO_627 (O_627,N_8727,N_8531);
xnor UO_628 (O_628,N_9424,N_8757);
xnor UO_629 (O_629,N_9499,N_8752);
nand UO_630 (O_630,N_8665,N_7576);
nand UO_631 (O_631,N_7537,N_9905);
nor UO_632 (O_632,N_7915,N_8764);
nor UO_633 (O_633,N_7996,N_8758);
nand UO_634 (O_634,N_9937,N_9766);
nand UO_635 (O_635,N_9325,N_7760);
xnor UO_636 (O_636,N_8732,N_9309);
xor UO_637 (O_637,N_8375,N_9144);
nor UO_638 (O_638,N_9678,N_8479);
nor UO_639 (O_639,N_9397,N_8366);
xor UO_640 (O_640,N_9069,N_8771);
nand UO_641 (O_641,N_9671,N_8147);
nor UO_642 (O_642,N_7909,N_9672);
and UO_643 (O_643,N_7503,N_9379);
or UO_644 (O_644,N_7999,N_9050);
nor UO_645 (O_645,N_7960,N_9686);
nor UO_646 (O_646,N_9637,N_9650);
xor UO_647 (O_647,N_9119,N_8987);
nor UO_648 (O_648,N_8773,N_8699);
nor UO_649 (O_649,N_8288,N_9156);
nor UO_650 (O_650,N_9968,N_9172);
xor UO_651 (O_651,N_8516,N_9025);
nand UO_652 (O_652,N_9657,N_9197);
xor UO_653 (O_653,N_9338,N_8811);
nand UO_654 (O_654,N_8640,N_9100);
nor UO_655 (O_655,N_8653,N_8132);
and UO_656 (O_656,N_9383,N_9462);
nor UO_657 (O_657,N_8982,N_8797);
nor UO_658 (O_658,N_9210,N_9744);
xor UO_659 (O_659,N_8933,N_8227);
xor UO_660 (O_660,N_9929,N_8535);
xor UO_661 (O_661,N_8840,N_7881);
or UO_662 (O_662,N_8371,N_9341);
nor UO_663 (O_663,N_7965,N_9355);
or UO_664 (O_664,N_9145,N_8928);
xnor UO_665 (O_665,N_7670,N_8865);
xor UO_666 (O_666,N_9980,N_7794);
or UO_667 (O_667,N_7604,N_9942);
nor UO_668 (O_668,N_8435,N_7958);
nand UO_669 (O_669,N_9860,N_9042);
and UO_670 (O_670,N_9827,N_7968);
xnor UO_671 (O_671,N_9186,N_8154);
nand UO_672 (O_672,N_7707,N_7930);
xnor UO_673 (O_673,N_9928,N_9675);
nand UO_674 (O_674,N_8753,N_8627);
and UO_675 (O_675,N_8212,N_8974);
nand UO_676 (O_676,N_7801,N_9787);
xnor UO_677 (O_677,N_9818,N_8939);
xor UO_678 (O_678,N_8344,N_8256);
xnor UO_679 (O_679,N_8157,N_7610);
xnor UO_680 (O_680,N_9460,N_9506);
xnor UO_681 (O_681,N_8870,N_8786);
nand UO_682 (O_682,N_9833,N_8037);
and UO_683 (O_683,N_8033,N_9435);
nor UO_684 (O_684,N_8225,N_8611);
xnor UO_685 (O_685,N_9347,N_9117);
and UO_686 (O_686,N_9385,N_9669);
nor UO_687 (O_687,N_7984,N_8083);
or UO_688 (O_688,N_9033,N_8907);
and UO_689 (O_689,N_8163,N_7910);
nor UO_690 (O_690,N_9798,N_9251);
or UO_691 (O_691,N_8981,N_9733);
nor UO_692 (O_692,N_9414,N_9505);
or UO_693 (O_693,N_8523,N_8591);
nor UO_694 (O_694,N_9760,N_9714);
nand UO_695 (O_695,N_8054,N_8140);
and UO_696 (O_696,N_9550,N_8367);
nor UO_697 (O_697,N_9674,N_7552);
nand UO_698 (O_698,N_9999,N_9343);
nor UO_699 (O_699,N_9525,N_8784);
nor UO_700 (O_700,N_8956,N_8692);
xnor UO_701 (O_701,N_9020,N_9597);
xnor UO_702 (O_702,N_7998,N_7797);
or UO_703 (O_703,N_9741,N_8553);
nor UO_704 (O_704,N_9365,N_9400);
or UO_705 (O_705,N_9337,N_7505);
nand UO_706 (O_706,N_8166,N_9078);
nand UO_707 (O_707,N_9831,N_8971);
nand UO_708 (O_708,N_9829,N_7888);
or UO_709 (O_709,N_8491,N_8609);
xor UO_710 (O_710,N_7788,N_9551);
and UO_711 (O_711,N_8759,N_7515);
or UO_712 (O_712,N_8137,N_9611);
nand UO_713 (O_713,N_7875,N_8992);
nand UO_714 (O_714,N_8524,N_8792);
or UO_715 (O_715,N_9194,N_9443);
and UO_716 (O_716,N_7973,N_9949);
or UO_717 (O_717,N_9211,N_8086);
or UO_718 (O_718,N_7921,N_7977);
or UO_719 (O_719,N_8654,N_8871);
nand UO_720 (O_720,N_9310,N_9162);
xor UO_721 (O_721,N_9384,N_9921);
nor UO_722 (O_722,N_7914,N_9983);
xnor UO_723 (O_723,N_8615,N_7654);
and UO_724 (O_724,N_9800,N_7522);
and UO_725 (O_725,N_9510,N_9114);
xnor UO_726 (O_726,N_9811,N_9237);
and UO_727 (O_727,N_9256,N_7837);
nand UO_728 (O_728,N_8772,N_9447);
or UO_729 (O_729,N_7986,N_8457);
nand UO_730 (O_730,N_7842,N_9974);
xnor UO_731 (O_731,N_9016,N_7589);
xor UO_732 (O_732,N_9625,N_9009);
and UO_733 (O_733,N_9904,N_9102);
xor UO_734 (O_734,N_7694,N_9897);
xor UO_735 (O_735,N_9351,N_9616);
or UO_736 (O_736,N_9863,N_9627);
nor UO_737 (O_737,N_8526,N_8538);
and UO_738 (O_738,N_8504,N_8461);
nand UO_739 (O_739,N_8528,N_8262);
or UO_740 (O_740,N_8045,N_8919);
nand UO_741 (O_741,N_7761,N_9131);
nor UO_742 (O_742,N_7833,N_7980);
xor UO_743 (O_743,N_7735,N_9051);
or UO_744 (O_744,N_8374,N_9062);
and UO_745 (O_745,N_7966,N_9795);
nand UO_746 (O_746,N_8585,N_9641);
and UO_747 (O_747,N_9876,N_8399);
nand UO_748 (O_748,N_9924,N_9814);
nand UO_749 (O_749,N_7508,N_8127);
nand UO_750 (O_750,N_9586,N_9965);
nor UO_751 (O_751,N_9032,N_9191);
and UO_752 (O_752,N_8021,N_9168);
nand UO_753 (O_753,N_9770,N_8275);
nor UO_754 (O_754,N_7516,N_9420);
nor UO_755 (O_755,N_9808,N_7629);
nor UO_756 (O_756,N_9266,N_8539);
or UO_757 (O_757,N_7702,N_8257);
nand UO_758 (O_758,N_8990,N_8238);
nor UO_759 (O_759,N_7953,N_7774);
nand UO_760 (O_760,N_8302,N_8354);
xor UO_761 (O_761,N_9104,N_9068);
nand UO_762 (O_762,N_9339,N_9841);
and UO_763 (O_763,N_9476,N_9440);
nor UO_764 (O_764,N_9542,N_9067);
nand UO_765 (O_765,N_8053,N_9279);
nand UO_766 (O_766,N_9792,N_9881);
or UO_767 (O_767,N_8549,N_8080);
nor UO_768 (O_768,N_9076,N_8483);
and UO_769 (O_769,N_9724,N_7994);
and UO_770 (O_770,N_8236,N_9035);
and UO_771 (O_771,N_8798,N_7903);
nor UO_772 (O_772,N_7538,N_8681);
nand UO_773 (O_773,N_8423,N_9626);
or UO_774 (O_774,N_7916,N_9070);
nand UO_775 (O_775,N_8406,N_7571);
xnor UO_776 (O_776,N_9305,N_9249);
xnor UO_777 (O_777,N_8913,N_7546);
xor UO_778 (O_778,N_8534,N_7831);
xnor UO_779 (O_779,N_8473,N_9654);
and UO_780 (O_780,N_8682,N_7591);
or UO_781 (O_781,N_8233,N_9594);
nor UO_782 (O_782,N_9336,N_8581);
nand UO_783 (O_783,N_8594,N_9610);
xor UO_784 (O_784,N_9189,N_8736);
or UO_785 (O_785,N_8812,N_9456);
xor UO_786 (O_786,N_7621,N_9150);
xnor UO_787 (O_787,N_7835,N_7771);
xor UO_788 (O_788,N_8734,N_9781);
nor UO_789 (O_789,N_9774,N_8316);
nor UO_790 (O_790,N_8486,N_8195);
or UO_791 (O_791,N_9776,N_8861);
or UO_792 (O_792,N_7836,N_8030);
and UO_793 (O_793,N_8087,N_8119);
xor UO_794 (O_794,N_9095,N_9958);
xnor UO_795 (O_795,N_7514,N_8103);
or UO_796 (O_796,N_9198,N_9868);
nor UO_797 (O_797,N_7624,N_9624);
nand UO_798 (O_798,N_8322,N_7992);
nor UO_799 (O_799,N_8172,N_9005);
and UO_800 (O_800,N_9565,N_8890);
and UO_801 (O_801,N_9345,N_9732);
nand UO_802 (O_802,N_9867,N_7517);
and UO_803 (O_803,N_8942,N_7744);
and UO_804 (O_804,N_8405,N_9085);
and UO_805 (O_805,N_9176,N_7632);
nor UO_806 (O_806,N_8324,N_8741);
nor UO_807 (O_807,N_9448,N_9569);
xor UO_808 (O_808,N_7830,N_8742);
or UO_809 (O_809,N_9064,N_9047);
and UO_810 (O_810,N_8345,N_8305);
xor UO_811 (O_811,N_8108,N_8529);
and UO_812 (O_812,N_7847,N_9185);
nand UO_813 (O_813,N_8024,N_8924);
nor UO_814 (O_814,N_8403,N_7907);
nand UO_815 (O_815,N_8079,N_8408);
nor UO_816 (O_816,N_7991,N_8425);
nor UO_817 (O_817,N_7626,N_7770);
and UO_818 (O_818,N_9738,N_9135);
or UO_819 (O_819,N_7645,N_7929);
nor UO_820 (O_820,N_9126,N_8139);
and UO_821 (O_821,N_7558,N_9507);
nand UO_822 (O_822,N_8072,N_8874);
xnor UO_823 (O_823,N_8559,N_8805);
xnor UO_824 (O_824,N_9081,N_9547);
xor UO_825 (O_825,N_7504,N_8629);
xnor UO_826 (O_826,N_8955,N_8713);
xnor UO_827 (O_827,N_8587,N_9990);
and UO_828 (O_828,N_9791,N_9855);
or UO_829 (O_829,N_8477,N_7565);
or UO_830 (O_830,N_7773,N_8026);
nand UO_831 (O_831,N_7817,N_8738);
nand UO_832 (O_832,N_9789,N_8303);
xor UO_833 (O_833,N_9996,N_7686);
or UO_834 (O_834,N_8838,N_7906);
xnor UO_835 (O_835,N_8472,N_7913);
or UO_836 (O_836,N_9927,N_8593);
xor UO_837 (O_837,N_8590,N_9825);
xor UO_838 (O_838,N_9982,N_7510);
or UO_839 (O_839,N_8698,N_8232);
and UO_840 (O_840,N_7557,N_9956);
xor UO_841 (O_841,N_8744,N_8433);
and UO_842 (O_842,N_9321,N_8497);
xor UO_843 (O_843,N_9060,N_8286);
nor UO_844 (O_844,N_8429,N_9430);
xor UO_845 (O_845,N_8512,N_8911);
nand UO_846 (O_846,N_9136,N_8007);
or UO_847 (O_847,N_9484,N_8719);
nor UO_848 (O_848,N_9821,N_9213);
and UO_849 (O_849,N_9094,N_7798);
nor UO_850 (O_850,N_8875,N_9314);
nand UO_851 (O_851,N_8097,N_9763);
nand UO_852 (O_852,N_7777,N_7997);
and UO_853 (O_853,N_8237,N_8807);
and UO_854 (O_854,N_9368,N_9801);
xor UO_855 (O_855,N_9138,N_9613);
xnor UO_856 (O_856,N_9503,N_8806);
xnor UO_857 (O_857,N_8887,N_8438);
or UO_858 (O_858,N_9694,N_7611);
nor UO_859 (O_859,N_9118,N_7748);
xor UO_860 (O_860,N_9803,N_8733);
xnor UO_861 (O_861,N_7787,N_9173);
nand UO_862 (O_862,N_9349,N_8935);
nor UO_863 (O_863,N_9967,N_9285);
or UO_864 (O_864,N_9879,N_9441);
nand UO_865 (O_865,N_9786,N_7964);
and UO_866 (O_866,N_9636,N_9203);
and UO_867 (O_867,N_9587,N_8533);
and UO_868 (O_868,N_9288,N_9286);
and UO_869 (O_869,N_9931,N_7931);
xor UO_870 (O_870,N_8883,N_9019);
and UO_871 (O_871,N_9725,N_7872);
or UO_872 (O_872,N_9008,N_7563);
xor UO_873 (O_873,N_9071,N_8506);
xor UO_874 (O_874,N_9011,N_9453);
and UO_875 (O_875,N_9601,N_8596);
or UO_876 (O_876,N_8813,N_9234);
nor UO_877 (O_877,N_9848,N_8431);
xnor UO_878 (O_878,N_9018,N_8775);
nand UO_879 (O_879,N_9560,N_8267);
xor UO_880 (O_880,N_9169,N_8765);
nand UO_881 (O_881,N_8409,N_8975);
nand UO_882 (O_882,N_9097,N_9761);
nand UO_883 (O_883,N_8357,N_8358);
and UO_884 (O_884,N_9264,N_8926);
nor UO_885 (O_885,N_7766,N_9959);
nor UO_886 (O_886,N_7969,N_8614);
or UO_887 (O_887,N_8122,N_9482);
xor UO_888 (O_888,N_7883,N_8003);
nand UO_889 (O_889,N_8944,N_9708);
xnor UO_890 (O_890,N_7945,N_9793);
nand UO_891 (O_891,N_8617,N_9971);
xor UO_892 (O_892,N_8229,N_8503);
nor UO_893 (O_893,N_8632,N_8561);
or UO_894 (O_894,N_8934,N_8416);
nor UO_895 (O_895,N_9683,N_9158);
nand UO_896 (O_896,N_9890,N_8950);
or UO_897 (O_897,N_8458,N_8670);
or UO_898 (O_898,N_7657,N_8621);
and UO_899 (O_899,N_8264,N_8489);
xor UO_900 (O_900,N_8488,N_8965);
nor UO_901 (O_901,N_9231,N_9159);
nor UO_902 (O_902,N_9026,N_7852);
nand UO_903 (O_903,N_9606,N_8377);
nand UO_904 (O_904,N_9350,N_8662);
nor UO_905 (O_905,N_8829,N_9985);
and UO_906 (O_906,N_8966,N_9684);
and UO_907 (O_907,N_8360,N_7922);
or UO_908 (O_908,N_9852,N_9945);
and UO_909 (O_909,N_7981,N_8648);
nand UO_910 (O_910,N_7561,N_9181);
or UO_911 (O_911,N_9209,N_9588);
or UO_912 (O_912,N_9709,N_9970);
xnor UO_913 (O_913,N_8943,N_8170);
nor UO_914 (O_914,N_8949,N_8001);
or UO_915 (O_915,N_8872,N_9895);
or UO_916 (O_916,N_9098,N_7532);
xnor UO_917 (O_917,N_8471,N_7722);
or UO_918 (O_918,N_8337,N_7651);
nand UO_919 (O_919,N_7978,N_9953);
and UO_920 (O_920,N_9075,N_8612);
nor UO_921 (O_921,N_9544,N_9406);
nor UO_922 (O_922,N_8004,N_9366);
nor UO_923 (O_923,N_8973,N_8062);
nor UO_924 (O_924,N_7806,N_9001);
nand UO_925 (O_925,N_8989,N_9632);
xnor UO_926 (O_926,N_8391,N_7974);
or UO_927 (O_927,N_9913,N_7581);
or UO_928 (O_928,N_8825,N_8547);
xor UO_929 (O_929,N_7739,N_9207);
and UO_930 (O_930,N_9043,N_7919);
and UO_931 (O_931,N_9259,N_8351);
nor UO_932 (O_932,N_9041,N_7948);
xor UO_933 (O_933,N_8544,N_8217);
nand UO_934 (O_934,N_9617,N_7925);
nor UO_935 (O_935,N_8750,N_8073);
and UO_936 (O_936,N_7987,N_8828);
xor UO_937 (O_937,N_9152,N_8996);
and UO_938 (O_938,N_8994,N_8852);
nand UO_939 (O_939,N_8841,N_8378);
or UO_940 (O_940,N_8474,N_9853);
xor UO_941 (O_941,N_8901,N_9582);
and UO_942 (O_942,N_7956,N_7719);
nand UO_943 (O_943,N_9332,N_8616);
nand UO_944 (O_944,N_8940,N_9405);
or UO_945 (O_945,N_7869,N_7821);
nor UO_946 (O_946,N_9367,N_9268);
nand UO_947 (O_947,N_9530,N_9892);
and UO_948 (O_948,N_8600,N_9619);
nand UO_949 (O_949,N_8027,N_9446);
and UO_950 (O_950,N_9580,N_9933);
xnor UO_951 (O_951,N_8029,N_7699);
or UO_952 (O_952,N_9994,N_8444);
and UO_953 (O_953,N_9782,N_9856);
and UO_954 (O_954,N_7818,N_8379);
xor UO_955 (O_955,N_9871,N_8723);
or UO_956 (O_956,N_7663,N_9487);
xor UO_957 (O_957,N_7717,N_9330);
nor UO_958 (O_958,N_9621,N_8035);
nor UO_959 (O_959,N_9287,N_8100);
nor UO_960 (O_960,N_7924,N_8755);
and UO_961 (O_961,N_9865,N_9088);
nand UO_962 (O_962,N_8582,N_9148);
and UO_963 (O_963,N_8824,N_8019);
nor UO_964 (O_964,N_9485,N_8424);
xnor UO_965 (O_965,N_8052,N_9630);
or UO_966 (O_966,N_8446,N_9103);
nor UO_967 (O_967,N_7871,N_7733);
and UO_968 (O_968,N_8066,N_7666);
nand UO_969 (O_969,N_8386,N_9682);
or UO_970 (O_970,N_9864,N_9908);
xor UO_971 (O_971,N_8396,N_9219);
nor UO_972 (O_972,N_7764,N_7619);
and UO_973 (O_973,N_8658,N_7778);
xnor UO_974 (O_974,N_9087,N_7946);
nor UO_975 (O_975,N_8562,N_9469);
or UO_976 (O_976,N_7609,N_9716);
nor UO_977 (O_977,N_7615,N_8903);
and UO_978 (O_978,N_9002,N_7697);
xnor UO_979 (O_979,N_9822,N_8210);
or UO_980 (O_980,N_8191,N_8703);
nor UO_981 (O_981,N_9358,N_9883);
and UO_982 (O_982,N_8381,N_8605);
or UO_983 (O_983,N_9519,N_8962);
and UO_984 (O_984,N_9914,N_7859);
nor UO_985 (O_985,N_7846,N_8126);
nor UO_986 (O_986,N_7634,N_7724);
nand UO_987 (O_987,N_9421,N_8576);
xor UO_988 (O_988,N_9024,N_8383);
and UO_989 (O_989,N_9804,N_8090);
nor UO_990 (O_990,N_8442,N_9091);
xnor UO_991 (O_991,N_7734,N_8521);
nor UO_992 (O_992,N_7825,N_8404);
nor UO_993 (O_993,N_9298,N_9504);
xnor UO_994 (O_994,N_9240,N_9873);
nand UO_995 (O_995,N_8700,N_8247);
xor UO_996 (O_996,N_9534,N_9535);
nor UO_997 (O_997,N_8683,N_9736);
nand UO_998 (O_998,N_9215,N_8279);
nor UO_999 (O_999,N_8664,N_8064);
nand UO_1000 (O_1000,N_7656,N_9634);
xnor UO_1001 (O_1001,N_8710,N_7687);
or UO_1002 (O_1002,N_9436,N_8908);
or UO_1003 (O_1003,N_7675,N_8015);
nor UO_1004 (O_1004,N_8696,N_7742);
and UO_1005 (O_1005,N_8844,N_8159);
xor UO_1006 (O_1006,N_9870,N_9952);
nor UO_1007 (O_1007,N_8010,N_8678);
xor UO_1008 (O_1008,N_8910,N_7506);
and UO_1009 (O_1009,N_7647,N_8339);
or UO_1010 (O_1010,N_8296,N_9566);
and UO_1011 (O_1011,N_8167,N_7711);
or UO_1012 (O_1012,N_7577,N_8720);
and UO_1013 (O_1013,N_9880,N_8863);
xnor UO_1014 (O_1014,N_7580,N_9728);
nand UO_1015 (O_1015,N_8967,N_9438);
xor UO_1016 (O_1016,N_8308,N_8493);
and UO_1017 (O_1017,N_8626,N_7763);
nand UO_1018 (O_1018,N_9004,N_8898);
nor UO_1019 (O_1019,N_9773,N_9700);
nand UO_1020 (O_1020,N_8846,N_8290);
xor UO_1021 (O_1021,N_7848,N_8603);
nand UO_1022 (O_1022,N_9401,N_7701);
nor UO_1023 (O_1023,N_9984,N_7751);
nor UO_1024 (O_1024,N_8951,N_9615);
nor UO_1025 (O_1025,N_7827,N_8686);
xnor UO_1026 (O_1026,N_9160,N_7868);
or UO_1027 (O_1027,N_8148,N_8832);
xnor UO_1028 (O_1028,N_8704,N_9697);
nor UO_1029 (O_1029,N_8070,N_8754);
xor UO_1030 (O_1030,N_8255,N_7936);
nand UO_1031 (O_1031,N_9936,N_8779);
and UO_1032 (O_1032,N_9567,N_9331);
xnor UO_1033 (O_1033,N_8036,N_8123);
or UO_1034 (O_1034,N_8023,N_9235);
xor UO_1035 (O_1035,N_7573,N_8954);
and UO_1036 (O_1036,N_8920,N_8259);
nand UO_1037 (O_1037,N_8715,N_9445);
xor UO_1038 (O_1038,N_8777,N_9989);
xnor UO_1039 (O_1039,N_9301,N_8417);
and UO_1040 (O_1040,N_9178,N_7709);
nor UO_1041 (O_1041,N_8051,N_9842);
or UO_1042 (O_1042,N_7943,N_7541);
nand UO_1043 (O_1043,N_8082,N_7618);
nand UO_1044 (O_1044,N_8254,N_7904);
or UO_1045 (O_1045,N_7790,N_8860);
nand UO_1046 (O_1046,N_9419,N_9919);
or UO_1047 (O_1047,N_9797,N_7754);
xor UO_1048 (O_1048,N_7608,N_9576);
or UO_1049 (O_1049,N_8831,N_9635);
nor UO_1050 (O_1050,N_8342,N_9975);
nand UO_1051 (O_1051,N_7643,N_8332);
nor UO_1052 (O_1052,N_7649,N_9652);
nor UO_1053 (O_1053,N_7635,N_9910);
or UO_1054 (O_1054,N_9375,N_8785);
nand UO_1055 (O_1055,N_8688,N_8554);
xor UO_1056 (O_1056,N_7759,N_8478);
xor UO_1057 (O_1057,N_9313,N_7664);
or UO_1058 (O_1058,N_9000,N_7812);
nand UO_1059 (O_1059,N_9149,N_8845);
or UO_1060 (O_1060,N_9608,N_8153);
nand UO_1061 (O_1061,N_8283,N_9729);
xnor UO_1062 (O_1062,N_8826,N_8192);
or UO_1063 (O_1063,N_8960,N_8271);
and UO_1064 (O_1064,N_7838,N_7834);
nand UO_1065 (O_1065,N_9556,N_8325);
and UO_1066 (O_1066,N_9570,N_9464);
or UO_1067 (O_1067,N_8739,N_7971);
or UO_1068 (O_1068,N_8321,N_9206);
nor UO_1069 (O_1069,N_9263,N_8984);
nor UO_1070 (O_1070,N_7633,N_9517);
nor UO_1071 (O_1071,N_9407,N_9007);
or UO_1072 (O_1072,N_9377,N_8515);
nor UO_1073 (O_1073,N_7866,N_9107);
or UO_1074 (O_1074,N_7650,N_9618);
and UO_1075 (O_1075,N_8211,N_8599);
xor UO_1076 (O_1076,N_8782,N_8623);
xnor UO_1077 (O_1077,N_7513,N_8341);
and UO_1078 (O_1078,N_7696,N_8595);
nand UO_1079 (O_1079,N_8889,N_8618);
nand UO_1080 (O_1080,N_9704,N_8188);
and UO_1081 (O_1081,N_8116,N_9778);
xnor UO_1082 (O_1082,N_8964,N_7809);
xnor UO_1083 (O_1083,N_8827,N_7899);
xor UO_1084 (O_1084,N_8411,N_9935);
or UO_1085 (O_1085,N_9947,N_9122);
nand UO_1086 (O_1086,N_8945,N_7937);
nand UO_1087 (O_1087,N_8270,N_8028);
nor UO_1088 (O_1088,N_9090,N_9651);
nor UO_1089 (O_1089,N_9054,N_8065);
or UO_1090 (O_1090,N_7743,N_7901);
nor UO_1091 (O_1091,N_9602,N_9882);
xnor UO_1092 (O_1092,N_9604,N_7894);
nor UO_1093 (O_1093,N_8501,N_9466);
nand UO_1094 (O_1094,N_9320,N_9596);
and UO_1095 (O_1095,N_7511,N_9099);
or UO_1096 (O_1096,N_8146,N_8570);
xnor UO_1097 (O_1097,N_9346,N_8467);
nand UO_1098 (O_1098,N_9557,N_9900);
or UO_1099 (O_1099,N_7829,N_9681);
nor UO_1100 (O_1100,N_9663,N_9437);
or UO_1101 (O_1101,N_8780,N_9307);
nand UO_1102 (O_1102,N_9918,N_9299);
nor UO_1103 (O_1103,N_9370,N_8592);
xor UO_1104 (O_1104,N_9518,N_8380);
nand UO_1105 (O_1105,N_9699,N_7844);
nor UO_1106 (O_1106,N_9739,N_8636);
nand UO_1107 (O_1107,N_7574,N_8921);
and UO_1108 (O_1108,N_9901,N_7957);
nand UO_1109 (O_1109,N_7661,N_9520);
xnor UO_1110 (O_1110,N_9101,N_8093);
and UO_1111 (O_1111,N_7768,N_9473);
or UO_1112 (O_1112,N_9134,N_8025);
xnor UO_1113 (O_1113,N_7642,N_7679);
nor UO_1114 (O_1114,N_8289,N_9481);
and UO_1115 (O_1115,N_8394,N_8177);
and UO_1116 (O_1116,N_7692,N_9995);
nor UO_1117 (O_1117,N_7857,N_7815);
and UO_1118 (O_1118,N_9891,N_8463);
nor UO_1119 (O_1119,N_8641,N_8372);
and UO_1120 (O_1120,N_8976,N_7740);
xnor UO_1121 (O_1121,N_9966,N_9951);
or UO_1122 (O_1122,N_9894,N_9623);
nor UO_1123 (O_1123,N_9745,N_9434);
nand UO_1124 (O_1124,N_9754,N_9371);
xnor UO_1125 (O_1125,N_8436,N_8071);
nand UO_1126 (O_1126,N_9659,N_8415);
xnor UO_1127 (O_1127,N_7507,N_8450);
and UO_1128 (O_1128,N_7665,N_8580);
or UO_1129 (O_1129,N_9642,N_9907);
nand UO_1130 (O_1130,N_7853,N_9721);
nor UO_1131 (O_1131,N_7527,N_9467);
nor UO_1132 (O_1132,N_7712,N_8421);
nor UO_1133 (O_1133,N_9416,N_9538);
or UO_1134 (O_1134,N_8936,N_9906);
xnor UO_1135 (O_1135,N_8017,N_8552);
nand UO_1136 (O_1136,N_7803,N_9221);
or UO_1137 (O_1137,N_7772,N_9247);
xnor UO_1138 (O_1138,N_8313,N_8502);
and UO_1139 (O_1139,N_9449,N_9648);
nor UO_1140 (O_1140,N_9165,N_8799);
and UO_1141 (O_1141,N_8039,N_7640);
and UO_1142 (O_1142,N_9948,N_8820);
xor UO_1143 (O_1143,N_9629,N_7746);
nor UO_1144 (O_1144,N_8635,N_8414);
nor UO_1145 (O_1145,N_9326,N_8445);
or UO_1146 (O_1146,N_8518,N_8854);
or UO_1147 (O_1147,N_7843,N_7824);
xor UO_1148 (O_1148,N_7886,N_9083);
or UO_1149 (O_1149,N_8091,N_8189);
or UO_1150 (O_1150,N_7539,N_9698);
and UO_1151 (O_1151,N_9442,N_9163);
xnor UO_1152 (O_1152,N_7902,N_8352);
or UO_1153 (O_1153,N_8656,N_8537);
xnor UO_1154 (O_1154,N_9184,N_7535);
nor UO_1155 (O_1155,N_8044,N_8661);
xor UO_1156 (O_1156,N_7613,N_8466);
or UO_1157 (O_1157,N_9059,N_9747);
xnor UO_1158 (O_1158,N_9228,N_9089);
nor UO_1159 (O_1159,N_7781,N_8740);
and UO_1160 (O_1160,N_8485,N_9817);
or UO_1161 (O_1161,N_9707,N_9241);
or UO_1162 (O_1162,N_9779,N_8707);
nand UO_1163 (O_1163,N_7601,N_9048);
nand UO_1164 (O_1164,N_7940,N_7706);
and UO_1165 (O_1165,N_8645,N_9639);
xnor UO_1166 (O_1166,N_8774,N_8957);
xor UO_1167 (O_1167,N_8312,N_9512);
and UO_1168 (O_1168,N_8885,N_9887);
or UO_1169 (O_1169,N_9561,N_9872);
and UO_1170 (O_1170,N_8056,N_7547);
or UO_1171 (O_1171,N_7502,N_7590);
nand UO_1172 (O_1172,N_9711,N_9603);
or UO_1173 (O_1173,N_8701,N_8465);
nand UO_1174 (O_1174,N_9316,N_9128);
nor UO_1175 (O_1175,N_7562,N_8133);
and UO_1176 (O_1176,N_8168,N_9772);
and UO_1177 (O_1177,N_9854,N_9283);
nand UO_1178 (O_1178,N_7874,N_7900);
nor UO_1179 (O_1179,N_8078,N_8916);
and UO_1180 (O_1180,N_8969,N_8922);
and UO_1181 (O_1181,N_7758,N_8031);
nand UO_1182 (O_1182,N_9425,N_9666);
nand UO_1183 (O_1183,N_9412,N_9849);
nor UO_1184 (O_1184,N_8098,N_8282);
nand UO_1185 (O_1185,N_9762,N_9696);
nand UO_1186 (O_1186,N_7622,N_7864);
nand UO_1187 (O_1187,N_9459,N_7967);
and UO_1188 (O_1188,N_9749,N_9730);
or UO_1189 (O_1189,N_8767,N_8983);
and UO_1190 (O_1190,N_9964,N_7713);
or UO_1191 (O_1191,N_8222,N_9802);
xor UO_1192 (O_1192,N_7698,N_8185);
or UO_1193 (O_1193,N_8747,N_9631);
and UO_1194 (O_1194,N_9497,N_9254);
nand UO_1195 (O_1195,N_8193,N_9693);
or UO_1196 (O_1196,N_8319,N_7979);
nor UO_1197 (O_1197,N_7804,N_8948);
nor UO_1198 (O_1198,N_9955,N_8131);
xnor UO_1199 (O_1199,N_9223,N_8413);
nor UO_1200 (O_1200,N_8968,N_7512);
nand UO_1201 (O_1201,N_9344,N_9113);
or UO_1202 (O_1202,N_9086,N_8109);
and UO_1203 (O_1203,N_7856,N_9369);
or UO_1204 (O_1204,N_8235,N_8207);
nor UO_1205 (O_1205,N_8398,N_8644);
and UO_1206 (O_1206,N_9354,N_8647);
and UO_1207 (O_1207,N_9262,N_8507);
or UO_1208 (O_1208,N_8735,N_9571);
or UO_1209 (O_1209,N_9217,N_8451);
or UO_1210 (O_1210,N_9735,N_9549);
and UO_1211 (O_1211,N_9893,N_9417);
nor UO_1212 (O_1212,N_7606,N_8441);
nand UO_1213 (O_1213,N_8204,N_7593);
nand UO_1214 (O_1214,N_8136,N_8634);
nand UO_1215 (O_1215,N_9915,N_9061);
xnor UO_1216 (O_1216,N_8334,N_9532);
xnor UO_1217 (O_1217,N_7961,N_8743);
nor UO_1218 (O_1218,N_7660,N_8746);
nand UO_1219 (O_1219,N_8912,N_9238);
nand UO_1220 (O_1220,N_9130,N_9932);
xor UO_1221 (O_1221,N_7672,N_7767);
xnor UO_1222 (O_1222,N_9862,N_9734);
nor UO_1223 (O_1223,N_7873,N_8058);
nor UO_1224 (O_1224,N_8075,N_9261);
nor UO_1225 (O_1225,N_9423,N_9656);
xnor UO_1226 (O_1226,N_9474,N_7603);
and UO_1227 (O_1227,N_8046,N_8822);
and UO_1228 (O_1228,N_9676,N_9986);
nor UO_1229 (O_1229,N_7814,N_9843);
xor UO_1230 (O_1230,N_7898,N_9522);
nand UO_1231 (O_1231,N_8816,N_8333);
nor UO_1232 (O_1232,N_8336,N_9477);
and UO_1233 (O_1233,N_8329,N_9805);
xor UO_1234 (O_1234,N_9812,N_9265);
nand UO_1235 (O_1235,N_9690,N_7988);
and UO_1236 (O_1236,N_8349,N_8390);
xnor UO_1237 (O_1237,N_8274,N_7550);
or UO_1238 (O_1238,N_7947,N_8675);
and UO_1239 (O_1239,N_8527,N_8804);
nand UO_1240 (O_1240,N_8356,N_8452);
nand UO_1241 (O_1241,N_8057,N_9572);
xor UO_1242 (O_1242,N_8790,N_7905);
xor UO_1243 (O_1243,N_9080,N_8749);
or UO_1244 (O_1244,N_9465,N_9537);
or UO_1245 (O_1245,N_8253,N_9155);
xnor UO_1246 (O_1246,N_9850,N_8684);
xor UO_1247 (O_1247,N_8214,N_7529);
nand UO_1248 (O_1248,N_8258,N_8628);
and UO_1249 (O_1249,N_9120,N_8293);
or UO_1250 (O_1250,N_8588,N_9607);
xnor UO_1251 (O_1251,N_9894,N_8196);
nand UO_1252 (O_1252,N_8573,N_9865);
xnor UO_1253 (O_1253,N_9147,N_8164);
and UO_1254 (O_1254,N_8816,N_9983);
or UO_1255 (O_1255,N_8779,N_7919);
and UO_1256 (O_1256,N_7694,N_8172);
and UO_1257 (O_1257,N_8377,N_7828);
and UO_1258 (O_1258,N_9340,N_9745);
nor UO_1259 (O_1259,N_9997,N_8219);
xor UO_1260 (O_1260,N_9640,N_9497);
nand UO_1261 (O_1261,N_8318,N_8384);
nor UO_1262 (O_1262,N_9921,N_7703);
and UO_1263 (O_1263,N_9747,N_9953);
and UO_1264 (O_1264,N_8338,N_8402);
or UO_1265 (O_1265,N_8539,N_8609);
nor UO_1266 (O_1266,N_8863,N_8762);
nand UO_1267 (O_1267,N_9717,N_8243);
nor UO_1268 (O_1268,N_7816,N_8653);
and UO_1269 (O_1269,N_7578,N_8178);
xnor UO_1270 (O_1270,N_8548,N_8058);
or UO_1271 (O_1271,N_7777,N_9302);
and UO_1272 (O_1272,N_8150,N_8428);
or UO_1273 (O_1273,N_8156,N_7667);
nand UO_1274 (O_1274,N_8935,N_9835);
or UO_1275 (O_1275,N_9280,N_9522);
nor UO_1276 (O_1276,N_9727,N_7742);
and UO_1277 (O_1277,N_9125,N_7629);
nor UO_1278 (O_1278,N_9169,N_9451);
nand UO_1279 (O_1279,N_9899,N_7538);
nor UO_1280 (O_1280,N_7862,N_9899);
nand UO_1281 (O_1281,N_9691,N_7747);
and UO_1282 (O_1282,N_9024,N_9143);
and UO_1283 (O_1283,N_7505,N_9029);
nand UO_1284 (O_1284,N_7773,N_8478);
nor UO_1285 (O_1285,N_7648,N_8217);
xnor UO_1286 (O_1286,N_9403,N_8739);
and UO_1287 (O_1287,N_7873,N_9265);
nor UO_1288 (O_1288,N_7791,N_9791);
nand UO_1289 (O_1289,N_7913,N_8068);
and UO_1290 (O_1290,N_8752,N_8646);
or UO_1291 (O_1291,N_8166,N_7782);
xor UO_1292 (O_1292,N_8864,N_9390);
nand UO_1293 (O_1293,N_9687,N_9343);
or UO_1294 (O_1294,N_9847,N_8194);
nor UO_1295 (O_1295,N_8762,N_9645);
nor UO_1296 (O_1296,N_8489,N_7750);
nor UO_1297 (O_1297,N_9771,N_8838);
or UO_1298 (O_1298,N_8289,N_8744);
and UO_1299 (O_1299,N_8972,N_8687);
nor UO_1300 (O_1300,N_9925,N_9677);
nor UO_1301 (O_1301,N_8893,N_8574);
xor UO_1302 (O_1302,N_8837,N_8819);
or UO_1303 (O_1303,N_9970,N_9512);
nor UO_1304 (O_1304,N_9391,N_8608);
or UO_1305 (O_1305,N_8095,N_7519);
and UO_1306 (O_1306,N_7799,N_9542);
nor UO_1307 (O_1307,N_7955,N_9256);
xor UO_1308 (O_1308,N_8035,N_9331);
or UO_1309 (O_1309,N_7751,N_7558);
nand UO_1310 (O_1310,N_9717,N_9561);
nand UO_1311 (O_1311,N_9965,N_9985);
xor UO_1312 (O_1312,N_9066,N_8995);
or UO_1313 (O_1313,N_9367,N_9457);
or UO_1314 (O_1314,N_9191,N_8952);
xnor UO_1315 (O_1315,N_7678,N_9049);
xnor UO_1316 (O_1316,N_9295,N_9142);
xnor UO_1317 (O_1317,N_9950,N_9713);
nor UO_1318 (O_1318,N_9747,N_9721);
nand UO_1319 (O_1319,N_9089,N_8227);
xor UO_1320 (O_1320,N_9393,N_9667);
nor UO_1321 (O_1321,N_9937,N_8123);
and UO_1322 (O_1322,N_9193,N_9950);
nor UO_1323 (O_1323,N_9490,N_9445);
nand UO_1324 (O_1324,N_8103,N_8785);
or UO_1325 (O_1325,N_9784,N_9692);
nor UO_1326 (O_1326,N_8121,N_8137);
or UO_1327 (O_1327,N_9606,N_8346);
and UO_1328 (O_1328,N_9826,N_8427);
xor UO_1329 (O_1329,N_7965,N_9331);
xor UO_1330 (O_1330,N_8249,N_8839);
xnor UO_1331 (O_1331,N_9182,N_9644);
nand UO_1332 (O_1332,N_8572,N_9653);
xnor UO_1333 (O_1333,N_7672,N_7663);
nor UO_1334 (O_1334,N_9076,N_9027);
nor UO_1335 (O_1335,N_9104,N_8903);
and UO_1336 (O_1336,N_8973,N_9665);
nor UO_1337 (O_1337,N_9530,N_9736);
or UO_1338 (O_1338,N_8416,N_8586);
or UO_1339 (O_1339,N_9191,N_9450);
nand UO_1340 (O_1340,N_8036,N_9918);
nand UO_1341 (O_1341,N_7814,N_8358);
and UO_1342 (O_1342,N_9892,N_8952);
nand UO_1343 (O_1343,N_8386,N_7713);
or UO_1344 (O_1344,N_8079,N_9331);
and UO_1345 (O_1345,N_8121,N_9393);
xor UO_1346 (O_1346,N_9981,N_8786);
nand UO_1347 (O_1347,N_8636,N_7636);
or UO_1348 (O_1348,N_8605,N_8785);
xnor UO_1349 (O_1349,N_9823,N_9718);
xor UO_1350 (O_1350,N_8440,N_8163);
xnor UO_1351 (O_1351,N_7774,N_8547);
xor UO_1352 (O_1352,N_8118,N_9705);
and UO_1353 (O_1353,N_7894,N_9940);
or UO_1354 (O_1354,N_9078,N_7986);
xnor UO_1355 (O_1355,N_9998,N_8917);
nor UO_1356 (O_1356,N_9902,N_7971);
nor UO_1357 (O_1357,N_8784,N_8636);
xor UO_1358 (O_1358,N_9777,N_7707);
and UO_1359 (O_1359,N_7635,N_7701);
xor UO_1360 (O_1360,N_8553,N_7772);
or UO_1361 (O_1361,N_9361,N_9100);
nor UO_1362 (O_1362,N_7827,N_9027);
nor UO_1363 (O_1363,N_8424,N_9897);
nor UO_1364 (O_1364,N_9265,N_8138);
and UO_1365 (O_1365,N_7993,N_7633);
nand UO_1366 (O_1366,N_8899,N_9656);
xor UO_1367 (O_1367,N_7952,N_8721);
nand UO_1368 (O_1368,N_9062,N_8439);
nor UO_1369 (O_1369,N_9800,N_9070);
xor UO_1370 (O_1370,N_7598,N_8663);
xnor UO_1371 (O_1371,N_7719,N_8553);
nand UO_1372 (O_1372,N_8295,N_8691);
and UO_1373 (O_1373,N_8290,N_8838);
and UO_1374 (O_1374,N_9617,N_9702);
nor UO_1375 (O_1375,N_7942,N_7936);
nand UO_1376 (O_1376,N_8148,N_8548);
or UO_1377 (O_1377,N_8136,N_9882);
and UO_1378 (O_1378,N_7866,N_8074);
or UO_1379 (O_1379,N_8061,N_7793);
xor UO_1380 (O_1380,N_8023,N_8680);
nor UO_1381 (O_1381,N_8599,N_7503);
nor UO_1382 (O_1382,N_9488,N_9119);
nand UO_1383 (O_1383,N_9995,N_9525);
nor UO_1384 (O_1384,N_9187,N_9469);
xnor UO_1385 (O_1385,N_8478,N_8477);
nor UO_1386 (O_1386,N_9126,N_8261);
or UO_1387 (O_1387,N_8932,N_9424);
or UO_1388 (O_1388,N_9637,N_9214);
xnor UO_1389 (O_1389,N_8761,N_7824);
and UO_1390 (O_1390,N_9720,N_9938);
and UO_1391 (O_1391,N_7864,N_8527);
nor UO_1392 (O_1392,N_8990,N_7844);
xnor UO_1393 (O_1393,N_8296,N_7633);
and UO_1394 (O_1394,N_7770,N_8914);
nand UO_1395 (O_1395,N_8475,N_8993);
or UO_1396 (O_1396,N_8173,N_8592);
or UO_1397 (O_1397,N_7870,N_9565);
nor UO_1398 (O_1398,N_8331,N_8063);
nor UO_1399 (O_1399,N_8109,N_9508);
xor UO_1400 (O_1400,N_9840,N_8539);
nand UO_1401 (O_1401,N_8300,N_9589);
xor UO_1402 (O_1402,N_8212,N_8194);
nand UO_1403 (O_1403,N_9727,N_9502);
nor UO_1404 (O_1404,N_9952,N_8624);
and UO_1405 (O_1405,N_9403,N_9892);
or UO_1406 (O_1406,N_9154,N_9067);
nor UO_1407 (O_1407,N_9862,N_9106);
nand UO_1408 (O_1408,N_9809,N_7509);
and UO_1409 (O_1409,N_9367,N_9396);
nand UO_1410 (O_1410,N_7503,N_8992);
nand UO_1411 (O_1411,N_8813,N_9252);
nand UO_1412 (O_1412,N_8199,N_8727);
or UO_1413 (O_1413,N_9061,N_9085);
xnor UO_1414 (O_1414,N_8752,N_8236);
xnor UO_1415 (O_1415,N_7604,N_9796);
or UO_1416 (O_1416,N_7834,N_7875);
xor UO_1417 (O_1417,N_8997,N_8402);
and UO_1418 (O_1418,N_8636,N_8655);
nand UO_1419 (O_1419,N_8849,N_9246);
nand UO_1420 (O_1420,N_7615,N_8472);
and UO_1421 (O_1421,N_8801,N_7759);
nand UO_1422 (O_1422,N_9722,N_7676);
nand UO_1423 (O_1423,N_8051,N_8402);
nand UO_1424 (O_1424,N_8989,N_8752);
nor UO_1425 (O_1425,N_8321,N_8802);
nand UO_1426 (O_1426,N_9160,N_8889);
and UO_1427 (O_1427,N_9683,N_9182);
and UO_1428 (O_1428,N_8494,N_8178);
and UO_1429 (O_1429,N_8633,N_7743);
and UO_1430 (O_1430,N_9748,N_8493);
or UO_1431 (O_1431,N_7960,N_7756);
xor UO_1432 (O_1432,N_9129,N_9064);
and UO_1433 (O_1433,N_9795,N_8882);
and UO_1434 (O_1434,N_9780,N_9329);
or UO_1435 (O_1435,N_7630,N_8760);
nand UO_1436 (O_1436,N_8077,N_7844);
and UO_1437 (O_1437,N_7719,N_8671);
or UO_1438 (O_1438,N_9300,N_7986);
or UO_1439 (O_1439,N_8448,N_8580);
or UO_1440 (O_1440,N_7584,N_7577);
xnor UO_1441 (O_1441,N_9653,N_9422);
nand UO_1442 (O_1442,N_8853,N_7589);
and UO_1443 (O_1443,N_8382,N_9074);
nand UO_1444 (O_1444,N_8329,N_8556);
nor UO_1445 (O_1445,N_8396,N_8064);
or UO_1446 (O_1446,N_9041,N_9446);
and UO_1447 (O_1447,N_9544,N_9647);
and UO_1448 (O_1448,N_8382,N_7862);
nor UO_1449 (O_1449,N_9065,N_7852);
or UO_1450 (O_1450,N_9163,N_8272);
nor UO_1451 (O_1451,N_9275,N_8321);
and UO_1452 (O_1452,N_7773,N_9911);
nor UO_1453 (O_1453,N_9804,N_7925);
nor UO_1454 (O_1454,N_8498,N_8582);
nand UO_1455 (O_1455,N_7538,N_9051);
xnor UO_1456 (O_1456,N_9033,N_8254);
nand UO_1457 (O_1457,N_7758,N_9355);
nor UO_1458 (O_1458,N_7523,N_9421);
or UO_1459 (O_1459,N_7657,N_9435);
xor UO_1460 (O_1460,N_8902,N_7799);
nand UO_1461 (O_1461,N_7771,N_7652);
nand UO_1462 (O_1462,N_8242,N_8417);
xnor UO_1463 (O_1463,N_8087,N_7798);
or UO_1464 (O_1464,N_8927,N_9604);
or UO_1465 (O_1465,N_8778,N_9608);
nor UO_1466 (O_1466,N_8942,N_7883);
xor UO_1467 (O_1467,N_8496,N_9921);
or UO_1468 (O_1468,N_9685,N_9860);
xnor UO_1469 (O_1469,N_8810,N_8431);
and UO_1470 (O_1470,N_9288,N_9984);
nor UO_1471 (O_1471,N_7666,N_8464);
or UO_1472 (O_1472,N_9242,N_9072);
xor UO_1473 (O_1473,N_7687,N_8196);
and UO_1474 (O_1474,N_8403,N_8962);
nor UO_1475 (O_1475,N_9260,N_9976);
nor UO_1476 (O_1476,N_7884,N_9989);
or UO_1477 (O_1477,N_8374,N_7605);
nand UO_1478 (O_1478,N_9961,N_7609);
or UO_1479 (O_1479,N_8916,N_9081);
or UO_1480 (O_1480,N_7504,N_9118);
nor UO_1481 (O_1481,N_7629,N_9823);
and UO_1482 (O_1482,N_8468,N_9315);
and UO_1483 (O_1483,N_8822,N_9930);
or UO_1484 (O_1484,N_9059,N_9173);
or UO_1485 (O_1485,N_8339,N_8817);
xnor UO_1486 (O_1486,N_8783,N_8422);
nor UO_1487 (O_1487,N_9686,N_9556);
or UO_1488 (O_1488,N_7592,N_7513);
nor UO_1489 (O_1489,N_8071,N_9871);
or UO_1490 (O_1490,N_7664,N_7982);
xnor UO_1491 (O_1491,N_8546,N_9721);
nor UO_1492 (O_1492,N_8172,N_8649);
nor UO_1493 (O_1493,N_8759,N_7815);
and UO_1494 (O_1494,N_7967,N_8479);
and UO_1495 (O_1495,N_9005,N_8229);
and UO_1496 (O_1496,N_9314,N_7924);
nand UO_1497 (O_1497,N_8411,N_8280);
and UO_1498 (O_1498,N_9468,N_7734);
xor UO_1499 (O_1499,N_8436,N_8350);
endmodule