module basic_750_5000_1000_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_24,In_496);
nor U1 (N_1,In_95,In_114);
xnor U2 (N_2,In_579,In_376);
nor U3 (N_3,In_655,In_200);
nor U4 (N_4,In_585,In_662);
or U5 (N_5,In_122,In_718);
nor U6 (N_6,In_423,In_635);
or U7 (N_7,In_168,In_648);
or U8 (N_8,In_76,In_747);
nor U9 (N_9,In_347,In_1);
and U10 (N_10,In_152,In_279);
and U11 (N_11,In_393,In_64);
xnor U12 (N_12,In_36,In_333);
xor U13 (N_13,In_621,In_177);
nor U14 (N_14,In_241,In_437);
or U15 (N_15,In_238,In_69);
and U16 (N_16,In_10,In_120);
xnor U17 (N_17,In_361,In_464);
and U18 (N_18,In_391,In_703);
and U19 (N_19,In_426,In_429);
xnor U20 (N_20,In_11,In_22);
nor U21 (N_21,In_631,In_477);
nor U22 (N_22,In_296,In_157);
and U23 (N_23,In_615,In_276);
and U24 (N_24,In_127,In_206);
xnor U25 (N_25,In_215,In_328);
xnor U26 (N_26,In_102,In_711);
nor U27 (N_27,In_715,In_189);
xnor U28 (N_28,In_85,In_399);
xnor U29 (N_29,In_123,In_449);
or U30 (N_30,In_367,In_534);
xor U31 (N_31,In_281,In_269);
or U32 (N_32,In_691,In_560);
nand U33 (N_33,In_21,In_221);
and U34 (N_34,In_724,In_664);
nor U35 (N_35,In_596,In_125);
xnor U36 (N_36,In_388,In_167);
nand U37 (N_37,In_197,In_435);
xnor U38 (N_38,In_681,In_278);
or U39 (N_39,In_433,In_143);
nand U40 (N_40,In_96,In_667);
and U41 (N_41,In_366,In_561);
or U42 (N_42,In_663,In_587);
xor U43 (N_43,In_682,In_4);
or U44 (N_44,In_352,In_522);
xor U45 (N_45,In_29,In_387);
nand U46 (N_46,In_533,In_503);
or U47 (N_47,In_484,In_458);
or U48 (N_48,In_285,In_68);
nor U49 (N_49,In_583,In_306);
nand U50 (N_50,In_12,In_271);
or U51 (N_51,In_629,In_566);
or U52 (N_52,In_686,In_551);
nand U53 (N_53,In_268,In_636);
xor U54 (N_54,In_705,In_644);
or U55 (N_55,In_625,In_498);
nand U56 (N_56,In_160,In_670);
or U57 (N_57,In_385,In_599);
nor U58 (N_58,In_372,In_505);
or U59 (N_59,In_94,In_148);
nor U60 (N_60,In_603,In_267);
nor U61 (N_61,In_612,In_698);
and U62 (N_62,In_424,In_547);
xor U63 (N_63,In_33,In_440);
nor U64 (N_64,In_744,In_261);
or U65 (N_65,In_730,In_39);
nand U66 (N_66,In_702,In_256);
nor U67 (N_67,In_677,In_617);
or U68 (N_68,In_77,In_719);
xor U69 (N_69,In_444,In_133);
nor U70 (N_70,In_526,In_601);
xnor U71 (N_71,In_332,In_700);
or U72 (N_72,In_312,In_574);
or U73 (N_73,In_161,In_548);
and U74 (N_74,In_354,In_90);
or U75 (N_75,In_380,In_51);
nand U76 (N_76,In_473,In_78);
nor U77 (N_77,In_340,In_604);
nand U78 (N_78,In_84,In_89);
or U79 (N_79,In_214,In_371);
nor U80 (N_80,In_497,In_334);
nand U81 (N_81,In_243,In_519);
xor U82 (N_82,In_112,In_182);
or U83 (N_83,In_139,In_493);
nand U84 (N_84,In_582,In_618);
and U85 (N_85,In_362,In_186);
nand U86 (N_86,In_672,In_417);
xor U87 (N_87,In_729,In_156);
nand U88 (N_88,In_485,In_309);
and U89 (N_89,In_198,In_145);
and U90 (N_90,In_460,In_209);
nor U91 (N_91,In_442,In_502);
and U92 (N_92,In_27,In_301);
and U93 (N_93,In_746,In_652);
or U94 (N_94,In_263,In_174);
xnor U95 (N_95,In_646,In_556);
nand U96 (N_96,In_171,In_568);
nor U97 (N_97,In_250,In_48);
xor U98 (N_98,In_410,In_588);
xnor U99 (N_99,In_723,In_557);
nor U100 (N_100,In_97,N_53);
and U101 (N_101,N_25,N_41);
xnor U102 (N_102,In_654,In_419);
xnor U103 (N_103,In_420,In_331);
xor U104 (N_104,In_181,In_126);
nand U105 (N_105,In_313,In_398);
or U106 (N_106,In_20,In_675);
nor U107 (N_107,N_5,In_541);
nor U108 (N_108,N_81,In_740);
xnor U109 (N_109,In_219,In_297);
nor U110 (N_110,In_273,In_343);
xnor U111 (N_111,N_36,In_111);
or U112 (N_112,In_222,N_24);
xor U113 (N_113,In_188,N_0);
and U114 (N_114,N_50,In_247);
and U115 (N_115,In_627,In_733);
and U116 (N_116,In_734,In_359);
xor U117 (N_117,In_514,In_100);
nor U118 (N_118,N_21,In_315);
nor U119 (N_119,N_79,In_725);
nor U120 (N_120,In_213,In_592);
xor U121 (N_121,In_205,In_71);
and U122 (N_122,In_350,In_735);
and U123 (N_123,In_300,In_580);
xnor U124 (N_124,N_94,In_314);
nor U125 (N_125,In_134,In_290);
xor U126 (N_126,In_693,In_369);
or U127 (N_127,N_16,N_51);
nor U128 (N_128,In_244,N_60);
nand U129 (N_129,In_465,N_97);
or U130 (N_130,In_228,In_259);
nor U131 (N_131,In_607,In_82);
nor U132 (N_132,In_402,In_469);
nor U133 (N_133,In_248,In_706);
nand U134 (N_134,In_235,N_70);
xnor U135 (N_135,N_71,N_23);
and U136 (N_136,In_397,N_88);
nor U137 (N_137,In_620,In_738);
nand U138 (N_138,In_748,In_395);
and U139 (N_139,N_67,In_633);
nor U140 (N_140,In_119,In_728);
nor U141 (N_141,In_147,In_688);
or U142 (N_142,In_418,In_598);
or U143 (N_143,In_572,In_683);
and U144 (N_144,In_479,In_637);
nand U145 (N_145,In_517,In_216);
or U146 (N_146,In_710,In_478);
nand U147 (N_147,In_737,In_491);
xor U148 (N_148,In_378,In_379);
xnor U149 (N_149,N_73,N_12);
or U150 (N_150,In_310,In_258);
nand U151 (N_151,In_431,In_645);
nor U152 (N_152,In_195,N_59);
xnor U153 (N_153,N_9,In_470);
xor U154 (N_154,In_689,In_146);
or U155 (N_155,In_55,In_443);
or U156 (N_156,In_613,In_344);
or U157 (N_157,In_499,In_712);
and U158 (N_158,In_628,In_660);
or U159 (N_159,N_63,In_50);
nor U160 (N_160,In_377,In_179);
or U161 (N_161,In_428,In_292);
nor U162 (N_162,N_17,In_448);
and U163 (N_163,In_708,N_26);
and U164 (N_164,In_321,In_394);
nor U165 (N_165,In_294,In_230);
and U166 (N_166,In_150,In_9);
and U167 (N_167,In_511,In_743);
nand U168 (N_168,In_529,In_674);
nand U169 (N_169,In_208,In_446);
and U170 (N_170,In_600,In_62);
nor U171 (N_171,In_293,In_8);
xnor U172 (N_172,In_202,In_2);
and U173 (N_173,N_90,In_25);
nand U174 (N_174,N_10,In_178);
or U175 (N_175,In_573,N_87);
or U176 (N_176,In_638,In_158);
nand U177 (N_177,In_121,In_454);
xnor U178 (N_178,In_404,In_468);
or U179 (N_179,In_83,In_282);
or U180 (N_180,In_162,In_166);
or U181 (N_181,In_389,In_709);
xor U182 (N_182,In_327,In_501);
nand U183 (N_183,In_357,In_647);
nor U184 (N_184,In_384,In_254);
nor U185 (N_185,In_322,In_16);
xnor U186 (N_186,In_319,In_155);
nor U187 (N_187,In_521,In_461);
or U188 (N_188,In_260,In_690);
or U189 (N_189,In_425,In_323);
or U190 (N_190,In_184,N_39);
or U191 (N_191,N_6,In_575);
nor U192 (N_192,N_75,N_76);
and U193 (N_193,In_91,In_581);
nand U194 (N_194,In_642,N_48);
xnor U195 (N_195,In_661,In_317);
nand U196 (N_196,In_272,In_251);
or U197 (N_197,N_78,In_236);
nor U198 (N_198,N_46,In_353);
xnor U199 (N_199,N_28,In_237);
nand U200 (N_200,N_133,In_164);
xor U201 (N_201,N_102,N_2);
nand U202 (N_202,N_158,In_624);
or U203 (N_203,In_298,N_86);
xor U204 (N_204,N_135,In_577);
nor U205 (N_205,In_467,In_274);
and U206 (N_206,In_515,In_539);
nand U207 (N_207,In_203,In_109);
xor U208 (N_208,In_679,N_145);
or U209 (N_209,N_138,In_584);
and U210 (N_210,N_136,In_509);
xor U211 (N_211,N_159,In_640);
nand U212 (N_212,N_22,In_318);
nand U213 (N_213,In_373,In_749);
nor U214 (N_214,In_54,In_459);
or U215 (N_215,N_99,In_14);
or U216 (N_216,In_540,N_113);
nand U217 (N_217,In_481,In_360);
nor U218 (N_218,In_500,N_15);
xnor U219 (N_219,N_171,In_563);
xor U220 (N_220,N_84,In_531);
xnor U221 (N_221,In_530,In_490);
and U222 (N_222,In_28,In_597);
nor U223 (N_223,In_714,N_196);
nand U224 (N_224,In_717,In_452);
or U225 (N_225,N_144,In_80);
nor U226 (N_226,In_41,In_320);
nor U227 (N_227,In_193,N_176);
and U228 (N_228,In_427,In_349);
and U229 (N_229,In_245,In_665);
xor U230 (N_230,In_538,N_197);
nand U231 (N_231,In_694,In_308);
and U232 (N_232,In_239,In_673);
nand U233 (N_233,N_33,In_255);
nor U234 (N_234,In_716,In_187);
xor U235 (N_235,N_77,In_422);
or U236 (N_236,In_98,In_0);
xnor U237 (N_237,N_111,In_475);
and U238 (N_238,In_136,N_92);
nor U239 (N_239,In_669,In_436);
and U240 (N_240,In_450,N_146);
xnor U241 (N_241,In_535,In_508);
nor U242 (N_242,In_34,In_159);
nor U243 (N_243,In_512,In_288);
or U244 (N_244,N_89,In_138);
xnor U245 (N_245,In_47,N_30);
nand U246 (N_246,In_396,In_546);
nand U247 (N_247,In_336,In_257);
and U248 (N_248,In_558,In_18);
nor U249 (N_249,In_565,N_147);
xor U250 (N_250,N_31,In_52);
nand U251 (N_251,In_616,N_143);
nand U252 (N_252,In_564,In_544);
or U253 (N_253,N_115,In_741);
nand U254 (N_254,N_98,In_576);
nor U255 (N_255,In_40,In_345);
or U256 (N_256,N_20,In_742);
nor U257 (N_257,N_19,In_386);
xor U258 (N_258,N_172,In_286);
nor U259 (N_259,N_69,In_365);
xnor U260 (N_260,In_264,N_120);
nand U261 (N_261,In_571,In_233);
or U262 (N_262,N_139,In_57);
and U263 (N_263,N_168,In_439);
xnor U264 (N_264,In_381,N_104);
nor U265 (N_265,In_270,In_593);
nand U266 (N_266,In_676,In_370);
nor U267 (N_267,In_651,In_110);
nand U268 (N_268,In_523,In_720);
nand U269 (N_269,N_126,In_390);
xor U270 (N_270,In_229,In_170);
or U271 (N_271,In_262,In_45);
xnor U272 (N_272,N_61,In_65);
xor U273 (N_273,In_494,In_329);
nor U274 (N_274,In_400,In_207);
or U275 (N_275,In_364,In_441);
nor U276 (N_276,In_639,In_731);
nor U277 (N_277,In_619,In_545);
or U278 (N_278,In_602,N_38);
nor U279 (N_279,N_198,In_346);
nor U280 (N_280,In_226,In_103);
and U281 (N_281,N_184,N_192);
xnor U282 (N_282,In_56,In_697);
and U283 (N_283,In_144,In_32);
nand U284 (N_284,In_480,In_445);
xnor U285 (N_285,N_177,In_630);
and U286 (N_286,N_72,In_299);
nor U287 (N_287,N_13,In_727);
nand U288 (N_288,N_167,In_252);
or U289 (N_289,In_295,N_42);
xnor U290 (N_290,N_124,In_153);
or U291 (N_291,N_175,N_85);
or U292 (N_292,N_153,In_552);
nand U293 (N_293,In_185,N_44);
nand U294 (N_294,In_524,N_45);
xor U295 (N_295,N_150,In_659);
nor U296 (N_296,In_289,In_72);
and U297 (N_297,In_92,In_374);
and U298 (N_298,In_283,In_223);
nand U299 (N_299,In_23,N_160);
and U300 (N_300,In_492,In_430);
nor U301 (N_301,N_29,In_43);
and U302 (N_302,N_93,In_456);
xnor U303 (N_303,In_457,In_721);
xnor U304 (N_304,In_307,N_261);
or U305 (N_305,N_246,In_46);
nor U306 (N_306,N_66,N_278);
nor U307 (N_307,In_31,In_337);
or U308 (N_308,In_190,In_93);
nor U309 (N_309,N_211,In_108);
xor U310 (N_310,In_405,N_166);
and U311 (N_311,N_83,In_438);
nand U312 (N_312,In_474,N_117);
or U313 (N_313,In_53,N_274);
or U314 (N_314,N_47,In_7);
or U315 (N_315,N_258,N_239);
or U316 (N_316,N_154,In_699);
nor U317 (N_317,N_82,In_30);
xnor U318 (N_318,N_269,N_125);
and U319 (N_319,In_507,N_188);
nor U320 (N_320,N_164,In_658);
and U321 (N_321,In_192,In_634);
nor U322 (N_322,In_671,In_104);
nor U323 (N_323,In_348,In_382);
xor U324 (N_324,N_242,In_284);
nand U325 (N_325,N_18,N_286);
nor U326 (N_326,In_506,N_1);
and U327 (N_327,In_489,In_113);
and U328 (N_328,In_586,N_249);
nor U329 (N_329,N_265,N_244);
nor U330 (N_330,N_245,N_11);
nor U331 (N_331,N_37,In_305);
and U332 (N_332,N_226,N_230);
and U333 (N_333,In_246,N_56);
or U334 (N_334,N_199,In_49);
xor U335 (N_335,N_200,In_356);
and U336 (N_336,In_632,N_212);
xor U337 (N_337,N_141,In_19);
and U338 (N_338,In_38,In_623);
xnor U339 (N_339,In_176,N_225);
and U340 (N_340,In_101,In_154);
nand U341 (N_341,N_137,N_259);
or U342 (N_342,N_279,In_218);
or U343 (N_343,In_684,In_518);
xor U344 (N_344,In_657,In_696);
nand U345 (N_345,In_453,In_463);
xnor U346 (N_346,N_263,N_287);
nand U347 (N_347,In_668,In_105);
or U348 (N_348,N_96,In_513);
xnor U349 (N_349,In_211,In_118);
nor U350 (N_350,In_392,N_290);
xnor U351 (N_351,In_42,In_537);
nand U352 (N_352,In_471,In_61);
or U353 (N_353,N_299,In_86);
or U354 (N_354,In_324,In_415);
and U355 (N_355,N_224,N_110);
nand U356 (N_356,In_525,In_401);
nand U357 (N_357,In_736,In_726);
xnor U358 (N_358,N_251,In_482);
nor U359 (N_359,In_253,In_363);
xor U360 (N_360,N_202,In_641);
xnor U361 (N_361,N_194,N_223);
nor U362 (N_362,N_221,In_74);
and U363 (N_363,N_169,N_100);
xor U364 (N_364,N_227,N_285);
nand U365 (N_365,N_178,In_653);
or U366 (N_366,In_131,N_254);
or U367 (N_367,In_70,N_49);
nor U368 (N_368,N_151,In_291);
xor U369 (N_369,In_17,In_549);
or U370 (N_370,N_91,In_416);
nor U371 (N_371,In_73,N_165);
nand U372 (N_372,N_101,In_212);
and U373 (N_373,N_204,In_680);
xor U374 (N_374,N_255,N_119);
xor U375 (N_375,In_687,N_74);
and U376 (N_376,N_27,N_182);
and U377 (N_377,In_466,In_60);
and U378 (N_378,N_121,N_268);
nor U379 (N_379,In_649,In_304);
and U380 (N_380,In_67,In_210);
xor U381 (N_381,In_149,N_229);
or U382 (N_382,N_213,N_173);
and U383 (N_383,In_358,In_342);
and U384 (N_384,N_40,N_284);
and U385 (N_385,In_594,In_326);
or U386 (N_386,N_253,In_383);
nor U387 (N_387,In_194,In_462);
and U388 (N_388,N_114,In_739);
xor U389 (N_389,N_216,N_209);
and U390 (N_390,In_707,In_81);
or U391 (N_391,In_63,N_106);
nor U392 (N_392,N_203,N_233);
xnor U393 (N_393,N_4,In_234);
nor U394 (N_394,In_87,In_472);
and U395 (N_395,In_614,In_407);
and U396 (N_396,N_130,N_118);
nor U397 (N_397,N_272,In_220);
xnor U398 (N_398,N_220,N_162);
nor U399 (N_399,In_589,In_58);
nand U400 (N_400,N_122,In_590);
and U401 (N_401,N_381,N_257);
xor U402 (N_402,In_341,N_127);
nor U403 (N_403,In_406,In_495);
nand U404 (N_404,N_306,N_382);
nor U405 (N_405,In_570,N_250);
nand U406 (N_406,In_595,N_264);
nor U407 (N_407,N_252,In_142);
nor U408 (N_408,N_148,N_237);
and U409 (N_409,N_132,In_559);
nor U410 (N_410,In_231,N_366);
nor U411 (N_411,N_310,N_3);
xor U412 (N_412,In_510,N_95);
nor U413 (N_413,In_330,N_330);
nor U414 (N_414,N_383,In_191);
nand U415 (N_415,N_387,N_329);
nor U416 (N_416,N_368,In_129);
and U417 (N_417,N_14,N_58);
or U418 (N_418,N_8,N_300);
or U419 (N_419,In_745,N_241);
nand U420 (N_420,N_345,N_236);
nor U421 (N_421,In_695,In_550);
or U422 (N_422,N_103,In_303);
or U423 (N_423,N_195,N_363);
or U424 (N_424,N_65,N_354);
nor U425 (N_425,N_57,In_339);
or U426 (N_426,In_280,N_358);
xnor U427 (N_427,N_396,N_332);
nor U428 (N_428,N_340,N_315);
nand U429 (N_429,N_108,N_334);
nor U430 (N_430,N_314,In_163);
or U431 (N_431,N_276,N_327);
and U432 (N_432,In_232,In_66);
xnor U433 (N_433,N_301,In_451);
nand U434 (N_434,N_302,N_292);
nor U435 (N_435,N_398,N_222);
and U436 (N_436,In_240,In_606);
nand U437 (N_437,In_701,N_228);
and U438 (N_438,N_107,N_238);
nor U439 (N_439,In_183,In_555);
and U440 (N_440,N_336,In_553);
and U441 (N_441,N_325,N_350);
and U442 (N_442,In_224,In_408);
nor U443 (N_443,N_281,N_185);
or U444 (N_444,In_542,N_123);
nand U445 (N_445,In_486,N_392);
and U446 (N_446,N_273,In_578);
or U447 (N_447,In_335,N_189);
and U448 (N_448,In_527,N_134);
and U449 (N_449,In_137,N_347);
xor U450 (N_450,In_609,In_713);
nor U451 (N_451,In_106,N_378);
or U452 (N_452,N_361,N_397);
and U453 (N_453,N_109,N_357);
nand U454 (N_454,N_112,N_105);
or U455 (N_455,In_591,In_528);
and U456 (N_456,N_320,In_227);
nand U457 (N_457,N_293,In_685);
and U458 (N_458,N_296,N_260);
nand U459 (N_459,N_288,In_562);
or U460 (N_460,N_232,N_142);
nor U461 (N_461,N_355,N_393);
and U462 (N_462,In_455,In_554);
and U463 (N_463,In_75,N_215);
and U464 (N_464,In_277,In_59);
and U465 (N_465,N_389,N_64);
or U466 (N_466,N_342,N_348);
nand U467 (N_467,N_283,N_266);
and U468 (N_468,N_304,In_421);
nand U469 (N_469,In_249,N_156);
nand U470 (N_470,N_262,N_179);
or U471 (N_471,In_704,In_117);
nand U472 (N_472,In_516,N_186);
or U473 (N_473,In_569,N_360);
and U474 (N_474,In_355,N_312);
and U475 (N_475,N_234,N_370);
nand U476 (N_476,In_128,N_384);
and U477 (N_477,N_386,N_68);
nor U478 (N_478,In_37,In_151);
and U479 (N_479,N_271,N_337);
and U480 (N_480,N_149,N_240);
xnor U481 (N_481,In_666,N_206);
or U482 (N_482,In_532,In_650);
nor U483 (N_483,In_504,N_128);
xnor U484 (N_484,N_54,N_309);
and U485 (N_485,In_622,In_180);
xor U486 (N_486,In_169,N_359);
nand U487 (N_487,In_325,N_322);
xnor U488 (N_488,N_181,In_225);
and U489 (N_489,N_328,N_210);
xnor U490 (N_490,In_5,In_626);
or U491 (N_491,In_656,In_165);
nor U492 (N_492,N_339,In_351);
nand U493 (N_493,In_316,N_338);
nor U494 (N_494,N_218,In_88);
nand U495 (N_495,In_487,N_362);
or U496 (N_496,N_380,N_344);
or U497 (N_497,N_391,In_199);
and U498 (N_498,N_80,N_289);
nor U499 (N_499,N_207,In_79);
nand U500 (N_500,N_372,In_266);
xor U501 (N_501,N_441,N_493);
nor U502 (N_502,N_307,In_432);
xnor U503 (N_503,N_62,N_356);
or U504 (N_504,N_410,N_129);
nand U505 (N_505,N_457,N_463);
nor U506 (N_506,In_140,In_132);
nand U507 (N_507,N_219,N_416);
nor U508 (N_508,N_313,In_26);
nor U509 (N_509,In_414,N_388);
nor U510 (N_510,N_399,N_294);
or U511 (N_511,N_433,In_412);
or U512 (N_512,N_321,N_427);
nor U513 (N_513,N_445,N_485);
nand U514 (N_514,N_367,N_498);
xor U515 (N_515,N_495,N_152);
and U516 (N_516,N_174,N_163);
and U517 (N_517,In_368,N_235);
and U518 (N_518,In_275,N_419);
or U519 (N_519,N_319,N_373);
nand U520 (N_520,N_407,In_175);
and U521 (N_521,N_365,N_180);
or U522 (N_522,N_484,N_418);
xnor U523 (N_523,N_465,In_567);
nor U524 (N_524,In_172,N_461);
xor U525 (N_525,N_295,In_434);
nand U526 (N_526,N_217,N_401);
and U527 (N_527,N_455,N_424);
xor U528 (N_528,N_420,N_297);
nand U529 (N_529,N_324,N_435);
nor U530 (N_530,In_115,N_458);
or U531 (N_531,N_476,N_415);
or U532 (N_532,N_402,In_483);
xor U533 (N_533,N_375,N_448);
nor U534 (N_534,N_349,N_187);
nor U535 (N_535,N_335,In_116);
nand U536 (N_536,In_13,In_643);
or U537 (N_537,In_536,N_479);
xor U538 (N_538,N_477,N_369);
or U539 (N_539,N_499,N_472);
nor U540 (N_540,N_446,In_44);
and U541 (N_541,In_375,N_406);
nor U542 (N_542,N_376,N_417);
nor U543 (N_543,N_277,N_183);
nor U544 (N_544,N_413,N_459);
nand U545 (N_545,N_483,In_543);
and U546 (N_546,N_374,In_409);
and U547 (N_547,N_492,N_341);
and U548 (N_548,N_468,In_413);
or U549 (N_549,N_323,N_32);
or U550 (N_550,N_496,N_161);
xor U551 (N_551,N_403,In_722);
nand U552 (N_552,N_478,In_35);
xor U553 (N_553,N_390,N_308);
or U554 (N_554,N_43,In_265);
and U555 (N_555,N_7,N_425);
nor U556 (N_556,N_469,N_298);
and U557 (N_557,In_135,N_491);
nand U558 (N_558,N_275,N_414);
and U559 (N_559,In_6,In_217);
and U560 (N_560,In_3,N_201);
or U561 (N_561,N_466,N_405);
xnor U562 (N_562,N_473,N_411);
nor U563 (N_563,In_411,N_432);
nor U564 (N_564,N_352,N_450);
nor U565 (N_565,N_474,In_520);
nand U566 (N_566,N_467,N_475);
nand U567 (N_567,N_434,N_426);
xnor U568 (N_568,N_243,N_205);
and U569 (N_569,N_303,N_482);
nand U570 (N_570,In_692,In_15);
or U571 (N_571,N_346,N_379);
or U572 (N_572,N_247,N_460);
nor U573 (N_573,N_462,In_201);
nor U574 (N_574,N_436,N_55);
xnor U575 (N_575,N_423,N_439);
or U576 (N_576,N_452,N_140);
nand U577 (N_577,In_311,N_193);
or U578 (N_578,In_338,N_451);
nand U579 (N_579,N_282,In_196);
nand U580 (N_580,N_170,N_480);
nand U581 (N_581,N_422,N_494);
or U582 (N_582,N_214,N_421);
nor U583 (N_583,N_305,In_447);
nor U584 (N_584,N_116,N_431);
and U585 (N_585,N_34,N_442);
and U586 (N_586,N_443,N_444);
and U587 (N_587,N_489,N_437);
xor U588 (N_588,N_394,N_280);
or U589 (N_589,N_471,N_248);
or U590 (N_590,N_464,N_430);
xnor U591 (N_591,N_481,N_311);
xor U592 (N_592,N_333,N_404);
nor U593 (N_593,N_488,In_204);
or U594 (N_594,N_456,N_316);
or U595 (N_595,N_191,N_35);
and U596 (N_596,N_270,N_429);
or U597 (N_597,N_400,N_131);
xor U598 (N_598,In_610,In_403);
and U599 (N_599,In_173,N_438);
nor U600 (N_600,N_515,N_517);
nor U601 (N_601,N_505,N_533);
and U602 (N_602,N_518,N_537);
or U603 (N_603,N_267,N_509);
nor U604 (N_604,N_497,N_502);
and U605 (N_605,N_584,N_590);
nand U606 (N_606,N_371,N_291);
nand U607 (N_607,N_528,N_507);
or U608 (N_608,N_532,N_155);
nor U609 (N_609,N_583,N_587);
or U610 (N_610,N_557,N_351);
or U611 (N_611,N_560,N_526);
and U612 (N_612,N_556,N_412);
nand U613 (N_613,N_545,N_501);
nor U614 (N_614,N_364,N_231);
or U615 (N_615,N_552,N_520);
and U616 (N_616,In_476,N_486);
nand U617 (N_617,N_52,N_551);
or U618 (N_618,In_678,N_454);
nor U619 (N_619,N_487,N_599);
and U620 (N_620,N_554,N_588);
or U621 (N_621,N_508,In_287);
nor U622 (N_622,N_385,N_593);
xnor U623 (N_623,N_563,N_585);
nor U624 (N_624,N_566,In_99);
or U625 (N_625,N_589,N_565);
nor U626 (N_626,In_242,N_256);
nand U627 (N_627,N_535,N_544);
nand U628 (N_628,N_574,N_577);
nor U629 (N_629,N_572,N_546);
xnor U630 (N_630,N_470,N_447);
xor U631 (N_631,N_428,N_536);
nor U632 (N_632,N_208,In_107);
xnor U633 (N_633,N_449,N_569);
nor U634 (N_634,N_564,N_512);
and U635 (N_635,N_558,In_611);
nor U636 (N_636,N_539,N_504);
or U637 (N_637,N_561,N_595);
nand U638 (N_638,N_562,N_519);
nor U639 (N_639,N_567,N_594);
or U640 (N_640,N_506,N_453);
nor U641 (N_641,N_503,N_576);
nor U642 (N_642,N_550,N_591);
or U643 (N_643,In_302,N_513);
xnor U644 (N_644,N_331,N_580);
and U645 (N_645,N_409,N_317);
nand U646 (N_646,N_573,N_559);
nor U647 (N_647,N_395,N_527);
and U648 (N_648,N_579,N_524);
nand U649 (N_649,N_326,N_514);
or U650 (N_650,N_440,N_523);
xor U651 (N_651,N_547,N_343);
and U652 (N_652,N_522,In_608);
and U653 (N_653,N_353,N_490);
nand U654 (N_654,N_571,N_553);
nor U655 (N_655,N_568,In_130);
nor U656 (N_656,N_521,N_530);
or U657 (N_657,N_529,N_540);
or U658 (N_658,N_549,N_596);
and U659 (N_659,N_582,N_510);
xnor U660 (N_660,N_500,N_531);
or U661 (N_661,N_575,N_408);
xnor U662 (N_662,N_516,N_555);
nand U663 (N_663,In_141,N_511);
nor U664 (N_664,N_586,N_541);
or U665 (N_665,N_157,N_190);
and U666 (N_666,N_548,N_542);
nor U667 (N_667,N_592,N_598);
or U668 (N_668,N_525,In_732);
or U669 (N_669,In_124,N_578);
nor U670 (N_670,N_597,In_605);
nand U671 (N_671,N_534,N_543);
nor U672 (N_672,N_318,N_377);
nor U673 (N_673,In_488,N_570);
or U674 (N_674,N_581,N_538);
nand U675 (N_675,N_569,In_302);
or U676 (N_676,N_504,N_525);
and U677 (N_677,N_542,N_554);
nand U678 (N_678,N_395,N_497);
and U679 (N_679,N_470,In_107);
or U680 (N_680,N_589,N_447);
and U681 (N_681,N_524,N_440);
xor U682 (N_682,N_343,N_552);
nand U683 (N_683,In_476,N_554);
and U684 (N_684,N_559,N_486);
nand U685 (N_685,N_502,N_371);
and U686 (N_686,N_578,N_540);
and U687 (N_687,N_534,N_157);
or U688 (N_688,N_574,N_208);
or U689 (N_689,In_488,N_534);
nor U690 (N_690,N_539,N_564);
xnor U691 (N_691,N_515,N_534);
or U692 (N_692,N_577,N_507);
xnor U693 (N_693,N_584,N_554);
or U694 (N_694,N_541,N_506);
nand U695 (N_695,N_562,N_598);
and U696 (N_696,N_553,N_597);
nand U697 (N_697,N_544,N_256);
or U698 (N_698,N_521,In_732);
xnor U699 (N_699,N_583,N_516);
and U700 (N_700,N_679,N_628);
and U701 (N_701,N_618,N_687);
and U702 (N_702,N_600,N_665);
nand U703 (N_703,N_623,N_682);
xnor U704 (N_704,N_672,N_694);
nand U705 (N_705,N_678,N_627);
or U706 (N_706,N_673,N_692);
nand U707 (N_707,N_622,N_651);
xnor U708 (N_708,N_609,N_698);
and U709 (N_709,N_624,N_656);
nor U710 (N_710,N_680,N_607);
xor U711 (N_711,N_625,N_630);
nor U712 (N_712,N_615,N_657);
nand U713 (N_713,N_614,N_668);
nand U714 (N_714,N_638,N_636);
and U715 (N_715,N_635,N_613);
and U716 (N_716,N_670,N_608);
nor U717 (N_717,N_642,N_641);
and U718 (N_718,N_683,N_617);
or U719 (N_719,N_691,N_659);
nand U720 (N_720,N_626,N_681);
xor U721 (N_721,N_649,N_652);
nand U722 (N_722,N_629,N_640);
xnor U723 (N_723,N_660,N_633);
and U724 (N_724,N_695,N_654);
and U725 (N_725,N_612,N_690);
or U726 (N_726,N_655,N_699);
nor U727 (N_727,N_647,N_646);
xnor U728 (N_728,N_664,N_685);
xnor U729 (N_729,N_643,N_604);
and U730 (N_730,N_666,N_697);
and U731 (N_731,N_661,N_639);
xnor U732 (N_732,N_601,N_603);
xor U733 (N_733,N_620,N_644);
and U734 (N_734,N_631,N_650);
nor U735 (N_735,N_610,N_663);
nand U736 (N_736,N_696,N_653);
nor U737 (N_737,N_619,N_634);
and U738 (N_738,N_667,N_669);
nand U739 (N_739,N_606,N_676);
nor U740 (N_740,N_688,N_611);
nor U741 (N_741,N_616,N_632);
or U742 (N_742,N_671,N_602);
xor U743 (N_743,N_675,N_689);
nor U744 (N_744,N_677,N_662);
or U745 (N_745,N_621,N_637);
or U746 (N_746,N_645,N_605);
xor U747 (N_747,N_686,N_674);
nor U748 (N_748,N_684,N_693);
or U749 (N_749,N_648,N_658);
or U750 (N_750,N_682,N_641);
nand U751 (N_751,N_670,N_682);
nand U752 (N_752,N_690,N_644);
xor U753 (N_753,N_687,N_604);
xor U754 (N_754,N_625,N_615);
nor U755 (N_755,N_627,N_605);
or U756 (N_756,N_636,N_668);
nand U757 (N_757,N_691,N_681);
nor U758 (N_758,N_633,N_666);
xor U759 (N_759,N_688,N_628);
xor U760 (N_760,N_612,N_692);
and U761 (N_761,N_649,N_658);
xnor U762 (N_762,N_641,N_616);
nor U763 (N_763,N_644,N_673);
nor U764 (N_764,N_605,N_688);
and U765 (N_765,N_683,N_618);
or U766 (N_766,N_691,N_671);
nor U767 (N_767,N_674,N_668);
nor U768 (N_768,N_635,N_631);
nor U769 (N_769,N_691,N_664);
nand U770 (N_770,N_631,N_654);
xor U771 (N_771,N_610,N_673);
or U772 (N_772,N_623,N_663);
xor U773 (N_773,N_650,N_610);
xor U774 (N_774,N_685,N_643);
nor U775 (N_775,N_640,N_667);
nor U776 (N_776,N_612,N_656);
or U777 (N_777,N_678,N_635);
xnor U778 (N_778,N_669,N_664);
or U779 (N_779,N_601,N_690);
or U780 (N_780,N_610,N_658);
or U781 (N_781,N_650,N_680);
and U782 (N_782,N_610,N_668);
and U783 (N_783,N_692,N_614);
nor U784 (N_784,N_621,N_668);
xnor U785 (N_785,N_629,N_613);
xnor U786 (N_786,N_679,N_668);
and U787 (N_787,N_678,N_618);
xor U788 (N_788,N_659,N_617);
and U789 (N_789,N_618,N_635);
and U790 (N_790,N_629,N_682);
nand U791 (N_791,N_617,N_612);
nand U792 (N_792,N_633,N_622);
and U793 (N_793,N_614,N_629);
xor U794 (N_794,N_671,N_666);
or U795 (N_795,N_686,N_675);
or U796 (N_796,N_667,N_650);
nor U797 (N_797,N_696,N_608);
nor U798 (N_798,N_644,N_693);
nand U799 (N_799,N_650,N_693);
nand U800 (N_800,N_704,N_719);
or U801 (N_801,N_769,N_757);
or U802 (N_802,N_773,N_727);
nor U803 (N_803,N_706,N_708);
nand U804 (N_804,N_754,N_718);
nand U805 (N_805,N_794,N_790);
and U806 (N_806,N_796,N_781);
nor U807 (N_807,N_797,N_793);
or U808 (N_808,N_785,N_783);
nor U809 (N_809,N_782,N_721);
xnor U810 (N_810,N_733,N_788);
nor U811 (N_811,N_759,N_760);
and U812 (N_812,N_772,N_776);
nor U813 (N_813,N_724,N_770);
nand U814 (N_814,N_710,N_712);
and U815 (N_815,N_742,N_778);
or U816 (N_816,N_745,N_777);
nor U817 (N_817,N_743,N_722);
xnor U818 (N_818,N_736,N_780);
xor U819 (N_819,N_730,N_746);
nand U820 (N_820,N_753,N_735);
and U821 (N_821,N_734,N_707);
or U822 (N_822,N_747,N_786);
xnor U823 (N_823,N_729,N_715);
and U824 (N_824,N_728,N_779);
and U825 (N_825,N_752,N_762);
nand U826 (N_826,N_768,N_787);
xnor U827 (N_827,N_720,N_774);
or U828 (N_828,N_748,N_744);
nand U829 (N_829,N_767,N_761);
nor U830 (N_830,N_758,N_765);
nor U831 (N_831,N_741,N_750);
or U832 (N_832,N_725,N_732);
nand U833 (N_833,N_701,N_763);
nand U834 (N_834,N_751,N_700);
xor U835 (N_835,N_749,N_795);
nand U836 (N_836,N_705,N_731);
or U837 (N_837,N_723,N_766);
nand U838 (N_838,N_702,N_775);
xnor U839 (N_839,N_756,N_717);
nor U840 (N_840,N_791,N_792);
and U841 (N_841,N_771,N_739);
nand U842 (N_842,N_709,N_737);
nand U843 (N_843,N_799,N_798);
and U844 (N_844,N_784,N_755);
and U845 (N_845,N_714,N_703);
nor U846 (N_846,N_738,N_716);
or U847 (N_847,N_764,N_711);
or U848 (N_848,N_726,N_740);
and U849 (N_849,N_789,N_713);
xor U850 (N_850,N_788,N_780);
nor U851 (N_851,N_768,N_722);
or U852 (N_852,N_767,N_781);
nor U853 (N_853,N_706,N_796);
and U854 (N_854,N_700,N_705);
and U855 (N_855,N_796,N_729);
or U856 (N_856,N_792,N_706);
nand U857 (N_857,N_754,N_721);
nand U858 (N_858,N_732,N_755);
nand U859 (N_859,N_749,N_700);
nand U860 (N_860,N_771,N_781);
and U861 (N_861,N_756,N_791);
and U862 (N_862,N_729,N_762);
and U863 (N_863,N_793,N_777);
nor U864 (N_864,N_714,N_735);
nor U865 (N_865,N_725,N_748);
nand U866 (N_866,N_773,N_747);
nor U867 (N_867,N_706,N_740);
nor U868 (N_868,N_725,N_790);
xor U869 (N_869,N_740,N_765);
nor U870 (N_870,N_776,N_771);
and U871 (N_871,N_702,N_786);
and U872 (N_872,N_724,N_736);
nand U873 (N_873,N_713,N_719);
or U874 (N_874,N_786,N_763);
or U875 (N_875,N_779,N_741);
nor U876 (N_876,N_781,N_714);
and U877 (N_877,N_747,N_791);
xnor U878 (N_878,N_747,N_732);
nand U879 (N_879,N_731,N_727);
xnor U880 (N_880,N_735,N_785);
nor U881 (N_881,N_784,N_797);
xor U882 (N_882,N_763,N_764);
nand U883 (N_883,N_787,N_712);
xor U884 (N_884,N_785,N_799);
and U885 (N_885,N_721,N_737);
nor U886 (N_886,N_786,N_751);
nor U887 (N_887,N_777,N_797);
and U888 (N_888,N_782,N_702);
nand U889 (N_889,N_772,N_783);
xnor U890 (N_890,N_702,N_758);
and U891 (N_891,N_747,N_709);
xor U892 (N_892,N_758,N_708);
nand U893 (N_893,N_788,N_717);
nand U894 (N_894,N_730,N_760);
or U895 (N_895,N_753,N_779);
nor U896 (N_896,N_711,N_772);
and U897 (N_897,N_777,N_764);
nand U898 (N_898,N_738,N_729);
xnor U899 (N_899,N_727,N_706);
xnor U900 (N_900,N_826,N_811);
xor U901 (N_901,N_804,N_848);
xnor U902 (N_902,N_899,N_810);
nand U903 (N_903,N_877,N_830);
xnor U904 (N_904,N_854,N_871);
nand U905 (N_905,N_829,N_824);
or U906 (N_906,N_890,N_894);
nand U907 (N_907,N_858,N_815);
xnor U908 (N_908,N_878,N_885);
or U909 (N_909,N_816,N_880);
xor U910 (N_910,N_835,N_882);
or U911 (N_911,N_813,N_841);
nand U912 (N_912,N_853,N_801);
or U913 (N_913,N_846,N_812);
xnor U914 (N_914,N_895,N_837);
and U915 (N_915,N_870,N_827);
nor U916 (N_916,N_807,N_856);
or U917 (N_917,N_867,N_819);
xnor U918 (N_918,N_891,N_898);
xnor U919 (N_919,N_863,N_893);
nor U920 (N_920,N_874,N_820);
or U921 (N_921,N_821,N_855);
and U922 (N_922,N_873,N_888);
xor U923 (N_923,N_845,N_865);
and U924 (N_924,N_886,N_809);
xnor U925 (N_925,N_866,N_875);
xnor U926 (N_926,N_857,N_862);
and U927 (N_927,N_800,N_818);
or U928 (N_928,N_817,N_850);
nor U929 (N_929,N_842,N_897);
or U930 (N_930,N_802,N_831);
nand U931 (N_931,N_822,N_843);
nor U932 (N_932,N_840,N_806);
xor U933 (N_933,N_864,N_814);
nor U934 (N_934,N_838,N_808);
or U935 (N_935,N_889,N_896);
nor U936 (N_936,N_847,N_860);
nand U937 (N_937,N_828,N_872);
and U938 (N_938,N_832,N_892);
or U939 (N_939,N_839,N_849);
nand U940 (N_940,N_879,N_861);
nor U941 (N_941,N_834,N_881);
xnor U942 (N_942,N_833,N_883);
nand U943 (N_943,N_876,N_823);
and U944 (N_944,N_805,N_887);
nand U945 (N_945,N_852,N_836);
xnor U946 (N_946,N_825,N_869);
and U947 (N_947,N_851,N_884);
nand U948 (N_948,N_868,N_859);
and U949 (N_949,N_844,N_803);
or U950 (N_950,N_894,N_893);
and U951 (N_951,N_836,N_879);
and U952 (N_952,N_873,N_880);
nor U953 (N_953,N_878,N_803);
xor U954 (N_954,N_831,N_832);
and U955 (N_955,N_828,N_890);
nor U956 (N_956,N_849,N_816);
or U957 (N_957,N_855,N_837);
or U958 (N_958,N_831,N_805);
and U959 (N_959,N_885,N_805);
nor U960 (N_960,N_881,N_817);
or U961 (N_961,N_850,N_828);
nand U962 (N_962,N_885,N_844);
or U963 (N_963,N_876,N_897);
and U964 (N_964,N_833,N_899);
nor U965 (N_965,N_856,N_881);
xor U966 (N_966,N_879,N_806);
and U967 (N_967,N_829,N_804);
nand U968 (N_968,N_885,N_803);
or U969 (N_969,N_899,N_848);
xnor U970 (N_970,N_889,N_825);
xor U971 (N_971,N_812,N_882);
or U972 (N_972,N_874,N_891);
xor U973 (N_973,N_807,N_851);
nor U974 (N_974,N_811,N_880);
xnor U975 (N_975,N_841,N_889);
nor U976 (N_976,N_873,N_802);
or U977 (N_977,N_896,N_856);
or U978 (N_978,N_881,N_829);
nand U979 (N_979,N_852,N_884);
or U980 (N_980,N_887,N_854);
or U981 (N_981,N_835,N_870);
nor U982 (N_982,N_893,N_840);
xnor U983 (N_983,N_831,N_827);
or U984 (N_984,N_859,N_827);
xor U985 (N_985,N_857,N_895);
nor U986 (N_986,N_891,N_838);
nand U987 (N_987,N_860,N_800);
nor U988 (N_988,N_893,N_888);
nor U989 (N_989,N_856,N_878);
or U990 (N_990,N_858,N_897);
nor U991 (N_991,N_896,N_843);
or U992 (N_992,N_880,N_866);
and U993 (N_993,N_853,N_856);
and U994 (N_994,N_890,N_820);
or U995 (N_995,N_862,N_874);
xnor U996 (N_996,N_866,N_809);
nand U997 (N_997,N_855,N_836);
nand U998 (N_998,N_834,N_887);
nand U999 (N_999,N_894,N_838);
nand U1000 (N_1000,N_992,N_973);
or U1001 (N_1001,N_943,N_921);
or U1002 (N_1002,N_966,N_914);
or U1003 (N_1003,N_977,N_938);
or U1004 (N_1004,N_906,N_956);
and U1005 (N_1005,N_912,N_922);
nor U1006 (N_1006,N_945,N_994);
or U1007 (N_1007,N_931,N_975);
nor U1008 (N_1008,N_930,N_902);
or U1009 (N_1009,N_952,N_988);
nand U1010 (N_1010,N_911,N_927);
xnor U1011 (N_1011,N_995,N_909);
xnor U1012 (N_1012,N_913,N_946);
nor U1013 (N_1013,N_993,N_900);
and U1014 (N_1014,N_949,N_939);
and U1015 (N_1015,N_967,N_915);
and U1016 (N_1016,N_903,N_942);
nor U1017 (N_1017,N_983,N_934);
nor U1018 (N_1018,N_971,N_985);
nand U1019 (N_1019,N_987,N_964);
or U1020 (N_1020,N_959,N_996);
nand U1021 (N_1021,N_910,N_950);
nand U1022 (N_1022,N_955,N_908);
xor U1023 (N_1023,N_974,N_907);
or U1024 (N_1024,N_986,N_941);
or U1025 (N_1025,N_976,N_933);
nand U1026 (N_1026,N_961,N_929);
or U1027 (N_1027,N_953,N_969);
xor U1028 (N_1028,N_924,N_965);
nor U1029 (N_1029,N_984,N_937);
nor U1030 (N_1030,N_999,N_962);
or U1031 (N_1031,N_936,N_919);
xnor U1032 (N_1032,N_917,N_970);
and U1033 (N_1033,N_947,N_905);
nor U1034 (N_1034,N_923,N_957);
and U1035 (N_1035,N_979,N_997);
xor U1036 (N_1036,N_972,N_920);
or U1037 (N_1037,N_940,N_998);
and U1038 (N_1038,N_948,N_916);
xor U1039 (N_1039,N_960,N_932);
and U1040 (N_1040,N_963,N_926);
xor U1041 (N_1041,N_918,N_944);
or U1042 (N_1042,N_990,N_951);
and U1043 (N_1043,N_901,N_978);
xor U1044 (N_1044,N_991,N_928);
and U1045 (N_1045,N_981,N_958);
nor U1046 (N_1046,N_935,N_954);
xor U1047 (N_1047,N_968,N_980);
nand U1048 (N_1048,N_982,N_989);
nor U1049 (N_1049,N_925,N_904);
nand U1050 (N_1050,N_965,N_910);
and U1051 (N_1051,N_971,N_975);
xor U1052 (N_1052,N_946,N_961);
or U1053 (N_1053,N_913,N_928);
or U1054 (N_1054,N_997,N_924);
or U1055 (N_1055,N_977,N_993);
xnor U1056 (N_1056,N_901,N_981);
or U1057 (N_1057,N_991,N_906);
nor U1058 (N_1058,N_954,N_924);
nor U1059 (N_1059,N_958,N_930);
or U1060 (N_1060,N_935,N_951);
nand U1061 (N_1061,N_960,N_971);
nand U1062 (N_1062,N_958,N_901);
nand U1063 (N_1063,N_998,N_994);
xnor U1064 (N_1064,N_983,N_972);
and U1065 (N_1065,N_980,N_967);
nor U1066 (N_1066,N_917,N_944);
xnor U1067 (N_1067,N_920,N_983);
and U1068 (N_1068,N_932,N_969);
or U1069 (N_1069,N_957,N_924);
nand U1070 (N_1070,N_940,N_914);
nor U1071 (N_1071,N_955,N_909);
xor U1072 (N_1072,N_934,N_966);
xnor U1073 (N_1073,N_971,N_944);
xnor U1074 (N_1074,N_938,N_978);
xor U1075 (N_1075,N_970,N_939);
xor U1076 (N_1076,N_972,N_927);
or U1077 (N_1077,N_999,N_936);
nand U1078 (N_1078,N_920,N_919);
or U1079 (N_1079,N_976,N_996);
nand U1080 (N_1080,N_984,N_947);
and U1081 (N_1081,N_937,N_913);
nand U1082 (N_1082,N_945,N_978);
and U1083 (N_1083,N_964,N_974);
nor U1084 (N_1084,N_943,N_998);
or U1085 (N_1085,N_950,N_937);
nor U1086 (N_1086,N_904,N_910);
xnor U1087 (N_1087,N_950,N_903);
xnor U1088 (N_1088,N_987,N_949);
nor U1089 (N_1089,N_915,N_906);
or U1090 (N_1090,N_904,N_978);
or U1091 (N_1091,N_993,N_965);
or U1092 (N_1092,N_998,N_915);
or U1093 (N_1093,N_941,N_902);
xor U1094 (N_1094,N_985,N_915);
nor U1095 (N_1095,N_905,N_953);
nand U1096 (N_1096,N_905,N_935);
nand U1097 (N_1097,N_972,N_903);
nor U1098 (N_1098,N_923,N_993);
or U1099 (N_1099,N_909,N_921);
or U1100 (N_1100,N_1058,N_1056);
nor U1101 (N_1101,N_1097,N_1034);
nor U1102 (N_1102,N_1008,N_1043);
nand U1103 (N_1103,N_1082,N_1032);
nand U1104 (N_1104,N_1071,N_1072);
nor U1105 (N_1105,N_1054,N_1070);
xnor U1106 (N_1106,N_1083,N_1010);
or U1107 (N_1107,N_1003,N_1027);
xor U1108 (N_1108,N_1041,N_1051);
nor U1109 (N_1109,N_1020,N_1085);
nor U1110 (N_1110,N_1060,N_1087);
xor U1111 (N_1111,N_1007,N_1049);
nand U1112 (N_1112,N_1013,N_1055);
nor U1113 (N_1113,N_1098,N_1042);
nor U1114 (N_1114,N_1053,N_1033);
nand U1115 (N_1115,N_1036,N_1014);
nor U1116 (N_1116,N_1073,N_1066);
or U1117 (N_1117,N_1018,N_1057);
and U1118 (N_1118,N_1040,N_1099);
nor U1119 (N_1119,N_1076,N_1001);
nand U1120 (N_1120,N_1022,N_1062);
or U1121 (N_1121,N_1024,N_1045);
nor U1122 (N_1122,N_1074,N_1038);
nand U1123 (N_1123,N_1086,N_1088);
and U1124 (N_1124,N_1080,N_1005);
or U1125 (N_1125,N_1046,N_1048);
nand U1126 (N_1126,N_1090,N_1016);
xnor U1127 (N_1127,N_1019,N_1079);
and U1128 (N_1128,N_1077,N_1068);
xnor U1129 (N_1129,N_1026,N_1065);
nor U1130 (N_1130,N_1091,N_1067);
and U1131 (N_1131,N_1030,N_1061);
or U1132 (N_1132,N_1064,N_1006);
nor U1133 (N_1133,N_1028,N_1063);
xnor U1134 (N_1134,N_1017,N_1047);
or U1135 (N_1135,N_1012,N_1095);
and U1136 (N_1136,N_1052,N_1029);
nand U1137 (N_1137,N_1035,N_1011);
nand U1138 (N_1138,N_1015,N_1094);
nor U1139 (N_1139,N_1092,N_1069);
or U1140 (N_1140,N_1002,N_1089);
nand U1141 (N_1141,N_1081,N_1009);
xnor U1142 (N_1142,N_1000,N_1025);
or U1143 (N_1143,N_1004,N_1050);
or U1144 (N_1144,N_1021,N_1075);
nor U1145 (N_1145,N_1039,N_1031);
nand U1146 (N_1146,N_1037,N_1096);
nor U1147 (N_1147,N_1093,N_1084);
and U1148 (N_1148,N_1078,N_1023);
xnor U1149 (N_1149,N_1059,N_1044);
or U1150 (N_1150,N_1015,N_1062);
nor U1151 (N_1151,N_1003,N_1065);
nor U1152 (N_1152,N_1051,N_1037);
nand U1153 (N_1153,N_1062,N_1068);
or U1154 (N_1154,N_1069,N_1059);
nand U1155 (N_1155,N_1038,N_1009);
nand U1156 (N_1156,N_1092,N_1052);
or U1157 (N_1157,N_1041,N_1049);
or U1158 (N_1158,N_1079,N_1064);
and U1159 (N_1159,N_1022,N_1013);
nor U1160 (N_1160,N_1070,N_1064);
and U1161 (N_1161,N_1077,N_1023);
xor U1162 (N_1162,N_1075,N_1041);
nor U1163 (N_1163,N_1083,N_1013);
nand U1164 (N_1164,N_1051,N_1046);
or U1165 (N_1165,N_1014,N_1073);
nand U1166 (N_1166,N_1049,N_1058);
xnor U1167 (N_1167,N_1095,N_1042);
xor U1168 (N_1168,N_1046,N_1054);
nor U1169 (N_1169,N_1004,N_1076);
or U1170 (N_1170,N_1011,N_1015);
xnor U1171 (N_1171,N_1009,N_1055);
and U1172 (N_1172,N_1087,N_1054);
xor U1173 (N_1173,N_1043,N_1091);
nor U1174 (N_1174,N_1091,N_1068);
xor U1175 (N_1175,N_1009,N_1049);
and U1176 (N_1176,N_1089,N_1046);
nand U1177 (N_1177,N_1048,N_1085);
nor U1178 (N_1178,N_1069,N_1072);
and U1179 (N_1179,N_1083,N_1038);
and U1180 (N_1180,N_1064,N_1021);
and U1181 (N_1181,N_1033,N_1057);
nand U1182 (N_1182,N_1054,N_1090);
nor U1183 (N_1183,N_1004,N_1002);
or U1184 (N_1184,N_1006,N_1017);
nand U1185 (N_1185,N_1013,N_1074);
and U1186 (N_1186,N_1084,N_1025);
nor U1187 (N_1187,N_1075,N_1074);
xor U1188 (N_1188,N_1045,N_1020);
xnor U1189 (N_1189,N_1021,N_1026);
nand U1190 (N_1190,N_1032,N_1014);
xor U1191 (N_1191,N_1029,N_1054);
or U1192 (N_1192,N_1068,N_1015);
and U1193 (N_1193,N_1065,N_1088);
or U1194 (N_1194,N_1099,N_1019);
or U1195 (N_1195,N_1003,N_1062);
and U1196 (N_1196,N_1062,N_1098);
and U1197 (N_1197,N_1065,N_1038);
and U1198 (N_1198,N_1077,N_1052);
xnor U1199 (N_1199,N_1060,N_1091);
xor U1200 (N_1200,N_1119,N_1100);
xnor U1201 (N_1201,N_1120,N_1174);
nor U1202 (N_1202,N_1175,N_1136);
or U1203 (N_1203,N_1146,N_1138);
nor U1204 (N_1204,N_1177,N_1110);
nand U1205 (N_1205,N_1158,N_1162);
nand U1206 (N_1206,N_1141,N_1147);
nor U1207 (N_1207,N_1169,N_1170);
and U1208 (N_1208,N_1160,N_1133);
or U1209 (N_1209,N_1184,N_1124);
nor U1210 (N_1210,N_1135,N_1176);
and U1211 (N_1211,N_1156,N_1191);
nand U1212 (N_1212,N_1151,N_1145);
nor U1213 (N_1213,N_1101,N_1104);
xor U1214 (N_1214,N_1164,N_1168);
or U1215 (N_1215,N_1103,N_1139);
nor U1216 (N_1216,N_1123,N_1140);
nor U1217 (N_1217,N_1107,N_1152);
nor U1218 (N_1218,N_1114,N_1149);
xnor U1219 (N_1219,N_1112,N_1129);
xor U1220 (N_1220,N_1148,N_1127);
nor U1221 (N_1221,N_1179,N_1125);
and U1222 (N_1222,N_1116,N_1187);
or U1223 (N_1223,N_1131,N_1159);
xor U1224 (N_1224,N_1157,N_1189);
xor U1225 (N_1225,N_1144,N_1113);
xor U1226 (N_1226,N_1134,N_1143);
xor U1227 (N_1227,N_1183,N_1106);
and U1228 (N_1228,N_1171,N_1172);
or U1229 (N_1229,N_1163,N_1128);
xnor U1230 (N_1230,N_1192,N_1193);
xnor U1231 (N_1231,N_1108,N_1130);
xnor U1232 (N_1232,N_1150,N_1195);
and U1233 (N_1233,N_1199,N_1167);
nand U1234 (N_1234,N_1197,N_1194);
nor U1235 (N_1235,N_1165,N_1186);
or U1236 (N_1236,N_1173,N_1126);
nor U1237 (N_1237,N_1105,N_1153);
or U1238 (N_1238,N_1122,N_1109);
and U1239 (N_1239,N_1154,N_1155);
xor U1240 (N_1240,N_1196,N_1188);
nand U1241 (N_1241,N_1182,N_1180);
xnor U1242 (N_1242,N_1185,N_1117);
xnor U1243 (N_1243,N_1132,N_1198);
or U1244 (N_1244,N_1178,N_1121);
and U1245 (N_1245,N_1181,N_1115);
xor U1246 (N_1246,N_1161,N_1102);
or U1247 (N_1247,N_1137,N_1118);
xor U1248 (N_1248,N_1166,N_1111);
and U1249 (N_1249,N_1142,N_1190);
xnor U1250 (N_1250,N_1184,N_1176);
xor U1251 (N_1251,N_1176,N_1168);
and U1252 (N_1252,N_1176,N_1116);
or U1253 (N_1253,N_1192,N_1156);
or U1254 (N_1254,N_1173,N_1111);
nand U1255 (N_1255,N_1140,N_1114);
nor U1256 (N_1256,N_1158,N_1133);
and U1257 (N_1257,N_1124,N_1132);
nand U1258 (N_1258,N_1173,N_1148);
xor U1259 (N_1259,N_1110,N_1179);
and U1260 (N_1260,N_1194,N_1166);
xor U1261 (N_1261,N_1125,N_1127);
nor U1262 (N_1262,N_1103,N_1115);
and U1263 (N_1263,N_1125,N_1158);
or U1264 (N_1264,N_1139,N_1115);
xor U1265 (N_1265,N_1107,N_1151);
nand U1266 (N_1266,N_1100,N_1146);
xor U1267 (N_1267,N_1136,N_1107);
xor U1268 (N_1268,N_1107,N_1163);
nor U1269 (N_1269,N_1186,N_1135);
xnor U1270 (N_1270,N_1133,N_1145);
nand U1271 (N_1271,N_1147,N_1117);
and U1272 (N_1272,N_1140,N_1158);
or U1273 (N_1273,N_1111,N_1152);
nand U1274 (N_1274,N_1170,N_1114);
nor U1275 (N_1275,N_1166,N_1193);
xor U1276 (N_1276,N_1146,N_1197);
and U1277 (N_1277,N_1158,N_1153);
xor U1278 (N_1278,N_1107,N_1157);
nor U1279 (N_1279,N_1165,N_1110);
or U1280 (N_1280,N_1103,N_1122);
nand U1281 (N_1281,N_1173,N_1199);
nor U1282 (N_1282,N_1151,N_1167);
or U1283 (N_1283,N_1146,N_1128);
or U1284 (N_1284,N_1180,N_1118);
nand U1285 (N_1285,N_1178,N_1135);
nor U1286 (N_1286,N_1153,N_1156);
xnor U1287 (N_1287,N_1164,N_1177);
xnor U1288 (N_1288,N_1170,N_1163);
or U1289 (N_1289,N_1147,N_1193);
and U1290 (N_1290,N_1113,N_1150);
nand U1291 (N_1291,N_1142,N_1137);
nor U1292 (N_1292,N_1117,N_1146);
or U1293 (N_1293,N_1167,N_1113);
nor U1294 (N_1294,N_1128,N_1107);
or U1295 (N_1295,N_1172,N_1135);
and U1296 (N_1296,N_1160,N_1197);
nor U1297 (N_1297,N_1184,N_1160);
nand U1298 (N_1298,N_1118,N_1145);
nand U1299 (N_1299,N_1166,N_1131);
xor U1300 (N_1300,N_1292,N_1224);
or U1301 (N_1301,N_1218,N_1272);
xnor U1302 (N_1302,N_1246,N_1273);
nand U1303 (N_1303,N_1275,N_1241);
and U1304 (N_1304,N_1238,N_1298);
xor U1305 (N_1305,N_1261,N_1269);
and U1306 (N_1306,N_1229,N_1287);
nor U1307 (N_1307,N_1281,N_1256);
nor U1308 (N_1308,N_1235,N_1236);
or U1309 (N_1309,N_1286,N_1203);
and U1310 (N_1310,N_1240,N_1289);
nand U1311 (N_1311,N_1265,N_1262);
nor U1312 (N_1312,N_1253,N_1290);
nor U1313 (N_1313,N_1234,N_1245);
or U1314 (N_1314,N_1202,N_1264);
nor U1315 (N_1315,N_1255,N_1200);
nor U1316 (N_1316,N_1209,N_1222);
nor U1317 (N_1317,N_1284,N_1214);
nand U1318 (N_1318,N_1276,N_1211);
and U1319 (N_1319,N_1233,N_1288);
or U1320 (N_1320,N_1257,N_1250);
nor U1321 (N_1321,N_1299,N_1213);
nor U1322 (N_1322,N_1219,N_1242);
xnor U1323 (N_1323,N_1205,N_1201);
nand U1324 (N_1324,N_1283,N_1267);
and U1325 (N_1325,N_1279,N_1268);
nand U1326 (N_1326,N_1207,N_1231);
nand U1327 (N_1327,N_1223,N_1252);
nand U1328 (N_1328,N_1293,N_1295);
or U1329 (N_1329,N_1285,N_1260);
nand U1330 (N_1330,N_1212,N_1258);
nor U1331 (N_1331,N_1291,N_1274);
xnor U1332 (N_1332,N_1225,N_1280);
xor U1333 (N_1333,N_1277,N_1206);
or U1334 (N_1334,N_1249,N_1228);
or U1335 (N_1335,N_1271,N_1208);
xor U1336 (N_1336,N_1232,N_1251);
nor U1337 (N_1337,N_1270,N_1230);
nand U1338 (N_1338,N_1220,N_1216);
and U1339 (N_1339,N_1294,N_1217);
or U1340 (N_1340,N_1215,N_1297);
or U1341 (N_1341,N_1259,N_1226);
nor U1342 (N_1342,N_1244,N_1204);
xnor U1343 (N_1343,N_1247,N_1263);
nor U1344 (N_1344,N_1296,N_1221);
and U1345 (N_1345,N_1239,N_1282);
xnor U1346 (N_1346,N_1227,N_1243);
or U1347 (N_1347,N_1266,N_1210);
xnor U1348 (N_1348,N_1248,N_1254);
or U1349 (N_1349,N_1278,N_1237);
and U1350 (N_1350,N_1291,N_1224);
and U1351 (N_1351,N_1215,N_1200);
nor U1352 (N_1352,N_1262,N_1299);
xor U1353 (N_1353,N_1292,N_1228);
nor U1354 (N_1354,N_1284,N_1222);
or U1355 (N_1355,N_1241,N_1272);
nor U1356 (N_1356,N_1249,N_1247);
xor U1357 (N_1357,N_1252,N_1251);
nand U1358 (N_1358,N_1233,N_1230);
nand U1359 (N_1359,N_1216,N_1204);
and U1360 (N_1360,N_1209,N_1285);
nor U1361 (N_1361,N_1299,N_1222);
nand U1362 (N_1362,N_1279,N_1257);
xnor U1363 (N_1363,N_1260,N_1292);
or U1364 (N_1364,N_1289,N_1282);
and U1365 (N_1365,N_1249,N_1238);
or U1366 (N_1366,N_1266,N_1274);
xnor U1367 (N_1367,N_1203,N_1207);
or U1368 (N_1368,N_1247,N_1230);
nor U1369 (N_1369,N_1230,N_1296);
xnor U1370 (N_1370,N_1230,N_1256);
or U1371 (N_1371,N_1255,N_1296);
or U1372 (N_1372,N_1256,N_1263);
nand U1373 (N_1373,N_1216,N_1241);
nor U1374 (N_1374,N_1263,N_1273);
nor U1375 (N_1375,N_1219,N_1287);
xor U1376 (N_1376,N_1258,N_1213);
and U1377 (N_1377,N_1243,N_1223);
or U1378 (N_1378,N_1238,N_1263);
and U1379 (N_1379,N_1242,N_1251);
nor U1380 (N_1380,N_1236,N_1263);
and U1381 (N_1381,N_1232,N_1240);
xor U1382 (N_1382,N_1244,N_1222);
nor U1383 (N_1383,N_1218,N_1231);
nor U1384 (N_1384,N_1212,N_1285);
nand U1385 (N_1385,N_1204,N_1262);
xor U1386 (N_1386,N_1270,N_1293);
xor U1387 (N_1387,N_1211,N_1246);
nand U1388 (N_1388,N_1225,N_1276);
nand U1389 (N_1389,N_1279,N_1265);
nand U1390 (N_1390,N_1227,N_1215);
xnor U1391 (N_1391,N_1226,N_1201);
nand U1392 (N_1392,N_1250,N_1266);
and U1393 (N_1393,N_1254,N_1260);
or U1394 (N_1394,N_1285,N_1204);
and U1395 (N_1395,N_1230,N_1215);
or U1396 (N_1396,N_1232,N_1260);
nand U1397 (N_1397,N_1282,N_1214);
nand U1398 (N_1398,N_1284,N_1297);
or U1399 (N_1399,N_1237,N_1246);
nor U1400 (N_1400,N_1337,N_1331);
xor U1401 (N_1401,N_1397,N_1332);
nor U1402 (N_1402,N_1318,N_1364);
nor U1403 (N_1403,N_1323,N_1328);
and U1404 (N_1404,N_1391,N_1381);
nand U1405 (N_1405,N_1359,N_1349);
and U1406 (N_1406,N_1375,N_1321);
xnor U1407 (N_1407,N_1304,N_1394);
or U1408 (N_1408,N_1392,N_1372);
xnor U1409 (N_1409,N_1358,N_1361);
nor U1410 (N_1410,N_1386,N_1312);
nand U1411 (N_1411,N_1336,N_1308);
and U1412 (N_1412,N_1384,N_1313);
xnor U1413 (N_1413,N_1302,N_1379);
and U1414 (N_1414,N_1368,N_1345);
or U1415 (N_1415,N_1377,N_1398);
nor U1416 (N_1416,N_1356,N_1388);
or U1417 (N_1417,N_1393,N_1351);
nand U1418 (N_1418,N_1396,N_1348);
nand U1419 (N_1419,N_1362,N_1366);
or U1420 (N_1420,N_1319,N_1346);
xnor U1421 (N_1421,N_1307,N_1353);
nand U1422 (N_1422,N_1340,N_1326);
nand U1423 (N_1423,N_1335,N_1324);
or U1424 (N_1424,N_1343,N_1378);
or U1425 (N_1425,N_1342,N_1320);
and U1426 (N_1426,N_1310,N_1373);
xor U1427 (N_1427,N_1333,N_1352);
nand U1428 (N_1428,N_1360,N_1370);
nand U1429 (N_1429,N_1382,N_1322);
nand U1430 (N_1430,N_1330,N_1306);
and U1431 (N_1431,N_1363,N_1327);
xnor U1432 (N_1432,N_1341,N_1399);
and U1433 (N_1433,N_1367,N_1315);
xor U1434 (N_1434,N_1311,N_1303);
and U1435 (N_1435,N_1354,N_1329);
nor U1436 (N_1436,N_1395,N_1357);
nand U1437 (N_1437,N_1389,N_1390);
and U1438 (N_1438,N_1338,N_1339);
nor U1439 (N_1439,N_1316,N_1380);
or U1440 (N_1440,N_1376,N_1371);
nor U1441 (N_1441,N_1383,N_1387);
and U1442 (N_1442,N_1347,N_1344);
nor U1443 (N_1443,N_1325,N_1355);
xnor U1444 (N_1444,N_1369,N_1305);
nor U1445 (N_1445,N_1309,N_1385);
and U1446 (N_1446,N_1365,N_1301);
nor U1447 (N_1447,N_1300,N_1374);
nand U1448 (N_1448,N_1350,N_1317);
or U1449 (N_1449,N_1334,N_1314);
or U1450 (N_1450,N_1386,N_1346);
nand U1451 (N_1451,N_1303,N_1381);
xor U1452 (N_1452,N_1384,N_1335);
nand U1453 (N_1453,N_1356,N_1308);
and U1454 (N_1454,N_1399,N_1381);
xnor U1455 (N_1455,N_1305,N_1330);
nand U1456 (N_1456,N_1379,N_1305);
or U1457 (N_1457,N_1330,N_1332);
xnor U1458 (N_1458,N_1365,N_1325);
or U1459 (N_1459,N_1323,N_1359);
nand U1460 (N_1460,N_1349,N_1330);
or U1461 (N_1461,N_1360,N_1351);
nand U1462 (N_1462,N_1356,N_1324);
nand U1463 (N_1463,N_1381,N_1395);
nand U1464 (N_1464,N_1311,N_1364);
and U1465 (N_1465,N_1383,N_1374);
nor U1466 (N_1466,N_1325,N_1310);
or U1467 (N_1467,N_1302,N_1349);
nand U1468 (N_1468,N_1315,N_1333);
and U1469 (N_1469,N_1350,N_1320);
or U1470 (N_1470,N_1390,N_1336);
and U1471 (N_1471,N_1326,N_1338);
and U1472 (N_1472,N_1360,N_1391);
and U1473 (N_1473,N_1335,N_1361);
nor U1474 (N_1474,N_1393,N_1335);
nor U1475 (N_1475,N_1319,N_1370);
nand U1476 (N_1476,N_1314,N_1335);
and U1477 (N_1477,N_1332,N_1393);
nor U1478 (N_1478,N_1369,N_1329);
nor U1479 (N_1479,N_1368,N_1306);
nand U1480 (N_1480,N_1305,N_1347);
nor U1481 (N_1481,N_1389,N_1312);
and U1482 (N_1482,N_1374,N_1318);
nor U1483 (N_1483,N_1349,N_1345);
and U1484 (N_1484,N_1356,N_1320);
nor U1485 (N_1485,N_1303,N_1360);
xnor U1486 (N_1486,N_1355,N_1391);
or U1487 (N_1487,N_1317,N_1385);
nand U1488 (N_1488,N_1317,N_1347);
or U1489 (N_1489,N_1307,N_1363);
nor U1490 (N_1490,N_1397,N_1361);
and U1491 (N_1491,N_1355,N_1351);
nand U1492 (N_1492,N_1388,N_1393);
and U1493 (N_1493,N_1354,N_1394);
nand U1494 (N_1494,N_1399,N_1397);
nor U1495 (N_1495,N_1350,N_1372);
nand U1496 (N_1496,N_1360,N_1397);
and U1497 (N_1497,N_1376,N_1352);
xor U1498 (N_1498,N_1306,N_1399);
or U1499 (N_1499,N_1373,N_1331);
nor U1500 (N_1500,N_1466,N_1459);
nand U1501 (N_1501,N_1418,N_1401);
xnor U1502 (N_1502,N_1429,N_1438);
xor U1503 (N_1503,N_1468,N_1476);
and U1504 (N_1504,N_1417,N_1457);
or U1505 (N_1505,N_1400,N_1493);
nor U1506 (N_1506,N_1474,N_1483);
or U1507 (N_1507,N_1480,N_1463);
nand U1508 (N_1508,N_1470,N_1433);
nand U1509 (N_1509,N_1471,N_1426);
xor U1510 (N_1510,N_1447,N_1492);
nand U1511 (N_1511,N_1414,N_1427);
or U1512 (N_1512,N_1448,N_1488);
nand U1513 (N_1513,N_1487,N_1443);
nor U1514 (N_1514,N_1444,N_1410);
and U1515 (N_1515,N_1415,N_1421);
nand U1516 (N_1516,N_1454,N_1412);
nor U1517 (N_1517,N_1440,N_1419);
and U1518 (N_1518,N_1481,N_1460);
or U1519 (N_1519,N_1450,N_1446);
xnor U1520 (N_1520,N_1409,N_1428);
and U1521 (N_1521,N_1431,N_1496);
nand U1522 (N_1522,N_1485,N_1462);
or U1523 (N_1523,N_1479,N_1456);
or U1524 (N_1524,N_1434,N_1445);
and U1525 (N_1525,N_1451,N_1472);
nand U1526 (N_1526,N_1477,N_1484);
nor U1527 (N_1527,N_1424,N_1402);
nand U1528 (N_1528,N_1413,N_1420);
xor U1529 (N_1529,N_1406,N_1422);
and U1530 (N_1530,N_1491,N_1408);
and U1531 (N_1531,N_1405,N_1494);
nor U1532 (N_1532,N_1497,N_1435);
nor U1533 (N_1533,N_1442,N_1478);
or U1534 (N_1534,N_1403,N_1439);
nand U1535 (N_1535,N_1489,N_1452);
nor U1536 (N_1536,N_1407,N_1455);
xnor U1537 (N_1537,N_1467,N_1458);
or U1538 (N_1538,N_1490,N_1436);
nor U1539 (N_1539,N_1441,N_1416);
and U1540 (N_1540,N_1453,N_1499);
or U1541 (N_1541,N_1475,N_1482);
xnor U1542 (N_1542,N_1430,N_1411);
nor U1543 (N_1543,N_1404,N_1473);
xnor U1544 (N_1544,N_1465,N_1461);
nor U1545 (N_1545,N_1498,N_1425);
nand U1546 (N_1546,N_1432,N_1495);
nor U1547 (N_1547,N_1464,N_1449);
nor U1548 (N_1548,N_1486,N_1469);
and U1549 (N_1549,N_1423,N_1437);
nor U1550 (N_1550,N_1464,N_1457);
and U1551 (N_1551,N_1483,N_1404);
xor U1552 (N_1552,N_1472,N_1443);
nand U1553 (N_1553,N_1412,N_1460);
and U1554 (N_1554,N_1493,N_1431);
xnor U1555 (N_1555,N_1419,N_1462);
xnor U1556 (N_1556,N_1471,N_1472);
or U1557 (N_1557,N_1471,N_1416);
nand U1558 (N_1558,N_1459,N_1448);
nand U1559 (N_1559,N_1418,N_1484);
xor U1560 (N_1560,N_1452,N_1478);
xnor U1561 (N_1561,N_1448,N_1469);
xor U1562 (N_1562,N_1430,N_1441);
and U1563 (N_1563,N_1456,N_1495);
nand U1564 (N_1564,N_1400,N_1444);
nor U1565 (N_1565,N_1495,N_1451);
and U1566 (N_1566,N_1499,N_1462);
nor U1567 (N_1567,N_1481,N_1499);
nand U1568 (N_1568,N_1492,N_1406);
or U1569 (N_1569,N_1499,N_1497);
or U1570 (N_1570,N_1404,N_1456);
nor U1571 (N_1571,N_1477,N_1447);
or U1572 (N_1572,N_1406,N_1459);
xnor U1573 (N_1573,N_1487,N_1431);
nor U1574 (N_1574,N_1462,N_1478);
nand U1575 (N_1575,N_1416,N_1456);
xor U1576 (N_1576,N_1405,N_1487);
nor U1577 (N_1577,N_1431,N_1418);
nand U1578 (N_1578,N_1471,N_1488);
nand U1579 (N_1579,N_1404,N_1409);
or U1580 (N_1580,N_1414,N_1458);
nand U1581 (N_1581,N_1456,N_1478);
or U1582 (N_1582,N_1424,N_1414);
xnor U1583 (N_1583,N_1419,N_1470);
xor U1584 (N_1584,N_1486,N_1499);
nor U1585 (N_1585,N_1443,N_1406);
nand U1586 (N_1586,N_1403,N_1493);
xnor U1587 (N_1587,N_1408,N_1474);
xor U1588 (N_1588,N_1491,N_1400);
nor U1589 (N_1589,N_1467,N_1486);
xnor U1590 (N_1590,N_1455,N_1468);
or U1591 (N_1591,N_1418,N_1406);
and U1592 (N_1592,N_1411,N_1477);
nor U1593 (N_1593,N_1435,N_1401);
xor U1594 (N_1594,N_1499,N_1478);
nand U1595 (N_1595,N_1441,N_1436);
and U1596 (N_1596,N_1445,N_1467);
or U1597 (N_1597,N_1471,N_1404);
xor U1598 (N_1598,N_1400,N_1482);
xnor U1599 (N_1599,N_1488,N_1453);
nor U1600 (N_1600,N_1566,N_1543);
and U1601 (N_1601,N_1521,N_1582);
or U1602 (N_1602,N_1514,N_1506);
nand U1603 (N_1603,N_1577,N_1551);
nand U1604 (N_1604,N_1547,N_1588);
or U1605 (N_1605,N_1584,N_1549);
nand U1606 (N_1606,N_1554,N_1541);
nor U1607 (N_1607,N_1574,N_1567);
nand U1608 (N_1608,N_1550,N_1500);
xnor U1609 (N_1609,N_1515,N_1508);
or U1610 (N_1610,N_1589,N_1568);
nand U1611 (N_1611,N_1520,N_1595);
xnor U1612 (N_1612,N_1538,N_1592);
and U1613 (N_1613,N_1539,N_1527);
and U1614 (N_1614,N_1572,N_1585);
nand U1615 (N_1615,N_1590,N_1507);
and U1616 (N_1616,N_1575,N_1502);
xor U1617 (N_1617,N_1571,N_1581);
nand U1618 (N_1618,N_1591,N_1501);
and U1619 (N_1619,N_1504,N_1557);
xnor U1620 (N_1620,N_1524,N_1594);
xnor U1621 (N_1621,N_1509,N_1556);
nor U1622 (N_1622,N_1573,N_1544);
nor U1623 (N_1623,N_1535,N_1516);
nand U1624 (N_1624,N_1540,N_1518);
xor U1625 (N_1625,N_1503,N_1526);
and U1626 (N_1626,N_1580,N_1596);
nand U1627 (N_1627,N_1576,N_1586);
or U1628 (N_1628,N_1548,N_1519);
and U1629 (N_1629,N_1545,N_1555);
and U1630 (N_1630,N_1579,N_1533);
xnor U1631 (N_1631,N_1562,N_1512);
nand U1632 (N_1632,N_1537,N_1510);
nand U1633 (N_1633,N_1513,N_1517);
and U1634 (N_1634,N_1597,N_1570);
xor U1635 (N_1635,N_1563,N_1569);
and U1636 (N_1636,N_1542,N_1525);
nand U1637 (N_1637,N_1553,N_1578);
xnor U1638 (N_1638,N_1558,N_1599);
or U1639 (N_1639,N_1565,N_1546);
nor U1640 (N_1640,N_1522,N_1587);
nor U1641 (N_1641,N_1561,N_1552);
xnor U1642 (N_1642,N_1530,N_1528);
nand U1643 (N_1643,N_1564,N_1534);
or U1644 (N_1644,N_1559,N_1536);
nand U1645 (N_1645,N_1560,N_1583);
xor U1646 (N_1646,N_1598,N_1511);
nand U1647 (N_1647,N_1531,N_1529);
and U1648 (N_1648,N_1505,N_1532);
nor U1649 (N_1649,N_1523,N_1593);
nor U1650 (N_1650,N_1556,N_1558);
xor U1651 (N_1651,N_1533,N_1545);
nand U1652 (N_1652,N_1507,N_1513);
nor U1653 (N_1653,N_1505,N_1507);
xnor U1654 (N_1654,N_1574,N_1504);
nor U1655 (N_1655,N_1538,N_1509);
xnor U1656 (N_1656,N_1559,N_1555);
and U1657 (N_1657,N_1576,N_1547);
and U1658 (N_1658,N_1570,N_1584);
nor U1659 (N_1659,N_1517,N_1593);
xor U1660 (N_1660,N_1503,N_1587);
or U1661 (N_1661,N_1554,N_1532);
nor U1662 (N_1662,N_1572,N_1567);
nor U1663 (N_1663,N_1505,N_1542);
nor U1664 (N_1664,N_1520,N_1597);
xnor U1665 (N_1665,N_1593,N_1502);
nor U1666 (N_1666,N_1543,N_1552);
nand U1667 (N_1667,N_1571,N_1556);
and U1668 (N_1668,N_1583,N_1524);
and U1669 (N_1669,N_1570,N_1544);
xnor U1670 (N_1670,N_1563,N_1571);
xnor U1671 (N_1671,N_1584,N_1508);
nand U1672 (N_1672,N_1525,N_1517);
or U1673 (N_1673,N_1575,N_1596);
xnor U1674 (N_1674,N_1520,N_1571);
xnor U1675 (N_1675,N_1514,N_1551);
or U1676 (N_1676,N_1521,N_1544);
nor U1677 (N_1677,N_1593,N_1586);
and U1678 (N_1678,N_1599,N_1506);
or U1679 (N_1679,N_1568,N_1565);
nand U1680 (N_1680,N_1521,N_1503);
xor U1681 (N_1681,N_1533,N_1527);
nand U1682 (N_1682,N_1564,N_1510);
nand U1683 (N_1683,N_1527,N_1576);
and U1684 (N_1684,N_1580,N_1517);
or U1685 (N_1685,N_1510,N_1509);
nor U1686 (N_1686,N_1514,N_1512);
xor U1687 (N_1687,N_1502,N_1594);
nand U1688 (N_1688,N_1599,N_1505);
xnor U1689 (N_1689,N_1578,N_1563);
nor U1690 (N_1690,N_1565,N_1572);
nand U1691 (N_1691,N_1525,N_1557);
or U1692 (N_1692,N_1593,N_1548);
xor U1693 (N_1693,N_1594,N_1529);
or U1694 (N_1694,N_1566,N_1538);
xnor U1695 (N_1695,N_1512,N_1575);
nor U1696 (N_1696,N_1507,N_1566);
xor U1697 (N_1697,N_1506,N_1592);
nor U1698 (N_1698,N_1589,N_1599);
or U1699 (N_1699,N_1582,N_1575);
nor U1700 (N_1700,N_1680,N_1654);
or U1701 (N_1701,N_1672,N_1613);
or U1702 (N_1702,N_1630,N_1645);
nor U1703 (N_1703,N_1643,N_1611);
and U1704 (N_1704,N_1658,N_1620);
nand U1705 (N_1705,N_1653,N_1605);
or U1706 (N_1706,N_1626,N_1675);
or U1707 (N_1707,N_1637,N_1689);
nor U1708 (N_1708,N_1679,N_1684);
xor U1709 (N_1709,N_1644,N_1667);
xnor U1710 (N_1710,N_1692,N_1625);
xor U1711 (N_1711,N_1603,N_1676);
or U1712 (N_1712,N_1685,N_1698);
xnor U1713 (N_1713,N_1641,N_1697);
and U1714 (N_1714,N_1622,N_1609);
nand U1715 (N_1715,N_1619,N_1628);
and U1716 (N_1716,N_1604,N_1694);
nand U1717 (N_1717,N_1607,N_1669);
nand U1718 (N_1718,N_1647,N_1633);
nand U1719 (N_1719,N_1612,N_1664);
or U1720 (N_1720,N_1677,N_1652);
xnor U1721 (N_1721,N_1606,N_1615);
nand U1722 (N_1722,N_1659,N_1656);
or U1723 (N_1723,N_1649,N_1693);
nor U1724 (N_1724,N_1690,N_1617);
xnor U1725 (N_1725,N_1678,N_1651);
nand U1726 (N_1726,N_1682,N_1660);
nor U1727 (N_1727,N_1668,N_1663);
nor U1728 (N_1728,N_1686,N_1688);
and U1729 (N_1729,N_1635,N_1618);
xor U1730 (N_1730,N_1638,N_1632);
and U1731 (N_1731,N_1691,N_1699);
or U1732 (N_1732,N_1616,N_1634);
nor U1733 (N_1733,N_1665,N_1601);
nand U1734 (N_1734,N_1623,N_1642);
or U1735 (N_1735,N_1610,N_1614);
xnor U1736 (N_1736,N_1671,N_1648);
nor U1737 (N_1737,N_1602,N_1639);
xnor U1738 (N_1738,N_1673,N_1636);
and U1739 (N_1739,N_1624,N_1683);
and U1740 (N_1740,N_1687,N_1608);
nand U1741 (N_1741,N_1629,N_1650);
and U1742 (N_1742,N_1600,N_1661);
nand U1743 (N_1743,N_1655,N_1640);
or U1744 (N_1744,N_1662,N_1681);
and U1745 (N_1745,N_1631,N_1627);
nor U1746 (N_1746,N_1674,N_1646);
or U1747 (N_1747,N_1670,N_1696);
and U1748 (N_1748,N_1621,N_1666);
and U1749 (N_1749,N_1657,N_1695);
nand U1750 (N_1750,N_1688,N_1648);
nand U1751 (N_1751,N_1609,N_1601);
or U1752 (N_1752,N_1609,N_1611);
nand U1753 (N_1753,N_1635,N_1619);
nand U1754 (N_1754,N_1666,N_1664);
and U1755 (N_1755,N_1607,N_1629);
and U1756 (N_1756,N_1692,N_1666);
and U1757 (N_1757,N_1679,N_1637);
xnor U1758 (N_1758,N_1627,N_1628);
nor U1759 (N_1759,N_1615,N_1627);
nand U1760 (N_1760,N_1614,N_1659);
or U1761 (N_1761,N_1677,N_1601);
xnor U1762 (N_1762,N_1683,N_1684);
and U1763 (N_1763,N_1663,N_1619);
or U1764 (N_1764,N_1676,N_1696);
nor U1765 (N_1765,N_1684,N_1640);
xor U1766 (N_1766,N_1669,N_1660);
or U1767 (N_1767,N_1626,N_1665);
and U1768 (N_1768,N_1605,N_1651);
and U1769 (N_1769,N_1605,N_1609);
xnor U1770 (N_1770,N_1697,N_1667);
xnor U1771 (N_1771,N_1661,N_1692);
nand U1772 (N_1772,N_1690,N_1636);
nand U1773 (N_1773,N_1674,N_1657);
nor U1774 (N_1774,N_1614,N_1693);
xnor U1775 (N_1775,N_1696,N_1603);
nand U1776 (N_1776,N_1622,N_1663);
and U1777 (N_1777,N_1626,N_1602);
xor U1778 (N_1778,N_1661,N_1606);
or U1779 (N_1779,N_1640,N_1657);
xnor U1780 (N_1780,N_1639,N_1628);
nand U1781 (N_1781,N_1664,N_1682);
or U1782 (N_1782,N_1641,N_1613);
or U1783 (N_1783,N_1635,N_1685);
nand U1784 (N_1784,N_1662,N_1626);
nand U1785 (N_1785,N_1669,N_1623);
xor U1786 (N_1786,N_1648,N_1600);
and U1787 (N_1787,N_1689,N_1664);
xnor U1788 (N_1788,N_1631,N_1658);
nand U1789 (N_1789,N_1646,N_1636);
xor U1790 (N_1790,N_1633,N_1644);
and U1791 (N_1791,N_1690,N_1606);
nand U1792 (N_1792,N_1678,N_1689);
and U1793 (N_1793,N_1608,N_1632);
nand U1794 (N_1794,N_1638,N_1656);
or U1795 (N_1795,N_1644,N_1600);
xor U1796 (N_1796,N_1676,N_1626);
nand U1797 (N_1797,N_1672,N_1639);
xnor U1798 (N_1798,N_1604,N_1662);
or U1799 (N_1799,N_1649,N_1692);
xnor U1800 (N_1800,N_1716,N_1747);
xnor U1801 (N_1801,N_1714,N_1727);
xor U1802 (N_1802,N_1769,N_1742);
nor U1803 (N_1803,N_1775,N_1713);
nor U1804 (N_1804,N_1728,N_1796);
nand U1805 (N_1805,N_1785,N_1740);
nor U1806 (N_1806,N_1758,N_1704);
nor U1807 (N_1807,N_1770,N_1710);
nand U1808 (N_1808,N_1746,N_1783);
xor U1809 (N_1809,N_1767,N_1763);
nor U1810 (N_1810,N_1781,N_1735);
xnor U1811 (N_1811,N_1755,N_1779);
nor U1812 (N_1812,N_1792,N_1777);
nor U1813 (N_1813,N_1753,N_1745);
xnor U1814 (N_1814,N_1737,N_1705);
and U1815 (N_1815,N_1778,N_1720);
xor U1816 (N_1816,N_1751,N_1797);
and U1817 (N_1817,N_1773,N_1738);
nand U1818 (N_1818,N_1765,N_1717);
and U1819 (N_1819,N_1799,N_1776);
or U1820 (N_1820,N_1774,N_1701);
xnor U1821 (N_1821,N_1757,N_1721);
and U1822 (N_1822,N_1739,N_1726);
or U1823 (N_1823,N_1760,N_1748);
nand U1824 (N_1824,N_1752,N_1787);
and U1825 (N_1825,N_1708,N_1772);
nand U1826 (N_1826,N_1741,N_1707);
nor U1827 (N_1827,N_1718,N_1729);
nor U1828 (N_1828,N_1768,N_1761);
nor U1829 (N_1829,N_1703,N_1711);
xnor U1830 (N_1830,N_1788,N_1731);
and U1831 (N_1831,N_1749,N_1790);
and U1832 (N_1832,N_1789,N_1730);
and U1833 (N_1833,N_1733,N_1702);
and U1834 (N_1834,N_1744,N_1732);
nor U1835 (N_1835,N_1719,N_1723);
nand U1836 (N_1836,N_1736,N_1771);
or U1837 (N_1837,N_1793,N_1795);
or U1838 (N_1838,N_1715,N_1743);
nand U1839 (N_1839,N_1700,N_1725);
and U1840 (N_1840,N_1734,N_1759);
and U1841 (N_1841,N_1786,N_1706);
and U1842 (N_1842,N_1762,N_1784);
nor U1843 (N_1843,N_1754,N_1750);
or U1844 (N_1844,N_1709,N_1794);
xor U1845 (N_1845,N_1712,N_1798);
nor U1846 (N_1846,N_1782,N_1780);
and U1847 (N_1847,N_1724,N_1756);
xor U1848 (N_1848,N_1764,N_1791);
nand U1849 (N_1849,N_1722,N_1766);
nor U1850 (N_1850,N_1759,N_1714);
or U1851 (N_1851,N_1732,N_1703);
and U1852 (N_1852,N_1711,N_1718);
xor U1853 (N_1853,N_1768,N_1758);
xor U1854 (N_1854,N_1777,N_1726);
and U1855 (N_1855,N_1784,N_1738);
nand U1856 (N_1856,N_1737,N_1722);
and U1857 (N_1857,N_1778,N_1799);
nor U1858 (N_1858,N_1749,N_1753);
xor U1859 (N_1859,N_1700,N_1754);
or U1860 (N_1860,N_1748,N_1765);
or U1861 (N_1861,N_1744,N_1719);
nor U1862 (N_1862,N_1798,N_1784);
nand U1863 (N_1863,N_1730,N_1778);
and U1864 (N_1864,N_1722,N_1758);
or U1865 (N_1865,N_1740,N_1784);
and U1866 (N_1866,N_1732,N_1773);
and U1867 (N_1867,N_1746,N_1762);
xor U1868 (N_1868,N_1702,N_1758);
nor U1869 (N_1869,N_1762,N_1788);
xnor U1870 (N_1870,N_1710,N_1797);
nand U1871 (N_1871,N_1761,N_1780);
nand U1872 (N_1872,N_1717,N_1772);
nor U1873 (N_1873,N_1708,N_1700);
nor U1874 (N_1874,N_1797,N_1746);
and U1875 (N_1875,N_1733,N_1701);
nand U1876 (N_1876,N_1783,N_1768);
xnor U1877 (N_1877,N_1769,N_1783);
xor U1878 (N_1878,N_1709,N_1742);
nand U1879 (N_1879,N_1737,N_1758);
nand U1880 (N_1880,N_1798,N_1751);
and U1881 (N_1881,N_1736,N_1775);
nand U1882 (N_1882,N_1766,N_1782);
nor U1883 (N_1883,N_1736,N_1743);
xor U1884 (N_1884,N_1712,N_1742);
and U1885 (N_1885,N_1716,N_1728);
and U1886 (N_1886,N_1771,N_1765);
and U1887 (N_1887,N_1723,N_1754);
xor U1888 (N_1888,N_1759,N_1797);
nand U1889 (N_1889,N_1769,N_1718);
or U1890 (N_1890,N_1719,N_1753);
and U1891 (N_1891,N_1771,N_1734);
or U1892 (N_1892,N_1715,N_1723);
nor U1893 (N_1893,N_1728,N_1719);
nand U1894 (N_1894,N_1758,N_1785);
or U1895 (N_1895,N_1763,N_1728);
nand U1896 (N_1896,N_1769,N_1700);
nor U1897 (N_1897,N_1768,N_1727);
xnor U1898 (N_1898,N_1717,N_1737);
and U1899 (N_1899,N_1759,N_1785);
xnor U1900 (N_1900,N_1811,N_1849);
and U1901 (N_1901,N_1805,N_1877);
xor U1902 (N_1902,N_1874,N_1886);
nand U1903 (N_1903,N_1885,N_1856);
nand U1904 (N_1904,N_1875,N_1847);
nand U1905 (N_1905,N_1881,N_1825);
nor U1906 (N_1906,N_1841,N_1837);
nand U1907 (N_1907,N_1860,N_1895);
nor U1908 (N_1908,N_1870,N_1899);
or U1909 (N_1909,N_1884,N_1894);
xnor U1910 (N_1910,N_1867,N_1810);
xor U1911 (N_1911,N_1812,N_1862);
and U1912 (N_1912,N_1802,N_1815);
or U1913 (N_1913,N_1829,N_1889);
xor U1914 (N_1914,N_1830,N_1844);
or U1915 (N_1915,N_1868,N_1819);
or U1916 (N_1916,N_1861,N_1817);
nor U1917 (N_1917,N_1808,N_1846);
nor U1918 (N_1918,N_1851,N_1831);
nand U1919 (N_1919,N_1807,N_1833);
xnor U1920 (N_1920,N_1854,N_1800);
or U1921 (N_1921,N_1863,N_1865);
or U1922 (N_1922,N_1835,N_1891);
nor U1923 (N_1923,N_1855,N_1823);
and U1924 (N_1924,N_1878,N_1820);
nor U1925 (N_1925,N_1834,N_1821);
xor U1926 (N_1926,N_1896,N_1848);
and U1927 (N_1927,N_1818,N_1857);
xor U1928 (N_1928,N_1828,N_1879);
nor U1929 (N_1929,N_1826,N_1883);
and U1930 (N_1930,N_1801,N_1845);
or U1931 (N_1931,N_1809,N_1814);
or U1932 (N_1932,N_1840,N_1866);
and U1933 (N_1933,N_1838,N_1893);
or U1934 (N_1934,N_1880,N_1804);
or U1935 (N_1935,N_1842,N_1897);
nor U1936 (N_1936,N_1892,N_1887);
or U1937 (N_1937,N_1803,N_1832);
xnor U1938 (N_1938,N_1836,N_1852);
and U1939 (N_1939,N_1871,N_1824);
nand U1940 (N_1940,N_1850,N_1859);
nand U1941 (N_1941,N_1822,N_1858);
and U1942 (N_1942,N_1898,N_1888);
and U1943 (N_1943,N_1816,N_1843);
and U1944 (N_1944,N_1876,N_1890);
and U1945 (N_1945,N_1813,N_1806);
xnor U1946 (N_1946,N_1839,N_1864);
nand U1947 (N_1947,N_1873,N_1869);
and U1948 (N_1948,N_1882,N_1872);
and U1949 (N_1949,N_1853,N_1827);
or U1950 (N_1950,N_1814,N_1808);
and U1951 (N_1951,N_1802,N_1870);
nor U1952 (N_1952,N_1866,N_1873);
or U1953 (N_1953,N_1850,N_1838);
nand U1954 (N_1954,N_1803,N_1837);
nand U1955 (N_1955,N_1890,N_1886);
and U1956 (N_1956,N_1866,N_1844);
and U1957 (N_1957,N_1830,N_1820);
and U1958 (N_1958,N_1846,N_1825);
and U1959 (N_1959,N_1872,N_1831);
and U1960 (N_1960,N_1820,N_1800);
xnor U1961 (N_1961,N_1868,N_1887);
and U1962 (N_1962,N_1854,N_1825);
and U1963 (N_1963,N_1812,N_1823);
nor U1964 (N_1964,N_1858,N_1803);
xnor U1965 (N_1965,N_1841,N_1897);
or U1966 (N_1966,N_1863,N_1818);
xor U1967 (N_1967,N_1800,N_1899);
nor U1968 (N_1968,N_1825,N_1820);
or U1969 (N_1969,N_1837,N_1849);
or U1970 (N_1970,N_1852,N_1822);
nor U1971 (N_1971,N_1873,N_1839);
and U1972 (N_1972,N_1842,N_1828);
and U1973 (N_1973,N_1811,N_1893);
nor U1974 (N_1974,N_1822,N_1896);
xnor U1975 (N_1975,N_1875,N_1879);
and U1976 (N_1976,N_1829,N_1830);
xor U1977 (N_1977,N_1891,N_1865);
or U1978 (N_1978,N_1894,N_1837);
nor U1979 (N_1979,N_1881,N_1868);
nand U1980 (N_1980,N_1814,N_1851);
or U1981 (N_1981,N_1838,N_1806);
xor U1982 (N_1982,N_1878,N_1890);
nand U1983 (N_1983,N_1846,N_1856);
nand U1984 (N_1984,N_1849,N_1878);
and U1985 (N_1985,N_1815,N_1811);
or U1986 (N_1986,N_1885,N_1837);
nor U1987 (N_1987,N_1806,N_1829);
nor U1988 (N_1988,N_1803,N_1893);
and U1989 (N_1989,N_1887,N_1891);
or U1990 (N_1990,N_1895,N_1827);
or U1991 (N_1991,N_1898,N_1823);
and U1992 (N_1992,N_1876,N_1819);
and U1993 (N_1993,N_1818,N_1866);
or U1994 (N_1994,N_1858,N_1897);
xnor U1995 (N_1995,N_1816,N_1821);
or U1996 (N_1996,N_1871,N_1855);
and U1997 (N_1997,N_1867,N_1827);
nor U1998 (N_1998,N_1800,N_1862);
or U1999 (N_1999,N_1893,N_1852);
and U2000 (N_2000,N_1998,N_1948);
or U2001 (N_2001,N_1918,N_1988);
nor U2002 (N_2002,N_1965,N_1956);
and U2003 (N_2003,N_1963,N_1986);
nor U2004 (N_2004,N_1919,N_1913);
nor U2005 (N_2005,N_1983,N_1962);
and U2006 (N_2006,N_1984,N_1908);
nand U2007 (N_2007,N_1941,N_1991);
or U2008 (N_2008,N_1905,N_1935);
and U2009 (N_2009,N_1926,N_1915);
and U2010 (N_2010,N_1902,N_1987);
nand U2011 (N_2011,N_1976,N_1955);
or U2012 (N_2012,N_1909,N_1932);
and U2013 (N_2013,N_1917,N_1901);
xor U2014 (N_2014,N_1922,N_1927);
nand U2015 (N_2015,N_1989,N_1959);
xnor U2016 (N_2016,N_1904,N_1907);
or U2017 (N_2017,N_1993,N_1929);
and U2018 (N_2018,N_1930,N_1958);
or U2019 (N_2019,N_1971,N_1949);
nand U2020 (N_2020,N_1960,N_1972);
xnor U2021 (N_2021,N_1966,N_1954);
nor U2022 (N_2022,N_1931,N_1934);
nand U2023 (N_2023,N_1937,N_1923);
and U2024 (N_2024,N_1974,N_1985);
or U2025 (N_2025,N_1910,N_1967);
or U2026 (N_2026,N_1903,N_1933);
nor U2027 (N_2027,N_1978,N_1975);
nand U2028 (N_2028,N_1951,N_1921);
nor U2029 (N_2029,N_1906,N_1914);
or U2030 (N_2030,N_1995,N_1977);
or U2031 (N_2031,N_1964,N_1911);
or U2032 (N_2032,N_1996,N_1969);
nand U2033 (N_2033,N_1912,N_1982);
nor U2034 (N_2034,N_1945,N_1953);
or U2035 (N_2035,N_1939,N_1968);
nand U2036 (N_2036,N_1920,N_1961);
or U2037 (N_2037,N_1900,N_1947);
nor U2038 (N_2038,N_1999,N_1938);
xor U2039 (N_2039,N_1940,N_1943);
nor U2040 (N_2040,N_1980,N_1925);
and U2041 (N_2041,N_1928,N_1950);
nor U2042 (N_2042,N_1979,N_1997);
nand U2043 (N_2043,N_1973,N_1994);
and U2044 (N_2044,N_1936,N_1924);
and U2045 (N_2045,N_1992,N_1946);
nand U2046 (N_2046,N_1981,N_1952);
xor U2047 (N_2047,N_1957,N_1990);
xnor U2048 (N_2048,N_1942,N_1916);
nor U2049 (N_2049,N_1944,N_1970);
nand U2050 (N_2050,N_1931,N_1946);
or U2051 (N_2051,N_1985,N_1958);
xor U2052 (N_2052,N_1951,N_1978);
nand U2053 (N_2053,N_1903,N_1965);
xnor U2054 (N_2054,N_1941,N_1932);
xor U2055 (N_2055,N_1904,N_1980);
xnor U2056 (N_2056,N_1922,N_1940);
and U2057 (N_2057,N_1922,N_1925);
xor U2058 (N_2058,N_1983,N_1925);
nor U2059 (N_2059,N_1917,N_1938);
nand U2060 (N_2060,N_1951,N_1977);
nor U2061 (N_2061,N_1978,N_1962);
nor U2062 (N_2062,N_1962,N_1923);
nor U2063 (N_2063,N_1901,N_1964);
or U2064 (N_2064,N_1906,N_1957);
nand U2065 (N_2065,N_1902,N_1979);
and U2066 (N_2066,N_1992,N_1929);
nand U2067 (N_2067,N_1982,N_1981);
or U2068 (N_2068,N_1943,N_1916);
xor U2069 (N_2069,N_1927,N_1977);
nand U2070 (N_2070,N_1924,N_1948);
and U2071 (N_2071,N_1966,N_1990);
or U2072 (N_2072,N_1982,N_1920);
xor U2073 (N_2073,N_1991,N_1911);
and U2074 (N_2074,N_1922,N_1966);
and U2075 (N_2075,N_1908,N_1955);
nor U2076 (N_2076,N_1965,N_1915);
xor U2077 (N_2077,N_1941,N_1907);
nor U2078 (N_2078,N_1929,N_1954);
xor U2079 (N_2079,N_1933,N_1931);
nand U2080 (N_2080,N_1977,N_1916);
xnor U2081 (N_2081,N_1969,N_1919);
or U2082 (N_2082,N_1949,N_1998);
or U2083 (N_2083,N_1907,N_1902);
nand U2084 (N_2084,N_1966,N_1970);
nand U2085 (N_2085,N_1917,N_1984);
xnor U2086 (N_2086,N_1960,N_1906);
nand U2087 (N_2087,N_1963,N_1931);
nand U2088 (N_2088,N_1942,N_1912);
or U2089 (N_2089,N_1973,N_1985);
and U2090 (N_2090,N_1901,N_1990);
or U2091 (N_2091,N_1915,N_1921);
nor U2092 (N_2092,N_1958,N_1989);
or U2093 (N_2093,N_1979,N_1968);
nand U2094 (N_2094,N_1961,N_1973);
xor U2095 (N_2095,N_1935,N_1919);
and U2096 (N_2096,N_1903,N_1971);
nor U2097 (N_2097,N_1963,N_1949);
xor U2098 (N_2098,N_1956,N_1959);
and U2099 (N_2099,N_1926,N_1962);
or U2100 (N_2100,N_2052,N_2064);
nor U2101 (N_2101,N_2025,N_2012);
and U2102 (N_2102,N_2071,N_2048);
and U2103 (N_2103,N_2077,N_2010);
nor U2104 (N_2104,N_2021,N_2070);
nand U2105 (N_2105,N_2060,N_2041);
nor U2106 (N_2106,N_2024,N_2005);
or U2107 (N_2107,N_2098,N_2069);
and U2108 (N_2108,N_2013,N_2009);
nand U2109 (N_2109,N_2072,N_2056);
or U2110 (N_2110,N_2006,N_2081);
and U2111 (N_2111,N_2037,N_2089);
xor U2112 (N_2112,N_2020,N_2090);
nor U2113 (N_2113,N_2082,N_2046);
or U2114 (N_2114,N_2044,N_2093);
nand U2115 (N_2115,N_2022,N_2000);
and U2116 (N_2116,N_2080,N_2017);
or U2117 (N_2117,N_2066,N_2067);
nor U2118 (N_2118,N_2073,N_2008);
nor U2119 (N_2119,N_2062,N_2087);
or U2120 (N_2120,N_2027,N_2032);
xnor U2121 (N_2121,N_2031,N_2034);
nor U2122 (N_2122,N_2038,N_2086);
nand U2123 (N_2123,N_2035,N_2026);
and U2124 (N_2124,N_2014,N_2097);
xnor U2125 (N_2125,N_2047,N_2059);
nand U2126 (N_2126,N_2078,N_2099);
nor U2127 (N_2127,N_2039,N_2053);
nand U2128 (N_2128,N_2088,N_2084);
or U2129 (N_2129,N_2045,N_2076);
and U2130 (N_2130,N_2043,N_2095);
and U2131 (N_2131,N_2040,N_2015);
or U2132 (N_2132,N_2050,N_2019);
nand U2133 (N_2133,N_2018,N_2091);
nand U2134 (N_2134,N_2001,N_2063);
xor U2135 (N_2135,N_2030,N_2051);
nand U2136 (N_2136,N_2002,N_2068);
or U2137 (N_2137,N_2094,N_2054);
and U2138 (N_2138,N_2074,N_2028);
and U2139 (N_2139,N_2061,N_2079);
nor U2140 (N_2140,N_2058,N_2023);
nor U2141 (N_2141,N_2075,N_2085);
or U2142 (N_2142,N_2055,N_2029);
nor U2143 (N_2143,N_2011,N_2057);
or U2144 (N_2144,N_2096,N_2036);
and U2145 (N_2145,N_2042,N_2016);
or U2146 (N_2146,N_2003,N_2083);
xnor U2147 (N_2147,N_2033,N_2049);
and U2148 (N_2148,N_2065,N_2007);
nor U2149 (N_2149,N_2004,N_2092);
or U2150 (N_2150,N_2098,N_2001);
nand U2151 (N_2151,N_2018,N_2052);
xnor U2152 (N_2152,N_2071,N_2023);
nor U2153 (N_2153,N_2022,N_2016);
nand U2154 (N_2154,N_2071,N_2091);
and U2155 (N_2155,N_2017,N_2075);
or U2156 (N_2156,N_2047,N_2078);
or U2157 (N_2157,N_2008,N_2090);
or U2158 (N_2158,N_2094,N_2034);
nor U2159 (N_2159,N_2056,N_2050);
nand U2160 (N_2160,N_2007,N_2078);
nand U2161 (N_2161,N_2015,N_2095);
xor U2162 (N_2162,N_2001,N_2039);
nand U2163 (N_2163,N_2022,N_2086);
xor U2164 (N_2164,N_2050,N_2093);
and U2165 (N_2165,N_2045,N_2052);
nand U2166 (N_2166,N_2021,N_2044);
nor U2167 (N_2167,N_2007,N_2068);
nor U2168 (N_2168,N_2044,N_2018);
or U2169 (N_2169,N_2025,N_2000);
and U2170 (N_2170,N_2064,N_2003);
or U2171 (N_2171,N_2003,N_2070);
or U2172 (N_2172,N_2086,N_2005);
xnor U2173 (N_2173,N_2041,N_2075);
or U2174 (N_2174,N_2074,N_2049);
and U2175 (N_2175,N_2060,N_2095);
xor U2176 (N_2176,N_2099,N_2041);
and U2177 (N_2177,N_2064,N_2088);
or U2178 (N_2178,N_2081,N_2059);
nand U2179 (N_2179,N_2093,N_2091);
nand U2180 (N_2180,N_2070,N_2094);
xor U2181 (N_2181,N_2088,N_2086);
xnor U2182 (N_2182,N_2046,N_2063);
or U2183 (N_2183,N_2071,N_2041);
nor U2184 (N_2184,N_2086,N_2000);
or U2185 (N_2185,N_2009,N_2031);
nor U2186 (N_2186,N_2028,N_2039);
and U2187 (N_2187,N_2006,N_2030);
or U2188 (N_2188,N_2078,N_2002);
nor U2189 (N_2189,N_2088,N_2005);
or U2190 (N_2190,N_2025,N_2067);
or U2191 (N_2191,N_2048,N_2083);
or U2192 (N_2192,N_2037,N_2018);
or U2193 (N_2193,N_2031,N_2076);
xnor U2194 (N_2194,N_2072,N_2013);
and U2195 (N_2195,N_2005,N_2052);
nand U2196 (N_2196,N_2021,N_2009);
and U2197 (N_2197,N_2074,N_2050);
nor U2198 (N_2198,N_2020,N_2004);
or U2199 (N_2199,N_2058,N_2077);
or U2200 (N_2200,N_2110,N_2178);
and U2201 (N_2201,N_2136,N_2166);
nand U2202 (N_2202,N_2113,N_2126);
xor U2203 (N_2203,N_2112,N_2135);
and U2204 (N_2204,N_2124,N_2109);
nand U2205 (N_2205,N_2105,N_2107);
nand U2206 (N_2206,N_2171,N_2102);
xor U2207 (N_2207,N_2174,N_2150);
and U2208 (N_2208,N_2153,N_2188);
nor U2209 (N_2209,N_2182,N_2156);
nor U2210 (N_2210,N_2148,N_2139);
and U2211 (N_2211,N_2123,N_2196);
and U2212 (N_2212,N_2147,N_2121);
nor U2213 (N_2213,N_2194,N_2193);
nand U2214 (N_2214,N_2151,N_2131);
xor U2215 (N_2215,N_2164,N_2160);
and U2216 (N_2216,N_2108,N_2140);
xor U2217 (N_2217,N_2168,N_2119);
or U2218 (N_2218,N_2169,N_2125);
nor U2219 (N_2219,N_2159,N_2143);
xnor U2220 (N_2220,N_2176,N_2155);
xnor U2221 (N_2221,N_2116,N_2197);
and U2222 (N_2222,N_2185,N_2120);
nor U2223 (N_2223,N_2138,N_2158);
nor U2224 (N_2224,N_2130,N_2111);
or U2225 (N_2225,N_2122,N_2161);
and U2226 (N_2226,N_2129,N_2104);
and U2227 (N_2227,N_2144,N_2180);
and U2228 (N_2228,N_2134,N_2141);
nand U2229 (N_2229,N_2157,N_2179);
or U2230 (N_2230,N_2106,N_2142);
or U2231 (N_2231,N_2177,N_2167);
or U2232 (N_2232,N_2137,N_2175);
and U2233 (N_2233,N_2115,N_2118);
or U2234 (N_2234,N_2170,N_2128);
xnor U2235 (N_2235,N_2152,N_2100);
nand U2236 (N_2236,N_2186,N_2132);
and U2237 (N_2237,N_2198,N_2199);
nor U2238 (N_2238,N_2189,N_2190);
nor U2239 (N_2239,N_2162,N_2187);
nor U2240 (N_2240,N_2154,N_2149);
and U2241 (N_2241,N_2127,N_2114);
nand U2242 (N_2242,N_2145,N_2172);
nand U2243 (N_2243,N_2103,N_2183);
and U2244 (N_2244,N_2117,N_2184);
or U2245 (N_2245,N_2101,N_2133);
and U2246 (N_2246,N_2195,N_2163);
and U2247 (N_2247,N_2173,N_2181);
nor U2248 (N_2248,N_2192,N_2165);
and U2249 (N_2249,N_2146,N_2191);
xor U2250 (N_2250,N_2161,N_2181);
nor U2251 (N_2251,N_2142,N_2143);
and U2252 (N_2252,N_2149,N_2122);
xnor U2253 (N_2253,N_2189,N_2117);
xnor U2254 (N_2254,N_2129,N_2179);
and U2255 (N_2255,N_2169,N_2167);
nor U2256 (N_2256,N_2131,N_2167);
xnor U2257 (N_2257,N_2131,N_2120);
xnor U2258 (N_2258,N_2154,N_2125);
or U2259 (N_2259,N_2158,N_2170);
nand U2260 (N_2260,N_2147,N_2130);
xor U2261 (N_2261,N_2184,N_2194);
or U2262 (N_2262,N_2123,N_2177);
xor U2263 (N_2263,N_2120,N_2153);
xnor U2264 (N_2264,N_2177,N_2155);
or U2265 (N_2265,N_2166,N_2127);
xnor U2266 (N_2266,N_2183,N_2186);
nand U2267 (N_2267,N_2149,N_2119);
nand U2268 (N_2268,N_2192,N_2129);
or U2269 (N_2269,N_2171,N_2111);
nor U2270 (N_2270,N_2110,N_2194);
and U2271 (N_2271,N_2198,N_2161);
nor U2272 (N_2272,N_2166,N_2102);
and U2273 (N_2273,N_2165,N_2162);
xor U2274 (N_2274,N_2145,N_2121);
nand U2275 (N_2275,N_2184,N_2192);
and U2276 (N_2276,N_2128,N_2109);
nor U2277 (N_2277,N_2101,N_2188);
xnor U2278 (N_2278,N_2113,N_2152);
nand U2279 (N_2279,N_2141,N_2199);
or U2280 (N_2280,N_2106,N_2152);
nor U2281 (N_2281,N_2108,N_2189);
nor U2282 (N_2282,N_2141,N_2110);
and U2283 (N_2283,N_2107,N_2181);
or U2284 (N_2284,N_2130,N_2119);
nand U2285 (N_2285,N_2184,N_2128);
or U2286 (N_2286,N_2126,N_2180);
nor U2287 (N_2287,N_2179,N_2112);
nor U2288 (N_2288,N_2140,N_2155);
nand U2289 (N_2289,N_2118,N_2133);
and U2290 (N_2290,N_2121,N_2148);
nand U2291 (N_2291,N_2108,N_2181);
nor U2292 (N_2292,N_2149,N_2105);
xnor U2293 (N_2293,N_2111,N_2172);
or U2294 (N_2294,N_2104,N_2185);
nor U2295 (N_2295,N_2140,N_2139);
nor U2296 (N_2296,N_2144,N_2123);
and U2297 (N_2297,N_2155,N_2165);
xnor U2298 (N_2298,N_2197,N_2145);
and U2299 (N_2299,N_2107,N_2184);
or U2300 (N_2300,N_2278,N_2289);
xnor U2301 (N_2301,N_2207,N_2273);
or U2302 (N_2302,N_2269,N_2218);
nor U2303 (N_2303,N_2214,N_2291);
and U2304 (N_2304,N_2243,N_2279);
xnor U2305 (N_2305,N_2249,N_2275);
nor U2306 (N_2306,N_2290,N_2211);
or U2307 (N_2307,N_2298,N_2282);
and U2308 (N_2308,N_2236,N_2216);
or U2309 (N_2309,N_2229,N_2256);
nand U2310 (N_2310,N_2208,N_2297);
or U2311 (N_2311,N_2260,N_2253);
xnor U2312 (N_2312,N_2259,N_2213);
nand U2313 (N_2313,N_2222,N_2251);
or U2314 (N_2314,N_2266,N_2294);
xnor U2315 (N_2315,N_2257,N_2201);
or U2316 (N_2316,N_2234,N_2202);
or U2317 (N_2317,N_2239,N_2223);
and U2318 (N_2318,N_2241,N_2295);
and U2319 (N_2319,N_2258,N_2244);
and U2320 (N_2320,N_2235,N_2232);
nand U2321 (N_2321,N_2287,N_2203);
and U2322 (N_2322,N_2267,N_2272);
nor U2323 (N_2323,N_2250,N_2228);
or U2324 (N_2324,N_2224,N_2271);
nand U2325 (N_2325,N_2219,N_2225);
and U2326 (N_2326,N_2263,N_2215);
and U2327 (N_2327,N_2237,N_2220);
or U2328 (N_2328,N_2265,N_2264);
xor U2329 (N_2329,N_2240,N_2284);
and U2330 (N_2330,N_2230,N_2288);
or U2331 (N_2331,N_2247,N_2217);
and U2332 (N_2332,N_2200,N_2261);
and U2333 (N_2333,N_2212,N_2268);
nor U2334 (N_2334,N_2231,N_2281);
or U2335 (N_2335,N_2204,N_2238);
xor U2336 (N_2336,N_2274,N_2248);
or U2337 (N_2337,N_2252,N_2245);
nand U2338 (N_2338,N_2262,N_2270);
or U2339 (N_2339,N_2221,N_2296);
nand U2340 (N_2340,N_2242,N_2299);
nand U2341 (N_2341,N_2255,N_2254);
nand U2342 (N_2342,N_2277,N_2209);
nor U2343 (N_2343,N_2280,N_2276);
xnor U2344 (N_2344,N_2285,N_2227);
xor U2345 (N_2345,N_2293,N_2292);
nand U2346 (N_2346,N_2226,N_2205);
xnor U2347 (N_2347,N_2210,N_2283);
nand U2348 (N_2348,N_2233,N_2246);
xnor U2349 (N_2349,N_2206,N_2286);
nand U2350 (N_2350,N_2211,N_2236);
nor U2351 (N_2351,N_2270,N_2203);
xnor U2352 (N_2352,N_2206,N_2290);
xor U2353 (N_2353,N_2220,N_2274);
and U2354 (N_2354,N_2251,N_2273);
nor U2355 (N_2355,N_2289,N_2249);
nor U2356 (N_2356,N_2245,N_2278);
nand U2357 (N_2357,N_2222,N_2214);
or U2358 (N_2358,N_2286,N_2214);
nor U2359 (N_2359,N_2246,N_2298);
or U2360 (N_2360,N_2235,N_2269);
nand U2361 (N_2361,N_2279,N_2273);
xnor U2362 (N_2362,N_2261,N_2278);
nand U2363 (N_2363,N_2216,N_2288);
or U2364 (N_2364,N_2296,N_2248);
nor U2365 (N_2365,N_2230,N_2287);
or U2366 (N_2366,N_2286,N_2287);
and U2367 (N_2367,N_2288,N_2210);
or U2368 (N_2368,N_2269,N_2280);
nand U2369 (N_2369,N_2288,N_2212);
nor U2370 (N_2370,N_2293,N_2260);
nand U2371 (N_2371,N_2280,N_2263);
and U2372 (N_2372,N_2286,N_2237);
and U2373 (N_2373,N_2208,N_2286);
nand U2374 (N_2374,N_2218,N_2273);
or U2375 (N_2375,N_2287,N_2209);
or U2376 (N_2376,N_2278,N_2249);
nor U2377 (N_2377,N_2285,N_2287);
nand U2378 (N_2378,N_2256,N_2217);
nand U2379 (N_2379,N_2216,N_2299);
nand U2380 (N_2380,N_2275,N_2211);
and U2381 (N_2381,N_2211,N_2262);
nand U2382 (N_2382,N_2207,N_2227);
nand U2383 (N_2383,N_2278,N_2228);
and U2384 (N_2384,N_2208,N_2220);
or U2385 (N_2385,N_2250,N_2288);
or U2386 (N_2386,N_2223,N_2292);
and U2387 (N_2387,N_2279,N_2201);
xnor U2388 (N_2388,N_2221,N_2255);
nand U2389 (N_2389,N_2293,N_2296);
nor U2390 (N_2390,N_2297,N_2236);
xnor U2391 (N_2391,N_2279,N_2267);
nand U2392 (N_2392,N_2295,N_2213);
nand U2393 (N_2393,N_2207,N_2239);
and U2394 (N_2394,N_2231,N_2277);
nand U2395 (N_2395,N_2283,N_2242);
nand U2396 (N_2396,N_2292,N_2287);
nand U2397 (N_2397,N_2261,N_2282);
or U2398 (N_2398,N_2284,N_2290);
nand U2399 (N_2399,N_2217,N_2271);
nor U2400 (N_2400,N_2374,N_2339);
nor U2401 (N_2401,N_2366,N_2306);
or U2402 (N_2402,N_2346,N_2361);
nor U2403 (N_2403,N_2364,N_2349);
nand U2404 (N_2404,N_2344,N_2300);
and U2405 (N_2405,N_2367,N_2304);
xor U2406 (N_2406,N_2336,N_2390);
nor U2407 (N_2407,N_2312,N_2382);
nor U2408 (N_2408,N_2386,N_2393);
and U2409 (N_2409,N_2314,N_2325);
nand U2410 (N_2410,N_2397,N_2381);
nor U2411 (N_2411,N_2353,N_2370);
nand U2412 (N_2412,N_2396,N_2387);
xor U2413 (N_2413,N_2332,N_2376);
nand U2414 (N_2414,N_2362,N_2391);
and U2415 (N_2415,N_2347,N_2340);
or U2416 (N_2416,N_2319,N_2389);
nand U2417 (N_2417,N_2323,N_2365);
or U2418 (N_2418,N_2392,N_2348);
nor U2419 (N_2419,N_2357,N_2302);
nor U2420 (N_2420,N_2341,N_2310);
and U2421 (N_2421,N_2379,N_2345);
xor U2422 (N_2422,N_2315,N_2373);
and U2423 (N_2423,N_2317,N_2399);
or U2424 (N_2424,N_2395,N_2354);
nand U2425 (N_2425,N_2305,N_2383);
or U2426 (N_2426,N_2311,N_2372);
nand U2427 (N_2427,N_2309,N_2359);
and U2428 (N_2428,N_2356,N_2351);
nor U2429 (N_2429,N_2375,N_2355);
nor U2430 (N_2430,N_2394,N_2360);
xnor U2431 (N_2431,N_2385,N_2338);
or U2432 (N_2432,N_2398,N_2380);
nor U2433 (N_2433,N_2331,N_2377);
or U2434 (N_2434,N_2350,N_2328);
or U2435 (N_2435,N_2321,N_2368);
nand U2436 (N_2436,N_2320,N_2333);
nand U2437 (N_2437,N_2307,N_2334);
or U2438 (N_2438,N_2322,N_2303);
and U2439 (N_2439,N_2313,N_2384);
nor U2440 (N_2440,N_2343,N_2329);
and U2441 (N_2441,N_2301,N_2318);
nand U2442 (N_2442,N_2316,N_2335);
xnor U2443 (N_2443,N_2330,N_2337);
nor U2444 (N_2444,N_2358,N_2363);
and U2445 (N_2445,N_2388,N_2342);
and U2446 (N_2446,N_2352,N_2327);
or U2447 (N_2447,N_2308,N_2324);
or U2448 (N_2448,N_2378,N_2326);
nand U2449 (N_2449,N_2369,N_2371);
nand U2450 (N_2450,N_2392,N_2399);
nand U2451 (N_2451,N_2378,N_2352);
or U2452 (N_2452,N_2312,N_2346);
xnor U2453 (N_2453,N_2384,N_2322);
xor U2454 (N_2454,N_2318,N_2331);
and U2455 (N_2455,N_2379,N_2347);
or U2456 (N_2456,N_2375,N_2319);
xnor U2457 (N_2457,N_2350,N_2396);
xor U2458 (N_2458,N_2386,N_2312);
xor U2459 (N_2459,N_2368,N_2332);
nor U2460 (N_2460,N_2342,N_2306);
xnor U2461 (N_2461,N_2339,N_2353);
and U2462 (N_2462,N_2306,N_2321);
or U2463 (N_2463,N_2348,N_2342);
or U2464 (N_2464,N_2379,N_2310);
and U2465 (N_2465,N_2353,N_2313);
and U2466 (N_2466,N_2364,N_2312);
nand U2467 (N_2467,N_2396,N_2308);
nand U2468 (N_2468,N_2369,N_2302);
nor U2469 (N_2469,N_2335,N_2387);
xor U2470 (N_2470,N_2318,N_2357);
nor U2471 (N_2471,N_2322,N_2358);
and U2472 (N_2472,N_2327,N_2311);
xnor U2473 (N_2473,N_2379,N_2348);
nor U2474 (N_2474,N_2370,N_2360);
nand U2475 (N_2475,N_2355,N_2397);
or U2476 (N_2476,N_2327,N_2312);
and U2477 (N_2477,N_2386,N_2302);
xor U2478 (N_2478,N_2339,N_2383);
or U2479 (N_2479,N_2399,N_2394);
and U2480 (N_2480,N_2343,N_2385);
xor U2481 (N_2481,N_2337,N_2392);
nand U2482 (N_2482,N_2364,N_2335);
and U2483 (N_2483,N_2379,N_2383);
nand U2484 (N_2484,N_2365,N_2396);
and U2485 (N_2485,N_2346,N_2377);
and U2486 (N_2486,N_2321,N_2340);
xor U2487 (N_2487,N_2302,N_2313);
nand U2488 (N_2488,N_2309,N_2334);
nand U2489 (N_2489,N_2302,N_2355);
xnor U2490 (N_2490,N_2340,N_2364);
nor U2491 (N_2491,N_2333,N_2397);
and U2492 (N_2492,N_2346,N_2376);
and U2493 (N_2493,N_2389,N_2323);
nor U2494 (N_2494,N_2337,N_2387);
and U2495 (N_2495,N_2311,N_2380);
and U2496 (N_2496,N_2331,N_2312);
nand U2497 (N_2497,N_2327,N_2381);
nor U2498 (N_2498,N_2339,N_2307);
nor U2499 (N_2499,N_2331,N_2382);
xor U2500 (N_2500,N_2496,N_2442);
nor U2501 (N_2501,N_2414,N_2450);
xor U2502 (N_2502,N_2446,N_2474);
nand U2503 (N_2503,N_2437,N_2457);
nand U2504 (N_2504,N_2430,N_2472);
and U2505 (N_2505,N_2425,N_2486);
nor U2506 (N_2506,N_2477,N_2440);
nor U2507 (N_2507,N_2408,N_2498);
or U2508 (N_2508,N_2417,N_2497);
nor U2509 (N_2509,N_2462,N_2484);
nor U2510 (N_2510,N_2470,N_2493);
and U2511 (N_2511,N_2404,N_2494);
xor U2512 (N_2512,N_2433,N_2490);
and U2513 (N_2513,N_2482,N_2464);
nand U2514 (N_2514,N_2471,N_2405);
or U2515 (N_2515,N_2469,N_2420);
xnor U2516 (N_2516,N_2441,N_2439);
or U2517 (N_2517,N_2410,N_2436);
nor U2518 (N_2518,N_2427,N_2489);
and U2519 (N_2519,N_2435,N_2478);
and U2520 (N_2520,N_2495,N_2468);
nand U2521 (N_2521,N_2456,N_2480);
xnor U2522 (N_2522,N_2455,N_2445);
nand U2523 (N_2523,N_2466,N_2403);
xor U2524 (N_2524,N_2447,N_2473);
and U2525 (N_2525,N_2487,N_2434);
or U2526 (N_2526,N_2407,N_2421);
and U2527 (N_2527,N_2492,N_2481);
nor U2528 (N_2528,N_2443,N_2451);
nand U2529 (N_2529,N_2406,N_2475);
and U2530 (N_2530,N_2461,N_2409);
and U2531 (N_2531,N_2454,N_2423);
and U2532 (N_2532,N_2449,N_2415);
nand U2533 (N_2533,N_2432,N_2453);
nor U2534 (N_2534,N_2460,N_2438);
xnor U2535 (N_2535,N_2465,N_2428);
and U2536 (N_2536,N_2444,N_2483);
nand U2537 (N_2537,N_2459,N_2416);
xnor U2538 (N_2538,N_2431,N_2452);
nor U2539 (N_2539,N_2491,N_2401);
xnor U2540 (N_2540,N_2485,N_2412);
and U2541 (N_2541,N_2424,N_2488);
nor U2542 (N_2542,N_2476,N_2411);
and U2543 (N_2543,N_2479,N_2448);
or U2544 (N_2544,N_2429,N_2467);
xnor U2545 (N_2545,N_2458,N_2463);
xor U2546 (N_2546,N_2402,N_2422);
and U2547 (N_2547,N_2413,N_2418);
nor U2548 (N_2548,N_2499,N_2400);
nor U2549 (N_2549,N_2419,N_2426);
xor U2550 (N_2550,N_2409,N_2454);
xor U2551 (N_2551,N_2416,N_2468);
nand U2552 (N_2552,N_2458,N_2419);
nand U2553 (N_2553,N_2418,N_2412);
xnor U2554 (N_2554,N_2430,N_2439);
and U2555 (N_2555,N_2460,N_2424);
nand U2556 (N_2556,N_2423,N_2485);
xnor U2557 (N_2557,N_2451,N_2468);
nor U2558 (N_2558,N_2494,N_2487);
xor U2559 (N_2559,N_2411,N_2480);
or U2560 (N_2560,N_2401,N_2445);
nor U2561 (N_2561,N_2418,N_2496);
nor U2562 (N_2562,N_2438,N_2489);
nor U2563 (N_2563,N_2428,N_2480);
or U2564 (N_2564,N_2463,N_2417);
nand U2565 (N_2565,N_2426,N_2450);
nor U2566 (N_2566,N_2488,N_2472);
or U2567 (N_2567,N_2470,N_2483);
and U2568 (N_2568,N_2427,N_2421);
xnor U2569 (N_2569,N_2484,N_2429);
or U2570 (N_2570,N_2477,N_2468);
nand U2571 (N_2571,N_2434,N_2444);
or U2572 (N_2572,N_2470,N_2465);
nand U2573 (N_2573,N_2417,N_2423);
nor U2574 (N_2574,N_2404,N_2471);
and U2575 (N_2575,N_2452,N_2458);
xnor U2576 (N_2576,N_2417,N_2465);
nor U2577 (N_2577,N_2477,N_2421);
nand U2578 (N_2578,N_2458,N_2472);
xor U2579 (N_2579,N_2476,N_2494);
nor U2580 (N_2580,N_2456,N_2423);
xnor U2581 (N_2581,N_2408,N_2489);
nand U2582 (N_2582,N_2451,N_2490);
and U2583 (N_2583,N_2482,N_2404);
xor U2584 (N_2584,N_2432,N_2493);
nand U2585 (N_2585,N_2421,N_2468);
nand U2586 (N_2586,N_2485,N_2415);
nor U2587 (N_2587,N_2430,N_2489);
xnor U2588 (N_2588,N_2457,N_2484);
xor U2589 (N_2589,N_2407,N_2420);
nand U2590 (N_2590,N_2459,N_2406);
nor U2591 (N_2591,N_2400,N_2407);
and U2592 (N_2592,N_2478,N_2465);
nor U2593 (N_2593,N_2421,N_2419);
and U2594 (N_2594,N_2405,N_2469);
xnor U2595 (N_2595,N_2460,N_2426);
nor U2596 (N_2596,N_2436,N_2449);
or U2597 (N_2597,N_2486,N_2404);
or U2598 (N_2598,N_2463,N_2422);
nor U2599 (N_2599,N_2422,N_2434);
and U2600 (N_2600,N_2542,N_2552);
xor U2601 (N_2601,N_2521,N_2514);
and U2602 (N_2602,N_2528,N_2513);
or U2603 (N_2603,N_2595,N_2527);
and U2604 (N_2604,N_2579,N_2570);
nor U2605 (N_2605,N_2532,N_2564);
nand U2606 (N_2606,N_2501,N_2573);
nand U2607 (N_2607,N_2547,N_2529);
nand U2608 (N_2608,N_2538,N_2554);
xnor U2609 (N_2609,N_2559,N_2525);
or U2610 (N_2610,N_2523,N_2586);
nor U2611 (N_2611,N_2583,N_2534);
xor U2612 (N_2612,N_2537,N_2593);
and U2613 (N_2613,N_2594,N_2578);
and U2614 (N_2614,N_2535,N_2591);
nand U2615 (N_2615,N_2510,N_2571);
xor U2616 (N_2616,N_2533,N_2545);
nor U2617 (N_2617,N_2546,N_2589);
xnor U2618 (N_2618,N_2508,N_2590);
xnor U2619 (N_2619,N_2543,N_2530);
nor U2620 (N_2620,N_2516,N_2574);
nor U2621 (N_2621,N_2520,N_2575);
and U2622 (N_2622,N_2522,N_2585);
nor U2623 (N_2623,N_2592,N_2568);
xor U2624 (N_2624,N_2563,N_2597);
or U2625 (N_2625,N_2567,N_2582);
nor U2626 (N_2626,N_2507,N_2556);
xor U2627 (N_2627,N_2549,N_2548);
or U2628 (N_2628,N_2544,N_2515);
nand U2629 (N_2629,N_2511,N_2524);
or U2630 (N_2630,N_2557,N_2531);
and U2631 (N_2631,N_2512,N_2550);
or U2632 (N_2632,N_2598,N_2541);
nand U2633 (N_2633,N_2518,N_2569);
or U2634 (N_2634,N_2503,N_2519);
xor U2635 (N_2635,N_2565,N_2536);
nand U2636 (N_2636,N_2558,N_2504);
nor U2637 (N_2637,N_2584,N_2588);
or U2638 (N_2638,N_2566,N_2555);
xnor U2639 (N_2639,N_2540,N_2572);
xnor U2640 (N_2640,N_2561,N_2596);
nand U2641 (N_2641,N_2553,N_2509);
or U2642 (N_2642,N_2577,N_2587);
or U2643 (N_2643,N_2551,N_2506);
nand U2644 (N_2644,N_2500,N_2581);
xnor U2645 (N_2645,N_2502,N_2576);
nand U2646 (N_2646,N_2560,N_2526);
or U2647 (N_2647,N_2562,N_2517);
nand U2648 (N_2648,N_2505,N_2580);
nor U2649 (N_2649,N_2539,N_2599);
nand U2650 (N_2650,N_2535,N_2540);
or U2651 (N_2651,N_2572,N_2576);
or U2652 (N_2652,N_2523,N_2539);
xor U2653 (N_2653,N_2506,N_2520);
nor U2654 (N_2654,N_2540,N_2514);
nand U2655 (N_2655,N_2552,N_2508);
nor U2656 (N_2656,N_2545,N_2596);
and U2657 (N_2657,N_2575,N_2571);
xor U2658 (N_2658,N_2586,N_2528);
nor U2659 (N_2659,N_2568,N_2544);
and U2660 (N_2660,N_2586,N_2505);
or U2661 (N_2661,N_2584,N_2593);
nor U2662 (N_2662,N_2590,N_2598);
and U2663 (N_2663,N_2520,N_2511);
nor U2664 (N_2664,N_2514,N_2505);
and U2665 (N_2665,N_2554,N_2523);
or U2666 (N_2666,N_2575,N_2534);
nand U2667 (N_2667,N_2538,N_2566);
nor U2668 (N_2668,N_2565,N_2527);
xor U2669 (N_2669,N_2552,N_2574);
nor U2670 (N_2670,N_2524,N_2584);
xor U2671 (N_2671,N_2556,N_2528);
nor U2672 (N_2672,N_2583,N_2516);
or U2673 (N_2673,N_2560,N_2539);
nand U2674 (N_2674,N_2585,N_2546);
nand U2675 (N_2675,N_2561,N_2556);
or U2676 (N_2676,N_2553,N_2564);
nor U2677 (N_2677,N_2519,N_2539);
or U2678 (N_2678,N_2565,N_2594);
and U2679 (N_2679,N_2538,N_2597);
nand U2680 (N_2680,N_2580,N_2546);
or U2681 (N_2681,N_2537,N_2547);
xnor U2682 (N_2682,N_2507,N_2563);
and U2683 (N_2683,N_2543,N_2550);
or U2684 (N_2684,N_2507,N_2578);
xor U2685 (N_2685,N_2512,N_2564);
nand U2686 (N_2686,N_2550,N_2589);
and U2687 (N_2687,N_2544,N_2534);
or U2688 (N_2688,N_2502,N_2595);
xnor U2689 (N_2689,N_2570,N_2508);
and U2690 (N_2690,N_2507,N_2594);
or U2691 (N_2691,N_2578,N_2551);
nand U2692 (N_2692,N_2567,N_2592);
nor U2693 (N_2693,N_2582,N_2537);
and U2694 (N_2694,N_2594,N_2563);
or U2695 (N_2695,N_2561,N_2577);
and U2696 (N_2696,N_2547,N_2562);
nor U2697 (N_2697,N_2501,N_2504);
nand U2698 (N_2698,N_2546,N_2506);
nand U2699 (N_2699,N_2530,N_2541);
nand U2700 (N_2700,N_2653,N_2695);
or U2701 (N_2701,N_2691,N_2675);
nor U2702 (N_2702,N_2628,N_2619);
nand U2703 (N_2703,N_2625,N_2638);
or U2704 (N_2704,N_2613,N_2698);
and U2705 (N_2705,N_2615,N_2665);
nor U2706 (N_2706,N_2602,N_2692);
or U2707 (N_2707,N_2664,N_2643);
nand U2708 (N_2708,N_2603,N_2608);
or U2709 (N_2709,N_2681,N_2611);
nand U2710 (N_2710,N_2690,N_2662);
nand U2711 (N_2711,N_2609,N_2630);
and U2712 (N_2712,N_2605,N_2655);
xor U2713 (N_2713,N_2677,N_2672);
or U2714 (N_2714,N_2657,N_2612);
or U2715 (N_2715,N_2601,N_2680);
and U2716 (N_2716,N_2624,N_2682);
nand U2717 (N_2717,N_2699,N_2614);
and U2718 (N_2718,N_2641,N_2634);
xnor U2719 (N_2719,N_2600,N_2652);
nor U2720 (N_2720,N_2660,N_2658);
and U2721 (N_2721,N_2696,N_2647);
and U2722 (N_2722,N_2642,N_2623);
xor U2723 (N_2723,N_2659,N_2693);
or U2724 (N_2724,N_2648,N_2636);
or U2725 (N_2725,N_2631,N_2678);
xnor U2726 (N_2726,N_2651,N_2670);
and U2727 (N_2727,N_2667,N_2694);
or U2728 (N_2728,N_2635,N_2687);
nor U2729 (N_2729,N_2661,N_2688);
xnor U2730 (N_2730,N_2686,N_2645);
or U2731 (N_2731,N_2666,N_2640);
or U2732 (N_2732,N_2673,N_2679);
and U2733 (N_2733,N_2644,N_2654);
nor U2734 (N_2734,N_2633,N_2650);
and U2735 (N_2735,N_2626,N_2646);
xnor U2736 (N_2736,N_2617,N_2656);
or U2737 (N_2737,N_2676,N_2668);
nor U2738 (N_2738,N_2606,N_2683);
or U2739 (N_2739,N_2620,N_2639);
nor U2740 (N_2740,N_2671,N_2685);
and U2741 (N_2741,N_2697,N_2663);
xor U2742 (N_2742,N_2616,N_2610);
and U2743 (N_2743,N_2632,N_2622);
nand U2744 (N_2744,N_2637,N_2684);
nor U2745 (N_2745,N_2649,N_2618);
or U2746 (N_2746,N_2621,N_2669);
nor U2747 (N_2747,N_2607,N_2627);
xor U2748 (N_2748,N_2629,N_2674);
and U2749 (N_2749,N_2604,N_2689);
or U2750 (N_2750,N_2665,N_2622);
and U2751 (N_2751,N_2614,N_2694);
xnor U2752 (N_2752,N_2647,N_2688);
nor U2753 (N_2753,N_2600,N_2653);
xnor U2754 (N_2754,N_2690,N_2689);
xnor U2755 (N_2755,N_2620,N_2675);
nand U2756 (N_2756,N_2600,N_2612);
or U2757 (N_2757,N_2663,N_2654);
and U2758 (N_2758,N_2692,N_2665);
nor U2759 (N_2759,N_2664,N_2651);
or U2760 (N_2760,N_2689,N_2646);
and U2761 (N_2761,N_2631,N_2685);
or U2762 (N_2762,N_2630,N_2696);
nor U2763 (N_2763,N_2618,N_2662);
and U2764 (N_2764,N_2643,N_2637);
nand U2765 (N_2765,N_2649,N_2619);
and U2766 (N_2766,N_2665,N_2693);
xor U2767 (N_2767,N_2692,N_2613);
xnor U2768 (N_2768,N_2686,N_2644);
xnor U2769 (N_2769,N_2642,N_2606);
and U2770 (N_2770,N_2644,N_2649);
xnor U2771 (N_2771,N_2630,N_2632);
and U2772 (N_2772,N_2654,N_2695);
and U2773 (N_2773,N_2646,N_2675);
nand U2774 (N_2774,N_2609,N_2677);
nand U2775 (N_2775,N_2661,N_2625);
or U2776 (N_2776,N_2632,N_2685);
xor U2777 (N_2777,N_2694,N_2656);
and U2778 (N_2778,N_2675,N_2665);
or U2779 (N_2779,N_2694,N_2651);
and U2780 (N_2780,N_2679,N_2664);
and U2781 (N_2781,N_2618,N_2691);
nand U2782 (N_2782,N_2695,N_2688);
nor U2783 (N_2783,N_2686,N_2624);
nor U2784 (N_2784,N_2609,N_2645);
nor U2785 (N_2785,N_2606,N_2660);
or U2786 (N_2786,N_2685,N_2629);
nor U2787 (N_2787,N_2609,N_2666);
nor U2788 (N_2788,N_2670,N_2603);
nor U2789 (N_2789,N_2659,N_2684);
nand U2790 (N_2790,N_2615,N_2683);
or U2791 (N_2791,N_2641,N_2652);
xnor U2792 (N_2792,N_2648,N_2630);
and U2793 (N_2793,N_2692,N_2696);
or U2794 (N_2794,N_2614,N_2669);
xnor U2795 (N_2795,N_2613,N_2694);
nor U2796 (N_2796,N_2614,N_2665);
nor U2797 (N_2797,N_2609,N_2675);
nor U2798 (N_2798,N_2690,N_2628);
nand U2799 (N_2799,N_2631,N_2690);
xor U2800 (N_2800,N_2793,N_2781);
and U2801 (N_2801,N_2741,N_2757);
nor U2802 (N_2802,N_2724,N_2768);
or U2803 (N_2803,N_2705,N_2771);
xor U2804 (N_2804,N_2790,N_2745);
nor U2805 (N_2805,N_2716,N_2719);
xor U2806 (N_2806,N_2775,N_2730);
nor U2807 (N_2807,N_2792,N_2780);
xor U2808 (N_2808,N_2795,N_2782);
and U2809 (N_2809,N_2744,N_2772);
or U2810 (N_2810,N_2788,N_2785);
xnor U2811 (N_2811,N_2715,N_2706);
xor U2812 (N_2812,N_2787,N_2753);
or U2813 (N_2813,N_2764,N_2798);
or U2814 (N_2814,N_2770,N_2761);
xor U2815 (N_2815,N_2769,N_2742);
nor U2816 (N_2816,N_2739,N_2709);
or U2817 (N_2817,N_2784,N_2794);
xor U2818 (N_2818,N_2754,N_2731);
or U2819 (N_2819,N_2763,N_2776);
or U2820 (N_2820,N_2701,N_2735);
nor U2821 (N_2821,N_2760,N_2750);
and U2822 (N_2822,N_2796,N_2756);
xor U2823 (N_2823,N_2729,N_2762);
nor U2824 (N_2824,N_2710,N_2728);
nor U2825 (N_2825,N_2778,N_2789);
nor U2826 (N_2826,N_2767,N_2717);
nand U2827 (N_2827,N_2725,N_2783);
and U2828 (N_2828,N_2747,N_2743);
nand U2829 (N_2829,N_2774,N_2714);
xnor U2830 (N_2830,N_2732,N_2777);
xnor U2831 (N_2831,N_2713,N_2726);
nand U2832 (N_2832,N_2702,N_2736);
nand U2833 (N_2833,N_2765,N_2720);
and U2834 (N_2834,N_2700,N_2738);
or U2835 (N_2835,N_2759,N_2799);
nor U2836 (N_2836,N_2734,N_2727);
or U2837 (N_2837,N_2786,N_2797);
and U2838 (N_2838,N_2718,N_2749);
nor U2839 (N_2839,N_2748,N_2791);
xor U2840 (N_2840,N_2751,N_2755);
or U2841 (N_2841,N_2708,N_2703);
and U2842 (N_2842,N_2773,N_2733);
nand U2843 (N_2843,N_2723,N_2758);
and U2844 (N_2844,N_2737,N_2711);
or U2845 (N_2845,N_2752,N_2722);
xor U2846 (N_2846,N_2721,N_2766);
and U2847 (N_2847,N_2779,N_2707);
xnor U2848 (N_2848,N_2704,N_2712);
nand U2849 (N_2849,N_2740,N_2746);
and U2850 (N_2850,N_2710,N_2733);
nand U2851 (N_2851,N_2794,N_2795);
or U2852 (N_2852,N_2782,N_2789);
nor U2853 (N_2853,N_2721,N_2705);
and U2854 (N_2854,N_2750,N_2741);
nor U2855 (N_2855,N_2776,N_2725);
xor U2856 (N_2856,N_2727,N_2705);
xor U2857 (N_2857,N_2714,N_2752);
nor U2858 (N_2858,N_2754,N_2719);
or U2859 (N_2859,N_2710,N_2797);
nor U2860 (N_2860,N_2714,N_2777);
and U2861 (N_2861,N_2797,N_2793);
or U2862 (N_2862,N_2745,N_2775);
nand U2863 (N_2863,N_2784,N_2782);
or U2864 (N_2864,N_2761,N_2768);
or U2865 (N_2865,N_2761,N_2719);
nor U2866 (N_2866,N_2729,N_2727);
nor U2867 (N_2867,N_2785,N_2750);
xnor U2868 (N_2868,N_2746,N_2773);
xor U2869 (N_2869,N_2708,N_2719);
or U2870 (N_2870,N_2730,N_2717);
nor U2871 (N_2871,N_2730,N_2737);
and U2872 (N_2872,N_2737,N_2772);
xor U2873 (N_2873,N_2778,N_2779);
xor U2874 (N_2874,N_2788,N_2753);
and U2875 (N_2875,N_2742,N_2727);
and U2876 (N_2876,N_2748,N_2708);
or U2877 (N_2877,N_2792,N_2700);
or U2878 (N_2878,N_2768,N_2742);
xnor U2879 (N_2879,N_2704,N_2708);
nand U2880 (N_2880,N_2730,N_2702);
nor U2881 (N_2881,N_2753,N_2701);
or U2882 (N_2882,N_2797,N_2791);
and U2883 (N_2883,N_2713,N_2740);
xor U2884 (N_2884,N_2703,N_2799);
or U2885 (N_2885,N_2743,N_2737);
or U2886 (N_2886,N_2781,N_2715);
and U2887 (N_2887,N_2796,N_2735);
or U2888 (N_2888,N_2702,N_2780);
and U2889 (N_2889,N_2793,N_2760);
or U2890 (N_2890,N_2732,N_2783);
nor U2891 (N_2891,N_2738,N_2790);
xnor U2892 (N_2892,N_2773,N_2771);
or U2893 (N_2893,N_2776,N_2741);
nand U2894 (N_2894,N_2750,N_2702);
xor U2895 (N_2895,N_2703,N_2783);
nand U2896 (N_2896,N_2752,N_2796);
xnor U2897 (N_2897,N_2704,N_2784);
xnor U2898 (N_2898,N_2767,N_2739);
nor U2899 (N_2899,N_2750,N_2773);
and U2900 (N_2900,N_2886,N_2805);
or U2901 (N_2901,N_2815,N_2887);
nand U2902 (N_2902,N_2807,N_2800);
and U2903 (N_2903,N_2846,N_2810);
and U2904 (N_2904,N_2814,N_2879);
nand U2905 (N_2905,N_2889,N_2861);
xnor U2906 (N_2906,N_2851,N_2874);
and U2907 (N_2907,N_2897,N_2863);
or U2908 (N_2908,N_2820,N_2848);
and U2909 (N_2909,N_2894,N_2839);
and U2910 (N_2910,N_2817,N_2806);
or U2911 (N_2911,N_2836,N_2808);
and U2912 (N_2912,N_2816,N_2843);
or U2913 (N_2913,N_2804,N_2835);
and U2914 (N_2914,N_2838,N_2827);
nand U2915 (N_2915,N_2802,N_2898);
xnor U2916 (N_2916,N_2882,N_2825);
xnor U2917 (N_2917,N_2855,N_2883);
xnor U2918 (N_2918,N_2842,N_2828);
or U2919 (N_2919,N_2875,N_2840);
xor U2920 (N_2920,N_2858,N_2864);
xnor U2921 (N_2921,N_2803,N_2892);
or U2922 (N_2922,N_2852,N_2818);
or U2923 (N_2923,N_2826,N_2868);
xor U2924 (N_2924,N_2878,N_2896);
or U2925 (N_2925,N_2873,N_2860);
nand U2926 (N_2926,N_2819,N_2844);
and U2927 (N_2927,N_2823,N_2821);
nand U2928 (N_2928,N_2811,N_2831);
and U2929 (N_2929,N_2881,N_2893);
and U2930 (N_2930,N_2862,N_2877);
and U2931 (N_2931,N_2841,N_2872);
nor U2932 (N_2932,N_2869,N_2870);
or U2933 (N_2933,N_2890,N_2834);
or U2934 (N_2934,N_2809,N_2884);
xnor U2935 (N_2935,N_2880,N_2833);
xor U2936 (N_2936,N_2876,N_2871);
xnor U2937 (N_2937,N_2857,N_2899);
or U2938 (N_2938,N_2885,N_2837);
nor U2939 (N_2939,N_2824,N_2854);
nor U2940 (N_2940,N_2856,N_2891);
or U2941 (N_2941,N_2895,N_2801);
xor U2942 (N_2942,N_2866,N_2830);
nor U2943 (N_2943,N_2812,N_2859);
xor U2944 (N_2944,N_2849,N_2829);
nand U2945 (N_2945,N_2865,N_2822);
and U2946 (N_2946,N_2832,N_2867);
xor U2947 (N_2947,N_2853,N_2847);
or U2948 (N_2948,N_2813,N_2845);
nor U2949 (N_2949,N_2850,N_2888);
and U2950 (N_2950,N_2890,N_2887);
and U2951 (N_2951,N_2881,N_2862);
and U2952 (N_2952,N_2832,N_2890);
or U2953 (N_2953,N_2811,N_2886);
and U2954 (N_2954,N_2874,N_2885);
nor U2955 (N_2955,N_2808,N_2834);
and U2956 (N_2956,N_2858,N_2867);
or U2957 (N_2957,N_2815,N_2855);
nand U2958 (N_2958,N_2873,N_2844);
nand U2959 (N_2959,N_2813,N_2818);
or U2960 (N_2960,N_2853,N_2843);
or U2961 (N_2961,N_2873,N_2800);
or U2962 (N_2962,N_2827,N_2800);
nor U2963 (N_2963,N_2879,N_2806);
or U2964 (N_2964,N_2827,N_2832);
nor U2965 (N_2965,N_2884,N_2850);
or U2966 (N_2966,N_2868,N_2869);
nor U2967 (N_2967,N_2859,N_2800);
nand U2968 (N_2968,N_2824,N_2828);
or U2969 (N_2969,N_2882,N_2843);
and U2970 (N_2970,N_2871,N_2893);
nor U2971 (N_2971,N_2810,N_2889);
or U2972 (N_2972,N_2827,N_2822);
nand U2973 (N_2973,N_2800,N_2871);
or U2974 (N_2974,N_2888,N_2838);
or U2975 (N_2975,N_2847,N_2890);
nand U2976 (N_2976,N_2846,N_2855);
nor U2977 (N_2977,N_2821,N_2879);
and U2978 (N_2978,N_2824,N_2862);
or U2979 (N_2979,N_2838,N_2884);
and U2980 (N_2980,N_2805,N_2834);
and U2981 (N_2981,N_2838,N_2832);
or U2982 (N_2982,N_2846,N_2826);
and U2983 (N_2983,N_2860,N_2839);
or U2984 (N_2984,N_2809,N_2855);
xor U2985 (N_2985,N_2861,N_2856);
and U2986 (N_2986,N_2886,N_2894);
and U2987 (N_2987,N_2891,N_2849);
nor U2988 (N_2988,N_2848,N_2822);
nor U2989 (N_2989,N_2890,N_2843);
nor U2990 (N_2990,N_2801,N_2881);
and U2991 (N_2991,N_2822,N_2874);
and U2992 (N_2992,N_2823,N_2826);
nand U2993 (N_2993,N_2824,N_2883);
nand U2994 (N_2994,N_2885,N_2875);
nor U2995 (N_2995,N_2846,N_2866);
nand U2996 (N_2996,N_2840,N_2882);
or U2997 (N_2997,N_2817,N_2893);
nor U2998 (N_2998,N_2801,N_2886);
or U2999 (N_2999,N_2876,N_2849);
and U3000 (N_3000,N_2914,N_2912);
nor U3001 (N_3001,N_2906,N_2989);
or U3002 (N_3002,N_2939,N_2902);
nor U3003 (N_3003,N_2997,N_2901);
and U3004 (N_3004,N_2941,N_2938);
xor U3005 (N_3005,N_2961,N_2958);
nand U3006 (N_3006,N_2983,N_2991);
nand U3007 (N_3007,N_2976,N_2969);
and U3008 (N_3008,N_2920,N_2949);
xnor U3009 (N_3009,N_2927,N_2911);
nor U3010 (N_3010,N_2947,N_2979);
nor U3011 (N_3011,N_2951,N_2913);
nor U3012 (N_3012,N_2972,N_2974);
nor U3013 (N_3013,N_2928,N_2978);
nor U3014 (N_3014,N_2904,N_2909);
and U3015 (N_3015,N_2937,N_2999);
nor U3016 (N_3016,N_2995,N_2998);
xnor U3017 (N_3017,N_2944,N_2964);
nand U3018 (N_3018,N_2953,N_2971);
and U3019 (N_3019,N_2903,N_2933);
nand U3020 (N_3020,N_2988,N_2929);
or U3021 (N_3021,N_2984,N_2955);
and U3022 (N_3022,N_2919,N_2977);
nor U3023 (N_3023,N_2946,N_2948);
xor U3024 (N_3024,N_2918,N_2963);
nand U3025 (N_3025,N_2923,N_2952);
and U3026 (N_3026,N_2966,N_2985);
nor U3027 (N_3027,N_2956,N_2930);
nor U3028 (N_3028,N_2996,N_2987);
xor U3029 (N_3029,N_2954,N_2926);
nor U3030 (N_3030,N_2916,N_2960);
nor U3031 (N_3031,N_2950,N_2915);
xnor U3032 (N_3032,N_2982,N_2965);
and U3033 (N_3033,N_2917,N_2921);
nand U3034 (N_3034,N_2970,N_2968);
or U3035 (N_3035,N_2900,N_2967);
nor U3036 (N_3036,N_2994,N_2993);
or U3037 (N_3037,N_2935,N_2905);
nor U3038 (N_3038,N_2910,N_2936);
and U3039 (N_3039,N_2975,N_2934);
or U3040 (N_3040,N_2962,N_2980);
nand U3041 (N_3041,N_2943,N_2940);
and U3042 (N_3042,N_2959,N_2986);
and U3043 (N_3043,N_2990,N_2931);
or U3044 (N_3044,N_2942,N_2945);
xor U3045 (N_3045,N_2932,N_2924);
or U3046 (N_3046,N_2957,N_2925);
nor U3047 (N_3047,N_2907,N_2981);
xnor U3048 (N_3048,N_2973,N_2922);
nor U3049 (N_3049,N_2992,N_2908);
xor U3050 (N_3050,N_2921,N_2980);
or U3051 (N_3051,N_2975,N_2935);
xor U3052 (N_3052,N_2912,N_2996);
nand U3053 (N_3053,N_2920,N_2993);
and U3054 (N_3054,N_2904,N_2969);
xnor U3055 (N_3055,N_2918,N_2916);
or U3056 (N_3056,N_2964,N_2986);
or U3057 (N_3057,N_2994,N_2988);
and U3058 (N_3058,N_2930,N_2937);
xor U3059 (N_3059,N_2963,N_2939);
nand U3060 (N_3060,N_2906,N_2943);
and U3061 (N_3061,N_2906,N_2973);
nor U3062 (N_3062,N_2926,N_2960);
xnor U3063 (N_3063,N_2999,N_2924);
xor U3064 (N_3064,N_2934,N_2990);
nand U3065 (N_3065,N_2935,N_2902);
or U3066 (N_3066,N_2967,N_2912);
xnor U3067 (N_3067,N_2958,N_2908);
and U3068 (N_3068,N_2974,N_2967);
nor U3069 (N_3069,N_2941,N_2989);
nor U3070 (N_3070,N_2941,N_2964);
nor U3071 (N_3071,N_2988,N_2962);
nand U3072 (N_3072,N_2919,N_2987);
xor U3073 (N_3073,N_2954,N_2915);
or U3074 (N_3074,N_2994,N_2909);
nor U3075 (N_3075,N_2960,N_2989);
nor U3076 (N_3076,N_2920,N_2924);
nor U3077 (N_3077,N_2927,N_2929);
nor U3078 (N_3078,N_2955,N_2961);
nand U3079 (N_3079,N_2940,N_2915);
nor U3080 (N_3080,N_2966,N_2987);
and U3081 (N_3081,N_2976,N_2913);
xnor U3082 (N_3082,N_2972,N_2901);
and U3083 (N_3083,N_2943,N_2929);
xor U3084 (N_3084,N_2958,N_2906);
nand U3085 (N_3085,N_2982,N_2916);
or U3086 (N_3086,N_2935,N_2984);
or U3087 (N_3087,N_2954,N_2925);
and U3088 (N_3088,N_2929,N_2984);
nand U3089 (N_3089,N_2996,N_2903);
xor U3090 (N_3090,N_2984,N_2946);
xnor U3091 (N_3091,N_2942,N_2990);
xor U3092 (N_3092,N_2943,N_2989);
or U3093 (N_3093,N_2981,N_2955);
or U3094 (N_3094,N_2937,N_2964);
nor U3095 (N_3095,N_2969,N_2980);
nor U3096 (N_3096,N_2916,N_2942);
nand U3097 (N_3097,N_2911,N_2948);
or U3098 (N_3098,N_2978,N_2941);
xor U3099 (N_3099,N_2986,N_2953);
xor U3100 (N_3100,N_3038,N_3096);
xnor U3101 (N_3101,N_3075,N_3048);
nor U3102 (N_3102,N_3025,N_3089);
or U3103 (N_3103,N_3024,N_3018);
xnor U3104 (N_3104,N_3019,N_3031);
nand U3105 (N_3105,N_3091,N_3028);
nand U3106 (N_3106,N_3065,N_3036);
and U3107 (N_3107,N_3084,N_3078);
nor U3108 (N_3108,N_3087,N_3030);
and U3109 (N_3109,N_3016,N_3098);
or U3110 (N_3110,N_3070,N_3034);
nand U3111 (N_3111,N_3040,N_3077);
xor U3112 (N_3112,N_3097,N_3041);
or U3113 (N_3113,N_3014,N_3085);
or U3114 (N_3114,N_3023,N_3076);
nand U3115 (N_3115,N_3003,N_3061);
nand U3116 (N_3116,N_3063,N_3073);
and U3117 (N_3117,N_3022,N_3064);
or U3118 (N_3118,N_3039,N_3050);
nor U3119 (N_3119,N_3035,N_3049);
or U3120 (N_3120,N_3037,N_3008);
nand U3121 (N_3121,N_3046,N_3043);
and U3122 (N_3122,N_3010,N_3099);
nand U3123 (N_3123,N_3042,N_3072);
or U3124 (N_3124,N_3068,N_3090);
xor U3125 (N_3125,N_3000,N_3088);
nand U3126 (N_3126,N_3007,N_3006);
nand U3127 (N_3127,N_3067,N_3059);
nand U3128 (N_3128,N_3071,N_3029);
or U3129 (N_3129,N_3047,N_3079);
xor U3130 (N_3130,N_3045,N_3086);
nor U3131 (N_3131,N_3001,N_3095);
xor U3132 (N_3132,N_3094,N_3082);
or U3133 (N_3133,N_3056,N_3062);
and U3134 (N_3134,N_3069,N_3012);
nand U3135 (N_3135,N_3058,N_3032);
xnor U3136 (N_3136,N_3080,N_3011);
and U3137 (N_3137,N_3017,N_3004);
or U3138 (N_3138,N_3020,N_3033);
nand U3139 (N_3139,N_3066,N_3054);
nor U3140 (N_3140,N_3002,N_3005);
xor U3141 (N_3141,N_3053,N_3013);
and U3142 (N_3142,N_3027,N_3083);
or U3143 (N_3143,N_3051,N_3093);
nor U3144 (N_3144,N_3015,N_3081);
nand U3145 (N_3145,N_3057,N_3009);
or U3146 (N_3146,N_3092,N_3060);
nand U3147 (N_3147,N_3044,N_3021);
nor U3148 (N_3148,N_3074,N_3052);
xor U3149 (N_3149,N_3026,N_3055);
and U3150 (N_3150,N_3062,N_3028);
nor U3151 (N_3151,N_3057,N_3023);
nor U3152 (N_3152,N_3075,N_3092);
and U3153 (N_3153,N_3002,N_3025);
and U3154 (N_3154,N_3084,N_3095);
nand U3155 (N_3155,N_3050,N_3001);
nand U3156 (N_3156,N_3032,N_3034);
or U3157 (N_3157,N_3020,N_3030);
xor U3158 (N_3158,N_3060,N_3013);
nor U3159 (N_3159,N_3005,N_3043);
xor U3160 (N_3160,N_3051,N_3052);
xor U3161 (N_3161,N_3055,N_3041);
nand U3162 (N_3162,N_3025,N_3027);
nor U3163 (N_3163,N_3097,N_3074);
nand U3164 (N_3164,N_3002,N_3087);
nand U3165 (N_3165,N_3015,N_3013);
and U3166 (N_3166,N_3090,N_3060);
nor U3167 (N_3167,N_3004,N_3088);
and U3168 (N_3168,N_3080,N_3084);
or U3169 (N_3169,N_3068,N_3029);
nand U3170 (N_3170,N_3071,N_3063);
and U3171 (N_3171,N_3090,N_3083);
nor U3172 (N_3172,N_3021,N_3082);
and U3173 (N_3173,N_3090,N_3035);
xnor U3174 (N_3174,N_3031,N_3012);
nand U3175 (N_3175,N_3043,N_3077);
or U3176 (N_3176,N_3093,N_3066);
nor U3177 (N_3177,N_3062,N_3035);
nand U3178 (N_3178,N_3097,N_3019);
xor U3179 (N_3179,N_3007,N_3077);
and U3180 (N_3180,N_3040,N_3032);
or U3181 (N_3181,N_3015,N_3083);
or U3182 (N_3182,N_3095,N_3059);
nor U3183 (N_3183,N_3077,N_3071);
and U3184 (N_3184,N_3013,N_3080);
nor U3185 (N_3185,N_3036,N_3083);
nand U3186 (N_3186,N_3077,N_3039);
xor U3187 (N_3187,N_3070,N_3041);
and U3188 (N_3188,N_3062,N_3018);
nand U3189 (N_3189,N_3021,N_3054);
nor U3190 (N_3190,N_3044,N_3031);
xor U3191 (N_3191,N_3049,N_3023);
or U3192 (N_3192,N_3009,N_3040);
nor U3193 (N_3193,N_3026,N_3025);
xnor U3194 (N_3194,N_3094,N_3050);
xor U3195 (N_3195,N_3023,N_3091);
or U3196 (N_3196,N_3073,N_3026);
xor U3197 (N_3197,N_3056,N_3009);
nand U3198 (N_3198,N_3067,N_3017);
nor U3199 (N_3199,N_3001,N_3073);
xnor U3200 (N_3200,N_3111,N_3121);
nor U3201 (N_3201,N_3138,N_3186);
nor U3202 (N_3202,N_3146,N_3159);
nor U3203 (N_3203,N_3127,N_3134);
xnor U3204 (N_3204,N_3101,N_3113);
or U3205 (N_3205,N_3118,N_3175);
or U3206 (N_3206,N_3135,N_3158);
nor U3207 (N_3207,N_3173,N_3116);
xnor U3208 (N_3208,N_3161,N_3130);
and U3209 (N_3209,N_3176,N_3107);
nor U3210 (N_3210,N_3165,N_3122);
nand U3211 (N_3211,N_3126,N_3151);
or U3212 (N_3212,N_3199,N_3196);
nand U3213 (N_3213,N_3168,N_3166);
nor U3214 (N_3214,N_3109,N_3124);
nand U3215 (N_3215,N_3189,N_3147);
nand U3216 (N_3216,N_3190,N_3160);
xor U3217 (N_3217,N_3155,N_3100);
and U3218 (N_3218,N_3184,N_3174);
or U3219 (N_3219,N_3178,N_3110);
xor U3220 (N_3220,N_3195,N_3164);
nor U3221 (N_3221,N_3150,N_3177);
xor U3222 (N_3222,N_3163,N_3180);
or U3223 (N_3223,N_3115,N_3132);
nand U3224 (N_3224,N_3137,N_3167);
nor U3225 (N_3225,N_3171,N_3198);
or U3226 (N_3226,N_3152,N_3191);
and U3227 (N_3227,N_3153,N_3103);
nand U3228 (N_3228,N_3154,N_3106);
nor U3229 (N_3229,N_3120,N_3162);
nor U3230 (N_3230,N_3123,N_3143);
nand U3231 (N_3231,N_3185,N_3192);
xor U3232 (N_3232,N_3187,N_3170);
nor U3233 (N_3233,N_3157,N_3193);
and U3234 (N_3234,N_3125,N_3181);
xnor U3235 (N_3235,N_3182,N_3114);
nor U3236 (N_3236,N_3188,N_3179);
and U3237 (N_3237,N_3129,N_3128);
xnor U3238 (N_3238,N_3145,N_3131);
and U3239 (N_3239,N_3136,N_3139);
nand U3240 (N_3240,N_3169,N_3149);
xnor U3241 (N_3241,N_3133,N_3112);
nand U3242 (N_3242,N_3108,N_3141);
nor U3243 (N_3243,N_3144,N_3172);
or U3244 (N_3244,N_3142,N_3183);
nor U3245 (N_3245,N_3117,N_3156);
or U3246 (N_3246,N_3104,N_3102);
xor U3247 (N_3247,N_3148,N_3197);
and U3248 (N_3248,N_3119,N_3194);
xnor U3249 (N_3249,N_3140,N_3105);
or U3250 (N_3250,N_3184,N_3194);
or U3251 (N_3251,N_3117,N_3116);
nand U3252 (N_3252,N_3167,N_3171);
nor U3253 (N_3253,N_3143,N_3112);
nor U3254 (N_3254,N_3128,N_3162);
nor U3255 (N_3255,N_3132,N_3119);
nor U3256 (N_3256,N_3123,N_3117);
nor U3257 (N_3257,N_3107,N_3194);
and U3258 (N_3258,N_3174,N_3157);
and U3259 (N_3259,N_3180,N_3115);
or U3260 (N_3260,N_3196,N_3193);
xnor U3261 (N_3261,N_3109,N_3130);
and U3262 (N_3262,N_3145,N_3116);
xnor U3263 (N_3263,N_3116,N_3129);
nand U3264 (N_3264,N_3180,N_3154);
nor U3265 (N_3265,N_3155,N_3160);
nor U3266 (N_3266,N_3142,N_3173);
xor U3267 (N_3267,N_3169,N_3152);
nand U3268 (N_3268,N_3165,N_3175);
and U3269 (N_3269,N_3189,N_3144);
or U3270 (N_3270,N_3180,N_3108);
or U3271 (N_3271,N_3142,N_3139);
nand U3272 (N_3272,N_3159,N_3152);
nor U3273 (N_3273,N_3162,N_3142);
or U3274 (N_3274,N_3131,N_3106);
or U3275 (N_3275,N_3133,N_3192);
nand U3276 (N_3276,N_3154,N_3177);
nand U3277 (N_3277,N_3120,N_3157);
nand U3278 (N_3278,N_3140,N_3126);
or U3279 (N_3279,N_3107,N_3154);
or U3280 (N_3280,N_3129,N_3115);
and U3281 (N_3281,N_3130,N_3166);
nand U3282 (N_3282,N_3162,N_3194);
nor U3283 (N_3283,N_3147,N_3179);
and U3284 (N_3284,N_3157,N_3127);
or U3285 (N_3285,N_3156,N_3122);
or U3286 (N_3286,N_3117,N_3110);
nor U3287 (N_3287,N_3103,N_3140);
xor U3288 (N_3288,N_3192,N_3110);
nand U3289 (N_3289,N_3170,N_3179);
nor U3290 (N_3290,N_3106,N_3137);
nor U3291 (N_3291,N_3169,N_3178);
xor U3292 (N_3292,N_3153,N_3150);
and U3293 (N_3293,N_3146,N_3184);
or U3294 (N_3294,N_3123,N_3163);
nand U3295 (N_3295,N_3108,N_3153);
nand U3296 (N_3296,N_3139,N_3104);
or U3297 (N_3297,N_3172,N_3126);
and U3298 (N_3298,N_3142,N_3158);
and U3299 (N_3299,N_3180,N_3199);
nand U3300 (N_3300,N_3275,N_3213);
xnor U3301 (N_3301,N_3227,N_3287);
nor U3302 (N_3302,N_3209,N_3214);
xor U3303 (N_3303,N_3242,N_3247);
nor U3304 (N_3304,N_3230,N_3284);
and U3305 (N_3305,N_3286,N_3244);
and U3306 (N_3306,N_3257,N_3238);
nor U3307 (N_3307,N_3277,N_3218);
and U3308 (N_3308,N_3228,N_3215);
and U3309 (N_3309,N_3240,N_3296);
nand U3310 (N_3310,N_3288,N_3256);
or U3311 (N_3311,N_3269,N_3272);
and U3312 (N_3312,N_3236,N_3252);
and U3313 (N_3313,N_3262,N_3232);
and U3314 (N_3314,N_3205,N_3276);
nand U3315 (N_3315,N_3229,N_3204);
or U3316 (N_3316,N_3251,N_3285);
xnor U3317 (N_3317,N_3221,N_3239);
or U3318 (N_3318,N_3267,N_3294);
xor U3319 (N_3319,N_3261,N_3278);
and U3320 (N_3320,N_3270,N_3297);
nand U3321 (N_3321,N_3233,N_3219);
or U3322 (N_3322,N_3206,N_3279);
and U3323 (N_3323,N_3241,N_3217);
and U3324 (N_3324,N_3225,N_3282);
and U3325 (N_3325,N_3211,N_3200);
xnor U3326 (N_3326,N_3243,N_3290);
or U3327 (N_3327,N_3299,N_3203);
or U3328 (N_3328,N_3255,N_3268);
nor U3329 (N_3329,N_3246,N_3281);
nor U3330 (N_3330,N_3210,N_3292);
and U3331 (N_3331,N_3259,N_3298);
nand U3332 (N_3332,N_3216,N_3264);
or U3333 (N_3333,N_3291,N_3235);
or U3334 (N_3334,N_3283,N_3212);
and U3335 (N_3335,N_3245,N_3266);
nand U3336 (N_3336,N_3224,N_3253);
nor U3337 (N_3337,N_3207,N_3208);
xor U3338 (N_3338,N_3271,N_3280);
nor U3339 (N_3339,N_3295,N_3234);
or U3340 (N_3340,N_3254,N_3274);
and U3341 (N_3341,N_3220,N_3263);
and U3342 (N_3342,N_3265,N_3258);
nand U3343 (N_3343,N_3202,N_3222);
nor U3344 (N_3344,N_3248,N_3260);
or U3345 (N_3345,N_3250,N_3273);
nor U3346 (N_3346,N_3249,N_3226);
or U3347 (N_3347,N_3289,N_3231);
and U3348 (N_3348,N_3201,N_3293);
nand U3349 (N_3349,N_3237,N_3223);
and U3350 (N_3350,N_3206,N_3232);
or U3351 (N_3351,N_3297,N_3267);
or U3352 (N_3352,N_3203,N_3279);
nor U3353 (N_3353,N_3285,N_3289);
nor U3354 (N_3354,N_3247,N_3238);
and U3355 (N_3355,N_3228,N_3292);
xnor U3356 (N_3356,N_3218,N_3282);
xor U3357 (N_3357,N_3273,N_3242);
and U3358 (N_3358,N_3239,N_3289);
xnor U3359 (N_3359,N_3217,N_3246);
and U3360 (N_3360,N_3287,N_3226);
xnor U3361 (N_3361,N_3244,N_3260);
nor U3362 (N_3362,N_3255,N_3286);
or U3363 (N_3363,N_3209,N_3283);
nor U3364 (N_3364,N_3268,N_3269);
and U3365 (N_3365,N_3256,N_3278);
nand U3366 (N_3366,N_3297,N_3280);
xor U3367 (N_3367,N_3239,N_3271);
or U3368 (N_3368,N_3230,N_3239);
nor U3369 (N_3369,N_3255,N_3220);
and U3370 (N_3370,N_3298,N_3204);
nor U3371 (N_3371,N_3287,N_3277);
xor U3372 (N_3372,N_3231,N_3211);
nor U3373 (N_3373,N_3248,N_3213);
xnor U3374 (N_3374,N_3232,N_3221);
nand U3375 (N_3375,N_3291,N_3214);
nor U3376 (N_3376,N_3289,N_3220);
and U3377 (N_3377,N_3204,N_3214);
xor U3378 (N_3378,N_3255,N_3259);
or U3379 (N_3379,N_3280,N_3268);
nor U3380 (N_3380,N_3235,N_3268);
and U3381 (N_3381,N_3249,N_3246);
xor U3382 (N_3382,N_3274,N_3220);
or U3383 (N_3383,N_3292,N_3274);
nor U3384 (N_3384,N_3296,N_3208);
nor U3385 (N_3385,N_3263,N_3232);
nand U3386 (N_3386,N_3291,N_3299);
nor U3387 (N_3387,N_3263,N_3267);
nand U3388 (N_3388,N_3225,N_3276);
xnor U3389 (N_3389,N_3215,N_3275);
or U3390 (N_3390,N_3200,N_3271);
nand U3391 (N_3391,N_3247,N_3287);
nand U3392 (N_3392,N_3281,N_3259);
or U3393 (N_3393,N_3287,N_3255);
xor U3394 (N_3394,N_3225,N_3253);
nor U3395 (N_3395,N_3270,N_3259);
and U3396 (N_3396,N_3224,N_3203);
nand U3397 (N_3397,N_3217,N_3286);
and U3398 (N_3398,N_3296,N_3201);
xnor U3399 (N_3399,N_3244,N_3246);
nor U3400 (N_3400,N_3392,N_3368);
or U3401 (N_3401,N_3335,N_3301);
or U3402 (N_3402,N_3320,N_3378);
xnor U3403 (N_3403,N_3307,N_3374);
nor U3404 (N_3404,N_3376,N_3321);
or U3405 (N_3405,N_3300,N_3397);
nor U3406 (N_3406,N_3346,N_3345);
nand U3407 (N_3407,N_3344,N_3361);
nor U3408 (N_3408,N_3351,N_3359);
nand U3409 (N_3409,N_3302,N_3303);
and U3410 (N_3410,N_3384,N_3387);
xor U3411 (N_3411,N_3339,N_3310);
and U3412 (N_3412,N_3356,N_3317);
or U3413 (N_3413,N_3375,N_3323);
xor U3414 (N_3414,N_3306,N_3362);
and U3415 (N_3415,N_3314,N_3324);
nand U3416 (N_3416,N_3367,N_3371);
nand U3417 (N_3417,N_3342,N_3395);
xor U3418 (N_3418,N_3372,N_3336);
and U3419 (N_3419,N_3364,N_3385);
and U3420 (N_3420,N_3322,N_3389);
xor U3421 (N_3421,N_3353,N_3329);
or U3422 (N_3422,N_3304,N_3341);
and U3423 (N_3423,N_3382,N_3366);
and U3424 (N_3424,N_3312,N_3338);
xnor U3425 (N_3425,N_3325,N_3348);
nor U3426 (N_3426,N_3370,N_3381);
nand U3427 (N_3427,N_3369,N_3358);
xnor U3428 (N_3428,N_3354,N_3305);
and U3429 (N_3429,N_3352,N_3363);
xor U3430 (N_3430,N_3343,N_3340);
nor U3431 (N_3431,N_3330,N_3337);
or U3432 (N_3432,N_3398,N_3328);
xnor U3433 (N_3433,N_3390,N_3327);
or U3434 (N_3434,N_3318,N_3388);
xor U3435 (N_3435,N_3386,N_3311);
and U3436 (N_3436,N_3355,N_3326);
and U3437 (N_3437,N_3357,N_3391);
nor U3438 (N_3438,N_3349,N_3393);
or U3439 (N_3439,N_3380,N_3394);
or U3440 (N_3440,N_3399,N_3334);
nand U3441 (N_3441,N_3373,N_3347);
nand U3442 (N_3442,N_3365,N_3309);
xor U3443 (N_3443,N_3333,N_3379);
nor U3444 (N_3444,N_3332,N_3360);
and U3445 (N_3445,N_3316,N_3308);
nand U3446 (N_3446,N_3383,N_3331);
nand U3447 (N_3447,N_3313,N_3315);
or U3448 (N_3448,N_3350,N_3319);
xor U3449 (N_3449,N_3396,N_3377);
nand U3450 (N_3450,N_3390,N_3393);
or U3451 (N_3451,N_3388,N_3391);
xnor U3452 (N_3452,N_3324,N_3362);
xnor U3453 (N_3453,N_3316,N_3376);
nand U3454 (N_3454,N_3327,N_3312);
and U3455 (N_3455,N_3384,N_3356);
xnor U3456 (N_3456,N_3349,N_3380);
xor U3457 (N_3457,N_3382,N_3353);
and U3458 (N_3458,N_3347,N_3344);
nor U3459 (N_3459,N_3309,N_3332);
and U3460 (N_3460,N_3352,N_3334);
nor U3461 (N_3461,N_3393,N_3359);
or U3462 (N_3462,N_3373,N_3385);
nand U3463 (N_3463,N_3388,N_3330);
nand U3464 (N_3464,N_3366,N_3388);
xnor U3465 (N_3465,N_3351,N_3375);
xor U3466 (N_3466,N_3378,N_3360);
nand U3467 (N_3467,N_3365,N_3311);
or U3468 (N_3468,N_3366,N_3362);
nand U3469 (N_3469,N_3336,N_3381);
nor U3470 (N_3470,N_3380,N_3375);
nand U3471 (N_3471,N_3337,N_3358);
nand U3472 (N_3472,N_3363,N_3327);
nand U3473 (N_3473,N_3364,N_3397);
and U3474 (N_3474,N_3305,N_3303);
or U3475 (N_3475,N_3316,N_3341);
nand U3476 (N_3476,N_3347,N_3329);
nor U3477 (N_3477,N_3335,N_3328);
or U3478 (N_3478,N_3352,N_3335);
xnor U3479 (N_3479,N_3368,N_3366);
or U3480 (N_3480,N_3343,N_3362);
nand U3481 (N_3481,N_3329,N_3396);
nand U3482 (N_3482,N_3367,N_3345);
and U3483 (N_3483,N_3310,N_3391);
and U3484 (N_3484,N_3326,N_3381);
and U3485 (N_3485,N_3351,N_3363);
xnor U3486 (N_3486,N_3313,N_3332);
nand U3487 (N_3487,N_3308,N_3351);
and U3488 (N_3488,N_3309,N_3349);
and U3489 (N_3489,N_3329,N_3318);
and U3490 (N_3490,N_3312,N_3317);
nor U3491 (N_3491,N_3300,N_3339);
nor U3492 (N_3492,N_3333,N_3332);
and U3493 (N_3493,N_3309,N_3388);
nand U3494 (N_3494,N_3309,N_3321);
nand U3495 (N_3495,N_3374,N_3310);
nand U3496 (N_3496,N_3395,N_3367);
or U3497 (N_3497,N_3388,N_3368);
nor U3498 (N_3498,N_3361,N_3339);
nand U3499 (N_3499,N_3366,N_3387);
xnor U3500 (N_3500,N_3478,N_3457);
xnor U3501 (N_3501,N_3487,N_3449);
and U3502 (N_3502,N_3465,N_3442);
nand U3503 (N_3503,N_3473,N_3472);
xor U3504 (N_3504,N_3480,N_3497);
and U3505 (N_3505,N_3440,N_3491);
xor U3506 (N_3506,N_3489,N_3410);
or U3507 (N_3507,N_3404,N_3488);
nor U3508 (N_3508,N_3405,N_3415);
nand U3509 (N_3509,N_3494,N_3427);
or U3510 (N_3510,N_3409,N_3458);
xnor U3511 (N_3511,N_3421,N_3466);
xnor U3512 (N_3512,N_3401,N_3485);
xor U3513 (N_3513,N_3419,N_3456);
or U3514 (N_3514,N_3486,N_3406);
nand U3515 (N_3515,N_3484,N_3423);
nor U3516 (N_3516,N_3495,N_3460);
nand U3517 (N_3517,N_3476,N_3499);
or U3518 (N_3518,N_3467,N_3453);
or U3519 (N_3519,N_3425,N_3413);
xor U3520 (N_3520,N_3437,N_3451);
or U3521 (N_3521,N_3429,N_3483);
and U3522 (N_3522,N_3412,N_3479);
nand U3523 (N_3523,N_3431,N_3403);
or U3524 (N_3524,N_3459,N_3475);
or U3525 (N_3525,N_3492,N_3493);
nand U3526 (N_3526,N_3496,N_3463);
nand U3527 (N_3527,N_3448,N_3481);
xor U3528 (N_3528,N_3420,N_3454);
and U3529 (N_3529,N_3470,N_3422);
nand U3530 (N_3530,N_3435,N_3468);
nand U3531 (N_3531,N_3434,N_3402);
and U3532 (N_3532,N_3436,N_3477);
or U3533 (N_3533,N_3464,N_3447);
and U3534 (N_3534,N_3439,N_3408);
and U3535 (N_3535,N_3445,N_3414);
nand U3536 (N_3536,N_3462,N_3407);
and U3537 (N_3537,N_3418,N_3444);
xnor U3538 (N_3538,N_3469,N_3424);
nand U3539 (N_3539,N_3416,N_3471);
xnor U3540 (N_3540,N_3482,N_3433);
and U3541 (N_3541,N_3438,N_3411);
nand U3542 (N_3542,N_3426,N_3443);
nand U3543 (N_3543,N_3400,N_3474);
or U3544 (N_3544,N_3432,N_3490);
and U3545 (N_3545,N_3446,N_3430);
nand U3546 (N_3546,N_3498,N_3450);
or U3547 (N_3547,N_3441,N_3455);
nor U3548 (N_3548,N_3452,N_3461);
and U3549 (N_3549,N_3428,N_3417);
or U3550 (N_3550,N_3401,N_3498);
and U3551 (N_3551,N_3415,N_3436);
and U3552 (N_3552,N_3470,N_3467);
and U3553 (N_3553,N_3415,N_3443);
nand U3554 (N_3554,N_3453,N_3465);
xor U3555 (N_3555,N_3446,N_3467);
and U3556 (N_3556,N_3432,N_3469);
or U3557 (N_3557,N_3412,N_3486);
nor U3558 (N_3558,N_3461,N_3499);
and U3559 (N_3559,N_3459,N_3439);
xor U3560 (N_3560,N_3422,N_3440);
nor U3561 (N_3561,N_3452,N_3438);
or U3562 (N_3562,N_3468,N_3410);
and U3563 (N_3563,N_3489,N_3413);
nand U3564 (N_3564,N_3401,N_3405);
xnor U3565 (N_3565,N_3404,N_3484);
and U3566 (N_3566,N_3436,N_3407);
or U3567 (N_3567,N_3405,N_3418);
nor U3568 (N_3568,N_3479,N_3445);
nand U3569 (N_3569,N_3409,N_3439);
and U3570 (N_3570,N_3486,N_3408);
xor U3571 (N_3571,N_3493,N_3444);
nand U3572 (N_3572,N_3412,N_3478);
nor U3573 (N_3573,N_3412,N_3495);
and U3574 (N_3574,N_3499,N_3418);
or U3575 (N_3575,N_3416,N_3406);
or U3576 (N_3576,N_3435,N_3472);
nor U3577 (N_3577,N_3424,N_3483);
nand U3578 (N_3578,N_3469,N_3460);
and U3579 (N_3579,N_3478,N_3488);
nor U3580 (N_3580,N_3474,N_3477);
and U3581 (N_3581,N_3467,N_3498);
nor U3582 (N_3582,N_3486,N_3429);
and U3583 (N_3583,N_3418,N_3457);
or U3584 (N_3584,N_3428,N_3487);
nand U3585 (N_3585,N_3427,N_3497);
nand U3586 (N_3586,N_3496,N_3466);
xnor U3587 (N_3587,N_3404,N_3412);
xnor U3588 (N_3588,N_3464,N_3489);
nor U3589 (N_3589,N_3458,N_3423);
or U3590 (N_3590,N_3415,N_3484);
and U3591 (N_3591,N_3426,N_3480);
nor U3592 (N_3592,N_3422,N_3496);
nor U3593 (N_3593,N_3476,N_3412);
xnor U3594 (N_3594,N_3422,N_3416);
nor U3595 (N_3595,N_3462,N_3412);
xnor U3596 (N_3596,N_3425,N_3481);
and U3597 (N_3597,N_3455,N_3491);
nor U3598 (N_3598,N_3438,N_3422);
or U3599 (N_3599,N_3404,N_3444);
nand U3600 (N_3600,N_3503,N_3521);
xor U3601 (N_3601,N_3590,N_3575);
nor U3602 (N_3602,N_3509,N_3545);
nand U3603 (N_3603,N_3592,N_3570);
or U3604 (N_3604,N_3579,N_3569);
and U3605 (N_3605,N_3567,N_3500);
xnor U3606 (N_3606,N_3586,N_3513);
and U3607 (N_3607,N_3522,N_3534);
xnor U3608 (N_3608,N_3502,N_3559);
and U3609 (N_3609,N_3561,N_3504);
or U3610 (N_3610,N_3568,N_3566);
or U3611 (N_3611,N_3539,N_3557);
xnor U3612 (N_3612,N_3529,N_3542);
nand U3613 (N_3613,N_3519,N_3541);
nand U3614 (N_3614,N_3576,N_3511);
xnor U3615 (N_3615,N_3597,N_3540);
and U3616 (N_3616,N_3558,N_3585);
and U3617 (N_3617,N_3520,N_3584);
and U3618 (N_3618,N_3582,N_3581);
or U3619 (N_3619,N_3524,N_3554);
nand U3620 (N_3620,N_3572,N_3543);
xor U3621 (N_3621,N_3587,N_3514);
or U3622 (N_3622,N_3505,N_3591);
nor U3623 (N_3623,N_3555,N_3574);
and U3624 (N_3624,N_3538,N_3595);
or U3625 (N_3625,N_3544,N_3596);
or U3626 (N_3626,N_3512,N_3523);
or U3627 (N_3627,N_3527,N_3507);
or U3628 (N_3628,N_3550,N_3530);
or U3629 (N_3629,N_3526,N_3578);
and U3630 (N_3630,N_3549,N_3535);
nor U3631 (N_3631,N_3556,N_3537);
and U3632 (N_3632,N_3598,N_3563);
or U3633 (N_3633,N_3546,N_3548);
xnor U3634 (N_3634,N_3564,N_3501);
nand U3635 (N_3635,N_3518,N_3560);
or U3636 (N_3636,N_3547,N_3533);
xnor U3637 (N_3637,N_3583,N_3589);
xnor U3638 (N_3638,N_3508,N_3516);
or U3639 (N_3639,N_3594,N_3536);
nor U3640 (N_3640,N_3573,N_3506);
nor U3641 (N_3641,N_3577,N_3580);
and U3642 (N_3642,N_3525,N_3510);
xnor U3643 (N_3643,N_3532,N_3599);
and U3644 (N_3644,N_3551,N_3588);
xnor U3645 (N_3645,N_3553,N_3517);
nand U3646 (N_3646,N_3593,N_3565);
and U3647 (N_3647,N_3562,N_3571);
nor U3648 (N_3648,N_3552,N_3515);
or U3649 (N_3649,N_3528,N_3531);
nand U3650 (N_3650,N_3524,N_3564);
and U3651 (N_3651,N_3559,N_3580);
or U3652 (N_3652,N_3542,N_3534);
xor U3653 (N_3653,N_3500,N_3541);
xor U3654 (N_3654,N_3552,N_3597);
or U3655 (N_3655,N_3551,N_3562);
or U3656 (N_3656,N_3573,N_3544);
nor U3657 (N_3657,N_3541,N_3510);
or U3658 (N_3658,N_3531,N_3522);
nor U3659 (N_3659,N_3564,N_3578);
or U3660 (N_3660,N_3554,N_3583);
xor U3661 (N_3661,N_3519,N_3543);
or U3662 (N_3662,N_3543,N_3551);
and U3663 (N_3663,N_3593,N_3589);
nand U3664 (N_3664,N_3505,N_3552);
xor U3665 (N_3665,N_3582,N_3593);
and U3666 (N_3666,N_3549,N_3546);
or U3667 (N_3667,N_3577,N_3583);
xor U3668 (N_3668,N_3585,N_3582);
and U3669 (N_3669,N_3561,N_3559);
and U3670 (N_3670,N_3553,N_3591);
nor U3671 (N_3671,N_3530,N_3581);
or U3672 (N_3672,N_3543,N_3529);
nand U3673 (N_3673,N_3548,N_3545);
xor U3674 (N_3674,N_3596,N_3594);
or U3675 (N_3675,N_3529,N_3586);
or U3676 (N_3676,N_3560,N_3540);
nand U3677 (N_3677,N_3524,N_3518);
or U3678 (N_3678,N_3566,N_3527);
or U3679 (N_3679,N_3536,N_3532);
nor U3680 (N_3680,N_3521,N_3546);
or U3681 (N_3681,N_3558,N_3563);
or U3682 (N_3682,N_3574,N_3579);
or U3683 (N_3683,N_3585,N_3505);
and U3684 (N_3684,N_3542,N_3597);
xnor U3685 (N_3685,N_3545,N_3536);
or U3686 (N_3686,N_3503,N_3545);
or U3687 (N_3687,N_3501,N_3531);
xor U3688 (N_3688,N_3580,N_3575);
xor U3689 (N_3689,N_3569,N_3503);
and U3690 (N_3690,N_3571,N_3533);
nand U3691 (N_3691,N_3590,N_3589);
or U3692 (N_3692,N_3537,N_3593);
nand U3693 (N_3693,N_3599,N_3525);
nor U3694 (N_3694,N_3575,N_3536);
xnor U3695 (N_3695,N_3557,N_3575);
and U3696 (N_3696,N_3504,N_3516);
nand U3697 (N_3697,N_3521,N_3583);
nor U3698 (N_3698,N_3567,N_3562);
nand U3699 (N_3699,N_3535,N_3558);
or U3700 (N_3700,N_3614,N_3601);
nand U3701 (N_3701,N_3615,N_3622);
and U3702 (N_3702,N_3645,N_3671);
xor U3703 (N_3703,N_3684,N_3696);
xor U3704 (N_3704,N_3647,N_3649);
nor U3705 (N_3705,N_3655,N_3692);
xor U3706 (N_3706,N_3687,N_3642);
nand U3707 (N_3707,N_3619,N_3634);
xnor U3708 (N_3708,N_3659,N_3676);
and U3709 (N_3709,N_3626,N_3613);
nor U3710 (N_3710,N_3653,N_3610);
nor U3711 (N_3711,N_3678,N_3636);
and U3712 (N_3712,N_3606,N_3677);
xnor U3713 (N_3713,N_3685,N_3637);
nor U3714 (N_3714,N_3621,N_3603);
nor U3715 (N_3715,N_3640,N_3608);
nor U3716 (N_3716,N_3666,N_3632);
xnor U3717 (N_3717,N_3664,N_3699);
and U3718 (N_3718,N_3646,N_3688);
or U3719 (N_3719,N_3697,N_3600);
nand U3720 (N_3720,N_3698,N_3695);
or U3721 (N_3721,N_3656,N_3611);
xnor U3722 (N_3722,N_3639,N_3650);
or U3723 (N_3723,N_3660,N_3612);
nor U3724 (N_3724,N_3690,N_3641);
xnor U3725 (N_3725,N_3651,N_3682);
or U3726 (N_3726,N_3617,N_3691);
nand U3727 (N_3727,N_3668,N_3672);
xnor U3728 (N_3728,N_3643,N_3654);
nor U3729 (N_3729,N_3635,N_3662);
xor U3730 (N_3730,N_3616,N_3675);
or U3731 (N_3731,N_3629,N_3674);
xnor U3732 (N_3732,N_3658,N_3638);
xor U3733 (N_3733,N_3657,N_3683);
xnor U3734 (N_3734,N_3631,N_3689);
xnor U3735 (N_3735,N_3667,N_3665);
and U3736 (N_3736,N_3680,N_3644);
nor U3737 (N_3737,N_3670,N_3628);
nor U3738 (N_3738,N_3624,N_3679);
nand U3739 (N_3739,N_3620,N_3669);
nor U3740 (N_3740,N_3681,N_3694);
or U3741 (N_3741,N_3627,N_3648);
xnor U3742 (N_3742,N_3661,N_3673);
nor U3743 (N_3743,N_3602,N_3663);
nand U3744 (N_3744,N_3633,N_3618);
nand U3745 (N_3745,N_3623,N_3630);
xnor U3746 (N_3746,N_3607,N_3686);
nor U3747 (N_3747,N_3604,N_3693);
nor U3748 (N_3748,N_3652,N_3605);
xnor U3749 (N_3749,N_3625,N_3609);
nor U3750 (N_3750,N_3666,N_3620);
and U3751 (N_3751,N_3649,N_3664);
nor U3752 (N_3752,N_3667,N_3652);
or U3753 (N_3753,N_3611,N_3642);
xor U3754 (N_3754,N_3641,N_3692);
nor U3755 (N_3755,N_3661,N_3624);
or U3756 (N_3756,N_3605,N_3641);
xnor U3757 (N_3757,N_3634,N_3665);
nand U3758 (N_3758,N_3629,N_3691);
or U3759 (N_3759,N_3689,N_3605);
or U3760 (N_3760,N_3630,N_3697);
nand U3761 (N_3761,N_3635,N_3675);
or U3762 (N_3762,N_3630,N_3671);
xnor U3763 (N_3763,N_3616,N_3689);
or U3764 (N_3764,N_3676,N_3688);
nand U3765 (N_3765,N_3660,N_3683);
and U3766 (N_3766,N_3648,N_3660);
and U3767 (N_3767,N_3617,N_3616);
xnor U3768 (N_3768,N_3673,N_3657);
xor U3769 (N_3769,N_3618,N_3681);
or U3770 (N_3770,N_3615,N_3684);
or U3771 (N_3771,N_3678,N_3653);
xor U3772 (N_3772,N_3621,N_3639);
xnor U3773 (N_3773,N_3699,N_3636);
nor U3774 (N_3774,N_3623,N_3608);
nand U3775 (N_3775,N_3690,N_3673);
nor U3776 (N_3776,N_3604,N_3638);
and U3777 (N_3777,N_3668,N_3695);
nand U3778 (N_3778,N_3605,N_3645);
xnor U3779 (N_3779,N_3625,N_3646);
xnor U3780 (N_3780,N_3627,N_3605);
xor U3781 (N_3781,N_3631,N_3668);
or U3782 (N_3782,N_3679,N_3696);
nand U3783 (N_3783,N_3686,N_3615);
or U3784 (N_3784,N_3650,N_3696);
nor U3785 (N_3785,N_3620,N_3678);
and U3786 (N_3786,N_3684,N_3613);
and U3787 (N_3787,N_3694,N_3636);
or U3788 (N_3788,N_3658,N_3624);
nor U3789 (N_3789,N_3660,N_3677);
xor U3790 (N_3790,N_3677,N_3618);
and U3791 (N_3791,N_3699,N_3606);
and U3792 (N_3792,N_3646,N_3632);
xor U3793 (N_3793,N_3681,N_3669);
or U3794 (N_3794,N_3600,N_3691);
and U3795 (N_3795,N_3603,N_3666);
and U3796 (N_3796,N_3650,N_3613);
nand U3797 (N_3797,N_3697,N_3675);
and U3798 (N_3798,N_3640,N_3663);
and U3799 (N_3799,N_3663,N_3693);
xor U3800 (N_3800,N_3736,N_3766);
nand U3801 (N_3801,N_3776,N_3788);
or U3802 (N_3802,N_3727,N_3738);
nand U3803 (N_3803,N_3743,N_3799);
and U3804 (N_3804,N_3791,N_3744);
nand U3805 (N_3805,N_3704,N_3707);
nand U3806 (N_3806,N_3781,N_3760);
or U3807 (N_3807,N_3767,N_3762);
or U3808 (N_3808,N_3732,N_3759);
xnor U3809 (N_3809,N_3726,N_3792);
and U3810 (N_3810,N_3752,N_3740);
xor U3811 (N_3811,N_3742,N_3722);
or U3812 (N_3812,N_3782,N_3772);
xor U3813 (N_3813,N_3710,N_3769);
nand U3814 (N_3814,N_3790,N_3797);
nor U3815 (N_3815,N_3783,N_3715);
xnor U3816 (N_3816,N_3739,N_3785);
or U3817 (N_3817,N_3729,N_3764);
xnor U3818 (N_3818,N_3702,N_3789);
nor U3819 (N_3819,N_3784,N_3737);
and U3820 (N_3820,N_3757,N_3765);
nor U3821 (N_3821,N_3712,N_3771);
nor U3822 (N_3822,N_3754,N_3773);
and U3823 (N_3823,N_3787,N_3711);
nor U3824 (N_3824,N_3793,N_3731);
nand U3825 (N_3825,N_3706,N_3700);
and U3826 (N_3826,N_3705,N_3794);
or U3827 (N_3827,N_3774,N_3786);
or U3828 (N_3828,N_3723,N_3708);
nor U3829 (N_3829,N_3770,N_3703);
nand U3830 (N_3830,N_3717,N_3749);
xor U3831 (N_3831,N_3756,N_3780);
or U3832 (N_3832,N_3758,N_3720);
xor U3833 (N_3833,N_3718,N_3746);
nand U3834 (N_3834,N_3778,N_3798);
xor U3835 (N_3835,N_3735,N_3777);
xor U3836 (N_3836,N_3747,N_3775);
xor U3837 (N_3837,N_3714,N_3728);
and U3838 (N_3838,N_3730,N_3751);
xor U3839 (N_3839,N_3753,N_3745);
nand U3840 (N_3840,N_3733,N_3721);
nor U3841 (N_3841,N_3748,N_3725);
nor U3842 (N_3842,N_3734,N_3761);
and U3843 (N_3843,N_3724,N_3768);
xor U3844 (N_3844,N_3750,N_3741);
or U3845 (N_3845,N_3709,N_3763);
nor U3846 (N_3846,N_3779,N_3701);
nand U3847 (N_3847,N_3713,N_3716);
and U3848 (N_3848,N_3795,N_3796);
nand U3849 (N_3849,N_3755,N_3719);
nor U3850 (N_3850,N_3714,N_3722);
nor U3851 (N_3851,N_3701,N_3791);
or U3852 (N_3852,N_3783,N_3795);
nor U3853 (N_3853,N_3703,N_3731);
nor U3854 (N_3854,N_3798,N_3728);
and U3855 (N_3855,N_3742,N_3797);
nor U3856 (N_3856,N_3760,N_3706);
and U3857 (N_3857,N_3713,N_3732);
nor U3858 (N_3858,N_3782,N_3750);
nor U3859 (N_3859,N_3706,N_3781);
nor U3860 (N_3860,N_3740,N_3771);
nor U3861 (N_3861,N_3775,N_3716);
xor U3862 (N_3862,N_3758,N_3793);
nand U3863 (N_3863,N_3777,N_3752);
nand U3864 (N_3864,N_3738,N_3705);
nand U3865 (N_3865,N_3719,N_3718);
nor U3866 (N_3866,N_3773,N_3788);
xnor U3867 (N_3867,N_3799,N_3763);
and U3868 (N_3868,N_3728,N_3723);
and U3869 (N_3869,N_3706,N_3707);
or U3870 (N_3870,N_3797,N_3709);
and U3871 (N_3871,N_3749,N_3781);
xor U3872 (N_3872,N_3723,N_3730);
nor U3873 (N_3873,N_3777,N_3762);
nand U3874 (N_3874,N_3719,N_3732);
and U3875 (N_3875,N_3719,N_3780);
nor U3876 (N_3876,N_3773,N_3736);
xor U3877 (N_3877,N_3713,N_3717);
xnor U3878 (N_3878,N_3799,N_3716);
nand U3879 (N_3879,N_3759,N_3727);
or U3880 (N_3880,N_3711,N_3755);
nor U3881 (N_3881,N_3765,N_3702);
nor U3882 (N_3882,N_3703,N_3717);
nor U3883 (N_3883,N_3716,N_3777);
or U3884 (N_3884,N_3725,N_3723);
or U3885 (N_3885,N_3706,N_3725);
xor U3886 (N_3886,N_3759,N_3706);
nand U3887 (N_3887,N_3715,N_3726);
nand U3888 (N_3888,N_3755,N_3772);
nor U3889 (N_3889,N_3722,N_3751);
nand U3890 (N_3890,N_3723,N_3735);
nor U3891 (N_3891,N_3751,N_3780);
nor U3892 (N_3892,N_3737,N_3742);
nand U3893 (N_3893,N_3757,N_3777);
nand U3894 (N_3894,N_3776,N_3764);
xor U3895 (N_3895,N_3774,N_3770);
or U3896 (N_3896,N_3716,N_3732);
or U3897 (N_3897,N_3765,N_3785);
nand U3898 (N_3898,N_3777,N_3737);
or U3899 (N_3899,N_3768,N_3782);
nor U3900 (N_3900,N_3839,N_3837);
xnor U3901 (N_3901,N_3823,N_3887);
and U3902 (N_3902,N_3878,N_3853);
or U3903 (N_3903,N_3804,N_3840);
or U3904 (N_3904,N_3884,N_3820);
xor U3905 (N_3905,N_3812,N_3838);
and U3906 (N_3906,N_3847,N_3825);
xor U3907 (N_3907,N_3886,N_3885);
nor U3908 (N_3908,N_3810,N_3828);
or U3909 (N_3909,N_3818,N_3861);
nor U3910 (N_3910,N_3831,N_3873);
nand U3911 (N_3911,N_3835,N_3892);
nor U3912 (N_3912,N_3832,N_3864);
nand U3913 (N_3913,N_3846,N_3800);
nand U3914 (N_3914,N_3852,N_3868);
nand U3915 (N_3915,N_3808,N_3859);
nand U3916 (N_3916,N_3856,N_3890);
nor U3917 (N_3917,N_3865,N_3894);
and U3918 (N_3918,N_3851,N_3869);
or U3919 (N_3919,N_3872,N_3821);
or U3920 (N_3920,N_3814,N_3858);
nor U3921 (N_3921,N_3888,N_3866);
xnor U3922 (N_3922,N_3898,N_3874);
nor U3923 (N_3923,N_3845,N_3819);
or U3924 (N_3924,N_3850,N_3809);
and U3925 (N_3925,N_3867,N_3803);
nor U3926 (N_3926,N_3870,N_3824);
nand U3927 (N_3927,N_3816,N_3876);
and U3928 (N_3928,N_3879,N_3813);
and U3929 (N_3929,N_3855,N_3801);
and U3930 (N_3930,N_3889,N_3834);
xor U3931 (N_3931,N_3871,N_3875);
nor U3932 (N_3932,N_3848,N_3815);
and U3933 (N_3933,N_3897,N_3807);
nand U3934 (N_3934,N_3822,N_3811);
nand U3935 (N_3935,N_3882,N_3844);
or U3936 (N_3936,N_3843,N_3817);
nor U3937 (N_3937,N_3880,N_3863);
nor U3938 (N_3938,N_3877,N_3806);
or U3939 (N_3939,N_3805,N_3896);
or U3940 (N_3940,N_3802,N_3895);
and U3941 (N_3941,N_3860,N_3836);
nand U3942 (N_3942,N_3830,N_3849);
xnor U3943 (N_3943,N_3857,N_3881);
nand U3944 (N_3944,N_3899,N_3891);
or U3945 (N_3945,N_3842,N_3829);
and U3946 (N_3946,N_3893,N_3862);
and U3947 (N_3947,N_3827,N_3883);
or U3948 (N_3948,N_3826,N_3841);
and U3949 (N_3949,N_3833,N_3854);
xor U3950 (N_3950,N_3814,N_3891);
or U3951 (N_3951,N_3818,N_3849);
nand U3952 (N_3952,N_3887,N_3874);
or U3953 (N_3953,N_3814,N_3881);
nand U3954 (N_3954,N_3886,N_3898);
nand U3955 (N_3955,N_3831,N_3805);
and U3956 (N_3956,N_3882,N_3828);
or U3957 (N_3957,N_3857,N_3843);
and U3958 (N_3958,N_3873,N_3854);
nor U3959 (N_3959,N_3832,N_3873);
xor U3960 (N_3960,N_3885,N_3832);
xnor U3961 (N_3961,N_3844,N_3848);
and U3962 (N_3962,N_3854,N_3879);
nand U3963 (N_3963,N_3817,N_3810);
and U3964 (N_3964,N_3820,N_3850);
or U3965 (N_3965,N_3816,N_3862);
nand U3966 (N_3966,N_3833,N_3815);
and U3967 (N_3967,N_3859,N_3849);
nor U3968 (N_3968,N_3827,N_3849);
and U3969 (N_3969,N_3834,N_3810);
nand U3970 (N_3970,N_3855,N_3817);
nor U3971 (N_3971,N_3824,N_3875);
xnor U3972 (N_3972,N_3837,N_3823);
and U3973 (N_3973,N_3812,N_3836);
nand U3974 (N_3974,N_3830,N_3811);
or U3975 (N_3975,N_3879,N_3844);
nand U3976 (N_3976,N_3828,N_3868);
and U3977 (N_3977,N_3814,N_3834);
nor U3978 (N_3978,N_3870,N_3812);
xnor U3979 (N_3979,N_3835,N_3815);
xnor U3980 (N_3980,N_3835,N_3822);
nand U3981 (N_3981,N_3832,N_3846);
nand U3982 (N_3982,N_3879,N_3831);
or U3983 (N_3983,N_3889,N_3853);
xor U3984 (N_3984,N_3844,N_3864);
nand U3985 (N_3985,N_3810,N_3869);
or U3986 (N_3986,N_3888,N_3876);
xor U3987 (N_3987,N_3819,N_3826);
or U3988 (N_3988,N_3848,N_3849);
xor U3989 (N_3989,N_3895,N_3801);
and U3990 (N_3990,N_3863,N_3868);
nor U3991 (N_3991,N_3852,N_3805);
nor U3992 (N_3992,N_3838,N_3800);
nand U3993 (N_3993,N_3824,N_3893);
and U3994 (N_3994,N_3865,N_3808);
nand U3995 (N_3995,N_3874,N_3877);
xor U3996 (N_3996,N_3896,N_3853);
nand U3997 (N_3997,N_3818,N_3808);
or U3998 (N_3998,N_3851,N_3821);
xor U3999 (N_3999,N_3829,N_3824);
and U4000 (N_4000,N_3929,N_3946);
or U4001 (N_4001,N_3952,N_3996);
and U4002 (N_4002,N_3992,N_3913);
nor U4003 (N_4003,N_3908,N_3937);
nand U4004 (N_4004,N_3991,N_3950);
and U4005 (N_4005,N_3940,N_3907);
nand U4006 (N_4006,N_3973,N_3949);
and U4007 (N_4007,N_3919,N_3927);
or U4008 (N_4008,N_3921,N_3944);
xnor U4009 (N_4009,N_3982,N_3928);
xnor U4010 (N_4010,N_3926,N_3904);
xor U4011 (N_4011,N_3900,N_3988);
or U4012 (N_4012,N_3964,N_3920);
or U4013 (N_4013,N_3972,N_3958);
nand U4014 (N_4014,N_3984,N_3995);
nand U4015 (N_4015,N_3971,N_3934);
nor U4016 (N_4016,N_3918,N_3911);
nor U4017 (N_4017,N_3922,N_3987);
xnor U4018 (N_4018,N_3909,N_3974);
nand U4019 (N_4019,N_3917,N_3943);
xnor U4020 (N_4020,N_3967,N_3914);
or U4021 (N_4021,N_3925,N_3941);
nor U4022 (N_4022,N_3989,N_3936);
nand U4023 (N_4023,N_3986,N_3965);
nor U4024 (N_4024,N_3968,N_3997);
nand U4025 (N_4025,N_3977,N_3933);
nand U4026 (N_4026,N_3956,N_3978);
and U4027 (N_4027,N_3970,N_3985);
xnor U4028 (N_4028,N_3905,N_3955);
or U4029 (N_4029,N_3999,N_3980);
or U4030 (N_4030,N_3923,N_3932);
nor U4031 (N_4031,N_3912,N_3959);
nand U4032 (N_4032,N_3942,N_3993);
xor U4033 (N_4033,N_3963,N_3961);
nor U4034 (N_4034,N_3906,N_3990);
xnor U4035 (N_4035,N_3969,N_3903);
nand U4036 (N_4036,N_3998,N_3957);
and U4037 (N_4037,N_3938,N_3945);
nor U4038 (N_4038,N_3915,N_3947);
xnor U4039 (N_4039,N_3975,N_3939);
nor U4040 (N_4040,N_3948,N_3976);
or U4041 (N_4041,N_3960,N_3979);
nand U4042 (N_4042,N_3951,N_3902);
and U4043 (N_4043,N_3924,N_3966);
nor U4044 (N_4044,N_3983,N_3935);
and U4045 (N_4045,N_3916,N_3953);
nand U4046 (N_4046,N_3962,N_3931);
and U4047 (N_4047,N_3901,N_3981);
nand U4048 (N_4048,N_3910,N_3930);
nor U4049 (N_4049,N_3994,N_3954);
and U4050 (N_4050,N_3991,N_3939);
or U4051 (N_4051,N_3985,N_3940);
nand U4052 (N_4052,N_3983,N_3919);
xor U4053 (N_4053,N_3980,N_3944);
xor U4054 (N_4054,N_3906,N_3907);
nand U4055 (N_4055,N_3936,N_3906);
xnor U4056 (N_4056,N_3935,N_3982);
and U4057 (N_4057,N_3964,N_3907);
or U4058 (N_4058,N_3944,N_3962);
and U4059 (N_4059,N_3927,N_3911);
nand U4060 (N_4060,N_3915,N_3901);
or U4061 (N_4061,N_3939,N_3914);
nor U4062 (N_4062,N_3956,N_3935);
nor U4063 (N_4063,N_3901,N_3920);
xor U4064 (N_4064,N_3993,N_3988);
nand U4065 (N_4065,N_3915,N_3946);
xnor U4066 (N_4066,N_3918,N_3944);
nand U4067 (N_4067,N_3973,N_3971);
xnor U4068 (N_4068,N_3956,N_3936);
and U4069 (N_4069,N_3999,N_3955);
and U4070 (N_4070,N_3938,N_3937);
nand U4071 (N_4071,N_3938,N_3921);
nor U4072 (N_4072,N_3943,N_3936);
nand U4073 (N_4073,N_3996,N_3908);
xor U4074 (N_4074,N_3980,N_3970);
xor U4075 (N_4075,N_3925,N_3942);
and U4076 (N_4076,N_3964,N_3971);
nand U4077 (N_4077,N_3914,N_3913);
nand U4078 (N_4078,N_3945,N_3921);
nor U4079 (N_4079,N_3901,N_3924);
nand U4080 (N_4080,N_3989,N_3991);
and U4081 (N_4081,N_3947,N_3936);
or U4082 (N_4082,N_3998,N_3980);
xnor U4083 (N_4083,N_3919,N_3962);
xor U4084 (N_4084,N_3964,N_3973);
or U4085 (N_4085,N_3910,N_3949);
or U4086 (N_4086,N_3954,N_3972);
nor U4087 (N_4087,N_3981,N_3924);
nand U4088 (N_4088,N_3994,N_3965);
or U4089 (N_4089,N_3986,N_3961);
nor U4090 (N_4090,N_3916,N_3946);
xnor U4091 (N_4091,N_3924,N_3951);
xnor U4092 (N_4092,N_3922,N_3930);
xnor U4093 (N_4093,N_3998,N_3920);
xor U4094 (N_4094,N_3944,N_3910);
xor U4095 (N_4095,N_3926,N_3929);
or U4096 (N_4096,N_3982,N_3922);
nand U4097 (N_4097,N_3988,N_3965);
nor U4098 (N_4098,N_3902,N_3900);
nand U4099 (N_4099,N_3980,N_3946);
nor U4100 (N_4100,N_4061,N_4056);
or U4101 (N_4101,N_4060,N_4016);
xor U4102 (N_4102,N_4088,N_4027);
xnor U4103 (N_4103,N_4033,N_4058);
xnor U4104 (N_4104,N_4077,N_4003);
and U4105 (N_4105,N_4073,N_4086);
xor U4106 (N_4106,N_4085,N_4024);
and U4107 (N_4107,N_4072,N_4097);
and U4108 (N_4108,N_4047,N_4000);
xnor U4109 (N_4109,N_4042,N_4028);
nand U4110 (N_4110,N_4032,N_4075);
or U4111 (N_4111,N_4049,N_4011);
nor U4112 (N_4112,N_4019,N_4092);
or U4113 (N_4113,N_4029,N_4002);
nand U4114 (N_4114,N_4017,N_4043);
or U4115 (N_4115,N_4021,N_4052);
or U4116 (N_4116,N_4083,N_4026);
or U4117 (N_4117,N_4091,N_4015);
and U4118 (N_4118,N_4065,N_4053);
xnor U4119 (N_4119,N_4045,N_4054);
and U4120 (N_4120,N_4035,N_4009);
nand U4121 (N_4121,N_4025,N_4068);
xor U4122 (N_4122,N_4023,N_4006);
or U4123 (N_4123,N_4051,N_4041);
or U4124 (N_4124,N_4071,N_4008);
or U4125 (N_4125,N_4096,N_4076);
nand U4126 (N_4126,N_4046,N_4036);
and U4127 (N_4127,N_4022,N_4067);
nor U4128 (N_4128,N_4087,N_4099);
nand U4129 (N_4129,N_4037,N_4090);
nor U4130 (N_4130,N_4004,N_4062);
nand U4131 (N_4131,N_4095,N_4034);
nand U4132 (N_4132,N_4078,N_4066);
or U4133 (N_4133,N_4082,N_4079);
and U4134 (N_4134,N_4069,N_4044);
xnor U4135 (N_4135,N_4081,N_4093);
or U4136 (N_4136,N_4031,N_4055);
nor U4137 (N_4137,N_4030,N_4098);
xor U4138 (N_4138,N_4074,N_4059);
or U4139 (N_4139,N_4057,N_4001);
or U4140 (N_4140,N_4040,N_4070);
and U4141 (N_4141,N_4064,N_4013);
nand U4142 (N_4142,N_4094,N_4063);
and U4143 (N_4143,N_4014,N_4039);
nor U4144 (N_4144,N_4084,N_4050);
and U4145 (N_4145,N_4080,N_4048);
xnor U4146 (N_4146,N_4089,N_4038);
nand U4147 (N_4147,N_4010,N_4005);
or U4148 (N_4148,N_4007,N_4020);
nand U4149 (N_4149,N_4012,N_4018);
nand U4150 (N_4150,N_4058,N_4090);
xor U4151 (N_4151,N_4041,N_4043);
xnor U4152 (N_4152,N_4083,N_4063);
nand U4153 (N_4153,N_4098,N_4019);
nand U4154 (N_4154,N_4092,N_4056);
xor U4155 (N_4155,N_4060,N_4074);
nand U4156 (N_4156,N_4063,N_4020);
and U4157 (N_4157,N_4013,N_4010);
or U4158 (N_4158,N_4019,N_4071);
and U4159 (N_4159,N_4059,N_4037);
nand U4160 (N_4160,N_4086,N_4042);
nand U4161 (N_4161,N_4012,N_4059);
or U4162 (N_4162,N_4053,N_4039);
nor U4163 (N_4163,N_4068,N_4061);
nand U4164 (N_4164,N_4081,N_4055);
and U4165 (N_4165,N_4011,N_4074);
xnor U4166 (N_4166,N_4041,N_4076);
nand U4167 (N_4167,N_4037,N_4098);
nor U4168 (N_4168,N_4093,N_4063);
xnor U4169 (N_4169,N_4020,N_4009);
nor U4170 (N_4170,N_4094,N_4026);
or U4171 (N_4171,N_4074,N_4099);
or U4172 (N_4172,N_4070,N_4015);
or U4173 (N_4173,N_4005,N_4095);
nand U4174 (N_4174,N_4082,N_4013);
nor U4175 (N_4175,N_4050,N_4047);
and U4176 (N_4176,N_4010,N_4089);
and U4177 (N_4177,N_4042,N_4056);
nand U4178 (N_4178,N_4017,N_4021);
xor U4179 (N_4179,N_4059,N_4094);
nor U4180 (N_4180,N_4094,N_4055);
nor U4181 (N_4181,N_4036,N_4082);
or U4182 (N_4182,N_4085,N_4064);
and U4183 (N_4183,N_4008,N_4027);
nor U4184 (N_4184,N_4091,N_4011);
and U4185 (N_4185,N_4003,N_4011);
nor U4186 (N_4186,N_4006,N_4015);
or U4187 (N_4187,N_4077,N_4021);
nand U4188 (N_4188,N_4070,N_4061);
or U4189 (N_4189,N_4079,N_4066);
nor U4190 (N_4190,N_4052,N_4031);
xor U4191 (N_4191,N_4064,N_4033);
and U4192 (N_4192,N_4075,N_4028);
or U4193 (N_4193,N_4060,N_4043);
or U4194 (N_4194,N_4062,N_4061);
or U4195 (N_4195,N_4039,N_4060);
xnor U4196 (N_4196,N_4068,N_4085);
nor U4197 (N_4197,N_4070,N_4051);
or U4198 (N_4198,N_4072,N_4019);
nand U4199 (N_4199,N_4060,N_4067);
or U4200 (N_4200,N_4113,N_4156);
xor U4201 (N_4201,N_4116,N_4163);
or U4202 (N_4202,N_4111,N_4138);
xnor U4203 (N_4203,N_4188,N_4140);
nand U4204 (N_4204,N_4150,N_4133);
or U4205 (N_4205,N_4160,N_4165);
xnor U4206 (N_4206,N_4182,N_4159);
xor U4207 (N_4207,N_4142,N_4139);
xor U4208 (N_4208,N_4124,N_4167);
or U4209 (N_4209,N_4171,N_4101);
or U4210 (N_4210,N_4131,N_4105);
or U4211 (N_4211,N_4197,N_4191);
or U4212 (N_4212,N_4157,N_4164);
xnor U4213 (N_4213,N_4178,N_4189);
nor U4214 (N_4214,N_4155,N_4172);
xor U4215 (N_4215,N_4198,N_4106);
or U4216 (N_4216,N_4103,N_4100);
xnor U4217 (N_4217,N_4153,N_4122);
xnor U4218 (N_4218,N_4173,N_4104);
nand U4219 (N_4219,N_4115,N_4126);
xor U4220 (N_4220,N_4174,N_4166);
and U4221 (N_4221,N_4127,N_4125);
xnor U4222 (N_4222,N_4162,N_4137);
xor U4223 (N_4223,N_4107,N_4154);
nand U4224 (N_4224,N_4194,N_4168);
xor U4225 (N_4225,N_4192,N_4141);
and U4226 (N_4226,N_4144,N_4169);
nand U4227 (N_4227,N_4187,N_4143);
xnor U4228 (N_4228,N_4110,N_4185);
xnor U4229 (N_4229,N_4193,N_4190);
nor U4230 (N_4230,N_4136,N_4176);
nand U4231 (N_4231,N_4180,N_4161);
and U4232 (N_4232,N_4119,N_4108);
nand U4233 (N_4233,N_4152,N_4151);
or U4234 (N_4234,N_4120,N_4118);
nand U4235 (N_4235,N_4184,N_4132);
or U4236 (N_4236,N_4117,N_4121);
or U4237 (N_4237,N_4112,N_4145);
nand U4238 (N_4238,N_4149,N_4186);
nor U4239 (N_4239,N_4146,N_4128);
or U4240 (N_4240,N_4179,N_4129);
and U4241 (N_4241,N_4177,N_4109);
or U4242 (N_4242,N_4147,N_4134);
nor U4243 (N_4243,N_4158,N_4135);
or U4244 (N_4244,N_4196,N_4175);
nand U4245 (N_4245,N_4148,N_4199);
or U4246 (N_4246,N_4130,N_4195);
xor U4247 (N_4247,N_4181,N_4183);
nor U4248 (N_4248,N_4170,N_4102);
or U4249 (N_4249,N_4114,N_4123);
nand U4250 (N_4250,N_4137,N_4187);
xnor U4251 (N_4251,N_4130,N_4134);
nor U4252 (N_4252,N_4182,N_4180);
xnor U4253 (N_4253,N_4113,N_4103);
or U4254 (N_4254,N_4160,N_4147);
nor U4255 (N_4255,N_4125,N_4139);
or U4256 (N_4256,N_4148,N_4130);
nand U4257 (N_4257,N_4192,N_4179);
and U4258 (N_4258,N_4145,N_4118);
xor U4259 (N_4259,N_4156,N_4158);
and U4260 (N_4260,N_4180,N_4160);
nand U4261 (N_4261,N_4126,N_4136);
and U4262 (N_4262,N_4125,N_4133);
xor U4263 (N_4263,N_4181,N_4152);
xnor U4264 (N_4264,N_4105,N_4119);
or U4265 (N_4265,N_4193,N_4137);
nor U4266 (N_4266,N_4173,N_4126);
nor U4267 (N_4267,N_4178,N_4150);
or U4268 (N_4268,N_4158,N_4186);
or U4269 (N_4269,N_4170,N_4100);
xor U4270 (N_4270,N_4116,N_4108);
or U4271 (N_4271,N_4137,N_4183);
xnor U4272 (N_4272,N_4195,N_4122);
nand U4273 (N_4273,N_4189,N_4197);
and U4274 (N_4274,N_4131,N_4139);
nand U4275 (N_4275,N_4119,N_4169);
and U4276 (N_4276,N_4197,N_4140);
and U4277 (N_4277,N_4119,N_4195);
or U4278 (N_4278,N_4145,N_4162);
or U4279 (N_4279,N_4186,N_4110);
nand U4280 (N_4280,N_4144,N_4110);
nand U4281 (N_4281,N_4176,N_4110);
and U4282 (N_4282,N_4107,N_4175);
nor U4283 (N_4283,N_4130,N_4122);
xor U4284 (N_4284,N_4146,N_4186);
nor U4285 (N_4285,N_4164,N_4172);
nor U4286 (N_4286,N_4131,N_4159);
nor U4287 (N_4287,N_4157,N_4123);
or U4288 (N_4288,N_4133,N_4148);
and U4289 (N_4289,N_4194,N_4124);
nand U4290 (N_4290,N_4167,N_4198);
nor U4291 (N_4291,N_4116,N_4118);
or U4292 (N_4292,N_4141,N_4197);
xor U4293 (N_4293,N_4182,N_4102);
nand U4294 (N_4294,N_4171,N_4152);
nor U4295 (N_4295,N_4125,N_4164);
and U4296 (N_4296,N_4141,N_4198);
or U4297 (N_4297,N_4120,N_4185);
xor U4298 (N_4298,N_4151,N_4178);
xor U4299 (N_4299,N_4118,N_4143);
or U4300 (N_4300,N_4208,N_4255);
nand U4301 (N_4301,N_4254,N_4266);
xnor U4302 (N_4302,N_4220,N_4200);
xor U4303 (N_4303,N_4232,N_4219);
or U4304 (N_4304,N_4221,N_4214);
xor U4305 (N_4305,N_4263,N_4217);
nor U4306 (N_4306,N_4216,N_4239);
and U4307 (N_4307,N_4241,N_4279);
nor U4308 (N_4308,N_4284,N_4223);
nand U4309 (N_4309,N_4298,N_4209);
and U4310 (N_4310,N_4294,N_4240);
nand U4311 (N_4311,N_4233,N_4229);
nand U4312 (N_4312,N_4280,N_4268);
nor U4313 (N_4313,N_4274,N_4215);
xor U4314 (N_4314,N_4291,N_4258);
nor U4315 (N_4315,N_4297,N_4287);
nor U4316 (N_4316,N_4234,N_4289);
xnor U4317 (N_4317,N_4210,N_4276);
or U4318 (N_4318,N_4295,N_4231);
and U4319 (N_4319,N_4265,N_4222);
or U4320 (N_4320,N_4253,N_4299);
or U4321 (N_4321,N_4246,N_4251);
nand U4322 (N_4322,N_4278,N_4247);
and U4323 (N_4323,N_4260,N_4269);
and U4324 (N_4324,N_4249,N_4248);
xor U4325 (N_4325,N_4267,N_4252);
nand U4326 (N_4326,N_4238,N_4245);
or U4327 (N_4327,N_4250,N_4224);
xnor U4328 (N_4328,N_4257,N_4275);
nor U4329 (N_4329,N_4259,N_4270);
xnor U4330 (N_4330,N_4264,N_4226);
or U4331 (N_4331,N_4218,N_4286);
xor U4332 (N_4332,N_4242,N_4293);
nor U4333 (N_4333,N_4227,N_4206);
nand U4334 (N_4334,N_4235,N_4262);
nor U4335 (N_4335,N_4285,N_4230);
nand U4336 (N_4336,N_4281,N_4272);
xor U4337 (N_4337,N_4292,N_4256);
nand U4338 (N_4338,N_4243,N_4271);
and U4339 (N_4339,N_4211,N_4282);
xnor U4340 (N_4340,N_4204,N_4296);
or U4341 (N_4341,N_4288,N_4261);
nor U4342 (N_4342,N_4228,N_4237);
nand U4343 (N_4343,N_4225,N_4207);
and U4344 (N_4344,N_4290,N_4203);
or U4345 (N_4345,N_4205,N_4202);
xnor U4346 (N_4346,N_4283,N_4236);
and U4347 (N_4347,N_4277,N_4273);
or U4348 (N_4348,N_4213,N_4201);
nand U4349 (N_4349,N_4244,N_4212);
and U4350 (N_4350,N_4282,N_4262);
nor U4351 (N_4351,N_4232,N_4217);
xor U4352 (N_4352,N_4250,N_4229);
nor U4353 (N_4353,N_4260,N_4263);
nand U4354 (N_4354,N_4240,N_4232);
nor U4355 (N_4355,N_4298,N_4212);
and U4356 (N_4356,N_4260,N_4258);
nor U4357 (N_4357,N_4263,N_4232);
or U4358 (N_4358,N_4220,N_4240);
and U4359 (N_4359,N_4212,N_4285);
or U4360 (N_4360,N_4210,N_4240);
xor U4361 (N_4361,N_4255,N_4271);
and U4362 (N_4362,N_4271,N_4241);
nand U4363 (N_4363,N_4234,N_4295);
or U4364 (N_4364,N_4263,N_4243);
nand U4365 (N_4365,N_4224,N_4242);
and U4366 (N_4366,N_4210,N_4242);
nor U4367 (N_4367,N_4214,N_4255);
or U4368 (N_4368,N_4292,N_4209);
xor U4369 (N_4369,N_4204,N_4208);
nand U4370 (N_4370,N_4281,N_4249);
nor U4371 (N_4371,N_4214,N_4259);
and U4372 (N_4372,N_4268,N_4245);
and U4373 (N_4373,N_4292,N_4220);
nor U4374 (N_4374,N_4299,N_4244);
xnor U4375 (N_4375,N_4268,N_4273);
and U4376 (N_4376,N_4296,N_4209);
and U4377 (N_4377,N_4222,N_4286);
xnor U4378 (N_4378,N_4268,N_4200);
nor U4379 (N_4379,N_4200,N_4213);
or U4380 (N_4380,N_4214,N_4204);
nand U4381 (N_4381,N_4237,N_4232);
and U4382 (N_4382,N_4266,N_4210);
and U4383 (N_4383,N_4260,N_4299);
nand U4384 (N_4384,N_4248,N_4298);
nand U4385 (N_4385,N_4272,N_4280);
and U4386 (N_4386,N_4262,N_4213);
nand U4387 (N_4387,N_4249,N_4215);
xor U4388 (N_4388,N_4220,N_4238);
nand U4389 (N_4389,N_4295,N_4220);
nor U4390 (N_4390,N_4259,N_4211);
and U4391 (N_4391,N_4282,N_4298);
nor U4392 (N_4392,N_4201,N_4280);
and U4393 (N_4393,N_4259,N_4227);
and U4394 (N_4394,N_4219,N_4249);
or U4395 (N_4395,N_4292,N_4240);
nand U4396 (N_4396,N_4228,N_4207);
or U4397 (N_4397,N_4278,N_4273);
nor U4398 (N_4398,N_4226,N_4201);
nor U4399 (N_4399,N_4201,N_4263);
and U4400 (N_4400,N_4339,N_4369);
nand U4401 (N_4401,N_4309,N_4336);
nand U4402 (N_4402,N_4341,N_4385);
xnor U4403 (N_4403,N_4329,N_4313);
nand U4404 (N_4404,N_4316,N_4320);
and U4405 (N_4405,N_4330,N_4315);
nor U4406 (N_4406,N_4378,N_4311);
nor U4407 (N_4407,N_4344,N_4383);
or U4408 (N_4408,N_4331,N_4363);
xor U4409 (N_4409,N_4353,N_4332);
nor U4410 (N_4410,N_4349,N_4308);
xor U4411 (N_4411,N_4372,N_4347);
nor U4412 (N_4412,N_4328,N_4312);
nand U4413 (N_4413,N_4374,N_4322);
nand U4414 (N_4414,N_4395,N_4396);
nand U4415 (N_4415,N_4394,N_4376);
and U4416 (N_4416,N_4381,N_4305);
nor U4417 (N_4417,N_4398,N_4327);
xor U4418 (N_4418,N_4338,N_4364);
xnor U4419 (N_4419,N_4384,N_4355);
and U4420 (N_4420,N_4388,N_4342);
xnor U4421 (N_4421,N_4324,N_4345);
nand U4422 (N_4422,N_4368,N_4362);
nand U4423 (N_4423,N_4340,N_4386);
nand U4424 (N_4424,N_4300,N_4371);
xnor U4425 (N_4425,N_4357,N_4318);
nor U4426 (N_4426,N_4354,N_4301);
nor U4427 (N_4427,N_4333,N_4399);
or U4428 (N_4428,N_4302,N_4377);
nand U4429 (N_4429,N_4310,N_4325);
nor U4430 (N_4430,N_4379,N_4307);
nor U4431 (N_4431,N_4350,N_4387);
nand U4432 (N_4432,N_4382,N_4389);
and U4433 (N_4433,N_4346,N_4392);
nand U4434 (N_4434,N_4317,N_4359);
nor U4435 (N_4435,N_4314,N_4380);
or U4436 (N_4436,N_4303,N_4360);
xor U4437 (N_4437,N_4358,N_4306);
xnor U4438 (N_4438,N_4390,N_4326);
xor U4439 (N_4439,N_4352,N_4356);
and U4440 (N_4440,N_4304,N_4391);
xnor U4441 (N_4441,N_4393,N_4375);
nor U4442 (N_4442,N_4323,N_4321);
and U4443 (N_4443,N_4365,N_4367);
or U4444 (N_4444,N_4319,N_4343);
and U4445 (N_4445,N_4366,N_4351);
xor U4446 (N_4446,N_4361,N_4373);
and U4447 (N_4447,N_4334,N_4370);
nor U4448 (N_4448,N_4397,N_4348);
and U4449 (N_4449,N_4335,N_4337);
xor U4450 (N_4450,N_4302,N_4308);
xor U4451 (N_4451,N_4365,N_4370);
or U4452 (N_4452,N_4329,N_4385);
or U4453 (N_4453,N_4307,N_4321);
and U4454 (N_4454,N_4390,N_4368);
and U4455 (N_4455,N_4304,N_4370);
or U4456 (N_4456,N_4353,N_4339);
nand U4457 (N_4457,N_4376,N_4309);
or U4458 (N_4458,N_4334,N_4302);
nand U4459 (N_4459,N_4341,N_4314);
or U4460 (N_4460,N_4364,N_4312);
or U4461 (N_4461,N_4346,N_4319);
nor U4462 (N_4462,N_4345,N_4394);
or U4463 (N_4463,N_4328,N_4393);
nand U4464 (N_4464,N_4386,N_4362);
or U4465 (N_4465,N_4319,N_4311);
nor U4466 (N_4466,N_4377,N_4336);
xnor U4467 (N_4467,N_4328,N_4372);
xnor U4468 (N_4468,N_4349,N_4314);
nand U4469 (N_4469,N_4357,N_4337);
and U4470 (N_4470,N_4380,N_4347);
nand U4471 (N_4471,N_4392,N_4319);
and U4472 (N_4472,N_4394,N_4304);
nor U4473 (N_4473,N_4307,N_4323);
nor U4474 (N_4474,N_4302,N_4365);
or U4475 (N_4475,N_4378,N_4313);
xor U4476 (N_4476,N_4338,N_4349);
or U4477 (N_4477,N_4394,N_4368);
nand U4478 (N_4478,N_4373,N_4367);
nor U4479 (N_4479,N_4320,N_4394);
and U4480 (N_4480,N_4300,N_4394);
nand U4481 (N_4481,N_4395,N_4372);
xnor U4482 (N_4482,N_4385,N_4349);
nand U4483 (N_4483,N_4372,N_4390);
xnor U4484 (N_4484,N_4364,N_4390);
and U4485 (N_4485,N_4396,N_4389);
nor U4486 (N_4486,N_4365,N_4311);
or U4487 (N_4487,N_4357,N_4322);
or U4488 (N_4488,N_4329,N_4380);
nand U4489 (N_4489,N_4395,N_4373);
nand U4490 (N_4490,N_4337,N_4323);
and U4491 (N_4491,N_4336,N_4333);
nor U4492 (N_4492,N_4347,N_4338);
xnor U4493 (N_4493,N_4309,N_4346);
and U4494 (N_4494,N_4306,N_4310);
xor U4495 (N_4495,N_4350,N_4327);
xor U4496 (N_4496,N_4317,N_4337);
xor U4497 (N_4497,N_4312,N_4398);
and U4498 (N_4498,N_4356,N_4376);
xnor U4499 (N_4499,N_4343,N_4302);
or U4500 (N_4500,N_4492,N_4448);
nand U4501 (N_4501,N_4421,N_4409);
nor U4502 (N_4502,N_4472,N_4445);
or U4503 (N_4503,N_4452,N_4474);
xnor U4504 (N_4504,N_4483,N_4429);
and U4505 (N_4505,N_4426,N_4420);
xor U4506 (N_4506,N_4488,N_4415);
or U4507 (N_4507,N_4471,N_4428);
and U4508 (N_4508,N_4437,N_4411);
xor U4509 (N_4509,N_4425,N_4436);
xor U4510 (N_4510,N_4458,N_4493);
or U4511 (N_4511,N_4439,N_4406);
nor U4512 (N_4512,N_4449,N_4480);
nand U4513 (N_4513,N_4435,N_4431);
xnor U4514 (N_4514,N_4497,N_4401);
nor U4515 (N_4515,N_4487,N_4499);
nand U4516 (N_4516,N_4418,N_4491);
or U4517 (N_4517,N_4404,N_4402);
nor U4518 (N_4518,N_4476,N_4454);
and U4519 (N_4519,N_4423,N_4486);
and U4520 (N_4520,N_4478,N_4419);
nor U4521 (N_4521,N_4457,N_4447);
or U4522 (N_4522,N_4417,N_4412);
nor U4523 (N_4523,N_4468,N_4496);
or U4524 (N_4524,N_4408,N_4432);
nor U4525 (N_4525,N_4450,N_4430);
or U4526 (N_4526,N_4455,N_4462);
and U4527 (N_4527,N_4407,N_4442);
and U4528 (N_4528,N_4466,N_4498);
or U4529 (N_4529,N_4461,N_4405);
and U4530 (N_4530,N_4460,N_4410);
nand U4531 (N_4531,N_4427,N_4459);
or U4532 (N_4532,N_4414,N_4469);
xnor U4533 (N_4533,N_4453,N_4464);
or U4534 (N_4534,N_4441,N_4470);
and U4535 (N_4535,N_4400,N_4463);
and U4536 (N_4536,N_4403,N_4440);
nor U4537 (N_4537,N_4494,N_4465);
nand U4538 (N_4538,N_4484,N_4475);
or U4539 (N_4539,N_4446,N_4481);
or U4540 (N_4540,N_4467,N_4451);
xor U4541 (N_4541,N_4434,N_4490);
xor U4542 (N_4542,N_4443,N_4485);
nand U4543 (N_4543,N_4473,N_4456);
or U4544 (N_4544,N_4495,N_4433);
or U4545 (N_4545,N_4479,N_4422);
xnor U4546 (N_4546,N_4424,N_4482);
or U4547 (N_4547,N_4477,N_4416);
or U4548 (N_4548,N_4438,N_4413);
and U4549 (N_4549,N_4444,N_4489);
nor U4550 (N_4550,N_4492,N_4440);
or U4551 (N_4551,N_4462,N_4410);
xnor U4552 (N_4552,N_4415,N_4442);
or U4553 (N_4553,N_4446,N_4453);
or U4554 (N_4554,N_4400,N_4454);
or U4555 (N_4555,N_4490,N_4488);
or U4556 (N_4556,N_4419,N_4488);
and U4557 (N_4557,N_4492,N_4449);
or U4558 (N_4558,N_4476,N_4425);
xnor U4559 (N_4559,N_4420,N_4468);
nand U4560 (N_4560,N_4487,N_4429);
or U4561 (N_4561,N_4426,N_4464);
or U4562 (N_4562,N_4497,N_4460);
or U4563 (N_4563,N_4481,N_4468);
nand U4564 (N_4564,N_4445,N_4478);
and U4565 (N_4565,N_4411,N_4407);
xor U4566 (N_4566,N_4449,N_4488);
xnor U4567 (N_4567,N_4426,N_4454);
and U4568 (N_4568,N_4470,N_4424);
nand U4569 (N_4569,N_4418,N_4419);
or U4570 (N_4570,N_4458,N_4407);
and U4571 (N_4571,N_4485,N_4494);
and U4572 (N_4572,N_4458,N_4495);
and U4573 (N_4573,N_4431,N_4485);
and U4574 (N_4574,N_4449,N_4481);
nand U4575 (N_4575,N_4443,N_4419);
and U4576 (N_4576,N_4447,N_4414);
or U4577 (N_4577,N_4494,N_4417);
xor U4578 (N_4578,N_4417,N_4449);
xnor U4579 (N_4579,N_4476,N_4410);
xnor U4580 (N_4580,N_4424,N_4443);
xnor U4581 (N_4581,N_4411,N_4440);
xnor U4582 (N_4582,N_4485,N_4472);
or U4583 (N_4583,N_4475,N_4470);
nand U4584 (N_4584,N_4425,N_4440);
or U4585 (N_4585,N_4421,N_4420);
and U4586 (N_4586,N_4470,N_4497);
xnor U4587 (N_4587,N_4450,N_4473);
or U4588 (N_4588,N_4467,N_4447);
and U4589 (N_4589,N_4499,N_4463);
and U4590 (N_4590,N_4465,N_4445);
or U4591 (N_4591,N_4455,N_4497);
xnor U4592 (N_4592,N_4457,N_4490);
and U4593 (N_4593,N_4490,N_4428);
xor U4594 (N_4594,N_4460,N_4455);
and U4595 (N_4595,N_4421,N_4491);
and U4596 (N_4596,N_4444,N_4427);
xor U4597 (N_4597,N_4465,N_4483);
and U4598 (N_4598,N_4487,N_4484);
or U4599 (N_4599,N_4458,N_4421);
or U4600 (N_4600,N_4522,N_4598);
and U4601 (N_4601,N_4590,N_4523);
nor U4602 (N_4602,N_4554,N_4504);
nand U4603 (N_4603,N_4579,N_4545);
and U4604 (N_4604,N_4509,N_4515);
nand U4605 (N_4605,N_4533,N_4596);
xor U4606 (N_4606,N_4539,N_4501);
or U4607 (N_4607,N_4593,N_4546);
nand U4608 (N_4608,N_4537,N_4525);
or U4609 (N_4609,N_4551,N_4578);
or U4610 (N_4610,N_4585,N_4550);
or U4611 (N_4611,N_4548,N_4524);
nand U4612 (N_4612,N_4594,N_4583);
or U4613 (N_4613,N_4587,N_4544);
or U4614 (N_4614,N_4572,N_4507);
xnor U4615 (N_4615,N_4516,N_4529);
and U4616 (N_4616,N_4518,N_4592);
and U4617 (N_4617,N_4506,N_4560);
nand U4618 (N_4618,N_4595,N_4556);
xor U4619 (N_4619,N_4588,N_4532);
nor U4620 (N_4620,N_4512,N_4564);
nor U4621 (N_4621,N_4530,N_4520);
or U4622 (N_4622,N_4575,N_4535);
xnor U4623 (N_4623,N_4511,N_4569);
nor U4624 (N_4624,N_4568,N_4527);
nor U4625 (N_4625,N_4528,N_4508);
nor U4626 (N_4626,N_4536,N_4517);
and U4627 (N_4627,N_4514,N_4555);
nand U4628 (N_4628,N_4599,N_4543);
xor U4629 (N_4629,N_4589,N_4573);
or U4630 (N_4630,N_4552,N_4577);
and U4631 (N_4631,N_4553,N_4584);
nor U4632 (N_4632,N_4591,N_4566);
nor U4633 (N_4633,N_4576,N_4559);
nand U4634 (N_4634,N_4538,N_4563);
xnor U4635 (N_4635,N_4510,N_4505);
and U4636 (N_4636,N_4541,N_4574);
or U4637 (N_4637,N_4503,N_4557);
nor U4638 (N_4638,N_4570,N_4526);
nor U4639 (N_4639,N_4502,N_4597);
or U4640 (N_4640,N_4571,N_4581);
and U4641 (N_4641,N_4567,N_4582);
xor U4642 (N_4642,N_4521,N_4513);
nand U4643 (N_4643,N_4540,N_4547);
nor U4644 (N_4644,N_4558,N_4565);
or U4645 (N_4645,N_4586,N_4542);
nor U4646 (N_4646,N_4562,N_4519);
nor U4647 (N_4647,N_4534,N_4580);
nand U4648 (N_4648,N_4531,N_4549);
and U4649 (N_4649,N_4500,N_4561);
and U4650 (N_4650,N_4512,N_4505);
and U4651 (N_4651,N_4588,N_4581);
xnor U4652 (N_4652,N_4554,N_4521);
nand U4653 (N_4653,N_4598,N_4529);
nand U4654 (N_4654,N_4504,N_4501);
xnor U4655 (N_4655,N_4558,N_4578);
xnor U4656 (N_4656,N_4544,N_4548);
or U4657 (N_4657,N_4507,N_4532);
xnor U4658 (N_4658,N_4530,N_4534);
nor U4659 (N_4659,N_4551,N_4598);
nand U4660 (N_4660,N_4565,N_4508);
nor U4661 (N_4661,N_4597,N_4588);
or U4662 (N_4662,N_4539,N_4551);
xnor U4663 (N_4663,N_4580,N_4562);
or U4664 (N_4664,N_4511,N_4513);
xor U4665 (N_4665,N_4557,N_4548);
and U4666 (N_4666,N_4503,N_4536);
or U4667 (N_4667,N_4548,N_4540);
and U4668 (N_4668,N_4577,N_4548);
and U4669 (N_4669,N_4506,N_4517);
xor U4670 (N_4670,N_4596,N_4586);
nor U4671 (N_4671,N_4595,N_4534);
and U4672 (N_4672,N_4525,N_4555);
nor U4673 (N_4673,N_4567,N_4504);
xor U4674 (N_4674,N_4592,N_4552);
nor U4675 (N_4675,N_4500,N_4573);
or U4676 (N_4676,N_4527,N_4567);
nor U4677 (N_4677,N_4597,N_4567);
xor U4678 (N_4678,N_4567,N_4543);
nand U4679 (N_4679,N_4562,N_4553);
or U4680 (N_4680,N_4566,N_4509);
nand U4681 (N_4681,N_4517,N_4568);
nor U4682 (N_4682,N_4598,N_4581);
nand U4683 (N_4683,N_4543,N_4582);
and U4684 (N_4684,N_4590,N_4517);
and U4685 (N_4685,N_4509,N_4582);
xnor U4686 (N_4686,N_4592,N_4523);
xnor U4687 (N_4687,N_4531,N_4581);
or U4688 (N_4688,N_4580,N_4528);
nand U4689 (N_4689,N_4572,N_4584);
nor U4690 (N_4690,N_4515,N_4533);
or U4691 (N_4691,N_4509,N_4579);
nor U4692 (N_4692,N_4539,N_4522);
and U4693 (N_4693,N_4516,N_4506);
and U4694 (N_4694,N_4586,N_4583);
or U4695 (N_4695,N_4504,N_4523);
and U4696 (N_4696,N_4584,N_4575);
or U4697 (N_4697,N_4512,N_4561);
and U4698 (N_4698,N_4581,N_4510);
and U4699 (N_4699,N_4502,N_4585);
nor U4700 (N_4700,N_4647,N_4660);
xnor U4701 (N_4701,N_4661,N_4646);
or U4702 (N_4702,N_4695,N_4685);
xor U4703 (N_4703,N_4652,N_4689);
xnor U4704 (N_4704,N_4635,N_4672);
nor U4705 (N_4705,N_4617,N_4669);
nor U4706 (N_4706,N_4633,N_4693);
nand U4707 (N_4707,N_4602,N_4632);
nand U4708 (N_4708,N_4600,N_4682);
or U4709 (N_4709,N_4607,N_4696);
nor U4710 (N_4710,N_4653,N_4666);
and U4711 (N_4711,N_4681,N_4609);
nand U4712 (N_4712,N_4658,N_4676);
xor U4713 (N_4713,N_4615,N_4637);
nor U4714 (N_4714,N_4625,N_4662);
xor U4715 (N_4715,N_4616,N_4640);
nor U4716 (N_4716,N_4678,N_4697);
xnor U4717 (N_4717,N_4606,N_4684);
or U4718 (N_4718,N_4611,N_4673);
nor U4719 (N_4719,N_4654,N_4649);
and U4720 (N_4720,N_4601,N_4644);
xnor U4721 (N_4721,N_4664,N_4604);
nand U4722 (N_4722,N_4671,N_4688);
nor U4723 (N_4723,N_4623,N_4641);
or U4724 (N_4724,N_4659,N_4613);
nand U4725 (N_4725,N_4603,N_4618);
nor U4726 (N_4726,N_4624,N_4614);
nor U4727 (N_4727,N_4663,N_4619);
xor U4728 (N_4728,N_4698,N_4639);
xnor U4729 (N_4729,N_4656,N_4627);
and U4730 (N_4730,N_4638,N_4621);
nand U4731 (N_4731,N_4629,N_4612);
xor U4732 (N_4732,N_4683,N_4605);
xor U4733 (N_4733,N_4634,N_4657);
and U4734 (N_4734,N_4648,N_4626);
nor U4735 (N_4735,N_4691,N_4665);
nor U4736 (N_4736,N_4642,N_4674);
xnor U4737 (N_4737,N_4677,N_4631);
and U4738 (N_4738,N_4670,N_4643);
and U4739 (N_4739,N_4699,N_4622);
xnor U4740 (N_4740,N_4668,N_4680);
xor U4741 (N_4741,N_4655,N_4608);
xor U4742 (N_4742,N_4636,N_4628);
nand U4743 (N_4743,N_4667,N_4651);
xor U4744 (N_4744,N_4650,N_4675);
xor U4745 (N_4745,N_4679,N_4692);
xnor U4746 (N_4746,N_4690,N_4620);
or U4747 (N_4747,N_4610,N_4686);
and U4748 (N_4748,N_4645,N_4687);
nand U4749 (N_4749,N_4630,N_4694);
nand U4750 (N_4750,N_4636,N_4654);
nor U4751 (N_4751,N_4655,N_4629);
xnor U4752 (N_4752,N_4658,N_4678);
or U4753 (N_4753,N_4600,N_4671);
and U4754 (N_4754,N_4629,N_4639);
nor U4755 (N_4755,N_4664,N_4614);
and U4756 (N_4756,N_4683,N_4674);
nor U4757 (N_4757,N_4629,N_4602);
xor U4758 (N_4758,N_4668,N_4698);
nand U4759 (N_4759,N_4633,N_4612);
nor U4760 (N_4760,N_4612,N_4658);
or U4761 (N_4761,N_4650,N_4615);
nor U4762 (N_4762,N_4613,N_4629);
nor U4763 (N_4763,N_4600,N_4642);
nand U4764 (N_4764,N_4699,N_4680);
or U4765 (N_4765,N_4656,N_4650);
and U4766 (N_4766,N_4649,N_4679);
nor U4767 (N_4767,N_4625,N_4655);
or U4768 (N_4768,N_4633,N_4675);
or U4769 (N_4769,N_4636,N_4655);
and U4770 (N_4770,N_4608,N_4640);
and U4771 (N_4771,N_4670,N_4610);
or U4772 (N_4772,N_4680,N_4650);
or U4773 (N_4773,N_4663,N_4681);
and U4774 (N_4774,N_4617,N_4647);
nor U4775 (N_4775,N_4626,N_4664);
nand U4776 (N_4776,N_4607,N_4676);
xor U4777 (N_4777,N_4652,N_4697);
or U4778 (N_4778,N_4699,N_4629);
and U4779 (N_4779,N_4641,N_4627);
nand U4780 (N_4780,N_4619,N_4631);
nand U4781 (N_4781,N_4636,N_4626);
nand U4782 (N_4782,N_4676,N_4605);
xor U4783 (N_4783,N_4638,N_4606);
or U4784 (N_4784,N_4617,N_4633);
nand U4785 (N_4785,N_4646,N_4622);
and U4786 (N_4786,N_4688,N_4638);
and U4787 (N_4787,N_4632,N_4616);
or U4788 (N_4788,N_4691,N_4650);
nor U4789 (N_4789,N_4674,N_4677);
nand U4790 (N_4790,N_4623,N_4664);
or U4791 (N_4791,N_4634,N_4690);
or U4792 (N_4792,N_4673,N_4667);
nand U4793 (N_4793,N_4644,N_4693);
nand U4794 (N_4794,N_4638,N_4637);
xnor U4795 (N_4795,N_4629,N_4620);
nand U4796 (N_4796,N_4678,N_4634);
or U4797 (N_4797,N_4603,N_4664);
nor U4798 (N_4798,N_4613,N_4626);
nor U4799 (N_4799,N_4678,N_4609);
and U4800 (N_4800,N_4745,N_4732);
nand U4801 (N_4801,N_4739,N_4767);
xor U4802 (N_4802,N_4753,N_4709);
or U4803 (N_4803,N_4774,N_4791);
nor U4804 (N_4804,N_4746,N_4733);
or U4805 (N_4805,N_4797,N_4758);
xor U4806 (N_4806,N_4705,N_4723);
nand U4807 (N_4807,N_4725,N_4764);
and U4808 (N_4808,N_4757,N_4773);
nor U4809 (N_4809,N_4783,N_4728);
nor U4810 (N_4810,N_4780,N_4787);
xnor U4811 (N_4811,N_4776,N_4765);
nor U4812 (N_4812,N_4798,N_4768);
or U4813 (N_4813,N_4740,N_4715);
and U4814 (N_4814,N_4789,N_4735);
xor U4815 (N_4815,N_4754,N_4730);
nand U4816 (N_4816,N_4755,N_4790);
or U4817 (N_4817,N_4786,N_4788);
or U4818 (N_4818,N_4763,N_4748);
and U4819 (N_4819,N_4731,N_4793);
and U4820 (N_4820,N_4741,N_4703);
nor U4821 (N_4821,N_4749,N_4770);
xor U4822 (N_4822,N_4714,N_4782);
nand U4823 (N_4823,N_4704,N_4772);
nand U4824 (N_4824,N_4759,N_4794);
and U4825 (N_4825,N_4760,N_4707);
or U4826 (N_4826,N_4799,N_4779);
nor U4827 (N_4827,N_4750,N_4752);
or U4828 (N_4828,N_4766,N_4751);
and U4829 (N_4829,N_4747,N_4712);
nor U4830 (N_4830,N_4784,N_4706);
xor U4831 (N_4831,N_4775,N_4734);
nand U4832 (N_4832,N_4771,N_4700);
nand U4833 (N_4833,N_4769,N_4701);
or U4834 (N_4834,N_4719,N_4724);
or U4835 (N_4835,N_4796,N_4729);
and U4836 (N_4836,N_4708,N_4762);
xnor U4837 (N_4837,N_4702,N_4718);
or U4838 (N_4838,N_4710,N_4722);
or U4839 (N_4839,N_4743,N_4713);
nor U4840 (N_4840,N_4717,N_4727);
or U4841 (N_4841,N_4737,N_4726);
or U4842 (N_4842,N_4777,N_4761);
nor U4843 (N_4843,N_4711,N_4736);
xnor U4844 (N_4844,N_4781,N_4792);
and U4845 (N_4845,N_4778,N_4721);
or U4846 (N_4846,N_4795,N_4756);
nand U4847 (N_4847,N_4716,N_4720);
xor U4848 (N_4848,N_4744,N_4738);
nand U4849 (N_4849,N_4785,N_4742);
xor U4850 (N_4850,N_4738,N_4731);
nor U4851 (N_4851,N_4782,N_4707);
nor U4852 (N_4852,N_4778,N_4759);
xor U4853 (N_4853,N_4788,N_4746);
xnor U4854 (N_4854,N_4707,N_4719);
nor U4855 (N_4855,N_4756,N_4746);
xor U4856 (N_4856,N_4755,N_4711);
and U4857 (N_4857,N_4707,N_4781);
nor U4858 (N_4858,N_4731,N_4790);
xor U4859 (N_4859,N_4766,N_4763);
or U4860 (N_4860,N_4781,N_4778);
xor U4861 (N_4861,N_4720,N_4724);
nor U4862 (N_4862,N_4776,N_4714);
nor U4863 (N_4863,N_4734,N_4760);
nand U4864 (N_4864,N_4789,N_4774);
or U4865 (N_4865,N_4766,N_4781);
and U4866 (N_4866,N_4756,N_4702);
nor U4867 (N_4867,N_4726,N_4787);
nand U4868 (N_4868,N_4709,N_4734);
and U4869 (N_4869,N_4761,N_4737);
xor U4870 (N_4870,N_4721,N_4755);
nand U4871 (N_4871,N_4738,N_4704);
or U4872 (N_4872,N_4794,N_4713);
or U4873 (N_4873,N_4726,N_4793);
nand U4874 (N_4874,N_4718,N_4700);
nand U4875 (N_4875,N_4769,N_4778);
and U4876 (N_4876,N_4703,N_4764);
xnor U4877 (N_4877,N_4777,N_4738);
nand U4878 (N_4878,N_4795,N_4752);
xor U4879 (N_4879,N_4728,N_4770);
or U4880 (N_4880,N_4776,N_4710);
and U4881 (N_4881,N_4753,N_4726);
nand U4882 (N_4882,N_4797,N_4713);
xnor U4883 (N_4883,N_4799,N_4798);
nand U4884 (N_4884,N_4754,N_4792);
nand U4885 (N_4885,N_4756,N_4743);
xor U4886 (N_4886,N_4791,N_4763);
or U4887 (N_4887,N_4775,N_4731);
or U4888 (N_4888,N_4739,N_4706);
or U4889 (N_4889,N_4770,N_4726);
and U4890 (N_4890,N_4718,N_4778);
and U4891 (N_4891,N_4733,N_4727);
and U4892 (N_4892,N_4718,N_4750);
nand U4893 (N_4893,N_4771,N_4750);
and U4894 (N_4894,N_4706,N_4779);
and U4895 (N_4895,N_4735,N_4722);
nor U4896 (N_4896,N_4787,N_4788);
xor U4897 (N_4897,N_4795,N_4721);
xnor U4898 (N_4898,N_4779,N_4728);
xnor U4899 (N_4899,N_4707,N_4780);
nor U4900 (N_4900,N_4886,N_4892);
nand U4901 (N_4901,N_4868,N_4816);
and U4902 (N_4902,N_4802,N_4844);
xnor U4903 (N_4903,N_4846,N_4888);
nor U4904 (N_4904,N_4869,N_4831);
and U4905 (N_4905,N_4884,N_4890);
xnor U4906 (N_4906,N_4847,N_4861);
xnor U4907 (N_4907,N_4879,N_4842);
or U4908 (N_4908,N_4824,N_4829);
or U4909 (N_4909,N_4838,N_4867);
nor U4910 (N_4910,N_4817,N_4894);
nor U4911 (N_4911,N_4833,N_4828);
and U4912 (N_4912,N_4864,N_4836);
or U4913 (N_4913,N_4819,N_4812);
nor U4914 (N_4914,N_4880,N_4889);
xor U4915 (N_4915,N_4810,N_4878);
xnor U4916 (N_4916,N_4805,N_4808);
nand U4917 (N_4917,N_4804,N_4809);
nor U4918 (N_4918,N_4863,N_4811);
xor U4919 (N_4919,N_4870,N_4893);
nor U4920 (N_4920,N_4815,N_4848);
or U4921 (N_4921,N_4840,N_4849);
xnor U4922 (N_4922,N_4800,N_4837);
nand U4923 (N_4923,N_4898,N_4881);
and U4924 (N_4924,N_4841,N_4851);
nand U4925 (N_4925,N_4859,N_4803);
nor U4926 (N_4926,N_4806,N_4856);
nor U4927 (N_4927,N_4875,N_4818);
and U4928 (N_4928,N_4855,N_4822);
or U4929 (N_4929,N_4896,N_4865);
nor U4930 (N_4930,N_4862,N_4895);
or U4931 (N_4931,N_4839,N_4823);
or U4932 (N_4932,N_4877,N_4882);
nor U4933 (N_4933,N_4852,N_4897);
nor U4934 (N_4934,N_4891,N_4845);
nor U4935 (N_4935,N_4820,N_4827);
and U4936 (N_4936,N_4813,N_4854);
or U4937 (N_4937,N_4872,N_4874);
nor U4938 (N_4938,N_4834,N_4899);
nor U4939 (N_4939,N_4858,N_4843);
or U4940 (N_4940,N_4807,N_4830);
nand U4941 (N_4941,N_4826,N_4821);
or U4942 (N_4942,N_4885,N_4825);
nand U4943 (N_4943,N_4857,N_4883);
or U4944 (N_4944,N_4887,N_4801);
xnor U4945 (N_4945,N_4835,N_4814);
nand U4946 (N_4946,N_4860,N_4876);
or U4947 (N_4947,N_4853,N_4832);
xor U4948 (N_4948,N_4871,N_4866);
nand U4949 (N_4949,N_4873,N_4850);
xor U4950 (N_4950,N_4806,N_4838);
nand U4951 (N_4951,N_4881,N_4855);
xnor U4952 (N_4952,N_4875,N_4889);
nand U4953 (N_4953,N_4803,N_4833);
and U4954 (N_4954,N_4896,N_4844);
nand U4955 (N_4955,N_4851,N_4829);
and U4956 (N_4956,N_4838,N_4845);
and U4957 (N_4957,N_4876,N_4843);
nor U4958 (N_4958,N_4813,N_4836);
or U4959 (N_4959,N_4889,N_4801);
nand U4960 (N_4960,N_4803,N_4881);
and U4961 (N_4961,N_4887,N_4859);
and U4962 (N_4962,N_4884,N_4895);
xor U4963 (N_4963,N_4869,N_4849);
or U4964 (N_4964,N_4872,N_4886);
and U4965 (N_4965,N_4832,N_4881);
or U4966 (N_4966,N_4883,N_4870);
or U4967 (N_4967,N_4802,N_4813);
xor U4968 (N_4968,N_4846,N_4836);
nand U4969 (N_4969,N_4841,N_4882);
or U4970 (N_4970,N_4881,N_4857);
and U4971 (N_4971,N_4867,N_4851);
or U4972 (N_4972,N_4836,N_4820);
and U4973 (N_4973,N_4867,N_4819);
nand U4974 (N_4974,N_4817,N_4809);
nor U4975 (N_4975,N_4862,N_4834);
nor U4976 (N_4976,N_4850,N_4822);
xnor U4977 (N_4977,N_4816,N_4815);
nand U4978 (N_4978,N_4824,N_4804);
and U4979 (N_4979,N_4815,N_4870);
or U4980 (N_4980,N_4835,N_4869);
or U4981 (N_4981,N_4891,N_4894);
or U4982 (N_4982,N_4816,N_4823);
xor U4983 (N_4983,N_4857,N_4844);
xor U4984 (N_4984,N_4867,N_4804);
and U4985 (N_4985,N_4883,N_4823);
or U4986 (N_4986,N_4828,N_4868);
xor U4987 (N_4987,N_4851,N_4881);
nand U4988 (N_4988,N_4807,N_4887);
and U4989 (N_4989,N_4802,N_4889);
xor U4990 (N_4990,N_4872,N_4825);
xnor U4991 (N_4991,N_4862,N_4824);
and U4992 (N_4992,N_4882,N_4811);
nand U4993 (N_4993,N_4825,N_4831);
and U4994 (N_4994,N_4876,N_4889);
and U4995 (N_4995,N_4891,N_4806);
nor U4996 (N_4996,N_4878,N_4884);
xnor U4997 (N_4997,N_4804,N_4869);
nand U4998 (N_4998,N_4850,N_4899);
nand U4999 (N_4999,N_4865,N_4860);
or UO_0 (O_0,N_4929,N_4956);
nand UO_1 (O_1,N_4930,N_4991);
xnor UO_2 (O_2,N_4920,N_4962);
or UO_3 (O_3,N_4985,N_4901);
xnor UO_4 (O_4,N_4937,N_4910);
nor UO_5 (O_5,N_4940,N_4931);
xor UO_6 (O_6,N_4996,N_4928);
and UO_7 (O_7,N_4993,N_4968);
xnor UO_8 (O_8,N_4925,N_4947);
xor UO_9 (O_9,N_4951,N_4994);
xnor UO_10 (O_10,N_4907,N_4953);
and UO_11 (O_11,N_4960,N_4981);
xnor UO_12 (O_12,N_4913,N_4946);
nor UO_13 (O_13,N_4914,N_4954);
nand UO_14 (O_14,N_4926,N_4978);
nor UO_15 (O_15,N_4967,N_4927);
xor UO_16 (O_16,N_4963,N_4952);
nor UO_17 (O_17,N_4966,N_4992);
or UO_18 (O_18,N_4906,N_4948);
nand UO_19 (O_19,N_4902,N_4934);
and UO_20 (O_20,N_4904,N_4916);
xnor UO_21 (O_21,N_4945,N_4932);
nand UO_22 (O_22,N_4998,N_4908);
and UO_23 (O_23,N_4923,N_4957);
or UO_24 (O_24,N_4989,N_4961);
and UO_25 (O_25,N_4964,N_4941);
xor UO_26 (O_26,N_4976,N_4944);
xnor UO_27 (O_27,N_4972,N_4917);
nor UO_28 (O_28,N_4900,N_4988);
or UO_29 (O_29,N_4958,N_4979);
and UO_30 (O_30,N_4915,N_4975);
or UO_31 (O_31,N_4942,N_4903);
nand UO_32 (O_32,N_4933,N_4936);
xor UO_33 (O_33,N_4924,N_4939);
and UO_34 (O_34,N_4922,N_4921);
nand UO_35 (O_35,N_4909,N_4943);
nand UO_36 (O_36,N_4984,N_4970);
and UO_37 (O_37,N_4986,N_4997);
or UO_38 (O_38,N_4949,N_4982);
nand UO_39 (O_39,N_4990,N_4911);
nand UO_40 (O_40,N_4980,N_4999);
nor UO_41 (O_41,N_4973,N_4918);
or UO_42 (O_42,N_4974,N_4938);
nand UO_43 (O_43,N_4955,N_4971);
or UO_44 (O_44,N_4919,N_4935);
and UO_45 (O_45,N_4995,N_4987);
nand UO_46 (O_46,N_4905,N_4965);
or UO_47 (O_47,N_4959,N_4950);
nor UO_48 (O_48,N_4977,N_4912);
nor UO_49 (O_49,N_4969,N_4983);
nand UO_50 (O_50,N_4988,N_4981);
and UO_51 (O_51,N_4999,N_4969);
nand UO_52 (O_52,N_4965,N_4948);
or UO_53 (O_53,N_4949,N_4968);
nor UO_54 (O_54,N_4966,N_4927);
and UO_55 (O_55,N_4912,N_4998);
nor UO_56 (O_56,N_4939,N_4954);
or UO_57 (O_57,N_4995,N_4962);
nor UO_58 (O_58,N_4982,N_4905);
nand UO_59 (O_59,N_4901,N_4908);
xor UO_60 (O_60,N_4947,N_4990);
or UO_61 (O_61,N_4985,N_4937);
and UO_62 (O_62,N_4916,N_4953);
nand UO_63 (O_63,N_4920,N_4929);
and UO_64 (O_64,N_4981,N_4941);
and UO_65 (O_65,N_4901,N_4935);
xor UO_66 (O_66,N_4927,N_4971);
and UO_67 (O_67,N_4932,N_4943);
nor UO_68 (O_68,N_4952,N_4940);
nand UO_69 (O_69,N_4981,N_4909);
nand UO_70 (O_70,N_4962,N_4942);
nand UO_71 (O_71,N_4962,N_4986);
or UO_72 (O_72,N_4928,N_4916);
nand UO_73 (O_73,N_4972,N_4977);
and UO_74 (O_74,N_4945,N_4970);
xnor UO_75 (O_75,N_4937,N_4909);
and UO_76 (O_76,N_4935,N_4925);
nor UO_77 (O_77,N_4979,N_4904);
xor UO_78 (O_78,N_4905,N_4987);
nand UO_79 (O_79,N_4935,N_4963);
xnor UO_80 (O_80,N_4987,N_4999);
nor UO_81 (O_81,N_4919,N_4962);
xor UO_82 (O_82,N_4983,N_4910);
xor UO_83 (O_83,N_4982,N_4934);
xor UO_84 (O_84,N_4911,N_4950);
and UO_85 (O_85,N_4925,N_4945);
nand UO_86 (O_86,N_4990,N_4915);
and UO_87 (O_87,N_4944,N_4995);
and UO_88 (O_88,N_4915,N_4927);
nand UO_89 (O_89,N_4922,N_4900);
nand UO_90 (O_90,N_4959,N_4962);
nand UO_91 (O_91,N_4929,N_4963);
nor UO_92 (O_92,N_4910,N_4915);
nand UO_93 (O_93,N_4948,N_4989);
or UO_94 (O_94,N_4964,N_4948);
or UO_95 (O_95,N_4952,N_4982);
xor UO_96 (O_96,N_4972,N_4915);
nand UO_97 (O_97,N_4930,N_4923);
xor UO_98 (O_98,N_4949,N_4902);
and UO_99 (O_99,N_4915,N_4912);
nor UO_100 (O_100,N_4981,N_4976);
or UO_101 (O_101,N_4967,N_4925);
and UO_102 (O_102,N_4907,N_4937);
xnor UO_103 (O_103,N_4909,N_4970);
or UO_104 (O_104,N_4942,N_4998);
nor UO_105 (O_105,N_4942,N_4946);
nor UO_106 (O_106,N_4996,N_4917);
nand UO_107 (O_107,N_4987,N_4933);
or UO_108 (O_108,N_4997,N_4934);
and UO_109 (O_109,N_4984,N_4914);
nor UO_110 (O_110,N_4933,N_4917);
or UO_111 (O_111,N_4990,N_4910);
or UO_112 (O_112,N_4952,N_4906);
nor UO_113 (O_113,N_4910,N_4981);
nor UO_114 (O_114,N_4911,N_4988);
or UO_115 (O_115,N_4978,N_4982);
and UO_116 (O_116,N_4913,N_4982);
nor UO_117 (O_117,N_4993,N_4920);
nand UO_118 (O_118,N_4966,N_4977);
or UO_119 (O_119,N_4995,N_4963);
or UO_120 (O_120,N_4950,N_4970);
xor UO_121 (O_121,N_4969,N_4939);
nand UO_122 (O_122,N_4933,N_4982);
nand UO_123 (O_123,N_4962,N_4937);
and UO_124 (O_124,N_4963,N_4949);
nand UO_125 (O_125,N_4952,N_4923);
and UO_126 (O_126,N_4926,N_4928);
and UO_127 (O_127,N_4988,N_4973);
xnor UO_128 (O_128,N_4915,N_4932);
or UO_129 (O_129,N_4908,N_4966);
nand UO_130 (O_130,N_4949,N_4907);
nand UO_131 (O_131,N_4927,N_4976);
nand UO_132 (O_132,N_4945,N_4923);
and UO_133 (O_133,N_4969,N_4991);
nor UO_134 (O_134,N_4952,N_4946);
nor UO_135 (O_135,N_4990,N_4977);
nor UO_136 (O_136,N_4908,N_4915);
nor UO_137 (O_137,N_4967,N_4988);
and UO_138 (O_138,N_4942,N_4980);
and UO_139 (O_139,N_4947,N_4999);
nand UO_140 (O_140,N_4928,N_4934);
and UO_141 (O_141,N_4918,N_4969);
or UO_142 (O_142,N_4909,N_4925);
xor UO_143 (O_143,N_4911,N_4918);
nand UO_144 (O_144,N_4918,N_4950);
and UO_145 (O_145,N_4990,N_4972);
nand UO_146 (O_146,N_4991,N_4937);
or UO_147 (O_147,N_4971,N_4936);
or UO_148 (O_148,N_4973,N_4920);
nor UO_149 (O_149,N_4910,N_4906);
nand UO_150 (O_150,N_4952,N_4987);
or UO_151 (O_151,N_4995,N_4946);
nor UO_152 (O_152,N_4985,N_4986);
nand UO_153 (O_153,N_4932,N_4958);
xor UO_154 (O_154,N_4931,N_4971);
xnor UO_155 (O_155,N_4903,N_4941);
and UO_156 (O_156,N_4976,N_4967);
nand UO_157 (O_157,N_4991,N_4912);
and UO_158 (O_158,N_4913,N_4992);
nor UO_159 (O_159,N_4985,N_4990);
nor UO_160 (O_160,N_4970,N_4982);
nand UO_161 (O_161,N_4925,N_4937);
xor UO_162 (O_162,N_4904,N_4976);
or UO_163 (O_163,N_4918,N_4925);
and UO_164 (O_164,N_4914,N_4905);
nor UO_165 (O_165,N_4928,N_4963);
nor UO_166 (O_166,N_4983,N_4945);
and UO_167 (O_167,N_4991,N_4910);
nand UO_168 (O_168,N_4906,N_4994);
or UO_169 (O_169,N_4920,N_4995);
nor UO_170 (O_170,N_4935,N_4956);
nand UO_171 (O_171,N_4943,N_4956);
and UO_172 (O_172,N_4976,N_4914);
or UO_173 (O_173,N_4924,N_4952);
xnor UO_174 (O_174,N_4970,N_4930);
or UO_175 (O_175,N_4921,N_4929);
nor UO_176 (O_176,N_4956,N_4907);
nand UO_177 (O_177,N_4995,N_4927);
nor UO_178 (O_178,N_4932,N_4965);
xor UO_179 (O_179,N_4978,N_4986);
and UO_180 (O_180,N_4992,N_4932);
xnor UO_181 (O_181,N_4989,N_4968);
or UO_182 (O_182,N_4953,N_4918);
and UO_183 (O_183,N_4917,N_4920);
or UO_184 (O_184,N_4999,N_4977);
or UO_185 (O_185,N_4937,N_4945);
or UO_186 (O_186,N_4986,N_4982);
or UO_187 (O_187,N_4989,N_4995);
or UO_188 (O_188,N_4997,N_4973);
xor UO_189 (O_189,N_4978,N_4924);
or UO_190 (O_190,N_4995,N_4921);
or UO_191 (O_191,N_4947,N_4987);
nor UO_192 (O_192,N_4989,N_4930);
and UO_193 (O_193,N_4912,N_4968);
nor UO_194 (O_194,N_4924,N_4970);
or UO_195 (O_195,N_4952,N_4975);
nor UO_196 (O_196,N_4910,N_4940);
or UO_197 (O_197,N_4913,N_4920);
or UO_198 (O_198,N_4997,N_4950);
nand UO_199 (O_199,N_4946,N_4962);
nand UO_200 (O_200,N_4957,N_4995);
xor UO_201 (O_201,N_4977,N_4934);
or UO_202 (O_202,N_4934,N_4976);
and UO_203 (O_203,N_4939,N_4996);
xnor UO_204 (O_204,N_4900,N_4923);
nand UO_205 (O_205,N_4917,N_4994);
and UO_206 (O_206,N_4927,N_4941);
or UO_207 (O_207,N_4953,N_4926);
and UO_208 (O_208,N_4994,N_4938);
nor UO_209 (O_209,N_4926,N_4907);
xor UO_210 (O_210,N_4971,N_4962);
xor UO_211 (O_211,N_4930,N_4981);
nand UO_212 (O_212,N_4913,N_4964);
and UO_213 (O_213,N_4941,N_4902);
xnor UO_214 (O_214,N_4941,N_4984);
nor UO_215 (O_215,N_4951,N_4943);
nor UO_216 (O_216,N_4946,N_4908);
or UO_217 (O_217,N_4987,N_4969);
or UO_218 (O_218,N_4955,N_4905);
and UO_219 (O_219,N_4954,N_4930);
xor UO_220 (O_220,N_4983,N_4970);
nand UO_221 (O_221,N_4984,N_4965);
and UO_222 (O_222,N_4927,N_4932);
xor UO_223 (O_223,N_4971,N_4922);
and UO_224 (O_224,N_4990,N_4962);
nand UO_225 (O_225,N_4932,N_4952);
xnor UO_226 (O_226,N_4959,N_4954);
nor UO_227 (O_227,N_4975,N_4970);
or UO_228 (O_228,N_4971,N_4964);
and UO_229 (O_229,N_4967,N_4978);
and UO_230 (O_230,N_4920,N_4906);
and UO_231 (O_231,N_4991,N_4977);
or UO_232 (O_232,N_4938,N_4901);
xor UO_233 (O_233,N_4935,N_4924);
or UO_234 (O_234,N_4911,N_4980);
and UO_235 (O_235,N_4912,N_4952);
nor UO_236 (O_236,N_4944,N_4962);
nand UO_237 (O_237,N_4949,N_4979);
xnor UO_238 (O_238,N_4972,N_4901);
or UO_239 (O_239,N_4932,N_4997);
or UO_240 (O_240,N_4998,N_4957);
or UO_241 (O_241,N_4980,N_4910);
and UO_242 (O_242,N_4942,N_4968);
nand UO_243 (O_243,N_4958,N_4982);
nand UO_244 (O_244,N_4923,N_4985);
xnor UO_245 (O_245,N_4994,N_4992);
nand UO_246 (O_246,N_4936,N_4974);
and UO_247 (O_247,N_4972,N_4957);
and UO_248 (O_248,N_4904,N_4991);
or UO_249 (O_249,N_4911,N_4964);
xor UO_250 (O_250,N_4967,N_4935);
or UO_251 (O_251,N_4936,N_4960);
nand UO_252 (O_252,N_4918,N_4939);
nand UO_253 (O_253,N_4992,N_4976);
and UO_254 (O_254,N_4924,N_4923);
and UO_255 (O_255,N_4969,N_4943);
nor UO_256 (O_256,N_4909,N_4919);
nor UO_257 (O_257,N_4930,N_4985);
nand UO_258 (O_258,N_4941,N_4951);
nand UO_259 (O_259,N_4935,N_4979);
nand UO_260 (O_260,N_4938,N_4934);
and UO_261 (O_261,N_4995,N_4901);
and UO_262 (O_262,N_4908,N_4916);
and UO_263 (O_263,N_4913,N_4999);
xnor UO_264 (O_264,N_4959,N_4984);
xnor UO_265 (O_265,N_4988,N_4906);
nor UO_266 (O_266,N_4953,N_4973);
nor UO_267 (O_267,N_4999,N_4993);
and UO_268 (O_268,N_4903,N_4906);
and UO_269 (O_269,N_4909,N_4917);
or UO_270 (O_270,N_4930,N_4933);
or UO_271 (O_271,N_4971,N_4904);
nand UO_272 (O_272,N_4993,N_4980);
xor UO_273 (O_273,N_4953,N_4911);
nand UO_274 (O_274,N_4916,N_4985);
nand UO_275 (O_275,N_4943,N_4995);
and UO_276 (O_276,N_4933,N_4999);
nand UO_277 (O_277,N_4942,N_4927);
or UO_278 (O_278,N_4927,N_4926);
nand UO_279 (O_279,N_4941,N_4906);
nand UO_280 (O_280,N_4941,N_4969);
and UO_281 (O_281,N_4998,N_4979);
nand UO_282 (O_282,N_4992,N_4957);
nand UO_283 (O_283,N_4972,N_4979);
nor UO_284 (O_284,N_4914,N_4993);
nor UO_285 (O_285,N_4915,N_4939);
and UO_286 (O_286,N_4937,N_4932);
and UO_287 (O_287,N_4902,N_4914);
nand UO_288 (O_288,N_4902,N_4999);
xor UO_289 (O_289,N_4927,N_4978);
or UO_290 (O_290,N_4915,N_4978);
nand UO_291 (O_291,N_4917,N_4949);
nand UO_292 (O_292,N_4907,N_4910);
nand UO_293 (O_293,N_4919,N_4910);
or UO_294 (O_294,N_4973,N_4967);
nor UO_295 (O_295,N_4982,N_4964);
nor UO_296 (O_296,N_4948,N_4971);
xnor UO_297 (O_297,N_4999,N_4963);
nor UO_298 (O_298,N_4969,N_4957);
xor UO_299 (O_299,N_4923,N_4954);
xnor UO_300 (O_300,N_4992,N_4970);
or UO_301 (O_301,N_4907,N_4957);
nor UO_302 (O_302,N_4996,N_4902);
nand UO_303 (O_303,N_4900,N_4965);
and UO_304 (O_304,N_4942,N_4948);
nor UO_305 (O_305,N_4974,N_4931);
xnor UO_306 (O_306,N_4948,N_4921);
or UO_307 (O_307,N_4928,N_4945);
nand UO_308 (O_308,N_4921,N_4942);
or UO_309 (O_309,N_4955,N_4993);
nor UO_310 (O_310,N_4902,N_4971);
and UO_311 (O_311,N_4979,N_4906);
nand UO_312 (O_312,N_4921,N_4985);
nand UO_313 (O_313,N_4954,N_4926);
nand UO_314 (O_314,N_4950,N_4948);
or UO_315 (O_315,N_4963,N_4972);
xor UO_316 (O_316,N_4996,N_4911);
xnor UO_317 (O_317,N_4930,N_4968);
nand UO_318 (O_318,N_4980,N_4967);
nand UO_319 (O_319,N_4925,N_4955);
and UO_320 (O_320,N_4935,N_4931);
xor UO_321 (O_321,N_4988,N_4954);
xor UO_322 (O_322,N_4976,N_4961);
or UO_323 (O_323,N_4943,N_4998);
nor UO_324 (O_324,N_4999,N_4974);
nor UO_325 (O_325,N_4959,N_4944);
nand UO_326 (O_326,N_4983,N_4922);
nand UO_327 (O_327,N_4978,N_4912);
nand UO_328 (O_328,N_4992,N_4954);
nor UO_329 (O_329,N_4942,N_4963);
xnor UO_330 (O_330,N_4997,N_4951);
xnor UO_331 (O_331,N_4968,N_4953);
nand UO_332 (O_332,N_4983,N_4964);
xor UO_333 (O_333,N_4955,N_4908);
or UO_334 (O_334,N_4932,N_4986);
nand UO_335 (O_335,N_4948,N_4991);
and UO_336 (O_336,N_4939,N_4937);
and UO_337 (O_337,N_4907,N_4974);
or UO_338 (O_338,N_4942,N_4984);
and UO_339 (O_339,N_4959,N_4974);
or UO_340 (O_340,N_4912,N_4967);
and UO_341 (O_341,N_4936,N_4935);
nand UO_342 (O_342,N_4957,N_4913);
and UO_343 (O_343,N_4984,N_4938);
xnor UO_344 (O_344,N_4946,N_4935);
nand UO_345 (O_345,N_4905,N_4951);
xor UO_346 (O_346,N_4982,N_4999);
nand UO_347 (O_347,N_4936,N_4982);
nand UO_348 (O_348,N_4902,N_4935);
xnor UO_349 (O_349,N_4907,N_4927);
xnor UO_350 (O_350,N_4917,N_4995);
and UO_351 (O_351,N_4938,N_4900);
xor UO_352 (O_352,N_4965,N_4910);
nand UO_353 (O_353,N_4984,N_4918);
xor UO_354 (O_354,N_4953,N_4943);
and UO_355 (O_355,N_4939,N_4932);
and UO_356 (O_356,N_4967,N_4934);
nor UO_357 (O_357,N_4920,N_4997);
nand UO_358 (O_358,N_4950,N_4933);
and UO_359 (O_359,N_4942,N_4982);
xnor UO_360 (O_360,N_4977,N_4917);
xnor UO_361 (O_361,N_4945,N_4977);
and UO_362 (O_362,N_4956,N_4955);
nand UO_363 (O_363,N_4970,N_4995);
xnor UO_364 (O_364,N_4954,N_4952);
and UO_365 (O_365,N_4997,N_4906);
nor UO_366 (O_366,N_4911,N_4927);
xor UO_367 (O_367,N_4918,N_4904);
xor UO_368 (O_368,N_4936,N_4964);
or UO_369 (O_369,N_4944,N_4980);
or UO_370 (O_370,N_4976,N_4919);
nand UO_371 (O_371,N_4929,N_4982);
nand UO_372 (O_372,N_4916,N_4946);
and UO_373 (O_373,N_4961,N_4994);
nand UO_374 (O_374,N_4963,N_4985);
or UO_375 (O_375,N_4949,N_4960);
xor UO_376 (O_376,N_4921,N_4907);
nor UO_377 (O_377,N_4956,N_4934);
nand UO_378 (O_378,N_4996,N_4975);
or UO_379 (O_379,N_4911,N_4926);
xor UO_380 (O_380,N_4998,N_4944);
nand UO_381 (O_381,N_4912,N_4950);
or UO_382 (O_382,N_4973,N_4904);
or UO_383 (O_383,N_4974,N_4954);
nand UO_384 (O_384,N_4969,N_4944);
xnor UO_385 (O_385,N_4932,N_4994);
nor UO_386 (O_386,N_4992,N_4963);
and UO_387 (O_387,N_4984,N_4931);
and UO_388 (O_388,N_4946,N_4907);
xor UO_389 (O_389,N_4920,N_4983);
nand UO_390 (O_390,N_4958,N_4919);
nand UO_391 (O_391,N_4951,N_4974);
nand UO_392 (O_392,N_4928,N_4910);
xnor UO_393 (O_393,N_4903,N_4982);
and UO_394 (O_394,N_4932,N_4941);
or UO_395 (O_395,N_4957,N_4963);
or UO_396 (O_396,N_4960,N_4903);
and UO_397 (O_397,N_4919,N_4934);
or UO_398 (O_398,N_4900,N_4992);
nand UO_399 (O_399,N_4923,N_4964);
and UO_400 (O_400,N_4962,N_4901);
and UO_401 (O_401,N_4955,N_4974);
and UO_402 (O_402,N_4920,N_4977);
or UO_403 (O_403,N_4915,N_4961);
nor UO_404 (O_404,N_4977,N_4919);
nor UO_405 (O_405,N_4981,N_4911);
or UO_406 (O_406,N_4912,N_4909);
and UO_407 (O_407,N_4902,N_4977);
and UO_408 (O_408,N_4986,N_4937);
and UO_409 (O_409,N_4953,N_4914);
nand UO_410 (O_410,N_4983,N_4988);
nand UO_411 (O_411,N_4956,N_4986);
or UO_412 (O_412,N_4901,N_4948);
or UO_413 (O_413,N_4965,N_4964);
xor UO_414 (O_414,N_4940,N_4966);
nor UO_415 (O_415,N_4908,N_4919);
nand UO_416 (O_416,N_4917,N_4903);
and UO_417 (O_417,N_4999,N_4991);
nand UO_418 (O_418,N_4970,N_4903);
or UO_419 (O_419,N_4932,N_4923);
nand UO_420 (O_420,N_4931,N_4970);
or UO_421 (O_421,N_4969,N_4900);
and UO_422 (O_422,N_4986,N_4902);
nor UO_423 (O_423,N_4993,N_4949);
or UO_424 (O_424,N_4956,N_4940);
nand UO_425 (O_425,N_4947,N_4933);
and UO_426 (O_426,N_4901,N_4903);
nor UO_427 (O_427,N_4985,N_4917);
nor UO_428 (O_428,N_4930,N_4975);
xor UO_429 (O_429,N_4982,N_4907);
or UO_430 (O_430,N_4985,N_4992);
or UO_431 (O_431,N_4904,N_4997);
xnor UO_432 (O_432,N_4953,N_4955);
nand UO_433 (O_433,N_4939,N_4917);
nand UO_434 (O_434,N_4948,N_4961);
or UO_435 (O_435,N_4969,N_4961);
or UO_436 (O_436,N_4996,N_4993);
and UO_437 (O_437,N_4938,N_4925);
nand UO_438 (O_438,N_4972,N_4929);
xnor UO_439 (O_439,N_4901,N_4933);
xor UO_440 (O_440,N_4982,N_4924);
and UO_441 (O_441,N_4951,N_4914);
and UO_442 (O_442,N_4997,N_4931);
xnor UO_443 (O_443,N_4900,N_4926);
nor UO_444 (O_444,N_4943,N_4980);
and UO_445 (O_445,N_4913,N_4998);
or UO_446 (O_446,N_4912,N_4962);
or UO_447 (O_447,N_4921,N_4978);
and UO_448 (O_448,N_4981,N_4985);
nor UO_449 (O_449,N_4905,N_4981);
nor UO_450 (O_450,N_4954,N_4961);
nor UO_451 (O_451,N_4995,N_4912);
or UO_452 (O_452,N_4960,N_4902);
or UO_453 (O_453,N_4957,N_4928);
nand UO_454 (O_454,N_4941,N_4982);
nor UO_455 (O_455,N_4933,N_4972);
nand UO_456 (O_456,N_4904,N_4900);
xor UO_457 (O_457,N_4967,N_4904);
and UO_458 (O_458,N_4979,N_4944);
nor UO_459 (O_459,N_4972,N_4959);
or UO_460 (O_460,N_4913,N_4934);
nand UO_461 (O_461,N_4959,N_4973);
nand UO_462 (O_462,N_4919,N_4997);
and UO_463 (O_463,N_4984,N_4904);
or UO_464 (O_464,N_4972,N_4908);
and UO_465 (O_465,N_4976,N_4945);
nand UO_466 (O_466,N_4965,N_4970);
nor UO_467 (O_467,N_4952,N_4922);
or UO_468 (O_468,N_4951,N_4922);
xor UO_469 (O_469,N_4918,N_4972);
and UO_470 (O_470,N_4925,N_4981);
or UO_471 (O_471,N_4954,N_4986);
and UO_472 (O_472,N_4974,N_4900);
nor UO_473 (O_473,N_4917,N_4958);
xor UO_474 (O_474,N_4938,N_4902);
xnor UO_475 (O_475,N_4940,N_4908);
xor UO_476 (O_476,N_4954,N_4955);
xor UO_477 (O_477,N_4939,N_4997);
nand UO_478 (O_478,N_4904,N_4974);
or UO_479 (O_479,N_4992,N_4920);
nand UO_480 (O_480,N_4944,N_4909);
nand UO_481 (O_481,N_4937,N_4950);
nand UO_482 (O_482,N_4934,N_4905);
and UO_483 (O_483,N_4922,N_4903);
nor UO_484 (O_484,N_4967,N_4983);
xor UO_485 (O_485,N_4920,N_4971);
or UO_486 (O_486,N_4984,N_4975);
xnor UO_487 (O_487,N_4938,N_4992);
and UO_488 (O_488,N_4956,N_4996);
or UO_489 (O_489,N_4952,N_4992);
or UO_490 (O_490,N_4973,N_4983);
and UO_491 (O_491,N_4926,N_4971);
and UO_492 (O_492,N_4952,N_4961);
xnor UO_493 (O_493,N_4974,N_4928);
and UO_494 (O_494,N_4981,N_4907);
nand UO_495 (O_495,N_4903,N_4921);
and UO_496 (O_496,N_4900,N_4957);
nand UO_497 (O_497,N_4903,N_4997);
or UO_498 (O_498,N_4948,N_4977);
xor UO_499 (O_499,N_4973,N_4900);
nand UO_500 (O_500,N_4916,N_4982);
nand UO_501 (O_501,N_4917,N_4973);
xor UO_502 (O_502,N_4900,N_4940);
xnor UO_503 (O_503,N_4985,N_4911);
and UO_504 (O_504,N_4917,N_4928);
or UO_505 (O_505,N_4948,N_4986);
and UO_506 (O_506,N_4974,N_4991);
nor UO_507 (O_507,N_4992,N_4941);
xnor UO_508 (O_508,N_4918,N_4908);
nand UO_509 (O_509,N_4936,N_4938);
xor UO_510 (O_510,N_4947,N_4980);
xor UO_511 (O_511,N_4964,N_4963);
and UO_512 (O_512,N_4919,N_4955);
nand UO_513 (O_513,N_4936,N_4942);
and UO_514 (O_514,N_4963,N_4906);
or UO_515 (O_515,N_4940,N_4927);
and UO_516 (O_516,N_4975,N_4922);
or UO_517 (O_517,N_4949,N_4984);
and UO_518 (O_518,N_4974,N_4944);
or UO_519 (O_519,N_4976,N_4937);
nand UO_520 (O_520,N_4929,N_4939);
nand UO_521 (O_521,N_4921,N_4937);
or UO_522 (O_522,N_4933,N_4902);
and UO_523 (O_523,N_4984,N_4994);
or UO_524 (O_524,N_4952,N_4991);
xnor UO_525 (O_525,N_4933,N_4955);
and UO_526 (O_526,N_4967,N_4997);
nor UO_527 (O_527,N_4910,N_4927);
xnor UO_528 (O_528,N_4991,N_4918);
or UO_529 (O_529,N_4979,N_4909);
nor UO_530 (O_530,N_4980,N_4946);
nand UO_531 (O_531,N_4996,N_4930);
xor UO_532 (O_532,N_4924,N_4944);
and UO_533 (O_533,N_4995,N_4960);
or UO_534 (O_534,N_4996,N_4994);
xnor UO_535 (O_535,N_4927,N_4972);
nand UO_536 (O_536,N_4936,N_4908);
xnor UO_537 (O_537,N_4996,N_4979);
xnor UO_538 (O_538,N_4955,N_4946);
nand UO_539 (O_539,N_4948,N_4902);
nand UO_540 (O_540,N_4983,N_4915);
and UO_541 (O_541,N_4965,N_4935);
and UO_542 (O_542,N_4909,N_4991);
xnor UO_543 (O_543,N_4993,N_4992);
or UO_544 (O_544,N_4924,N_4926);
xor UO_545 (O_545,N_4971,N_4934);
xor UO_546 (O_546,N_4918,N_4926);
nor UO_547 (O_547,N_4916,N_4915);
nand UO_548 (O_548,N_4935,N_4998);
nor UO_549 (O_549,N_4969,N_4917);
nand UO_550 (O_550,N_4938,N_4970);
xnor UO_551 (O_551,N_4916,N_4941);
or UO_552 (O_552,N_4976,N_4943);
nor UO_553 (O_553,N_4983,N_4982);
xnor UO_554 (O_554,N_4950,N_4982);
nand UO_555 (O_555,N_4987,N_4941);
xor UO_556 (O_556,N_4933,N_4944);
nand UO_557 (O_557,N_4925,N_4944);
nor UO_558 (O_558,N_4993,N_4938);
xor UO_559 (O_559,N_4925,N_4958);
xor UO_560 (O_560,N_4943,N_4929);
xor UO_561 (O_561,N_4940,N_4982);
nor UO_562 (O_562,N_4963,N_4986);
xnor UO_563 (O_563,N_4984,N_4990);
nor UO_564 (O_564,N_4920,N_4964);
and UO_565 (O_565,N_4910,N_4938);
or UO_566 (O_566,N_4951,N_4971);
xnor UO_567 (O_567,N_4949,N_4923);
xnor UO_568 (O_568,N_4907,N_4975);
or UO_569 (O_569,N_4983,N_4952);
xor UO_570 (O_570,N_4972,N_4920);
or UO_571 (O_571,N_4943,N_4990);
or UO_572 (O_572,N_4970,N_4923);
or UO_573 (O_573,N_4922,N_4948);
nor UO_574 (O_574,N_4933,N_4990);
nand UO_575 (O_575,N_4923,N_4959);
xor UO_576 (O_576,N_4951,N_4916);
nor UO_577 (O_577,N_4951,N_4906);
or UO_578 (O_578,N_4926,N_4999);
xor UO_579 (O_579,N_4939,N_4990);
and UO_580 (O_580,N_4972,N_4904);
and UO_581 (O_581,N_4937,N_4987);
xnor UO_582 (O_582,N_4943,N_4927);
nor UO_583 (O_583,N_4918,N_4927);
or UO_584 (O_584,N_4900,N_4972);
or UO_585 (O_585,N_4902,N_4923);
nor UO_586 (O_586,N_4999,N_4920);
and UO_587 (O_587,N_4973,N_4901);
nand UO_588 (O_588,N_4930,N_4909);
nor UO_589 (O_589,N_4900,N_4946);
xnor UO_590 (O_590,N_4904,N_4950);
xnor UO_591 (O_591,N_4902,N_4962);
or UO_592 (O_592,N_4926,N_4955);
nand UO_593 (O_593,N_4951,N_4930);
nor UO_594 (O_594,N_4900,N_4911);
nand UO_595 (O_595,N_4904,N_4901);
nor UO_596 (O_596,N_4922,N_4996);
or UO_597 (O_597,N_4919,N_4994);
and UO_598 (O_598,N_4961,N_4926);
and UO_599 (O_599,N_4915,N_4952);
nand UO_600 (O_600,N_4998,N_4931);
nor UO_601 (O_601,N_4990,N_4946);
and UO_602 (O_602,N_4946,N_4969);
and UO_603 (O_603,N_4915,N_4995);
or UO_604 (O_604,N_4991,N_4996);
nor UO_605 (O_605,N_4955,N_4966);
nand UO_606 (O_606,N_4993,N_4998);
nor UO_607 (O_607,N_4909,N_4920);
xnor UO_608 (O_608,N_4995,N_4978);
nand UO_609 (O_609,N_4928,N_4973);
or UO_610 (O_610,N_4995,N_4905);
nor UO_611 (O_611,N_4964,N_4980);
xnor UO_612 (O_612,N_4947,N_4910);
and UO_613 (O_613,N_4952,N_4934);
xnor UO_614 (O_614,N_4910,N_4961);
nand UO_615 (O_615,N_4922,N_4981);
xor UO_616 (O_616,N_4918,N_4948);
or UO_617 (O_617,N_4964,N_4912);
xnor UO_618 (O_618,N_4920,N_4918);
and UO_619 (O_619,N_4993,N_4997);
and UO_620 (O_620,N_4907,N_4932);
or UO_621 (O_621,N_4992,N_4921);
or UO_622 (O_622,N_4952,N_4947);
xnor UO_623 (O_623,N_4936,N_4951);
or UO_624 (O_624,N_4991,N_4919);
xor UO_625 (O_625,N_4994,N_4948);
nand UO_626 (O_626,N_4951,N_4969);
and UO_627 (O_627,N_4970,N_4925);
nor UO_628 (O_628,N_4937,N_4918);
xnor UO_629 (O_629,N_4939,N_4907);
xor UO_630 (O_630,N_4919,N_4959);
nor UO_631 (O_631,N_4975,N_4978);
and UO_632 (O_632,N_4928,N_4956);
nand UO_633 (O_633,N_4998,N_4907);
nand UO_634 (O_634,N_4903,N_4933);
nor UO_635 (O_635,N_4909,N_4945);
nand UO_636 (O_636,N_4936,N_4924);
nand UO_637 (O_637,N_4956,N_4988);
and UO_638 (O_638,N_4964,N_4938);
nor UO_639 (O_639,N_4981,N_4923);
nor UO_640 (O_640,N_4961,N_4906);
or UO_641 (O_641,N_4939,N_4935);
xnor UO_642 (O_642,N_4935,N_4990);
nand UO_643 (O_643,N_4912,N_4910);
xor UO_644 (O_644,N_4928,N_4975);
and UO_645 (O_645,N_4920,N_4926);
nor UO_646 (O_646,N_4918,N_4902);
xnor UO_647 (O_647,N_4921,N_4963);
nor UO_648 (O_648,N_4953,N_4908);
nand UO_649 (O_649,N_4949,N_4904);
and UO_650 (O_650,N_4944,N_4939);
or UO_651 (O_651,N_4927,N_4977);
and UO_652 (O_652,N_4953,N_4929);
xor UO_653 (O_653,N_4995,N_4983);
xor UO_654 (O_654,N_4983,N_4993);
xor UO_655 (O_655,N_4968,N_4972);
nand UO_656 (O_656,N_4999,N_4990);
or UO_657 (O_657,N_4938,N_4917);
nor UO_658 (O_658,N_4929,N_4914);
nor UO_659 (O_659,N_4928,N_4999);
nor UO_660 (O_660,N_4956,N_4972);
nand UO_661 (O_661,N_4950,N_4979);
and UO_662 (O_662,N_4955,N_4988);
or UO_663 (O_663,N_4959,N_4924);
nand UO_664 (O_664,N_4983,N_4901);
nor UO_665 (O_665,N_4994,N_4915);
or UO_666 (O_666,N_4960,N_4958);
xor UO_667 (O_667,N_4958,N_4901);
xor UO_668 (O_668,N_4924,N_4905);
and UO_669 (O_669,N_4940,N_4989);
and UO_670 (O_670,N_4918,N_4962);
nor UO_671 (O_671,N_4918,N_4943);
and UO_672 (O_672,N_4993,N_4924);
and UO_673 (O_673,N_4945,N_4964);
or UO_674 (O_674,N_4947,N_4909);
nand UO_675 (O_675,N_4927,N_4955);
nor UO_676 (O_676,N_4935,N_4903);
nor UO_677 (O_677,N_4979,N_4955);
nand UO_678 (O_678,N_4933,N_4934);
xor UO_679 (O_679,N_4959,N_4980);
or UO_680 (O_680,N_4909,N_4939);
nor UO_681 (O_681,N_4964,N_4957);
xor UO_682 (O_682,N_4933,N_4969);
or UO_683 (O_683,N_4961,N_4987);
or UO_684 (O_684,N_4992,N_4908);
nand UO_685 (O_685,N_4998,N_4938);
xnor UO_686 (O_686,N_4989,N_4925);
and UO_687 (O_687,N_4947,N_4946);
nand UO_688 (O_688,N_4922,N_4961);
xor UO_689 (O_689,N_4946,N_4948);
xnor UO_690 (O_690,N_4978,N_4946);
or UO_691 (O_691,N_4923,N_4971);
nand UO_692 (O_692,N_4929,N_4989);
nand UO_693 (O_693,N_4931,N_4924);
and UO_694 (O_694,N_4900,N_4995);
nor UO_695 (O_695,N_4909,N_4929);
xnor UO_696 (O_696,N_4944,N_4992);
nand UO_697 (O_697,N_4972,N_4960);
and UO_698 (O_698,N_4932,N_4960);
nor UO_699 (O_699,N_4975,N_4994);
xnor UO_700 (O_700,N_4966,N_4960);
or UO_701 (O_701,N_4969,N_4909);
and UO_702 (O_702,N_4944,N_4915);
xnor UO_703 (O_703,N_4904,N_4941);
xnor UO_704 (O_704,N_4963,N_4945);
nor UO_705 (O_705,N_4988,N_4932);
and UO_706 (O_706,N_4974,N_4933);
xnor UO_707 (O_707,N_4950,N_4976);
nor UO_708 (O_708,N_4998,N_4909);
or UO_709 (O_709,N_4930,N_4944);
nand UO_710 (O_710,N_4970,N_4900);
nor UO_711 (O_711,N_4910,N_4967);
and UO_712 (O_712,N_4961,N_4951);
nor UO_713 (O_713,N_4990,N_4944);
nor UO_714 (O_714,N_4959,N_4981);
nor UO_715 (O_715,N_4960,N_4913);
nand UO_716 (O_716,N_4938,N_4977);
and UO_717 (O_717,N_4941,N_4930);
and UO_718 (O_718,N_4932,N_4956);
or UO_719 (O_719,N_4976,N_4909);
or UO_720 (O_720,N_4996,N_4950);
nand UO_721 (O_721,N_4948,N_4903);
nor UO_722 (O_722,N_4943,N_4950);
or UO_723 (O_723,N_4992,N_4965);
and UO_724 (O_724,N_4938,N_4907);
nor UO_725 (O_725,N_4990,N_4996);
and UO_726 (O_726,N_4990,N_4928);
or UO_727 (O_727,N_4958,N_4969);
nor UO_728 (O_728,N_4948,N_4968);
or UO_729 (O_729,N_4972,N_4967);
nor UO_730 (O_730,N_4997,N_4982);
xnor UO_731 (O_731,N_4999,N_4966);
or UO_732 (O_732,N_4956,N_4944);
xnor UO_733 (O_733,N_4912,N_4980);
xnor UO_734 (O_734,N_4980,N_4974);
xnor UO_735 (O_735,N_4967,N_4950);
or UO_736 (O_736,N_4946,N_4999);
and UO_737 (O_737,N_4930,N_4901);
and UO_738 (O_738,N_4956,N_4973);
nand UO_739 (O_739,N_4947,N_4970);
or UO_740 (O_740,N_4952,N_4969);
or UO_741 (O_741,N_4954,N_4903);
and UO_742 (O_742,N_4942,N_4909);
xnor UO_743 (O_743,N_4927,N_4929);
nor UO_744 (O_744,N_4959,N_4951);
nor UO_745 (O_745,N_4988,N_4961);
nand UO_746 (O_746,N_4972,N_4993);
nand UO_747 (O_747,N_4947,N_4995);
and UO_748 (O_748,N_4923,N_4979);
xor UO_749 (O_749,N_4994,N_4944);
nand UO_750 (O_750,N_4986,N_4910);
xnor UO_751 (O_751,N_4983,N_4927);
xnor UO_752 (O_752,N_4982,N_4915);
xnor UO_753 (O_753,N_4915,N_4955);
nand UO_754 (O_754,N_4900,N_4994);
nand UO_755 (O_755,N_4990,N_4975);
nor UO_756 (O_756,N_4954,N_4944);
nor UO_757 (O_757,N_4955,N_4961);
or UO_758 (O_758,N_4984,N_4935);
nor UO_759 (O_759,N_4928,N_4949);
or UO_760 (O_760,N_4905,N_4900);
nand UO_761 (O_761,N_4987,N_4928);
or UO_762 (O_762,N_4947,N_4978);
or UO_763 (O_763,N_4934,N_4922);
nand UO_764 (O_764,N_4914,N_4969);
or UO_765 (O_765,N_4923,N_4921);
xnor UO_766 (O_766,N_4945,N_4965);
nand UO_767 (O_767,N_4951,N_4902);
xor UO_768 (O_768,N_4937,N_4942);
nor UO_769 (O_769,N_4971,N_4976);
xnor UO_770 (O_770,N_4997,N_4942);
or UO_771 (O_771,N_4950,N_4913);
and UO_772 (O_772,N_4903,N_4959);
nand UO_773 (O_773,N_4903,N_4956);
xnor UO_774 (O_774,N_4961,N_4966);
and UO_775 (O_775,N_4962,N_4948);
xor UO_776 (O_776,N_4977,N_4936);
nor UO_777 (O_777,N_4971,N_4915);
or UO_778 (O_778,N_4999,N_4931);
nor UO_779 (O_779,N_4982,N_4960);
and UO_780 (O_780,N_4988,N_4992);
xor UO_781 (O_781,N_4945,N_4926);
nor UO_782 (O_782,N_4959,N_4985);
nand UO_783 (O_783,N_4966,N_4957);
nor UO_784 (O_784,N_4965,N_4980);
and UO_785 (O_785,N_4929,N_4994);
or UO_786 (O_786,N_4915,N_4945);
or UO_787 (O_787,N_4906,N_4914);
xor UO_788 (O_788,N_4989,N_4926);
and UO_789 (O_789,N_4973,N_4964);
nor UO_790 (O_790,N_4929,N_4951);
or UO_791 (O_791,N_4988,N_4964);
or UO_792 (O_792,N_4929,N_4996);
nand UO_793 (O_793,N_4914,N_4924);
and UO_794 (O_794,N_4931,N_4996);
nor UO_795 (O_795,N_4926,N_4980);
nand UO_796 (O_796,N_4986,N_4928);
xnor UO_797 (O_797,N_4956,N_4961);
nor UO_798 (O_798,N_4972,N_4999);
nand UO_799 (O_799,N_4958,N_4971);
xnor UO_800 (O_800,N_4932,N_4918);
xnor UO_801 (O_801,N_4971,N_4995);
nor UO_802 (O_802,N_4983,N_4900);
nand UO_803 (O_803,N_4934,N_4940);
nand UO_804 (O_804,N_4939,N_4994);
nor UO_805 (O_805,N_4994,N_4987);
xor UO_806 (O_806,N_4970,N_4991);
or UO_807 (O_807,N_4941,N_4961);
nand UO_808 (O_808,N_4966,N_4935);
or UO_809 (O_809,N_4962,N_4954);
nand UO_810 (O_810,N_4923,N_4914);
xnor UO_811 (O_811,N_4955,N_4968);
and UO_812 (O_812,N_4926,N_4940);
or UO_813 (O_813,N_4964,N_4991);
or UO_814 (O_814,N_4995,N_4975);
or UO_815 (O_815,N_4950,N_4932);
nand UO_816 (O_816,N_4906,N_4991);
and UO_817 (O_817,N_4940,N_4971);
or UO_818 (O_818,N_4939,N_4948);
nor UO_819 (O_819,N_4905,N_4985);
nor UO_820 (O_820,N_4955,N_4917);
nand UO_821 (O_821,N_4965,N_4959);
nor UO_822 (O_822,N_4948,N_4917);
and UO_823 (O_823,N_4950,N_4935);
xnor UO_824 (O_824,N_4936,N_4994);
nor UO_825 (O_825,N_4993,N_4909);
nand UO_826 (O_826,N_4944,N_4963);
xnor UO_827 (O_827,N_4993,N_4953);
nor UO_828 (O_828,N_4988,N_4901);
nor UO_829 (O_829,N_4959,N_4902);
nand UO_830 (O_830,N_4905,N_4986);
nor UO_831 (O_831,N_4967,N_4921);
and UO_832 (O_832,N_4938,N_4908);
nor UO_833 (O_833,N_4997,N_4912);
and UO_834 (O_834,N_4985,N_4924);
and UO_835 (O_835,N_4936,N_4993);
nand UO_836 (O_836,N_4980,N_4998);
nand UO_837 (O_837,N_4986,N_4913);
nor UO_838 (O_838,N_4930,N_4958);
or UO_839 (O_839,N_4928,N_4981);
xnor UO_840 (O_840,N_4978,N_4959);
or UO_841 (O_841,N_4905,N_4979);
nand UO_842 (O_842,N_4962,N_4936);
or UO_843 (O_843,N_4951,N_4944);
xor UO_844 (O_844,N_4942,N_4971);
xor UO_845 (O_845,N_4935,N_4954);
nor UO_846 (O_846,N_4930,N_4916);
or UO_847 (O_847,N_4955,N_4939);
and UO_848 (O_848,N_4921,N_4981);
xnor UO_849 (O_849,N_4963,N_4910);
nand UO_850 (O_850,N_4916,N_4907);
or UO_851 (O_851,N_4943,N_4959);
and UO_852 (O_852,N_4991,N_4951);
or UO_853 (O_853,N_4910,N_4931);
or UO_854 (O_854,N_4901,N_4981);
nor UO_855 (O_855,N_4987,N_4925);
xor UO_856 (O_856,N_4992,N_4949);
nor UO_857 (O_857,N_4948,N_4963);
nand UO_858 (O_858,N_4970,N_4904);
nand UO_859 (O_859,N_4906,N_4964);
nand UO_860 (O_860,N_4938,N_4971);
nand UO_861 (O_861,N_4939,N_4912);
and UO_862 (O_862,N_4992,N_4905);
and UO_863 (O_863,N_4907,N_4948);
nor UO_864 (O_864,N_4993,N_4961);
nand UO_865 (O_865,N_4909,N_4966);
nor UO_866 (O_866,N_4951,N_4949);
or UO_867 (O_867,N_4960,N_4925);
nor UO_868 (O_868,N_4979,N_4934);
and UO_869 (O_869,N_4937,N_4964);
and UO_870 (O_870,N_4949,N_4975);
and UO_871 (O_871,N_4960,N_4974);
or UO_872 (O_872,N_4961,N_4939);
nor UO_873 (O_873,N_4954,N_4983);
and UO_874 (O_874,N_4913,N_4991);
or UO_875 (O_875,N_4930,N_4900);
and UO_876 (O_876,N_4912,N_4902);
xnor UO_877 (O_877,N_4964,N_4944);
and UO_878 (O_878,N_4918,N_4999);
nor UO_879 (O_879,N_4949,N_4947);
or UO_880 (O_880,N_4931,N_4985);
xor UO_881 (O_881,N_4940,N_4976);
nor UO_882 (O_882,N_4901,N_4970);
xnor UO_883 (O_883,N_4933,N_4978);
nand UO_884 (O_884,N_4954,N_4912);
xnor UO_885 (O_885,N_4914,N_4943);
xor UO_886 (O_886,N_4968,N_4920);
or UO_887 (O_887,N_4988,N_4971);
xnor UO_888 (O_888,N_4977,N_4914);
and UO_889 (O_889,N_4970,N_4955);
nand UO_890 (O_890,N_4964,N_4900);
and UO_891 (O_891,N_4942,N_4956);
or UO_892 (O_892,N_4959,N_4929);
nor UO_893 (O_893,N_4961,N_4903);
xor UO_894 (O_894,N_4934,N_4968);
nor UO_895 (O_895,N_4970,N_4994);
xor UO_896 (O_896,N_4913,N_4963);
xnor UO_897 (O_897,N_4911,N_4924);
nor UO_898 (O_898,N_4977,N_4980);
or UO_899 (O_899,N_4922,N_4910);
nand UO_900 (O_900,N_4989,N_4906);
and UO_901 (O_901,N_4922,N_4935);
and UO_902 (O_902,N_4942,N_4976);
or UO_903 (O_903,N_4937,N_4957);
nor UO_904 (O_904,N_4964,N_4908);
and UO_905 (O_905,N_4939,N_4988);
nand UO_906 (O_906,N_4967,N_4917);
and UO_907 (O_907,N_4942,N_4914);
nor UO_908 (O_908,N_4947,N_4976);
nor UO_909 (O_909,N_4900,N_4928);
xor UO_910 (O_910,N_4981,N_4916);
nor UO_911 (O_911,N_4975,N_4934);
or UO_912 (O_912,N_4940,N_4975);
nand UO_913 (O_913,N_4927,N_4991);
nand UO_914 (O_914,N_4970,N_4922);
or UO_915 (O_915,N_4954,N_4978);
nand UO_916 (O_916,N_4969,N_4938);
and UO_917 (O_917,N_4900,N_4967);
xor UO_918 (O_918,N_4971,N_4982);
nand UO_919 (O_919,N_4915,N_4911);
and UO_920 (O_920,N_4916,N_4920);
and UO_921 (O_921,N_4993,N_4963);
or UO_922 (O_922,N_4916,N_4992);
and UO_923 (O_923,N_4997,N_4966);
and UO_924 (O_924,N_4902,N_4903);
nor UO_925 (O_925,N_4917,N_4902);
or UO_926 (O_926,N_4949,N_4957);
nand UO_927 (O_927,N_4939,N_4963);
nand UO_928 (O_928,N_4998,N_4905);
and UO_929 (O_929,N_4947,N_4984);
nor UO_930 (O_930,N_4910,N_4952);
or UO_931 (O_931,N_4954,N_4993);
xor UO_932 (O_932,N_4928,N_4964);
or UO_933 (O_933,N_4912,N_4971);
and UO_934 (O_934,N_4932,N_4975);
nand UO_935 (O_935,N_4956,N_4980);
nor UO_936 (O_936,N_4996,N_4955);
and UO_937 (O_937,N_4975,N_4956);
nand UO_938 (O_938,N_4980,N_4990);
xnor UO_939 (O_939,N_4990,N_4956);
xnor UO_940 (O_940,N_4995,N_4952);
and UO_941 (O_941,N_4964,N_4917);
nor UO_942 (O_942,N_4954,N_4982);
and UO_943 (O_943,N_4997,N_4909);
or UO_944 (O_944,N_4928,N_4935);
and UO_945 (O_945,N_4943,N_4900);
nor UO_946 (O_946,N_4905,N_4960);
nor UO_947 (O_947,N_4962,N_4905);
xnor UO_948 (O_948,N_4929,N_4975);
nor UO_949 (O_949,N_4987,N_4990);
nand UO_950 (O_950,N_4906,N_4996);
nor UO_951 (O_951,N_4966,N_4981);
nand UO_952 (O_952,N_4907,N_4978);
and UO_953 (O_953,N_4983,N_4908);
and UO_954 (O_954,N_4992,N_4919);
and UO_955 (O_955,N_4978,N_4969);
or UO_956 (O_956,N_4956,N_4946);
xnor UO_957 (O_957,N_4984,N_4973);
and UO_958 (O_958,N_4931,N_4976);
xnor UO_959 (O_959,N_4914,N_4909);
or UO_960 (O_960,N_4992,N_4973);
nor UO_961 (O_961,N_4929,N_4966);
nand UO_962 (O_962,N_4925,N_4983);
xor UO_963 (O_963,N_4906,N_4912);
nand UO_964 (O_964,N_4916,N_4971);
or UO_965 (O_965,N_4990,N_4908);
nor UO_966 (O_966,N_4928,N_4976);
or UO_967 (O_967,N_4978,N_4952);
nand UO_968 (O_968,N_4985,N_4995);
or UO_969 (O_969,N_4957,N_4933);
or UO_970 (O_970,N_4931,N_4955);
or UO_971 (O_971,N_4934,N_4931);
xnor UO_972 (O_972,N_4924,N_4916);
or UO_973 (O_973,N_4992,N_4928);
nand UO_974 (O_974,N_4972,N_4952);
nor UO_975 (O_975,N_4936,N_4916);
nor UO_976 (O_976,N_4989,N_4960);
nand UO_977 (O_977,N_4944,N_4926);
and UO_978 (O_978,N_4991,N_4980);
xor UO_979 (O_979,N_4982,N_4956);
nor UO_980 (O_980,N_4986,N_4950);
and UO_981 (O_981,N_4918,N_4946);
xor UO_982 (O_982,N_4920,N_4931);
or UO_983 (O_983,N_4991,N_4929);
xnor UO_984 (O_984,N_4927,N_4956);
or UO_985 (O_985,N_4994,N_4995);
and UO_986 (O_986,N_4930,N_4995);
xor UO_987 (O_987,N_4962,N_4981);
xor UO_988 (O_988,N_4997,N_4929);
nand UO_989 (O_989,N_4934,N_4901);
nor UO_990 (O_990,N_4954,N_4938);
and UO_991 (O_991,N_4906,N_4968);
nand UO_992 (O_992,N_4993,N_4917);
nand UO_993 (O_993,N_4904,N_4935);
xor UO_994 (O_994,N_4958,N_4972);
or UO_995 (O_995,N_4975,N_4919);
xnor UO_996 (O_996,N_4924,N_4940);
and UO_997 (O_997,N_4940,N_4907);
xnor UO_998 (O_998,N_4945,N_4934);
nand UO_999 (O_999,N_4903,N_4938);
endmodule