module basic_1500_15000_2000_3_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10014,N_10016,N_10017,N_10019,N_10020,N_10022,N_10023,N_10024,N_10025,N_10026,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10045,N_10046,N_10048,N_10051,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10081,N_10082,N_10083,N_10085,N_10086,N_10087,N_10089,N_10091,N_10092,N_10094,N_10095,N_10096,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10107,N_10108,N_10110,N_10112,N_10113,N_10114,N_10115,N_10116,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10125,N_10126,N_10127,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10161,N_10163,N_10165,N_10166,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10180,N_10181,N_10182,N_10183,N_10185,N_10186,N_10187,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10201,N_10203,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10225,N_10226,N_10227,N_10229,N_10230,N_10231,N_10234,N_10235,N_10236,N_10238,N_10241,N_10243,N_10244,N_10245,N_10246,N_10248,N_10249,N_10250,N_10251,N_10253,N_10254,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10269,N_10271,N_10273,N_10274,N_10275,N_10276,N_10278,N_10280,N_10281,N_10282,N_10283,N_10285,N_10286,N_10287,N_10293,N_10294,N_10296,N_10297,N_10301,N_10303,N_10304,N_10307,N_10308,N_10309,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10339,N_10340,N_10341,N_10342,N_10344,N_10345,N_10346,N_10347,N_10349,N_10353,N_10355,N_10356,N_10357,N_10358,N_10359,N_10361,N_10362,N_10363,N_10364,N_10365,N_10369,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10387,N_10388,N_10389,N_10390,N_10391,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10401,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10410,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10422,N_10423,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10455,N_10456,N_10457,N_10458,N_10459,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10485,N_10486,N_10489,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10513,N_10515,N_10517,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10531,N_10535,N_10536,N_10538,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10561,N_10563,N_10564,N_10565,N_10566,N_10569,N_10570,N_10571,N_10572,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10588,N_10589,N_10591,N_10592,N_10593,N_10595,N_10596,N_10597,N_10598,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10607,N_10609,N_10610,N_10611,N_10612,N_10613,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10652,N_10653,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10683,N_10685,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10701,N_10702,N_10704,N_10705,N_10706,N_10708,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10725,N_10726,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10736,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10747,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10791,N_10792,N_10793,N_10795,N_10796,N_10797,N_10799,N_10800,N_10802,N_10803,N_10804,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10813,N_10814,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10844,N_10845,N_10846,N_10848,N_10849,N_10850,N_10851,N_10853,N_10854,N_10855,N_10856,N_10857,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10877,N_10878,N_10879,N_10880,N_10882,N_10883,N_10884,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10904,N_10905,N_10906,N_10909,N_10911,N_10912,N_10913,N_10916,N_10917,N_10918,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10936,N_10938,N_10939,N_10940,N_10945,N_10946,N_10947,N_10949,N_10950,N_10951,N_10952,N_10953,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10963,N_10964,N_10966,N_10967,N_10968,N_10969,N_10970,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11010,N_11011,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11025,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11055,N_11058,N_11059,N_11060,N_11061,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11076,N_11077,N_11078,N_11079,N_11080,N_11082,N_11083,N_11085,N_11086,N_11087,N_11088,N_11090,N_11092,N_11093,N_11094,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11112,N_11113,N_11114,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11124,N_11125,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11134,N_11135,N_11137,N_11138,N_11139,N_11141,N_11142,N_11143,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11156,N_11157,N_11158,N_11159,N_11160,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11170,N_11171,N_11172,N_11174,N_11175,N_11176,N_11177,N_11178,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11188,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11203,N_11204,N_11205,N_11206,N_11209,N_11210,N_11211,N_11212,N_11214,N_11215,N_11216,N_11217,N_11218,N_11221,N_11222,N_11223,N_11224,N_11226,N_11227,N_11228,N_11229,N_11231,N_11232,N_11233,N_11235,N_11236,N_11237,N_11239,N_11240,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11254,N_11255,N_11256,N_11257,N_11258,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11275,N_11278,N_11279,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11289,N_11290,N_11291,N_11292,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11312,N_11315,N_11318,N_11319,N_11320,N_11322,N_11323,N_11325,N_11326,N_11327,N_11329,N_11330,N_11331,N_11332,N_11333,N_11335,N_11338,N_11339,N_11340,N_11342,N_11343,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11353,N_11356,N_11358,N_11359,N_11361,N_11363,N_11364,N_11365,N_11366,N_11367,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11379,N_11380,N_11381,N_11384,N_11385,N_11387,N_11388,N_11389,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11400,N_11401,N_11402,N_11404,N_11405,N_11406,N_11407,N_11408,N_11410,N_11411,N_11412,N_11413,N_11414,N_11416,N_11420,N_11421,N_11422,N_11423,N_11425,N_11426,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11455,N_11456,N_11457,N_11458,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11470,N_11471,N_11472,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11522,N_11523,N_11525,N_11526,N_11527,N_11530,N_11531,N_11533,N_11534,N_11535,N_11536,N_11537,N_11539,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11559,N_11560,N_11561,N_11562,N_11563,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11577,N_11578,N_11579,N_11581,N_11583,N_11584,N_11585,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11598,N_11599,N_11600,N_11601,N_11604,N_11606,N_11607,N_11608,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11629,N_11630,N_11634,N_11635,N_11636,N_11637,N_11638,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11655,N_11656,N_11657,N_11660,N_11662,N_11664,N_11665,N_11667,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11690,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11710,N_11711,N_11712,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11721,N_11723,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11732,N_11734,N_11735,N_11737,N_11738,N_11739,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11749,N_11750,N_11751,N_11753,N_11754,N_11755,N_11756,N_11757,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11768,N_11769,N_11771,N_11772,N_11773,N_11774,N_11775,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11785,N_11787,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11805,N_11807,N_11812,N_11813,N_11814,N_11816,N_11817,N_11818,N_11819,N_11820,N_11823,N_11824,N_11825,N_11828,N_11829,N_11832,N_11833,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11843,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11868,N_11869,N_11870,N_11872,N_11873,N_11874,N_11876,N_11878,N_11879,N_11880,N_11882,N_11883,N_11884,N_11885,N_11886,N_11888,N_11890,N_11891,N_11892,N_11893,N_11894,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11929,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11940,N_11941,N_11944,N_11945,N_11946,N_11949,N_11950,N_11953,N_11954,N_11955,N_11956,N_11957,N_11959,N_11961,N_11962,N_11963,N_11964,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11983,N_11984,N_11985,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11999,N_12000,N_12001,N_12003,N_12004,N_12005,N_12007,N_12008,N_12010,N_12011,N_12012,N_12013,N_12015,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12035,N_12038,N_12039,N_12040,N_12042,N_12043,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12059,N_12060,N_12061,N_12063,N_12064,N_12065,N_12066,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12087,N_12088,N_12089,N_12090,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12103,N_12104,N_12105,N_12106,N_12107,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12128,N_12129,N_12130,N_12131,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12159,N_12160,N_12162,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12172,N_12173,N_12174,N_12177,N_12178,N_12179,N_12180,N_12181,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12220,N_12222,N_12223,N_12224,N_12226,N_12227,N_12229,N_12230,N_12232,N_12235,N_12236,N_12237,N_12238,N_12240,N_12241,N_12242,N_12243,N_12245,N_12246,N_12249,N_12250,N_12251,N_12253,N_12255,N_12257,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12278,N_12279,N_12280,N_12282,N_12283,N_12287,N_12289,N_12290,N_12291,N_12294,N_12296,N_12298,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12308,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12318,N_12319,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12341,N_12342,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12364,N_12365,N_12366,N_12368,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12426,N_12427,N_12428,N_12429,N_12432,N_12433,N_12434,N_12435,N_12436,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12451,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12461,N_12463,N_12464,N_12465,N_12467,N_12468,N_12469,N_12470,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12480,N_12481,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12494,N_12497,N_12498,N_12500,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12531,N_12533,N_12534,N_12535,N_12536,N_12537,N_12540,N_12542,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12554,N_12555,N_12556,N_12557,N_12558,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12586,N_12587,N_12588,N_12590,N_12591,N_12592,N_12595,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12605,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12616,N_12618,N_12619,N_12620,N_12621,N_12622,N_12624,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12637,N_12639,N_12640,N_12641,N_12642,N_12643,N_12645,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12661,N_12662,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12677,N_12678,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12689,N_12690,N_12691,N_12692,N_12693,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12715,N_12717,N_12718,N_12719,N_12720,N_12722,N_12723,N_12724,N_12725,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12740,N_12741,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12751,N_12752,N_12753,N_12754,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12766,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12777,N_12778,N_12779,N_12780,N_12782,N_12783,N_12784,N_12786,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12813,N_12817,N_12818,N_12819,N_12820,N_12821,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12855,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12872,N_12873,N_12874,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12888,N_12889,N_12891,N_12892,N_12893,N_12894,N_12897,N_12898,N_12899,N_12900,N_12901,N_12903,N_12905,N_12908,N_12909,N_12910,N_12911,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12927,N_12928,N_12929,N_12930,N_12933,N_12934,N_12935,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12954,N_12956,N_12958,N_12960,N_12962,N_12964,N_12965,N_12967,N_12969,N_12970,N_12971,N_12973,N_12974,N_12975,N_12978,N_12980,N_12981,N_12982,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12992,N_12993,N_12994,N_12996,N_12997,N_12998,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13010,N_13011,N_13013,N_13014,N_13015,N_13016,N_13017,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13039,N_13040,N_13041,N_13043,N_13044,N_13045,N_13046,N_13048,N_13050,N_13052,N_13053,N_13054,N_13056,N_13058,N_13059,N_13060,N_13062,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13076,N_13077,N_13078,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13093,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13123,N_13124,N_13125,N_13126,N_13128,N_13129,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13142,N_13146,N_13149,N_13150,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13160,N_13161,N_13162,N_13163,N_13166,N_13168,N_13169,N_13170,N_13171,N_13172,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13187,N_13188,N_13189,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13204,N_13205,N_13206,N_13207,N_13208,N_13210,N_13211,N_13212,N_13213,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13224,N_13225,N_13226,N_13227,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13236,N_13237,N_13238,N_13240,N_13241,N_13242,N_13244,N_13245,N_13246,N_13247,N_13248,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13275,N_13276,N_13277,N_13279,N_13281,N_13282,N_13283,N_13285,N_13286,N_13287,N_13289,N_13290,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13299,N_13300,N_13301,N_13302,N_13303,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13312,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13352,N_13353,N_13354,N_13355,N_13357,N_13358,N_13359,N_13361,N_13362,N_13363,N_13364,N_13365,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13375,N_13376,N_13377,N_13378,N_13379,N_13381,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13392,N_13393,N_13394,N_13395,N_13397,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13409,N_13410,N_13411,N_13412,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13431,N_13432,N_13433,N_13434,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13459,N_13461,N_13462,N_13463,N_13465,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13498,N_13499,N_13501,N_13502,N_13503,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13518,N_13519,N_13520,N_13521,N_13523,N_13524,N_13525,N_13526,N_13527,N_13529,N_13530,N_13531,N_13533,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13545,N_13546,N_13547,N_13548,N_13549,N_13551,N_13552,N_13553,N_13554,N_13555,N_13557,N_13558,N_13559,N_13561,N_13562,N_13564,N_13565,N_13567,N_13568,N_13570,N_13571,N_13572,N_13573,N_13575,N_13576,N_13577,N_13578,N_13580,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13600,N_13601,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13615,N_13617,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13626,N_13627,N_13628,N_13629,N_13631,N_13632,N_13633,N_13634,N_13635,N_13637,N_13638,N_13640,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13650,N_13651,N_13652,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13672,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13681,N_13682,N_13683,N_13684,N_13685,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13702,N_13703,N_13704,N_13705,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13716,N_13718,N_13719,N_13720,N_13721,N_13723,N_13724,N_13725,N_13728,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13744,N_13745,N_13747,N_13748,N_13750,N_13751,N_13752,N_13754,N_13756,N_13757,N_13759,N_13760,N_13761,N_13762,N_13764,N_13765,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13778,N_13779,N_13780,N_13782,N_13784,N_13785,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13796,N_13797,N_13798,N_13799,N_13800,N_13802,N_13803,N_13804,N_13805,N_13806,N_13809,N_13810,N_13812,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13821,N_13822,N_13823,N_13825,N_13826,N_13827,N_13829,N_13830,N_13831,N_13832,N_13833,N_13835,N_13836,N_13837,N_13838,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13853,N_13854,N_13855,N_13856,N_13857,N_13859,N_13860,N_13861,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13872,N_13873,N_13875,N_13879,N_13880,N_13881,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13904,N_13906,N_13907,N_13909,N_13910,N_13911,N_13913,N_13916,N_13917,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13935,N_13937,N_13938,N_13939,N_13940,N_13942,N_13943,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13959,N_13960,N_13962,N_13963,N_13964,N_13965,N_13966,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13989,N_13991,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14004,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14017,N_14022,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14032,N_14033,N_14034,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14044,N_14045,N_14046,N_14048,N_14049,N_14050,N_14052,N_14053,N_14055,N_14056,N_14057,N_14058,N_14059,N_14061,N_14062,N_14063,N_14064,N_14065,N_14067,N_14068,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14106,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14117,N_14118,N_14119,N_14120,N_14121,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14132,N_14133,N_14134,N_14135,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14146,N_14147,N_14148,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14157,N_14158,N_14160,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14172,N_14174,N_14175,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14185,N_14186,N_14188,N_14189,N_14190,N_14191,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14219,N_14220,N_14221,N_14223,N_14226,N_14229,N_14230,N_14231,N_14232,N_14234,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14244,N_14245,N_14247,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14257,N_14258,N_14259,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14280,N_14281,N_14282,N_14283,N_14284,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14298,N_14299,N_14302,N_14303,N_14304,N_14306,N_14307,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14321,N_14322,N_14323,N_14324,N_14325,N_14327,N_14328,N_14329,N_14330,N_14331,N_14334,N_14335,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14380,N_14381,N_14384,N_14385,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14412,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14486,N_14487,N_14488,N_14490,N_14491,N_14492,N_14493,N_14494,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14504,N_14505,N_14506,N_14507,N_14509,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14523,N_14524,N_14525,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14536,N_14537,N_14538,N_14539,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14548,N_14549,N_14550,N_14551,N_14554,N_14555,N_14557,N_14558,N_14559,N_14561,N_14562,N_14564,N_14566,N_14567,N_14568,N_14569,N_14571,N_14573,N_14574,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14598,N_14599,N_14601,N_14602,N_14603,N_14606,N_14607,N_14608,N_14609,N_14612,N_14613,N_14614,N_14616,N_14617,N_14618,N_14619,N_14621,N_14623,N_14624,N_14626,N_14627,N_14628,N_14629,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14647,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14661,N_14662,N_14663,N_14664,N_14665,N_14668,N_14669,N_14670,N_14671,N_14672,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14708,N_14709,N_14711,N_14712,N_14713,N_14714,N_14716,N_14717,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14731,N_14733,N_14735,N_14736,N_14737,N_14740,N_14741,N_14743,N_14744,N_14745,N_14746,N_14748,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14776,N_14777,N_14778,N_14781,N_14783,N_14784,N_14785,N_14786,N_14787,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14799,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14828,N_14830,N_14831,N_14832,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14860,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14888,N_14889,N_14890,N_14891,N_14893,N_14894,N_14895,N_14896,N_14898,N_14902,N_14903,N_14904,N_14905,N_14907,N_14908,N_14909,N_14910,N_14911,N_14913,N_14914,N_14915,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14933,N_14934,N_14935,N_14939,N_14940,N_14942,N_14943,N_14944,N_14945,N_14947,N_14948,N_14950,N_14951,N_14953,N_14954,N_14955,N_14956,N_14957,N_14960,N_14961,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14983,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998;
nor U0 (N_0,In_1167,In_522);
xnor U1 (N_1,In_513,In_120);
and U2 (N_2,In_1472,In_955);
nor U3 (N_3,In_1255,In_348);
nand U4 (N_4,In_1334,In_182);
and U5 (N_5,In_1498,In_503);
nor U6 (N_6,In_127,In_99);
nor U7 (N_7,In_740,In_1205);
or U8 (N_8,In_1406,In_536);
and U9 (N_9,In_1471,In_1478);
and U10 (N_10,In_1149,In_710);
or U11 (N_11,In_17,In_628);
and U12 (N_12,In_27,In_92);
and U13 (N_13,In_1147,In_666);
nor U14 (N_14,In_922,In_1151);
or U15 (N_15,In_163,In_546);
xor U16 (N_16,In_688,In_266);
nor U17 (N_17,In_971,In_68);
nor U18 (N_18,In_1320,In_1392);
nand U19 (N_19,In_178,In_586);
or U20 (N_20,In_1459,In_743);
nand U21 (N_21,In_1409,In_129);
and U22 (N_22,In_36,In_515);
or U23 (N_23,In_1068,In_1097);
nor U24 (N_24,In_984,In_772);
nor U25 (N_25,In_78,In_899);
and U26 (N_26,In_359,In_1190);
nor U27 (N_27,In_254,In_1186);
nand U28 (N_28,In_1202,In_470);
and U29 (N_29,In_564,In_638);
or U30 (N_30,In_57,In_237);
xnor U31 (N_31,In_1483,In_953);
and U32 (N_32,In_103,In_623);
nand U33 (N_33,In_1163,In_1364);
nand U34 (N_34,In_1236,In_1142);
or U35 (N_35,In_1239,In_1323);
nor U36 (N_36,In_555,In_770);
and U37 (N_37,In_136,In_818);
and U38 (N_38,In_1177,In_1073);
or U39 (N_39,In_323,In_1494);
and U40 (N_40,In_872,In_862);
nor U41 (N_41,In_833,In_433);
or U42 (N_42,In_1380,In_232);
nor U43 (N_43,In_1252,In_22);
nand U44 (N_44,In_475,In_1160);
or U45 (N_45,In_287,In_1442);
nor U46 (N_46,In_734,In_914);
nor U47 (N_47,In_45,In_1088);
nand U48 (N_48,In_1183,In_1074);
nor U49 (N_49,In_680,In_542);
or U50 (N_50,In_262,In_183);
and U51 (N_51,In_72,In_437);
nor U52 (N_52,In_419,In_428);
or U53 (N_53,In_530,In_873);
xor U54 (N_54,In_1455,In_987);
or U55 (N_55,In_435,In_1187);
nor U56 (N_56,In_1017,In_1340);
and U57 (N_57,In_253,In_297);
nor U58 (N_58,In_844,In_1185);
nor U59 (N_59,In_375,In_1264);
nand U60 (N_60,In_658,In_753);
or U61 (N_61,In_936,In_401);
nor U62 (N_62,In_87,In_979);
nor U63 (N_63,In_440,In_1032);
and U64 (N_64,In_1371,In_74);
xnor U65 (N_65,In_400,In_1369);
or U66 (N_66,In_209,In_1055);
xnor U67 (N_67,In_248,In_134);
nand U68 (N_68,In_0,In_538);
or U69 (N_69,In_1019,In_1121);
nand U70 (N_70,In_1069,In_1287);
or U71 (N_71,In_1404,In_1056);
or U72 (N_72,In_1384,In_620);
nor U73 (N_73,In_1026,In_594);
nand U74 (N_74,In_365,In_1028);
or U75 (N_75,In_100,In_12);
nand U76 (N_76,In_892,In_793);
nand U77 (N_77,In_829,In_723);
and U78 (N_78,In_865,In_289);
nor U79 (N_79,In_1100,In_112);
nor U80 (N_80,In_114,In_630);
and U81 (N_81,In_618,In_337);
or U82 (N_82,In_669,In_343);
nor U83 (N_83,In_33,In_921);
nand U84 (N_84,In_1157,In_1411);
or U85 (N_85,In_77,In_367);
nor U86 (N_86,In_958,In_529);
nor U87 (N_87,In_1221,In_1214);
or U88 (N_88,In_1436,In_644);
xor U89 (N_89,In_215,In_1112);
xor U90 (N_90,In_117,In_1085);
nor U91 (N_91,In_1417,In_1398);
and U92 (N_92,In_1363,In_1253);
xor U93 (N_93,In_60,In_1388);
and U94 (N_94,In_1152,In_205);
nor U95 (N_95,In_1440,In_1022);
and U96 (N_96,In_1269,In_482);
xor U97 (N_97,In_430,In_465);
nand U98 (N_98,In_229,In_251);
nand U99 (N_99,In_523,In_742);
or U100 (N_100,In_1222,In_1424);
and U101 (N_101,In_1219,In_1496);
nand U102 (N_102,In_1378,In_224);
nor U103 (N_103,In_1465,In_131);
xor U104 (N_104,In_764,In_445);
nor U105 (N_105,In_600,In_149);
and U106 (N_106,In_1002,In_654);
nand U107 (N_107,In_826,In_1171);
or U108 (N_108,In_1332,In_30);
nand U109 (N_109,In_53,In_518);
nand U110 (N_110,In_50,In_382);
and U111 (N_111,In_24,In_992);
or U112 (N_112,In_1191,In_1141);
nand U113 (N_113,In_878,In_402);
nor U114 (N_114,In_714,In_115);
or U115 (N_115,In_990,In_1449);
nand U116 (N_116,In_64,In_242);
xnor U117 (N_117,In_1128,In_413);
and U118 (N_118,In_632,In_1107);
nand U119 (N_119,In_1006,In_827);
nand U120 (N_120,In_1244,In_1220);
and U121 (N_121,In_1397,In_369);
or U122 (N_122,In_1053,In_1210);
nor U123 (N_123,In_81,In_212);
xnor U124 (N_124,In_752,In_791);
and U125 (N_125,In_1135,In_496);
xor U126 (N_126,In_962,In_520);
nor U127 (N_127,In_493,In_6);
xor U128 (N_128,In_106,In_1482);
nand U129 (N_129,In_1102,In_1289);
nor U130 (N_130,In_1086,In_1230);
or U131 (N_131,In_436,In_569);
or U132 (N_132,In_142,In_1276);
nor U133 (N_133,In_549,In_611);
nand U134 (N_134,In_1401,In_143);
and U135 (N_135,In_1412,In_1432);
and U136 (N_136,In_606,In_1103);
nor U137 (N_137,In_1217,In_338);
nor U138 (N_138,In_155,In_422);
and U139 (N_139,In_633,In_952);
and U140 (N_140,In_1418,In_788);
and U141 (N_141,In_1415,In_257);
and U142 (N_142,In_874,In_959);
and U143 (N_143,In_656,In_1194);
nor U144 (N_144,In_659,In_901);
or U145 (N_145,In_741,In_1297);
nand U146 (N_146,In_657,In_179);
or U147 (N_147,In_198,In_38);
and U148 (N_148,In_676,In_1036);
nor U149 (N_149,In_755,In_1350);
nand U150 (N_150,In_341,In_1109);
nand U151 (N_151,In_974,In_245);
nor U152 (N_152,In_614,In_394);
and U153 (N_153,In_662,In_1473);
nand U154 (N_154,In_47,In_1093);
nor U155 (N_155,In_146,In_381);
and U156 (N_156,In_1313,In_41);
nor U157 (N_157,In_98,In_1416);
or U158 (N_158,In_746,In_870);
or U159 (N_159,In_647,In_1427);
and U160 (N_160,In_28,In_1360);
nand U161 (N_161,In_769,In_1108);
nand U162 (N_162,In_605,In_565);
xor U163 (N_163,In_466,In_598);
xnor U164 (N_164,In_333,In_780);
nand U165 (N_165,In_383,In_1327);
nand U166 (N_166,In_222,In_977);
or U167 (N_167,In_54,In_1084);
nand U168 (N_168,In_843,In_619);
xor U169 (N_169,In_849,In_84);
and U170 (N_170,In_1296,In_691);
and U171 (N_171,In_227,In_1386);
or U172 (N_172,In_582,In_290);
nor U173 (N_173,In_514,In_532);
xor U174 (N_174,In_1458,In_559);
nand U175 (N_175,In_312,In_983);
nor U176 (N_176,In_882,In_732);
xnor U177 (N_177,In_1265,In_686);
nor U178 (N_178,In_562,In_1037);
nand U179 (N_179,In_1242,In_145);
and U180 (N_180,In_1051,In_181);
and U181 (N_181,In_492,In_5);
and U182 (N_182,In_1329,In_1351);
nor U183 (N_183,In_853,In_889);
nor U184 (N_184,In_761,In_247);
and U185 (N_185,In_1080,In_525);
and U186 (N_186,In_684,In_458);
and U187 (N_187,In_1487,In_1039);
xnor U188 (N_188,In_264,In_331);
or U189 (N_189,In_792,In_560);
or U190 (N_190,In_185,In_840);
or U191 (N_191,In_776,In_403);
or U192 (N_192,In_794,In_1389);
or U193 (N_193,In_351,In_858);
and U194 (N_194,In_697,In_527);
nor U195 (N_195,In_352,In_122);
and U196 (N_196,In_86,In_912);
or U197 (N_197,In_1308,In_167);
and U198 (N_198,In_968,In_1333);
nor U199 (N_199,In_67,In_507);
nor U200 (N_200,In_616,In_576);
and U201 (N_201,In_378,In_276);
or U202 (N_202,In_602,In_293);
or U203 (N_203,In_766,In_411);
or U204 (N_204,In_1326,In_926);
and U205 (N_205,In_1198,In_228);
nor U206 (N_206,In_231,In_377);
nor U207 (N_207,In_720,In_1435);
or U208 (N_208,In_281,In_1305);
nor U209 (N_209,In_808,In_1425);
or U210 (N_210,In_485,In_1035);
or U211 (N_211,In_854,In_226);
and U212 (N_212,In_613,In_510);
and U213 (N_213,In_1270,In_386);
nand U214 (N_214,In_587,In_1481);
or U215 (N_215,In_705,In_762);
nor U216 (N_216,In_1126,In_932);
or U217 (N_217,In_345,In_478);
nor U218 (N_218,In_756,In_144);
and U219 (N_219,In_700,In_497);
or U220 (N_220,In_636,In_828);
xnor U221 (N_221,In_21,In_1490);
or U222 (N_222,In_671,In_151);
nand U223 (N_223,In_220,In_1224);
nor U224 (N_224,In_735,In_250);
and U225 (N_225,In_230,In_685);
nand U226 (N_226,In_1251,In_988);
nor U227 (N_227,In_1321,In_421);
and U228 (N_228,In_767,In_661);
and U229 (N_229,In_781,In_347);
or U230 (N_230,In_306,In_165);
xor U231 (N_231,In_550,In_1492);
or U232 (N_232,In_1235,In_730);
nand U233 (N_233,In_1294,In_573);
nand U234 (N_234,In_213,In_875);
nor U235 (N_235,In_831,In_1311);
xor U236 (N_236,In_1115,In_322);
nor U237 (N_237,In_1447,In_321);
nor U238 (N_238,In_408,In_773);
nand U239 (N_239,In_934,In_1315);
or U240 (N_240,In_123,In_102);
nor U241 (N_241,In_168,In_1402);
nand U242 (N_242,In_1286,In_1009);
and U243 (N_243,In_610,In_881);
xnor U244 (N_244,In_903,In_439);
nand U245 (N_245,In_1422,In_1199);
nor U246 (N_246,In_877,In_1010);
or U247 (N_247,In_689,In_211);
nor U248 (N_248,In_1310,In_1325);
nor U249 (N_249,In_374,In_362);
xor U250 (N_250,In_902,In_32);
and U251 (N_251,In_683,In_850);
or U252 (N_252,In_1113,In_815);
or U253 (N_253,In_687,In_947);
or U254 (N_254,In_1355,In_951);
and U255 (N_255,In_1124,In_911);
nor U256 (N_256,In_907,In_1248);
or U257 (N_257,In_1197,In_868);
nor U258 (N_258,In_82,In_982);
or U259 (N_259,In_1241,In_298);
or U260 (N_260,In_994,In_989);
and U261 (N_261,In_141,In_652);
or U262 (N_262,In_883,In_171);
nor U263 (N_263,In_790,In_137);
nand U264 (N_264,In_1366,In_324);
or U265 (N_265,In_942,In_512);
or U266 (N_266,In_477,In_797);
and U267 (N_267,In_310,In_246);
nand U268 (N_268,In_1451,In_787);
nor U269 (N_269,In_1144,In_52);
or U270 (N_270,In_1292,In_385);
nor U271 (N_271,In_916,In_217);
nand U272 (N_272,In_88,In_291);
nand U273 (N_273,In_414,In_800);
or U274 (N_274,In_1475,In_157);
xor U275 (N_275,In_488,In_370);
nor U276 (N_276,In_534,In_937);
nor U277 (N_277,In_837,In_1277);
nand U278 (N_278,In_501,In_132);
xor U279 (N_279,In_857,In_1118);
and U280 (N_280,In_577,In_929);
nor U281 (N_281,In_380,In_1493);
and U282 (N_282,In_296,In_716);
xor U283 (N_283,In_1405,In_601);
xnor U284 (N_284,In_272,In_682);
nand U285 (N_285,In_1046,In_1083);
nor U286 (N_286,In_1324,In_96);
nand U287 (N_287,In_1182,In_1175);
nor U288 (N_288,In_681,In_806);
or U289 (N_289,In_360,In_1131);
and U290 (N_290,In_1231,In_34);
and U291 (N_291,In_842,In_1279);
and U292 (N_292,In_139,In_471);
nor U293 (N_293,In_646,In_1400);
and U294 (N_294,In_1280,In_1314);
or U295 (N_295,In_830,In_268);
or U296 (N_296,In_1446,In_1489);
nand U297 (N_297,In_271,In_1072);
nor U298 (N_298,In_314,In_452);
and U299 (N_299,In_650,In_1030);
or U300 (N_300,In_739,In_923);
nand U301 (N_301,In_418,In_384);
or U302 (N_302,In_484,In_15);
nor U303 (N_303,In_234,In_480);
xor U304 (N_304,In_1052,In_166);
or U305 (N_305,In_94,In_1331);
nor U306 (N_306,In_1165,In_355);
nor U307 (N_307,In_125,In_591);
or U308 (N_308,In_1013,In_648);
or U309 (N_309,In_938,In_201);
nand U310 (N_310,In_590,In_1345);
nor U311 (N_311,In_282,In_824);
and U312 (N_312,In_1337,In_1419);
and U313 (N_313,In_778,In_1047);
or U314 (N_314,In_540,In_631);
nand U315 (N_315,In_941,In_1385);
and U316 (N_316,In_1353,In_803);
nor U317 (N_317,In_1025,In_107);
and U318 (N_318,In_1448,In_856);
and U319 (N_319,In_7,In_1007);
xor U320 (N_320,In_879,In_554);
nand U321 (N_321,In_93,In_1336);
or U322 (N_322,In_1237,In_670);
and U323 (N_323,In_1259,In_1189);
or U324 (N_324,In_1499,In_1285);
nand U325 (N_325,In_1343,In_1300);
or U326 (N_326,In_1421,In_463);
nor U327 (N_327,In_18,In_285);
nor U328 (N_328,In_29,In_765);
nor U329 (N_329,In_1218,In_13);
or U330 (N_330,In_356,In_1127);
nor U331 (N_331,In_1024,In_1159);
nand U332 (N_332,In_801,In_561);
nand U333 (N_333,In_1257,In_802);
and U334 (N_334,In_195,In_19);
and U335 (N_335,In_785,In_880);
or U336 (N_336,In_986,In_438);
xnor U337 (N_337,In_749,In_1335);
nand U338 (N_338,In_249,In_1299);
nand U339 (N_339,In_197,In_845);
and U340 (N_340,In_69,In_1228);
nor U341 (N_341,In_1161,In_160);
or U342 (N_342,In_387,In_1431);
xor U343 (N_343,In_1322,In_617);
or U344 (N_344,In_733,In_420);
nor U345 (N_345,In_153,In_860);
or U346 (N_346,In_1208,In_404);
nor U347 (N_347,In_1145,In_138);
and U348 (N_348,In_396,In_164);
or U349 (N_349,In_1377,In_395);
or U350 (N_350,In_241,In_1078);
xnor U351 (N_351,In_894,In_442);
and U352 (N_352,In_1207,In_1203);
or U353 (N_353,In_1238,In_1172);
nor U354 (N_354,In_288,In_302);
nand U355 (N_355,In_311,In_431);
nor U356 (N_356,In_187,In_461);
xor U357 (N_357,In_604,In_1023);
or U358 (N_358,In_509,In_1463);
or U359 (N_359,In_1125,In_1129);
and U360 (N_360,In_66,In_583);
nand U361 (N_361,In_1428,In_317);
nor U362 (N_362,In_1266,In_11);
and U363 (N_363,In_1,In_494);
or U364 (N_364,In_1346,In_263);
nor U365 (N_365,In_1021,In_537);
nor U366 (N_366,In_61,In_219);
nor U367 (N_367,In_119,In_548);
nor U368 (N_368,In_1140,In_273);
nor U369 (N_369,In_159,In_1312);
nor U370 (N_370,In_978,In_468);
nor U371 (N_371,In_603,In_118);
or U372 (N_372,In_906,In_855);
nand U373 (N_373,In_90,In_1011);
nor U374 (N_374,In_960,In_1132);
and U375 (N_375,In_319,In_303);
nor U376 (N_376,In_981,In_320);
or U377 (N_377,In_1065,In_233);
and U378 (N_378,In_956,In_286);
nor U379 (N_379,In_128,In_775);
and U380 (N_380,In_1195,In_454);
and U381 (N_381,In_810,In_1354);
or U382 (N_382,In_731,In_1273);
or U383 (N_383,In_747,In_434);
or U384 (N_384,In_1077,In_1200);
nor U385 (N_385,In_1379,In_1034);
and U386 (N_386,In_1031,In_970);
xor U387 (N_387,In_8,In_474);
nand U388 (N_388,In_1291,In_771);
or U389 (N_389,In_909,In_1390);
or U390 (N_390,In_649,In_1133);
and U391 (N_391,In_725,In_10);
nor U392 (N_392,In_895,In_1049);
nor U393 (N_393,In_997,In_1423);
and U394 (N_394,In_235,In_949);
and U395 (N_395,In_698,In_161);
and U396 (N_396,In_244,In_998);
nor U397 (N_397,In_847,In_189);
nand U398 (N_398,In_722,In_736);
and U399 (N_399,In_1461,In_1318);
nand U400 (N_400,In_1123,In_713);
nand U401 (N_401,In_904,In_1048);
or U402 (N_402,In_609,In_1293);
nor U403 (N_403,In_950,In_318);
nand U404 (N_404,In_629,In_653);
and U405 (N_405,In_690,In_972);
or U406 (N_406,In_169,In_920);
xnor U407 (N_407,In_397,In_704);
or U408 (N_408,In_1303,In_531);
nor U409 (N_409,In_500,In_694);
or U410 (N_410,In_1283,In_1272);
nor U411 (N_411,In_332,In_1288);
or U412 (N_412,In_412,In_679);
or U413 (N_413,In_807,In_545);
or U414 (N_414,In_1383,In_1464);
and U415 (N_415,In_1263,In_483);
nand U416 (N_416,In_574,In_1064);
nor U417 (N_417,In_744,In_1096);
xor U418 (N_418,In_677,In_473);
and U419 (N_419,In_964,In_622);
nand U420 (N_420,In_425,In_1136);
nor U421 (N_421,In_31,In_1240);
and U422 (N_422,In_1184,In_63);
xnor U423 (N_423,In_267,In_864);
nor U424 (N_424,In_116,In_763);
or U425 (N_425,In_925,In_366);
nand U426 (N_426,In_1041,In_544);
or U427 (N_427,In_1382,In_643);
xnor U428 (N_428,In_729,In_626);
nand U429 (N_429,In_1268,In_1374);
and U430 (N_430,In_557,In_336);
or U431 (N_431,In_313,In_1066);
and U432 (N_432,In_265,In_274);
nand U433 (N_433,In_1348,In_1001);
or U434 (N_434,In_1196,In_627);
nor U435 (N_435,In_1437,In_1038);
nor U436 (N_436,In_593,In_1284);
nand U437 (N_437,In_1079,In_258);
and U438 (N_438,In_207,In_1488);
nor U439 (N_439,In_176,In_841);
nand U440 (N_440,In_1029,In_567);
nand U441 (N_441,In_1407,In_140);
nand U442 (N_442,In_221,In_1341);
nor U443 (N_443,In_640,In_777);
or U444 (N_444,In_204,In_1243);
nor U445 (N_445,In_1347,In_65);
or U446 (N_446,In_315,In_476);
and U447 (N_447,In_441,In_243);
nor U448 (N_448,In_502,In_696);
nor U449 (N_449,In_718,In_91);
xnor U450 (N_450,In_446,In_935);
nand U451 (N_451,In_641,In_748);
nor U452 (N_452,In_639,In_939);
xor U453 (N_453,In_1148,In_462);
or U454 (N_454,In_651,In_1178);
or U455 (N_455,In_43,In_1356);
and U456 (N_456,In_1063,In_852);
nor U457 (N_457,In_1414,In_457);
nor U458 (N_458,In_1062,In_1122);
and U459 (N_459,In_79,In_812);
and U460 (N_460,In_1391,In_1155);
and U461 (N_461,In_612,In_552);
or U462 (N_462,In_692,In_238);
nor U463 (N_463,In_240,In_721);
or U464 (N_464,In_1176,In_876);
and U465 (N_465,In_702,In_751);
xnor U466 (N_466,In_1054,In_1316);
nor U467 (N_467,In_933,In_1164);
nor U468 (N_468,In_239,In_719);
or U469 (N_469,In_379,In_162);
nor U470 (N_470,In_521,In_121);
and U471 (N_471,In_505,In_58);
or U472 (N_472,In_592,In_449);
nand U473 (N_473,In_760,In_177);
nor U474 (N_474,In_985,In_615);
nor U475 (N_475,In_40,In_727);
xnor U476 (N_476,In_105,In_202);
xnor U477 (N_477,In_961,In_832);
and U478 (N_478,In_194,In_568);
and U479 (N_479,In_173,In_539);
nor U480 (N_480,In_1469,In_342);
or U481 (N_481,In_861,In_796);
or U482 (N_482,In_1206,In_1370);
nand U483 (N_483,In_758,In_426);
nor U484 (N_484,In_275,In_1486);
nand U485 (N_485,In_135,In_417);
or U486 (N_486,In_415,In_675);
nor U487 (N_487,In_1480,In_1376);
and U488 (N_488,In_823,In_1095);
nand U489 (N_489,In_1452,In_456);
and U490 (N_490,In_642,In_711);
and U491 (N_491,In_1367,In_750);
nand U492 (N_492,In_1439,In_1004);
or U493 (N_493,In_1470,In_1005);
nand U494 (N_494,In_1250,In_1174);
and U495 (N_495,In_472,In_2);
or U496 (N_496,In_784,In_388);
or U497 (N_497,In_300,In_1227);
and U498 (N_498,In_851,In_1247);
nor U499 (N_499,In_1201,In_811);
nor U500 (N_500,In_890,In_1014);
nor U501 (N_501,In_821,In_1012);
nor U502 (N_502,In_506,In_1089);
nand U503 (N_503,In_451,In_133);
nor U504 (N_504,In_1290,In_225);
nor U505 (N_505,In_1000,In_1139);
nor U506 (N_506,In_1245,In_634);
and U507 (N_507,In_393,In_124);
or U508 (N_508,In_1111,In_795);
or U509 (N_509,In_364,In_1162);
xnor U510 (N_510,In_1495,In_208);
nor U511 (N_511,In_464,In_175);
and U512 (N_512,In_193,In_867);
nor U513 (N_513,In_871,In_1426);
nor U514 (N_514,In_1258,In_528);
and U515 (N_515,In_672,In_976);
nand U516 (N_516,In_1213,In_1403);
xnor U517 (N_517,In_1420,In_1075);
nand U518 (N_518,In_835,In_23);
or U519 (N_519,In_915,In_918);
nor U520 (N_520,In_919,In_190);
and U521 (N_521,In_834,In_101);
nand U522 (N_522,In_252,In_301);
nor U523 (N_523,In_1092,In_432);
or U524 (N_524,In_305,In_328);
or U525 (N_525,In_1295,In_1408);
nand U526 (N_526,In_1223,In_910);
xnor U527 (N_527,In_717,In_665);
nand U528 (N_528,In_89,In_368);
or U529 (N_529,In_1209,In_511);
or U530 (N_530,In_200,In_664);
or U531 (N_531,In_97,In_1429);
nor U532 (N_532,In_1352,In_798);
nand U533 (N_533,In_1395,In_1262);
nor U534 (N_534,In_55,In_754);
nand U535 (N_535,In_1307,In_1044);
xnor U536 (N_536,In_1444,In_1061);
nand U537 (N_537,In_1330,In_104);
nand U538 (N_538,In_695,In_16);
and U539 (N_539,In_9,In_498);
or U540 (N_540,In_353,In_490);
or U541 (N_541,In_398,In_1170);
or U542 (N_542,In_1474,In_126);
nand U543 (N_543,In_354,In_900);
xor U544 (N_544,In_269,In_579);
nand U545 (N_545,In_526,In_1274);
nor U546 (N_546,In_1154,In_846);
and U547 (N_547,In_152,In_1460);
or U548 (N_548,In_578,In_148);
nor U549 (N_549,In_261,In_973);
or U550 (N_550,In_358,In_391);
or U551 (N_551,In_980,In_817);
nand U552 (N_552,In_1137,In_330);
nor U553 (N_553,In_1339,In_1317);
nor U554 (N_554,In_673,In_668);
nand U555 (N_555,In_156,In_95);
or U556 (N_556,In_56,In_1090);
nand U557 (N_557,In_405,In_635);
nor U558 (N_558,In_809,In_556);
or U559 (N_559,In_693,In_1443);
nor U560 (N_560,In_150,In_885);
and U561 (N_561,In_524,In_931);
or U562 (N_562,In_307,In_996);
nor U563 (N_563,In_308,In_995);
nand U564 (N_564,In_1042,In_42);
or U565 (N_565,In_1180,In_663);
nand U566 (N_566,In_1119,In_350);
or U567 (N_567,In_825,In_667);
nand U568 (N_568,In_469,In_39);
xor U569 (N_569,In_1143,In_715);
and U570 (N_570,In_898,In_1267);
nor U571 (N_571,In_255,In_327);
or U572 (N_572,In_196,In_1484);
nor U573 (N_573,In_930,In_940);
and U574 (N_574,In_999,In_637);
nor U575 (N_575,In_1491,In_399);
xnor U576 (N_576,In_905,In_887);
nor U577 (N_577,In_349,In_1116);
nand U578 (N_578,In_814,In_280);
nor U579 (N_579,In_1438,In_563);
nand U580 (N_580,In_85,In_597);
nor U581 (N_581,In_35,In_75);
nor U582 (N_582,In_423,In_1076);
nor U583 (N_583,In_1045,In_479);
nor U584 (N_584,In_884,In_25);
or U585 (N_585,In_216,In_575);
or U586 (N_586,In_1226,In_499);
xor U587 (N_587,In_299,In_1454);
or U588 (N_588,In_80,In_708);
xor U589 (N_589,In_460,In_1302);
or U590 (N_590,In_816,In_1156);
or U591 (N_591,In_1058,In_113);
or U592 (N_592,In_838,In_203);
or U593 (N_593,In_924,In_14);
nand U594 (N_594,In_481,In_1158);
nand U595 (N_595,In_1104,In_295);
nor U596 (N_596,In_111,In_1479);
nor U597 (N_597,In_709,In_789);
or U598 (N_598,In_1188,In_158);
nand U599 (N_599,In_184,In_1453);
and U600 (N_600,In_572,In_256);
nand U601 (N_601,In_533,In_535);
and U602 (N_602,In_453,In_707);
xnor U603 (N_603,In_893,In_599);
and U604 (N_604,In_822,In_1192);
xnor U605 (N_605,In_975,In_1365);
nor U606 (N_606,In_1138,In_1173);
nor U607 (N_607,In_839,In_489);
xnor U608 (N_608,In_813,In_83);
or U609 (N_609,In_3,In_712);
or U610 (N_610,In_76,In_1134);
xor U611 (N_611,In_206,In_1033);
or U612 (N_612,In_588,In_191);
and U613 (N_613,In_109,In_585);
or U614 (N_614,In_674,In_277);
xor U615 (N_615,In_409,In_1070);
or U616 (N_616,In_48,In_1057);
nand U617 (N_617,In_154,In_1357);
and U618 (N_618,In_1396,In_1497);
nor U619 (N_619,In_897,In_260);
nor U620 (N_620,In_147,In_786);
and U621 (N_621,In_223,In_1169);
and U622 (N_622,In_1358,In_779);
nor U623 (N_623,In_1101,In_566);
or U624 (N_624,In_73,In_1462);
nand U625 (N_625,In_495,In_607);
or U626 (N_626,In_1445,In_1067);
nand U627 (N_627,In_745,In_410);
and U628 (N_628,In_270,In_1094);
nor U629 (N_629,In_655,In_963);
nand U630 (N_630,In_455,In_737);
and U631 (N_631,In_782,In_913);
or U632 (N_632,In_467,In_1399);
nand U633 (N_633,In_1372,In_1309);
nor U634 (N_634,In_424,In_863);
or U635 (N_635,In_703,In_1168);
nand U636 (N_636,In_660,In_284);
and U637 (N_637,In_1215,In_1081);
and U638 (N_638,In_236,In_1015);
nand U639 (N_639,In_1016,In_199);
and U640 (N_640,In_1328,In_279);
nor U641 (N_641,In_896,In_1359);
xnor U642 (N_642,In_108,In_1304);
and U643 (N_643,In_966,In_1110);
or U644 (N_644,In_1232,In_1071);
or U645 (N_645,In_407,In_20);
or U646 (N_646,In_888,In_450);
nor U647 (N_647,In_581,In_1485);
or U648 (N_648,In_1020,In_1393);
nor U649 (N_649,In_820,In_625);
and U650 (N_650,In_1433,In_768);
or U651 (N_651,In_1368,In_1059);
and U652 (N_652,In_1468,In_944);
and U653 (N_653,In_596,In_429);
nor U654 (N_654,In_361,In_357);
nor U655 (N_655,In_621,In_180);
and U656 (N_656,In_1099,In_701);
nor U657 (N_657,In_1301,In_948);
nand U658 (N_658,In_1003,In_416);
or U659 (N_659,In_1413,In_993);
nand U660 (N_660,In_508,In_1179);
nand U661 (N_661,In_943,In_325);
or U662 (N_662,In_848,In_558);
nand U663 (N_663,In_1150,In_1216);
or U664 (N_664,In_1234,In_427);
xnor U665 (N_665,In_957,In_51);
and U666 (N_666,In_71,In_340);
nand U667 (N_667,In_294,In_759);
xor U668 (N_668,In_62,In_392);
nor U669 (N_669,In_1260,In_1450);
nor U670 (N_670,In_580,In_70);
nor U671 (N_671,In_459,In_1278);
or U672 (N_672,In_1256,In_1275);
or U673 (N_673,In_170,In_59);
or U674 (N_674,In_946,In_491);
and U675 (N_675,In_869,In_836);
nor U676 (N_676,In_1430,In_886);
or U677 (N_677,In_44,In_965);
nor U678 (N_678,In_945,In_1193);
xor U679 (N_679,In_344,In_1466);
nor U680 (N_680,In_645,In_799);
nand U681 (N_681,In_504,In_309);
nand U682 (N_682,In_1282,In_1212);
or U683 (N_683,In_346,In_726);
or U684 (N_684,In_1467,In_541);
nand U685 (N_685,In_130,In_1027);
and U686 (N_686,In_1233,In_624);
nor U687 (N_687,In_1211,In_372);
and U688 (N_688,In_678,In_1306);
or U689 (N_689,In_292,In_1060);
nand U690 (N_690,In_486,In_1338);
xnor U691 (N_691,In_805,In_174);
and U692 (N_692,In_991,In_1298);
nand U693 (N_693,In_46,In_1114);
and U694 (N_694,In_571,In_214);
and U695 (N_695,In_371,In_283);
nor U696 (N_696,In_1040,In_738);
nand U697 (N_697,In_1106,In_259);
nand U698 (N_698,In_1456,In_570);
nor U699 (N_699,In_335,In_516);
nand U700 (N_700,In_804,In_774);
nand U701 (N_701,In_584,In_1477);
nand U702 (N_702,In_595,In_1130);
xor U703 (N_703,In_373,In_706);
or U704 (N_704,In_859,In_543);
xor U705 (N_705,In_547,In_1342);
xnor U706 (N_706,In_1225,In_1476);
nor U707 (N_707,In_1387,In_1181);
nor U708 (N_708,In_908,In_1381);
and U709 (N_709,In_699,In_917);
and U710 (N_710,In_1410,In_1153);
nand U711 (N_711,In_928,In_1457);
nand U712 (N_712,In_49,In_1434);
or U713 (N_713,In_443,In_1246);
nor U714 (N_714,In_1043,In_188);
and U715 (N_715,In_1098,In_1050);
nor U716 (N_716,In_954,In_1249);
and U717 (N_717,In_447,In_1361);
nor U718 (N_718,In_1018,In_1344);
nand U719 (N_719,In_927,In_1008);
or U720 (N_720,In_1254,In_551);
or U721 (N_721,In_376,In_866);
and U722 (N_722,In_757,In_1441);
or U723 (N_723,In_218,In_728);
and U724 (N_724,In_278,In_608);
xnor U725 (N_725,In_406,In_553);
and U726 (N_726,In_37,In_1394);
and U727 (N_727,In_110,In_487);
nor U728 (N_728,In_1166,In_819);
and U729 (N_729,In_1375,In_1362);
and U730 (N_730,In_1229,In_1117);
xnor U731 (N_731,In_967,In_326);
nor U732 (N_732,In_334,In_1087);
or U733 (N_733,In_363,In_589);
and U734 (N_734,In_783,In_192);
nand U735 (N_735,In_969,In_186);
xor U736 (N_736,In_1271,In_389);
or U737 (N_737,In_1281,In_1204);
and U738 (N_738,In_1146,In_519);
and U739 (N_739,In_172,In_26);
and U740 (N_740,In_304,In_448);
or U741 (N_741,In_316,In_1373);
or U742 (N_742,In_1105,In_891);
nand U743 (N_743,In_724,In_390);
xnor U744 (N_744,In_210,In_1261);
nand U745 (N_745,In_517,In_1120);
nand U746 (N_746,In_329,In_1091);
nor U747 (N_747,In_339,In_1082);
or U748 (N_748,In_444,In_4);
nor U749 (N_749,In_1349,In_1319);
nand U750 (N_750,In_995,In_526);
nand U751 (N_751,In_907,In_1126);
and U752 (N_752,In_39,In_1149);
or U753 (N_753,In_668,In_1147);
or U754 (N_754,In_561,In_142);
nand U755 (N_755,In_73,In_1082);
or U756 (N_756,In_338,In_1307);
or U757 (N_757,In_964,In_1031);
or U758 (N_758,In_885,In_1183);
nor U759 (N_759,In_1399,In_146);
xnor U760 (N_760,In_1042,In_1269);
nand U761 (N_761,In_331,In_919);
nand U762 (N_762,In_996,In_312);
nand U763 (N_763,In_938,In_544);
and U764 (N_764,In_763,In_1456);
xnor U765 (N_765,In_1457,In_479);
and U766 (N_766,In_27,In_876);
nor U767 (N_767,In_654,In_233);
or U768 (N_768,In_1211,In_732);
and U769 (N_769,In_1402,In_1242);
nor U770 (N_770,In_464,In_138);
or U771 (N_771,In_624,In_625);
nor U772 (N_772,In_2,In_1019);
nor U773 (N_773,In_39,In_1132);
xnor U774 (N_774,In_599,In_1425);
nand U775 (N_775,In_1112,In_270);
nand U776 (N_776,In_1026,In_105);
or U777 (N_777,In_221,In_862);
and U778 (N_778,In_997,In_1230);
nand U779 (N_779,In_1000,In_923);
or U780 (N_780,In_1083,In_1299);
nor U781 (N_781,In_1456,In_50);
nor U782 (N_782,In_611,In_678);
nand U783 (N_783,In_383,In_507);
xnor U784 (N_784,In_1299,In_801);
and U785 (N_785,In_678,In_133);
xor U786 (N_786,In_865,In_742);
nand U787 (N_787,In_693,In_902);
or U788 (N_788,In_1266,In_1247);
or U789 (N_789,In_196,In_867);
or U790 (N_790,In_1174,In_302);
nor U791 (N_791,In_126,In_267);
nor U792 (N_792,In_157,In_544);
or U793 (N_793,In_1460,In_261);
xor U794 (N_794,In_1070,In_1403);
xnor U795 (N_795,In_831,In_457);
nand U796 (N_796,In_113,In_1264);
and U797 (N_797,In_663,In_557);
and U798 (N_798,In_1285,In_391);
and U799 (N_799,In_257,In_221);
or U800 (N_800,In_103,In_647);
nor U801 (N_801,In_494,In_1049);
and U802 (N_802,In_90,In_575);
or U803 (N_803,In_490,In_522);
nor U804 (N_804,In_514,In_1031);
or U805 (N_805,In_705,In_340);
or U806 (N_806,In_917,In_1377);
and U807 (N_807,In_1087,In_468);
and U808 (N_808,In_613,In_1047);
nor U809 (N_809,In_123,In_11);
nand U810 (N_810,In_244,In_79);
and U811 (N_811,In_890,In_301);
nand U812 (N_812,In_834,In_866);
nor U813 (N_813,In_318,In_979);
nand U814 (N_814,In_169,In_1260);
nor U815 (N_815,In_429,In_564);
xnor U816 (N_816,In_846,In_912);
or U817 (N_817,In_1091,In_972);
or U818 (N_818,In_617,In_1291);
or U819 (N_819,In_537,In_44);
and U820 (N_820,In_1223,In_1181);
xor U821 (N_821,In_919,In_431);
and U822 (N_822,In_632,In_1408);
nor U823 (N_823,In_1393,In_744);
or U824 (N_824,In_1128,In_1238);
and U825 (N_825,In_933,In_1492);
nand U826 (N_826,In_1224,In_1404);
nand U827 (N_827,In_555,In_598);
nor U828 (N_828,In_472,In_618);
or U829 (N_829,In_548,In_1448);
xor U830 (N_830,In_465,In_1182);
nor U831 (N_831,In_129,In_453);
or U832 (N_832,In_1342,In_825);
nand U833 (N_833,In_1375,In_61);
nor U834 (N_834,In_1260,In_1453);
nor U835 (N_835,In_255,In_1205);
nor U836 (N_836,In_414,In_106);
nand U837 (N_837,In_450,In_312);
and U838 (N_838,In_1013,In_663);
nand U839 (N_839,In_1004,In_17);
nand U840 (N_840,In_262,In_32);
nor U841 (N_841,In_1288,In_443);
nor U842 (N_842,In_61,In_303);
and U843 (N_843,In_1363,In_296);
nor U844 (N_844,In_388,In_742);
nor U845 (N_845,In_629,In_656);
nand U846 (N_846,In_205,In_660);
nor U847 (N_847,In_969,In_324);
and U848 (N_848,In_1318,In_577);
nand U849 (N_849,In_107,In_94);
nor U850 (N_850,In_854,In_751);
nand U851 (N_851,In_957,In_932);
nor U852 (N_852,In_1466,In_466);
xnor U853 (N_853,In_566,In_1453);
nand U854 (N_854,In_1491,In_1140);
xnor U855 (N_855,In_1448,In_565);
and U856 (N_856,In_689,In_387);
and U857 (N_857,In_893,In_457);
xor U858 (N_858,In_1225,In_215);
and U859 (N_859,In_632,In_1099);
or U860 (N_860,In_1144,In_248);
and U861 (N_861,In_836,In_1116);
or U862 (N_862,In_343,In_1372);
or U863 (N_863,In_600,In_777);
or U864 (N_864,In_541,In_705);
nand U865 (N_865,In_1024,In_527);
or U866 (N_866,In_669,In_58);
nand U867 (N_867,In_1417,In_1333);
or U868 (N_868,In_865,In_1112);
nor U869 (N_869,In_1380,In_1143);
and U870 (N_870,In_555,In_448);
and U871 (N_871,In_246,In_11);
nor U872 (N_872,In_1357,In_67);
nor U873 (N_873,In_696,In_1238);
nor U874 (N_874,In_349,In_1296);
nand U875 (N_875,In_1498,In_974);
nand U876 (N_876,In_696,In_865);
nand U877 (N_877,In_941,In_1466);
nand U878 (N_878,In_768,In_1393);
and U879 (N_879,In_513,In_768);
or U880 (N_880,In_1421,In_876);
and U881 (N_881,In_133,In_1452);
nor U882 (N_882,In_1095,In_1438);
nor U883 (N_883,In_426,In_573);
nand U884 (N_884,In_1349,In_1279);
nor U885 (N_885,In_1,In_1325);
nand U886 (N_886,In_643,In_943);
nand U887 (N_887,In_867,In_622);
and U888 (N_888,In_1321,In_69);
xor U889 (N_889,In_352,In_1182);
or U890 (N_890,In_1481,In_829);
xnor U891 (N_891,In_393,In_961);
nand U892 (N_892,In_1157,In_1041);
and U893 (N_893,In_235,In_152);
xnor U894 (N_894,In_13,In_154);
or U895 (N_895,In_648,In_247);
xnor U896 (N_896,In_494,In_660);
or U897 (N_897,In_1443,In_705);
and U898 (N_898,In_80,In_1157);
or U899 (N_899,In_1393,In_1190);
and U900 (N_900,In_112,In_750);
or U901 (N_901,In_994,In_978);
nor U902 (N_902,In_1010,In_1139);
or U903 (N_903,In_745,In_239);
or U904 (N_904,In_213,In_1433);
nor U905 (N_905,In_903,In_271);
nand U906 (N_906,In_798,In_1415);
xor U907 (N_907,In_364,In_1247);
or U908 (N_908,In_333,In_625);
xor U909 (N_909,In_821,In_1271);
nand U910 (N_910,In_42,In_650);
nand U911 (N_911,In_699,In_1235);
nor U912 (N_912,In_447,In_804);
and U913 (N_913,In_5,In_1250);
and U914 (N_914,In_1351,In_911);
or U915 (N_915,In_917,In_1049);
nor U916 (N_916,In_157,In_436);
or U917 (N_917,In_267,In_1480);
and U918 (N_918,In_23,In_26);
nor U919 (N_919,In_798,In_1209);
and U920 (N_920,In_958,In_584);
or U921 (N_921,In_897,In_59);
nor U922 (N_922,In_363,In_174);
nor U923 (N_923,In_1487,In_1011);
and U924 (N_924,In_276,In_841);
or U925 (N_925,In_828,In_300);
or U926 (N_926,In_532,In_1284);
nor U927 (N_927,In_1471,In_1041);
nand U928 (N_928,In_58,In_736);
and U929 (N_929,In_1000,In_1092);
and U930 (N_930,In_884,In_576);
and U931 (N_931,In_395,In_1273);
nand U932 (N_932,In_437,In_633);
nand U933 (N_933,In_118,In_584);
nor U934 (N_934,In_392,In_1068);
and U935 (N_935,In_337,In_387);
nand U936 (N_936,In_498,In_540);
nand U937 (N_937,In_725,In_281);
nand U938 (N_938,In_464,In_249);
xnor U939 (N_939,In_682,In_983);
nand U940 (N_940,In_173,In_147);
and U941 (N_941,In_456,In_444);
and U942 (N_942,In_737,In_482);
nand U943 (N_943,In_302,In_562);
and U944 (N_944,In_395,In_330);
and U945 (N_945,In_1045,In_1264);
nor U946 (N_946,In_331,In_1135);
or U947 (N_947,In_461,In_118);
nor U948 (N_948,In_241,In_252);
and U949 (N_949,In_852,In_1217);
nand U950 (N_950,In_912,In_709);
xnor U951 (N_951,In_693,In_237);
and U952 (N_952,In_723,In_173);
nor U953 (N_953,In_1127,In_539);
and U954 (N_954,In_475,In_944);
and U955 (N_955,In_310,In_1215);
nor U956 (N_956,In_811,In_1361);
or U957 (N_957,In_142,In_1085);
or U958 (N_958,In_1050,In_1184);
and U959 (N_959,In_421,In_56);
nor U960 (N_960,In_996,In_159);
and U961 (N_961,In_54,In_28);
nand U962 (N_962,In_1350,In_480);
or U963 (N_963,In_280,In_7);
nor U964 (N_964,In_604,In_492);
and U965 (N_965,In_126,In_343);
xor U966 (N_966,In_899,In_893);
nor U967 (N_967,In_1064,In_5);
nand U968 (N_968,In_28,In_767);
nor U969 (N_969,In_822,In_1014);
or U970 (N_970,In_1190,In_896);
and U971 (N_971,In_543,In_254);
and U972 (N_972,In_638,In_295);
and U973 (N_973,In_1451,In_1364);
and U974 (N_974,In_424,In_391);
nor U975 (N_975,In_20,In_1048);
xnor U976 (N_976,In_1292,In_730);
nand U977 (N_977,In_181,In_1173);
or U978 (N_978,In_482,In_127);
or U979 (N_979,In_581,In_941);
nor U980 (N_980,In_1056,In_583);
xor U981 (N_981,In_337,In_653);
and U982 (N_982,In_1066,In_73);
and U983 (N_983,In_1401,In_47);
and U984 (N_984,In_761,In_756);
and U985 (N_985,In_1067,In_634);
xor U986 (N_986,In_1431,In_1151);
nor U987 (N_987,In_361,In_545);
and U988 (N_988,In_1037,In_147);
and U989 (N_989,In_351,In_834);
nor U990 (N_990,In_1161,In_1012);
nor U991 (N_991,In_1083,In_570);
or U992 (N_992,In_161,In_902);
nor U993 (N_993,In_1298,In_738);
nor U994 (N_994,In_299,In_547);
or U995 (N_995,In_455,In_597);
nand U996 (N_996,In_185,In_697);
and U997 (N_997,In_180,In_208);
and U998 (N_998,In_1088,In_489);
or U999 (N_999,In_1182,In_602);
nand U1000 (N_1000,In_254,In_443);
xnor U1001 (N_1001,In_1257,In_19);
xor U1002 (N_1002,In_1052,In_1064);
or U1003 (N_1003,In_1480,In_1145);
or U1004 (N_1004,In_201,In_1385);
and U1005 (N_1005,In_904,In_1446);
or U1006 (N_1006,In_574,In_1223);
nand U1007 (N_1007,In_399,In_1132);
nand U1008 (N_1008,In_925,In_268);
nor U1009 (N_1009,In_27,In_1380);
nor U1010 (N_1010,In_118,In_327);
or U1011 (N_1011,In_379,In_4);
or U1012 (N_1012,In_275,In_1122);
nand U1013 (N_1013,In_1070,In_373);
and U1014 (N_1014,In_317,In_22);
and U1015 (N_1015,In_1221,In_336);
and U1016 (N_1016,In_1259,In_988);
and U1017 (N_1017,In_0,In_638);
and U1018 (N_1018,In_209,In_872);
or U1019 (N_1019,In_997,In_1105);
nand U1020 (N_1020,In_1339,In_1272);
and U1021 (N_1021,In_731,In_388);
or U1022 (N_1022,In_564,In_696);
or U1023 (N_1023,In_347,In_284);
or U1024 (N_1024,In_325,In_937);
and U1025 (N_1025,In_271,In_1195);
nand U1026 (N_1026,In_554,In_942);
and U1027 (N_1027,In_824,In_1082);
nand U1028 (N_1028,In_1361,In_1217);
or U1029 (N_1029,In_188,In_962);
xnor U1030 (N_1030,In_604,In_908);
or U1031 (N_1031,In_1252,In_637);
or U1032 (N_1032,In_146,In_56);
nor U1033 (N_1033,In_1045,In_944);
xor U1034 (N_1034,In_201,In_126);
and U1035 (N_1035,In_1404,In_154);
or U1036 (N_1036,In_758,In_328);
xnor U1037 (N_1037,In_741,In_1184);
or U1038 (N_1038,In_644,In_157);
nor U1039 (N_1039,In_168,In_799);
nor U1040 (N_1040,In_215,In_1021);
or U1041 (N_1041,In_392,In_1395);
nor U1042 (N_1042,In_825,In_765);
nor U1043 (N_1043,In_996,In_411);
or U1044 (N_1044,In_485,In_652);
nor U1045 (N_1045,In_679,In_550);
nor U1046 (N_1046,In_1310,In_423);
nor U1047 (N_1047,In_950,In_1220);
and U1048 (N_1048,In_464,In_93);
and U1049 (N_1049,In_453,In_30);
nand U1050 (N_1050,In_1242,In_437);
nor U1051 (N_1051,In_1193,In_1479);
and U1052 (N_1052,In_682,In_1241);
and U1053 (N_1053,In_611,In_1070);
nor U1054 (N_1054,In_1383,In_257);
nor U1055 (N_1055,In_940,In_1288);
and U1056 (N_1056,In_565,In_337);
or U1057 (N_1057,In_1006,In_576);
nor U1058 (N_1058,In_1464,In_8);
nor U1059 (N_1059,In_1083,In_135);
nor U1060 (N_1060,In_985,In_207);
nand U1061 (N_1061,In_718,In_289);
nand U1062 (N_1062,In_4,In_621);
nor U1063 (N_1063,In_1030,In_1278);
nor U1064 (N_1064,In_614,In_992);
nand U1065 (N_1065,In_985,In_1398);
nor U1066 (N_1066,In_1227,In_898);
nand U1067 (N_1067,In_1097,In_1154);
or U1068 (N_1068,In_761,In_1078);
nand U1069 (N_1069,In_1449,In_1127);
nor U1070 (N_1070,In_1401,In_1319);
nand U1071 (N_1071,In_643,In_1137);
and U1072 (N_1072,In_988,In_529);
nand U1073 (N_1073,In_1018,In_1015);
xor U1074 (N_1074,In_643,In_601);
and U1075 (N_1075,In_289,In_1481);
nand U1076 (N_1076,In_1271,In_555);
or U1077 (N_1077,In_868,In_503);
and U1078 (N_1078,In_259,In_663);
or U1079 (N_1079,In_1104,In_711);
nor U1080 (N_1080,In_31,In_1302);
nor U1081 (N_1081,In_1129,In_539);
xnor U1082 (N_1082,In_1281,In_1425);
nand U1083 (N_1083,In_457,In_1238);
nand U1084 (N_1084,In_294,In_116);
or U1085 (N_1085,In_1202,In_85);
or U1086 (N_1086,In_1135,In_285);
or U1087 (N_1087,In_99,In_1247);
nor U1088 (N_1088,In_752,In_130);
nand U1089 (N_1089,In_475,In_129);
nand U1090 (N_1090,In_384,In_1201);
or U1091 (N_1091,In_125,In_85);
nor U1092 (N_1092,In_823,In_805);
and U1093 (N_1093,In_1178,In_1276);
and U1094 (N_1094,In_945,In_758);
and U1095 (N_1095,In_627,In_189);
nand U1096 (N_1096,In_825,In_1103);
nor U1097 (N_1097,In_1358,In_796);
xor U1098 (N_1098,In_1208,In_208);
nand U1099 (N_1099,In_286,In_631);
or U1100 (N_1100,In_1453,In_271);
nor U1101 (N_1101,In_421,In_315);
nor U1102 (N_1102,In_1491,In_1114);
nor U1103 (N_1103,In_596,In_215);
and U1104 (N_1104,In_700,In_989);
nand U1105 (N_1105,In_35,In_592);
nand U1106 (N_1106,In_143,In_665);
or U1107 (N_1107,In_1340,In_527);
and U1108 (N_1108,In_697,In_119);
and U1109 (N_1109,In_694,In_883);
nand U1110 (N_1110,In_860,In_1316);
and U1111 (N_1111,In_1322,In_676);
and U1112 (N_1112,In_1136,In_705);
or U1113 (N_1113,In_327,In_1133);
or U1114 (N_1114,In_1174,In_823);
or U1115 (N_1115,In_1196,In_1393);
nand U1116 (N_1116,In_1489,In_52);
nor U1117 (N_1117,In_173,In_1193);
nor U1118 (N_1118,In_585,In_637);
nor U1119 (N_1119,In_198,In_520);
nor U1120 (N_1120,In_964,In_721);
nand U1121 (N_1121,In_731,In_732);
xor U1122 (N_1122,In_318,In_1145);
nand U1123 (N_1123,In_1041,In_696);
nor U1124 (N_1124,In_1065,In_1158);
or U1125 (N_1125,In_348,In_528);
and U1126 (N_1126,In_867,In_1370);
and U1127 (N_1127,In_586,In_1443);
or U1128 (N_1128,In_990,In_887);
xnor U1129 (N_1129,In_379,In_1269);
nand U1130 (N_1130,In_1246,In_813);
and U1131 (N_1131,In_187,In_202);
nor U1132 (N_1132,In_1282,In_976);
nor U1133 (N_1133,In_296,In_527);
nand U1134 (N_1134,In_1215,In_1379);
nand U1135 (N_1135,In_499,In_874);
nor U1136 (N_1136,In_615,In_1141);
xnor U1137 (N_1137,In_389,In_917);
or U1138 (N_1138,In_861,In_1417);
and U1139 (N_1139,In_592,In_1063);
nor U1140 (N_1140,In_320,In_143);
and U1141 (N_1141,In_620,In_1050);
nand U1142 (N_1142,In_307,In_1188);
and U1143 (N_1143,In_285,In_333);
nand U1144 (N_1144,In_196,In_424);
and U1145 (N_1145,In_1416,In_1109);
nand U1146 (N_1146,In_624,In_60);
and U1147 (N_1147,In_455,In_477);
and U1148 (N_1148,In_650,In_762);
or U1149 (N_1149,In_798,In_1306);
nor U1150 (N_1150,In_697,In_0);
nor U1151 (N_1151,In_625,In_150);
nand U1152 (N_1152,In_1461,In_230);
nor U1153 (N_1153,In_1066,In_1195);
or U1154 (N_1154,In_1459,In_908);
nor U1155 (N_1155,In_914,In_875);
or U1156 (N_1156,In_1493,In_276);
and U1157 (N_1157,In_1186,In_265);
nor U1158 (N_1158,In_1407,In_1346);
or U1159 (N_1159,In_668,In_622);
and U1160 (N_1160,In_1075,In_265);
nor U1161 (N_1161,In_1352,In_1122);
nor U1162 (N_1162,In_1421,In_733);
and U1163 (N_1163,In_1365,In_600);
or U1164 (N_1164,In_466,In_336);
and U1165 (N_1165,In_187,In_666);
xor U1166 (N_1166,In_372,In_349);
xnor U1167 (N_1167,In_886,In_185);
or U1168 (N_1168,In_994,In_832);
and U1169 (N_1169,In_454,In_891);
nor U1170 (N_1170,In_320,In_211);
nand U1171 (N_1171,In_71,In_198);
and U1172 (N_1172,In_517,In_987);
nor U1173 (N_1173,In_554,In_66);
nor U1174 (N_1174,In_908,In_1061);
or U1175 (N_1175,In_768,In_628);
and U1176 (N_1176,In_654,In_660);
nor U1177 (N_1177,In_227,In_1171);
or U1178 (N_1178,In_433,In_558);
or U1179 (N_1179,In_1164,In_162);
nor U1180 (N_1180,In_1355,In_1068);
and U1181 (N_1181,In_889,In_666);
nand U1182 (N_1182,In_1013,In_1337);
and U1183 (N_1183,In_840,In_477);
nand U1184 (N_1184,In_341,In_574);
or U1185 (N_1185,In_1138,In_1220);
and U1186 (N_1186,In_873,In_297);
and U1187 (N_1187,In_1405,In_888);
xnor U1188 (N_1188,In_486,In_948);
nor U1189 (N_1189,In_660,In_842);
or U1190 (N_1190,In_1052,In_1345);
nand U1191 (N_1191,In_90,In_1135);
nor U1192 (N_1192,In_1326,In_907);
and U1193 (N_1193,In_984,In_1492);
and U1194 (N_1194,In_1455,In_350);
nor U1195 (N_1195,In_381,In_161);
or U1196 (N_1196,In_1232,In_297);
xnor U1197 (N_1197,In_59,In_934);
or U1198 (N_1198,In_385,In_1165);
and U1199 (N_1199,In_1278,In_1150);
nor U1200 (N_1200,In_953,In_1293);
or U1201 (N_1201,In_803,In_628);
or U1202 (N_1202,In_1349,In_1369);
nor U1203 (N_1203,In_1039,In_1156);
nor U1204 (N_1204,In_859,In_1245);
and U1205 (N_1205,In_79,In_477);
nand U1206 (N_1206,In_1281,In_352);
nand U1207 (N_1207,In_363,In_1077);
and U1208 (N_1208,In_1265,In_195);
or U1209 (N_1209,In_144,In_147);
or U1210 (N_1210,In_1277,In_703);
or U1211 (N_1211,In_1389,In_727);
or U1212 (N_1212,In_433,In_455);
and U1213 (N_1213,In_363,In_1360);
and U1214 (N_1214,In_877,In_167);
nor U1215 (N_1215,In_1450,In_211);
and U1216 (N_1216,In_631,In_893);
or U1217 (N_1217,In_1119,In_8);
or U1218 (N_1218,In_417,In_479);
nor U1219 (N_1219,In_290,In_210);
nor U1220 (N_1220,In_970,In_1289);
and U1221 (N_1221,In_55,In_431);
nor U1222 (N_1222,In_1085,In_529);
and U1223 (N_1223,In_1234,In_764);
nand U1224 (N_1224,In_646,In_191);
and U1225 (N_1225,In_239,In_809);
and U1226 (N_1226,In_1247,In_74);
or U1227 (N_1227,In_129,In_979);
xor U1228 (N_1228,In_756,In_1214);
or U1229 (N_1229,In_101,In_1452);
nor U1230 (N_1230,In_820,In_851);
xnor U1231 (N_1231,In_821,In_1236);
and U1232 (N_1232,In_1050,In_1412);
xor U1233 (N_1233,In_405,In_958);
or U1234 (N_1234,In_61,In_703);
nor U1235 (N_1235,In_1141,In_259);
nor U1236 (N_1236,In_703,In_1118);
or U1237 (N_1237,In_236,In_258);
xor U1238 (N_1238,In_570,In_532);
or U1239 (N_1239,In_1188,In_1392);
nand U1240 (N_1240,In_1374,In_146);
nand U1241 (N_1241,In_179,In_84);
nand U1242 (N_1242,In_33,In_23);
nor U1243 (N_1243,In_852,In_865);
and U1244 (N_1244,In_663,In_1157);
nand U1245 (N_1245,In_1071,In_994);
and U1246 (N_1246,In_1336,In_1086);
and U1247 (N_1247,In_328,In_590);
and U1248 (N_1248,In_697,In_475);
or U1249 (N_1249,In_6,In_1047);
xor U1250 (N_1250,In_864,In_31);
nand U1251 (N_1251,In_435,In_528);
nand U1252 (N_1252,In_1162,In_543);
and U1253 (N_1253,In_676,In_1329);
xor U1254 (N_1254,In_1400,In_263);
nand U1255 (N_1255,In_603,In_1443);
nor U1256 (N_1256,In_1381,In_252);
nor U1257 (N_1257,In_54,In_589);
nand U1258 (N_1258,In_1379,In_725);
and U1259 (N_1259,In_1457,In_257);
xor U1260 (N_1260,In_818,In_224);
nand U1261 (N_1261,In_1198,In_336);
nor U1262 (N_1262,In_1230,In_1350);
and U1263 (N_1263,In_778,In_307);
nor U1264 (N_1264,In_278,In_1488);
or U1265 (N_1265,In_1342,In_332);
nor U1266 (N_1266,In_1352,In_264);
and U1267 (N_1267,In_227,In_1089);
nor U1268 (N_1268,In_600,In_998);
and U1269 (N_1269,In_1032,In_68);
nor U1270 (N_1270,In_351,In_905);
nor U1271 (N_1271,In_220,In_1276);
nor U1272 (N_1272,In_135,In_1233);
nor U1273 (N_1273,In_308,In_646);
nand U1274 (N_1274,In_843,In_384);
and U1275 (N_1275,In_1033,In_865);
xor U1276 (N_1276,In_528,In_293);
nor U1277 (N_1277,In_1327,In_534);
and U1278 (N_1278,In_710,In_143);
xor U1279 (N_1279,In_430,In_388);
or U1280 (N_1280,In_173,In_151);
and U1281 (N_1281,In_359,In_1393);
nor U1282 (N_1282,In_766,In_59);
nor U1283 (N_1283,In_640,In_142);
and U1284 (N_1284,In_1333,In_164);
nand U1285 (N_1285,In_1228,In_1154);
xnor U1286 (N_1286,In_1319,In_483);
and U1287 (N_1287,In_414,In_1128);
or U1288 (N_1288,In_1221,In_328);
and U1289 (N_1289,In_1084,In_1300);
or U1290 (N_1290,In_656,In_951);
nor U1291 (N_1291,In_1436,In_39);
nand U1292 (N_1292,In_266,In_1077);
nor U1293 (N_1293,In_609,In_432);
xnor U1294 (N_1294,In_286,In_821);
xnor U1295 (N_1295,In_561,In_1495);
nor U1296 (N_1296,In_174,In_964);
or U1297 (N_1297,In_1085,In_390);
nand U1298 (N_1298,In_724,In_1139);
nand U1299 (N_1299,In_375,In_1461);
nor U1300 (N_1300,In_1261,In_583);
xor U1301 (N_1301,In_885,In_1357);
or U1302 (N_1302,In_714,In_255);
or U1303 (N_1303,In_287,In_87);
nor U1304 (N_1304,In_1190,In_908);
nor U1305 (N_1305,In_1445,In_1267);
nor U1306 (N_1306,In_1232,In_31);
and U1307 (N_1307,In_1091,In_265);
or U1308 (N_1308,In_915,In_1384);
xnor U1309 (N_1309,In_261,In_1402);
and U1310 (N_1310,In_297,In_1409);
or U1311 (N_1311,In_564,In_1422);
nor U1312 (N_1312,In_544,In_1116);
nor U1313 (N_1313,In_388,In_467);
nand U1314 (N_1314,In_1114,In_825);
nor U1315 (N_1315,In_110,In_1102);
or U1316 (N_1316,In_452,In_1173);
nor U1317 (N_1317,In_509,In_531);
nand U1318 (N_1318,In_1058,In_578);
nor U1319 (N_1319,In_893,In_1059);
or U1320 (N_1320,In_654,In_646);
and U1321 (N_1321,In_9,In_92);
and U1322 (N_1322,In_1412,In_289);
nand U1323 (N_1323,In_281,In_548);
nand U1324 (N_1324,In_510,In_1009);
or U1325 (N_1325,In_993,In_1072);
and U1326 (N_1326,In_398,In_1365);
or U1327 (N_1327,In_625,In_1129);
nor U1328 (N_1328,In_896,In_542);
xnor U1329 (N_1329,In_232,In_855);
and U1330 (N_1330,In_1047,In_721);
nand U1331 (N_1331,In_578,In_140);
and U1332 (N_1332,In_1336,In_164);
nand U1333 (N_1333,In_306,In_556);
or U1334 (N_1334,In_734,In_1250);
nor U1335 (N_1335,In_1384,In_778);
nor U1336 (N_1336,In_786,In_1498);
and U1337 (N_1337,In_983,In_574);
and U1338 (N_1338,In_1143,In_1448);
nor U1339 (N_1339,In_1359,In_957);
xnor U1340 (N_1340,In_290,In_1199);
nor U1341 (N_1341,In_1479,In_629);
or U1342 (N_1342,In_1386,In_520);
nor U1343 (N_1343,In_491,In_1464);
nand U1344 (N_1344,In_1114,In_400);
and U1345 (N_1345,In_12,In_511);
xor U1346 (N_1346,In_43,In_103);
nand U1347 (N_1347,In_177,In_151);
nor U1348 (N_1348,In_1277,In_294);
xnor U1349 (N_1349,In_277,In_1424);
nor U1350 (N_1350,In_1044,In_374);
and U1351 (N_1351,In_38,In_184);
nor U1352 (N_1352,In_346,In_1421);
nor U1353 (N_1353,In_24,In_553);
xor U1354 (N_1354,In_93,In_327);
and U1355 (N_1355,In_329,In_446);
nor U1356 (N_1356,In_688,In_135);
nor U1357 (N_1357,In_998,In_383);
nor U1358 (N_1358,In_412,In_1414);
nand U1359 (N_1359,In_653,In_1436);
nor U1360 (N_1360,In_1113,In_1264);
and U1361 (N_1361,In_1302,In_302);
or U1362 (N_1362,In_781,In_464);
nand U1363 (N_1363,In_657,In_221);
and U1364 (N_1364,In_97,In_133);
nor U1365 (N_1365,In_1071,In_304);
xnor U1366 (N_1366,In_953,In_1157);
nor U1367 (N_1367,In_1472,In_53);
nor U1368 (N_1368,In_1350,In_561);
nand U1369 (N_1369,In_1232,In_611);
xor U1370 (N_1370,In_89,In_589);
nand U1371 (N_1371,In_1360,In_512);
xor U1372 (N_1372,In_1397,In_551);
or U1373 (N_1373,In_707,In_91);
and U1374 (N_1374,In_451,In_1421);
and U1375 (N_1375,In_1244,In_710);
nor U1376 (N_1376,In_16,In_37);
and U1377 (N_1377,In_1337,In_613);
or U1378 (N_1378,In_1363,In_242);
nand U1379 (N_1379,In_420,In_615);
and U1380 (N_1380,In_146,In_1439);
or U1381 (N_1381,In_838,In_312);
nand U1382 (N_1382,In_854,In_676);
or U1383 (N_1383,In_929,In_1450);
and U1384 (N_1384,In_892,In_250);
and U1385 (N_1385,In_261,In_1280);
and U1386 (N_1386,In_656,In_830);
nor U1387 (N_1387,In_1051,In_732);
and U1388 (N_1388,In_965,In_177);
nor U1389 (N_1389,In_925,In_125);
xnor U1390 (N_1390,In_1076,In_1059);
nor U1391 (N_1391,In_109,In_580);
nor U1392 (N_1392,In_1492,In_459);
and U1393 (N_1393,In_550,In_602);
xnor U1394 (N_1394,In_416,In_540);
and U1395 (N_1395,In_718,In_1325);
or U1396 (N_1396,In_1412,In_187);
and U1397 (N_1397,In_1127,In_346);
and U1398 (N_1398,In_173,In_1);
or U1399 (N_1399,In_1203,In_1117);
or U1400 (N_1400,In_139,In_948);
and U1401 (N_1401,In_1446,In_1006);
and U1402 (N_1402,In_1454,In_555);
and U1403 (N_1403,In_1129,In_1102);
nor U1404 (N_1404,In_613,In_80);
nor U1405 (N_1405,In_44,In_156);
and U1406 (N_1406,In_753,In_508);
nor U1407 (N_1407,In_101,In_988);
and U1408 (N_1408,In_1202,In_704);
or U1409 (N_1409,In_1033,In_843);
or U1410 (N_1410,In_663,In_845);
nor U1411 (N_1411,In_7,In_121);
nand U1412 (N_1412,In_130,In_669);
or U1413 (N_1413,In_721,In_260);
nand U1414 (N_1414,In_368,In_159);
and U1415 (N_1415,In_639,In_1032);
or U1416 (N_1416,In_801,In_1407);
and U1417 (N_1417,In_1110,In_1478);
and U1418 (N_1418,In_674,In_273);
nor U1419 (N_1419,In_11,In_1063);
nor U1420 (N_1420,In_578,In_263);
nand U1421 (N_1421,In_388,In_816);
nand U1422 (N_1422,In_1233,In_954);
and U1423 (N_1423,In_1415,In_1319);
nor U1424 (N_1424,In_967,In_582);
xor U1425 (N_1425,In_1142,In_841);
or U1426 (N_1426,In_838,In_4);
and U1427 (N_1427,In_333,In_644);
nand U1428 (N_1428,In_1371,In_348);
or U1429 (N_1429,In_96,In_1095);
and U1430 (N_1430,In_374,In_1290);
and U1431 (N_1431,In_575,In_348);
nor U1432 (N_1432,In_1060,In_1145);
nand U1433 (N_1433,In_1279,In_503);
and U1434 (N_1434,In_983,In_585);
xor U1435 (N_1435,In_619,In_1386);
nand U1436 (N_1436,In_869,In_942);
and U1437 (N_1437,In_167,In_297);
xor U1438 (N_1438,In_233,In_171);
nor U1439 (N_1439,In_1399,In_691);
nor U1440 (N_1440,In_1415,In_942);
or U1441 (N_1441,In_318,In_69);
nor U1442 (N_1442,In_256,In_242);
nor U1443 (N_1443,In_622,In_1003);
and U1444 (N_1444,In_290,In_663);
and U1445 (N_1445,In_1166,In_1176);
and U1446 (N_1446,In_378,In_76);
nand U1447 (N_1447,In_1371,In_190);
xnor U1448 (N_1448,In_1165,In_1309);
xnor U1449 (N_1449,In_141,In_1404);
nor U1450 (N_1450,In_830,In_508);
nand U1451 (N_1451,In_818,In_510);
nor U1452 (N_1452,In_650,In_1483);
xor U1453 (N_1453,In_1137,In_849);
or U1454 (N_1454,In_203,In_780);
nor U1455 (N_1455,In_975,In_1190);
and U1456 (N_1456,In_669,In_1008);
xnor U1457 (N_1457,In_414,In_599);
nand U1458 (N_1458,In_888,In_671);
or U1459 (N_1459,In_1091,In_1201);
or U1460 (N_1460,In_436,In_500);
nor U1461 (N_1461,In_1164,In_804);
nand U1462 (N_1462,In_1186,In_1211);
xor U1463 (N_1463,In_398,In_1024);
nand U1464 (N_1464,In_667,In_1063);
or U1465 (N_1465,In_1028,In_587);
or U1466 (N_1466,In_927,In_1313);
nor U1467 (N_1467,In_1359,In_1436);
and U1468 (N_1468,In_331,In_48);
nand U1469 (N_1469,In_1142,In_203);
or U1470 (N_1470,In_192,In_1323);
nand U1471 (N_1471,In_574,In_1034);
and U1472 (N_1472,In_182,In_909);
or U1473 (N_1473,In_1298,In_857);
xor U1474 (N_1474,In_1114,In_961);
or U1475 (N_1475,In_1217,In_949);
nand U1476 (N_1476,In_788,In_440);
or U1477 (N_1477,In_1090,In_1038);
xnor U1478 (N_1478,In_723,In_149);
or U1479 (N_1479,In_578,In_1048);
or U1480 (N_1480,In_1070,In_471);
xor U1481 (N_1481,In_991,In_381);
nand U1482 (N_1482,In_668,In_676);
nor U1483 (N_1483,In_1298,In_191);
nor U1484 (N_1484,In_1454,In_397);
and U1485 (N_1485,In_62,In_851);
nand U1486 (N_1486,In_122,In_505);
and U1487 (N_1487,In_156,In_588);
or U1488 (N_1488,In_1484,In_865);
nand U1489 (N_1489,In_487,In_1375);
nand U1490 (N_1490,In_1196,In_879);
and U1491 (N_1491,In_692,In_772);
nor U1492 (N_1492,In_545,In_1281);
or U1493 (N_1493,In_631,In_1471);
xnor U1494 (N_1494,In_783,In_1334);
or U1495 (N_1495,In_852,In_519);
and U1496 (N_1496,In_174,In_490);
nand U1497 (N_1497,In_468,In_374);
nor U1498 (N_1498,In_320,In_1021);
or U1499 (N_1499,In_13,In_775);
and U1500 (N_1500,In_834,In_1338);
and U1501 (N_1501,In_1073,In_794);
nor U1502 (N_1502,In_367,In_371);
nand U1503 (N_1503,In_908,In_601);
nor U1504 (N_1504,In_908,In_1369);
nand U1505 (N_1505,In_1076,In_1070);
and U1506 (N_1506,In_1065,In_1495);
nor U1507 (N_1507,In_73,In_998);
or U1508 (N_1508,In_42,In_1047);
nor U1509 (N_1509,In_213,In_1276);
and U1510 (N_1510,In_1205,In_854);
nor U1511 (N_1511,In_533,In_312);
and U1512 (N_1512,In_864,In_845);
nand U1513 (N_1513,In_1004,In_1160);
or U1514 (N_1514,In_77,In_1131);
nor U1515 (N_1515,In_246,In_81);
and U1516 (N_1516,In_321,In_1258);
or U1517 (N_1517,In_1372,In_1455);
and U1518 (N_1518,In_708,In_280);
nand U1519 (N_1519,In_259,In_69);
or U1520 (N_1520,In_886,In_1435);
xor U1521 (N_1521,In_1405,In_369);
nand U1522 (N_1522,In_1423,In_584);
nor U1523 (N_1523,In_1035,In_1306);
or U1524 (N_1524,In_1220,In_309);
xor U1525 (N_1525,In_11,In_997);
nand U1526 (N_1526,In_962,In_1170);
nand U1527 (N_1527,In_1481,In_1419);
nand U1528 (N_1528,In_731,In_565);
nor U1529 (N_1529,In_1006,In_966);
or U1530 (N_1530,In_888,In_595);
xor U1531 (N_1531,In_1183,In_1025);
nand U1532 (N_1532,In_964,In_1216);
and U1533 (N_1533,In_1309,In_206);
nand U1534 (N_1534,In_990,In_113);
or U1535 (N_1535,In_269,In_681);
xor U1536 (N_1536,In_1007,In_634);
nand U1537 (N_1537,In_769,In_1156);
nor U1538 (N_1538,In_362,In_1051);
and U1539 (N_1539,In_46,In_1325);
nand U1540 (N_1540,In_1393,In_534);
xnor U1541 (N_1541,In_1006,In_800);
or U1542 (N_1542,In_1396,In_129);
nor U1543 (N_1543,In_356,In_284);
nor U1544 (N_1544,In_512,In_424);
nand U1545 (N_1545,In_528,In_126);
xor U1546 (N_1546,In_502,In_722);
and U1547 (N_1547,In_1151,In_616);
and U1548 (N_1548,In_1265,In_1131);
or U1549 (N_1549,In_406,In_1219);
xor U1550 (N_1550,In_1151,In_1326);
or U1551 (N_1551,In_167,In_796);
nor U1552 (N_1552,In_296,In_726);
or U1553 (N_1553,In_22,In_200);
nor U1554 (N_1554,In_167,In_1408);
or U1555 (N_1555,In_1273,In_1070);
nor U1556 (N_1556,In_993,In_564);
xnor U1557 (N_1557,In_1372,In_961);
and U1558 (N_1558,In_882,In_893);
and U1559 (N_1559,In_1470,In_903);
nand U1560 (N_1560,In_234,In_48);
or U1561 (N_1561,In_948,In_401);
xnor U1562 (N_1562,In_722,In_482);
nor U1563 (N_1563,In_1429,In_107);
or U1564 (N_1564,In_1270,In_1477);
and U1565 (N_1565,In_1058,In_110);
or U1566 (N_1566,In_239,In_838);
nor U1567 (N_1567,In_539,In_624);
nand U1568 (N_1568,In_41,In_311);
xor U1569 (N_1569,In_953,In_952);
xnor U1570 (N_1570,In_1044,In_613);
nor U1571 (N_1571,In_68,In_362);
or U1572 (N_1572,In_914,In_576);
and U1573 (N_1573,In_1151,In_584);
nor U1574 (N_1574,In_1129,In_1244);
nor U1575 (N_1575,In_1388,In_884);
and U1576 (N_1576,In_591,In_1467);
nand U1577 (N_1577,In_1008,In_622);
nor U1578 (N_1578,In_528,In_643);
and U1579 (N_1579,In_1057,In_1396);
nor U1580 (N_1580,In_1386,In_168);
and U1581 (N_1581,In_923,In_744);
or U1582 (N_1582,In_689,In_717);
xnor U1583 (N_1583,In_439,In_924);
and U1584 (N_1584,In_1273,In_467);
and U1585 (N_1585,In_1290,In_983);
xnor U1586 (N_1586,In_286,In_1253);
xor U1587 (N_1587,In_744,In_1460);
or U1588 (N_1588,In_1215,In_1278);
nand U1589 (N_1589,In_562,In_94);
nor U1590 (N_1590,In_1281,In_163);
xor U1591 (N_1591,In_823,In_78);
nor U1592 (N_1592,In_526,In_665);
xor U1593 (N_1593,In_1470,In_633);
and U1594 (N_1594,In_405,In_1348);
and U1595 (N_1595,In_1021,In_1357);
nand U1596 (N_1596,In_1206,In_248);
or U1597 (N_1597,In_1048,In_1203);
nor U1598 (N_1598,In_372,In_497);
or U1599 (N_1599,In_92,In_280);
nand U1600 (N_1600,In_912,In_1307);
and U1601 (N_1601,In_517,In_702);
nor U1602 (N_1602,In_677,In_676);
nand U1603 (N_1603,In_1350,In_1096);
nand U1604 (N_1604,In_882,In_553);
xor U1605 (N_1605,In_997,In_724);
and U1606 (N_1606,In_1311,In_1340);
nand U1607 (N_1607,In_539,In_1460);
nor U1608 (N_1608,In_1180,In_1076);
or U1609 (N_1609,In_784,In_585);
and U1610 (N_1610,In_731,In_652);
nor U1611 (N_1611,In_795,In_1187);
or U1612 (N_1612,In_759,In_182);
or U1613 (N_1613,In_1478,In_517);
or U1614 (N_1614,In_378,In_382);
or U1615 (N_1615,In_1050,In_1465);
nor U1616 (N_1616,In_238,In_946);
or U1617 (N_1617,In_42,In_731);
and U1618 (N_1618,In_617,In_1464);
and U1619 (N_1619,In_890,In_1369);
nor U1620 (N_1620,In_991,In_542);
or U1621 (N_1621,In_177,In_23);
nor U1622 (N_1622,In_18,In_1270);
nand U1623 (N_1623,In_845,In_521);
or U1624 (N_1624,In_673,In_806);
or U1625 (N_1625,In_753,In_648);
or U1626 (N_1626,In_686,In_587);
nand U1627 (N_1627,In_814,In_1458);
nor U1628 (N_1628,In_917,In_1365);
or U1629 (N_1629,In_491,In_984);
nand U1630 (N_1630,In_557,In_203);
nand U1631 (N_1631,In_274,In_1498);
nand U1632 (N_1632,In_875,In_789);
or U1633 (N_1633,In_501,In_1089);
nor U1634 (N_1634,In_1472,In_840);
and U1635 (N_1635,In_375,In_372);
or U1636 (N_1636,In_1434,In_1199);
and U1637 (N_1637,In_168,In_439);
or U1638 (N_1638,In_1277,In_895);
or U1639 (N_1639,In_56,In_243);
nand U1640 (N_1640,In_706,In_602);
and U1641 (N_1641,In_1059,In_721);
and U1642 (N_1642,In_484,In_296);
nor U1643 (N_1643,In_752,In_936);
nor U1644 (N_1644,In_1373,In_824);
and U1645 (N_1645,In_629,In_347);
or U1646 (N_1646,In_902,In_145);
nand U1647 (N_1647,In_250,In_57);
or U1648 (N_1648,In_3,In_318);
nand U1649 (N_1649,In_766,In_238);
xor U1650 (N_1650,In_238,In_1339);
nand U1651 (N_1651,In_432,In_1409);
nor U1652 (N_1652,In_485,In_1149);
and U1653 (N_1653,In_673,In_830);
nand U1654 (N_1654,In_829,In_1399);
nand U1655 (N_1655,In_859,In_775);
and U1656 (N_1656,In_1099,In_510);
or U1657 (N_1657,In_681,In_821);
nor U1658 (N_1658,In_836,In_1081);
nand U1659 (N_1659,In_1041,In_519);
nand U1660 (N_1660,In_717,In_132);
nor U1661 (N_1661,In_687,In_1213);
nor U1662 (N_1662,In_247,In_434);
or U1663 (N_1663,In_133,In_875);
or U1664 (N_1664,In_705,In_979);
or U1665 (N_1665,In_158,In_226);
nand U1666 (N_1666,In_482,In_1291);
nor U1667 (N_1667,In_509,In_1349);
nor U1668 (N_1668,In_637,In_779);
nor U1669 (N_1669,In_744,In_915);
and U1670 (N_1670,In_496,In_504);
and U1671 (N_1671,In_472,In_181);
nor U1672 (N_1672,In_120,In_72);
nand U1673 (N_1673,In_454,In_195);
nor U1674 (N_1674,In_49,In_50);
nor U1675 (N_1675,In_989,In_1085);
nand U1676 (N_1676,In_1139,In_174);
or U1677 (N_1677,In_1126,In_1073);
or U1678 (N_1678,In_54,In_1463);
and U1679 (N_1679,In_1094,In_948);
or U1680 (N_1680,In_242,In_3);
and U1681 (N_1681,In_1215,In_63);
or U1682 (N_1682,In_1005,In_1078);
nor U1683 (N_1683,In_873,In_127);
nand U1684 (N_1684,In_894,In_509);
nand U1685 (N_1685,In_1402,In_462);
xnor U1686 (N_1686,In_1056,In_1499);
or U1687 (N_1687,In_19,In_1117);
or U1688 (N_1688,In_829,In_481);
nand U1689 (N_1689,In_498,In_1286);
and U1690 (N_1690,In_1428,In_973);
nor U1691 (N_1691,In_1381,In_193);
nor U1692 (N_1692,In_93,In_672);
nor U1693 (N_1693,In_14,In_741);
nor U1694 (N_1694,In_1424,In_305);
or U1695 (N_1695,In_1421,In_917);
nand U1696 (N_1696,In_977,In_888);
nor U1697 (N_1697,In_1185,In_1408);
nor U1698 (N_1698,In_388,In_946);
nand U1699 (N_1699,In_1398,In_858);
xor U1700 (N_1700,In_274,In_185);
or U1701 (N_1701,In_60,In_126);
xor U1702 (N_1702,In_144,In_1171);
nand U1703 (N_1703,In_1163,In_1207);
nand U1704 (N_1704,In_714,In_858);
and U1705 (N_1705,In_1398,In_826);
nor U1706 (N_1706,In_1446,In_63);
nor U1707 (N_1707,In_1358,In_1218);
nand U1708 (N_1708,In_709,In_264);
nor U1709 (N_1709,In_1221,In_190);
and U1710 (N_1710,In_1439,In_929);
and U1711 (N_1711,In_280,In_148);
and U1712 (N_1712,In_637,In_1345);
or U1713 (N_1713,In_170,In_104);
nand U1714 (N_1714,In_632,In_1065);
nand U1715 (N_1715,In_861,In_759);
xor U1716 (N_1716,In_749,In_763);
and U1717 (N_1717,In_1079,In_1085);
and U1718 (N_1718,In_1284,In_377);
or U1719 (N_1719,In_313,In_166);
nand U1720 (N_1720,In_738,In_945);
nor U1721 (N_1721,In_1101,In_266);
nor U1722 (N_1722,In_311,In_985);
and U1723 (N_1723,In_637,In_440);
nand U1724 (N_1724,In_790,In_1090);
nor U1725 (N_1725,In_473,In_698);
or U1726 (N_1726,In_297,In_1431);
xor U1727 (N_1727,In_1307,In_1317);
or U1728 (N_1728,In_461,In_682);
or U1729 (N_1729,In_1116,In_1039);
or U1730 (N_1730,In_587,In_471);
nor U1731 (N_1731,In_128,In_855);
or U1732 (N_1732,In_137,In_1373);
or U1733 (N_1733,In_565,In_1254);
xor U1734 (N_1734,In_561,In_162);
nand U1735 (N_1735,In_826,In_1133);
and U1736 (N_1736,In_1388,In_659);
or U1737 (N_1737,In_67,In_989);
and U1738 (N_1738,In_1287,In_1486);
and U1739 (N_1739,In_543,In_334);
or U1740 (N_1740,In_670,In_1487);
nor U1741 (N_1741,In_73,In_398);
and U1742 (N_1742,In_329,In_784);
or U1743 (N_1743,In_890,In_156);
xnor U1744 (N_1744,In_1443,In_84);
or U1745 (N_1745,In_47,In_283);
or U1746 (N_1746,In_1340,In_835);
or U1747 (N_1747,In_970,In_1075);
nand U1748 (N_1748,In_1365,In_401);
and U1749 (N_1749,In_905,In_192);
xnor U1750 (N_1750,In_1006,In_1291);
and U1751 (N_1751,In_752,In_564);
or U1752 (N_1752,In_611,In_627);
nor U1753 (N_1753,In_240,In_859);
nor U1754 (N_1754,In_638,In_1181);
nor U1755 (N_1755,In_692,In_516);
nand U1756 (N_1756,In_954,In_1080);
nand U1757 (N_1757,In_879,In_183);
or U1758 (N_1758,In_744,In_956);
or U1759 (N_1759,In_703,In_341);
nor U1760 (N_1760,In_1005,In_53);
and U1761 (N_1761,In_303,In_169);
nand U1762 (N_1762,In_691,In_211);
and U1763 (N_1763,In_1297,In_1364);
nor U1764 (N_1764,In_186,In_1369);
and U1765 (N_1765,In_1371,In_142);
nand U1766 (N_1766,In_197,In_1375);
and U1767 (N_1767,In_64,In_421);
and U1768 (N_1768,In_546,In_1474);
nand U1769 (N_1769,In_322,In_1074);
or U1770 (N_1770,In_910,In_631);
or U1771 (N_1771,In_115,In_40);
nand U1772 (N_1772,In_1284,In_1452);
nand U1773 (N_1773,In_850,In_185);
nor U1774 (N_1774,In_1067,In_206);
nor U1775 (N_1775,In_558,In_420);
and U1776 (N_1776,In_391,In_1383);
nand U1777 (N_1777,In_1257,In_445);
and U1778 (N_1778,In_289,In_1261);
or U1779 (N_1779,In_1355,In_237);
nor U1780 (N_1780,In_811,In_657);
and U1781 (N_1781,In_937,In_765);
and U1782 (N_1782,In_959,In_963);
and U1783 (N_1783,In_978,In_464);
nand U1784 (N_1784,In_1305,In_1067);
or U1785 (N_1785,In_1048,In_1113);
nand U1786 (N_1786,In_1229,In_440);
xnor U1787 (N_1787,In_242,In_840);
nand U1788 (N_1788,In_219,In_209);
and U1789 (N_1789,In_853,In_917);
nand U1790 (N_1790,In_364,In_467);
xor U1791 (N_1791,In_1446,In_949);
nand U1792 (N_1792,In_265,In_480);
nor U1793 (N_1793,In_251,In_1385);
and U1794 (N_1794,In_242,In_81);
nor U1795 (N_1795,In_635,In_561);
nand U1796 (N_1796,In_486,In_806);
nand U1797 (N_1797,In_148,In_548);
nor U1798 (N_1798,In_787,In_626);
nand U1799 (N_1799,In_1098,In_699);
nand U1800 (N_1800,In_1326,In_1344);
or U1801 (N_1801,In_1138,In_150);
nor U1802 (N_1802,In_635,In_186);
nor U1803 (N_1803,In_369,In_1061);
and U1804 (N_1804,In_90,In_1091);
nor U1805 (N_1805,In_334,In_524);
nor U1806 (N_1806,In_49,In_940);
nor U1807 (N_1807,In_312,In_1222);
and U1808 (N_1808,In_1050,In_1391);
nor U1809 (N_1809,In_1441,In_1048);
or U1810 (N_1810,In_1417,In_1141);
and U1811 (N_1811,In_1134,In_691);
nor U1812 (N_1812,In_1067,In_337);
nand U1813 (N_1813,In_1051,In_1358);
nor U1814 (N_1814,In_220,In_852);
or U1815 (N_1815,In_1060,In_1036);
nand U1816 (N_1816,In_1167,In_28);
or U1817 (N_1817,In_305,In_963);
nor U1818 (N_1818,In_1402,In_23);
nor U1819 (N_1819,In_64,In_1003);
or U1820 (N_1820,In_1431,In_321);
nor U1821 (N_1821,In_188,In_175);
and U1822 (N_1822,In_654,In_868);
nor U1823 (N_1823,In_46,In_1341);
or U1824 (N_1824,In_1441,In_1230);
xnor U1825 (N_1825,In_273,In_234);
nand U1826 (N_1826,In_764,In_382);
and U1827 (N_1827,In_757,In_486);
and U1828 (N_1828,In_1227,In_488);
nand U1829 (N_1829,In_542,In_395);
or U1830 (N_1830,In_367,In_766);
or U1831 (N_1831,In_456,In_1403);
or U1832 (N_1832,In_1104,In_1406);
nand U1833 (N_1833,In_652,In_796);
nor U1834 (N_1834,In_890,In_1253);
nand U1835 (N_1835,In_881,In_331);
and U1836 (N_1836,In_1200,In_1175);
nand U1837 (N_1837,In_474,In_668);
nand U1838 (N_1838,In_299,In_779);
nand U1839 (N_1839,In_442,In_1225);
nand U1840 (N_1840,In_464,In_1258);
or U1841 (N_1841,In_352,In_1365);
nand U1842 (N_1842,In_50,In_451);
nor U1843 (N_1843,In_768,In_216);
or U1844 (N_1844,In_1491,In_995);
nand U1845 (N_1845,In_54,In_931);
nor U1846 (N_1846,In_1420,In_225);
and U1847 (N_1847,In_237,In_415);
nor U1848 (N_1848,In_229,In_1071);
xnor U1849 (N_1849,In_662,In_982);
nor U1850 (N_1850,In_1093,In_571);
and U1851 (N_1851,In_448,In_1038);
and U1852 (N_1852,In_740,In_650);
nand U1853 (N_1853,In_188,In_1385);
nor U1854 (N_1854,In_415,In_1435);
nand U1855 (N_1855,In_303,In_1384);
nor U1856 (N_1856,In_788,In_1412);
nand U1857 (N_1857,In_109,In_1389);
nor U1858 (N_1858,In_547,In_1035);
and U1859 (N_1859,In_209,In_1274);
xor U1860 (N_1860,In_1219,In_1375);
nor U1861 (N_1861,In_906,In_329);
and U1862 (N_1862,In_87,In_1204);
nor U1863 (N_1863,In_489,In_1329);
nand U1864 (N_1864,In_1379,In_1366);
nand U1865 (N_1865,In_725,In_1094);
or U1866 (N_1866,In_340,In_510);
nor U1867 (N_1867,In_70,In_1326);
xnor U1868 (N_1868,In_527,In_657);
or U1869 (N_1869,In_666,In_102);
or U1870 (N_1870,In_111,In_480);
and U1871 (N_1871,In_1023,In_1094);
xor U1872 (N_1872,In_1406,In_1317);
nand U1873 (N_1873,In_1059,In_638);
and U1874 (N_1874,In_753,In_1222);
and U1875 (N_1875,In_1412,In_385);
or U1876 (N_1876,In_1240,In_1415);
or U1877 (N_1877,In_1211,In_1201);
nor U1878 (N_1878,In_1200,In_193);
or U1879 (N_1879,In_898,In_254);
nor U1880 (N_1880,In_1051,In_530);
nor U1881 (N_1881,In_1184,In_627);
and U1882 (N_1882,In_786,In_970);
or U1883 (N_1883,In_640,In_521);
or U1884 (N_1884,In_55,In_151);
and U1885 (N_1885,In_667,In_1382);
or U1886 (N_1886,In_1207,In_413);
xnor U1887 (N_1887,In_1451,In_333);
and U1888 (N_1888,In_1489,In_21);
nand U1889 (N_1889,In_823,In_115);
xnor U1890 (N_1890,In_1172,In_713);
nor U1891 (N_1891,In_911,In_244);
xnor U1892 (N_1892,In_1406,In_959);
or U1893 (N_1893,In_1089,In_553);
and U1894 (N_1894,In_1109,In_759);
and U1895 (N_1895,In_412,In_561);
or U1896 (N_1896,In_939,In_656);
nor U1897 (N_1897,In_1403,In_1400);
nand U1898 (N_1898,In_487,In_316);
and U1899 (N_1899,In_1306,In_841);
or U1900 (N_1900,In_1346,In_994);
xor U1901 (N_1901,In_1380,In_984);
xor U1902 (N_1902,In_809,In_1061);
nor U1903 (N_1903,In_532,In_180);
xnor U1904 (N_1904,In_412,In_1234);
nand U1905 (N_1905,In_1203,In_1417);
xnor U1906 (N_1906,In_1061,In_1440);
and U1907 (N_1907,In_535,In_117);
nand U1908 (N_1908,In_805,In_291);
and U1909 (N_1909,In_340,In_1179);
or U1910 (N_1910,In_970,In_430);
or U1911 (N_1911,In_780,In_459);
or U1912 (N_1912,In_1469,In_380);
nor U1913 (N_1913,In_508,In_94);
or U1914 (N_1914,In_514,In_1011);
nor U1915 (N_1915,In_1013,In_135);
and U1916 (N_1916,In_528,In_1184);
or U1917 (N_1917,In_19,In_225);
or U1918 (N_1918,In_794,In_274);
nand U1919 (N_1919,In_1247,In_824);
nor U1920 (N_1920,In_836,In_1008);
or U1921 (N_1921,In_86,In_80);
nor U1922 (N_1922,In_1459,In_1443);
nand U1923 (N_1923,In_452,In_1320);
or U1924 (N_1924,In_655,In_703);
xnor U1925 (N_1925,In_1014,In_144);
xnor U1926 (N_1926,In_1299,In_947);
or U1927 (N_1927,In_845,In_1267);
and U1928 (N_1928,In_432,In_726);
nor U1929 (N_1929,In_1291,In_820);
nand U1930 (N_1930,In_1463,In_144);
and U1931 (N_1931,In_737,In_1009);
nor U1932 (N_1932,In_1076,In_956);
xnor U1933 (N_1933,In_1193,In_316);
nor U1934 (N_1934,In_33,In_183);
nor U1935 (N_1935,In_1095,In_1397);
nor U1936 (N_1936,In_499,In_863);
nand U1937 (N_1937,In_1014,In_45);
and U1938 (N_1938,In_1115,In_1174);
and U1939 (N_1939,In_489,In_151);
nand U1940 (N_1940,In_873,In_1307);
nor U1941 (N_1941,In_398,In_216);
and U1942 (N_1942,In_869,In_168);
or U1943 (N_1943,In_996,In_441);
and U1944 (N_1944,In_975,In_509);
nor U1945 (N_1945,In_1108,In_1266);
nor U1946 (N_1946,In_611,In_482);
nor U1947 (N_1947,In_897,In_1096);
or U1948 (N_1948,In_695,In_1163);
and U1949 (N_1949,In_66,In_578);
nor U1950 (N_1950,In_1431,In_116);
and U1951 (N_1951,In_1008,In_1066);
nor U1952 (N_1952,In_73,In_26);
nor U1953 (N_1953,In_1166,In_1459);
xor U1954 (N_1954,In_1059,In_968);
nor U1955 (N_1955,In_1469,In_589);
nand U1956 (N_1956,In_513,In_1225);
or U1957 (N_1957,In_1072,In_36);
nand U1958 (N_1958,In_475,In_1211);
xor U1959 (N_1959,In_1158,In_333);
nor U1960 (N_1960,In_667,In_1431);
or U1961 (N_1961,In_345,In_1447);
and U1962 (N_1962,In_873,In_876);
nand U1963 (N_1963,In_159,In_1490);
and U1964 (N_1964,In_635,In_359);
nand U1965 (N_1965,In_845,In_648);
and U1966 (N_1966,In_837,In_776);
or U1967 (N_1967,In_378,In_827);
nor U1968 (N_1968,In_951,In_1494);
or U1969 (N_1969,In_1424,In_461);
or U1970 (N_1970,In_1263,In_44);
and U1971 (N_1971,In_708,In_1112);
nor U1972 (N_1972,In_1487,In_825);
or U1973 (N_1973,In_1111,In_1091);
nand U1974 (N_1974,In_608,In_762);
nor U1975 (N_1975,In_764,In_493);
nand U1976 (N_1976,In_683,In_1088);
and U1977 (N_1977,In_598,In_575);
or U1978 (N_1978,In_1304,In_1271);
nor U1979 (N_1979,In_774,In_458);
and U1980 (N_1980,In_1166,In_1475);
or U1981 (N_1981,In_1441,In_1120);
or U1982 (N_1982,In_1414,In_1299);
nand U1983 (N_1983,In_291,In_197);
or U1984 (N_1984,In_950,In_273);
xnor U1985 (N_1985,In_22,In_823);
nor U1986 (N_1986,In_733,In_47);
nand U1987 (N_1987,In_1153,In_1211);
and U1988 (N_1988,In_1226,In_714);
nor U1989 (N_1989,In_106,In_694);
xnor U1990 (N_1990,In_1445,In_297);
and U1991 (N_1991,In_308,In_1045);
and U1992 (N_1992,In_540,In_709);
nor U1993 (N_1993,In_1046,In_1236);
nand U1994 (N_1994,In_455,In_1242);
nand U1995 (N_1995,In_985,In_1065);
or U1996 (N_1996,In_1020,In_278);
nor U1997 (N_1997,In_760,In_1270);
and U1998 (N_1998,In_392,In_729);
nor U1999 (N_1999,In_905,In_1055);
or U2000 (N_2000,In_471,In_98);
and U2001 (N_2001,In_569,In_640);
nor U2002 (N_2002,In_378,In_165);
nor U2003 (N_2003,In_738,In_165);
nor U2004 (N_2004,In_860,In_388);
and U2005 (N_2005,In_279,In_1368);
nor U2006 (N_2006,In_995,In_130);
nor U2007 (N_2007,In_1369,In_1182);
or U2008 (N_2008,In_381,In_1218);
nand U2009 (N_2009,In_119,In_554);
or U2010 (N_2010,In_1303,In_279);
xnor U2011 (N_2011,In_1033,In_1316);
nand U2012 (N_2012,In_671,In_569);
or U2013 (N_2013,In_665,In_681);
nand U2014 (N_2014,In_1068,In_633);
nor U2015 (N_2015,In_215,In_1059);
or U2016 (N_2016,In_1433,In_737);
or U2017 (N_2017,In_885,In_685);
xor U2018 (N_2018,In_403,In_496);
nor U2019 (N_2019,In_325,In_1497);
or U2020 (N_2020,In_1474,In_255);
nor U2021 (N_2021,In_141,In_484);
or U2022 (N_2022,In_129,In_958);
nor U2023 (N_2023,In_1222,In_188);
or U2024 (N_2024,In_190,In_737);
nand U2025 (N_2025,In_1362,In_451);
nand U2026 (N_2026,In_1370,In_673);
xnor U2027 (N_2027,In_903,In_45);
and U2028 (N_2028,In_924,In_394);
and U2029 (N_2029,In_116,In_1261);
or U2030 (N_2030,In_1347,In_666);
and U2031 (N_2031,In_1006,In_666);
nor U2032 (N_2032,In_1235,In_724);
nand U2033 (N_2033,In_410,In_754);
nor U2034 (N_2034,In_384,In_959);
xnor U2035 (N_2035,In_1480,In_134);
or U2036 (N_2036,In_1072,In_1481);
nor U2037 (N_2037,In_655,In_356);
and U2038 (N_2038,In_422,In_490);
or U2039 (N_2039,In_295,In_1131);
nand U2040 (N_2040,In_507,In_541);
and U2041 (N_2041,In_629,In_1401);
and U2042 (N_2042,In_260,In_1208);
xor U2043 (N_2043,In_1011,In_77);
and U2044 (N_2044,In_356,In_516);
or U2045 (N_2045,In_135,In_728);
nand U2046 (N_2046,In_111,In_1168);
nand U2047 (N_2047,In_885,In_1344);
or U2048 (N_2048,In_846,In_623);
nor U2049 (N_2049,In_690,In_807);
and U2050 (N_2050,In_951,In_499);
and U2051 (N_2051,In_1288,In_840);
and U2052 (N_2052,In_859,In_1122);
xor U2053 (N_2053,In_413,In_872);
or U2054 (N_2054,In_655,In_645);
nand U2055 (N_2055,In_1326,In_1190);
or U2056 (N_2056,In_190,In_504);
nor U2057 (N_2057,In_668,In_113);
or U2058 (N_2058,In_559,In_467);
or U2059 (N_2059,In_1415,In_1350);
and U2060 (N_2060,In_906,In_983);
and U2061 (N_2061,In_1388,In_906);
or U2062 (N_2062,In_1104,In_667);
and U2063 (N_2063,In_12,In_1101);
nor U2064 (N_2064,In_720,In_603);
xnor U2065 (N_2065,In_1459,In_99);
or U2066 (N_2066,In_1003,In_1201);
or U2067 (N_2067,In_1002,In_12);
nand U2068 (N_2068,In_1472,In_512);
or U2069 (N_2069,In_151,In_1317);
or U2070 (N_2070,In_23,In_1010);
nor U2071 (N_2071,In_189,In_1309);
nor U2072 (N_2072,In_1232,In_1142);
and U2073 (N_2073,In_47,In_1412);
or U2074 (N_2074,In_654,In_1024);
and U2075 (N_2075,In_144,In_156);
nor U2076 (N_2076,In_331,In_878);
nor U2077 (N_2077,In_934,In_538);
nand U2078 (N_2078,In_503,In_362);
nor U2079 (N_2079,In_1466,In_724);
or U2080 (N_2080,In_949,In_528);
nand U2081 (N_2081,In_97,In_12);
nor U2082 (N_2082,In_852,In_378);
nor U2083 (N_2083,In_735,In_328);
nand U2084 (N_2084,In_121,In_1478);
and U2085 (N_2085,In_1022,In_503);
and U2086 (N_2086,In_354,In_733);
xnor U2087 (N_2087,In_1146,In_746);
xnor U2088 (N_2088,In_132,In_455);
nor U2089 (N_2089,In_557,In_96);
and U2090 (N_2090,In_423,In_1081);
and U2091 (N_2091,In_818,In_86);
and U2092 (N_2092,In_1400,In_1468);
nor U2093 (N_2093,In_312,In_1390);
nor U2094 (N_2094,In_1294,In_252);
or U2095 (N_2095,In_1446,In_272);
xor U2096 (N_2096,In_1454,In_1144);
nand U2097 (N_2097,In_1204,In_1456);
nand U2098 (N_2098,In_1269,In_23);
and U2099 (N_2099,In_1243,In_481);
nor U2100 (N_2100,In_1229,In_67);
nor U2101 (N_2101,In_1065,In_302);
or U2102 (N_2102,In_1093,In_731);
xor U2103 (N_2103,In_82,In_1347);
nand U2104 (N_2104,In_905,In_1399);
and U2105 (N_2105,In_276,In_937);
and U2106 (N_2106,In_1166,In_1144);
nand U2107 (N_2107,In_1339,In_293);
or U2108 (N_2108,In_881,In_340);
or U2109 (N_2109,In_1492,In_1083);
nor U2110 (N_2110,In_1411,In_86);
nor U2111 (N_2111,In_328,In_804);
and U2112 (N_2112,In_415,In_988);
or U2113 (N_2113,In_1,In_419);
nand U2114 (N_2114,In_1336,In_485);
or U2115 (N_2115,In_399,In_507);
and U2116 (N_2116,In_43,In_943);
nor U2117 (N_2117,In_1277,In_1275);
or U2118 (N_2118,In_1126,In_645);
or U2119 (N_2119,In_621,In_885);
nand U2120 (N_2120,In_743,In_1410);
nand U2121 (N_2121,In_31,In_1385);
or U2122 (N_2122,In_1497,In_1087);
nand U2123 (N_2123,In_693,In_1192);
xor U2124 (N_2124,In_672,In_1335);
nand U2125 (N_2125,In_1072,In_41);
nor U2126 (N_2126,In_1488,In_113);
nand U2127 (N_2127,In_917,In_1437);
nand U2128 (N_2128,In_216,In_430);
or U2129 (N_2129,In_582,In_1353);
xor U2130 (N_2130,In_190,In_899);
or U2131 (N_2131,In_762,In_582);
or U2132 (N_2132,In_1497,In_835);
and U2133 (N_2133,In_353,In_292);
and U2134 (N_2134,In_266,In_595);
nor U2135 (N_2135,In_727,In_635);
nand U2136 (N_2136,In_1036,In_1029);
or U2137 (N_2137,In_517,In_849);
xnor U2138 (N_2138,In_1003,In_1031);
nand U2139 (N_2139,In_596,In_294);
nor U2140 (N_2140,In_184,In_1069);
or U2141 (N_2141,In_21,In_833);
nand U2142 (N_2142,In_288,In_1453);
or U2143 (N_2143,In_898,In_640);
and U2144 (N_2144,In_268,In_361);
and U2145 (N_2145,In_1093,In_638);
nor U2146 (N_2146,In_201,In_931);
and U2147 (N_2147,In_744,In_1235);
nand U2148 (N_2148,In_1319,In_1216);
and U2149 (N_2149,In_1172,In_922);
or U2150 (N_2150,In_1007,In_1432);
or U2151 (N_2151,In_187,In_810);
nand U2152 (N_2152,In_1280,In_1367);
xor U2153 (N_2153,In_458,In_518);
and U2154 (N_2154,In_798,In_626);
xor U2155 (N_2155,In_20,In_979);
and U2156 (N_2156,In_650,In_390);
or U2157 (N_2157,In_1101,In_1244);
nand U2158 (N_2158,In_1050,In_52);
nand U2159 (N_2159,In_1411,In_1107);
and U2160 (N_2160,In_921,In_509);
or U2161 (N_2161,In_869,In_1306);
nand U2162 (N_2162,In_369,In_657);
and U2163 (N_2163,In_1287,In_1378);
nand U2164 (N_2164,In_33,In_806);
or U2165 (N_2165,In_762,In_1339);
nor U2166 (N_2166,In_443,In_1041);
or U2167 (N_2167,In_1096,In_388);
or U2168 (N_2168,In_29,In_593);
nor U2169 (N_2169,In_893,In_1171);
nand U2170 (N_2170,In_364,In_1154);
or U2171 (N_2171,In_336,In_280);
xor U2172 (N_2172,In_1205,In_1180);
and U2173 (N_2173,In_1254,In_638);
xnor U2174 (N_2174,In_1153,In_113);
nand U2175 (N_2175,In_980,In_1437);
and U2176 (N_2176,In_1240,In_1212);
or U2177 (N_2177,In_728,In_773);
nor U2178 (N_2178,In_476,In_600);
nor U2179 (N_2179,In_620,In_1221);
nor U2180 (N_2180,In_529,In_26);
nor U2181 (N_2181,In_131,In_1148);
nand U2182 (N_2182,In_1252,In_896);
xnor U2183 (N_2183,In_213,In_1460);
or U2184 (N_2184,In_988,In_1233);
or U2185 (N_2185,In_120,In_850);
nor U2186 (N_2186,In_582,In_1222);
nand U2187 (N_2187,In_699,In_522);
nor U2188 (N_2188,In_1070,In_52);
nor U2189 (N_2189,In_583,In_973);
nor U2190 (N_2190,In_859,In_871);
nor U2191 (N_2191,In_484,In_358);
nor U2192 (N_2192,In_1037,In_1035);
nor U2193 (N_2193,In_52,In_73);
or U2194 (N_2194,In_564,In_1055);
nor U2195 (N_2195,In_468,In_156);
or U2196 (N_2196,In_205,In_217);
and U2197 (N_2197,In_1310,In_328);
nor U2198 (N_2198,In_805,In_1005);
or U2199 (N_2199,In_431,In_405);
nor U2200 (N_2200,In_74,In_902);
and U2201 (N_2201,In_886,In_1334);
and U2202 (N_2202,In_211,In_1041);
nand U2203 (N_2203,In_370,In_1289);
nand U2204 (N_2204,In_39,In_1039);
xor U2205 (N_2205,In_383,In_1195);
nor U2206 (N_2206,In_205,In_592);
and U2207 (N_2207,In_631,In_417);
nor U2208 (N_2208,In_689,In_1207);
xnor U2209 (N_2209,In_1388,In_398);
or U2210 (N_2210,In_1331,In_797);
or U2211 (N_2211,In_98,In_782);
nor U2212 (N_2212,In_761,In_1293);
or U2213 (N_2213,In_568,In_223);
nand U2214 (N_2214,In_1366,In_183);
nand U2215 (N_2215,In_485,In_749);
or U2216 (N_2216,In_1121,In_1450);
and U2217 (N_2217,In_403,In_110);
xnor U2218 (N_2218,In_75,In_468);
nor U2219 (N_2219,In_1259,In_458);
nor U2220 (N_2220,In_787,In_911);
and U2221 (N_2221,In_1236,In_177);
nand U2222 (N_2222,In_1301,In_888);
nor U2223 (N_2223,In_592,In_1381);
nand U2224 (N_2224,In_30,In_742);
and U2225 (N_2225,In_1220,In_60);
or U2226 (N_2226,In_601,In_733);
or U2227 (N_2227,In_562,In_660);
nor U2228 (N_2228,In_1497,In_498);
or U2229 (N_2229,In_585,In_418);
nor U2230 (N_2230,In_139,In_301);
nor U2231 (N_2231,In_410,In_256);
nor U2232 (N_2232,In_749,In_1110);
nor U2233 (N_2233,In_1114,In_94);
nand U2234 (N_2234,In_341,In_342);
and U2235 (N_2235,In_676,In_1363);
nand U2236 (N_2236,In_335,In_492);
nand U2237 (N_2237,In_1098,In_421);
and U2238 (N_2238,In_1255,In_346);
nor U2239 (N_2239,In_127,In_1256);
nor U2240 (N_2240,In_1077,In_1177);
nand U2241 (N_2241,In_30,In_719);
and U2242 (N_2242,In_596,In_782);
nand U2243 (N_2243,In_713,In_1195);
nand U2244 (N_2244,In_401,In_306);
nand U2245 (N_2245,In_342,In_904);
nand U2246 (N_2246,In_135,In_304);
nand U2247 (N_2247,In_763,In_1002);
or U2248 (N_2248,In_103,In_52);
nand U2249 (N_2249,In_356,In_1417);
or U2250 (N_2250,In_120,In_1208);
and U2251 (N_2251,In_513,In_1252);
nand U2252 (N_2252,In_262,In_23);
and U2253 (N_2253,In_104,In_1139);
nand U2254 (N_2254,In_720,In_1415);
nor U2255 (N_2255,In_195,In_1432);
or U2256 (N_2256,In_238,In_114);
xor U2257 (N_2257,In_1433,In_1405);
nor U2258 (N_2258,In_1477,In_1028);
and U2259 (N_2259,In_724,In_1407);
nand U2260 (N_2260,In_281,In_411);
or U2261 (N_2261,In_481,In_1321);
nand U2262 (N_2262,In_1264,In_583);
nor U2263 (N_2263,In_423,In_338);
and U2264 (N_2264,In_712,In_760);
and U2265 (N_2265,In_1393,In_390);
nor U2266 (N_2266,In_619,In_1326);
or U2267 (N_2267,In_497,In_139);
or U2268 (N_2268,In_1000,In_638);
nand U2269 (N_2269,In_664,In_765);
xnor U2270 (N_2270,In_359,In_1093);
nor U2271 (N_2271,In_1476,In_167);
and U2272 (N_2272,In_1096,In_636);
nand U2273 (N_2273,In_698,In_887);
nor U2274 (N_2274,In_1174,In_703);
nor U2275 (N_2275,In_825,In_126);
and U2276 (N_2276,In_92,In_1199);
nor U2277 (N_2277,In_1172,In_985);
or U2278 (N_2278,In_1003,In_1100);
and U2279 (N_2279,In_19,In_675);
nor U2280 (N_2280,In_647,In_256);
xnor U2281 (N_2281,In_302,In_430);
or U2282 (N_2282,In_1307,In_1449);
or U2283 (N_2283,In_588,In_1188);
nand U2284 (N_2284,In_1044,In_660);
nor U2285 (N_2285,In_1371,In_526);
or U2286 (N_2286,In_1239,In_587);
nand U2287 (N_2287,In_373,In_1075);
nor U2288 (N_2288,In_330,In_488);
and U2289 (N_2289,In_881,In_424);
nor U2290 (N_2290,In_618,In_621);
or U2291 (N_2291,In_571,In_885);
nor U2292 (N_2292,In_1008,In_1408);
nor U2293 (N_2293,In_755,In_287);
nand U2294 (N_2294,In_227,In_1265);
nor U2295 (N_2295,In_18,In_1350);
or U2296 (N_2296,In_214,In_581);
nor U2297 (N_2297,In_1051,In_525);
nand U2298 (N_2298,In_1393,In_1299);
or U2299 (N_2299,In_908,In_743);
nand U2300 (N_2300,In_665,In_162);
nor U2301 (N_2301,In_124,In_473);
nand U2302 (N_2302,In_325,In_230);
or U2303 (N_2303,In_80,In_164);
xnor U2304 (N_2304,In_751,In_144);
and U2305 (N_2305,In_220,In_830);
nand U2306 (N_2306,In_811,In_347);
xnor U2307 (N_2307,In_786,In_634);
nor U2308 (N_2308,In_1337,In_992);
or U2309 (N_2309,In_779,In_49);
and U2310 (N_2310,In_235,In_669);
nor U2311 (N_2311,In_506,In_42);
nand U2312 (N_2312,In_954,In_112);
nor U2313 (N_2313,In_20,In_1288);
and U2314 (N_2314,In_236,In_1159);
xor U2315 (N_2315,In_337,In_734);
xor U2316 (N_2316,In_232,In_537);
nor U2317 (N_2317,In_753,In_213);
nor U2318 (N_2318,In_1264,In_106);
nor U2319 (N_2319,In_581,In_1436);
xor U2320 (N_2320,In_888,In_377);
or U2321 (N_2321,In_197,In_1264);
or U2322 (N_2322,In_973,In_1072);
and U2323 (N_2323,In_477,In_356);
and U2324 (N_2324,In_221,In_1442);
nor U2325 (N_2325,In_1402,In_536);
xor U2326 (N_2326,In_698,In_536);
or U2327 (N_2327,In_493,In_628);
xor U2328 (N_2328,In_1405,In_401);
nand U2329 (N_2329,In_287,In_1347);
or U2330 (N_2330,In_63,In_1476);
or U2331 (N_2331,In_768,In_118);
xnor U2332 (N_2332,In_268,In_255);
or U2333 (N_2333,In_63,In_50);
and U2334 (N_2334,In_922,In_246);
nor U2335 (N_2335,In_655,In_1073);
xnor U2336 (N_2336,In_335,In_76);
or U2337 (N_2337,In_1038,In_154);
or U2338 (N_2338,In_1026,In_822);
nand U2339 (N_2339,In_1069,In_1001);
and U2340 (N_2340,In_719,In_366);
and U2341 (N_2341,In_559,In_807);
and U2342 (N_2342,In_1086,In_698);
xor U2343 (N_2343,In_1048,In_860);
nand U2344 (N_2344,In_1247,In_853);
and U2345 (N_2345,In_832,In_1022);
nand U2346 (N_2346,In_172,In_513);
nor U2347 (N_2347,In_1237,In_460);
nand U2348 (N_2348,In_326,In_354);
and U2349 (N_2349,In_151,In_572);
nand U2350 (N_2350,In_25,In_1453);
xnor U2351 (N_2351,In_1031,In_279);
or U2352 (N_2352,In_55,In_779);
nor U2353 (N_2353,In_286,In_67);
nor U2354 (N_2354,In_605,In_380);
nor U2355 (N_2355,In_1131,In_170);
xor U2356 (N_2356,In_987,In_335);
and U2357 (N_2357,In_470,In_1102);
nand U2358 (N_2358,In_1403,In_541);
nand U2359 (N_2359,In_1362,In_873);
or U2360 (N_2360,In_1031,In_770);
and U2361 (N_2361,In_426,In_245);
nand U2362 (N_2362,In_8,In_1282);
and U2363 (N_2363,In_83,In_1015);
nor U2364 (N_2364,In_210,In_504);
xor U2365 (N_2365,In_974,In_465);
and U2366 (N_2366,In_350,In_1041);
and U2367 (N_2367,In_1434,In_1486);
and U2368 (N_2368,In_1435,In_1310);
nor U2369 (N_2369,In_56,In_602);
nand U2370 (N_2370,In_801,In_244);
xnor U2371 (N_2371,In_1159,In_726);
nand U2372 (N_2372,In_445,In_835);
nor U2373 (N_2373,In_1474,In_105);
nand U2374 (N_2374,In_1467,In_1429);
and U2375 (N_2375,In_74,In_854);
nand U2376 (N_2376,In_328,In_578);
nor U2377 (N_2377,In_364,In_598);
and U2378 (N_2378,In_253,In_809);
or U2379 (N_2379,In_1335,In_354);
nand U2380 (N_2380,In_1118,In_1454);
and U2381 (N_2381,In_662,In_756);
nor U2382 (N_2382,In_839,In_409);
xnor U2383 (N_2383,In_1329,In_940);
nor U2384 (N_2384,In_1234,In_1093);
xor U2385 (N_2385,In_681,In_1429);
and U2386 (N_2386,In_214,In_869);
or U2387 (N_2387,In_446,In_1223);
or U2388 (N_2388,In_458,In_1235);
or U2389 (N_2389,In_590,In_300);
nor U2390 (N_2390,In_412,In_1003);
or U2391 (N_2391,In_309,In_508);
or U2392 (N_2392,In_208,In_81);
nand U2393 (N_2393,In_344,In_181);
nand U2394 (N_2394,In_487,In_1101);
and U2395 (N_2395,In_1122,In_396);
nor U2396 (N_2396,In_1353,In_870);
or U2397 (N_2397,In_1044,In_1481);
or U2398 (N_2398,In_1015,In_1496);
or U2399 (N_2399,In_1005,In_849);
and U2400 (N_2400,In_167,In_1361);
and U2401 (N_2401,In_183,In_63);
or U2402 (N_2402,In_1394,In_609);
and U2403 (N_2403,In_1306,In_700);
and U2404 (N_2404,In_395,In_63);
or U2405 (N_2405,In_900,In_380);
and U2406 (N_2406,In_407,In_951);
and U2407 (N_2407,In_230,In_327);
nor U2408 (N_2408,In_638,In_304);
xnor U2409 (N_2409,In_187,In_112);
or U2410 (N_2410,In_804,In_1366);
and U2411 (N_2411,In_302,In_355);
or U2412 (N_2412,In_804,In_271);
nand U2413 (N_2413,In_345,In_178);
nand U2414 (N_2414,In_1244,In_1296);
or U2415 (N_2415,In_1057,In_1109);
nor U2416 (N_2416,In_49,In_1218);
nor U2417 (N_2417,In_1478,In_1167);
and U2418 (N_2418,In_68,In_983);
or U2419 (N_2419,In_807,In_100);
and U2420 (N_2420,In_453,In_1148);
and U2421 (N_2421,In_432,In_156);
or U2422 (N_2422,In_1200,In_117);
nor U2423 (N_2423,In_1252,In_1125);
or U2424 (N_2424,In_616,In_1035);
or U2425 (N_2425,In_935,In_253);
and U2426 (N_2426,In_1012,In_1037);
and U2427 (N_2427,In_624,In_50);
nand U2428 (N_2428,In_1392,In_546);
nor U2429 (N_2429,In_402,In_525);
nor U2430 (N_2430,In_1113,In_104);
nor U2431 (N_2431,In_1183,In_1481);
nor U2432 (N_2432,In_1418,In_1438);
nand U2433 (N_2433,In_1215,In_966);
or U2434 (N_2434,In_1289,In_1328);
nor U2435 (N_2435,In_886,In_148);
and U2436 (N_2436,In_1142,In_117);
nand U2437 (N_2437,In_1418,In_719);
nand U2438 (N_2438,In_1236,In_1211);
or U2439 (N_2439,In_279,In_1376);
or U2440 (N_2440,In_1200,In_931);
and U2441 (N_2441,In_560,In_1043);
nor U2442 (N_2442,In_944,In_1301);
and U2443 (N_2443,In_161,In_1344);
or U2444 (N_2444,In_39,In_1444);
or U2445 (N_2445,In_275,In_649);
and U2446 (N_2446,In_100,In_538);
nand U2447 (N_2447,In_448,In_1428);
and U2448 (N_2448,In_1276,In_742);
and U2449 (N_2449,In_713,In_488);
xor U2450 (N_2450,In_603,In_186);
and U2451 (N_2451,In_1162,In_672);
nand U2452 (N_2452,In_764,In_1336);
nor U2453 (N_2453,In_1471,In_288);
or U2454 (N_2454,In_867,In_1212);
and U2455 (N_2455,In_54,In_275);
nor U2456 (N_2456,In_1343,In_818);
or U2457 (N_2457,In_1427,In_1357);
and U2458 (N_2458,In_497,In_423);
or U2459 (N_2459,In_1239,In_674);
nor U2460 (N_2460,In_291,In_38);
nand U2461 (N_2461,In_1147,In_746);
or U2462 (N_2462,In_1226,In_189);
nor U2463 (N_2463,In_564,In_1339);
and U2464 (N_2464,In_712,In_1233);
nand U2465 (N_2465,In_967,In_1023);
nand U2466 (N_2466,In_1406,In_1106);
xor U2467 (N_2467,In_604,In_1412);
nor U2468 (N_2468,In_290,In_1230);
and U2469 (N_2469,In_98,In_140);
nor U2470 (N_2470,In_1062,In_264);
nand U2471 (N_2471,In_52,In_1049);
xnor U2472 (N_2472,In_1092,In_776);
and U2473 (N_2473,In_1488,In_810);
and U2474 (N_2474,In_214,In_157);
nor U2475 (N_2475,In_675,In_762);
or U2476 (N_2476,In_106,In_858);
nand U2477 (N_2477,In_553,In_1427);
nor U2478 (N_2478,In_494,In_863);
and U2479 (N_2479,In_932,In_1087);
and U2480 (N_2480,In_502,In_879);
or U2481 (N_2481,In_1278,In_248);
nor U2482 (N_2482,In_191,In_1405);
or U2483 (N_2483,In_811,In_601);
and U2484 (N_2484,In_248,In_437);
nor U2485 (N_2485,In_173,In_518);
xnor U2486 (N_2486,In_1143,In_38);
nand U2487 (N_2487,In_673,In_417);
and U2488 (N_2488,In_1374,In_200);
nor U2489 (N_2489,In_695,In_1042);
xnor U2490 (N_2490,In_710,In_1202);
nor U2491 (N_2491,In_641,In_735);
or U2492 (N_2492,In_1172,In_184);
or U2493 (N_2493,In_1055,In_53);
nor U2494 (N_2494,In_675,In_453);
or U2495 (N_2495,In_1,In_135);
xnor U2496 (N_2496,In_1137,In_1050);
nor U2497 (N_2497,In_869,In_4);
nand U2498 (N_2498,In_998,In_721);
xor U2499 (N_2499,In_200,In_853);
nor U2500 (N_2500,In_311,In_1426);
xnor U2501 (N_2501,In_140,In_1307);
nor U2502 (N_2502,In_609,In_379);
xnor U2503 (N_2503,In_1157,In_736);
or U2504 (N_2504,In_415,In_1108);
nor U2505 (N_2505,In_85,In_1283);
nor U2506 (N_2506,In_893,In_107);
nor U2507 (N_2507,In_394,In_128);
nor U2508 (N_2508,In_836,In_1234);
nor U2509 (N_2509,In_65,In_135);
and U2510 (N_2510,In_617,In_901);
or U2511 (N_2511,In_272,In_1253);
or U2512 (N_2512,In_1270,In_1063);
or U2513 (N_2513,In_205,In_820);
and U2514 (N_2514,In_198,In_519);
nor U2515 (N_2515,In_478,In_396);
and U2516 (N_2516,In_298,In_1242);
nand U2517 (N_2517,In_769,In_1356);
xnor U2518 (N_2518,In_336,In_1137);
and U2519 (N_2519,In_652,In_1397);
nor U2520 (N_2520,In_8,In_354);
or U2521 (N_2521,In_521,In_516);
xor U2522 (N_2522,In_310,In_913);
xnor U2523 (N_2523,In_49,In_65);
or U2524 (N_2524,In_314,In_869);
nor U2525 (N_2525,In_38,In_90);
nand U2526 (N_2526,In_499,In_701);
nor U2527 (N_2527,In_1145,In_163);
nand U2528 (N_2528,In_296,In_592);
and U2529 (N_2529,In_258,In_1343);
or U2530 (N_2530,In_1386,In_175);
xnor U2531 (N_2531,In_1384,In_1387);
and U2532 (N_2532,In_624,In_347);
or U2533 (N_2533,In_1369,In_1420);
nor U2534 (N_2534,In_1114,In_1041);
and U2535 (N_2535,In_885,In_1267);
nand U2536 (N_2536,In_854,In_1101);
and U2537 (N_2537,In_467,In_248);
or U2538 (N_2538,In_453,In_227);
or U2539 (N_2539,In_885,In_556);
nand U2540 (N_2540,In_625,In_78);
and U2541 (N_2541,In_287,In_72);
or U2542 (N_2542,In_764,In_1102);
nor U2543 (N_2543,In_946,In_708);
or U2544 (N_2544,In_1054,In_126);
nor U2545 (N_2545,In_584,In_883);
nand U2546 (N_2546,In_784,In_664);
or U2547 (N_2547,In_44,In_1240);
nand U2548 (N_2548,In_900,In_343);
and U2549 (N_2549,In_931,In_766);
nand U2550 (N_2550,In_17,In_239);
and U2551 (N_2551,In_215,In_918);
xnor U2552 (N_2552,In_481,In_1083);
and U2553 (N_2553,In_170,In_630);
nor U2554 (N_2554,In_399,In_527);
and U2555 (N_2555,In_1312,In_456);
nor U2556 (N_2556,In_741,In_387);
or U2557 (N_2557,In_280,In_1080);
and U2558 (N_2558,In_397,In_724);
and U2559 (N_2559,In_17,In_271);
nand U2560 (N_2560,In_713,In_936);
and U2561 (N_2561,In_292,In_597);
and U2562 (N_2562,In_212,In_880);
nand U2563 (N_2563,In_940,In_665);
nor U2564 (N_2564,In_423,In_175);
nand U2565 (N_2565,In_731,In_859);
xor U2566 (N_2566,In_426,In_1023);
or U2567 (N_2567,In_355,In_498);
or U2568 (N_2568,In_12,In_1086);
and U2569 (N_2569,In_750,In_507);
or U2570 (N_2570,In_1343,In_861);
and U2571 (N_2571,In_793,In_1164);
or U2572 (N_2572,In_1222,In_1074);
nand U2573 (N_2573,In_71,In_1421);
and U2574 (N_2574,In_1065,In_1218);
nor U2575 (N_2575,In_702,In_147);
and U2576 (N_2576,In_1115,In_128);
or U2577 (N_2577,In_52,In_1246);
xnor U2578 (N_2578,In_575,In_775);
or U2579 (N_2579,In_639,In_1343);
nor U2580 (N_2580,In_219,In_591);
and U2581 (N_2581,In_847,In_395);
or U2582 (N_2582,In_153,In_327);
nor U2583 (N_2583,In_187,In_843);
nor U2584 (N_2584,In_231,In_1425);
or U2585 (N_2585,In_158,In_795);
nor U2586 (N_2586,In_529,In_133);
and U2587 (N_2587,In_156,In_444);
and U2588 (N_2588,In_226,In_1258);
nand U2589 (N_2589,In_1408,In_432);
and U2590 (N_2590,In_1487,In_334);
and U2591 (N_2591,In_154,In_1436);
nand U2592 (N_2592,In_652,In_1012);
xnor U2593 (N_2593,In_122,In_1467);
nand U2594 (N_2594,In_893,In_1211);
nor U2595 (N_2595,In_208,In_971);
and U2596 (N_2596,In_149,In_300);
or U2597 (N_2597,In_1265,In_973);
or U2598 (N_2598,In_1389,In_1217);
xnor U2599 (N_2599,In_883,In_1243);
nor U2600 (N_2600,In_493,In_1031);
or U2601 (N_2601,In_692,In_77);
nand U2602 (N_2602,In_1173,In_211);
nand U2603 (N_2603,In_704,In_147);
xnor U2604 (N_2604,In_485,In_987);
nor U2605 (N_2605,In_499,In_1251);
or U2606 (N_2606,In_915,In_1209);
nor U2607 (N_2607,In_1004,In_207);
nor U2608 (N_2608,In_581,In_982);
nor U2609 (N_2609,In_1362,In_1012);
or U2610 (N_2610,In_197,In_13);
nor U2611 (N_2611,In_57,In_36);
nor U2612 (N_2612,In_796,In_585);
nor U2613 (N_2613,In_1289,In_171);
nand U2614 (N_2614,In_691,In_947);
xor U2615 (N_2615,In_33,In_694);
nor U2616 (N_2616,In_663,In_564);
nand U2617 (N_2617,In_1121,In_389);
nand U2618 (N_2618,In_697,In_1345);
nor U2619 (N_2619,In_96,In_774);
and U2620 (N_2620,In_1323,In_853);
xor U2621 (N_2621,In_878,In_993);
nor U2622 (N_2622,In_662,In_377);
nand U2623 (N_2623,In_792,In_221);
or U2624 (N_2624,In_1497,In_778);
nand U2625 (N_2625,In_878,In_1333);
xor U2626 (N_2626,In_833,In_466);
nand U2627 (N_2627,In_335,In_1495);
and U2628 (N_2628,In_493,In_1019);
nand U2629 (N_2629,In_763,In_399);
nor U2630 (N_2630,In_1182,In_1084);
or U2631 (N_2631,In_1447,In_1007);
and U2632 (N_2632,In_1104,In_1266);
or U2633 (N_2633,In_1076,In_1248);
and U2634 (N_2634,In_134,In_949);
nor U2635 (N_2635,In_435,In_1219);
nand U2636 (N_2636,In_687,In_711);
and U2637 (N_2637,In_1071,In_1017);
nor U2638 (N_2638,In_1340,In_585);
or U2639 (N_2639,In_354,In_77);
nand U2640 (N_2640,In_730,In_1178);
nand U2641 (N_2641,In_1425,In_1095);
or U2642 (N_2642,In_784,In_1450);
xnor U2643 (N_2643,In_662,In_956);
and U2644 (N_2644,In_1468,In_138);
nor U2645 (N_2645,In_375,In_1324);
or U2646 (N_2646,In_822,In_789);
nand U2647 (N_2647,In_1074,In_212);
or U2648 (N_2648,In_1123,In_718);
nand U2649 (N_2649,In_1384,In_656);
xor U2650 (N_2650,In_769,In_1097);
and U2651 (N_2651,In_803,In_731);
or U2652 (N_2652,In_1232,In_542);
xor U2653 (N_2653,In_1096,In_785);
nand U2654 (N_2654,In_1451,In_1446);
and U2655 (N_2655,In_1326,In_605);
and U2656 (N_2656,In_1016,In_390);
nand U2657 (N_2657,In_791,In_23);
and U2658 (N_2658,In_415,In_1444);
or U2659 (N_2659,In_40,In_1453);
nand U2660 (N_2660,In_564,In_78);
or U2661 (N_2661,In_418,In_503);
nand U2662 (N_2662,In_134,In_1044);
nor U2663 (N_2663,In_515,In_367);
and U2664 (N_2664,In_1261,In_1477);
nor U2665 (N_2665,In_476,In_235);
or U2666 (N_2666,In_1394,In_409);
and U2667 (N_2667,In_915,In_172);
nor U2668 (N_2668,In_132,In_1424);
nand U2669 (N_2669,In_551,In_1011);
or U2670 (N_2670,In_1494,In_32);
and U2671 (N_2671,In_351,In_1288);
nand U2672 (N_2672,In_790,In_1491);
nand U2673 (N_2673,In_320,In_383);
xnor U2674 (N_2674,In_331,In_662);
and U2675 (N_2675,In_209,In_1402);
and U2676 (N_2676,In_1115,In_1415);
nand U2677 (N_2677,In_90,In_1230);
nand U2678 (N_2678,In_996,In_183);
nand U2679 (N_2679,In_594,In_1080);
and U2680 (N_2680,In_91,In_287);
nor U2681 (N_2681,In_220,In_367);
and U2682 (N_2682,In_1064,In_386);
and U2683 (N_2683,In_265,In_126);
nand U2684 (N_2684,In_248,In_882);
nor U2685 (N_2685,In_429,In_608);
and U2686 (N_2686,In_705,In_247);
xnor U2687 (N_2687,In_1123,In_56);
or U2688 (N_2688,In_1005,In_652);
nor U2689 (N_2689,In_912,In_1240);
nor U2690 (N_2690,In_570,In_282);
nor U2691 (N_2691,In_243,In_4);
nand U2692 (N_2692,In_304,In_71);
and U2693 (N_2693,In_1120,In_79);
or U2694 (N_2694,In_789,In_1305);
and U2695 (N_2695,In_559,In_645);
and U2696 (N_2696,In_848,In_310);
and U2697 (N_2697,In_236,In_1303);
and U2698 (N_2698,In_1077,In_470);
nand U2699 (N_2699,In_1028,In_78);
or U2700 (N_2700,In_1276,In_861);
and U2701 (N_2701,In_337,In_148);
and U2702 (N_2702,In_906,In_1062);
or U2703 (N_2703,In_958,In_471);
or U2704 (N_2704,In_879,In_1357);
xor U2705 (N_2705,In_793,In_56);
or U2706 (N_2706,In_79,In_1087);
and U2707 (N_2707,In_1142,In_768);
nor U2708 (N_2708,In_1363,In_592);
nor U2709 (N_2709,In_649,In_720);
and U2710 (N_2710,In_1100,In_47);
nor U2711 (N_2711,In_548,In_1420);
nand U2712 (N_2712,In_359,In_708);
or U2713 (N_2713,In_1225,In_381);
or U2714 (N_2714,In_1330,In_418);
xnor U2715 (N_2715,In_321,In_295);
and U2716 (N_2716,In_229,In_882);
nand U2717 (N_2717,In_448,In_883);
nor U2718 (N_2718,In_1335,In_1049);
xor U2719 (N_2719,In_464,In_494);
and U2720 (N_2720,In_1265,In_1273);
nor U2721 (N_2721,In_1468,In_560);
or U2722 (N_2722,In_1310,In_559);
and U2723 (N_2723,In_441,In_1271);
or U2724 (N_2724,In_446,In_1240);
nor U2725 (N_2725,In_390,In_1319);
and U2726 (N_2726,In_794,In_1118);
nand U2727 (N_2727,In_1444,In_525);
and U2728 (N_2728,In_1148,In_477);
and U2729 (N_2729,In_43,In_127);
or U2730 (N_2730,In_1407,In_973);
xor U2731 (N_2731,In_954,In_980);
xnor U2732 (N_2732,In_948,In_1061);
xnor U2733 (N_2733,In_1232,In_1144);
xnor U2734 (N_2734,In_759,In_237);
or U2735 (N_2735,In_550,In_555);
and U2736 (N_2736,In_1326,In_143);
nor U2737 (N_2737,In_739,In_1407);
nor U2738 (N_2738,In_1447,In_1199);
or U2739 (N_2739,In_372,In_966);
nor U2740 (N_2740,In_853,In_1458);
and U2741 (N_2741,In_1159,In_131);
nand U2742 (N_2742,In_812,In_114);
nor U2743 (N_2743,In_542,In_1006);
and U2744 (N_2744,In_634,In_688);
nand U2745 (N_2745,In_955,In_826);
xnor U2746 (N_2746,In_1448,In_1337);
nand U2747 (N_2747,In_712,In_766);
and U2748 (N_2748,In_787,In_1268);
nand U2749 (N_2749,In_462,In_998);
nand U2750 (N_2750,In_989,In_1289);
or U2751 (N_2751,In_605,In_428);
nor U2752 (N_2752,In_316,In_1362);
nand U2753 (N_2753,In_534,In_975);
nand U2754 (N_2754,In_371,In_206);
nor U2755 (N_2755,In_1396,In_938);
and U2756 (N_2756,In_981,In_246);
nand U2757 (N_2757,In_886,In_59);
and U2758 (N_2758,In_1401,In_817);
or U2759 (N_2759,In_322,In_746);
nor U2760 (N_2760,In_1088,In_1408);
nand U2761 (N_2761,In_1208,In_17);
or U2762 (N_2762,In_349,In_1091);
nor U2763 (N_2763,In_649,In_851);
xor U2764 (N_2764,In_707,In_571);
xor U2765 (N_2765,In_615,In_510);
or U2766 (N_2766,In_154,In_1391);
xnor U2767 (N_2767,In_155,In_623);
nor U2768 (N_2768,In_947,In_1254);
nand U2769 (N_2769,In_522,In_232);
nor U2770 (N_2770,In_1047,In_1054);
xor U2771 (N_2771,In_649,In_316);
nand U2772 (N_2772,In_125,In_652);
nand U2773 (N_2773,In_265,In_1432);
nor U2774 (N_2774,In_1444,In_112);
nor U2775 (N_2775,In_371,In_1292);
or U2776 (N_2776,In_205,In_805);
nor U2777 (N_2777,In_485,In_29);
and U2778 (N_2778,In_620,In_635);
nor U2779 (N_2779,In_1352,In_321);
or U2780 (N_2780,In_448,In_1074);
nand U2781 (N_2781,In_161,In_1005);
nor U2782 (N_2782,In_1477,In_1134);
or U2783 (N_2783,In_510,In_428);
or U2784 (N_2784,In_1387,In_760);
and U2785 (N_2785,In_1147,In_419);
and U2786 (N_2786,In_704,In_1164);
or U2787 (N_2787,In_808,In_836);
and U2788 (N_2788,In_1227,In_1298);
nand U2789 (N_2789,In_99,In_1038);
nor U2790 (N_2790,In_565,In_350);
nand U2791 (N_2791,In_1445,In_659);
nand U2792 (N_2792,In_1297,In_653);
nor U2793 (N_2793,In_840,In_694);
nor U2794 (N_2794,In_1033,In_1207);
nand U2795 (N_2795,In_337,In_589);
or U2796 (N_2796,In_1155,In_332);
and U2797 (N_2797,In_1112,In_1320);
or U2798 (N_2798,In_572,In_1131);
nand U2799 (N_2799,In_690,In_888);
nand U2800 (N_2800,In_1422,In_726);
and U2801 (N_2801,In_309,In_400);
and U2802 (N_2802,In_112,In_26);
nand U2803 (N_2803,In_957,In_1201);
nor U2804 (N_2804,In_1379,In_31);
and U2805 (N_2805,In_1190,In_71);
nand U2806 (N_2806,In_704,In_903);
nand U2807 (N_2807,In_466,In_1110);
nor U2808 (N_2808,In_488,In_1313);
nor U2809 (N_2809,In_643,In_847);
and U2810 (N_2810,In_1276,In_1463);
or U2811 (N_2811,In_554,In_239);
or U2812 (N_2812,In_273,In_1226);
and U2813 (N_2813,In_516,In_1360);
or U2814 (N_2814,In_412,In_1499);
nand U2815 (N_2815,In_94,In_781);
nor U2816 (N_2816,In_1452,In_23);
or U2817 (N_2817,In_882,In_575);
or U2818 (N_2818,In_851,In_261);
xor U2819 (N_2819,In_786,In_1276);
nor U2820 (N_2820,In_1142,In_1259);
and U2821 (N_2821,In_984,In_965);
nor U2822 (N_2822,In_652,In_613);
and U2823 (N_2823,In_824,In_1225);
nand U2824 (N_2824,In_1438,In_1127);
nor U2825 (N_2825,In_729,In_154);
and U2826 (N_2826,In_1191,In_654);
nor U2827 (N_2827,In_1242,In_391);
and U2828 (N_2828,In_8,In_1173);
nand U2829 (N_2829,In_368,In_366);
xnor U2830 (N_2830,In_590,In_1033);
xnor U2831 (N_2831,In_788,In_1221);
nor U2832 (N_2832,In_921,In_1142);
or U2833 (N_2833,In_527,In_502);
or U2834 (N_2834,In_28,In_931);
and U2835 (N_2835,In_1344,In_844);
xnor U2836 (N_2836,In_565,In_449);
or U2837 (N_2837,In_1058,In_634);
nand U2838 (N_2838,In_933,In_1466);
nand U2839 (N_2839,In_368,In_103);
nand U2840 (N_2840,In_481,In_33);
or U2841 (N_2841,In_741,In_1309);
nor U2842 (N_2842,In_735,In_858);
and U2843 (N_2843,In_1439,In_1011);
nor U2844 (N_2844,In_60,In_1421);
nand U2845 (N_2845,In_1359,In_123);
or U2846 (N_2846,In_348,In_484);
and U2847 (N_2847,In_1472,In_306);
or U2848 (N_2848,In_234,In_271);
and U2849 (N_2849,In_1385,In_128);
nand U2850 (N_2850,In_682,In_1407);
or U2851 (N_2851,In_461,In_1065);
nor U2852 (N_2852,In_719,In_1360);
nor U2853 (N_2853,In_243,In_760);
nand U2854 (N_2854,In_645,In_348);
nor U2855 (N_2855,In_881,In_169);
nor U2856 (N_2856,In_535,In_112);
and U2857 (N_2857,In_1183,In_822);
or U2858 (N_2858,In_952,In_966);
nor U2859 (N_2859,In_996,In_603);
nor U2860 (N_2860,In_183,In_127);
or U2861 (N_2861,In_882,In_743);
or U2862 (N_2862,In_476,In_885);
xnor U2863 (N_2863,In_83,In_537);
nand U2864 (N_2864,In_799,In_902);
nand U2865 (N_2865,In_1000,In_633);
nor U2866 (N_2866,In_824,In_97);
or U2867 (N_2867,In_603,In_761);
nor U2868 (N_2868,In_1007,In_140);
xnor U2869 (N_2869,In_246,In_821);
and U2870 (N_2870,In_1132,In_1427);
nand U2871 (N_2871,In_1182,In_780);
xor U2872 (N_2872,In_721,In_1324);
nor U2873 (N_2873,In_1032,In_424);
and U2874 (N_2874,In_443,In_491);
nor U2875 (N_2875,In_1064,In_824);
and U2876 (N_2876,In_945,In_1306);
nor U2877 (N_2877,In_227,In_696);
xor U2878 (N_2878,In_1269,In_938);
xnor U2879 (N_2879,In_777,In_1255);
nor U2880 (N_2880,In_886,In_450);
and U2881 (N_2881,In_806,In_299);
xnor U2882 (N_2882,In_655,In_41);
nand U2883 (N_2883,In_1178,In_561);
nand U2884 (N_2884,In_305,In_1014);
and U2885 (N_2885,In_341,In_808);
nand U2886 (N_2886,In_494,In_1443);
nor U2887 (N_2887,In_1272,In_686);
nand U2888 (N_2888,In_492,In_83);
or U2889 (N_2889,In_1206,In_833);
and U2890 (N_2890,In_552,In_943);
nor U2891 (N_2891,In_291,In_1338);
or U2892 (N_2892,In_473,In_452);
nor U2893 (N_2893,In_263,In_592);
nand U2894 (N_2894,In_367,In_1111);
nor U2895 (N_2895,In_692,In_250);
and U2896 (N_2896,In_685,In_644);
nor U2897 (N_2897,In_1332,In_150);
nand U2898 (N_2898,In_403,In_22);
and U2899 (N_2899,In_1018,In_1029);
nand U2900 (N_2900,In_128,In_1103);
and U2901 (N_2901,In_437,In_522);
or U2902 (N_2902,In_203,In_261);
and U2903 (N_2903,In_121,In_15);
nor U2904 (N_2904,In_433,In_764);
or U2905 (N_2905,In_585,In_1007);
nand U2906 (N_2906,In_127,In_76);
xnor U2907 (N_2907,In_792,In_523);
nor U2908 (N_2908,In_932,In_809);
and U2909 (N_2909,In_267,In_409);
nand U2910 (N_2910,In_1013,In_310);
nor U2911 (N_2911,In_697,In_1211);
and U2912 (N_2912,In_647,In_5);
or U2913 (N_2913,In_127,In_195);
or U2914 (N_2914,In_482,In_71);
nand U2915 (N_2915,In_1098,In_567);
nand U2916 (N_2916,In_360,In_886);
nor U2917 (N_2917,In_769,In_1149);
or U2918 (N_2918,In_937,In_781);
or U2919 (N_2919,In_1002,In_1401);
nand U2920 (N_2920,In_586,In_344);
and U2921 (N_2921,In_1321,In_824);
nand U2922 (N_2922,In_557,In_592);
nand U2923 (N_2923,In_1038,In_1492);
and U2924 (N_2924,In_1299,In_980);
nor U2925 (N_2925,In_775,In_744);
xnor U2926 (N_2926,In_1009,In_104);
nand U2927 (N_2927,In_617,In_434);
or U2928 (N_2928,In_1333,In_1065);
and U2929 (N_2929,In_140,In_1164);
and U2930 (N_2930,In_231,In_563);
nand U2931 (N_2931,In_1110,In_1332);
or U2932 (N_2932,In_1337,In_165);
and U2933 (N_2933,In_881,In_495);
nor U2934 (N_2934,In_733,In_122);
or U2935 (N_2935,In_1361,In_554);
nor U2936 (N_2936,In_496,In_318);
or U2937 (N_2937,In_1463,In_1015);
or U2938 (N_2938,In_1341,In_209);
xor U2939 (N_2939,In_305,In_639);
nand U2940 (N_2940,In_315,In_1187);
nand U2941 (N_2941,In_1206,In_1237);
or U2942 (N_2942,In_509,In_1335);
or U2943 (N_2943,In_1195,In_259);
and U2944 (N_2944,In_587,In_921);
nor U2945 (N_2945,In_607,In_135);
xnor U2946 (N_2946,In_447,In_960);
nand U2947 (N_2947,In_1309,In_284);
nand U2948 (N_2948,In_380,In_887);
nor U2949 (N_2949,In_1143,In_892);
and U2950 (N_2950,In_290,In_626);
or U2951 (N_2951,In_584,In_351);
nor U2952 (N_2952,In_699,In_856);
nor U2953 (N_2953,In_182,In_846);
nor U2954 (N_2954,In_566,In_460);
or U2955 (N_2955,In_501,In_463);
nand U2956 (N_2956,In_293,In_181);
and U2957 (N_2957,In_1009,In_1258);
xnor U2958 (N_2958,In_152,In_231);
nor U2959 (N_2959,In_429,In_871);
nor U2960 (N_2960,In_1273,In_792);
and U2961 (N_2961,In_673,In_1142);
xor U2962 (N_2962,In_1269,In_432);
or U2963 (N_2963,In_308,In_1436);
or U2964 (N_2964,In_888,In_1204);
and U2965 (N_2965,In_168,In_1410);
nor U2966 (N_2966,In_918,In_190);
xnor U2967 (N_2967,In_553,In_982);
nand U2968 (N_2968,In_178,In_704);
nand U2969 (N_2969,In_1064,In_69);
or U2970 (N_2970,In_95,In_629);
nor U2971 (N_2971,In_244,In_574);
nand U2972 (N_2972,In_295,In_868);
nand U2973 (N_2973,In_1042,In_1399);
and U2974 (N_2974,In_663,In_362);
or U2975 (N_2975,In_164,In_442);
or U2976 (N_2976,In_992,In_786);
xor U2977 (N_2977,In_434,In_124);
or U2978 (N_2978,In_477,In_311);
or U2979 (N_2979,In_536,In_236);
and U2980 (N_2980,In_1460,In_1375);
nand U2981 (N_2981,In_890,In_71);
nand U2982 (N_2982,In_778,In_1449);
nand U2983 (N_2983,In_1099,In_466);
nor U2984 (N_2984,In_276,In_428);
nor U2985 (N_2985,In_986,In_285);
nand U2986 (N_2986,In_1200,In_360);
and U2987 (N_2987,In_603,In_590);
and U2988 (N_2988,In_1285,In_26);
or U2989 (N_2989,In_782,In_77);
or U2990 (N_2990,In_1091,In_807);
or U2991 (N_2991,In_478,In_690);
nand U2992 (N_2992,In_872,In_819);
and U2993 (N_2993,In_118,In_1287);
xnor U2994 (N_2994,In_1330,In_154);
and U2995 (N_2995,In_1217,In_1280);
and U2996 (N_2996,In_954,In_204);
and U2997 (N_2997,In_763,In_756);
nand U2998 (N_2998,In_735,In_471);
nand U2999 (N_2999,In_402,In_129);
or U3000 (N_3000,In_827,In_179);
or U3001 (N_3001,In_484,In_909);
or U3002 (N_3002,In_835,In_467);
nor U3003 (N_3003,In_939,In_940);
nor U3004 (N_3004,In_984,In_11);
or U3005 (N_3005,In_897,In_687);
and U3006 (N_3006,In_739,In_879);
nand U3007 (N_3007,In_163,In_1327);
nor U3008 (N_3008,In_750,In_908);
nand U3009 (N_3009,In_31,In_1102);
nor U3010 (N_3010,In_1025,In_133);
and U3011 (N_3011,In_40,In_585);
or U3012 (N_3012,In_1073,In_1168);
nand U3013 (N_3013,In_493,In_984);
or U3014 (N_3014,In_815,In_1068);
or U3015 (N_3015,In_397,In_1158);
and U3016 (N_3016,In_837,In_944);
and U3017 (N_3017,In_354,In_388);
xnor U3018 (N_3018,In_585,In_1227);
and U3019 (N_3019,In_772,In_773);
nand U3020 (N_3020,In_1243,In_541);
nand U3021 (N_3021,In_421,In_1397);
and U3022 (N_3022,In_567,In_20);
or U3023 (N_3023,In_338,In_487);
nor U3024 (N_3024,In_320,In_435);
nor U3025 (N_3025,In_1030,In_1343);
xnor U3026 (N_3026,In_447,In_494);
xor U3027 (N_3027,In_346,In_1400);
or U3028 (N_3028,In_406,In_1348);
nor U3029 (N_3029,In_1145,In_850);
and U3030 (N_3030,In_179,In_524);
nand U3031 (N_3031,In_62,In_262);
and U3032 (N_3032,In_410,In_1217);
or U3033 (N_3033,In_246,In_1260);
nor U3034 (N_3034,In_944,In_625);
nand U3035 (N_3035,In_1420,In_866);
nand U3036 (N_3036,In_122,In_1230);
and U3037 (N_3037,In_693,In_873);
nor U3038 (N_3038,In_93,In_1209);
nand U3039 (N_3039,In_479,In_530);
nor U3040 (N_3040,In_431,In_344);
and U3041 (N_3041,In_508,In_689);
or U3042 (N_3042,In_1164,In_863);
nor U3043 (N_3043,In_861,In_1169);
xor U3044 (N_3044,In_794,In_1275);
nand U3045 (N_3045,In_200,In_105);
nor U3046 (N_3046,In_621,In_1058);
nand U3047 (N_3047,In_261,In_1409);
and U3048 (N_3048,In_1151,In_344);
nand U3049 (N_3049,In_176,In_196);
nor U3050 (N_3050,In_1302,In_241);
or U3051 (N_3051,In_1255,In_662);
or U3052 (N_3052,In_71,In_1207);
nand U3053 (N_3053,In_891,In_691);
and U3054 (N_3054,In_722,In_1486);
or U3055 (N_3055,In_939,In_152);
and U3056 (N_3056,In_869,In_540);
or U3057 (N_3057,In_1186,In_1004);
and U3058 (N_3058,In_578,In_1345);
nor U3059 (N_3059,In_1348,In_374);
nor U3060 (N_3060,In_1143,In_424);
nand U3061 (N_3061,In_31,In_758);
nand U3062 (N_3062,In_131,In_371);
nor U3063 (N_3063,In_908,In_217);
or U3064 (N_3064,In_18,In_908);
nor U3065 (N_3065,In_485,In_763);
nand U3066 (N_3066,In_1465,In_424);
xnor U3067 (N_3067,In_243,In_178);
and U3068 (N_3068,In_432,In_475);
or U3069 (N_3069,In_1037,In_514);
or U3070 (N_3070,In_390,In_173);
or U3071 (N_3071,In_1036,In_311);
or U3072 (N_3072,In_714,In_1288);
or U3073 (N_3073,In_1150,In_1142);
and U3074 (N_3074,In_247,In_1076);
xnor U3075 (N_3075,In_76,In_826);
nor U3076 (N_3076,In_1464,In_508);
or U3077 (N_3077,In_899,In_1413);
nor U3078 (N_3078,In_170,In_1339);
and U3079 (N_3079,In_115,In_338);
and U3080 (N_3080,In_1101,In_751);
and U3081 (N_3081,In_921,In_794);
and U3082 (N_3082,In_683,In_1373);
nand U3083 (N_3083,In_1299,In_1219);
or U3084 (N_3084,In_93,In_240);
or U3085 (N_3085,In_125,In_923);
nand U3086 (N_3086,In_1091,In_190);
nand U3087 (N_3087,In_810,In_1063);
xor U3088 (N_3088,In_954,In_629);
or U3089 (N_3089,In_629,In_647);
nor U3090 (N_3090,In_1135,In_1116);
xnor U3091 (N_3091,In_1498,In_189);
nor U3092 (N_3092,In_122,In_305);
nor U3093 (N_3093,In_598,In_416);
or U3094 (N_3094,In_618,In_679);
nor U3095 (N_3095,In_743,In_483);
and U3096 (N_3096,In_100,In_640);
or U3097 (N_3097,In_3,In_1084);
and U3098 (N_3098,In_1317,In_1498);
nand U3099 (N_3099,In_1365,In_35);
and U3100 (N_3100,In_1110,In_65);
xnor U3101 (N_3101,In_193,In_1295);
or U3102 (N_3102,In_1306,In_950);
nand U3103 (N_3103,In_231,In_397);
or U3104 (N_3104,In_1354,In_803);
nand U3105 (N_3105,In_295,In_1149);
xnor U3106 (N_3106,In_894,In_955);
nand U3107 (N_3107,In_904,In_563);
nand U3108 (N_3108,In_783,In_954);
nand U3109 (N_3109,In_1462,In_8);
or U3110 (N_3110,In_309,In_359);
or U3111 (N_3111,In_5,In_1367);
nor U3112 (N_3112,In_605,In_767);
and U3113 (N_3113,In_1279,In_1274);
nand U3114 (N_3114,In_1340,In_128);
nand U3115 (N_3115,In_1259,In_208);
nand U3116 (N_3116,In_270,In_1126);
nand U3117 (N_3117,In_860,In_50);
and U3118 (N_3118,In_911,In_160);
xor U3119 (N_3119,In_1013,In_61);
nor U3120 (N_3120,In_531,In_1432);
and U3121 (N_3121,In_492,In_312);
nor U3122 (N_3122,In_682,In_114);
nand U3123 (N_3123,In_875,In_88);
nor U3124 (N_3124,In_224,In_662);
or U3125 (N_3125,In_603,In_245);
or U3126 (N_3126,In_485,In_617);
nor U3127 (N_3127,In_868,In_1025);
xnor U3128 (N_3128,In_393,In_722);
or U3129 (N_3129,In_556,In_60);
nor U3130 (N_3130,In_1419,In_595);
and U3131 (N_3131,In_1329,In_1064);
nand U3132 (N_3132,In_732,In_553);
or U3133 (N_3133,In_1132,In_571);
and U3134 (N_3134,In_1472,In_1196);
nand U3135 (N_3135,In_1106,In_633);
or U3136 (N_3136,In_404,In_757);
nand U3137 (N_3137,In_1381,In_1186);
or U3138 (N_3138,In_1037,In_416);
or U3139 (N_3139,In_476,In_1473);
xor U3140 (N_3140,In_581,In_559);
and U3141 (N_3141,In_791,In_1055);
nor U3142 (N_3142,In_1375,In_912);
nand U3143 (N_3143,In_1417,In_163);
or U3144 (N_3144,In_180,In_702);
xnor U3145 (N_3145,In_359,In_1236);
or U3146 (N_3146,In_1429,In_707);
and U3147 (N_3147,In_218,In_289);
nor U3148 (N_3148,In_392,In_23);
nand U3149 (N_3149,In_159,In_688);
nand U3150 (N_3150,In_596,In_1401);
nand U3151 (N_3151,In_661,In_47);
and U3152 (N_3152,In_705,In_735);
or U3153 (N_3153,In_75,In_1028);
xnor U3154 (N_3154,In_465,In_1490);
nor U3155 (N_3155,In_733,In_361);
and U3156 (N_3156,In_325,In_1456);
nand U3157 (N_3157,In_938,In_766);
xnor U3158 (N_3158,In_547,In_137);
xnor U3159 (N_3159,In_684,In_757);
nand U3160 (N_3160,In_1111,In_1462);
nand U3161 (N_3161,In_694,In_1499);
xor U3162 (N_3162,In_545,In_228);
or U3163 (N_3163,In_176,In_939);
nand U3164 (N_3164,In_1378,In_43);
nand U3165 (N_3165,In_800,In_194);
nand U3166 (N_3166,In_599,In_690);
or U3167 (N_3167,In_23,In_733);
xor U3168 (N_3168,In_1233,In_786);
nand U3169 (N_3169,In_769,In_1074);
or U3170 (N_3170,In_53,In_157);
nand U3171 (N_3171,In_1075,In_268);
nand U3172 (N_3172,In_472,In_211);
nor U3173 (N_3173,In_71,In_212);
nand U3174 (N_3174,In_1242,In_250);
xor U3175 (N_3175,In_931,In_426);
or U3176 (N_3176,In_610,In_1381);
or U3177 (N_3177,In_849,In_1460);
or U3178 (N_3178,In_737,In_1082);
and U3179 (N_3179,In_807,In_182);
or U3180 (N_3180,In_952,In_546);
and U3181 (N_3181,In_1288,In_203);
nor U3182 (N_3182,In_877,In_72);
nand U3183 (N_3183,In_329,In_820);
and U3184 (N_3184,In_706,In_1496);
xor U3185 (N_3185,In_1234,In_287);
or U3186 (N_3186,In_648,In_721);
and U3187 (N_3187,In_572,In_1247);
nor U3188 (N_3188,In_783,In_1414);
nor U3189 (N_3189,In_1126,In_1352);
nand U3190 (N_3190,In_556,In_405);
and U3191 (N_3191,In_960,In_1364);
nand U3192 (N_3192,In_559,In_710);
nand U3193 (N_3193,In_943,In_736);
and U3194 (N_3194,In_120,In_867);
or U3195 (N_3195,In_671,In_1189);
xor U3196 (N_3196,In_82,In_845);
xnor U3197 (N_3197,In_1418,In_347);
or U3198 (N_3198,In_377,In_459);
nand U3199 (N_3199,In_917,In_1216);
and U3200 (N_3200,In_972,In_844);
nand U3201 (N_3201,In_1250,In_87);
nand U3202 (N_3202,In_636,In_962);
or U3203 (N_3203,In_514,In_559);
and U3204 (N_3204,In_82,In_178);
nor U3205 (N_3205,In_802,In_417);
nor U3206 (N_3206,In_1330,In_1269);
nand U3207 (N_3207,In_1308,In_174);
and U3208 (N_3208,In_604,In_1150);
nor U3209 (N_3209,In_634,In_410);
or U3210 (N_3210,In_797,In_887);
or U3211 (N_3211,In_556,In_253);
or U3212 (N_3212,In_283,In_570);
nor U3213 (N_3213,In_450,In_53);
xnor U3214 (N_3214,In_1167,In_599);
or U3215 (N_3215,In_552,In_992);
or U3216 (N_3216,In_1020,In_1271);
or U3217 (N_3217,In_503,In_206);
nor U3218 (N_3218,In_1494,In_1026);
nor U3219 (N_3219,In_277,In_1282);
nor U3220 (N_3220,In_1002,In_259);
or U3221 (N_3221,In_1189,In_0);
and U3222 (N_3222,In_837,In_1264);
nor U3223 (N_3223,In_1016,In_509);
and U3224 (N_3224,In_509,In_523);
or U3225 (N_3225,In_473,In_363);
or U3226 (N_3226,In_1326,In_513);
xnor U3227 (N_3227,In_802,In_584);
and U3228 (N_3228,In_1225,In_401);
or U3229 (N_3229,In_965,In_1240);
xnor U3230 (N_3230,In_105,In_517);
xnor U3231 (N_3231,In_869,In_1334);
and U3232 (N_3232,In_863,In_835);
or U3233 (N_3233,In_878,In_1468);
nor U3234 (N_3234,In_530,In_703);
nor U3235 (N_3235,In_875,In_1114);
and U3236 (N_3236,In_1348,In_950);
or U3237 (N_3237,In_950,In_606);
or U3238 (N_3238,In_1472,In_532);
and U3239 (N_3239,In_0,In_1151);
and U3240 (N_3240,In_1429,In_359);
nand U3241 (N_3241,In_18,In_1257);
or U3242 (N_3242,In_1434,In_1074);
or U3243 (N_3243,In_1144,In_1369);
and U3244 (N_3244,In_71,In_822);
and U3245 (N_3245,In_783,In_793);
xor U3246 (N_3246,In_65,In_616);
nand U3247 (N_3247,In_395,In_69);
and U3248 (N_3248,In_1111,In_631);
or U3249 (N_3249,In_931,In_795);
or U3250 (N_3250,In_130,In_376);
xor U3251 (N_3251,In_1110,In_578);
nand U3252 (N_3252,In_2,In_200);
xnor U3253 (N_3253,In_1185,In_314);
nand U3254 (N_3254,In_778,In_1473);
nand U3255 (N_3255,In_174,In_661);
nand U3256 (N_3256,In_541,In_1111);
nor U3257 (N_3257,In_969,In_835);
nor U3258 (N_3258,In_416,In_888);
nor U3259 (N_3259,In_955,In_215);
nor U3260 (N_3260,In_324,In_114);
xnor U3261 (N_3261,In_884,In_631);
nor U3262 (N_3262,In_585,In_205);
nand U3263 (N_3263,In_1026,In_779);
and U3264 (N_3264,In_1402,In_1106);
nor U3265 (N_3265,In_124,In_1414);
nand U3266 (N_3266,In_1067,In_18);
nor U3267 (N_3267,In_494,In_317);
and U3268 (N_3268,In_608,In_873);
nand U3269 (N_3269,In_736,In_505);
nor U3270 (N_3270,In_17,In_778);
and U3271 (N_3271,In_581,In_539);
nor U3272 (N_3272,In_675,In_1219);
nand U3273 (N_3273,In_212,In_1293);
or U3274 (N_3274,In_681,In_752);
or U3275 (N_3275,In_704,In_792);
xor U3276 (N_3276,In_459,In_208);
and U3277 (N_3277,In_339,In_13);
and U3278 (N_3278,In_1414,In_1335);
or U3279 (N_3279,In_81,In_818);
nand U3280 (N_3280,In_759,In_28);
or U3281 (N_3281,In_1295,In_459);
nor U3282 (N_3282,In_968,In_996);
nand U3283 (N_3283,In_313,In_667);
nand U3284 (N_3284,In_329,In_894);
nand U3285 (N_3285,In_595,In_921);
or U3286 (N_3286,In_1139,In_1197);
and U3287 (N_3287,In_1303,In_38);
nand U3288 (N_3288,In_218,In_587);
or U3289 (N_3289,In_462,In_980);
xor U3290 (N_3290,In_1032,In_794);
or U3291 (N_3291,In_333,In_140);
nor U3292 (N_3292,In_1080,In_1069);
nor U3293 (N_3293,In_1455,In_498);
nor U3294 (N_3294,In_398,In_1038);
xnor U3295 (N_3295,In_1409,In_653);
and U3296 (N_3296,In_117,In_1292);
or U3297 (N_3297,In_1072,In_1025);
nor U3298 (N_3298,In_82,In_1244);
nand U3299 (N_3299,In_1025,In_405);
and U3300 (N_3300,In_303,In_56);
or U3301 (N_3301,In_479,In_576);
nor U3302 (N_3302,In_187,In_639);
nand U3303 (N_3303,In_1346,In_434);
or U3304 (N_3304,In_591,In_672);
nor U3305 (N_3305,In_569,In_854);
or U3306 (N_3306,In_366,In_82);
and U3307 (N_3307,In_1439,In_8);
and U3308 (N_3308,In_1483,In_1136);
xor U3309 (N_3309,In_53,In_214);
nor U3310 (N_3310,In_693,In_928);
and U3311 (N_3311,In_1065,In_1456);
and U3312 (N_3312,In_782,In_1181);
nor U3313 (N_3313,In_1277,In_166);
and U3314 (N_3314,In_694,In_885);
or U3315 (N_3315,In_801,In_110);
and U3316 (N_3316,In_906,In_1154);
or U3317 (N_3317,In_829,In_490);
nand U3318 (N_3318,In_453,In_1173);
nand U3319 (N_3319,In_581,In_574);
or U3320 (N_3320,In_667,In_458);
nand U3321 (N_3321,In_39,In_1372);
or U3322 (N_3322,In_676,In_770);
nor U3323 (N_3323,In_1189,In_387);
or U3324 (N_3324,In_548,In_590);
nor U3325 (N_3325,In_117,In_1348);
or U3326 (N_3326,In_409,In_1007);
or U3327 (N_3327,In_772,In_480);
or U3328 (N_3328,In_894,In_170);
xor U3329 (N_3329,In_1104,In_559);
and U3330 (N_3330,In_773,In_79);
and U3331 (N_3331,In_1153,In_1015);
xor U3332 (N_3332,In_809,In_576);
and U3333 (N_3333,In_952,In_103);
or U3334 (N_3334,In_391,In_1275);
nand U3335 (N_3335,In_1284,In_546);
or U3336 (N_3336,In_1448,In_1282);
or U3337 (N_3337,In_994,In_508);
nand U3338 (N_3338,In_1177,In_431);
nor U3339 (N_3339,In_1074,In_134);
or U3340 (N_3340,In_1131,In_490);
and U3341 (N_3341,In_621,In_1247);
nor U3342 (N_3342,In_257,In_576);
and U3343 (N_3343,In_745,In_486);
nor U3344 (N_3344,In_519,In_775);
nor U3345 (N_3345,In_1203,In_473);
nand U3346 (N_3346,In_96,In_599);
or U3347 (N_3347,In_79,In_333);
nand U3348 (N_3348,In_679,In_834);
xor U3349 (N_3349,In_956,In_119);
nand U3350 (N_3350,In_818,In_1209);
nand U3351 (N_3351,In_469,In_60);
nor U3352 (N_3352,In_1019,In_398);
nor U3353 (N_3353,In_764,In_505);
nor U3354 (N_3354,In_713,In_1135);
or U3355 (N_3355,In_892,In_379);
or U3356 (N_3356,In_385,In_474);
or U3357 (N_3357,In_162,In_808);
nor U3358 (N_3358,In_958,In_913);
and U3359 (N_3359,In_288,In_1398);
and U3360 (N_3360,In_233,In_1269);
nand U3361 (N_3361,In_18,In_583);
nor U3362 (N_3362,In_895,In_317);
nand U3363 (N_3363,In_1467,In_424);
nand U3364 (N_3364,In_1320,In_1458);
or U3365 (N_3365,In_590,In_205);
nor U3366 (N_3366,In_832,In_709);
or U3367 (N_3367,In_1167,In_1068);
nand U3368 (N_3368,In_1335,In_224);
nor U3369 (N_3369,In_326,In_557);
nand U3370 (N_3370,In_1146,In_426);
nor U3371 (N_3371,In_1006,In_985);
and U3372 (N_3372,In_697,In_706);
nor U3373 (N_3373,In_766,In_439);
and U3374 (N_3374,In_412,In_1342);
xnor U3375 (N_3375,In_1449,In_749);
or U3376 (N_3376,In_367,In_383);
and U3377 (N_3377,In_1236,In_1226);
and U3378 (N_3378,In_1102,In_1308);
nand U3379 (N_3379,In_475,In_1336);
nor U3380 (N_3380,In_82,In_1416);
nor U3381 (N_3381,In_287,In_824);
nand U3382 (N_3382,In_899,In_466);
nand U3383 (N_3383,In_29,In_92);
and U3384 (N_3384,In_383,In_660);
nor U3385 (N_3385,In_882,In_538);
nor U3386 (N_3386,In_734,In_1003);
or U3387 (N_3387,In_1278,In_1003);
or U3388 (N_3388,In_949,In_117);
nand U3389 (N_3389,In_403,In_873);
nand U3390 (N_3390,In_1053,In_856);
nand U3391 (N_3391,In_310,In_553);
or U3392 (N_3392,In_767,In_463);
nand U3393 (N_3393,In_1018,In_682);
or U3394 (N_3394,In_162,In_981);
or U3395 (N_3395,In_1482,In_1015);
nor U3396 (N_3396,In_363,In_375);
and U3397 (N_3397,In_484,In_611);
or U3398 (N_3398,In_627,In_1321);
nor U3399 (N_3399,In_1358,In_119);
or U3400 (N_3400,In_440,In_402);
nand U3401 (N_3401,In_870,In_303);
nor U3402 (N_3402,In_780,In_1199);
nor U3403 (N_3403,In_1469,In_1161);
xor U3404 (N_3404,In_289,In_1053);
nand U3405 (N_3405,In_1234,In_1236);
or U3406 (N_3406,In_442,In_923);
or U3407 (N_3407,In_1357,In_367);
or U3408 (N_3408,In_814,In_1134);
nor U3409 (N_3409,In_920,In_1070);
nand U3410 (N_3410,In_1434,In_1240);
nand U3411 (N_3411,In_25,In_267);
xor U3412 (N_3412,In_609,In_1409);
nand U3413 (N_3413,In_439,In_1282);
nor U3414 (N_3414,In_1195,In_147);
and U3415 (N_3415,In_540,In_660);
or U3416 (N_3416,In_831,In_103);
xor U3417 (N_3417,In_517,In_1178);
nor U3418 (N_3418,In_1373,In_443);
or U3419 (N_3419,In_789,In_1067);
nand U3420 (N_3420,In_1113,In_1476);
nand U3421 (N_3421,In_1128,In_929);
and U3422 (N_3422,In_322,In_1237);
nand U3423 (N_3423,In_1362,In_1487);
nand U3424 (N_3424,In_1079,In_1204);
nand U3425 (N_3425,In_626,In_1236);
or U3426 (N_3426,In_462,In_632);
and U3427 (N_3427,In_965,In_212);
nand U3428 (N_3428,In_76,In_834);
nor U3429 (N_3429,In_835,In_184);
and U3430 (N_3430,In_204,In_1107);
and U3431 (N_3431,In_1188,In_118);
and U3432 (N_3432,In_1445,In_14);
and U3433 (N_3433,In_1437,In_962);
nor U3434 (N_3434,In_644,In_1458);
nand U3435 (N_3435,In_787,In_1053);
or U3436 (N_3436,In_94,In_505);
or U3437 (N_3437,In_858,In_1388);
and U3438 (N_3438,In_604,In_968);
or U3439 (N_3439,In_1368,In_732);
nand U3440 (N_3440,In_171,In_1046);
or U3441 (N_3441,In_655,In_1489);
nor U3442 (N_3442,In_1128,In_1112);
and U3443 (N_3443,In_240,In_1081);
xor U3444 (N_3444,In_430,In_213);
and U3445 (N_3445,In_236,In_1077);
and U3446 (N_3446,In_966,In_566);
or U3447 (N_3447,In_581,In_457);
nor U3448 (N_3448,In_1132,In_690);
xor U3449 (N_3449,In_368,In_875);
nand U3450 (N_3450,In_382,In_667);
nor U3451 (N_3451,In_974,In_669);
xnor U3452 (N_3452,In_246,In_1150);
nor U3453 (N_3453,In_742,In_1135);
or U3454 (N_3454,In_44,In_719);
or U3455 (N_3455,In_523,In_74);
nand U3456 (N_3456,In_106,In_1467);
nand U3457 (N_3457,In_543,In_280);
nor U3458 (N_3458,In_321,In_681);
xnor U3459 (N_3459,In_45,In_433);
and U3460 (N_3460,In_206,In_586);
and U3461 (N_3461,In_332,In_898);
nor U3462 (N_3462,In_109,In_463);
or U3463 (N_3463,In_1484,In_518);
nand U3464 (N_3464,In_970,In_767);
nor U3465 (N_3465,In_208,In_140);
xnor U3466 (N_3466,In_768,In_16);
or U3467 (N_3467,In_198,In_1009);
and U3468 (N_3468,In_1174,In_567);
or U3469 (N_3469,In_168,In_48);
nor U3470 (N_3470,In_944,In_1398);
xnor U3471 (N_3471,In_610,In_204);
nor U3472 (N_3472,In_1226,In_324);
and U3473 (N_3473,In_217,In_324);
or U3474 (N_3474,In_1295,In_859);
or U3475 (N_3475,In_188,In_387);
and U3476 (N_3476,In_1000,In_618);
nor U3477 (N_3477,In_1110,In_982);
nand U3478 (N_3478,In_42,In_423);
and U3479 (N_3479,In_92,In_1191);
nor U3480 (N_3480,In_1126,In_1152);
and U3481 (N_3481,In_609,In_445);
and U3482 (N_3482,In_25,In_1022);
xnor U3483 (N_3483,In_1366,In_179);
and U3484 (N_3484,In_737,In_1158);
nor U3485 (N_3485,In_1462,In_460);
and U3486 (N_3486,In_116,In_1151);
nand U3487 (N_3487,In_1009,In_597);
nand U3488 (N_3488,In_162,In_624);
or U3489 (N_3489,In_230,In_1039);
nand U3490 (N_3490,In_1101,In_725);
nand U3491 (N_3491,In_1457,In_1345);
and U3492 (N_3492,In_664,In_469);
and U3493 (N_3493,In_481,In_288);
and U3494 (N_3494,In_1438,In_746);
xor U3495 (N_3495,In_117,In_79);
nand U3496 (N_3496,In_1399,In_867);
nor U3497 (N_3497,In_1381,In_989);
nor U3498 (N_3498,In_970,In_246);
nor U3499 (N_3499,In_434,In_144);
xnor U3500 (N_3500,In_823,In_82);
nor U3501 (N_3501,In_777,In_548);
or U3502 (N_3502,In_1382,In_957);
and U3503 (N_3503,In_399,In_208);
nand U3504 (N_3504,In_1014,In_1069);
and U3505 (N_3505,In_1421,In_976);
nand U3506 (N_3506,In_402,In_1242);
and U3507 (N_3507,In_228,In_825);
or U3508 (N_3508,In_73,In_784);
nand U3509 (N_3509,In_283,In_417);
xnor U3510 (N_3510,In_277,In_12);
and U3511 (N_3511,In_493,In_597);
or U3512 (N_3512,In_289,In_885);
nand U3513 (N_3513,In_3,In_674);
nand U3514 (N_3514,In_1074,In_722);
and U3515 (N_3515,In_1139,In_1060);
or U3516 (N_3516,In_719,In_306);
and U3517 (N_3517,In_495,In_843);
nand U3518 (N_3518,In_167,In_323);
nand U3519 (N_3519,In_740,In_795);
nor U3520 (N_3520,In_334,In_1030);
nand U3521 (N_3521,In_233,In_12);
and U3522 (N_3522,In_223,In_252);
and U3523 (N_3523,In_1372,In_814);
and U3524 (N_3524,In_235,In_802);
or U3525 (N_3525,In_1426,In_207);
and U3526 (N_3526,In_1322,In_314);
nand U3527 (N_3527,In_1189,In_1197);
or U3528 (N_3528,In_1073,In_94);
and U3529 (N_3529,In_119,In_1274);
xnor U3530 (N_3530,In_825,In_398);
xor U3531 (N_3531,In_1298,In_414);
nor U3532 (N_3532,In_378,In_634);
or U3533 (N_3533,In_841,In_942);
and U3534 (N_3534,In_1056,In_183);
nand U3535 (N_3535,In_348,In_510);
xor U3536 (N_3536,In_1184,In_693);
nand U3537 (N_3537,In_485,In_1470);
and U3538 (N_3538,In_174,In_311);
and U3539 (N_3539,In_1178,In_1231);
nand U3540 (N_3540,In_1478,In_395);
or U3541 (N_3541,In_1095,In_1406);
xor U3542 (N_3542,In_686,In_1428);
nor U3543 (N_3543,In_859,In_23);
or U3544 (N_3544,In_1404,In_900);
and U3545 (N_3545,In_1271,In_1157);
nand U3546 (N_3546,In_581,In_756);
or U3547 (N_3547,In_551,In_1359);
nor U3548 (N_3548,In_820,In_531);
and U3549 (N_3549,In_1417,In_893);
nand U3550 (N_3550,In_587,In_786);
nand U3551 (N_3551,In_1399,In_1417);
and U3552 (N_3552,In_1164,In_1355);
or U3553 (N_3553,In_1261,In_1318);
xnor U3554 (N_3554,In_883,In_501);
and U3555 (N_3555,In_211,In_31);
and U3556 (N_3556,In_782,In_491);
nor U3557 (N_3557,In_481,In_796);
or U3558 (N_3558,In_1263,In_1454);
and U3559 (N_3559,In_101,In_1437);
nand U3560 (N_3560,In_760,In_341);
and U3561 (N_3561,In_186,In_122);
nand U3562 (N_3562,In_1226,In_305);
nor U3563 (N_3563,In_262,In_922);
xnor U3564 (N_3564,In_1118,In_996);
xor U3565 (N_3565,In_725,In_188);
nand U3566 (N_3566,In_1144,In_69);
nand U3567 (N_3567,In_142,In_995);
or U3568 (N_3568,In_824,In_210);
and U3569 (N_3569,In_925,In_760);
or U3570 (N_3570,In_1129,In_269);
nand U3571 (N_3571,In_440,In_141);
nand U3572 (N_3572,In_225,In_535);
nor U3573 (N_3573,In_660,In_212);
or U3574 (N_3574,In_1263,In_1365);
and U3575 (N_3575,In_1287,In_754);
nand U3576 (N_3576,In_1093,In_832);
or U3577 (N_3577,In_605,In_1127);
or U3578 (N_3578,In_587,In_543);
and U3579 (N_3579,In_987,In_468);
nor U3580 (N_3580,In_321,In_81);
and U3581 (N_3581,In_1361,In_137);
nor U3582 (N_3582,In_952,In_1293);
or U3583 (N_3583,In_705,In_400);
and U3584 (N_3584,In_980,In_1330);
nor U3585 (N_3585,In_515,In_1055);
and U3586 (N_3586,In_672,In_321);
or U3587 (N_3587,In_922,In_1467);
or U3588 (N_3588,In_1450,In_319);
nor U3589 (N_3589,In_616,In_27);
and U3590 (N_3590,In_859,In_1383);
and U3591 (N_3591,In_1030,In_930);
or U3592 (N_3592,In_179,In_857);
and U3593 (N_3593,In_166,In_269);
or U3594 (N_3594,In_1331,In_112);
xor U3595 (N_3595,In_1456,In_481);
and U3596 (N_3596,In_1398,In_1308);
or U3597 (N_3597,In_433,In_1098);
xnor U3598 (N_3598,In_1189,In_1394);
nor U3599 (N_3599,In_1293,In_1092);
or U3600 (N_3600,In_1444,In_403);
and U3601 (N_3601,In_249,In_1314);
nor U3602 (N_3602,In_1063,In_83);
or U3603 (N_3603,In_767,In_1118);
and U3604 (N_3604,In_210,In_134);
nand U3605 (N_3605,In_947,In_697);
nand U3606 (N_3606,In_142,In_182);
nor U3607 (N_3607,In_711,In_267);
or U3608 (N_3608,In_1426,In_1478);
and U3609 (N_3609,In_491,In_1160);
or U3610 (N_3610,In_968,In_879);
or U3611 (N_3611,In_1185,In_119);
or U3612 (N_3612,In_779,In_1231);
nor U3613 (N_3613,In_721,In_1172);
nand U3614 (N_3614,In_240,In_1370);
and U3615 (N_3615,In_1185,In_1227);
nand U3616 (N_3616,In_1182,In_495);
and U3617 (N_3617,In_925,In_835);
nand U3618 (N_3618,In_1469,In_1368);
nor U3619 (N_3619,In_1300,In_1269);
or U3620 (N_3620,In_504,In_807);
and U3621 (N_3621,In_586,In_673);
or U3622 (N_3622,In_1140,In_333);
nor U3623 (N_3623,In_1452,In_460);
or U3624 (N_3624,In_1234,In_1266);
nor U3625 (N_3625,In_564,In_940);
and U3626 (N_3626,In_410,In_661);
and U3627 (N_3627,In_912,In_708);
xnor U3628 (N_3628,In_157,In_1467);
and U3629 (N_3629,In_1390,In_771);
nor U3630 (N_3630,In_1154,In_981);
or U3631 (N_3631,In_997,In_184);
xor U3632 (N_3632,In_794,In_131);
nor U3633 (N_3633,In_237,In_734);
or U3634 (N_3634,In_878,In_542);
and U3635 (N_3635,In_658,In_302);
or U3636 (N_3636,In_140,In_628);
and U3637 (N_3637,In_553,In_845);
and U3638 (N_3638,In_58,In_1111);
nand U3639 (N_3639,In_119,In_367);
or U3640 (N_3640,In_186,In_212);
or U3641 (N_3641,In_1072,In_315);
nor U3642 (N_3642,In_690,In_199);
xor U3643 (N_3643,In_925,In_392);
nand U3644 (N_3644,In_33,In_853);
nand U3645 (N_3645,In_107,In_436);
or U3646 (N_3646,In_985,In_955);
nand U3647 (N_3647,In_1493,In_141);
nor U3648 (N_3648,In_973,In_1011);
or U3649 (N_3649,In_1047,In_1136);
and U3650 (N_3650,In_393,In_467);
nor U3651 (N_3651,In_284,In_281);
nand U3652 (N_3652,In_181,In_561);
nand U3653 (N_3653,In_453,In_1044);
and U3654 (N_3654,In_705,In_1276);
or U3655 (N_3655,In_257,In_1168);
nor U3656 (N_3656,In_844,In_319);
or U3657 (N_3657,In_211,In_565);
nor U3658 (N_3658,In_142,In_1486);
nand U3659 (N_3659,In_1485,In_103);
nand U3660 (N_3660,In_1342,In_1206);
or U3661 (N_3661,In_845,In_675);
or U3662 (N_3662,In_137,In_128);
or U3663 (N_3663,In_838,In_1152);
or U3664 (N_3664,In_105,In_1110);
and U3665 (N_3665,In_828,In_1301);
or U3666 (N_3666,In_830,In_1136);
nand U3667 (N_3667,In_614,In_844);
or U3668 (N_3668,In_250,In_147);
or U3669 (N_3669,In_295,In_245);
and U3670 (N_3670,In_1257,In_486);
nand U3671 (N_3671,In_1012,In_1338);
nor U3672 (N_3672,In_848,In_1017);
nand U3673 (N_3673,In_529,In_1454);
nor U3674 (N_3674,In_313,In_256);
and U3675 (N_3675,In_750,In_204);
or U3676 (N_3676,In_736,In_1127);
and U3677 (N_3677,In_103,In_1083);
nand U3678 (N_3678,In_876,In_383);
nor U3679 (N_3679,In_32,In_1486);
nor U3680 (N_3680,In_1045,In_70);
nand U3681 (N_3681,In_1302,In_1191);
and U3682 (N_3682,In_1275,In_33);
or U3683 (N_3683,In_1261,In_91);
nor U3684 (N_3684,In_481,In_880);
nor U3685 (N_3685,In_396,In_465);
nor U3686 (N_3686,In_140,In_480);
nand U3687 (N_3687,In_1463,In_596);
and U3688 (N_3688,In_1283,In_1210);
nor U3689 (N_3689,In_1379,In_887);
or U3690 (N_3690,In_75,In_100);
nand U3691 (N_3691,In_1326,In_875);
xor U3692 (N_3692,In_1229,In_1067);
or U3693 (N_3693,In_307,In_1038);
nand U3694 (N_3694,In_955,In_1279);
nor U3695 (N_3695,In_929,In_700);
and U3696 (N_3696,In_462,In_1314);
nor U3697 (N_3697,In_1359,In_662);
and U3698 (N_3698,In_1360,In_10);
nor U3699 (N_3699,In_541,In_1461);
and U3700 (N_3700,In_1449,In_552);
nor U3701 (N_3701,In_573,In_475);
xnor U3702 (N_3702,In_1357,In_810);
nand U3703 (N_3703,In_1104,In_922);
nand U3704 (N_3704,In_522,In_116);
and U3705 (N_3705,In_492,In_603);
nor U3706 (N_3706,In_926,In_857);
or U3707 (N_3707,In_406,In_1371);
nand U3708 (N_3708,In_34,In_989);
and U3709 (N_3709,In_759,In_1386);
nor U3710 (N_3710,In_277,In_1045);
and U3711 (N_3711,In_26,In_163);
xnor U3712 (N_3712,In_1249,In_1256);
xnor U3713 (N_3713,In_1331,In_116);
nand U3714 (N_3714,In_1366,In_854);
nor U3715 (N_3715,In_1435,In_267);
nor U3716 (N_3716,In_1094,In_507);
nand U3717 (N_3717,In_45,In_1365);
xnor U3718 (N_3718,In_535,In_220);
nand U3719 (N_3719,In_1417,In_1241);
and U3720 (N_3720,In_1260,In_1127);
or U3721 (N_3721,In_937,In_84);
xnor U3722 (N_3722,In_37,In_681);
and U3723 (N_3723,In_824,In_472);
and U3724 (N_3724,In_800,In_491);
nor U3725 (N_3725,In_153,In_371);
or U3726 (N_3726,In_1133,In_1467);
or U3727 (N_3727,In_895,In_1138);
nor U3728 (N_3728,In_569,In_52);
xor U3729 (N_3729,In_594,In_917);
or U3730 (N_3730,In_44,In_726);
or U3731 (N_3731,In_606,In_494);
or U3732 (N_3732,In_355,In_850);
and U3733 (N_3733,In_1162,In_612);
nor U3734 (N_3734,In_1020,In_1418);
and U3735 (N_3735,In_1372,In_1131);
and U3736 (N_3736,In_1218,In_885);
or U3737 (N_3737,In_446,In_942);
nand U3738 (N_3738,In_543,In_943);
nand U3739 (N_3739,In_555,In_35);
nand U3740 (N_3740,In_502,In_147);
or U3741 (N_3741,In_302,In_383);
or U3742 (N_3742,In_118,In_990);
or U3743 (N_3743,In_475,In_1097);
nand U3744 (N_3744,In_1185,In_735);
nand U3745 (N_3745,In_562,In_1017);
nand U3746 (N_3746,In_1420,In_537);
nand U3747 (N_3747,In_225,In_1296);
nand U3748 (N_3748,In_847,In_390);
or U3749 (N_3749,In_1349,In_695);
nor U3750 (N_3750,In_281,In_1368);
xnor U3751 (N_3751,In_946,In_424);
nand U3752 (N_3752,In_48,In_815);
nor U3753 (N_3753,In_150,In_1084);
xnor U3754 (N_3754,In_1201,In_973);
and U3755 (N_3755,In_200,In_836);
nand U3756 (N_3756,In_1014,In_379);
or U3757 (N_3757,In_1262,In_461);
and U3758 (N_3758,In_1313,In_343);
nand U3759 (N_3759,In_394,In_946);
or U3760 (N_3760,In_457,In_59);
and U3761 (N_3761,In_909,In_383);
or U3762 (N_3762,In_323,In_379);
or U3763 (N_3763,In_357,In_948);
or U3764 (N_3764,In_294,In_197);
and U3765 (N_3765,In_1445,In_162);
and U3766 (N_3766,In_464,In_501);
nor U3767 (N_3767,In_173,In_1096);
or U3768 (N_3768,In_31,In_691);
xor U3769 (N_3769,In_1203,In_894);
or U3770 (N_3770,In_1144,In_1455);
nor U3771 (N_3771,In_77,In_318);
or U3772 (N_3772,In_1013,In_427);
and U3773 (N_3773,In_1221,In_327);
or U3774 (N_3774,In_440,In_797);
or U3775 (N_3775,In_790,In_961);
nand U3776 (N_3776,In_1352,In_399);
or U3777 (N_3777,In_939,In_1430);
or U3778 (N_3778,In_1402,In_1029);
or U3779 (N_3779,In_91,In_1175);
or U3780 (N_3780,In_424,In_700);
or U3781 (N_3781,In_752,In_1129);
nor U3782 (N_3782,In_871,In_1118);
nand U3783 (N_3783,In_176,In_1201);
nand U3784 (N_3784,In_206,In_1148);
and U3785 (N_3785,In_377,In_186);
nand U3786 (N_3786,In_320,In_8);
nor U3787 (N_3787,In_1009,In_1303);
and U3788 (N_3788,In_907,In_936);
or U3789 (N_3789,In_222,In_1370);
nor U3790 (N_3790,In_433,In_58);
nor U3791 (N_3791,In_979,In_1460);
nand U3792 (N_3792,In_1153,In_334);
nor U3793 (N_3793,In_877,In_1125);
and U3794 (N_3794,In_1044,In_796);
nand U3795 (N_3795,In_1263,In_898);
and U3796 (N_3796,In_1162,In_1102);
or U3797 (N_3797,In_65,In_675);
nand U3798 (N_3798,In_462,In_983);
or U3799 (N_3799,In_355,In_323);
nand U3800 (N_3800,In_1344,In_955);
nor U3801 (N_3801,In_572,In_289);
xnor U3802 (N_3802,In_605,In_1252);
and U3803 (N_3803,In_316,In_1070);
or U3804 (N_3804,In_529,In_30);
xor U3805 (N_3805,In_565,In_408);
nand U3806 (N_3806,In_420,In_576);
xor U3807 (N_3807,In_875,In_437);
or U3808 (N_3808,In_420,In_550);
and U3809 (N_3809,In_961,In_25);
and U3810 (N_3810,In_401,In_1115);
nand U3811 (N_3811,In_410,In_791);
and U3812 (N_3812,In_363,In_800);
nand U3813 (N_3813,In_538,In_1295);
and U3814 (N_3814,In_705,In_1484);
and U3815 (N_3815,In_631,In_191);
nand U3816 (N_3816,In_1134,In_606);
and U3817 (N_3817,In_1379,In_34);
nor U3818 (N_3818,In_410,In_628);
and U3819 (N_3819,In_1168,In_786);
and U3820 (N_3820,In_1471,In_522);
or U3821 (N_3821,In_1073,In_1436);
nand U3822 (N_3822,In_300,In_1236);
xnor U3823 (N_3823,In_232,In_1082);
nand U3824 (N_3824,In_1074,In_1071);
xnor U3825 (N_3825,In_1192,In_1402);
or U3826 (N_3826,In_107,In_895);
and U3827 (N_3827,In_14,In_1187);
and U3828 (N_3828,In_1347,In_975);
or U3829 (N_3829,In_51,In_721);
and U3830 (N_3830,In_326,In_390);
and U3831 (N_3831,In_1260,In_863);
and U3832 (N_3832,In_676,In_1482);
and U3833 (N_3833,In_967,In_748);
nand U3834 (N_3834,In_1270,In_1114);
or U3835 (N_3835,In_394,In_996);
nand U3836 (N_3836,In_102,In_914);
xnor U3837 (N_3837,In_933,In_463);
and U3838 (N_3838,In_1199,In_755);
or U3839 (N_3839,In_1140,In_177);
nor U3840 (N_3840,In_702,In_1167);
nand U3841 (N_3841,In_94,In_99);
nor U3842 (N_3842,In_183,In_787);
nand U3843 (N_3843,In_159,In_596);
xor U3844 (N_3844,In_1242,In_1186);
nor U3845 (N_3845,In_1315,In_1327);
nand U3846 (N_3846,In_324,In_263);
or U3847 (N_3847,In_644,In_1226);
xor U3848 (N_3848,In_71,In_1099);
nand U3849 (N_3849,In_1039,In_200);
or U3850 (N_3850,In_1265,In_250);
and U3851 (N_3851,In_78,In_1013);
or U3852 (N_3852,In_443,In_997);
xor U3853 (N_3853,In_698,In_1315);
and U3854 (N_3854,In_929,In_162);
or U3855 (N_3855,In_288,In_758);
nor U3856 (N_3856,In_842,In_551);
and U3857 (N_3857,In_400,In_1227);
and U3858 (N_3858,In_1493,In_1309);
nand U3859 (N_3859,In_471,In_1123);
and U3860 (N_3860,In_763,In_679);
nor U3861 (N_3861,In_279,In_1499);
nand U3862 (N_3862,In_750,In_250);
or U3863 (N_3863,In_914,In_1056);
nor U3864 (N_3864,In_1015,In_812);
or U3865 (N_3865,In_855,In_446);
and U3866 (N_3866,In_1492,In_7);
nor U3867 (N_3867,In_234,In_1083);
or U3868 (N_3868,In_1167,In_1310);
xor U3869 (N_3869,In_157,In_47);
nand U3870 (N_3870,In_1018,In_9);
nor U3871 (N_3871,In_1429,In_1158);
or U3872 (N_3872,In_725,In_660);
or U3873 (N_3873,In_24,In_979);
nor U3874 (N_3874,In_1344,In_887);
xnor U3875 (N_3875,In_383,In_1044);
xnor U3876 (N_3876,In_1209,In_540);
or U3877 (N_3877,In_254,In_890);
or U3878 (N_3878,In_629,In_689);
nor U3879 (N_3879,In_1409,In_356);
nand U3880 (N_3880,In_268,In_929);
and U3881 (N_3881,In_1432,In_545);
xnor U3882 (N_3882,In_284,In_1247);
and U3883 (N_3883,In_504,In_660);
nand U3884 (N_3884,In_998,In_545);
and U3885 (N_3885,In_1312,In_388);
and U3886 (N_3886,In_571,In_266);
and U3887 (N_3887,In_427,In_619);
or U3888 (N_3888,In_353,In_1008);
or U3889 (N_3889,In_1394,In_1249);
or U3890 (N_3890,In_1455,In_1414);
nor U3891 (N_3891,In_1368,In_376);
or U3892 (N_3892,In_1032,In_711);
or U3893 (N_3893,In_4,In_3);
nand U3894 (N_3894,In_1068,In_1262);
nor U3895 (N_3895,In_1139,In_1131);
nand U3896 (N_3896,In_833,In_872);
nand U3897 (N_3897,In_1449,In_696);
nor U3898 (N_3898,In_290,In_1378);
or U3899 (N_3899,In_88,In_1193);
or U3900 (N_3900,In_1417,In_922);
or U3901 (N_3901,In_816,In_1270);
nor U3902 (N_3902,In_269,In_263);
nor U3903 (N_3903,In_21,In_1276);
xnor U3904 (N_3904,In_77,In_1406);
nor U3905 (N_3905,In_1202,In_89);
xor U3906 (N_3906,In_52,In_1416);
nand U3907 (N_3907,In_652,In_73);
or U3908 (N_3908,In_917,In_391);
nand U3909 (N_3909,In_861,In_1221);
or U3910 (N_3910,In_422,In_1092);
or U3911 (N_3911,In_1207,In_594);
nor U3912 (N_3912,In_1328,In_335);
and U3913 (N_3913,In_640,In_1152);
nor U3914 (N_3914,In_721,In_272);
nand U3915 (N_3915,In_356,In_695);
or U3916 (N_3916,In_347,In_437);
and U3917 (N_3917,In_1485,In_1341);
and U3918 (N_3918,In_1294,In_1168);
or U3919 (N_3919,In_68,In_391);
nor U3920 (N_3920,In_797,In_204);
nor U3921 (N_3921,In_253,In_202);
or U3922 (N_3922,In_571,In_1122);
nor U3923 (N_3923,In_560,In_1352);
nor U3924 (N_3924,In_955,In_1175);
nand U3925 (N_3925,In_238,In_779);
and U3926 (N_3926,In_202,In_485);
and U3927 (N_3927,In_64,In_987);
or U3928 (N_3928,In_521,In_117);
and U3929 (N_3929,In_828,In_1464);
or U3930 (N_3930,In_906,In_665);
or U3931 (N_3931,In_1387,In_997);
or U3932 (N_3932,In_1087,In_476);
xor U3933 (N_3933,In_460,In_746);
nand U3934 (N_3934,In_132,In_69);
and U3935 (N_3935,In_885,In_765);
nand U3936 (N_3936,In_246,In_472);
or U3937 (N_3937,In_575,In_1271);
nand U3938 (N_3938,In_610,In_387);
and U3939 (N_3939,In_734,In_818);
and U3940 (N_3940,In_209,In_1078);
nor U3941 (N_3941,In_142,In_1324);
nand U3942 (N_3942,In_80,In_1408);
nor U3943 (N_3943,In_1390,In_452);
and U3944 (N_3944,In_1132,In_1018);
nand U3945 (N_3945,In_1093,In_1386);
xnor U3946 (N_3946,In_779,In_225);
xor U3947 (N_3947,In_968,In_975);
nor U3948 (N_3948,In_1424,In_1004);
and U3949 (N_3949,In_1006,In_524);
and U3950 (N_3950,In_33,In_543);
and U3951 (N_3951,In_1332,In_1129);
nand U3952 (N_3952,In_349,In_432);
nand U3953 (N_3953,In_1,In_946);
or U3954 (N_3954,In_660,In_86);
or U3955 (N_3955,In_1398,In_1396);
or U3956 (N_3956,In_879,In_633);
or U3957 (N_3957,In_818,In_1430);
xor U3958 (N_3958,In_1173,In_886);
nand U3959 (N_3959,In_1208,In_741);
xnor U3960 (N_3960,In_1276,In_327);
nand U3961 (N_3961,In_183,In_949);
and U3962 (N_3962,In_532,In_176);
or U3963 (N_3963,In_864,In_1223);
or U3964 (N_3964,In_824,In_845);
xnor U3965 (N_3965,In_908,In_625);
or U3966 (N_3966,In_606,In_1306);
and U3967 (N_3967,In_1471,In_955);
and U3968 (N_3968,In_706,In_472);
nor U3969 (N_3969,In_951,In_238);
or U3970 (N_3970,In_1343,In_839);
and U3971 (N_3971,In_1079,In_710);
or U3972 (N_3972,In_153,In_987);
and U3973 (N_3973,In_167,In_18);
nand U3974 (N_3974,In_358,In_719);
nor U3975 (N_3975,In_1044,In_328);
and U3976 (N_3976,In_1305,In_655);
nand U3977 (N_3977,In_53,In_1021);
or U3978 (N_3978,In_618,In_644);
nand U3979 (N_3979,In_612,In_755);
nor U3980 (N_3980,In_1331,In_903);
nand U3981 (N_3981,In_1448,In_813);
nor U3982 (N_3982,In_650,In_427);
nand U3983 (N_3983,In_792,In_1325);
or U3984 (N_3984,In_52,In_537);
nand U3985 (N_3985,In_1280,In_31);
nor U3986 (N_3986,In_1101,In_649);
and U3987 (N_3987,In_197,In_1287);
and U3988 (N_3988,In_604,In_361);
nor U3989 (N_3989,In_1264,In_172);
or U3990 (N_3990,In_1402,In_97);
and U3991 (N_3991,In_667,In_1423);
and U3992 (N_3992,In_363,In_926);
or U3993 (N_3993,In_1212,In_129);
or U3994 (N_3994,In_296,In_223);
xor U3995 (N_3995,In_987,In_1365);
and U3996 (N_3996,In_916,In_908);
and U3997 (N_3997,In_934,In_434);
and U3998 (N_3998,In_342,In_655);
nor U3999 (N_3999,In_244,In_1293);
or U4000 (N_4000,In_695,In_625);
or U4001 (N_4001,In_390,In_267);
or U4002 (N_4002,In_306,In_23);
and U4003 (N_4003,In_713,In_1497);
and U4004 (N_4004,In_945,In_1311);
nor U4005 (N_4005,In_663,In_374);
nand U4006 (N_4006,In_544,In_1124);
nor U4007 (N_4007,In_5,In_669);
nand U4008 (N_4008,In_243,In_290);
and U4009 (N_4009,In_596,In_131);
xor U4010 (N_4010,In_773,In_489);
and U4011 (N_4011,In_1485,In_1144);
xnor U4012 (N_4012,In_300,In_1184);
or U4013 (N_4013,In_322,In_92);
nor U4014 (N_4014,In_424,In_348);
nand U4015 (N_4015,In_1076,In_222);
nand U4016 (N_4016,In_835,In_1212);
nor U4017 (N_4017,In_1347,In_511);
and U4018 (N_4018,In_1452,In_791);
or U4019 (N_4019,In_221,In_517);
nor U4020 (N_4020,In_842,In_1029);
or U4021 (N_4021,In_550,In_556);
nand U4022 (N_4022,In_809,In_1160);
and U4023 (N_4023,In_1311,In_197);
and U4024 (N_4024,In_300,In_981);
or U4025 (N_4025,In_1280,In_624);
nand U4026 (N_4026,In_383,In_23);
or U4027 (N_4027,In_415,In_486);
nand U4028 (N_4028,In_1120,In_768);
or U4029 (N_4029,In_792,In_1078);
and U4030 (N_4030,In_1247,In_1042);
or U4031 (N_4031,In_458,In_31);
xnor U4032 (N_4032,In_282,In_267);
or U4033 (N_4033,In_959,In_24);
and U4034 (N_4034,In_1077,In_107);
or U4035 (N_4035,In_203,In_1324);
xnor U4036 (N_4036,In_1319,In_207);
and U4037 (N_4037,In_909,In_727);
nor U4038 (N_4038,In_1191,In_196);
xor U4039 (N_4039,In_166,In_1118);
or U4040 (N_4040,In_709,In_223);
or U4041 (N_4041,In_318,In_1196);
xnor U4042 (N_4042,In_109,In_1351);
or U4043 (N_4043,In_731,In_330);
nor U4044 (N_4044,In_487,In_523);
nor U4045 (N_4045,In_1063,In_339);
and U4046 (N_4046,In_723,In_1125);
and U4047 (N_4047,In_935,In_1159);
nor U4048 (N_4048,In_1199,In_919);
nand U4049 (N_4049,In_1120,In_290);
nor U4050 (N_4050,In_332,In_305);
nand U4051 (N_4051,In_1362,In_1209);
and U4052 (N_4052,In_790,In_782);
nor U4053 (N_4053,In_37,In_1403);
or U4054 (N_4054,In_212,In_925);
nand U4055 (N_4055,In_501,In_1115);
and U4056 (N_4056,In_1048,In_1007);
and U4057 (N_4057,In_1282,In_512);
nand U4058 (N_4058,In_414,In_1124);
or U4059 (N_4059,In_1022,In_431);
nor U4060 (N_4060,In_59,In_90);
nor U4061 (N_4061,In_1335,In_1226);
and U4062 (N_4062,In_206,In_1011);
nor U4063 (N_4063,In_823,In_1033);
nor U4064 (N_4064,In_781,In_176);
xnor U4065 (N_4065,In_1102,In_245);
and U4066 (N_4066,In_203,In_1038);
xor U4067 (N_4067,In_765,In_171);
or U4068 (N_4068,In_1228,In_633);
nor U4069 (N_4069,In_683,In_1488);
nand U4070 (N_4070,In_431,In_1162);
nand U4071 (N_4071,In_1432,In_1140);
and U4072 (N_4072,In_1372,In_1296);
nor U4073 (N_4073,In_271,In_1296);
nor U4074 (N_4074,In_520,In_1366);
and U4075 (N_4075,In_1498,In_1226);
and U4076 (N_4076,In_1086,In_1240);
or U4077 (N_4077,In_106,In_321);
or U4078 (N_4078,In_711,In_397);
nand U4079 (N_4079,In_117,In_793);
nand U4080 (N_4080,In_11,In_873);
and U4081 (N_4081,In_1487,In_846);
nor U4082 (N_4082,In_1228,In_710);
nand U4083 (N_4083,In_445,In_1320);
nor U4084 (N_4084,In_1028,In_467);
nor U4085 (N_4085,In_392,In_504);
nor U4086 (N_4086,In_1153,In_784);
or U4087 (N_4087,In_321,In_348);
or U4088 (N_4088,In_1430,In_914);
and U4089 (N_4089,In_1229,In_492);
nor U4090 (N_4090,In_1031,In_694);
xor U4091 (N_4091,In_1493,In_375);
xor U4092 (N_4092,In_359,In_1476);
or U4093 (N_4093,In_874,In_613);
xnor U4094 (N_4094,In_1307,In_766);
nor U4095 (N_4095,In_857,In_748);
or U4096 (N_4096,In_231,In_1355);
or U4097 (N_4097,In_1332,In_1100);
nor U4098 (N_4098,In_302,In_662);
xor U4099 (N_4099,In_297,In_244);
nand U4100 (N_4100,In_536,In_837);
or U4101 (N_4101,In_19,In_1195);
nand U4102 (N_4102,In_1423,In_85);
nand U4103 (N_4103,In_1464,In_1133);
nor U4104 (N_4104,In_754,In_227);
and U4105 (N_4105,In_60,In_1255);
xor U4106 (N_4106,In_1482,In_724);
or U4107 (N_4107,In_887,In_1000);
and U4108 (N_4108,In_671,In_246);
nand U4109 (N_4109,In_481,In_1138);
nor U4110 (N_4110,In_884,In_1481);
and U4111 (N_4111,In_1420,In_257);
nor U4112 (N_4112,In_671,In_1085);
nand U4113 (N_4113,In_25,In_314);
nor U4114 (N_4114,In_1414,In_815);
or U4115 (N_4115,In_1216,In_1221);
or U4116 (N_4116,In_1119,In_949);
xor U4117 (N_4117,In_351,In_896);
nor U4118 (N_4118,In_443,In_128);
nor U4119 (N_4119,In_797,In_912);
nor U4120 (N_4120,In_1076,In_71);
xor U4121 (N_4121,In_1455,In_1005);
nor U4122 (N_4122,In_971,In_904);
nand U4123 (N_4123,In_673,In_677);
nand U4124 (N_4124,In_819,In_987);
xor U4125 (N_4125,In_678,In_1054);
nand U4126 (N_4126,In_663,In_354);
nor U4127 (N_4127,In_374,In_1050);
nand U4128 (N_4128,In_299,In_750);
nor U4129 (N_4129,In_1313,In_1251);
nor U4130 (N_4130,In_641,In_237);
or U4131 (N_4131,In_243,In_718);
or U4132 (N_4132,In_486,In_303);
nor U4133 (N_4133,In_821,In_522);
and U4134 (N_4134,In_1490,In_66);
nand U4135 (N_4135,In_1168,In_252);
and U4136 (N_4136,In_1095,In_595);
and U4137 (N_4137,In_23,In_507);
and U4138 (N_4138,In_499,In_1098);
and U4139 (N_4139,In_355,In_881);
or U4140 (N_4140,In_1401,In_105);
nand U4141 (N_4141,In_758,In_1499);
xnor U4142 (N_4142,In_1488,In_386);
and U4143 (N_4143,In_887,In_1340);
nand U4144 (N_4144,In_1412,In_956);
xor U4145 (N_4145,In_173,In_826);
or U4146 (N_4146,In_1385,In_1090);
nand U4147 (N_4147,In_266,In_1439);
nor U4148 (N_4148,In_616,In_1139);
nor U4149 (N_4149,In_1088,In_984);
xnor U4150 (N_4150,In_1337,In_481);
or U4151 (N_4151,In_674,In_1350);
and U4152 (N_4152,In_502,In_581);
nand U4153 (N_4153,In_392,In_644);
or U4154 (N_4154,In_127,In_946);
nor U4155 (N_4155,In_183,In_677);
or U4156 (N_4156,In_142,In_593);
nor U4157 (N_4157,In_572,In_652);
nand U4158 (N_4158,In_637,In_12);
nor U4159 (N_4159,In_933,In_596);
and U4160 (N_4160,In_953,In_451);
and U4161 (N_4161,In_1277,In_811);
nand U4162 (N_4162,In_532,In_619);
nand U4163 (N_4163,In_438,In_1350);
and U4164 (N_4164,In_1338,In_1345);
nor U4165 (N_4165,In_891,In_245);
nor U4166 (N_4166,In_14,In_543);
and U4167 (N_4167,In_790,In_1103);
and U4168 (N_4168,In_942,In_569);
and U4169 (N_4169,In_313,In_1444);
nand U4170 (N_4170,In_962,In_1268);
or U4171 (N_4171,In_1430,In_1249);
nor U4172 (N_4172,In_381,In_84);
and U4173 (N_4173,In_1271,In_992);
xor U4174 (N_4174,In_290,In_1060);
nand U4175 (N_4175,In_1198,In_386);
nand U4176 (N_4176,In_1008,In_578);
nand U4177 (N_4177,In_561,In_671);
nand U4178 (N_4178,In_1243,In_1405);
nor U4179 (N_4179,In_336,In_578);
nor U4180 (N_4180,In_674,In_1264);
xnor U4181 (N_4181,In_1238,In_811);
or U4182 (N_4182,In_454,In_247);
and U4183 (N_4183,In_361,In_962);
or U4184 (N_4184,In_908,In_744);
xor U4185 (N_4185,In_786,In_751);
xor U4186 (N_4186,In_296,In_980);
nand U4187 (N_4187,In_403,In_1419);
or U4188 (N_4188,In_1426,In_1198);
or U4189 (N_4189,In_1073,In_745);
xor U4190 (N_4190,In_1014,In_311);
nor U4191 (N_4191,In_539,In_233);
nor U4192 (N_4192,In_14,In_481);
and U4193 (N_4193,In_1066,In_232);
nand U4194 (N_4194,In_1346,In_1293);
nor U4195 (N_4195,In_1252,In_1414);
nor U4196 (N_4196,In_1351,In_1255);
xor U4197 (N_4197,In_1321,In_336);
nor U4198 (N_4198,In_280,In_1317);
and U4199 (N_4199,In_186,In_1495);
xnor U4200 (N_4200,In_1260,In_251);
and U4201 (N_4201,In_1291,In_445);
or U4202 (N_4202,In_685,In_208);
nor U4203 (N_4203,In_1276,In_689);
or U4204 (N_4204,In_1482,In_635);
nand U4205 (N_4205,In_851,In_916);
xor U4206 (N_4206,In_833,In_982);
nor U4207 (N_4207,In_425,In_871);
xnor U4208 (N_4208,In_1221,In_352);
nand U4209 (N_4209,In_381,In_1169);
nand U4210 (N_4210,In_988,In_961);
nor U4211 (N_4211,In_201,In_73);
xnor U4212 (N_4212,In_1189,In_27);
and U4213 (N_4213,In_1056,In_574);
and U4214 (N_4214,In_737,In_1411);
nor U4215 (N_4215,In_921,In_1341);
nand U4216 (N_4216,In_424,In_269);
or U4217 (N_4217,In_1430,In_104);
and U4218 (N_4218,In_67,In_1157);
and U4219 (N_4219,In_1424,In_1023);
nor U4220 (N_4220,In_1416,In_714);
nor U4221 (N_4221,In_427,In_1023);
or U4222 (N_4222,In_599,In_352);
and U4223 (N_4223,In_1214,In_476);
or U4224 (N_4224,In_14,In_278);
or U4225 (N_4225,In_1226,In_1067);
xnor U4226 (N_4226,In_969,In_85);
nand U4227 (N_4227,In_17,In_310);
xor U4228 (N_4228,In_49,In_1277);
nor U4229 (N_4229,In_1123,In_1468);
nor U4230 (N_4230,In_14,In_1180);
or U4231 (N_4231,In_404,In_451);
nand U4232 (N_4232,In_83,In_91);
nand U4233 (N_4233,In_655,In_646);
or U4234 (N_4234,In_1465,In_989);
nor U4235 (N_4235,In_882,In_426);
xnor U4236 (N_4236,In_413,In_778);
nor U4237 (N_4237,In_112,In_852);
nand U4238 (N_4238,In_1218,In_920);
and U4239 (N_4239,In_1058,In_842);
nor U4240 (N_4240,In_197,In_190);
and U4241 (N_4241,In_29,In_773);
and U4242 (N_4242,In_1315,In_1139);
nor U4243 (N_4243,In_1153,In_524);
or U4244 (N_4244,In_469,In_837);
xor U4245 (N_4245,In_430,In_662);
nand U4246 (N_4246,In_120,In_892);
xor U4247 (N_4247,In_1494,In_1357);
nand U4248 (N_4248,In_8,In_1054);
nor U4249 (N_4249,In_884,In_969);
or U4250 (N_4250,In_437,In_140);
or U4251 (N_4251,In_86,In_981);
xnor U4252 (N_4252,In_1122,In_85);
nand U4253 (N_4253,In_1328,In_723);
or U4254 (N_4254,In_1123,In_732);
and U4255 (N_4255,In_796,In_29);
and U4256 (N_4256,In_1299,In_1010);
or U4257 (N_4257,In_495,In_1116);
or U4258 (N_4258,In_1265,In_309);
or U4259 (N_4259,In_1424,In_971);
and U4260 (N_4260,In_110,In_384);
or U4261 (N_4261,In_1219,In_185);
nand U4262 (N_4262,In_1030,In_1240);
nor U4263 (N_4263,In_17,In_332);
xor U4264 (N_4264,In_1215,In_830);
nand U4265 (N_4265,In_1148,In_925);
or U4266 (N_4266,In_690,In_455);
nand U4267 (N_4267,In_738,In_222);
or U4268 (N_4268,In_1191,In_942);
nor U4269 (N_4269,In_834,In_378);
and U4270 (N_4270,In_433,In_174);
xor U4271 (N_4271,In_1183,In_989);
and U4272 (N_4272,In_1300,In_841);
and U4273 (N_4273,In_951,In_354);
or U4274 (N_4274,In_821,In_723);
xnor U4275 (N_4275,In_990,In_1203);
and U4276 (N_4276,In_282,In_1259);
nor U4277 (N_4277,In_44,In_258);
or U4278 (N_4278,In_771,In_485);
nor U4279 (N_4279,In_804,In_1273);
or U4280 (N_4280,In_342,In_1093);
or U4281 (N_4281,In_872,In_1416);
or U4282 (N_4282,In_589,In_223);
nand U4283 (N_4283,In_763,In_1111);
xnor U4284 (N_4284,In_437,In_379);
or U4285 (N_4285,In_771,In_57);
and U4286 (N_4286,In_842,In_1126);
nand U4287 (N_4287,In_243,In_502);
or U4288 (N_4288,In_114,In_1178);
nand U4289 (N_4289,In_216,In_713);
nor U4290 (N_4290,In_701,In_104);
nand U4291 (N_4291,In_942,In_758);
and U4292 (N_4292,In_850,In_1124);
or U4293 (N_4293,In_574,In_60);
nand U4294 (N_4294,In_416,In_831);
nor U4295 (N_4295,In_216,In_851);
nor U4296 (N_4296,In_289,In_390);
and U4297 (N_4297,In_332,In_110);
or U4298 (N_4298,In_637,In_632);
nor U4299 (N_4299,In_1096,In_1421);
nand U4300 (N_4300,In_226,In_798);
nor U4301 (N_4301,In_588,In_1218);
and U4302 (N_4302,In_140,In_1085);
nand U4303 (N_4303,In_470,In_826);
nand U4304 (N_4304,In_886,In_701);
and U4305 (N_4305,In_800,In_49);
and U4306 (N_4306,In_806,In_718);
nor U4307 (N_4307,In_1252,In_420);
nand U4308 (N_4308,In_1254,In_509);
xor U4309 (N_4309,In_627,In_1384);
and U4310 (N_4310,In_914,In_1183);
xnor U4311 (N_4311,In_554,In_232);
and U4312 (N_4312,In_375,In_768);
and U4313 (N_4313,In_855,In_213);
and U4314 (N_4314,In_1156,In_247);
nor U4315 (N_4315,In_251,In_934);
nor U4316 (N_4316,In_1038,In_880);
xnor U4317 (N_4317,In_48,In_1069);
and U4318 (N_4318,In_1152,In_570);
nor U4319 (N_4319,In_1429,In_118);
nand U4320 (N_4320,In_645,In_342);
and U4321 (N_4321,In_305,In_1332);
or U4322 (N_4322,In_1280,In_741);
xnor U4323 (N_4323,In_1021,In_1339);
nor U4324 (N_4324,In_729,In_295);
and U4325 (N_4325,In_986,In_1408);
or U4326 (N_4326,In_387,In_32);
or U4327 (N_4327,In_319,In_722);
nor U4328 (N_4328,In_611,In_490);
nand U4329 (N_4329,In_1447,In_1173);
xnor U4330 (N_4330,In_291,In_831);
or U4331 (N_4331,In_1420,In_1003);
and U4332 (N_4332,In_568,In_135);
or U4333 (N_4333,In_480,In_994);
nor U4334 (N_4334,In_945,In_860);
or U4335 (N_4335,In_591,In_141);
nor U4336 (N_4336,In_1064,In_980);
xnor U4337 (N_4337,In_970,In_784);
nor U4338 (N_4338,In_1419,In_722);
and U4339 (N_4339,In_1332,In_465);
nor U4340 (N_4340,In_713,In_486);
or U4341 (N_4341,In_851,In_826);
or U4342 (N_4342,In_1173,In_249);
or U4343 (N_4343,In_388,In_435);
or U4344 (N_4344,In_692,In_717);
nor U4345 (N_4345,In_421,In_259);
and U4346 (N_4346,In_1086,In_1187);
nand U4347 (N_4347,In_1218,In_485);
nand U4348 (N_4348,In_429,In_37);
nor U4349 (N_4349,In_590,In_201);
nand U4350 (N_4350,In_655,In_661);
or U4351 (N_4351,In_292,In_392);
xor U4352 (N_4352,In_679,In_1462);
or U4353 (N_4353,In_737,In_1037);
or U4354 (N_4354,In_143,In_1327);
nand U4355 (N_4355,In_1062,In_845);
and U4356 (N_4356,In_530,In_94);
xor U4357 (N_4357,In_890,In_7);
or U4358 (N_4358,In_275,In_301);
and U4359 (N_4359,In_1291,In_585);
nor U4360 (N_4360,In_1180,In_410);
xor U4361 (N_4361,In_145,In_758);
or U4362 (N_4362,In_1156,In_1289);
and U4363 (N_4363,In_77,In_200);
and U4364 (N_4364,In_813,In_1219);
nand U4365 (N_4365,In_114,In_964);
or U4366 (N_4366,In_593,In_312);
or U4367 (N_4367,In_428,In_514);
and U4368 (N_4368,In_392,In_896);
xor U4369 (N_4369,In_142,In_766);
or U4370 (N_4370,In_372,In_721);
xnor U4371 (N_4371,In_1042,In_1172);
nand U4372 (N_4372,In_655,In_1325);
and U4373 (N_4373,In_717,In_1038);
nand U4374 (N_4374,In_1423,In_1128);
or U4375 (N_4375,In_1218,In_860);
nor U4376 (N_4376,In_888,In_1275);
or U4377 (N_4377,In_998,In_945);
nor U4378 (N_4378,In_364,In_256);
nor U4379 (N_4379,In_195,In_1476);
xor U4380 (N_4380,In_1164,In_871);
or U4381 (N_4381,In_452,In_1434);
xor U4382 (N_4382,In_1392,In_871);
nor U4383 (N_4383,In_951,In_9);
nand U4384 (N_4384,In_481,In_193);
nor U4385 (N_4385,In_143,In_1190);
or U4386 (N_4386,In_265,In_798);
or U4387 (N_4387,In_598,In_321);
nor U4388 (N_4388,In_289,In_843);
nor U4389 (N_4389,In_190,In_139);
xnor U4390 (N_4390,In_596,In_705);
and U4391 (N_4391,In_411,In_990);
nand U4392 (N_4392,In_1181,In_985);
and U4393 (N_4393,In_107,In_1002);
nand U4394 (N_4394,In_851,In_686);
nor U4395 (N_4395,In_578,In_1215);
nand U4396 (N_4396,In_1221,In_700);
xnor U4397 (N_4397,In_1380,In_1314);
or U4398 (N_4398,In_557,In_1440);
and U4399 (N_4399,In_1323,In_136);
nor U4400 (N_4400,In_217,In_1224);
nor U4401 (N_4401,In_1027,In_253);
and U4402 (N_4402,In_715,In_505);
nand U4403 (N_4403,In_275,In_325);
nor U4404 (N_4404,In_467,In_264);
nand U4405 (N_4405,In_228,In_525);
and U4406 (N_4406,In_1281,In_359);
nand U4407 (N_4407,In_1416,In_1143);
or U4408 (N_4408,In_567,In_1175);
nor U4409 (N_4409,In_515,In_1441);
and U4410 (N_4410,In_560,In_1440);
and U4411 (N_4411,In_811,In_450);
or U4412 (N_4412,In_408,In_1203);
or U4413 (N_4413,In_1064,In_1161);
nor U4414 (N_4414,In_216,In_549);
nor U4415 (N_4415,In_749,In_220);
or U4416 (N_4416,In_1104,In_1192);
xor U4417 (N_4417,In_149,In_716);
xnor U4418 (N_4418,In_1032,In_1129);
nor U4419 (N_4419,In_1445,In_63);
or U4420 (N_4420,In_654,In_1300);
or U4421 (N_4421,In_325,In_955);
nor U4422 (N_4422,In_64,In_1172);
and U4423 (N_4423,In_461,In_643);
nor U4424 (N_4424,In_1398,In_981);
and U4425 (N_4425,In_712,In_338);
or U4426 (N_4426,In_725,In_369);
nor U4427 (N_4427,In_294,In_1209);
xor U4428 (N_4428,In_286,In_95);
nand U4429 (N_4429,In_139,In_1289);
nor U4430 (N_4430,In_851,In_982);
or U4431 (N_4431,In_76,In_1412);
nand U4432 (N_4432,In_1292,In_604);
nand U4433 (N_4433,In_1202,In_109);
and U4434 (N_4434,In_188,In_1339);
or U4435 (N_4435,In_46,In_1348);
or U4436 (N_4436,In_911,In_298);
nor U4437 (N_4437,In_1446,In_19);
and U4438 (N_4438,In_1317,In_1);
xor U4439 (N_4439,In_1221,In_30);
nand U4440 (N_4440,In_629,In_1471);
nand U4441 (N_4441,In_3,In_1352);
or U4442 (N_4442,In_702,In_977);
nor U4443 (N_4443,In_35,In_1164);
xor U4444 (N_4444,In_936,In_1059);
nor U4445 (N_4445,In_52,In_1036);
nor U4446 (N_4446,In_210,In_151);
and U4447 (N_4447,In_1244,In_643);
nand U4448 (N_4448,In_1215,In_476);
or U4449 (N_4449,In_337,In_77);
or U4450 (N_4450,In_281,In_1495);
nor U4451 (N_4451,In_370,In_276);
or U4452 (N_4452,In_919,In_683);
nor U4453 (N_4453,In_265,In_987);
and U4454 (N_4454,In_1044,In_92);
nand U4455 (N_4455,In_1399,In_45);
nor U4456 (N_4456,In_12,In_339);
xor U4457 (N_4457,In_167,In_391);
nor U4458 (N_4458,In_41,In_275);
nand U4459 (N_4459,In_707,In_1273);
xor U4460 (N_4460,In_1201,In_822);
nand U4461 (N_4461,In_3,In_1165);
or U4462 (N_4462,In_644,In_503);
and U4463 (N_4463,In_57,In_89);
nor U4464 (N_4464,In_728,In_1316);
nor U4465 (N_4465,In_460,In_981);
and U4466 (N_4466,In_568,In_588);
and U4467 (N_4467,In_1314,In_1282);
or U4468 (N_4468,In_718,In_304);
and U4469 (N_4469,In_890,In_739);
and U4470 (N_4470,In_582,In_1317);
xnor U4471 (N_4471,In_459,In_869);
nand U4472 (N_4472,In_1119,In_1448);
or U4473 (N_4473,In_184,In_1166);
or U4474 (N_4474,In_182,In_403);
nand U4475 (N_4475,In_240,In_968);
and U4476 (N_4476,In_467,In_4);
or U4477 (N_4477,In_877,In_85);
nor U4478 (N_4478,In_535,In_1239);
nor U4479 (N_4479,In_612,In_1028);
or U4480 (N_4480,In_1144,In_382);
and U4481 (N_4481,In_363,In_1205);
nor U4482 (N_4482,In_795,In_1129);
nand U4483 (N_4483,In_155,In_1026);
nor U4484 (N_4484,In_1192,In_960);
and U4485 (N_4485,In_884,In_910);
nand U4486 (N_4486,In_70,In_75);
xor U4487 (N_4487,In_1478,In_1343);
nor U4488 (N_4488,In_969,In_373);
nand U4489 (N_4489,In_635,In_1349);
or U4490 (N_4490,In_867,In_9);
and U4491 (N_4491,In_155,In_310);
nand U4492 (N_4492,In_719,In_182);
nor U4493 (N_4493,In_461,In_926);
nand U4494 (N_4494,In_24,In_934);
nor U4495 (N_4495,In_472,In_1337);
xor U4496 (N_4496,In_1058,In_641);
or U4497 (N_4497,In_483,In_376);
nor U4498 (N_4498,In_681,In_972);
and U4499 (N_4499,In_618,In_69);
or U4500 (N_4500,In_42,In_228);
nor U4501 (N_4501,In_758,In_330);
nand U4502 (N_4502,In_904,In_99);
or U4503 (N_4503,In_340,In_1495);
nor U4504 (N_4504,In_116,In_22);
nor U4505 (N_4505,In_44,In_1277);
and U4506 (N_4506,In_964,In_995);
or U4507 (N_4507,In_1246,In_544);
nand U4508 (N_4508,In_1183,In_555);
nand U4509 (N_4509,In_1230,In_111);
nand U4510 (N_4510,In_623,In_1415);
and U4511 (N_4511,In_270,In_559);
and U4512 (N_4512,In_372,In_984);
or U4513 (N_4513,In_268,In_579);
nand U4514 (N_4514,In_445,In_922);
nor U4515 (N_4515,In_1068,In_688);
nor U4516 (N_4516,In_391,In_696);
nand U4517 (N_4517,In_142,In_202);
or U4518 (N_4518,In_1314,In_450);
or U4519 (N_4519,In_1136,In_1370);
or U4520 (N_4520,In_40,In_885);
and U4521 (N_4521,In_245,In_491);
nor U4522 (N_4522,In_1321,In_788);
xnor U4523 (N_4523,In_327,In_432);
nand U4524 (N_4524,In_1200,In_1084);
or U4525 (N_4525,In_1014,In_1108);
xor U4526 (N_4526,In_1277,In_1479);
nand U4527 (N_4527,In_1110,In_879);
nor U4528 (N_4528,In_939,In_437);
or U4529 (N_4529,In_1098,In_843);
or U4530 (N_4530,In_771,In_826);
nand U4531 (N_4531,In_127,In_305);
nand U4532 (N_4532,In_308,In_421);
nor U4533 (N_4533,In_553,In_1289);
nand U4534 (N_4534,In_404,In_264);
or U4535 (N_4535,In_753,In_841);
or U4536 (N_4536,In_133,In_598);
nor U4537 (N_4537,In_1463,In_1466);
nor U4538 (N_4538,In_850,In_1233);
nand U4539 (N_4539,In_1086,In_1194);
xor U4540 (N_4540,In_1336,In_1277);
and U4541 (N_4541,In_1016,In_1147);
nor U4542 (N_4542,In_683,In_1029);
or U4543 (N_4543,In_1051,In_609);
and U4544 (N_4544,In_519,In_774);
nand U4545 (N_4545,In_262,In_783);
nor U4546 (N_4546,In_208,In_1263);
and U4547 (N_4547,In_132,In_720);
nor U4548 (N_4548,In_991,In_867);
nand U4549 (N_4549,In_62,In_104);
nor U4550 (N_4550,In_870,In_686);
xor U4551 (N_4551,In_208,In_815);
and U4552 (N_4552,In_431,In_1435);
or U4553 (N_4553,In_1162,In_127);
nand U4554 (N_4554,In_1218,In_753);
or U4555 (N_4555,In_1057,In_769);
or U4556 (N_4556,In_173,In_1491);
and U4557 (N_4557,In_520,In_1005);
nand U4558 (N_4558,In_491,In_192);
nor U4559 (N_4559,In_1349,In_651);
nand U4560 (N_4560,In_888,In_303);
or U4561 (N_4561,In_1332,In_193);
or U4562 (N_4562,In_604,In_1413);
xor U4563 (N_4563,In_258,In_1058);
nor U4564 (N_4564,In_407,In_18);
nand U4565 (N_4565,In_567,In_994);
nand U4566 (N_4566,In_497,In_639);
nor U4567 (N_4567,In_1472,In_1411);
xnor U4568 (N_4568,In_353,In_966);
or U4569 (N_4569,In_1437,In_785);
or U4570 (N_4570,In_950,In_435);
or U4571 (N_4571,In_466,In_461);
nor U4572 (N_4572,In_139,In_705);
or U4573 (N_4573,In_836,In_1407);
nand U4574 (N_4574,In_626,In_325);
or U4575 (N_4575,In_1468,In_1142);
nor U4576 (N_4576,In_141,In_64);
nor U4577 (N_4577,In_1218,In_740);
nand U4578 (N_4578,In_814,In_1174);
and U4579 (N_4579,In_549,In_764);
xnor U4580 (N_4580,In_643,In_437);
nor U4581 (N_4581,In_1285,In_1427);
nand U4582 (N_4582,In_288,In_422);
nand U4583 (N_4583,In_1309,In_858);
and U4584 (N_4584,In_600,In_1280);
and U4585 (N_4585,In_243,In_968);
xnor U4586 (N_4586,In_888,In_998);
nor U4587 (N_4587,In_1443,In_1136);
nand U4588 (N_4588,In_1090,In_49);
nand U4589 (N_4589,In_742,In_1278);
xnor U4590 (N_4590,In_136,In_950);
and U4591 (N_4591,In_87,In_98);
nor U4592 (N_4592,In_1233,In_619);
nor U4593 (N_4593,In_247,In_918);
or U4594 (N_4594,In_1243,In_335);
and U4595 (N_4595,In_1033,In_72);
or U4596 (N_4596,In_1183,In_880);
or U4597 (N_4597,In_691,In_802);
and U4598 (N_4598,In_434,In_321);
nor U4599 (N_4599,In_26,In_347);
nor U4600 (N_4600,In_1442,In_980);
or U4601 (N_4601,In_1497,In_306);
or U4602 (N_4602,In_187,In_902);
and U4603 (N_4603,In_970,In_1265);
and U4604 (N_4604,In_175,In_1330);
or U4605 (N_4605,In_995,In_1370);
nor U4606 (N_4606,In_1346,In_132);
or U4607 (N_4607,In_958,In_1401);
or U4608 (N_4608,In_696,In_1044);
nand U4609 (N_4609,In_748,In_557);
nor U4610 (N_4610,In_658,In_1260);
and U4611 (N_4611,In_1231,In_431);
nor U4612 (N_4612,In_1059,In_1212);
and U4613 (N_4613,In_1017,In_950);
nand U4614 (N_4614,In_613,In_1384);
and U4615 (N_4615,In_1464,In_1453);
nand U4616 (N_4616,In_1123,In_234);
nor U4617 (N_4617,In_738,In_1354);
nand U4618 (N_4618,In_1374,In_485);
or U4619 (N_4619,In_1124,In_1424);
and U4620 (N_4620,In_1291,In_636);
nand U4621 (N_4621,In_686,In_211);
and U4622 (N_4622,In_840,In_754);
and U4623 (N_4623,In_693,In_330);
or U4624 (N_4624,In_1053,In_662);
nor U4625 (N_4625,In_1123,In_973);
and U4626 (N_4626,In_210,In_783);
and U4627 (N_4627,In_464,In_484);
xnor U4628 (N_4628,In_237,In_68);
and U4629 (N_4629,In_451,In_600);
and U4630 (N_4630,In_1184,In_122);
and U4631 (N_4631,In_1345,In_1419);
nand U4632 (N_4632,In_1368,In_581);
xor U4633 (N_4633,In_66,In_31);
nand U4634 (N_4634,In_283,In_276);
and U4635 (N_4635,In_1123,In_678);
or U4636 (N_4636,In_881,In_134);
xor U4637 (N_4637,In_718,In_1336);
nor U4638 (N_4638,In_1270,In_408);
and U4639 (N_4639,In_88,In_718);
nor U4640 (N_4640,In_284,In_500);
nor U4641 (N_4641,In_1211,In_471);
or U4642 (N_4642,In_1114,In_1475);
or U4643 (N_4643,In_1165,In_499);
and U4644 (N_4644,In_1477,In_577);
or U4645 (N_4645,In_506,In_438);
nor U4646 (N_4646,In_1180,In_33);
xor U4647 (N_4647,In_1362,In_790);
nand U4648 (N_4648,In_421,In_534);
xor U4649 (N_4649,In_835,In_1136);
nand U4650 (N_4650,In_1364,In_1482);
or U4651 (N_4651,In_517,In_966);
and U4652 (N_4652,In_392,In_765);
nand U4653 (N_4653,In_1417,In_1260);
nand U4654 (N_4654,In_804,In_735);
and U4655 (N_4655,In_980,In_1172);
or U4656 (N_4656,In_1322,In_1488);
nand U4657 (N_4657,In_1427,In_552);
or U4658 (N_4658,In_624,In_306);
or U4659 (N_4659,In_1203,In_580);
nor U4660 (N_4660,In_1245,In_287);
nand U4661 (N_4661,In_890,In_801);
or U4662 (N_4662,In_414,In_672);
nor U4663 (N_4663,In_121,In_756);
and U4664 (N_4664,In_947,In_41);
and U4665 (N_4665,In_1406,In_618);
and U4666 (N_4666,In_590,In_1433);
nand U4667 (N_4667,In_988,In_391);
nor U4668 (N_4668,In_31,In_1147);
nand U4669 (N_4669,In_630,In_162);
and U4670 (N_4670,In_422,In_1020);
and U4671 (N_4671,In_1182,In_97);
nand U4672 (N_4672,In_236,In_469);
and U4673 (N_4673,In_1291,In_1327);
or U4674 (N_4674,In_1280,In_1461);
nor U4675 (N_4675,In_220,In_882);
or U4676 (N_4676,In_213,In_1424);
or U4677 (N_4677,In_914,In_893);
or U4678 (N_4678,In_308,In_1497);
or U4679 (N_4679,In_1055,In_1346);
nor U4680 (N_4680,In_1119,In_663);
or U4681 (N_4681,In_644,In_707);
nand U4682 (N_4682,In_245,In_980);
xor U4683 (N_4683,In_911,In_352);
xor U4684 (N_4684,In_605,In_1259);
xor U4685 (N_4685,In_1180,In_1155);
and U4686 (N_4686,In_893,In_901);
nand U4687 (N_4687,In_218,In_30);
xor U4688 (N_4688,In_1344,In_119);
nand U4689 (N_4689,In_548,In_561);
or U4690 (N_4690,In_918,In_186);
and U4691 (N_4691,In_684,In_863);
nor U4692 (N_4692,In_934,In_939);
and U4693 (N_4693,In_1244,In_154);
nor U4694 (N_4694,In_1097,In_801);
nor U4695 (N_4695,In_676,In_160);
or U4696 (N_4696,In_1068,In_1083);
nand U4697 (N_4697,In_1336,In_1404);
nand U4698 (N_4698,In_711,In_907);
xnor U4699 (N_4699,In_295,In_761);
and U4700 (N_4700,In_1030,In_1311);
nand U4701 (N_4701,In_1111,In_652);
nor U4702 (N_4702,In_876,In_1250);
nor U4703 (N_4703,In_413,In_393);
nand U4704 (N_4704,In_117,In_1039);
and U4705 (N_4705,In_642,In_145);
and U4706 (N_4706,In_1128,In_1412);
or U4707 (N_4707,In_152,In_442);
nand U4708 (N_4708,In_1366,In_274);
and U4709 (N_4709,In_408,In_1276);
nand U4710 (N_4710,In_1440,In_1011);
and U4711 (N_4711,In_1031,In_650);
and U4712 (N_4712,In_1109,In_601);
xnor U4713 (N_4713,In_212,In_641);
or U4714 (N_4714,In_1231,In_506);
nand U4715 (N_4715,In_71,In_352);
nor U4716 (N_4716,In_613,In_214);
and U4717 (N_4717,In_326,In_793);
and U4718 (N_4718,In_785,In_1310);
nor U4719 (N_4719,In_613,In_1096);
and U4720 (N_4720,In_105,In_418);
xor U4721 (N_4721,In_1253,In_1468);
and U4722 (N_4722,In_45,In_984);
and U4723 (N_4723,In_1000,In_463);
xnor U4724 (N_4724,In_986,In_1028);
and U4725 (N_4725,In_1100,In_74);
and U4726 (N_4726,In_592,In_350);
nand U4727 (N_4727,In_796,In_1441);
or U4728 (N_4728,In_1028,In_1112);
nor U4729 (N_4729,In_177,In_468);
nor U4730 (N_4730,In_1394,In_320);
or U4731 (N_4731,In_1397,In_1367);
xor U4732 (N_4732,In_1464,In_1343);
or U4733 (N_4733,In_854,In_1300);
nor U4734 (N_4734,In_595,In_1193);
and U4735 (N_4735,In_1319,In_498);
or U4736 (N_4736,In_433,In_1351);
or U4737 (N_4737,In_982,In_1457);
or U4738 (N_4738,In_1494,In_478);
and U4739 (N_4739,In_572,In_1193);
or U4740 (N_4740,In_1476,In_629);
nor U4741 (N_4741,In_973,In_704);
nand U4742 (N_4742,In_312,In_1006);
xor U4743 (N_4743,In_1203,In_1175);
and U4744 (N_4744,In_730,In_608);
or U4745 (N_4745,In_1278,In_316);
nand U4746 (N_4746,In_599,In_1325);
or U4747 (N_4747,In_933,In_1074);
nor U4748 (N_4748,In_278,In_156);
nor U4749 (N_4749,In_129,In_320);
or U4750 (N_4750,In_1497,In_1083);
or U4751 (N_4751,In_771,In_919);
nand U4752 (N_4752,In_52,In_211);
and U4753 (N_4753,In_106,In_258);
nor U4754 (N_4754,In_1026,In_506);
nand U4755 (N_4755,In_1182,In_237);
and U4756 (N_4756,In_1257,In_330);
or U4757 (N_4757,In_1371,In_1268);
nor U4758 (N_4758,In_879,In_686);
nor U4759 (N_4759,In_335,In_1138);
or U4760 (N_4760,In_692,In_491);
and U4761 (N_4761,In_966,In_1293);
nor U4762 (N_4762,In_550,In_1490);
and U4763 (N_4763,In_1479,In_470);
nand U4764 (N_4764,In_15,In_765);
and U4765 (N_4765,In_80,In_605);
and U4766 (N_4766,In_738,In_1240);
and U4767 (N_4767,In_101,In_1056);
and U4768 (N_4768,In_698,In_606);
nor U4769 (N_4769,In_274,In_743);
nor U4770 (N_4770,In_710,In_274);
nand U4771 (N_4771,In_606,In_701);
nand U4772 (N_4772,In_1244,In_1042);
nand U4773 (N_4773,In_1129,In_408);
nand U4774 (N_4774,In_695,In_483);
or U4775 (N_4775,In_311,In_587);
xnor U4776 (N_4776,In_342,In_1178);
nand U4777 (N_4777,In_1420,In_1014);
nor U4778 (N_4778,In_653,In_181);
nand U4779 (N_4779,In_1446,In_103);
and U4780 (N_4780,In_220,In_107);
and U4781 (N_4781,In_624,In_116);
nor U4782 (N_4782,In_40,In_385);
nor U4783 (N_4783,In_102,In_1385);
nand U4784 (N_4784,In_341,In_4);
or U4785 (N_4785,In_1486,In_256);
xor U4786 (N_4786,In_13,In_631);
or U4787 (N_4787,In_71,In_609);
or U4788 (N_4788,In_442,In_229);
nand U4789 (N_4789,In_543,In_933);
nor U4790 (N_4790,In_1342,In_592);
xor U4791 (N_4791,In_342,In_71);
xnor U4792 (N_4792,In_1193,In_213);
or U4793 (N_4793,In_743,In_254);
nor U4794 (N_4794,In_832,In_460);
nor U4795 (N_4795,In_915,In_722);
nand U4796 (N_4796,In_618,In_77);
and U4797 (N_4797,In_869,In_155);
xnor U4798 (N_4798,In_741,In_498);
or U4799 (N_4799,In_975,In_629);
nor U4800 (N_4800,In_348,In_297);
and U4801 (N_4801,In_177,In_76);
and U4802 (N_4802,In_1474,In_944);
nand U4803 (N_4803,In_272,In_369);
nor U4804 (N_4804,In_141,In_1227);
or U4805 (N_4805,In_583,In_59);
xor U4806 (N_4806,In_1327,In_287);
and U4807 (N_4807,In_350,In_463);
nor U4808 (N_4808,In_638,In_370);
and U4809 (N_4809,In_127,In_387);
xor U4810 (N_4810,In_802,In_171);
nand U4811 (N_4811,In_952,In_580);
or U4812 (N_4812,In_10,In_745);
and U4813 (N_4813,In_403,In_535);
xnor U4814 (N_4814,In_407,In_200);
or U4815 (N_4815,In_383,In_512);
nor U4816 (N_4816,In_828,In_1091);
and U4817 (N_4817,In_377,In_22);
or U4818 (N_4818,In_756,In_1129);
or U4819 (N_4819,In_460,In_728);
or U4820 (N_4820,In_679,In_1383);
and U4821 (N_4821,In_591,In_726);
xnor U4822 (N_4822,In_205,In_926);
nand U4823 (N_4823,In_582,In_1047);
nand U4824 (N_4824,In_1470,In_1011);
nand U4825 (N_4825,In_473,In_1312);
nand U4826 (N_4826,In_829,In_619);
xnor U4827 (N_4827,In_981,In_1183);
nand U4828 (N_4828,In_550,In_1164);
nand U4829 (N_4829,In_874,In_1111);
nand U4830 (N_4830,In_477,In_1478);
nor U4831 (N_4831,In_754,In_246);
nand U4832 (N_4832,In_1327,In_509);
and U4833 (N_4833,In_1041,In_914);
nor U4834 (N_4834,In_1210,In_308);
or U4835 (N_4835,In_599,In_1351);
nor U4836 (N_4836,In_937,In_230);
nor U4837 (N_4837,In_555,In_1368);
and U4838 (N_4838,In_893,In_399);
nor U4839 (N_4839,In_216,In_315);
and U4840 (N_4840,In_952,In_1431);
xnor U4841 (N_4841,In_360,In_1259);
nand U4842 (N_4842,In_512,In_248);
and U4843 (N_4843,In_487,In_1394);
nor U4844 (N_4844,In_628,In_1044);
xnor U4845 (N_4845,In_669,In_172);
and U4846 (N_4846,In_822,In_86);
xnor U4847 (N_4847,In_791,In_1051);
nand U4848 (N_4848,In_770,In_1330);
nand U4849 (N_4849,In_1431,In_830);
nand U4850 (N_4850,In_553,In_1005);
nand U4851 (N_4851,In_386,In_195);
nor U4852 (N_4852,In_1378,In_1187);
nor U4853 (N_4853,In_241,In_1301);
and U4854 (N_4854,In_758,In_1327);
nand U4855 (N_4855,In_107,In_1198);
nor U4856 (N_4856,In_179,In_1231);
xor U4857 (N_4857,In_803,In_525);
nand U4858 (N_4858,In_1310,In_763);
or U4859 (N_4859,In_36,In_1183);
xnor U4860 (N_4860,In_554,In_147);
nand U4861 (N_4861,In_575,In_915);
or U4862 (N_4862,In_182,In_757);
or U4863 (N_4863,In_1224,In_851);
or U4864 (N_4864,In_1485,In_214);
and U4865 (N_4865,In_533,In_17);
nor U4866 (N_4866,In_1316,In_1378);
and U4867 (N_4867,In_46,In_1293);
and U4868 (N_4868,In_359,In_72);
nor U4869 (N_4869,In_1098,In_1021);
or U4870 (N_4870,In_579,In_989);
xnor U4871 (N_4871,In_1245,In_826);
nor U4872 (N_4872,In_872,In_981);
and U4873 (N_4873,In_1104,In_771);
nor U4874 (N_4874,In_492,In_1307);
nor U4875 (N_4875,In_928,In_769);
nand U4876 (N_4876,In_1281,In_1169);
and U4877 (N_4877,In_345,In_524);
nor U4878 (N_4878,In_777,In_1344);
nand U4879 (N_4879,In_1151,In_1424);
and U4880 (N_4880,In_80,In_153);
nor U4881 (N_4881,In_342,In_459);
nor U4882 (N_4882,In_55,In_1267);
nand U4883 (N_4883,In_1066,In_57);
nor U4884 (N_4884,In_1304,In_1364);
and U4885 (N_4885,In_797,In_231);
xnor U4886 (N_4886,In_1149,In_644);
nand U4887 (N_4887,In_1146,In_803);
and U4888 (N_4888,In_275,In_326);
nor U4889 (N_4889,In_662,In_874);
nand U4890 (N_4890,In_1399,In_882);
xor U4891 (N_4891,In_971,In_1130);
and U4892 (N_4892,In_886,In_378);
or U4893 (N_4893,In_724,In_942);
nand U4894 (N_4894,In_30,In_784);
and U4895 (N_4895,In_708,In_895);
xnor U4896 (N_4896,In_678,In_55);
xnor U4897 (N_4897,In_836,In_608);
or U4898 (N_4898,In_58,In_808);
nor U4899 (N_4899,In_1180,In_646);
nor U4900 (N_4900,In_830,In_1161);
nor U4901 (N_4901,In_715,In_476);
nor U4902 (N_4902,In_1236,In_1001);
and U4903 (N_4903,In_66,In_631);
nand U4904 (N_4904,In_1470,In_885);
and U4905 (N_4905,In_85,In_10);
and U4906 (N_4906,In_349,In_263);
nor U4907 (N_4907,In_886,In_1011);
nor U4908 (N_4908,In_1217,In_108);
nand U4909 (N_4909,In_789,In_1494);
nor U4910 (N_4910,In_112,In_841);
nand U4911 (N_4911,In_366,In_780);
nand U4912 (N_4912,In_235,In_444);
or U4913 (N_4913,In_10,In_701);
nor U4914 (N_4914,In_954,In_782);
nor U4915 (N_4915,In_1285,In_983);
nor U4916 (N_4916,In_798,In_417);
nor U4917 (N_4917,In_29,In_684);
nor U4918 (N_4918,In_370,In_785);
nand U4919 (N_4919,In_501,In_465);
xor U4920 (N_4920,In_1321,In_608);
nor U4921 (N_4921,In_1428,In_394);
or U4922 (N_4922,In_1160,In_388);
and U4923 (N_4923,In_1075,In_1219);
nand U4924 (N_4924,In_1119,In_1031);
nor U4925 (N_4925,In_712,In_729);
nand U4926 (N_4926,In_1100,In_776);
nand U4927 (N_4927,In_281,In_1077);
xor U4928 (N_4928,In_65,In_1230);
and U4929 (N_4929,In_1392,In_311);
nor U4930 (N_4930,In_775,In_610);
nor U4931 (N_4931,In_275,In_883);
nor U4932 (N_4932,In_524,In_323);
and U4933 (N_4933,In_572,In_523);
and U4934 (N_4934,In_802,In_1150);
nand U4935 (N_4935,In_868,In_365);
nor U4936 (N_4936,In_740,In_575);
and U4937 (N_4937,In_573,In_724);
nand U4938 (N_4938,In_1169,In_58);
nor U4939 (N_4939,In_857,In_90);
nor U4940 (N_4940,In_1361,In_1385);
or U4941 (N_4941,In_681,In_1382);
xor U4942 (N_4942,In_515,In_1068);
nor U4943 (N_4943,In_1458,In_50);
nand U4944 (N_4944,In_595,In_194);
or U4945 (N_4945,In_326,In_1019);
nor U4946 (N_4946,In_571,In_1335);
or U4947 (N_4947,In_701,In_76);
nand U4948 (N_4948,In_1021,In_975);
nand U4949 (N_4949,In_236,In_625);
nor U4950 (N_4950,In_295,In_668);
nand U4951 (N_4951,In_47,In_1135);
or U4952 (N_4952,In_1346,In_765);
nand U4953 (N_4953,In_471,In_365);
xor U4954 (N_4954,In_1363,In_615);
or U4955 (N_4955,In_139,In_444);
or U4956 (N_4956,In_885,In_559);
and U4957 (N_4957,In_818,In_416);
nand U4958 (N_4958,In_364,In_208);
and U4959 (N_4959,In_1407,In_987);
nor U4960 (N_4960,In_1110,In_1271);
nor U4961 (N_4961,In_694,In_386);
xnor U4962 (N_4962,In_250,In_1480);
and U4963 (N_4963,In_359,In_1015);
and U4964 (N_4964,In_139,In_583);
and U4965 (N_4965,In_1123,In_20);
nor U4966 (N_4966,In_379,In_84);
or U4967 (N_4967,In_594,In_800);
or U4968 (N_4968,In_253,In_624);
nor U4969 (N_4969,In_703,In_1309);
xor U4970 (N_4970,In_143,In_1340);
or U4971 (N_4971,In_995,In_1006);
or U4972 (N_4972,In_254,In_1400);
and U4973 (N_4973,In_1008,In_485);
nor U4974 (N_4974,In_1284,In_463);
and U4975 (N_4975,In_817,In_1420);
nor U4976 (N_4976,In_489,In_308);
and U4977 (N_4977,In_560,In_150);
nor U4978 (N_4978,In_862,In_1005);
or U4979 (N_4979,In_1188,In_530);
and U4980 (N_4980,In_479,In_541);
or U4981 (N_4981,In_1499,In_1457);
nand U4982 (N_4982,In_505,In_154);
or U4983 (N_4983,In_165,In_1123);
nand U4984 (N_4984,In_955,In_447);
nand U4985 (N_4985,In_970,In_907);
nor U4986 (N_4986,In_646,In_1101);
xor U4987 (N_4987,In_91,In_1337);
and U4988 (N_4988,In_647,In_71);
and U4989 (N_4989,In_713,In_612);
and U4990 (N_4990,In_781,In_1305);
or U4991 (N_4991,In_963,In_1182);
nor U4992 (N_4992,In_809,In_634);
nand U4993 (N_4993,In_361,In_179);
nand U4994 (N_4994,In_895,In_523);
nor U4995 (N_4995,In_878,In_612);
nor U4996 (N_4996,In_201,In_741);
or U4997 (N_4997,In_1327,In_1074);
nor U4998 (N_4998,In_1128,In_445);
nor U4999 (N_4999,In_1412,In_148);
nand U5000 (N_5000,N_4355,N_3995);
nor U5001 (N_5001,N_4460,N_871);
nand U5002 (N_5002,N_1283,N_731);
and U5003 (N_5003,N_4114,N_2721);
nand U5004 (N_5004,N_2481,N_1463);
nor U5005 (N_5005,N_2769,N_3805);
nor U5006 (N_5006,N_1530,N_1426);
and U5007 (N_5007,N_941,N_225);
and U5008 (N_5008,N_3479,N_1121);
or U5009 (N_5009,N_4428,N_4280);
or U5010 (N_5010,N_1152,N_1851);
and U5011 (N_5011,N_3169,N_3411);
nor U5012 (N_5012,N_2646,N_3790);
xnor U5013 (N_5013,N_3903,N_1630);
xnor U5014 (N_5014,N_4394,N_1303);
xnor U5015 (N_5015,N_84,N_1313);
or U5016 (N_5016,N_1474,N_3308);
or U5017 (N_5017,N_2904,N_1963);
or U5018 (N_5018,N_3958,N_1904);
nor U5019 (N_5019,N_3293,N_541);
or U5020 (N_5020,N_3088,N_2622);
nand U5021 (N_5021,N_1064,N_750);
nor U5022 (N_5022,N_2147,N_3094);
nand U5023 (N_5023,N_2619,N_4604);
or U5024 (N_5024,N_2324,N_3077);
nor U5025 (N_5025,N_1621,N_4470);
or U5026 (N_5026,N_957,N_3609);
or U5027 (N_5027,N_105,N_2400);
nand U5028 (N_5028,N_2239,N_4313);
nand U5029 (N_5029,N_949,N_494);
or U5030 (N_5030,N_102,N_2033);
nor U5031 (N_5031,N_2060,N_4733);
nand U5032 (N_5032,N_2031,N_798);
and U5033 (N_5033,N_276,N_4501);
or U5034 (N_5034,N_3643,N_1437);
nor U5035 (N_5035,N_2449,N_470);
nor U5036 (N_5036,N_479,N_1113);
nand U5037 (N_5037,N_1031,N_2531);
or U5038 (N_5038,N_2885,N_2253);
nor U5039 (N_5039,N_1584,N_698);
nand U5040 (N_5040,N_3416,N_2386);
xnor U5041 (N_5041,N_1163,N_70);
nor U5042 (N_5042,N_625,N_4621);
nor U5043 (N_5043,N_2151,N_725);
nand U5044 (N_5044,N_4231,N_521);
xor U5045 (N_5045,N_744,N_751);
or U5046 (N_5046,N_637,N_4830);
or U5047 (N_5047,N_4268,N_4776);
nor U5048 (N_5048,N_621,N_4459);
nand U5049 (N_5049,N_415,N_4788);
nand U5050 (N_5050,N_1854,N_4796);
xor U5051 (N_5051,N_4906,N_962);
xor U5052 (N_5052,N_3567,N_4671);
nor U5053 (N_5053,N_4689,N_47);
nor U5054 (N_5054,N_3671,N_2550);
nor U5055 (N_5055,N_1914,N_2879);
nand U5056 (N_5056,N_431,N_2791);
nor U5057 (N_5057,N_2077,N_4082);
or U5058 (N_5058,N_627,N_2633);
or U5059 (N_5059,N_2698,N_3906);
and U5060 (N_5060,N_4681,N_1766);
and U5061 (N_5061,N_3905,N_1439);
nor U5062 (N_5062,N_1485,N_1716);
and U5063 (N_5063,N_1061,N_1883);
or U5064 (N_5064,N_4132,N_1550);
xor U5065 (N_5065,N_667,N_3371);
or U5066 (N_5066,N_3277,N_1098);
xor U5067 (N_5067,N_151,N_2639);
or U5068 (N_5068,N_2547,N_224);
nand U5069 (N_5069,N_3864,N_620);
and U5070 (N_5070,N_3190,N_1328);
or U5071 (N_5071,N_62,N_179);
nor U5072 (N_5072,N_2385,N_1398);
or U5073 (N_5073,N_2997,N_4543);
nand U5074 (N_5074,N_3737,N_86);
nand U5075 (N_5075,N_3355,N_15);
nand U5076 (N_5076,N_707,N_3381);
nor U5077 (N_5077,N_1724,N_2482);
nand U5078 (N_5078,N_1441,N_4287);
nand U5079 (N_5079,N_868,N_3276);
nand U5080 (N_5080,N_3608,N_3564);
or U5081 (N_5081,N_1862,N_1711);
xor U5082 (N_5082,N_4163,N_2659);
and U5083 (N_5083,N_531,N_2073);
nor U5084 (N_5084,N_4016,N_101);
or U5085 (N_5085,N_2264,N_4805);
nand U5086 (N_5086,N_1882,N_168);
or U5087 (N_5087,N_1381,N_1351);
xnor U5088 (N_5088,N_1772,N_2590);
nor U5089 (N_5089,N_3532,N_1105);
nor U5090 (N_5090,N_480,N_2676);
nor U5091 (N_5091,N_203,N_356);
nor U5092 (N_5092,N_8,N_4602);
xnor U5093 (N_5093,N_4263,N_3366);
and U5094 (N_5094,N_898,N_1989);
xor U5095 (N_5095,N_4236,N_2949);
nor U5096 (N_5096,N_1935,N_2971);
and U5097 (N_5097,N_443,N_2237);
or U5098 (N_5098,N_1145,N_742);
nor U5099 (N_5099,N_1785,N_40);
nor U5100 (N_5100,N_1449,N_4122);
or U5101 (N_5101,N_2412,N_797);
and U5102 (N_5102,N_97,N_1130);
or U5103 (N_5103,N_1401,N_2394);
and U5104 (N_5104,N_2198,N_2605);
or U5105 (N_5105,N_3358,N_1900);
nand U5106 (N_5106,N_2476,N_4749);
or U5107 (N_5107,N_3345,N_2323);
nor U5108 (N_5108,N_1305,N_3288);
nor U5109 (N_5109,N_3876,N_4932);
nand U5110 (N_5110,N_25,N_2325);
or U5111 (N_5111,N_4712,N_2133);
and U5112 (N_5112,N_4102,N_4870);
nor U5113 (N_5113,N_4068,N_2469);
nor U5114 (N_5114,N_807,N_4477);
or U5115 (N_5115,N_3114,N_1765);
or U5116 (N_5116,N_1033,N_1985);
or U5117 (N_5117,N_3710,N_4304);
or U5118 (N_5118,N_1206,N_4503);
nor U5119 (N_5119,N_410,N_1270);
nor U5120 (N_5120,N_2192,N_688);
nor U5121 (N_5121,N_3986,N_1216);
or U5122 (N_5122,N_4786,N_3880);
nor U5123 (N_5123,N_2629,N_4195);
nand U5124 (N_5124,N_2780,N_808);
nand U5125 (N_5125,N_1135,N_309);
and U5126 (N_5126,N_4869,N_4553);
nand U5127 (N_5127,N_788,N_2760);
and U5128 (N_5128,N_749,N_349);
and U5129 (N_5129,N_2947,N_1175);
or U5130 (N_5130,N_1660,N_3560);
or U5131 (N_5131,N_220,N_2085);
and U5132 (N_5132,N_2899,N_3705);
nand U5133 (N_5133,N_3550,N_3424);
nor U5134 (N_5134,N_4617,N_1694);
and U5135 (N_5135,N_635,N_4837);
nand U5136 (N_5136,N_4374,N_839);
xor U5137 (N_5137,N_614,N_230);
or U5138 (N_5138,N_1198,N_3573);
and U5139 (N_5139,N_3350,N_1);
nand U5140 (N_5140,N_2913,N_2078);
nor U5141 (N_5141,N_3212,N_2195);
and U5142 (N_5142,N_2992,N_3744);
or U5143 (N_5143,N_1992,N_2110);
nor U5144 (N_5144,N_4444,N_4532);
or U5145 (N_5145,N_3534,N_3193);
or U5146 (N_5146,N_4522,N_1495);
xor U5147 (N_5147,N_1295,N_558);
nor U5148 (N_5148,N_131,N_2);
or U5149 (N_5149,N_1492,N_640);
and U5150 (N_5150,N_3160,N_74);
nand U5151 (N_5151,N_2932,N_4357);
nor U5152 (N_5152,N_2082,N_2240);
nand U5153 (N_5153,N_1258,N_3227);
and U5154 (N_5154,N_607,N_4341);
nand U5155 (N_5155,N_3758,N_4884);
or U5156 (N_5156,N_1693,N_3156);
and U5157 (N_5157,N_2431,N_2361);
or U5158 (N_5158,N_3920,N_653);
xor U5159 (N_5159,N_2834,N_1170);
or U5160 (N_5160,N_3289,N_124);
xor U5161 (N_5161,N_1301,N_910);
and U5162 (N_5162,N_540,N_263);
or U5163 (N_5163,N_3523,N_2528);
and U5164 (N_5164,N_3654,N_4111);
and U5165 (N_5165,N_3976,N_4743);
or U5166 (N_5166,N_1435,N_3044);
nor U5167 (N_5167,N_774,N_3271);
nor U5168 (N_5168,N_1235,N_365);
nand U5169 (N_5169,N_4990,N_2084);
nor U5170 (N_5170,N_1897,N_1013);
nor U5171 (N_5171,N_4073,N_1060);
xnor U5172 (N_5172,N_2076,N_905);
or U5173 (N_5173,N_417,N_3809);
or U5174 (N_5174,N_4184,N_2847);
nor U5175 (N_5175,N_311,N_2812);
xor U5176 (N_5176,N_3446,N_2712);
and U5177 (N_5177,N_4953,N_3032);
nand U5178 (N_5178,N_3684,N_456);
and U5179 (N_5179,N_3461,N_3230);
nor U5180 (N_5180,N_2080,N_1611);
and U5181 (N_5181,N_854,N_119);
xnor U5182 (N_5182,N_1604,N_2214);
nand U5183 (N_5183,N_1497,N_1884);
nor U5184 (N_5184,N_2657,N_3804);
nand U5185 (N_5185,N_539,N_2223);
or U5186 (N_5186,N_1302,N_2774);
and U5187 (N_5187,N_69,N_1222);
nor U5188 (N_5188,N_1102,N_4027);
or U5189 (N_5189,N_1397,N_1643);
or U5190 (N_5190,N_1980,N_3788);
nor U5191 (N_5191,N_2785,N_256);
or U5192 (N_5192,N_505,N_1822);
or U5193 (N_5193,N_2532,N_1728);
or U5194 (N_5194,N_598,N_2108);
nor U5195 (N_5195,N_2287,N_1932);
nand U5196 (N_5196,N_4556,N_3448);
and U5197 (N_5197,N_3460,N_1419);
xnor U5198 (N_5198,N_3686,N_4598);
and U5199 (N_5199,N_827,N_3623);
nand U5200 (N_5200,N_4323,N_3727);
or U5201 (N_5201,N_1334,N_3228);
nand U5202 (N_5202,N_2813,N_819);
or U5203 (N_5203,N_719,N_1965);
nand U5204 (N_5204,N_1916,N_4438);
or U5205 (N_5205,N_1378,N_2015);
nand U5206 (N_5206,N_268,N_1590);
nand U5207 (N_5207,N_4996,N_1997);
and U5208 (N_5208,N_3085,N_4206);
or U5209 (N_5209,N_3102,N_4054);
xor U5210 (N_5210,N_3436,N_3848);
nand U5211 (N_5211,N_4573,N_4436);
nor U5212 (N_5212,N_1589,N_2357);
nand U5213 (N_5213,N_4004,N_2988);
xnor U5214 (N_5214,N_2683,N_4564);
nor U5215 (N_5215,N_32,N_4736);
or U5216 (N_5216,N_733,N_2610);
nor U5217 (N_5217,N_4478,N_932);
or U5218 (N_5218,N_4802,N_1934);
xor U5219 (N_5219,N_1583,N_3207);
and U5220 (N_5220,N_766,N_3721);
xnor U5221 (N_5221,N_670,N_4715);
xnor U5222 (N_5222,N_4216,N_1498);
xor U5223 (N_5223,N_3441,N_3041);
or U5224 (N_5224,N_1990,N_2091);
nand U5225 (N_5225,N_974,N_2565);
and U5226 (N_5226,N_2944,N_4220);
or U5227 (N_5227,N_1048,N_4845);
nor U5228 (N_5228,N_2472,N_4619);
nand U5229 (N_5229,N_3831,N_3291);
or U5230 (N_5230,N_1427,N_1591);
nand U5231 (N_5231,N_1114,N_474);
and U5232 (N_5232,N_1608,N_450);
xor U5233 (N_5233,N_4354,N_330);
and U5234 (N_5234,N_3312,N_3544);
and U5235 (N_5235,N_204,N_4711);
and U5236 (N_5236,N_1893,N_1768);
or U5237 (N_5237,N_202,N_2806);
and U5238 (N_5238,N_1204,N_4311);
or U5239 (N_5239,N_902,N_4259);
and U5240 (N_5240,N_99,N_136);
or U5241 (N_5241,N_2782,N_1058);
nand U5242 (N_5242,N_4207,N_4900);
and U5243 (N_5243,N_938,N_2345);
and U5244 (N_5244,N_2348,N_2632);
and U5245 (N_5245,N_3124,N_4062);
nor U5246 (N_5246,N_3470,N_3373);
nor U5247 (N_5247,N_4403,N_4511);
or U5248 (N_5248,N_4606,N_4199);
and U5249 (N_5249,N_872,N_2184);
or U5250 (N_5250,N_4187,N_2055);
and U5251 (N_5251,N_4169,N_874);
and U5252 (N_5252,N_4267,N_4437);
nor U5253 (N_5253,N_3249,N_896);
and U5254 (N_5254,N_1677,N_1653);
nand U5255 (N_5255,N_4235,N_3569);
and U5256 (N_5256,N_2097,N_4678);
nand U5257 (N_5257,N_4702,N_2373);
or U5258 (N_5258,N_2788,N_3430);
nor U5259 (N_5259,N_4792,N_170);
nor U5260 (N_5260,N_3642,N_4790);
or U5261 (N_5261,N_496,N_2766);
or U5262 (N_5262,N_712,N_2939);
nand U5263 (N_5263,N_2810,N_1244);
or U5264 (N_5264,N_880,N_4001);
nor U5265 (N_5265,N_1845,N_3216);
and U5266 (N_5266,N_4093,N_1015);
or U5267 (N_5267,N_3557,N_1407);
or U5268 (N_5268,N_1559,N_4322);
and U5269 (N_5269,N_3117,N_2648);
nor U5270 (N_5270,N_231,N_813);
or U5271 (N_5271,N_4258,N_2857);
and U5272 (N_5272,N_3887,N_2787);
nand U5273 (N_5273,N_2606,N_4347);
nor U5274 (N_5274,N_4411,N_924);
nand U5275 (N_5275,N_1007,N_2064);
xnor U5276 (N_5276,N_4363,N_3196);
nand U5277 (N_5277,N_3095,N_3636);
nor U5278 (N_5278,N_4964,N_3454);
or U5279 (N_5279,N_1730,N_3941);
or U5280 (N_5280,N_1176,N_4191);
nand U5281 (N_5281,N_21,N_300);
and U5282 (N_5282,N_3979,N_2587);
nand U5283 (N_5283,N_4423,N_2941);
and U5284 (N_5284,N_2797,N_3495);
nand U5285 (N_5285,N_718,N_3759);
nor U5286 (N_5286,N_526,N_4238);
and U5287 (N_5287,N_4105,N_2168);
nor U5288 (N_5288,N_2304,N_2370);
nor U5289 (N_5289,N_3586,N_948);
or U5290 (N_5290,N_4506,N_1137);
nand U5291 (N_5291,N_3064,N_2832);
nor U5292 (N_5292,N_4080,N_377);
nand U5293 (N_5293,N_3154,N_3106);
and U5294 (N_5294,N_1010,N_1734);
xnor U5295 (N_5295,N_911,N_1556);
nand U5296 (N_5296,N_3699,N_1018);
nor U5297 (N_5297,N_4889,N_1355);
and U5298 (N_5298,N_3731,N_1509);
nor U5299 (N_5299,N_2658,N_4464);
or U5300 (N_5300,N_1038,N_1518);
or U5301 (N_5301,N_1561,N_4410);
nand U5302 (N_5302,N_1852,N_3725);
nand U5303 (N_5303,N_4525,N_1760);
and U5304 (N_5304,N_1274,N_3997);
or U5305 (N_5305,N_4144,N_2756);
and U5306 (N_5306,N_1678,N_2169);
nor U5307 (N_5307,N_4659,N_2232);
and U5308 (N_5308,N_3224,N_2331);
and U5309 (N_5309,N_2501,N_3445);
or U5310 (N_5310,N_3932,N_3184);
nor U5311 (N_5311,N_4903,N_26);
nor U5312 (N_5312,N_869,N_4657);
xnor U5313 (N_5313,N_2896,N_4360);
or U5314 (N_5314,N_3015,N_2960);
nand U5315 (N_5315,N_3728,N_4721);
or U5316 (N_5316,N_1299,N_626);
and U5317 (N_5317,N_2354,N_4646);
or U5318 (N_5318,N_2196,N_838);
or U5319 (N_5319,N_3007,N_2305);
and U5320 (N_5320,N_3022,N_1679);
or U5321 (N_5321,N_1120,N_1710);
or U5322 (N_5322,N_4396,N_3859);
nand U5323 (N_5323,N_1720,N_1843);
nand U5324 (N_5324,N_3241,N_2961);
or U5325 (N_5325,N_3667,N_4502);
nor U5326 (N_5326,N_4116,N_841);
nand U5327 (N_5327,N_4457,N_3820);
and U5328 (N_5328,N_736,N_385);
and U5329 (N_5329,N_643,N_1903);
and U5330 (N_5330,N_3538,N_4233);
xor U5331 (N_5331,N_2966,N_950);
or U5332 (N_5332,N_3001,N_3084);
nor U5333 (N_5333,N_2667,N_4398);
or U5334 (N_5334,N_3339,N_1076);
or U5335 (N_5335,N_3695,N_116);
xor U5336 (N_5336,N_3428,N_4735);
xnor U5337 (N_5337,N_829,N_1316);
and U5338 (N_5338,N_816,N_2129);
and U5339 (N_5339,N_1784,N_2919);
and U5340 (N_5340,N_4050,N_4453);
nor U5341 (N_5341,N_407,N_3733);
xnor U5342 (N_5342,N_4078,N_3635);
nand U5343 (N_5343,N_2178,N_1895);
nor U5344 (N_5344,N_2863,N_1665);
or U5345 (N_5345,N_4250,N_4738);
nor U5346 (N_5346,N_4167,N_4387);
or U5347 (N_5347,N_4315,N_4645);
nor U5348 (N_5348,N_462,N_2146);
nand U5349 (N_5349,N_3622,N_1020);
or U5350 (N_5350,N_694,N_1309);
xnor U5351 (N_5351,N_4369,N_596);
nor U5352 (N_5352,N_4866,N_1464);
and U5353 (N_5353,N_4627,N_1063);
nand U5354 (N_5354,N_1229,N_4407);
and U5355 (N_5355,N_1578,N_963);
nor U5356 (N_5356,N_4641,N_3257);
and U5357 (N_5357,N_2871,N_1491);
and U5358 (N_5358,N_866,N_2350);
nand U5359 (N_5359,N_1131,N_1276);
and U5360 (N_5360,N_1291,N_1557);
or U5361 (N_5361,N_2808,N_1021);
nand U5362 (N_5362,N_4035,N_4538);
nor U5363 (N_5363,N_1178,N_1171);
nor U5364 (N_5364,N_4677,N_3414);
or U5365 (N_5365,N_4325,N_2319);
nand U5366 (N_5366,N_2407,N_361);
nor U5367 (N_5367,N_517,N_3045);
nor U5368 (N_5368,N_2881,N_3305);
xnor U5369 (N_5369,N_4230,N_2572);
and U5370 (N_5370,N_3043,N_2126);
and U5371 (N_5371,N_1826,N_1200);
nand U5372 (N_5372,N_3376,N_3130);
and U5373 (N_5373,N_3127,N_1800);
nor U5374 (N_5374,N_3128,N_446);
nand U5375 (N_5375,N_161,N_3899);
nand U5376 (N_5376,N_4512,N_4096);
or U5377 (N_5377,N_2526,N_916);
nand U5378 (N_5378,N_1109,N_4454);
and U5379 (N_5379,N_4772,N_1197);
and U5380 (N_5380,N_369,N_4079);
xor U5381 (N_5381,N_215,N_587);
or U5382 (N_5382,N_3583,N_2101);
xnor U5383 (N_5383,N_2041,N_4658);
nor U5384 (N_5384,N_793,N_1483);
nand U5385 (N_5385,N_128,N_2711);
nor U5386 (N_5386,N_2890,N_1953);
xnor U5387 (N_5387,N_3907,N_4368);
and U5388 (N_5388,N_3690,N_1233);
xor U5389 (N_5389,N_3256,N_1245);
nand U5390 (N_5390,N_3396,N_2674);
and U5391 (N_5391,N_3991,N_4585);
nand U5392 (N_5392,N_2784,N_3026);
nand U5393 (N_5393,N_3370,N_1575);
or U5394 (N_5394,N_4950,N_3808);
or U5395 (N_5395,N_1817,N_1874);
nor U5396 (N_5396,N_2404,N_803);
and U5397 (N_5397,N_4261,N_2490);
nand U5398 (N_5398,N_3529,N_4798);
or U5399 (N_5399,N_53,N_3222);
and U5400 (N_5400,N_4089,N_4388);
nand U5401 (N_5401,N_889,N_216);
nand U5402 (N_5402,N_3659,N_1855);
or U5403 (N_5403,N_3131,N_1538);
or U5404 (N_5404,N_1496,N_2705);
and U5405 (N_5405,N_673,N_3341);
or U5406 (N_5406,N_239,N_3774);
nand U5407 (N_5407,N_4265,N_3678);
nor U5408 (N_5408,N_2007,N_1991);
nand U5409 (N_5409,N_2545,N_3944);
nor U5410 (N_5410,N_524,N_509);
and U5411 (N_5411,N_137,N_2246);
nand U5412 (N_5412,N_4461,N_3218);
or U5413 (N_5413,N_4752,N_3136);
nor U5414 (N_5414,N_2173,N_2765);
xor U5415 (N_5415,N_2171,N_4956);
and U5416 (N_5416,N_3013,N_2737);
and U5417 (N_5417,N_2139,N_1467);
xnor U5418 (N_5418,N_4371,N_272);
xnor U5419 (N_5419,N_3992,N_632);
and U5420 (N_5420,N_223,N_2959);
and U5421 (N_5421,N_3650,N_3294);
xnor U5422 (N_5422,N_1902,N_281);
and U5423 (N_5423,N_1571,N_4320);
nor U5424 (N_5424,N_2625,N_2235);
and U5425 (N_5425,N_1090,N_1918);
nor U5426 (N_5426,N_2471,N_4375);
and U5427 (N_5427,N_2520,N_1599);
or U5428 (N_5428,N_453,N_2362);
or U5429 (N_5429,N_4800,N_1416);
nor U5430 (N_5430,N_3393,N_3679);
nor U5431 (N_5431,N_3913,N_730);
nand U5432 (N_5432,N_2145,N_3543);
or U5433 (N_5433,N_1465,N_1379);
and U5434 (N_5434,N_4056,N_2824);
or U5435 (N_5435,N_1196,N_4940);
xnor U5436 (N_5436,N_4516,N_2991);
nor U5437 (N_5437,N_994,N_112);
or U5438 (N_5438,N_391,N_1703);
nor U5439 (N_5439,N_993,N_4644);
nor U5440 (N_5440,N_1612,N_1527);
nor U5441 (N_5441,N_2853,N_3606);
and U5442 (N_5442,N_3665,N_394);
or U5443 (N_5443,N_3147,N_262);
or U5444 (N_5444,N_1181,N_2996);
nand U5445 (N_5445,N_3601,N_460);
nor U5446 (N_5446,N_2402,N_2174);
xnor U5447 (N_5447,N_115,N_3290);
or U5448 (N_5448,N_3498,N_3764);
or U5449 (N_5449,N_4890,N_2973);
and U5450 (N_5450,N_4673,N_4639);
nor U5451 (N_5451,N_1542,N_555);
nor U5452 (N_5452,N_3059,N_3740);
nor U5453 (N_5453,N_1146,N_1209);
nand U5454 (N_5454,N_2249,N_490);
nor U5455 (N_5455,N_721,N_3878);
nand U5456 (N_5456,N_381,N_138);
nand U5457 (N_5457,N_1238,N_3279);
nand U5458 (N_5458,N_1700,N_1016);
nor U5459 (N_5459,N_1144,N_3969);
and U5460 (N_5460,N_514,N_1969);
and U5461 (N_5461,N_4264,N_3476);
xor U5462 (N_5462,N_1383,N_1503);
nand U5463 (N_5463,N_2188,N_4819);
and U5464 (N_5464,N_95,N_2982);
nand U5465 (N_5465,N_897,N_1284);
nand U5466 (N_5466,N_4281,N_4651);
nand U5467 (N_5467,N_3359,N_3328);
nor U5468 (N_5468,N_3263,N_1634);
nor U5469 (N_5469,N_142,N_512);
nand U5470 (N_5470,N_2615,N_50);
and U5471 (N_5471,N_1415,N_2958);
nand U5472 (N_5472,N_3814,N_4620);
and U5473 (N_5473,N_2732,N_1096);
nand U5474 (N_5474,N_1025,N_3314);
and U5475 (N_5475,N_1567,N_4635);
xor U5476 (N_5476,N_2340,N_1977);
xor U5477 (N_5477,N_4352,N_4808);
or U5478 (N_5478,N_4888,N_498);
and U5479 (N_5479,N_421,N_1046);
and U5480 (N_5480,N_4134,N_2487);
nand U5481 (N_5481,N_912,N_4887);
and U5482 (N_5482,N_2928,N_2247);
and U5483 (N_5483,N_681,N_2314);
nand U5484 (N_5484,N_2075,N_3090);
xor U5485 (N_5485,N_3640,N_3912);
nand U5486 (N_5486,N_1788,N_4431);
and U5487 (N_5487,N_388,N_1227);
nor U5488 (N_5488,N_2533,N_2850);
xnor U5489 (N_5489,N_2742,N_3789);
nor U5490 (N_5490,N_1410,N_4365);
and U5491 (N_5491,N_4730,N_4085);
or U5492 (N_5492,N_171,N_292);
nand U5493 (N_5493,N_2855,N_3242);
nand U5494 (N_5494,N_3187,N_416);
nor U5495 (N_5495,N_4699,N_3431);
and U5496 (N_5496,N_3472,N_2470);
nand U5497 (N_5497,N_4070,N_560);
nand U5498 (N_5498,N_1733,N_1281);
and U5499 (N_5499,N_2926,N_265);
or U5500 (N_5500,N_2614,N_346);
nand U5501 (N_5501,N_483,N_3353);
and U5502 (N_5502,N_3687,N_1103);
nand U5503 (N_5503,N_1511,N_4013);
and U5504 (N_5504,N_4967,N_1252);
and U5505 (N_5505,N_1085,N_3922);
or U5506 (N_5506,N_858,N_1787);
xnor U5507 (N_5507,N_3151,N_1040);
xor U5508 (N_5508,N_4930,N_4928);
nor U5509 (N_5509,N_3828,N_3183);
nand U5510 (N_5510,N_4748,N_2187);
or U5511 (N_5511,N_104,N_1068);
nor U5512 (N_5512,N_2623,N_3491);
xor U5513 (N_5513,N_802,N_4024);
nor U5514 (N_5514,N_4954,N_2495);
nand U5515 (N_5515,N_700,N_1185);
xnor U5516 (N_5516,N_3463,N_691);
nand U5517 (N_5517,N_4146,N_879);
and U5518 (N_5518,N_2783,N_4504);
xnor U5519 (N_5519,N_37,N_4631);
xor U5520 (N_5520,N_1632,N_2444);
and U5521 (N_5521,N_779,N_4181);
nand U5522 (N_5522,N_3999,N_4270);
nand U5523 (N_5523,N_547,N_4210);
or U5524 (N_5524,N_1805,N_4708);
xor U5525 (N_5525,N_715,N_810);
nor U5526 (N_5526,N_4974,N_4192);
xor U5527 (N_5527,N_301,N_103);
nand U5528 (N_5528,N_3439,N_277);
and U5529 (N_5529,N_3852,N_4028);
and U5530 (N_5530,N_2210,N_2754);
or U5531 (N_5531,N_4066,N_2752);
nand U5532 (N_5532,N_2725,N_4117);
xor U5533 (N_5533,N_3115,N_4364);
and U5534 (N_5534,N_831,N_1619);
nor U5535 (N_5535,N_4650,N_293);
nand U5536 (N_5536,N_1246,N_3364);
and U5537 (N_5537,N_3046,N_2967);
xnor U5538 (N_5538,N_1210,N_457);
nor U5539 (N_5539,N_3258,N_3747);
and U5540 (N_5540,N_2775,N_2620);
or U5541 (N_5541,N_2036,N_3553);
or U5542 (N_5542,N_3404,N_1214);
or U5543 (N_5543,N_2128,N_72);
and U5544 (N_5544,N_1917,N_477);
xor U5545 (N_5545,N_93,N_3066);
and U5546 (N_5546,N_310,N_2248);
nor U5547 (N_5547,N_4959,N_4925);
nand U5548 (N_5548,N_2132,N_4562);
and U5549 (N_5549,N_4914,N_3772);
nand U5550 (N_5550,N_350,N_1240);
nor U5551 (N_5551,N_2138,N_353);
and U5552 (N_5552,N_1592,N_2087);
xor U5553 (N_5553,N_1566,N_3356);
and U5554 (N_5554,N_1620,N_1622);
xor U5555 (N_5555,N_354,N_2042);
or U5556 (N_5556,N_2956,N_3351);
xnor U5557 (N_5557,N_1369,N_4835);
nand U5558 (N_5558,N_1732,N_1709);
xor U5559 (N_5559,N_3818,N_3198);
and U5560 (N_5560,N_2460,N_3215);
nor U5561 (N_5561,N_2359,N_966);
nand U5562 (N_5562,N_760,N_4040);
nor U5563 (N_5563,N_4848,N_1774);
nor U5564 (N_5564,N_2258,N_3971);
and U5565 (N_5565,N_3327,N_4158);
nand U5566 (N_5566,N_557,N_1228);
nor U5567 (N_5567,N_352,N_3170);
and U5568 (N_5568,N_4613,N_882);
nand U5569 (N_5569,N_3611,N_10);
nand U5570 (N_5570,N_3607,N_1268);
nand U5571 (N_5571,N_2430,N_2978);
and U5572 (N_5572,N_1911,N_3137);
or U5573 (N_5573,N_1881,N_3802);
nor U5574 (N_5574,N_3579,N_3347);
nor U5575 (N_5575,N_1519,N_1073);
and U5576 (N_5576,N_411,N_120);
xnor U5577 (N_5577,N_45,N_2311);
nand U5578 (N_5578,N_2894,N_339);
nor U5579 (N_5579,N_1367,N_2523);
and U5580 (N_5580,N_4876,N_4787);
nand U5581 (N_5581,N_3896,N_3119);
nor U5582 (N_5582,N_4303,N_3452);
nand U5583 (N_5583,N_4878,N_3135);
and U5584 (N_5584,N_4321,N_3908);
or U5585 (N_5585,N_2994,N_4389);
or U5586 (N_5586,N_4841,N_3664);
nand U5587 (N_5587,N_2026,N_4472);
and U5588 (N_5588,N_4806,N_1502);
nor U5589 (N_5589,N_2159,N_1986);
nor U5590 (N_5590,N_4349,N_1071);
or U5591 (N_5591,N_3524,N_3838);
nor U5592 (N_5592,N_878,N_3420);
or U5593 (N_5593,N_825,N_3904);
nor U5594 (N_5594,N_1377,N_1646);
nand U5595 (N_5595,N_504,N_4186);
nor U5596 (N_5596,N_3400,N_1481);
nand U5597 (N_5597,N_1956,N_1972);
and U5598 (N_5598,N_419,N_373);
nand U5599 (N_5599,N_1866,N_536);
nand U5600 (N_5600,N_900,N_3781);
xnor U5601 (N_5601,N_611,N_4766);
and U5602 (N_5602,N_2493,N_2351);
or U5603 (N_5603,N_332,N_4530);
or U5604 (N_5604,N_723,N_2315);
nor U5605 (N_5605,N_2422,N_2024);
and U5606 (N_5606,N_3074,N_1809);
and U5607 (N_5607,N_2936,N_2029);
and U5608 (N_5608,N_507,N_4829);
and U5609 (N_5609,N_1512,N_606);
nor U5610 (N_5610,N_4307,N_4655);
nand U5611 (N_5611,N_111,N_342);
nand U5612 (N_5612,N_4276,N_2582);
and U5613 (N_5613,N_3743,N_2918);
nor U5614 (N_5614,N_3385,N_2274);
nor U5615 (N_5615,N_4409,N_33);
or U5616 (N_5616,N_2930,N_4190);
or U5617 (N_5617,N_3275,N_4667);
xnor U5618 (N_5618,N_4165,N_286);
and U5619 (N_5619,N_2089,N_2038);
and U5620 (N_5620,N_969,N_4185);
and U5621 (N_5621,N_3832,N_1594);
and U5622 (N_5622,N_619,N_3618);
and U5623 (N_5623,N_1231,N_1875);
and U5624 (N_5624,N_2047,N_3395);
or U5625 (N_5625,N_1263,N_4469);
nor U5626 (N_5626,N_4182,N_4960);
xnor U5627 (N_5627,N_2396,N_2751);
and U5628 (N_5628,N_1462,N_3845);
and U5629 (N_5629,N_1273,N_1782);
nand U5630 (N_5630,N_2937,N_4785);
or U5631 (N_5631,N_208,N_1028);
nor U5632 (N_5632,N_3036,N_2365);
xnor U5633 (N_5633,N_2183,N_2555);
or U5634 (N_5634,N_2035,N_1011);
or U5635 (N_5635,N_995,N_2332);
and U5636 (N_5636,N_3819,N_241);
nand U5637 (N_5637,N_2649,N_1487);
or U5638 (N_5638,N_1877,N_3739);
nand U5639 (N_5639,N_275,N_4160);
or U5640 (N_5640,N_3116,N_4640);
and U5641 (N_5641,N_436,N_3268);
nand U5642 (N_5642,N_338,N_2244);
nand U5643 (N_5643,N_964,N_122);
nor U5644 (N_5644,N_4778,N_4180);
nand U5645 (N_5645,N_3049,N_3317);
and U5646 (N_5646,N_3585,N_3011);
nand U5647 (N_5647,N_2250,N_915);
and U5648 (N_5648,N_3935,N_2778);
nand U5649 (N_5649,N_2288,N_3336);
nor U5650 (N_5650,N_4174,N_167);
nor U5651 (N_5651,N_3984,N_2330);
nor U5652 (N_5652,N_439,N_3703);
and U5653 (N_5653,N_1402,N_4832);
nand U5654 (N_5654,N_636,N_1208);
nor U5655 (N_5655,N_2229,N_3975);
nand U5656 (N_5656,N_4201,N_1104);
and U5657 (N_5657,N_55,N_3797);
nor U5658 (N_5658,N_42,N_317);
nand U5659 (N_5659,N_1645,N_4898);
nand U5660 (N_5660,N_3799,N_1009);
nor U5661 (N_5661,N_4414,N_3925);
and U5662 (N_5662,N_809,N_806);
and U5663 (N_5663,N_3039,N_2316);
or U5664 (N_5664,N_795,N_4723);
xnor U5665 (N_5665,N_988,N_2923);
xor U5666 (N_5666,N_3211,N_3326);
or U5667 (N_5667,N_2635,N_1535);
nand U5668 (N_5668,N_3722,N_383);
nand U5669 (N_5669,N_1674,N_1067);
xnor U5670 (N_5670,N_3697,N_219);
and U5671 (N_5671,N_4043,N_255);
and U5672 (N_5672,N_4611,N_3939);
nand U5673 (N_5673,N_4983,N_1588);
nor U5674 (N_5674,N_146,N_3536);
xor U5675 (N_5675,N_2764,N_3990);
or U5676 (N_5676,N_1999,N_4771);
nand U5677 (N_5677,N_630,N_1164);
xnor U5678 (N_5678,N_4329,N_572);
nor U5679 (N_5679,N_2140,N_3477);
nor U5680 (N_5680,N_2948,N_185);
nand U5681 (N_5681,N_2403,N_2356);
or U5682 (N_5682,N_1841,N_4045);
nand U5683 (N_5683,N_2612,N_4119);
nand U5684 (N_5684,N_4351,N_4840);
nand U5685 (N_5685,N_1952,N_4484);
nor U5686 (N_5686,N_895,N_1338);
nand U5687 (N_5687,N_2044,N_4107);
nor U5688 (N_5688,N_3274,N_4630);
nand U5689 (N_5689,N_959,N_3970);
or U5690 (N_5690,N_2728,N_3763);
and U5691 (N_5691,N_1905,N_2462);
and U5692 (N_5692,N_3429,N_550);
nor U5693 (N_5693,N_3709,N_3620);
nor U5694 (N_5694,N_663,N_3148);
or U5695 (N_5695,N_4698,N_973);
and U5696 (N_5696,N_2300,N_382);
nor U5697 (N_5697,N_862,N_181);
or U5698 (N_5698,N_2903,N_1345);
or U5699 (N_5699,N_3692,N_2056);
nand U5700 (N_5700,N_3019,N_2415);
and U5701 (N_5701,N_4548,N_234);
nor U5702 (N_5702,N_771,N_199);
or U5703 (N_5703,N_2999,N_1406);
or U5704 (N_5704,N_3514,N_3724);
nor U5705 (N_5705,N_818,N_1446);
nor U5706 (N_5706,N_1241,N_3178);
nand U5707 (N_5707,N_2155,N_3500);
nand U5708 (N_5708,N_3295,N_127);
xor U5709 (N_5709,N_4526,N_3633);
xnor U5710 (N_5710,N_4123,N_2580);
or U5711 (N_5711,N_4058,N_553);
nor U5712 (N_5712,N_367,N_2519);
nand U5713 (N_5713,N_2468,N_1955);
or U5714 (N_5714,N_1587,N_860);
nor U5715 (N_5715,N_1280,N_1339);
nand U5716 (N_5716,N_2588,N_3232);
and U5717 (N_5717,N_1318,N_1568);
nand U5718 (N_5718,N_1605,N_2448);
and U5719 (N_5719,N_3741,N_1865);
or U5720 (N_5720,N_289,N_1094);
nor U5721 (N_5721,N_489,N_565);
and U5722 (N_5722,N_1946,N_822);
nor U5723 (N_5723,N_3419,N_696);
or U5724 (N_5724,N_3929,N_3716);
nor U5725 (N_5725,N_3630,N_77);
nor U5726 (N_5726,N_1546,N_4087);
xor U5727 (N_5727,N_2616,N_4044);
nor U5728 (N_5728,N_145,N_684);
and U5729 (N_5729,N_3967,N_2800);
nand U5730 (N_5730,N_3158,N_3807);
nor U5731 (N_5731,N_4789,N_4282);
and U5732 (N_5732,N_2051,N_755);
nand U5733 (N_5733,N_3384,N_1161);
nand U5734 (N_5734,N_2142,N_1823);
and U5735 (N_5735,N_4716,N_1359);
nor U5736 (N_5736,N_196,N_1454);
nor U5737 (N_5737,N_513,N_358);
xor U5738 (N_5738,N_1032,N_4434);
nor U5739 (N_5739,N_3545,N_4125);
and U5740 (N_5740,N_2153,N_3021);
nor U5741 (N_5741,N_1942,N_2194);
xnor U5742 (N_5742,N_3843,N_4745);
and U5743 (N_5743,N_3185,N_1326);
nor U5744 (N_5744,N_1215,N_1167);
or U5745 (N_5745,N_562,N_1982);
or U5746 (N_5746,N_430,N_1656);
and U5747 (N_5747,N_4,N_843);
or U5748 (N_5748,N_4922,N_3647);
nor U5749 (N_5749,N_3316,N_2322);
xor U5750 (N_5750,N_2768,N_2296);
nor U5751 (N_5751,N_685,N_605);
and U5752 (N_5752,N_4850,N_2286);
and U5753 (N_5753,N_4683,N_3531);
and U5754 (N_5754,N_3286,N_658);
nor U5755 (N_5755,N_3854,N_2585);
or U5756 (N_5756,N_4337,N_4425);
or U5757 (N_5757,N_2477,N_4041);
and U5758 (N_5758,N_3837,N_3833);
and U5759 (N_5759,N_821,N_2164);
nor U5760 (N_5760,N_3040,N_4719);
nand U5761 (N_5761,N_1930,N_2445);
nand U5762 (N_5762,N_1501,N_772);
nor U5763 (N_5763,N_933,N_3765);
nor U5764 (N_5764,N_1565,N_4340);
nor U5765 (N_5765,N_1791,N_804);
or U5766 (N_5766,N_1835,N_1036);
and U5767 (N_5767,N_2436,N_998);
and U5768 (N_5768,N_2845,N_525);
nor U5769 (N_5769,N_2593,N_2355);
nor U5770 (N_5770,N_4704,N_218);
and U5771 (N_5771,N_4705,N_3700);
nor U5772 (N_5772,N_660,N_472);
or U5773 (N_5773,N_762,N_449);
or U5774 (N_5774,N_3950,N_2148);
nor U5775 (N_5775,N_4345,N_1931);
or U5776 (N_5776,N_1872,N_2701);
nand U5777 (N_5777,N_3450,N_3959);
nor U5778 (N_5778,N_4482,N_3502);
or U5779 (N_5779,N_1764,N_2020);
or U5780 (N_5780,N_1839,N_4072);
nor U5781 (N_5781,N_840,N_3005);
and U5782 (N_5782,N_438,N_4225);
nand U5783 (N_5783,N_2347,N_3881);
nor U5784 (N_5784,N_1601,N_4458);
nand U5785 (N_5785,N_333,N_2556);
nand U5786 (N_5786,N_4881,N_3815);
xnor U5787 (N_5787,N_4015,N_1148);
nor U5788 (N_5788,N_4034,N_3732);
nand U5789 (N_5789,N_156,N_835);
nor U5790 (N_5790,N_3693,N_3778);
or U5791 (N_5791,N_987,N_4463);
nand U5792 (N_5792,N_4196,N_2388);
xnor U5793 (N_5793,N_3836,N_2798);
and U5794 (N_5794,N_1133,N_2004);
or U5795 (N_5795,N_3417,N_1613);
or U5796 (N_5796,N_4251,N_1600);
and U5797 (N_5797,N_3978,N_4497);
nor U5798 (N_5798,N_422,N_2736);
or U5799 (N_5799,N_4594,N_1675);
nor U5800 (N_5800,N_2203,N_2391);
xnor U5801 (N_5801,N_3392,N_3259);
nor U5802 (N_5802,N_4252,N_1445);
nor U5803 (N_5803,N_3145,N_3631);
and U5804 (N_5804,N_1887,N_3399);
or U5805 (N_5805,N_397,N_1808);
or U5806 (N_5806,N_4933,N_746);
xor U5807 (N_5807,N_1737,N_2398);
xor U5808 (N_5808,N_3144,N_2935);
nor U5809 (N_5809,N_3480,N_1159);
nor U5810 (N_5810,N_4370,N_3829);
or U5811 (N_5811,N_4751,N_318);
nor U5812 (N_5812,N_1051,N_3683);
nand U5813 (N_5813,N_1745,N_3485);
nor U5814 (N_5814,N_390,N_1083);
and U5815 (N_5815,N_2335,N_759);
nor U5816 (N_5816,N_1069,N_502);
and U5817 (N_5817,N_4330,N_1414);
and U5818 (N_5818,N_522,N_1294);
xor U5819 (N_5819,N_2438,N_228);
xnor U5820 (N_5820,N_4031,N_3415);
xor U5821 (N_5821,N_4284,N_2878);
and U5822 (N_5822,N_4063,N_3598);
or U5823 (N_5823,N_4901,N_1234);
and U5824 (N_5824,N_4862,N_4255);
nor U5825 (N_5825,N_2828,N_1138);
nor U5826 (N_5826,N_545,N_1940);
nand U5827 (N_5827,N_402,N_2180);
nor U5828 (N_5828,N_3035,N_2691);
nand U5829 (N_5829,N_4624,N_4610);
nor U5830 (N_5830,N_92,N_3063);
nand U5831 (N_5831,N_1748,N_1350);
nor U5832 (N_5832,N_3118,N_767);
or U5833 (N_5833,N_4292,N_4399);
and U5834 (N_5834,N_3238,N_1433);
or U5835 (N_5835,N_1077,N_2189);
or U5836 (N_5836,N_599,N_2408);
nand U5837 (N_5837,N_71,N_892);
nor U5838 (N_5838,N_1998,N_4572);
and U5839 (N_5839,N_608,N_1458);
nor U5840 (N_5840,N_2897,N_716);
xnor U5841 (N_5841,N_325,N_266);
nor U5842 (N_5842,N_4874,N_1044);
or U5843 (N_5843,N_4777,N_4513);
or U5844 (N_5844,N_2929,N_2454);
nor U5845 (N_5845,N_2455,N_3200);
xor U5846 (N_5846,N_39,N_2427);
and U5847 (N_5847,N_3860,N_493);
xnor U5848 (N_5848,N_3467,N_3250);
xor U5849 (N_5849,N_1638,N_579);
nand U5850 (N_5850,N_727,N_4946);
nor U5851 (N_5851,N_2543,N_782);
or U5852 (N_5852,N_4492,N_616);
or U5853 (N_5853,N_985,N_4714);
nor U5854 (N_5854,N_2672,N_4025);
nor U5855 (N_5855,N_4958,N_1586);
or U5856 (N_5856,N_1471,N_1180);
nand U5857 (N_5857,N_13,N_4686);
and U5858 (N_5858,N_3020,N_2819);
nor U5859 (N_5859,N_4164,N_1042);
nand U5860 (N_5860,N_4090,N_3079);
or U5861 (N_5861,N_3672,N_227);
nand U5862 (N_5862,N_1562,N_2983);
or U5863 (N_5863,N_2360,N_1093);
or U5864 (N_5864,N_481,N_4285);
nor U5865 (N_5865,N_3194,N_713);
nor U5866 (N_5866,N_2513,N_3503);
nor U5867 (N_5867,N_1827,N_2830);
nand U5868 (N_5868,N_3745,N_3537);
and U5869 (N_5869,N_2423,N_4580);
nor U5870 (N_5870,N_4720,N_2114);
and U5871 (N_5871,N_2591,N_1658);
xor U5872 (N_5872,N_3546,N_3469);
nand U5873 (N_5873,N_4475,N_3752);
nand U5874 (N_5874,N_615,N_1898);
or U5875 (N_5875,N_4150,N_516);
nor U5876 (N_5876,N_1551,N_3552);
nand U5877 (N_5877,N_568,N_1676);
or U5878 (N_5878,N_765,N_4742);
nor U5879 (N_5879,N_4427,N_2979);
xor U5880 (N_5880,N_3776,N_921);
and U5881 (N_5881,N_515,N_488);
nor U5882 (N_5882,N_4549,N_741);
nor U5883 (N_5883,N_2746,N_800);
or U5884 (N_5884,N_501,N_2938);
nand U5885 (N_5885,N_61,N_4278);
nor U5886 (N_5886,N_601,N_3582);
and U5887 (N_5887,N_2854,N_1834);
xor U5888 (N_5888,N_3509,N_745);
xor U5889 (N_5889,N_3806,N_1248);
and U5890 (N_5890,N_965,N_1029);
and U5891 (N_5891,N_3239,N_2549);
and U5892 (N_5892,N_1603,N_250);
nor U5893 (N_5893,N_679,N_3270);
and U5894 (N_5894,N_217,N_1735);
nand U5895 (N_5895,N_4560,N_1370);
or U5896 (N_5896,N_4596,N_3749);
and U5897 (N_5897,N_1563,N_4688);
and U5898 (N_5898,N_3508,N_2856);
and U5899 (N_5899,N_80,N_2561);
and U5900 (N_5900,N_2410,N_3443);
nand U5901 (N_5901,N_628,N_177);
nand U5902 (N_5902,N_2285,N_1950);
xnor U5903 (N_5903,N_2862,N_1422);
or U5904 (N_5904,N_2213,N_304);
and U5905 (N_5905,N_3453,N_3352);
xor U5906 (N_5906,N_2916,N_589);
nor U5907 (N_5907,N_3173,N_1461);
nor U5908 (N_5908,N_4067,N_1668);
or U5909 (N_5909,N_3960,N_552);
and U5910 (N_5910,N_4680,N_538);
nand U5911 (N_5911,N_1721,N_4011);
nor U5912 (N_5912,N_4053,N_3974);
or U5913 (N_5913,N_2260,N_264);
nand U5914 (N_5914,N_1430,N_1290);
nor U5915 (N_5915,N_1024,N_2829);
nand U5916 (N_5916,N_3499,N_3987);
xnor U5917 (N_5917,N_783,N_3226);
or U5918 (N_5918,N_3576,N_1287);
nor U5919 (N_5919,N_3515,N_4938);
nor U5920 (N_5920,N_4851,N_2901);
or U5921 (N_5921,N_2718,N_4893);
or U5922 (N_5922,N_847,N_3645);
xor U5923 (N_5923,N_2776,N_4130);
nand U5924 (N_5924,N_3126,N_4854);
and U5925 (N_5925,N_815,N_1915);
or U5926 (N_5926,N_1913,N_243);
or U5927 (N_5927,N_4154,N_1293);
and U5928 (N_5928,N_2105,N_1026);
nor U5929 (N_5929,N_284,N_3367);
nor U5930 (N_5930,N_337,N_4534);
nand U5931 (N_5931,N_190,N_2478);
and U5932 (N_5932,N_3769,N_357);
and U5933 (N_5933,N_3530,N_3141);
and U5934 (N_5934,N_1780,N_1824);
or U5935 (N_5935,N_2900,N_4977);
or U5936 (N_5936,N_4533,N_1899);
nor U5937 (N_5937,N_2113,N_4763);
nor U5938 (N_5938,N_3231,N_4857);
nand U5939 (N_5939,N_4172,N_4194);
nand U5940 (N_5940,N_2738,N_970);
nor U5941 (N_5941,N_3323,N_3320);
or U5942 (N_5942,N_3738,N_3034);
xnor U5943 (N_5943,N_3089,N_343);
or U5944 (N_5944,N_374,N_537);
nor U5945 (N_5945,N_4214,N_2895);
nand U5946 (N_5946,N_2689,N_2483);
nor U5947 (N_5947,N_2722,N_478);
xor U5948 (N_5948,N_4661,N_861);
nor U5949 (N_5949,N_4666,N_984);
nor U5950 (N_5950,N_1775,N_4081);
and U5951 (N_5951,N_2714,N_1663);
and U5952 (N_5952,N_3670,N_4319);
nand U5953 (N_5953,N_1115,N_154);
nand U5954 (N_5954,N_3333,N_1070);
xor U5955 (N_5955,N_4426,N_3746);
nor U5956 (N_5956,N_492,N_2827);
nand U5957 (N_5957,N_4227,N_2094);
nor U5958 (N_5958,N_3780,N_2012);
and U5959 (N_5959,N_2517,N_2252);
nor U5960 (N_5960,N_2224,N_2974);
or U5961 (N_5961,N_1763,N_4612);
nor U5962 (N_5962,N_251,N_1373);
nand U5963 (N_5963,N_2602,N_257);
nor U5964 (N_5964,N_476,N_4676);
nand U5965 (N_5965,N_2222,N_4491);
nor U5966 (N_5966,N_3900,N_2611);
nand U5967 (N_5967,N_3426,N_2364);
nor U5968 (N_5968,N_4865,N_4827);
and U5969 (N_5969,N_3965,N_3785);
nand U5970 (N_5970,N_4653,N_1920);
nand U5971 (N_5971,N_4554,N_672);
nor U5972 (N_5972,N_4343,N_3835);
and U5973 (N_5973,N_2717,N_4769);
nand U5974 (N_5974,N_2310,N_1636);
xnor U5975 (N_5975,N_4249,N_4575);
nor U5976 (N_5976,N_2986,N_463);
and U5977 (N_5977,N_1499,N_937);
nor U5978 (N_5978,N_3931,N_4883);
and U5979 (N_5979,N_3047,N_1269);
and U5980 (N_5980,N_3111,N_3471);
xnor U5981 (N_5981,N_4886,N_4794);
and U5982 (N_5982,N_3104,N_1690);
and U5983 (N_5983,N_687,N_4725);
nand U5984 (N_5984,N_38,N_274);
nor U5985 (N_5985,N_2675,N_1205);
nor U5986 (N_5986,N_1948,N_4193);
or U5987 (N_5987,N_1975,N_4361);
nor U5988 (N_5988,N_2645,N_3157);
xor U5989 (N_5989,N_2157,N_1405);
or U5990 (N_5990,N_612,N_1968);
and U5991 (N_5991,N_711,N_4882);
xnor U5992 (N_5992,N_2050,N_954);
nor U5993 (N_5993,N_91,N_1797);
xor U5994 (N_5994,N_4217,N_4710);
nor U5995 (N_5995,N_1574,N_2685);
xnor U5996 (N_5996,N_3390,N_2706);
and U5997 (N_5997,N_209,N_2671);
nand U5998 (N_5998,N_3182,N_1279);
nand U5999 (N_5999,N_4843,N_341);
xor U6000 (N_6000,N_3600,N_1122);
nand U6001 (N_6001,N_2687,N_2710);
nor U6002 (N_6002,N_4138,N_425);
or U6003 (N_6003,N_1403,N_4703);
nand U6004 (N_6004,N_27,N_3101);
and U6005 (N_6005,N_646,N_2772);
nor U6006 (N_6006,N_4133,N_3521);
and U6007 (N_6007,N_2921,N_2104);
nor U6008 (N_6008,N_3541,N_4204);
nor U6009 (N_6009,N_1286,N_4254);
or U6010 (N_6010,N_3051,N_2665);
xor U6011 (N_6011,N_4801,N_1655);
xor U6012 (N_6012,N_2393,N_888);
nand U6013 (N_6013,N_3299,N_1545);
and U6014 (N_6014,N_2839,N_3943);
nor U6015 (N_6015,N_2381,N_2907);
and U6016 (N_6016,N_1879,N_4833);
nand U6017 (N_6017,N_1896,N_3217);
nor U6018 (N_6018,N_3570,N_3637);
nor U6019 (N_6019,N_4429,N_561);
or U6020 (N_6020,N_754,N_187);
nor U6021 (N_6021,N_909,N_3168);
xor U6022 (N_6022,N_418,N_1364);
nand U6023 (N_6023,N_3483,N_2272);
and U6024 (N_6024,N_3729,N_414);
and U6025 (N_6025,N_3786,N_2524);
nand U6026 (N_6026,N_152,N_4804);
and U6027 (N_6027,N_1798,N_3369);
nor U6028 (N_6028,N_639,N_1891);
or U6029 (N_6029,N_2419,N_4240);
or U6030 (N_6030,N_4121,N_1541);
nor U6031 (N_6031,N_320,N_2915);
or U6032 (N_6032,N_3338,N_3056);
nand U6033 (N_6033,N_4159,N_4218);
nand U6034 (N_6034,N_3590,N_885);
nand U6035 (N_6035,N_1084,N_2065);
nor U6036 (N_6036,N_2204,N_1387);
nand U6037 (N_6037,N_634,N_4260);
nor U6038 (N_6038,N_2418,N_3644);
nand U6039 (N_6039,N_4961,N_824);
or U6040 (N_6040,N_857,N_4795);
or U6041 (N_6041,N_661,N_4537);
nor U6042 (N_6042,N_287,N_2542);
and U6043 (N_6043,N_4510,N_4696);
nand U6044 (N_6044,N_139,N_4595);
xor U6045 (N_6045,N_2870,N_613);
xor U6046 (N_6046,N_64,N_1166);
nand U6047 (N_6047,N_952,N_468);
and U6048 (N_6048,N_3730,N_859);
nor U6049 (N_6049,N_1237,N_4039);
nor U6050 (N_6050,N_638,N_3889);
and U6051 (N_6051,N_3235,N_1981);
xor U6052 (N_6052,N_1212,N_1192);
nor U6053 (N_6053,N_3221,N_150);
xor U6054 (N_6054,N_4542,N_1194);
xor U6055 (N_6055,N_4445,N_530);
and U6056 (N_6056,N_364,N_2662);
and U6057 (N_6057,N_982,N_4687);
nor U6058 (N_6058,N_2071,N_2538);
or U6059 (N_6059,N_1941,N_2557);
or U6060 (N_6060,N_2200,N_426);
and U6061 (N_6061,N_2663,N_864);
nor U6062 (N_6062,N_2484,N_4951);
or U6063 (N_6063,N_1450,N_2177);
xnor U6064 (N_6064,N_1473,N_2626);
and U6065 (N_6065,N_518,N_81);
and U6066 (N_6066,N_1996,N_1987);
nand U6067 (N_6067,N_1516,N_1754);
or U6068 (N_6068,N_1816,N_708);
xnor U6069 (N_6069,N_4335,N_1844);
or U6070 (N_6070,N_1308,N_296);
nor U6071 (N_6071,N_3571,N_4729);
nand U6072 (N_6072,N_2209,N_4433);
xor U6073 (N_6073,N_2848,N_2045);
and U6074 (N_6074,N_4836,N_4183);
or U6075 (N_6075,N_3493,N_288);
nor U6076 (N_6076,N_2367,N_4505);
nor U6077 (N_6077,N_2241,N_2574);
or U6078 (N_6078,N_4591,N_1906);
nand U6079 (N_6079,N_979,N_3604);
or U6080 (N_6080,N_3562,N_3080);
and U6081 (N_6081,N_2864,N_4367);
or U6082 (N_6082,N_2589,N_3083);
and U6083 (N_6083,N_956,N_1199);
or U6084 (N_6084,N_3898,N_967);
nand U6085 (N_6085,N_4724,N_2368);
nor U6086 (N_6086,N_3186,N_76);
nor U6087 (N_6087,N_3099,N_655);
nand U6088 (N_6088,N_4170,N_3548);
nand U6089 (N_6089,N_1552,N_3464);
xor U6090 (N_6090,N_4980,N_4274);
or U6091 (N_6091,N_4202,N_4626);
and U6092 (N_6092,N_3773,N_1395);
and U6093 (N_6093,N_2034,N_2369);
and U6094 (N_6094,N_1544,N_253);
nor U6095 (N_6095,N_4740,N_4576);
nor U6096 (N_6096,N_1354,N_1521);
xor U6097 (N_6097,N_3966,N_66);
nor U6098 (N_6098,N_4880,N_3387);
nand U6099 (N_6099,N_3874,N_336);
and U6100 (N_6100,N_1087,N_3409);
or U6101 (N_6101,N_3624,N_2149);
nand U6102 (N_6102,N_2925,N_2320);
or U6103 (N_6103,N_4815,N_1747);
and U6104 (N_6104,N_4774,N_3977);
or U6105 (N_6105,N_3798,N_887);
xor U6106 (N_6106,N_913,N_523);
or U6107 (N_6107,N_781,N_1649);
or U6108 (N_6108,N_3161,N_4921);
nor U6109 (N_6109,N_2641,N_3886);
or U6110 (N_6110,N_2212,N_1842);
and U6111 (N_6111,N_852,N_1974);
nand U6112 (N_6112,N_4103,N_2578);
nand U6113 (N_6113,N_3757,N_836);
and U6114 (N_6114,N_1220,N_4291);
nor U6115 (N_6115,N_206,N_2181);
or U6116 (N_6116,N_3596,N_942);
and U6117 (N_6117,N_3482,N_4157);
nor U6118 (N_6118,N_2443,N_3734);
nand U6119 (N_6119,N_3662,N_4283);
nand U6120 (N_6120,N_2326,N_1796);
or U6121 (N_6121,N_4288,N_4242);
and U6122 (N_6122,N_1479,N_2057);
and U6123 (N_6123,N_4336,N_4467);
xor U6124 (N_6124,N_3070,N_380);
nor U6125 (N_6125,N_2753,N_2399);
or U6126 (N_6126,N_3010,N_3150);
xnor U6127 (N_6127,N_18,N_482);
nor U6128 (N_6128,N_4385,N_3923);
nor U6129 (N_6129,N_3914,N_570);
nor U6130 (N_6130,N_2660,N_4161);
nor U6131 (N_6131,N_4648,N_174);
nor U6132 (N_6132,N_4931,N_3213);
and U6133 (N_6133,N_1307,N_2280);
and U6134 (N_6134,N_2009,N_2409);
or U6135 (N_6135,N_197,N_686);
nor U6136 (N_6136,N_3071,N_3237);
nand U6137 (N_6137,N_975,N_1813);
nor U6138 (N_6138,N_1335,N_2048);
nand U6139 (N_6139,N_3418,N_1820);
nand U6140 (N_6140,N_114,N_3489);
and U6141 (N_6141,N_2498,N_2575);
and U6142 (N_6142,N_222,N_3199);
nand U6143 (N_6143,N_4047,N_2161);
or U6144 (N_6144,N_2124,N_2509);
xor U6145 (N_6145,N_1680,N_4757);
nand U6146 (N_6146,N_3917,N_3615);
nor U6147 (N_6147,N_4508,N_1871);
or U6148 (N_6148,N_2027,N_4128);
or U6149 (N_6149,N_4899,N_4713);
nand U6150 (N_6150,N_1292,N_1285);
and U6151 (N_6151,N_4366,N_1749);
or U6152 (N_6152,N_118,N_2461);
or U6153 (N_6153,N_3050,N_4558);
and U6154 (N_6154,N_4422,N_3689);
and U6155 (N_6155,N_4275,N_331);
xnor U6156 (N_6156,N_692,N_1086);
nand U6157 (N_6157,N_3949,N_3996);
xnor U6158 (N_6158,N_4818,N_2609);
nand U6159 (N_6159,N_1912,N_2003);
nor U6160 (N_6160,N_1298,N_1801);
nor U6161 (N_6161,N_875,N_2242);
nor U6162 (N_6162,N_3513,N_1943);
nand U6163 (N_6163,N_143,N_2451);
and U6164 (N_6164,N_1374,N_2053);
or U6165 (N_6165,N_953,N_3839);
nand U6166 (N_6166,N_4603,N_328);
or U6167 (N_6167,N_2818,N_1440);
or U6168 (N_6168,N_695,N_4987);
and U6169 (N_6169,N_1207,N_2503);
or U6170 (N_6170,N_2281,N_1659);
and U6171 (N_6171,N_2442,N_1111);
or U6172 (N_6172,N_3602,N_4498);
nand U6173 (N_6173,N_533,N_1828);
or U6174 (N_6174,N_117,N_1759);
and U6175 (N_6175,N_1947,N_3883);
nor U6176 (N_6176,N_3909,N_2627);
or U6177 (N_6177,N_4391,N_2851);
and U6178 (N_6178,N_2182,N_2755);
or U6179 (N_6179,N_1282,N_2724);
nand U6180 (N_6180,N_3948,N_1128);
nand U6181 (N_6181,N_4547,N_3750);
nor U6182 (N_6182,N_4483,N_2465);
nor U6183 (N_6183,N_675,N_2062);
and U6184 (N_6184,N_1304,N_648);
nor U6185 (N_6185,N_3527,N_3796);
nand U6186 (N_6186,N_1066,N_4139);
nand U6187 (N_6187,N_4277,N_484);
or U6188 (N_6188,N_4208,N_3708);
xnor U6189 (N_6189,N_1558,N_3272);
nor U6190 (N_6190,N_3937,N_3389);
xor U6191 (N_6191,N_3201,N_3533);
or U6192 (N_6192,N_1107,N_702);
nor U6193 (N_6193,N_662,N_2028);
xnor U6194 (N_6194,N_4153,N_2634);
or U6195 (N_6195,N_226,N_3132);
and U6196 (N_6196,N_4994,N_2425);
nor U6197 (N_6197,N_1596,N_1697);
xnor U6198 (N_6198,N_3073,N_4947);
xnor U6199 (N_6199,N_4982,N_4071);
nor U6200 (N_6200,N_3349,N_785);
nand U6201 (N_6201,N_680,N_3078);
and U6202 (N_6202,N_4535,N_2995);
nand U6203 (N_6203,N_1761,N_2965);
or U6204 (N_6204,N_3313,N_826);
nor U6205 (N_6205,N_1253,N_2815);
or U6206 (N_6206,N_2624,N_1012);
nor U6207 (N_6207,N_556,N_2777);
and U6208 (N_6208,N_3162,N_3953);
or U6209 (N_6209,N_500,N_2372);
nand U6210 (N_6210,N_1979,N_4177);
nand U6211 (N_6211,N_4448,N_2688);
and U6212 (N_6212,N_4141,N_1190);
or U6213 (N_6213,N_359,N_2117);
and U6214 (N_6214,N_245,N_3269);
xor U6215 (N_6215,N_2207,N_4571);
nand U6216 (N_6216,N_1560,N_4531);
nor U6217 (N_6217,N_2726,N_3176);
and U6218 (N_6218,N_3363,N_1129);
and U6219 (N_6219,N_1531,N_1513);
nand U6220 (N_6220,N_2265,N_1524);
or U6221 (N_6221,N_4224,N_4544);
or U6222 (N_6222,N_3956,N_188);
and U6223 (N_6223,N_4393,N_1065);
or U6224 (N_6224,N_1376,N_4809);
or U6225 (N_6225,N_1886,N_2293);
xnor U6226 (N_6226,N_4455,N_475);
nor U6227 (N_6227,N_886,N_345);
nand U6228 (N_6228,N_1954,N_2516);
nor U6229 (N_6229,N_2255,N_3895);
and U6230 (N_6230,N_1352,N_3713);
nor U6231 (N_6231,N_3646,N_928);
nor U6232 (N_6232,N_291,N_2277);
nand U6233 (N_6233,N_1030,N_3302);
nand U6234 (N_6234,N_1526,N_4605);
and U6235 (N_6235,N_4069,N_249);
and U6236 (N_6236,N_3412,N_1386);
nor U6237 (N_6237,N_4084,N_2748);
or U6238 (N_6238,N_2892,N_732);
and U6239 (N_6239,N_3264,N_4248);
nor U6240 (N_6240,N_133,N_3065);
nor U6241 (N_6241,N_4781,N_4003);
nor U6242 (N_6242,N_4166,N_2823);
xnor U6243 (N_6243,N_3189,N_2115);
nand U6244 (N_6244,N_3857,N_321);
nand U6245 (N_6245,N_2584,N_2866);
nand U6246 (N_6246,N_2417,N_1472);
nor U6247 (N_6247,N_2413,N_1297);
and U6248 (N_6248,N_2165,N_566);
nand U6249 (N_6249,N_2030,N_485);
or U6250 (N_6250,N_1110,N_1825);
nor U6251 (N_6251,N_4988,N_2761);
nand U6252 (N_6252,N_3629,N_465);
nor U6253 (N_6253,N_4018,N_2291);
and U6254 (N_6254,N_3180,N_1310);
nand U6255 (N_6255,N_4920,N_2522);
and U6256 (N_6256,N_1846,N_240);
xor U6257 (N_6257,N_4332,N_444);
or U6258 (N_6258,N_323,N_3890);
or U6259 (N_6259,N_1014,N_1255);
and U6260 (N_6260,N_1795,N_2284);
or U6261 (N_6261,N_2160,N_4846);
or U6262 (N_6262,N_34,N_3850);
or U6263 (N_6263,N_3777,N_2758);
and U6264 (N_6264,N_3287,N_4149);
nor U6265 (N_6265,N_1812,N_2317);
or U6266 (N_6266,N_4509,N_2859);
or U6267 (N_6267,N_4607,N_2891);
nand U6268 (N_6268,N_4652,N_4435);
and U6269 (N_6269,N_528,N_2872);
or U6270 (N_6270,N_3594,N_3782);
nor U6271 (N_6271,N_1776,N_4927);
nor U6272 (N_6272,N_4008,N_883);
or U6273 (N_6273,N_4014,N_3174);
nand U6274 (N_6274,N_3002,N_4059);
nand U6275 (N_6275,N_4590,N_4136);
nor U6276 (N_6276,N_1296,N_1360);
and U6277 (N_6277,N_3715,N_4487);
nor U6278 (N_6278,N_441,N_1958);
nor U6279 (N_6279,N_690,N_280);
nand U6280 (N_6280,N_2902,N_927);
nand U6281 (N_6281,N_2820,N_2202);
xnor U6282 (N_6282,N_3588,N_3980);
nor U6283 (N_6283,N_575,N_4998);
nand U6284 (N_6284,N_1236,N_2416);
and U6285 (N_6285,N_3243,N_1173);
or U6286 (N_6286,N_2677,N_1254);
and U6287 (N_6287,N_1049,N_2107);
xnor U6288 (N_6288,N_1022,N_302);
and U6289 (N_6289,N_3166,N_1325);
or U6290 (N_6290,N_3421,N_2912);
nand U6291 (N_6291,N_4446,N_4257);
or U6292 (N_6292,N_3870,N_4112);
or U6293 (N_6293,N_2840,N_2741);
or U6294 (N_6294,N_1349,N_571);
nand U6295 (N_6295,N_747,N_1100);
nand U6296 (N_6296,N_3487,N_58);
xnor U6297 (N_6297,N_4582,N_433);
nor U6298 (N_6298,N_582,N_1971);
and U6299 (N_6299,N_4091,N_2270);
nand U6300 (N_6300,N_1818,N_1162);
and U6301 (N_6301,N_3413,N_4418);
nor U6302 (N_6302,N_1195,N_2592);
xnor U6303 (N_6303,N_3267,N_108);
nand U6304 (N_6304,N_2826,N_1331);
nand U6305 (N_6305,N_2700,N_2577);
or U6306 (N_6306,N_4324,N_2014);
nand U6307 (N_6307,N_761,N_1259);
or U6308 (N_6308,N_4957,N_3163);
nand U6309 (N_6309,N_4152,N_1673);
nand U6310 (N_6310,N_4864,N_1919);
nand U6311 (N_6311,N_4515,N_212);
nand U6312 (N_6312,N_4342,N_1019);
nand U6313 (N_6313,N_4825,N_2514);
or U6314 (N_6314,N_1224,N_778);
nand U6315 (N_6315,N_940,N_3915);
or U6316 (N_6316,N_3244,N_4327);
and U6317 (N_6317,N_583,N_1389);
nor U6318 (N_6318,N_3869,N_720);
nand U6319 (N_6319,N_442,N_904);
or U6320 (N_6320,N_4828,N_437);
nand U6321 (N_6321,N_3575,N_4755);
xor U6322 (N_6322,N_922,N_3625);
nand U6323 (N_6323,N_4376,N_4115);
nand U6324 (N_6324,N_17,N_3179);
nand U6325 (N_6325,N_4807,N_997);
nor U6326 (N_6326,N_298,N_3304);
nor U6327 (N_6327,N_3626,N_4868);
or U6328 (N_6328,N_2670,N_2096);
nor U6329 (N_6329,N_4402,N_2032);
and U6330 (N_6330,N_3875,N_1964);
nand U6331 (N_6331,N_1380,N_2497);
nor U6332 (N_6332,N_2496,N_1625);
nand U6333 (N_6333,N_2521,N_3195);
or U6334 (N_6334,N_2205,N_1039);
nand U6335 (N_6335,N_1183,N_676);
or U6336 (N_6336,N_3840,N_3033);
nand U6337 (N_6337,N_4243,N_4118);
nand U6338 (N_6338,N_3888,N_424);
xor U6339 (N_6339,N_4494,N_3255);
nor U6340 (N_6340,N_3322,N_270);
xnor U6341 (N_6341,N_2299,N_3873);
nand U6342 (N_6342,N_2333,N_4306);
and U6343 (N_6343,N_2236,N_1347);
nor U6344 (N_6344,N_2704,N_1342);
and U6345 (N_6345,N_4289,N_845);
xor U6346 (N_6346,N_31,N_370);
nor U6347 (N_6347,N_768,N_780);
nand U6348 (N_6348,N_1850,N_3696);
and U6349 (N_6349,N_3748,N_4784);
xor U6350 (N_6350,N_876,N_3054);
nor U6351 (N_6351,N_1336,N_729);
and U6352 (N_6352,N_2763,N_4634);
nor U6353 (N_6353,N_396,N_1683);
nand U6354 (N_6354,N_543,N_3813);
xor U6355 (N_6355,N_4441,N_1688);
xor U6356 (N_6356,N_654,N_2757);
and U6357 (N_6357,N_1034,N_2429);
and U6358 (N_6358,N_2201,N_2170);
nand U6359 (N_6359,N_2380,N_548);
nand U6360 (N_6360,N_1510,N_4588);
and U6361 (N_6361,N_57,N_2199);
or U6362 (N_6362,N_2116,N_3849);
nor U6363 (N_6363,N_340,N_1731);
and U6364 (N_6364,N_1610,N_752);
nand U6365 (N_6365,N_4442,N_1267);
and U6366 (N_6366,N_1203,N_4709);
nand U6367 (N_6367,N_2786,N_2811);
nor U6368 (N_6368,N_4718,N_1616);
nor U6369 (N_6369,N_4462,N_3346);
and U6370 (N_6370,N_2655,N_1411);
or U6371 (N_6371,N_4762,N_2638);
xor U6372 (N_6372,N_1072,N_1408);
xnor U6373 (N_6373,N_2740,N_3879);
nor U6374 (N_6374,N_183,N_4593);
and U6375 (N_6375,N_992,N_2245);
or U6376 (N_6376,N_651,N_4913);
nand U6377 (N_6377,N_3565,N_4266);
xor U6378 (N_6378,N_906,N_2327);
and U6379 (N_6379,N_3076,N_823);
or U6380 (N_6380,N_2962,N_3817);
or U6381 (N_6381,N_4969,N_329);
nor U6382 (N_6382,N_4747,N_3842);
and U6383 (N_6383,N_3335,N_2702);
and U6384 (N_6384,N_1362,N_428);
and U6385 (N_6385,N_1744,N_4662);
or U6386 (N_6386,N_1723,N_1682);
or U6387 (N_6387,N_4129,N_2770);
or U6388 (N_6388,N_4831,N_4855);
nand U6389 (N_6389,N_4480,N_3675);
or U6390 (N_6390,N_671,N_401);
nor U6391 (N_6391,N_1385,N_2922);
nor U6392 (N_6392,N_657,N_1444);
nor U6393 (N_6393,N_3526,N_1361);
xnor U6394 (N_6394,N_3668,N_3053);
nor U6395 (N_6395,N_4468,N_1543);
nor U6396 (N_6396,N_2773,N_2301);
nand U6397 (N_6397,N_666,N_3129);
nor U6398 (N_6398,N_899,N_2642);
or U6399 (N_6399,N_4871,N_372);
nand U6400 (N_6400,N_2946,N_609);
nor U6401 (N_6401,N_4077,N_4761);
nand U6402 (N_6402,N_3027,N_3110);
nand U6403 (N_6403,N_189,N_376);
nor U6404 (N_6404,N_3325,N_3023);
nor U6405 (N_6405,N_3042,N_1789);
or U6406 (N_6406,N_757,N_207);
and U6407 (N_6407,N_2231,N_1186);
or U6408 (N_6408,N_4700,N_4100);
nand U6409 (N_6409,N_1201,N_2976);
nor U6410 (N_6410,N_920,N_4765);
or U6411 (N_6411,N_738,N_1779);
or U6412 (N_6412,N_348,N_2163);
and U6413 (N_6413,N_4952,N_4076);
and U6414 (N_6414,N_246,N_3726);
and U6415 (N_6415,N_811,N_4838);
nor U6416 (N_6416,N_2302,N_4649);
xnor U6417 (N_6417,N_1478,N_4955);
and U6418 (N_6418,N_164,N_3488);
nor U6419 (N_6419,N_1738,N_2220);
and U6420 (N_6420,N_2474,N_2066);
and U6421 (N_6421,N_4346,N_740);
nand U6422 (N_6422,N_404,N_1743);
and U6423 (N_6423,N_3539,N_1388);
nand U6424 (N_6424,N_180,N_2666);
or U6425 (N_6425,N_2491,N_2914);
and U6426 (N_6426,N_1452,N_3581);
or U6427 (N_6427,N_1717,N_23);
xor U6428 (N_6428,N_2822,N_1213);
or U6429 (N_6429,N_3474,N_4000);
or U6430 (N_6430,N_735,N_362);
nand U6431 (N_6431,N_4668,N_2841);
nor U6432 (N_6432,N_4110,N_2447);
nor U6433 (N_6433,N_3202,N_2537);
nand U6434 (N_6434,N_7,N_2111);
nand U6435 (N_6435,N_2162,N_3233);
and U6436 (N_6436,N_1081,N_4380);
or U6437 (N_6437,N_4456,N_2086);
and U6438 (N_6438,N_4706,N_2873);
xnor U6439 (N_6439,N_4579,N_0);
and U6440 (N_6440,N_1938,N_603);
and U6441 (N_6441,N_1413,N_4728);
and U6442 (N_6442,N_3052,N_917);
nand U6443 (N_6443,N_983,N_3800);
and U6444 (N_6444,N_3655,N_1966);
nand U6445 (N_6445,N_79,N_1685);
nor U6446 (N_6446,N_2068,N_1329);
or U6447 (N_6447,N_375,N_4768);
nor U6448 (N_6448,N_163,N_2464);
nor U6449 (N_6449,N_4753,N_2141);
nand U6450 (N_6450,N_4625,N_1878);
and U6451 (N_6451,N_448,N_384);
or U6452 (N_6452,N_4861,N_4328);
or U6453 (N_6453,N_67,N_3081);
nand U6454 (N_6454,N_2716,N_2336);
or U6455 (N_6455,N_3736,N_6);
xnor U6456 (N_6456,N_3862,N_3794);
and U6457 (N_6457,N_1687,N_3627);
or U6458 (N_6458,N_2268,N_3296);
and U6459 (N_6459,N_3707,N_326);
nand U6460 (N_6460,N_3379,N_2303);
nand U6461 (N_6461,N_4520,N_4583);
nor U6462 (N_6462,N_1614,N_812);
nor U6463 (N_6463,N_1607,N_1631);
or U6464 (N_6464,N_820,N_4397);
nor U6465 (N_6465,N_2981,N_2428);
nand U6466 (N_6466,N_3197,N_1438);
nand U6467 (N_6467,N_1261,N_3946);
nor U6468 (N_6468,N_4359,N_4142);
nor U6469 (N_6469,N_4219,N_2678);
nand U6470 (N_6470,N_580,N_4064);
and U6471 (N_6471,N_3599,N_4628);
nor U6472 (N_6472,N_4421,N_2283);
or U6473 (N_6473,N_2805,N_3830);
nor U6474 (N_6474,N_121,N_2618);
nor U6475 (N_6475,N_100,N_4290);
nor U6476 (N_6476,N_1951,N_3698);
and U6477 (N_6477,N_3551,N_3028);
xor U6478 (N_6478,N_1831,N_1704);
xnor U6479 (N_6479,N_1097,N_1319);
nand U6480 (N_6480,N_2987,N_2560);
nor U6481 (N_6481,N_563,N_1804);
nor U6482 (N_6482,N_1320,N_4143);
and U6483 (N_6483,N_2375,N_3149);
xnor U6484 (N_6484,N_313,N_3175);
nor U6485 (N_6485,N_192,N_4486);
and U6486 (N_6486,N_4156,N_4030);
and U6487 (N_6487,N_1225,N_2308);
or U6488 (N_6488,N_455,N_2566);
and U6489 (N_6489,N_3866,N_4555);
or U6490 (N_6490,N_891,N_2762);
or U6491 (N_6491,N_977,N_3768);
and U6492 (N_6492,N_4222,N_2102);
or U6493 (N_6493,N_503,N_1365);
nor U6494 (N_6494,N_3952,N_2809);
and U6495 (N_6495,N_4750,N_756);
or U6496 (N_6496,N_1275,N_2570);
and U6497 (N_6497,N_113,N_1671);
or U6498 (N_6498,N_2230,N_1876);
xnor U6499 (N_6499,N_4569,N_1477);
nor U6500 (N_6500,N_1451,N_2803);
or U6501 (N_6501,N_2767,N_3072);
nand U6502 (N_6502,N_4473,N_3504);
nor U6503 (N_6503,N_447,N_3613);
nand U6504 (N_6504,N_4443,N_2292);
or U6505 (N_6505,N_56,N_2318);
and U6506 (N_6506,N_4023,N_144);
nor U6507 (N_6507,N_3989,N_2506);
xnor U6508 (N_6508,N_1289,N_1936);
and U6509 (N_6509,N_2861,N_3004);
nand U6510 (N_6510,N_4803,N_647);
and U6511 (N_6511,N_3669,N_1540);
nor U6512 (N_6512,N_763,N_4853);
nand U6513 (N_6513,N_1448,N_4780);
or U6514 (N_6514,N_4333,N_2790);
and U6515 (N_6515,N_2597,N_4449);
and U6516 (N_6516,N_2825,N_2595);
nor U6517 (N_6517,N_586,N_4088);
nor U6518 (N_6518,N_737,N_4452);
and U6519 (N_6519,N_3337,N_2219);
nor U6520 (N_6520,N_3641,N_1396);
or U6521 (N_6521,N_1001,N_3167);
xor U6522 (N_6522,N_4638,N_3910);
and U6523 (N_6523,N_1095,N_3891);
nand U6524 (N_6524,N_3397,N_3240);
and U6525 (N_6525,N_2860,N_1707);
xor U6526 (N_6526,N_2573,N_4155);
and U6527 (N_6527,N_2807,N_3884);
or U6528 (N_6528,N_4212,N_1484);
or U6529 (N_6529,N_3205,N_4178);
nand U6530 (N_6530,N_1434,N_4859);
xor U6531 (N_6531,N_3386,N_3466);
or U6532 (N_6532,N_2505,N_4521);
or U6533 (N_6533,N_1157,N_1644);
and U6534 (N_6534,N_132,N_4012);
or U6535 (N_6535,N_945,N_946);
nor U6536 (N_6536,N_3191,N_4726);
or U6537 (N_6537,N_4094,N_4221);
or U6538 (N_6538,N_4296,N_1833);
nand U6539 (N_6539,N_3125,N_4507);
nor U6540 (N_6540,N_9,N_2176);
nor U6541 (N_6541,N_4493,N_184);
or U6542 (N_6542,N_1832,N_1486);
and U6543 (N_6543,N_2021,N_3735);
nand U6544 (N_6544,N_3146,N_3973);
and U6545 (N_6545,N_2313,N_2637);
and U6546 (N_6546,N_4856,N_4300);
nor U6547 (N_6547,N_3398,N_2276);
nand U6548 (N_6548,N_4392,N_4756);
or U6549 (N_6549,N_1507,N_907);
nand U6550 (N_6550,N_3801,N_83);
or U6551 (N_6551,N_4406,N_3954);
nor U6552 (N_6552,N_2221,N_1856);
and U6553 (N_6553,N_855,N_29);
and U6554 (N_6554,N_968,N_2640);
or U6555 (N_6555,N_1741,N_1053);
or U6556 (N_6556,N_487,N_305);
nor U6557 (N_6557,N_728,N_3927);
and U6558 (N_6558,N_4813,N_1970);
nand U6559 (N_6559,N_2290,N_269);
or U6560 (N_6560,N_551,N_4200);
nor U6561 (N_6561,N_4949,N_2143);
or U6562 (N_6562,N_2100,N_4232);
and U6563 (N_6563,N_2801,N_4295);
nand U6564 (N_6564,N_4083,N_2218);
nor U6565 (N_6565,N_939,N_299);
and U6566 (N_6566,N_1528,N_3382);
nor U6567 (N_6567,N_1223,N_2366);
nand U6568 (N_6568,N_506,N_629);
or U6569 (N_6569,N_4892,N_4009);
nor U6570 (N_6570,N_4314,N_3486);
nand U6571 (N_6571,N_3853,N_4665);
xnor U6572 (N_6572,N_1306,N_2271);
or U6573 (N_6573,N_125,N_2942);
nand U6574 (N_6574,N_2099,N_4362);
xor U6575 (N_6575,N_3936,N_3587);
or U6576 (N_6576,N_4858,N_3771);
xor U6577 (N_6577,N_1727,N_59);
nor U6578 (N_6578,N_1907,N_4424);
and U6579 (N_6579,N_3082,N_918);
and U6580 (N_6580,N_4592,N_617);
nor U6581 (N_6581,N_4584,N_2877);
nor U6582 (N_6582,N_2729,N_2289);
nor U6583 (N_6583,N_389,N_2379);
nand U6584 (N_6584,N_2975,N_3926);
nor U6585 (N_6585,N_1520,N_157);
and U6586 (N_6586,N_4741,N_656);
nand U6587 (N_6587,N_1921,N_4586);
and U6588 (N_6588,N_3663,N_307);
nand U6589 (N_6589,N_4500,N_4872);
nand U6590 (N_6590,N_4189,N_1043);
or U6591 (N_6591,N_1505,N_294);
or U6592 (N_6592,N_1959,N_2817);
or U6593 (N_6593,N_4986,N_1184);
and U6594 (N_6594,N_1149,N_3278);
nor U6595 (N_6595,N_4744,N_3578);
nor U6596 (N_6596,N_588,N_2680);
nor U6597 (N_6597,N_1617,N_1894);
xnor U6598 (N_6598,N_2563,N_355);
and U6599 (N_6599,N_258,N_1150);
or U6600 (N_6600,N_881,N_594);
nand U6601 (N_6601,N_4020,N_722);
nor U6602 (N_6602,N_4919,N_445);
or U6603 (N_6603,N_4989,N_1962);
and U6604 (N_6604,N_1988,N_3651);
nand U6605 (N_6605,N_434,N_3123);
nor U6606 (N_6606,N_1577,N_2109);
nor U6607 (N_6607,N_387,N_4943);
nand U6608 (N_6608,N_3589,N_532);
and U6609 (N_6609,N_4518,N_1108);
nor U6610 (N_6610,N_1757,N_4005);
nor U6611 (N_6611,N_1327,N_3203);
and U6612 (N_6612,N_2439,N_3319);
nor U6613 (N_6613,N_542,N_4057);
and U6614 (N_6614,N_650,N_2651);
nor U6615 (N_6615,N_3266,N_943);
nor U6616 (N_6616,N_3284,N_4126);
or U6617 (N_6617,N_870,N_4948);
xnor U6618 (N_6618,N_3962,N_4495);
nor U6619 (N_6619,N_4415,N_2233);
and U6620 (N_6620,N_499,N_1699);
and U6621 (N_6621,N_1399,N_3229);
nand U6622 (N_6622,N_753,N_2337);
and U6623 (N_6623,N_3595,N_1547);
nand U6624 (N_6624,N_2993,N_1815);
and U6625 (N_6625,N_830,N_2604);
and U6626 (N_6626,N_3134,N_3751);
or U6627 (N_6627,N_1888,N_2453);
and U6628 (N_6628,N_2266,N_3787);
or U6629 (N_6629,N_4812,N_4937);
or U6630 (N_6630,N_976,N_3855);
xor U6631 (N_6631,N_3093,N_4412);
or U6632 (N_6632,N_3657,N_1191);
nand U6633 (N_6633,N_2515,N_242);
nand U6634 (N_6634,N_4674,N_3300);
nor U6635 (N_6635,N_842,N_3408);
nand U6636 (N_6636,N_3402,N_379);
xnor U6637 (N_6637,N_3988,N_271);
nand U6638 (N_6638,N_1074,N_2342);
or U6639 (N_6639,N_4891,N_578);
and U6640 (N_6640,N_2559,N_2392);
xnor U6641 (N_6641,N_295,N_3762);
nor U6642 (N_6642,N_4934,N_2424);
or U6643 (N_6643,N_1642,N_2135);
or U6644 (N_6644,N_1532,N_3009);
and U6645 (N_6645,N_4450,N_4966);
xnor U6646 (N_6646,N_3087,N_4692);
nor U6647 (N_6647,N_3682,N_4654);
and U6648 (N_6648,N_2259,N_770);
nor U6649 (N_6649,N_1525,N_4113);
and U6650 (N_6650,N_3029,N_1099);
and U6651 (N_6651,N_1793,N_283);
nand U6652 (N_6652,N_3603,N_3516);
and U6653 (N_6653,N_3556,N_519);
nor U6654 (N_6654,N_2719,N_2836);
or U6655 (N_6655,N_3000,N_2985);
xnor U6656 (N_6656,N_4973,N_1106);
xor U6657 (N_6657,N_2598,N_743);
and U6658 (N_6658,N_1689,N_94);
nand U6659 (N_6659,N_1156,N_4021);
xnor U6660 (N_6660,N_3181,N_2262);
xor U6661 (N_6661,N_3983,N_4637);
nand U6662 (N_6662,N_1265,N_1549);
nor U6663 (N_6663,N_3204,N_2092);
nand U6664 (N_6664,N_1455,N_999);
nor U6665 (N_6665,N_3342,N_2426);
nand U6666 (N_6666,N_459,N_2739);
or U6667 (N_6667,N_3871,N_4567);
nand U6668 (N_6668,N_3375,N_4546);
nand U6669 (N_6669,N_989,N_1459);
xnor U6670 (N_6670,N_4578,N_546);
nor U6671 (N_6671,N_2927,N_1686);
and U6672 (N_6672,N_1924,N_259);
or U6673 (N_6673,N_3245,N_2294);
nor U6674 (N_6674,N_2972,N_4241);
nand U6675 (N_6675,N_4877,N_3220);
and U6676 (N_6676,N_3666,N_4029);
and U6677 (N_6677,N_3018,N_4145);
nand U6678 (N_6678,N_1790,N_4060);
nand U6679 (N_6679,N_4656,N_3311);
nor U6680 (N_6680,N_4975,N_14);
and U6681 (N_6681,N_1400,N_3206);
and U6682 (N_6682,N_4759,N_4907);
xor U6683 (N_6683,N_2743,N_3770);
and U6684 (N_6684,N_4566,N_3535);
and U6685 (N_6685,N_1088,N_4101);
xor U6686 (N_6686,N_178,N_2695);
or U6687 (N_6687,N_2329,N_3865);
nor U6688 (N_6688,N_4075,N_2088);
xor U6689 (N_6689,N_1392,N_600);
nor U6690 (N_6690,N_4529,N_36);
xnor U6691 (N_6691,N_559,N_2383);
and U6692 (N_6692,N_1366,N_2376);
nor U6693 (N_6693,N_4669,N_3484);
or U6694 (N_6694,N_642,N_1117);
or U6695 (N_6695,N_3406,N_2799);
and U6696 (N_6696,N_2554,N_2309);
or U6697 (N_6697,N_4239,N_4682);
nor U6698 (N_6698,N_1949,N_1147);
and U6699 (N_6699,N_703,N_3465);
nand U6700 (N_6700,N_4690,N_1811);
nor U6701 (N_6701,N_335,N_4962);
and U6702 (N_6702,N_126,N_210);
nand U6703 (N_6703,N_535,N_1508);
and U6704 (N_6704,N_4474,N_1777);
nand U6705 (N_6705,N_2581,N_2893);
or U6706 (N_6706,N_3928,N_2040);
xnor U6707 (N_6707,N_2440,N_2552);
xnor U6708 (N_6708,N_901,N_244);
or U6709 (N_6709,N_2562,N_4885);
nor U6710 (N_6710,N_3451,N_260);
and U6711 (N_6711,N_3109,N_4379);
and U6712 (N_6712,N_1944,N_1662);
and U6713 (N_6713,N_3378,N_1762);
or U6714 (N_6714,N_87,N_4223);
and U6715 (N_6715,N_3994,N_4816);
nor U6716 (N_6716,N_4382,N_3344);
or U6717 (N_6717,N_919,N_2630);
or U6718 (N_6718,N_2307,N_2390);
nor U6719 (N_6719,N_267,N_3661);
nand U6720 (N_6720,N_4055,N_3810);
and U6721 (N_6721,N_1880,N_4305);
nor U6722 (N_6722,N_2507,N_1713);
xor U6723 (N_6723,N_2953,N_934);
or U6724 (N_6724,N_4010,N_16);
and U6725 (N_6725,N_1581,N_1136);
xor U6726 (N_6726,N_1555,N_2387);
nor U6727 (N_6727,N_4731,N_4451);
nand U6728 (N_6728,N_1767,N_3964);
nand U6729 (N_6729,N_4065,N_769);
nor U6730 (N_6730,N_3685,N_1593);
nor U6731 (N_6731,N_1323,N_1739);
nor U6732 (N_6732,N_1041,N_3025);
and U6733 (N_6733,N_4847,N_273);
or U6734 (N_6734,N_4979,N_4908);
and U6735 (N_6735,N_2793,N_3058);
and U6736 (N_6736,N_3405,N_1423);
or U6737 (N_6737,N_1926,N_2708);
and U6738 (N_6738,N_3930,N_4684);
or U6739 (N_6739,N_1494,N_1078);
and U6740 (N_6740,N_4664,N_1177);
nor U6741 (N_6741,N_2463,N_2208);
and U6742 (N_6742,N_1340,N_4430);
nor U6743 (N_6743,N_2843,N_201);
or U6744 (N_6744,N_2571,N_2964);
nand U6745 (N_6745,N_1669,N_930);
or U6746 (N_6746,N_1217,N_403);
nand U6747 (N_6747,N_4823,N_3614);
nand U6748 (N_6748,N_644,N_2492);
nor U6749 (N_6749,N_4488,N_3851);
and U6750 (N_6750,N_4577,N_3060);
nor U6751 (N_6751,N_3767,N_1978);
and U6752 (N_6752,N_3826,N_3945);
nor U6753 (N_6753,N_3942,N_3048);
nor U6754 (N_6754,N_2257,N_2273);
or U6755 (N_6755,N_2920,N_4600);
or U6756 (N_6756,N_4310,N_3456);
nor U6757 (N_6757,N_4179,N_701);
nor U6758 (N_6758,N_1211,N_4019);
nor U6759 (N_6759,N_3283,N_3712);
nor U6760 (N_6760,N_1624,N_4609);
or U6761 (N_6761,N_2156,N_344);
nor U6762 (N_6762,N_4824,N_1193);
and U6763 (N_6763,N_4317,N_3841);
xor U6764 (N_6764,N_618,N_649);
and U6765 (N_6765,N_2074,N_1321);
nand U6766 (N_6766,N_2228,N_3691);
and U6767 (N_6767,N_4568,N_1537);
or U6768 (N_6768,N_2690,N_440);
and U6769 (N_6769,N_2734,N_1490);
or U6770 (N_6770,N_2594,N_773);
nor U6771 (N_6771,N_3343,N_1837);
or U6772 (N_6772,N_2852,N_4262);
nor U6773 (N_6773,N_1127,N_2512);
nor U6774 (N_6774,N_4476,N_4465);
nor U6775 (N_6775,N_2699,N_2267);
nor U6776 (N_6776,N_3827,N_3501);
nor U6777 (N_6777,N_3957,N_1691);
nor U6778 (N_6778,N_1585,N_3139);
nor U6779 (N_6779,N_194,N_1529);
xor U6780 (N_6780,N_1412,N_4294);
nor U6781 (N_6781,N_4541,N_497);
and U6782 (N_6782,N_2186,N_3742);
or U6783 (N_6783,N_1187,N_2043);
nor U6784 (N_6784,N_4782,N_1428);
nor U6785 (N_6785,N_4902,N_2473);
and U6786 (N_6786,N_3265,N_3561);
and U6787 (N_6787,N_3251,N_3014);
and U6788 (N_6788,N_1929,N_4002);
nand U6789 (N_6789,N_4237,N_877);
or U6790 (N_6790,N_3652,N_1836);
nor U6791 (N_6791,N_1892,N_2833);
or U6792 (N_6792,N_491,N_4162);
nor U6793 (N_6793,N_2954,N_2529);
nand U6794 (N_6794,N_2061,N_2643);
and U6795 (N_6795,N_4811,N_3940);
nand U6796 (N_6796,N_3449,N_4271);
nor U6797 (N_6797,N_2621,N_1718);
or U6798 (N_6798,N_2945,N_2459);
and U6799 (N_6799,N_2405,N_3433);
or U6800 (N_6800,N_1332,N_4860);
nor U6801 (N_6801,N_1867,N_4875);
nand U6802 (N_6802,N_1488,N_683);
or U6803 (N_6803,N_668,N_4140);
nor U6804 (N_6804,N_1736,N_4915);
nor U6805 (N_6805,N_22,N_3100);
and U6806 (N_6806,N_1553,N_972);
and U6807 (N_6807,N_2849,N_4642);
or U6808 (N_6808,N_85,N_1132);
or U6809 (N_6809,N_3038,N_2749);
nor U6810 (N_6810,N_3882,N_2070);
and U6811 (N_6811,N_2789,N_1995);
nor U6812 (N_6812,N_4395,N_1101);
nor U6813 (N_6813,N_848,N_2617);
or U6814 (N_6814,N_3494,N_2613);
and U6815 (N_6815,N_2095,N_4440);
xnor U6816 (N_6816,N_3234,N_2150);
xnor U6817 (N_6817,N_2206,N_1356);
or U6818 (N_6818,N_1708,N_158);
and U6819 (N_6819,N_1814,N_4022);
xor U6820 (N_6820,N_1633,N_2197);
or U6821 (N_6821,N_3694,N_1344);
and U6822 (N_6822,N_3673,N_4821);
or U6823 (N_6823,N_3511,N_467);
nand U6824 (N_6824,N_717,N_3863);
nand U6825 (N_6825,N_3329,N_2835);
nand U6826 (N_6826,N_2816,N_2433);
and U6827 (N_6827,N_1705,N_724);
and U6828 (N_6828,N_610,N_1670);
nor U6829 (N_6829,N_4727,N_1062);
xnor U6830 (N_6830,N_585,N_3717);
nor U6831 (N_6831,N_5,N_4198);
nor U6832 (N_6832,N_3067,N_1165);
and U6833 (N_6833,N_363,N_63);
and U6834 (N_6834,N_4244,N_3008);
or U6835 (N_6835,N_1092,N_3605);
xnor U6836 (N_6836,N_3246,N_3961);
nor U6837 (N_6837,N_1140,N_229);
nand U6838 (N_6838,N_1134,N_890);
or U6839 (N_6839,N_1751,N_4417);
nor U6840 (N_6840,N_764,N_2601);
and U6841 (N_6841,N_3377,N_4197);
or U6842 (N_6842,N_3152,N_2951);
nand U6843 (N_6843,N_2254,N_2353);
nand U6844 (N_6844,N_3214,N_1116);
nand U6845 (N_6845,N_748,N_89);
nand U6846 (N_6846,N_3261,N_2017);
nand U6847 (N_6847,N_4339,N_1424);
and U6848 (N_6848,N_4033,N_787);
nand U6849 (N_6849,N_3097,N_4496);
or U6850 (N_6850,N_4570,N_1554);
or U6851 (N_6851,N_2457,N_3756);
or U6852 (N_6852,N_2485,N_285);
nor U6853 (N_6853,N_1006,N_4309);
or U6854 (N_6854,N_2771,N_4622);
and U6855 (N_6855,N_3133,N_3823);
xor U6856 (N_6856,N_3459,N_3307);
nor U6857 (N_6857,N_469,N_4978);
nor U6858 (N_6858,N_1515,N_3610);
nor U6859 (N_6859,N_1243,N_581);
and U6860 (N_6860,N_1052,N_2709);
nand U6861 (N_6861,N_1993,N_1056);
xnor U6862 (N_6862,N_834,N_60);
nand U6863 (N_6863,N_4318,N_1476);
and U6864 (N_6864,N_2106,N_1756);
or U6865 (N_6865,N_955,N_2631);
or U6866 (N_6866,N_4519,N_853);
nor U6867 (N_6867,N_3918,N_665);
xor U6868 (N_6868,N_1810,N_12);
and U6869 (N_6869,N_235,N_429);
nor U6870 (N_6870,N_166,N_65);
xor U6871 (N_6871,N_1300,N_1266);
nor U6872 (N_6872,N_2499,N_4820);
or U6873 (N_6873,N_4992,N_2838);
nor U6874 (N_6874,N_3057,N_1860);
nor U6875 (N_6875,N_1315,N_1000);
nor U6876 (N_6876,N_1247,N_3982);
nand U6877 (N_6877,N_3919,N_4514);
and U6878 (N_6878,N_3506,N_3030);
xor U6879 (N_6879,N_395,N_3981);
nor U6880 (N_6880,N_3972,N_3775);
and U6881 (N_6881,N_1050,N_214);
nand U6882 (N_6882,N_3916,N_2282);
nor U6883 (N_6883,N_2673,N_4381);
nor U6884 (N_6884,N_2654,N_2858);
nor U6885 (N_6885,N_2119,N_1657);
or U6886 (N_6886,N_134,N_1456);
or U6887 (N_6887,N_2727,N_4432);
nor U6888 (N_6888,N_3171,N_3822);
or U6889 (N_6889,N_4793,N_2731);
or U6890 (N_6890,N_4485,N_2016);
xor U6891 (N_6891,N_2653,N_4557);
nand U6892 (N_6892,N_3055,N_4471);
and U6893 (N_6893,N_1696,N_1372);
or U6894 (N_6894,N_3591,N_2669);
or U6895 (N_6895,N_3103,N_2191);
xnor U6896 (N_6896,N_849,N_1418);
or U6897 (N_6897,N_786,N_4981);
nand U6898 (N_6898,N_1057,N_98);
nor U6899 (N_6899,N_3877,N_3208);
nand U6900 (N_6900,N_3677,N_4895);
nand U6901 (N_6901,N_2374,N_386);
nor U6902 (N_6902,N_3612,N_2489);
nor U6903 (N_6903,N_3512,N_2759);
nor U6904 (N_6904,N_1047,N_2579);
nor U6905 (N_6905,N_1470,N_2217);
xor U6906 (N_6906,N_1849,N_1384);
or U6907 (N_6907,N_4439,N_129);
nand U6908 (N_6908,N_46,N_4770);
nor U6909 (N_6909,N_1453,N_3062);
or U6910 (N_6910,N_3792,N_4106);
or U6911 (N_6911,N_777,N_4826);
nand U6912 (N_6912,N_4032,N_1242);
or U6913 (N_6913,N_2917,N_1807);
nand U6914 (N_6914,N_2295,N_2002);
xnor U6915 (N_6915,N_3496,N_2536);
and U6916 (N_6916,N_2990,N_508);
nor U6917 (N_6917,N_4758,N_3153);
nor U6918 (N_6918,N_54,N_1639);
or U6919 (N_6919,N_1783,N_2112);
nor U6920 (N_6920,N_4209,N_1853);
nand U6921 (N_6921,N_3811,N_4797);
or U6922 (N_6922,N_789,N_195);
nand U6923 (N_6923,N_3648,N_3593);
or U6924 (N_6924,N_4817,N_1870);
and U6925 (N_6925,N_4408,N_3192);
nand U6926 (N_6926,N_2525,N_1606);
and U6927 (N_6927,N_3321,N_4976);
nor U6928 (N_6928,N_4316,N_1534);
nand U6929 (N_6929,N_3391,N_4647);
or U6930 (N_6930,N_4286,N_2842);
nand U6931 (N_6931,N_3639,N_4879);
nand U6932 (N_6932,N_1802,N_2312);
or U6933 (N_6933,N_591,N_147);
or U6934 (N_6934,N_2576,N_3434);
or U6935 (N_6935,N_923,N_1729);
and U6936 (N_6936,N_739,N_3793);
or U6937 (N_6937,N_3159,N_3098);
nand U6938 (N_6938,N_44,N_846);
or U6939 (N_6939,N_2167,N_1317);
nor U6940 (N_6940,N_1357,N_2251);
nor U6941 (N_6941,N_41,N_3253);
nand U6942 (N_6942,N_4863,N_776);
nand U6943 (N_6943,N_3660,N_1393);
nor U6944 (N_6944,N_2019,N_1698);
nor U6945 (N_6945,N_248,N_4109);
or U6946 (N_6946,N_3951,N_4984);
xnor U6947 (N_6947,N_3547,N_2158);
or U6948 (N_6948,N_3566,N_4205);
or U6949 (N_6949,N_3821,N_2234);
and U6950 (N_6950,N_237,N_2298);
and U6951 (N_6951,N_1158,N_1431);
and U6952 (N_6952,N_1667,N_4791);
and U6953 (N_6953,N_3407,N_577);
and U6954 (N_6954,N_1746,N_3357);
nand U6955 (N_6955,N_1348,N_1910);
nand U6956 (N_6956,N_2720,N_3330);
nor U6957 (N_6957,N_1324,N_1937);
xor U6958 (N_6958,N_3248,N_2568);
nor U6959 (N_6959,N_4334,N_20);
nand U6960 (N_6960,N_2152,N_4168);
nand U6961 (N_6961,N_867,N_2535);
or U6962 (N_6962,N_4970,N_3236);
xor U6963 (N_6963,N_4608,N_1346);
and U6964 (N_6964,N_1681,N_2261);
or U6965 (N_6965,N_2344,N_4601);
nand U6966 (N_6966,N_4670,N_1188);
nor U6967 (N_6967,N_4916,N_4559);
nand U6968 (N_6968,N_1742,N_4481);
nor U6969 (N_6969,N_1651,N_590);
or U6970 (N_6970,N_659,N_947);
nor U6971 (N_6971,N_2263,N_4175);
nand U6972 (N_6972,N_1714,N_392);
nand U6973 (N_6973,N_929,N_2384);
and U6974 (N_6974,N_308,N_1595);
nor U6975 (N_6975,N_315,N_4234);
or U6976 (N_6976,N_4524,N_43);
and U6977 (N_6977,N_2952,N_198);
nand U6978 (N_6978,N_51,N_4312);
nand U6979 (N_6979,N_2599,N_567);
nor U6980 (N_6980,N_3462,N_1692);
and U6981 (N_6981,N_3332,N_3177);
nor U6982 (N_6982,N_2458,N_1312);
xnor U6983 (N_6983,N_693,N_279);
nand U6984 (N_6984,N_2395,N_4086);
nor U6985 (N_6985,N_2511,N_1961);
and U6986 (N_6986,N_799,N_2880);
nand U6987 (N_6987,N_3432,N_2504);
nand U6988 (N_6988,N_893,N_3490);
nor U6989 (N_6989,N_135,N_3113);
and U6990 (N_6990,N_631,N_2103);
or U6991 (N_6991,N_1311,N_4844);
nor U6992 (N_6992,N_191,N_3444);
nor U6993 (N_6993,N_4007,N_1489);
or U6994 (N_6994,N_1863,N_2940);
nor U6995 (N_6995,N_3096,N_2886);
nor U6996 (N_6996,N_4517,N_1750);
nor U6997 (N_6997,N_1629,N_2256);
nor U6998 (N_6998,N_3006,N_4783);
nor U6999 (N_6999,N_704,N_3549);
or U7000 (N_7000,N_1055,N_595);
xor U7001 (N_7001,N_2421,N_3473);
nor U7002 (N_7002,N_3455,N_4137);
nor U7003 (N_7003,N_4390,N_1443);
nand U7004 (N_7004,N_4048,N_4378);
and U7005 (N_7005,N_110,N_3619);
or U7006 (N_7006,N_3676,N_1239);
nor U7007 (N_7007,N_4926,N_4539);
or U7008 (N_7008,N_4732,N_35);
xnor U7009 (N_7009,N_1858,N_4924);
nand U7010 (N_7010,N_986,N_2389);
nor U7011 (N_7011,N_4945,N_3155);
nor U7012 (N_7012,N_160,N_4120);
and U7013 (N_7013,N_327,N_2127);
nand U7014 (N_7014,N_4852,N_2656);
nor U7015 (N_7015,N_2970,N_3933);
xnor U7016 (N_7016,N_3,N_4331);
or U7017 (N_7017,N_1829,N_2377);
and U7018 (N_7018,N_1375,N_3856);
nand U7019 (N_7019,N_3122,N_3143);
and U7020 (N_7020,N_2730,N_1582);
nor U7021 (N_7021,N_2121,N_2696);
and U7022 (N_7022,N_30,N_3638);
nand U7023 (N_7023,N_2884,N_2943);
and U7024 (N_7024,N_3617,N_2686);
nor U7025 (N_7025,N_3457,N_1548);
nand U7026 (N_7026,N_4499,N_699);
nand U7027 (N_7027,N_3262,N_2567);
nor U7028 (N_7028,N_3847,N_1314);
xor U7029 (N_7029,N_4308,N_1628);
and U7030 (N_7030,N_3911,N_1976);
and U7031 (N_7031,N_4909,N_3388);
xor U7032 (N_7032,N_2093,N_4615);
nand U7033 (N_7033,N_140,N_4972);
or U7034 (N_7034,N_2684,N_1151);
and U7035 (N_7035,N_3542,N_3481);
nand U7036 (N_7036,N_837,N_791);
and U7037 (N_7037,N_4540,N_1652);
nand U7038 (N_7038,N_2227,N_2130);
and U7039 (N_7039,N_1847,N_2796);
or U7040 (N_7040,N_427,N_3247);
xor U7041 (N_7041,N_3285,N_2000);
nand U7042 (N_7042,N_4939,N_981);
and U7043 (N_7043,N_3435,N_1037);
and U7044 (N_7044,N_1017,N_2225);
xor U7045 (N_7045,N_2343,N_2494);
or U7046 (N_7046,N_1722,N_2441);
nand U7047 (N_7047,N_1569,N_527);
or U7048 (N_7048,N_4565,N_96);
nand U7049 (N_7049,N_4131,N_2868);
and U7050 (N_7050,N_734,N_1564);
nor U7051 (N_7051,N_4413,N_3438);
nand U7052 (N_7052,N_2437,N_200);
and U7053 (N_7053,N_473,N_1579);
xor U7054 (N_7054,N_435,N_4447);
nor U7055 (N_7055,N_2957,N_1770);
nor U7056 (N_7056,N_3632,N_3121);
and U7057 (N_7057,N_3592,N_1598);
nand U7058 (N_7058,N_2211,N_2072);
nand U7059 (N_7059,N_3105,N_3394);
nor U7060 (N_7060,N_3361,N_2144);
nand U7061 (N_7061,N_4822,N_2647);
nand U7062 (N_7062,N_3993,N_2215);
nor U7063 (N_7063,N_3068,N_4099);
and U7064 (N_7064,N_4739,N_3017);
and U7065 (N_7065,N_1358,N_2279);
or U7066 (N_7066,N_233,N_282);
and U7067 (N_7067,N_2134,N_1927);
or U7068 (N_7068,N_1786,N_1202);
or U7069 (N_7069,N_1726,N_903);
nand U7070 (N_7070,N_865,N_261);
and U7071 (N_7071,N_1771,N_796);
or U7072 (N_7072,N_4905,N_1089);
or U7073 (N_7073,N_714,N_1119);
nor U7074 (N_7074,N_4124,N_2238);
or U7075 (N_7075,N_3517,N_1250);
or U7076 (N_7076,N_2867,N_850);
nor U7077 (N_7077,N_2874,N_3219);
and U7078 (N_7078,N_1221,N_1480);
or U7079 (N_7079,N_832,N_664);
and U7080 (N_7080,N_3816,N_4353);
and U7081 (N_7081,N_3704,N_1576);
and U7082 (N_7082,N_2980,N_2058);
nor U7083 (N_7083,N_674,N_1005);
and U7084 (N_7084,N_554,N_4929);
nor U7085 (N_7085,N_1967,N_3069);
and U7086 (N_7086,N_3427,N_3649);
nand U7087 (N_7087,N_2989,N_980);
nor U7088 (N_7088,N_312,N_4037);
nor U7089 (N_7089,N_2600,N_3858);
xnor U7090 (N_7090,N_2081,N_1857);
and U7091 (N_7091,N_3868,N_412);
nor U7092 (N_7092,N_49,N_4173);
nand U7093 (N_7093,N_2735,N_3766);
and U7094 (N_7094,N_2875,N_2681);
xor U7095 (N_7095,N_1174,N_2781);
xnor U7096 (N_7096,N_165,N_1654);
nand U7097 (N_7097,N_186,N_148);
nand U7098 (N_7098,N_2306,N_4618);
or U7099 (N_7099,N_454,N_3783);
or U7100 (N_7100,N_1172,N_458);
nand U7101 (N_7101,N_1288,N_1394);
or U7102 (N_7102,N_290,N_2644);
nor U7103 (N_7103,N_534,N_2551);
or U7104 (N_7104,N_1409,N_2530);
and U7105 (N_7105,N_2414,N_3754);
or U7106 (N_7106,N_2668,N_1337);
or U7107 (N_7107,N_159,N_2480);
nand U7108 (N_7108,N_3273,N_4301);
and U7109 (N_7109,N_1080,N_297);
xor U7110 (N_7110,N_3901,N_3893);
nor U7111 (N_7111,N_805,N_2814);
nand U7112 (N_7112,N_4466,N_1035);
and U7113 (N_7113,N_4616,N_3292);
nor U7114 (N_7114,N_1960,N_1702);
nor U7115 (N_7115,N_4344,N_1803);
nor U7116 (N_7116,N_926,N_1124);
nor U7117 (N_7117,N_4384,N_1648);
or U7118 (N_7118,N_4707,N_278);
nor U7119 (N_7119,N_1740,N_544);
nor U7120 (N_7120,N_758,N_2650);
and U7121 (N_7121,N_584,N_1641);
or U7122 (N_7122,N_1864,N_2166);
and U7123 (N_7123,N_4523,N_1363);
or U7124 (N_7124,N_4849,N_1353);
and U7125 (N_7125,N_3824,N_1469);
or U7126 (N_7126,N_1602,N_2067);
xor U7127 (N_7127,N_4695,N_1425);
nor U7128 (N_7128,N_2564,N_3310);
xor U7129 (N_7129,N_3120,N_3681);
nand U7130 (N_7130,N_3107,N_4074);
and U7131 (N_7131,N_1262,N_1908);
nor U7132 (N_7132,N_2008,N_1848);
and U7133 (N_7133,N_4151,N_176);
nand U7134 (N_7134,N_1580,N_4896);
and U7135 (N_7135,N_511,N_2321);
or U7136 (N_7136,N_4229,N_1885);
nand U7137 (N_7137,N_1609,N_2652);
and U7138 (N_7138,N_4528,N_4051);
or U7139 (N_7139,N_4061,N_3301);
and U7140 (N_7140,N_347,N_2869);
and U7141 (N_7141,N_652,N_3559);
and U7142 (N_7142,N_2098,N_236);
xor U7143 (N_7143,N_4775,N_1457);
and U7144 (N_7144,N_3718,N_2911);
nand U7145 (N_7145,N_4326,N_1923);
and U7146 (N_7146,N_991,N_1504);
nor U7147 (N_7147,N_2802,N_1637);
and U7148 (N_7148,N_678,N_775);
or U7149 (N_7149,N_4386,N_3254);
and U7150 (N_7150,N_1695,N_169);
or U7151 (N_7151,N_2341,N_4660);
nand U7152 (N_7152,N_2011,N_3701);
and U7153 (N_7153,N_2693,N_3706);
nor U7154 (N_7154,N_3720,N_1142);
xor U7155 (N_7155,N_3380,N_4632);
and U7156 (N_7156,N_2120,N_1390);
nand U7157 (N_7157,N_4810,N_1769);
and U7158 (N_7158,N_4737,N_4754);
nand U7159 (N_7159,N_4701,N_3209);
xor U7160 (N_7160,N_193,N_3138);
or U7161 (N_7161,N_4338,N_1475);
and U7162 (N_7162,N_4298,N_645);
nor U7163 (N_7163,N_3616,N_2694);
nor U7164 (N_7164,N_4049,N_420);
nor U7165 (N_7165,N_1257,N_1627);
nand U7166 (N_7166,N_1219,N_1522);
and U7167 (N_7167,N_4561,N_4148);
and U7168 (N_7168,N_2243,N_2334);
and U7169 (N_7169,N_2608,N_4383);
and U7170 (N_7170,N_856,N_817);
nand U7171 (N_7171,N_2466,N_2172);
nor U7172 (N_7172,N_2794,N_1719);
nand U7173 (N_7173,N_2131,N_2006);
xor U7174 (N_7174,N_3628,N_3938);
nor U7175 (N_7175,N_4026,N_334);
and U7176 (N_7176,N_705,N_641);
and U7177 (N_7177,N_366,N_3507);
nor U7178 (N_7178,N_4272,N_4273);
nor U7179 (N_7179,N_3803,N_3223);
or U7180 (N_7180,N_88,N_4046);
xor U7181 (N_7181,N_2452,N_1466);
or U7182 (N_7182,N_3520,N_1230);
nor U7183 (N_7183,N_405,N_4873);
nor U7184 (N_7184,N_3374,N_4372);
and U7185 (N_7185,N_3172,N_2664);
nor U7186 (N_7186,N_3423,N_1794);
and U7187 (N_7187,N_1873,N_3525);
or U7188 (N_7188,N_82,N_2905);
nand U7189 (N_7189,N_4779,N_2837);
xnor U7190 (N_7190,N_4734,N_2955);
nor U7191 (N_7191,N_4527,N_3791);
and U7192 (N_7192,N_3897,N_1004);
and U7193 (N_7193,N_3861,N_3303);
or U7194 (N_7194,N_1664,N_4679);
and U7195 (N_7195,N_1249,N_4643);
and U7196 (N_7196,N_238,N_2831);
xor U7197 (N_7197,N_2049,N_884);
and U7198 (N_7198,N_2553,N_3297);
or U7199 (N_7199,N_1179,N_3372);
or U7200 (N_7200,N_2185,N_155);
or U7201 (N_7201,N_1773,N_1442);
nor U7202 (N_7202,N_604,N_4991);
or U7203 (N_7203,N_2349,N_1536);
and U7204 (N_7204,N_4038,N_4490);
nand U7205 (N_7205,N_4419,N_2544);
nor U7206 (N_7206,N_4623,N_2679);
nor U7207 (N_7207,N_4842,N_4092);
nand U7208 (N_7208,N_914,N_1182);
and U7209 (N_7209,N_592,N_1079);
and U7210 (N_7210,N_4489,N_576);
or U7211 (N_7211,N_2118,N_4597);
nand U7212 (N_7212,N_324,N_1792);
or U7213 (N_7213,N_3280,N_1141);
and U7214 (N_7214,N_1271,N_4420);
nor U7215 (N_7215,N_3210,N_1371);
and U7216 (N_7216,N_3318,N_1168);
nand U7217 (N_7217,N_2846,N_3360);
or U7218 (N_7218,N_2434,N_4400);
nor U7219 (N_7219,N_4302,N_2795);
nor U7220 (N_7220,N_2898,N_4675);
and U7221 (N_7221,N_2406,N_3674);
nor U7222 (N_7222,N_4052,N_3383);
and U7223 (N_7223,N_4589,N_1806);
nor U7224 (N_7224,N_3061,N_1264);
nand U7225 (N_7225,N_1436,N_2692);
or U7226 (N_7226,N_3714,N_2558);
nor U7227 (N_7227,N_2297,N_2358);
nand U7228 (N_7228,N_393,N_1155);
nor U7229 (N_7229,N_2968,N_4799);
or U7230 (N_7230,N_2022,N_951);
nor U7231 (N_7231,N_3437,N_3784);
or U7232 (N_7232,N_3475,N_1945);
nor U7233 (N_7233,N_1889,N_2432);
nand U7234 (N_7234,N_908,N_3497);
xor U7235 (N_7235,N_935,N_1618);
and U7236 (N_7236,N_130,N_2744);
or U7237 (N_7237,N_3519,N_1573);
or U7238 (N_7238,N_4108,N_573);
or U7239 (N_7239,N_4834,N_3091);
nand U7240 (N_7240,N_851,N_1160);
nand U7241 (N_7241,N_2977,N_4536);
nor U7242 (N_7242,N_1672,N_409);
xor U7243 (N_7243,N_1539,N_173);
and U7244 (N_7244,N_3580,N_1819);
nor U7245 (N_7245,N_1957,N_2534);
nand U7246 (N_7246,N_153,N_2909);
nand U7247 (N_7247,N_4213,N_1082);
nand U7248 (N_7248,N_4767,N_4215);
xnor U7249 (N_7249,N_2715,N_1460);
nand U7250 (N_7250,N_4551,N_1597);
and U7251 (N_7251,N_1640,N_828);
xor U7252 (N_7252,N_2122,N_2090);
and U7253 (N_7253,N_4245,N_1256);
nor U7254 (N_7254,N_3112,N_3540);
xnor U7255 (N_7255,N_1391,N_1493);
nand U7256 (N_7256,N_213,N_4348);
xnor U7257 (N_7257,N_1075,N_2661);
or U7258 (N_7258,N_4911,N_2934);
xor U7259 (N_7259,N_1626,N_1909);
nor U7260 (N_7260,N_2583,N_4764);
nor U7261 (N_7261,N_2420,N_4587);
nor U7262 (N_7262,N_360,N_4226);
and U7263 (N_7263,N_2510,N_710);
or U7264 (N_7264,N_3755,N_90);
and U7265 (N_7265,N_3281,N_1533);
or U7266 (N_7266,N_1706,N_1482);
nand U7267 (N_7267,N_368,N_2603);
nor U7268 (N_7268,N_4356,N_4985);
and U7269 (N_7269,N_107,N_2541);
nand U7270 (N_7270,N_351,N_1330);
and U7271 (N_7271,N_1368,N_3779);
nor U7272 (N_7272,N_1278,N_2546);
nand U7273 (N_7273,N_1154,N_1429);
nor U7274 (N_7274,N_2733,N_3597);
nand U7275 (N_7275,N_622,N_2707);
or U7276 (N_7276,N_2703,N_4147);
or U7277 (N_7277,N_172,N_4993);
and U7278 (N_7278,N_3680,N_833);
or U7279 (N_7279,N_2010,N_784);
xnor U7280 (N_7280,N_1869,N_4663);
nor U7281 (N_7281,N_3505,N_4760);
nor U7282 (N_7282,N_1933,N_2401);
or U7283 (N_7283,N_2984,N_624);
and U7284 (N_7284,N_4912,N_1523);
nand U7285 (N_7285,N_1615,N_529);
nand U7286 (N_7286,N_682,N_792);
nor U7287 (N_7287,N_4697,N_2779);
and U7288 (N_7288,N_689,N_221);
or U7289 (N_7289,N_3656,N_3334);
xor U7290 (N_7290,N_2328,N_3985);
and U7291 (N_7291,N_2539,N_3658);
and U7292 (N_7292,N_3401,N_2723);
and U7293 (N_7293,N_925,N_1778);
nand U7294 (N_7294,N_2275,N_669);
and U7295 (N_7295,N_706,N_3298);
or U7296 (N_7296,N_3518,N_3024);
and U7297 (N_7297,N_1169,N_3894);
nor U7298 (N_7298,N_19,N_2628);
nor U7299 (N_7299,N_1755,N_11);
nor U7300 (N_7300,N_2596,N_4545);
or U7301 (N_7301,N_1868,N_3140);
nor U7302 (N_7302,N_1417,N_1091);
nand U7303 (N_7303,N_4581,N_709);
nand U7304 (N_7304,N_844,N_4036);
nand U7305 (N_7305,N_894,N_1890);
nor U7306 (N_7306,N_322,N_1781);
and U7307 (N_7307,N_4894,N_1661);
and U7308 (N_7308,N_1045,N_3711);
and U7309 (N_7309,N_3442,N_1715);
and U7310 (N_7310,N_2713,N_4479);
or U7311 (N_7311,N_4897,N_2475);
or U7312 (N_7312,N_2697,N_3963);
xor U7313 (N_7313,N_48,N_3998);
and U7314 (N_7314,N_1341,N_371);
xor U7315 (N_7315,N_1922,N_466);
or U7316 (N_7316,N_3108,N_4941);
or U7317 (N_7317,N_423,N_726);
nand U7318 (N_7318,N_2745,N_1830);
xnor U7319 (N_7319,N_4171,N_3003);
or U7320 (N_7320,N_3365,N_2804);
nor U7321 (N_7321,N_2397,N_4968);
nor U7322 (N_7322,N_2969,N_2998);
and U7323 (N_7323,N_1343,N_162);
xnor U7324 (N_7324,N_2908,N_2479);
or U7325 (N_7325,N_3555,N_2887);
nand U7326 (N_7326,N_2059,N_1251);
nor U7327 (N_7327,N_464,N_2467);
nor U7328 (N_7328,N_2924,N_3968);
nand U7329 (N_7329,N_400,N_4773);
or U7330 (N_7330,N_2175,N_4246);
nand U7331 (N_7331,N_1218,N_2446);
and U7332 (N_7332,N_574,N_863);
and U7333 (N_7333,N_2411,N_2865);
and U7334 (N_7334,N_1517,N_3702);
nor U7335 (N_7335,N_1420,N_790);
xor U7336 (N_7336,N_2063,N_3458);
nor U7337 (N_7337,N_452,N_3340);
or U7338 (N_7338,N_1232,N_2136);
nand U7339 (N_7339,N_205,N_1901);
or U7340 (N_7340,N_1799,N_28);
nor U7341 (N_7341,N_3440,N_1572);
or U7342 (N_7342,N_801,N_1701);
xor U7343 (N_7343,N_252,N_3528);
or U7344 (N_7344,N_2052,N_3825);
and U7345 (N_7345,N_4935,N_247);
nor U7346 (N_7346,N_2882,N_1002);
and U7347 (N_7347,N_432,N_602);
and U7348 (N_7348,N_3309,N_3282);
or U7349 (N_7349,N_316,N_677);
and U7350 (N_7350,N_2269,N_3719);
nor U7351 (N_7351,N_1838,N_2069);
xor U7352 (N_7352,N_1635,N_3867);
nand U7353 (N_7353,N_1333,N_4910);
nor U7354 (N_7354,N_1260,N_413);
xor U7355 (N_7355,N_1126,N_4006);
and U7356 (N_7356,N_1861,N_3577);
nor U7357 (N_7357,N_2371,N_24);
or U7358 (N_7358,N_4188,N_2346);
or U7359 (N_7359,N_520,N_4691);
or U7360 (N_7360,N_1468,N_2382);
nor U7361 (N_7361,N_4999,N_3348);
or U7362 (N_7362,N_2540,N_794);
and U7363 (N_7363,N_2518,N_971);
nor U7364 (N_7364,N_306,N_1003);
nor U7365 (N_7365,N_3760,N_314);
or U7366 (N_7366,N_2910,N_549);
or U7367 (N_7367,N_1432,N_4203);
and U7368 (N_7368,N_3723,N_3554);
nor U7369 (N_7369,N_4401,N_1054);
nor U7370 (N_7370,N_3422,N_4944);
nand U7371 (N_7371,N_3086,N_2125);
xor U7372 (N_7372,N_4563,N_1821);
nor U7373 (N_7373,N_2378,N_1143);
xnor U7374 (N_7374,N_75,N_2083);
nand U7375 (N_7375,N_3142,N_2488);
nand U7376 (N_7376,N_3902,N_3447);
nor U7377 (N_7377,N_1840,N_3568);
and U7378 (N_7378,N_1322,N_1712);
or U7379 (N_7379,N_1514,N_944);
and U7380 (N_7380,N_1272,N_3164);
xor U7381 (N_7381,N_4971,N_990);
nor U7382 (N_7382,N_2046,N_3362);
nor U7383 (N_7383,N_1623,N_2450);
and U7384 (N_7384,N_2844,N_3324);
nor U7385 (N_7385,N_3934,N_2586);
or U7386 (N_7386,N_1008,N_3892);
nor U7387 (N_7387,N_2933,N_3492);
nand U7388 (N_7388,N_2548,N_2005);
or U7389 (N_7389,N_958,N_451);
and U7390 (N_7390,N_3574,N_182);
xnor U7391 (N_7391,N_211,N_1404);
or U7392 (N_7392,N_4942,N_232);
and U7393 (N_7393,N_73,N_4350);
nand U7394 (N_7394,N_1939,N_4904);
xnor U7395 (N_7395,N_3634,N_3872);
nand U7396 (N_7396,N_873,N_3260);
and U7397 (N_7397,N_1500,N_4247);
and U7398 (N_7398,N_4672,N_1189);
xor U7399 (N_7399,N_2883,N_2876);
nor U7400 (N_7400,N_4923,N_1153);
or U7401 (N_7401,N_2123,N_106);
and U7402 (N_7402,N_378,N_2486);
nor U7403 (N_7403,N_2906,N_4965);
nor U7404 (N_7404,N_1139,N_1112);
nor U7405 (N_7405,N_1666,N_1506);
nor U7406 (N_7406,N_3621,N_2950);
nand U7407 (N_7407,N_1647,N_1123);
and U7408 (N_7408,N_4550,N_1027);
xnor U7409 (N_7409,N_399,N_996);
nand U7410 (N_7410,N_4135,N_2607);
and U7411 (N_7411,N_123,N_2888);
nor U7412 (N_7412,N_175,N_2037);
and U7413 (N_7413,N_3037,N_4717);
or U7414 (N_7414,N_697,N_3331);
xnor U7415 (N_7415,N_68,N_2154);
nand U7416 (N_7416,N_2500,N_1447);
nand U7417 (N_7417,N_4599,N_254);
nand U7418 (N_7418,N_2636,N_2079);
nor U7419 (N_7419,N_303,N_3306);
nor U7420 (N_7420,N_1994,N_2193);
and U7421 (N_7421,N_4995,N_3812);
and U7422 (N_7422,N_1277,N_3795);
or U7423 (N_7423,N_2039,N_4917);
nand U7424 (N_7424,N_2338,N_4299);
nor U7425 (N_7425,N_564,N_2682);
nand U7426 (N_7426,N_3924,N_4867);
nand U7427 (N_7427,N_3846,N_814);
nor U7428 (N_7428,N_4377,N_3354);
nand U7429 (N_7429,N_2747,N_3368);
nand U7430 (N_7430,N_2963,N_3252);
and U7431 (N_7431,N_4405,N_978);
nand U7432 (N_7432,N_1570,N_4633);
nand U7433 (N_7433,N_2508,N_2352);
xor U7434 (N_7434,N_4963,N_2363);
nand U7435 (N_7435,N_597,N_2889);
and U7436 (N_7436,N_408,N_1753);
nor U7437 (N_7437,N_633,N_3921);
nor U7438 (N_7438,N_2750,N_1984);
nor U7439 (N_7439,N_3092,N_3834);
nand U7440 (N_7440,N_4746,N_4997);
and U7441 (N_7441,N_4839,N_3510);
nor U7442 (N_7442,N_3225,N_931);
nor U7443 (N_7443,N_2216,N_4127);
and U7444 (N_7444,N_3563,N_593);
nor U7445 (N_7445,N_623,N_4017);
nand U7446 (N_7446,N_319,N_3584);
or U7447 (N_7447,N_3753,N_4936);
nand U7448 (N_7448,N_2792,N_4685);
nor U7449 (N_7449,N_2931,N_3761);
or U7450 (N_7450,N_1684,N_1421);
nand U7451 (N_7451,N_3885,N_2013);
or U7452 (N_7452,N_2821,N_1928);
nand U7453 (N_7453,N_149,N_1859);
or U7454 (N_7454,N_1125,N_4228);
or U7455 (N_7455,N_2226,N_3947);
and U7456 (N_7456,N_4693,N_4253);
or U7457 (N_7457,N_2018,N_2569);
or U7458 (N_7458,N_398,N_1118);
or U7459 (N_7459,N_4636,N_2001);
nor U7460 (N_7460,N_4358,N_3425);
or U7461 (N_7461,N_961,N_3572);
or U7462 (N_7462,N_2023,N_1983);
and U7463 (N_7463,N_960,N_4269);
and U7464 (N_7464,N_3016,N_4104);
xnor U7465 (N_7465,N_3188,N_1925);
or U7466 (N_7466,N_4814,N_1725);
and U7467 (N_7467,N_1059,N_4211);
xnor U7468 (N_7468,N_2190,N_3012);
nand U7469 (N_7469,N_4176,N_3315);
nor U7470 (N_7470,N_2054,N_4918);
and U7471 (N_7471,N_495,N_4416);
and U7472 (N_7472,N_4297,N_3468);
nand U7473 (N_7473,N_3410,N_3558);
or U7474 (N_7474,N_1758,N_1023);
or U7475 (N_7475,N_2527,N_1226);
and U7476 (N_7476,N_3844,N_2137);
and U7477 (N_7477,N_4373,N_2179);
nand U7478 (N_7478,N_4042,N_471);
and U7479 (N_7479,N_1752,N_4574);
nor U7480 (N_7480,N_4256,N_2339);
or U7481 (N_7481,N_2502,N_1650);
nor U7482 (N_7482,N_3478,N_141);
nand U7483 (N_7483,N_4097,N_486);
and U7484 (N_7484,N_4404,N_3031);
or U7485 (N_7485,N_569,N_3955);
or U7486 (N_7486,N_3522,N_3688);
nand U7487 (N_7487,N_4614,N_52);
nor U7488 (N_7488,N_109,N_4293);
xor U7489 (N_7489,N_3165,N_406);
and U7490 (N_7490,N_1973,N_3653);
nand U7491 (N_7491,N_510,N_2025);
or U7492 (N_7492,N_4095,N_4629);
nor U7493 (N_7493,N_461,N_2456);
nand U7494 (N_7494,N_3403,N_4722);
nor U7495 (N_7495,N_78,N_4279);
and U7496 (N_7496,N_1382,N_4694);
nor U7497 (N_7497,N_4098,N_936);
and U7498 (N_7498,N_3075,N_4552);
xor U7499 (N_7499,N_2435,N_2278);
nor U7500 (N_7500,N_2616,N_4248);
nor U7501 (N_7501,N_4091,N_2123);
and U7502 (N_7502,N_2834,N_3829);
nand U7503 (N_7503,N_1264,N_1186);
or U7504 (N_7504,N_3301,N_877);
nand U7505 (N_7505,N_3043,N_970);
or U7506 (N_7506,N_4584,N_1711);
or U7507 (N_7507,N_4792,N_702);
or U7508 (N_7508,N_1450,N_3622);
or U7509 (N_7509,N_1082,N_866);
nand U7510 (N_7510,N_731,N_906);
nand U7511 (N_7511,N_3668,N_1119);
or U7512 (N_7512,N_2177,N_3749);
or U7513 (N_7513,N_3730,N_3400);
and U7514 (N_7514,N_436,N_1489);
nor U7515 (N_7515,N_1506,N_2847);
nand U7516 (N_7516,N_2734,N_1110);
nand U7517 (N_7517,N_382,N_2474);
nand U7518 (N_7518,N_1558,N_342);
or U7519 (N_7519,N_1467,N_4511);
or U7520 (N_7520,N_4730,N_4048);
nor U7521 (N_7521,N_2102,N_913);
or U7522 (N_7522,N_510,N_490);
nand U7523 (N_7523,N_1911,N_3520);
or U7524 (N_7524,N_3132,N_220);
xnor U7525 (N_7525,N_3181,N_1538);
or U7526 (N_7526,N_675,N_2450);
nor U7527 (N_7527,N_332,N_3650);
nor U7528 (N_7528,N_381,N_167);
nand U7529 (N_7529,N_3492,N_3272);
and U7530 (N_7530,N_738,N_3407);
nor U7531 (N_7531,N_4846,N_4095);
and U7532 (N_7532,N_4149,N_2371);
xnor U7533 (N_7533,N_936,N_3040);
and U7534 (N_7534,N_4083,N_1012);
xnor U7535 (N_7535,N_408,N_808);
nor U7536 (N_7536,N_2259,N_4210);
nor U7537 (N_7537,N_1006,N_3134);
and U7538 (N_7538,N_3455,N_494);
or U7539 (N_7539,N_2178,N_3517);
or U7540 (N_7540,N_1040,N_2255);
nor U7541 (N_7541,N_616,N_117);
xor U7542 (N_7542,N_3916,N_864);
or U7543 (N_7543,N_4905,N_2991);
nor U7544 (N_7544,N_3366,N_182);
and U7545 (N_7545,N_1822,N_3405);
and U7546 (N_7546,N_1635,N_4184);
or U7547 (N_7547,N_821,N_1260);
nand U7548 (N_7548,N_2294,N_2654);
nor U7549 (N_7549,N_2245,N_1678);
and U7550 (N_7550,N_3930,N_2269);
nor U7551 (N_7551,N_4250,N_4967);
and U7552 (N_7552,N_85,N_1322);
xor U7553 (N_7553,N_3123,N_3660);
nor U7554 (N_7554,N_2885,N_4274);
nand U7555 (N_7555,N_4860,N_493);
nand U7556 (N_7556,N_1748,N_783);
nand U7557 (N_7557,N_2951,N_115);
nand U7558 (N_7558,N_3397,N_3204);
or U7559 (N_7559,N_1106,N_2996);
nor U7560 (N_7560,N_4815,N_4397);
or U7561 (N_7561,N_2220,N_4836);
nand U7562 (N_7562,N_1836,N_947);
xnor U7563 (N_7563,N_2610,N_2449);
nand U7564 (N_7564,N_431,N_3257);
nand U7565 (N_7565,N_1923,N_2011);
nor U7566 (N_7566,N_4485,N_1183);
and U7567 (N_7567,N_2716,N_821);
and U7568 (N_7568,N_1818,N_658);
nand U7569 (N_7569,N_3575,N_3256);
and U7570 (N_7570,N_3357,N_282);
and U7571 (N_7571,N_661,N_2062);
nand U7572 (N_7572,N_3408,N_3479);
xor U7573 (N_7573,N_2250,N_1);
or U7574 (N_7574,N_1353,N_4966);
nand U7575 (N_7575,N_1462,N_1652);
or U7576 (N_7576,N_3602,N_2774);
or U7577 (N_7577,N_4951,N_2256);
or U7578 (N_7578,N_3251,N_3868);
nor U7579 (N_7579,N_2730,N_963);
and U7580 (N_7580,N_3167,N_1117);
and U7581 (N_7581,N_4104,N_2063);
nand U7582 (N_7582,N_914,N_1369);
or U7583 (N_7583,N_3728,N_4234);
nand U7584 (N_7584,N_2952,N_3870);
xor U7585 (N_7585,N_4173,N_118);
nor U7586 (N_7586,N_92,N_2482);
nand U7587 (N_7587,N_2977,N_1579);
nor U7588 (N_7588,N_3013,N_4579);
or U7589 (N_7589,N_2103,N_3297);
nor U7590 (N_7590,N_3095,N_272);
or U7591 (N_7591,N_301,N_2153);
and U7592 (N_7592,N_3797,N_473);
or U7593 (N_7593,N_742,N_338);
and U7594 (N_7594,N_321,N_2059);
nor U7595 (N_7595,N_1514,N_1092);
and U7596 (N_7596,N_1308,N_4861);
or U7597 (N_7597,N_4847,N_1974);
or U7598 (N_7598,N_3547,N_491);
and U7599 (N_7599,N_4663,N_173);
nand U7600 (N_7600,N_3725,N_855);
nand U7601 (N_7601,N_709,N_2323);
nor U7602 (N_7602,N_4671,N_3628);
nand U7603 (N_7603,N_2995,N_1449);
and U7604 (N_7604,N_4244,N_76);
nand U7605 (N_7605,N_1607,N_3469);
nand U7606 (N_7606,N_544,N_938);
and U7607 (N_7607,N_3222,N_139);
xor U7608 (N_7608,N_2608,N_1061);
xnor U7609 (N_7609,N_4651,N_3985);
or U7610 (N_7610,N_4776,N_2597);
nand U7611 (N_7611,N_4882,N_1334);
and U7612 (N_7612,N_3917,N_1852);
xnor U7613 (N_7613,N_470,N_216);
nand U7614 (N_7614,N_1841,N_3163);
nand U7615 (N_7615,N_3772,N_4709);
and U7616 (N_7616,N_4243,N_503);
or U7617 (N_7617,N_4794,N_3525);
nor U7618 (N_7618,N_3294,N_1246);
xnor U7619 (N_7619,N_3879,N_1033);
xor U7620 (N_7620,N_706,N_4368);
nor U7621 (N_7621,N_3906,N_1552);
nor U7622 (N_7622,N_1966,N_2516);
nand U7623 (N_7623,N_3405,N_4397);
and U7624 (N_7624,N_1343,N_4764);
xnor U7625 (N_7625,N_379,N_3093);
and U7626 (N_7626,N_487,N_4310);
or U7627 (N_7627,N_4413,N_4158);
nor U7628 (N_7628,N_4896,N_4508);
nor U7629 (N_7629,N_2541,N_1396);
or U7630 (N_7630,N_4308,N_1422);
and U7631 (N_7631,N_4269,N_318);
nand U7632 (N_7632,N_4949,N_1450);
and U7633 (N_7633,N_1813,N_3480);
or U7634 (N_7634,N_1618,N_1607);
nor U7635 (N_7635,N_1832,N_1191);
or U7636 (N_7636,N_3589,N_2216);
nand U7637 (N_7637,N_61,N_2728);
and U7638 (N_7638,N_4330,N_2165);
xor U7639 (N_7639,N_1670,N_3242);
or U7640 (N_7640,N_3458,N_2863);
nor U7641 (N_7641,N_2690,N_2976);
xor U7642 (N_7642,N_2052,N_1089);
nor U7643 (N_7643,N_168,N_3444);
or U7644 (N_7644,N_789,N_4427);
nor U7645 (N_7645,N_1834,N_4405);
and U7646 (N_7646,N_1050,N_1749);
or U7647 (N_7647,N_3659,N_1248);
or U7648 (N_7648,N_4435,N_3760);
or U7649 (N_7649,N_4344,N_4693);
and U7650 (N_7650,N_1473,N_4089);
nor U7651 (N_7651,N_502,N_40);
and U7652 (N_7652,N_3876,N_2912);
nand U7653 (N_7653,N_2069,N_3520);
nand U7654 (N_7654,N_3760,N_1972);
or U7655 (N_7655,N_2376,N_3713);
nor U7656 (N_7656,N_4608,N_783);
xnor U7657 (N_7657,N_2812,N_3770);
nor U7658 (N_7658,N_1562,N_4392);
and U7659 (N_7659,N_3674,N_2011);
nor U7660 (N_7660,N_4124,N_3603);
and U7661 (N_7661,N_3350,N_855);
nor U7662 (N_7662,N_2061,N_3713);
or U7663 (N_7663,N_2962,N_3019);
nor U7664 (N_7664,N_1332,N_1133);
nor U7665 (N_7665,N_51,N_2456);
nand U7666 (N_7666,N_3439,N_3031);
and U7667 (N_7667,N_4516,N_2906);
nor U7668 (N_7668,N_3626,N_3854);
nor U7669 (N_7669,N_3074,N_4064);
nand U7670 (N_7670,N_2596,N_381);
or U7671 (N_7671,N_4266,N_2281);
or U7672 (N_7672,N_452,N_2062);
nand U7673 (N_7673,N_4682,N_4076);
nand U7674 (N_7674,N_4014,N_4541);
xnor U7675 (N_7675,N_669,N_4950);
and U7676 (N_7676,N_2124,N_537);
xor U7677 (N_7677,N_3886,N_4387);
nor U7678 (N_7678,N_3634,N_4808);
nand U7679 (N_7679,N_3891,N_3336);
nand U7680 (N_7680,N_3524,N_1253);
xor U7681 (N_7681,N_1760,N_2706);
or U7682 (N_7682,N_4138,N_3276);
and U7683 (N_7683,N_3596,N_588);
xor U7684 (N_7684,N_3739,N_331);
or U7685 (N_7685,N_3358,N_3057);
xnor U7686 (N_7686,N_165,N_900);
nand U7687 (N_7687,N_2250,N_1026);
and U7688 (N_7688,N_3926,N_70);
and U7689 (N_7689,N_3472,N_3750);
and U7690 (N_7690,N_3375,N_3596);
and U7691 (N_7691,N_1722,N_3053);
nand U7692 (N_7692,N_1565,N_2672);
and U7693 (N_7693,N_515,N_4912);
xnor U7694 (N_7694,N_1356,N_4676);
or U7695 (N_7695,N_2395,N_190);
or U7696 (N_7696,N_4998,N_535);
and U7697 (N_7697,N_4975,N_1414);
or U7698 (N_7698,N_1789,N_4970);
nor U7699 (N_7699,N_2176,N_3034);
xor U7700 (N_7700,N_2960,N_2585);
nor U7701 (N_7701,N_4101,N_892);
or U7702 (N_7702,N_1778,N_1427);
and U7703 (N_7703,N_3952,N_2025);
xnor U7704 (N_7704,N_1002,N_1872);
or U7705 (N_7705,N_1245,N_4032);
and U7706 (N_7706,N_4681,N_2271);
or U7707 (N_7707,N_567,N_3536);
and U7708 (N_7708,N_4357,N_933);
and U7709 (N_7709,N_598,N_3993);
nor U7710 (N_7710,N_3632,N_1975);
xnor U7711 (N_7711,N_305,N_3709);
nor U7712 (N_7712,N_4561,N_4936);
nand U7713 (N_7713,N_2655,N_4954);
nand U7714 (N_7714,N_1043,N_952);
xor U7715 (N_7715,N_2400,N_3705);
nand U7716 (N_7716,N_1063,N_4831);
nor U7717 (N_7717,N_2603,N_1949);
or U7718 (N_7718,N_913,N_336);
nor U7719 (N_7719,N_4078,N_2280);
or U7720 (N_7720,N_887,N_3457);
nand U7721 (N_7721,N_3527,N_2377);
nor U7722 (N_7722,N_3788,N_124);
or U7723 (N_7723,N_936,N_2084);
nor U7724 (N_7724,N_3789,N_4202);
nand U7725 (N_7725,N_250,N_1544);
and U7726 (N_7726,N_3266,N_2318);
nor U7727 (N_7727,N_2711,N_1477);
or U7728 (N_7728,N_3723,N_3398);
or U7729 (N_7729,N_2687,N_715);
and U7730 (N_7730,N_3830,N_1285);
and U7731 (N_7731,N_1977,N_1076);
or U7732 (N_7732,N_532,N_1249);
nand U7733 (N_7733,N_2660,N_4251);
and U7734 (N_7734,N_2514,N_2902);
and U7735 (N_7735,N_1166,N_4603);
nor U7736 (N_7736,N_289,N_3904);
and U7737 (N_7737,N_2977,N_1483);
and U7738 (N_7738,N_4816,N_945);
and U7739 (N_7739,N_511,N_4217);
nand U7740 (N_7740,N_3246,N_1615);
nor U7741 (N_7741,N_4346,N_305);
nand U7742 (N_7742,N_3361,N_4366);
or U7743 (N_7743,N_1530,N_4649);
nand U7744 (N_7744,N_1652,N_1653);
nor U7745 (N_7745,N_3658,N_1447);
nand U7746 (N_7746,N_4399,N_3517);
and U7747 (N_7747,N_119,N_3488);
or U7748 (N_7748,N_4544,N_3150);
xnor U7749 (N_7749,N_2096,N_3789);
and U7750 (N_7750,N_3228,N_3604);
nor U7751 (N_7751,N_2814,N_691);
and U7752 (N_7752,N_1561,N_3298);
nor U7753 (N_7753,N_879,N_264);
nor U7754 (N_7754,N_2930,N_4427);
and U7755 (N_7755,N_2603,N_1983);
and U7756 (N_7756,N_120,N_4153);
nand U7757 (N_7757,N_1994,N_4285);
and U7758 (N_7758,N_374,N_4899);
xnor U7759 (N_7759,N_1036,N_103);
nand U7760 (N_7760,N_3905,N_1001);
nor U7761 (N_7761,N_4095,N_79);
or U7762 (N_7762,N_4846,N_3848);
nor U7763 (N_7763,N_179,N_3172);
or U7764 (N_7764,N_1187,N_2170);
nand U7765 (N_7765,N_1893,N_4440);
nor U7766 (N_7766,N_2401,N_2427);
xor U7767 (N_7767,N_975,N_606);
nor U7768 (N_7768,N_1059,N_1654);
and U7769 (N_7769,N_970,N_302);
nor U7770 (N_7770,N_984,N_3649);
or U7771 (N_7771,N_2696,N_676);
nor U7772 (N_7772,N_4243,N_4753);
xor U7773 (N_7773,N_816,N_3083);
and U7774 (N_7774,N_85,N_4556);
nand U7775 (N_7775,N_2877,N_3211);
nor U7776 (N_7776,N_3902,N_2386);
and U7777 (N_7777,N_3391,N_3658);
nand U7778 (N_7778,N_4222,N_1751);
nand U7779 (N_7779,N_1421,N_2723);
nor U7780 (N_7780,N_4701,N_2662);
xnor U7781 (N_7781,N_4894,N_2260);
and U7782 (N_7782,N_1943,N_730);
nand U7783 (N_7783,N_4803,N_1901);
nor U7784 (N_7784,N_2563,N_1751);
nor U7785 (N_7785,N_2202,N_4150);
and U7786 (N_7786,N_64,N_971);
nand U7787 (N_7787,N_3229,N_1677);
and U7788 (N_7788,N_1213,N_4455);
nor U7789 (N_7789,N_3713,N_4857);
and U7790 (N_7790,N_4252,N_4838);
and U7791 (N_7791,N_3344,N_3369);
and U7792 (N_7792,N_3524,N_4181);
and U7793 (N_7793,N_4693,N_4501);
nor U7794 (N_7794,N_2838,N_4989);
nor U7795 (N_7795,N_1343,N_2573);
or U7796 (N_7796,N_1179,N_3075);
nor U7797 (N_7797,N_4906,N_3647);
nand U7798 (N_7798,N_4411,N_106);
xnor U7799 (N_7799,N_4654,N_4115);
xnor U7800 (N_7800,N_1501,N_99);
nand U7801 (N_7801,N_3695,N_2520);
or U7802 (N_7802,N_2991,N_29);
and U7803 (N_7803,N_845,N_3118);
and U7804 (N_7804,N_1932,N_4912);
or U7805 (N_7805,N_2330,N_4601);
or U7806 (N_7806,N_4213,N_4830);
or U7807 (N_7807,N_3523,N_3296);
nor U7808 (N_7808,N_661,N_2075);
and U7809 (N_7809,N_952,N_2789);
xor U7810 (N_7810,N_3886,N_2920);
nand U7811 (N_7811,N_2701,N_4760);
or U7812 (N_7812,N_3788,N_1066);
nand U7813 (N_7813,N_1427,N_4653);
nand U7814 (N_7814,N_4286,N_4900);
nor U7815 (N_7815,N_4479,N_3690);
and U7816 (N_7816,N_4732,N_829);
and U7817 (N_7817,N_2171,N_3489);
xor U7818 (N_7818,N_3078,N_2808);
nand U7819 (N_7819,N_4021,N_1806);
or U7820 (N_7820,N_2989,N_573);
nor U7821 (N_7821,N_3635,N_2057);
or U7822 (N_7822,N_2645,N_2178);
xnor U7823 (N_7823,N_2626,N_2050);
and U7824 (N_7824,N_1602,N_4451);
nor U7825 (N_7825,N_126,N_4506);
and U7826 (N_7826,N_734,N_402);
and U7827 (N_7827,N_4986,N_3827);
nor U7828 (N_7828,N_692,N_636);
and U7829 (N_7829,N_4382,N_4761);
nor U7830 (N_7830,N_4461,N_4371);
nor U7831 (N_7831,N_4605,N_893);
nand U7832 (N_7832,N_4323,N_1469);
nand U7833 (N_7833,N_3014,N_2763);
or U7834 (N_7834,N_4713,N_3459);
or U7835 (N_7835,N_2260,N_4271);
nor U7836 (N_7836,N_1474,N_3783);
or U7837 (N_7837,N_218,N_909);
xnor U7838 (N_7838,N_3217,N_642);
xnor U7839 (N_7839,N_4225,N_4611);
nor U7840 (N_7840,N_1634,N_3551);
and U7841 (N_7841,N_3434,N_249);
xnor U7842 (N_7842,N_2521,N_4927);
nand U7843 (N_7843,N_1130,N_1324);
nor U7844 (N_7844,N_4048,N_2303);
or U7845 (N_7845,N_1194,N_344);
xor U7846 (N_7846,N_58,N_626);
nand U7847 (N_7847,N_2250,N_3757);
nand U7848 (N_7848,N_2712,N_705);
nand U7849 (N_7849,N_1372,N_529);
nor U7850 (N_7850,N_4449,N_1095);
xnor U7851 (N_7851,N_2449,N_2713);
or U7852 (N_7852,N_1998,N_609);
or U7853 (N_7853,N_1190,N_1033);
and U7854 (N_7854,N_1393,N_4177);
or U7855 (N_7855,N_1908,N_818);
or U7856 (N_7856,N_277,N_4415);
xor U7857 (N_7857,N_2904,N_3489);
nor U7858 (N_7858,N_4972,N_2499);
or U7859 (N_7859,N_1875,N_2147);
nor U7860 (N_7860,N_2026,N_2196);
or U7861 (N_7861,N_912,N_2580);
and U7862 (N_7862,N_1370,N_1540);
nand U7863 (N_7863,N_4845,N_2224);
nand U7864 (N_7864,N_4443,N_353);
and U7865 (N_7865,N_489,N_3304);
nor U7866 (N_7866,N_4291,N_2303);
nand U7867 (N_7867,N_4017,N_10);
or U7868 (N_7868,N_3857,N_4424);
or U7869 (N_7869,N_622,N_2666);
xnor U7870 (N_7870,N_582,N_2150);
nor U7871 (N_7871,N_1038,N_3409);
nor U7872 (N_7872,N_1652,N_601);
and U7873 (N_7873,N_2548,N_4619);
nand U7874 (N_7874,N_3276,N_3365);
nand U7875 (N_7875,N_3012,N_3257);
and U7876 (N_7876,N_1883,N_3356);
and U7877 (N_7877,N_3468,N_939);
or U7878 (N_7878,N_3947,N_1134);
or U7879 (N_7879,N_755,N_4895);
nor U7880 (N_7880,N_204,N_2187);
nand U7881 (N_7881,N_3906,N_2328);
nor U7882 (N_7882,N_1844,N_1728);
and U7883 (N_7883,N_2125,N_4550);
nand U7884 (N_7884,N_4243,N_1490);
nor U7885 (N_7885,N_3707,N_2635);
nor U7886 (N_7886,N_4426,N_2945);
xnor U7887 (N_7887,N_2037,N_2656);
nor U7888 (N_7888,N_4879,N_656);
and U7889 (N_7889,N_3653,N_1265);
xnor U7890 (N_7890,N_2589,N_1907);
nor U7891 (N_7891,N_3737,N_2841);
or U7892 (N_7892,N_4552,N_3452);
and U7893 (N_7893,N_4857,N_2689);
and U7894 (N_7894,N_2279,N_1855);
nor U7895 (N_7895,N_1571,N_913);
or U7896 (N_7896,N_691,N_2957);
nor U7897 (N_7897,N_4911,N_387);
and U7898 (N_7898,N_2194,N_1953);
nor U7899 (N_7899,N_644,N_4909);
nand U7900 (N_7900,N_4300,N_4730);
nor U7901 (N_7901,N_4796,N_3269);
xor U7902 (N_7902,N_4335,N_4388);
or U7903 (N_7903,N_2760,N_412);
nand U7904 (N_7904,N_1258,N_873);
or U7905 (N_7905,N_2122,N_4586);
or U7906 (N_7906,N_388,N_2619);
and U7907 (N_7907,N_1549,N_4144);
and U7908 (N_7908,N_3805,N_547);
or U7909 (N_7909,N_2051,N_3698);
or U7910 (N_7910,N_2895,N_2185);
xnor U7911 (N_7911,N_3272,N_410);
nand U7912 (N_7912,N_2833,N_1723);
nor U7913 (N_7913,N_504,N_4184);
nand U7914 (N_7914,N_3451,N_4109);
nor U7915 (N_7915,N_71,N_1096);
nor U7916 (N_7916,N_628,N_4467);
and U7917 (N_7917,N_3726,N_4905);
nand U7918 (N_7918,N_2521,N_535);
or U7919 (N_7919,N_4605,N_4876);
and U7920 (N_7920,N_1575,N_3890);
nand U7921 (N_7921,N_1918,N_4388);
xnor U7922 (N_7922,N_2969,N_4618);
nand U7923 (N_7923,N_4429,N_1625);
nor U7924 (N_7924,N_172,N_1880);
nand U7925 (N_7925,N_1442,N_2887);
xor U7926 (N_7926,N_3102,N_3438);
or U7927 (N_7927,N_1550,N_4504);
nand U7928 (N_7928,N_4687,N_180);
nor U7929 (N_7929,N_666,N_3331);
nor U7930 (N_7930,N_1312,N_2033);
or U7931 (N_7931,N_4537,N_214);
nand U7932 (N_7932,N_3714,N_877);
nand U7933 (N_7933,N_560,N_2182);
or U7934 (N_7934,N_2496,N_3611);
xnor U7935 (N_7935,N_2808,N_4838);
and U7936 (N_7936,N_3116,N_1113);
and U7937 (N_7937,N_3885,N_903);
or U7938 (N_7938,N_4812,N_1057);
and U7939 (N_7939,N_315,N_3476);
nor U7940 (N_7940,N_3204,N_2524);
nand U7941 (N_7941,N_2902,N_372);
nand U7942 (N_7942,N_3401,N_3573);
nor U7943 (N_7943,N_4719,N_312);
or U7944 (N_7944,N_4835,N_242);
nand U7945 (N_7945,N_2337,N_2033);
or U7946 (N_7946,N_3921,N_361);
nor U7947 (N_7947,N_3709,N_2473);
nor U7948 (N_7948,N_905,N_1192);
and U7949 (N_7949,N_3920,N_1639);
and U7950 (N_7950,N_4427,N_2047);
or U7951 (N_7951,N_495,N_4339);
nand U7952 (N_7952,N_1259,N_2344);
and U7953 (N_7953,N_3882,N_327);
or U7954 (N_7954,N_1850,N_1000);
nand U7955 (N_7955,N_3393,N_1816);
and U7956 (N_7956,N_4769,N_1750);
or U7957 (N_7957,N_4882,N_4249);
or U7958 (N_7958,N_3484,N_762);
nor U7959 (N_7959,N_4406,N_2990);
or U7960 (N_7960,N_4541,N_4103);
or U7961 (N_7961,N_392,N_2408);
nand U7962 (N_7962,N_13,N_582);
and U7963 (N_7963,N_3987,N_2775);
nor U7964 (N_7964,N_4873,N_3702);
nand U7965 (N_7965,N_644,N_611);
or U7966 (N_7966,N_4974,N_1248);
and U7967 (N_7967,N_831,N_3287);
nand U7968 (N_7968,N_3720,N_373);
nand U7969 (N_7969,N_2140,N_1582);
and U7970 (N_7970,N_3875,N_1796);
and U7971 (N_7971,N_1789,N_3841);
or U7972 (N_7972,N_2114,N_3991);
nand U7973 (N_7973,N_796,N_249);
nor U7974 (N_7974,N_2963,N_4131);
and U7975 (N_7975,N_2056,N_965);
nand U7976 (N_7976,N_1693,N_4477);
or U7977 (N_7977,N_3036,N_1829);
or U7978 (N_7978,N_4572,N_2928);
nand U7979 (N_7979,N_3319,N_3125);
nand U7980 (N_7980,N_3301,N_2137);
nor U7981 (N_7981,N_2455,N_3004);
and U7982 (N_7982,N_101,N_1753);
and U7983 (N_7983,N_3897,N_4520);
xor U7984 (N_7984,N_4054,N_3092);
and U7985 (N_7985,N_1180,N_1707);
and U7986 (N_7986,N_4850,N_948);
nand U7987 (N_7987,N_4544,N_4474);
nor U7988 (N_7988,N_3832,N_4868);
nand U7989 (N_7989,N_331,N_2457);
nor U7990 (N_7990,N_463,N_4197);
nand U7991 (N_7991,N_2368,N_2642);
nor U7992 (N_7992,N_507,N_3432);
nand U7993 (N_7993,N_1244,N_1860);
nor U7994 (N_7994,N_3915,N_2702);
and U7995 (N_7995,N_2021,N_2946);
xor U7996 (N_7996,N_1928,N_2308);
and U7997 (N_7997,N_2126,N_2388);
nand U7998 (N_7998,N_3636,N_3362);
xor U7999 (N_7999,N_1622,N_3681);
xnor U8000 (N_8000,N_2617,N_1867);
nor U8001 (N_8001,N_32,N_4201);
xor U8002 (N_8002,N_4665,N_4442);
nand U8003 (N_8003,N_551,N_4658);
nor U8004 (N_8004,N_4886,N_3837);
nand U8005 (N_8005,N_2816,N_4947);
or U8006 (N_8006,N_4839,N_3198);
or U8007 (N_8007,N_3269,N_2227);
and U8008 (N_8008,N_4412,N_4806);
xor U8009 (N_8009,N_2020,N_2102);
nor U8010 (N_8010,N_3520,N_3398);
and U8011 (N_8011,N_3138,N_2839);
nand U8012 (N_8012,N_3432,N_1875);
nand U8013 (N_8013,N_3627,N_3028);
nand U8014 (N_8014,N_4565,N_2861);
nand U8015 (N_8015,N_2861,N_3736);
nand U8016 (N_8016,N_47,N_738);
nor U8017 (N_8017,N_1554,N_293);
nor U8018 (N_8018,N_4309,N_2701);
xor U8019 (N_8019,N_3380,N_1812);
or U8020 (N_8020,N_844,N_1182);
or U8021 (N_8021,N_3226,N_694);
nand U8022 (N_8022,N_1063,N_650);
nand U8023 (N_8023,N_4340,N_328);
nor U8024 (N_8024,N_236,N_2137);
nand U8025 (N_8025,N_4191,N_456);
xnor U8026 (N_8026,N_688,N_3552);
nor U8027 (N_8027,N_1469,N_1109);
xor U8028 (N_8028,N_2444,N_3425);
and U8029 (N_8029,N_4064,N_4462);
and U8030 (N_8030,N_848,N_397);
or U8031 (N_8031,N_2689,N_2150);
or U8032 (N_8032,N_451,N_2264);
or U8033 (N_8033,N_2620,N_77);
and U8034 (N_8034,N_4962,N_2555);
or U8035 (N_8035,N_4734,N_867);
nand U8036 (N_8036,N_389,N_4241);
xor U8037 (N_8037,N_1042,N_4291);
nand U8038 (N_8038,N_2689,N_2619);
xnor U8039 (N_8039,N_487,N_2261);
nor U8040 (N_8040,N_348,N_626);
nand U8041 (N_8041,N_3311,N_1269);
and U8042 (N_8042,N_2115,N_2139);
nand U8043 (N_8043,N_4757,N_2306);
or U8044 (N_8044,N_3557,N_566);
nand U8045 (N_8045,N_4660,N_4124);
and U8046 (N_8046,N_2001,N_3368);
nand U8047 (N_8047,N_2845,N_912);
nor U8048 (N_8048,N_2904,N_147);
nor U8049 (N_8049,N_3910,N_237);
nor U8050 (N_8050,N_3217,N_2766);
nand U8051 (N_8051,N_2399,N_3320);
or U8052 (N_8052,N_135,N_1543);
or U8053 (N_8053,N_1491,N_796);
nand U8054 (N_8054,N_1091,N_2906);
nor U8055 (N_8055,N_4397,N_1455);
nand U8056 (N_8056,N_2608,N_2616);
nor U8057 (N_8057,N_2999,N_555);
or U8058 (N_8058,N_2121,N_878);
and U8059 (N_8059,N_2861,N_2091);
nor U8060 (N_8060,N_2765,N_3124);
or U8061 (N_8061,N_4939,N_2191);
or U8062 (N_8062,N_56,N_2474);
nor U8063 (N_8063,N_1702,N_512);
or U8064 (N_8064,N_2380,N_1044);
and U8065 (N_8065,N_114,N_2433);
and U8066 (N_8066,N_196,N_1352);
and U8067 (N_8067,N_2725,N_4685);
nor U8068 (N_8068,N_358,N_2668);
nand U8069 (N_8069,N_1760,N_4848);
or U8070 (N_8070,N_3755,N_21);
nand U8071 (N_8071,N_771,N_2128);
or U8072 (N_8072,N_1167,N_2690);
or U8073 (N_8073,N_1028,N_1026);
nand U8074 (N_8074,N_990,N_4668);
or U8075 (N_8075,N_1541,N_4626);
and U8076 (N_8076,N_3003,N_937);
nor U8077 (N_8077,N_2862,N_3852);
nor U8078 (N_8078,N_1794,N_4894);
nor U8079 (N_8079,N_674,N_3096);
and U8080 (N_8080,N_1731,N_1649);
nor U8081 (N_8081,N_3034,N_1129);
and U8082 (N_8082,N_3159,N_2635);
nand U8083 (N_8083,N_2599,N_810);
nand U8084 (N_8084,N_1515,N_3305);
nor U8085 (N_8085,N_101,N_1088);
and U8086 (N_8086,N_3666,N_4432);
nor U8087 (N_8087,N_3853,N_2041);
nand U8088 (N_8088,N_874,N_3869);
and U8089 (N_8089,N_3585,N_709);
or U8090 (N_8090,N_4101,N_2970);
nand U8091 (N_8091,N_2349,N_1502);
and U8092 (N_8092,N_3536,N_4904);
xor U8093 (N_8093,N_3003,N_4242);
xor U8094 (N_8094,N_2388,N_4058);
xor U8095 (N_8095,N_1976,N_2982);
and U8096 (N_8096,N_3195,N_4110);
nand U8097 (N_8097,N_4828,N_3707);
nand U8098 (N_8098,N_2786,N_561);
or U8099 (N_8099,N_4407,N_2119);
nand U8100 (N_8100,N_3518,N_4540);
nor U8101 (N_8101,N_2438,N_2432);
nand U8102 (N_8102,N_4960,N_1832);
or U8103 (N_8103,N_4694,N_1306);
nand U8104 (N_8104,N_3443,N_4033);
or U8105 (N_8105,N_1696,N_3048);
or U8106 (N_8106,N_4134,N_320);
and U8107 (N_8107,N_4120,N_1);
nor U8108 (N_8108,N_4400,N_1888);
nand U8109 (N_8109,N_2522,N_959);
nand U8110 (N_8110,N_1151,N_2771);
and U8111 (N_8111,N_4022,N_605);
and U8112 (N_8112,N_4055,N_4960);
nor U8113 (N_8113,N_1224,N_2633);
xor U8114 (N_8114,N_961,N_1775);
nand U8115 (N_8115,N_1565,N_398);
and U8116 (N_8116,N_2256,N_1126);
nand U8117 (N_8117,N_2174,N_678);
nand U8118 (N_8118,N_1117,N_4178);
nor U8119 (N_8119,N_2729,N_2078);
or U8120 (N_8120,N_676,N_4698);
nand U8121 (N_8121,N_3316,N_4209);
nand U8122 (N_8122,N_2570,N_4318);
nor U8123 (N_8123,N_2898,N_2180);
or U8124 (N_8124,N_862,N_4139);
nor U8125 (N_8125,N_3684,N_2781);
nor U8126 (N_8126,N_3832,N_1034);
and U8127 (N_8127,N_3923,N_4365);
nand U8128 (N_8128,N_572,N_537);
nand U8129 (N_8129,N_1087,N_374);
or U8130 (N_8130,N_1682,N_3930);
nor U8131 (N_8131,N_1952,N_60);
or U8132 (N_8132,N_2565,N_3527);
or U8133 (N_8133,N_1176,N_1338);
nand U8134 (N_8134,N_2927,N_4459);
and U8135 (N_8135,N_4926,N_2665);
xor U8136 (N_8136,N_985,N_3246);
or U8137 (N_8137,N_3263,N_4484);
and U8138 (N_8138,N_2070,N_3244);
nand U8139 (N_8139,N_4755,N_364);
and U8140 (N_8140,N_168,N_572);
nand U8141 (N_8141,N_3865,N_1833);
nand U8142 (N_8142,N_2053,N_2536);
nor U8143 (N_8143,N_3471,N_4485);
nand U8144 (N_8144,N_4683,N_1154);
xor U8145 (N_8145,N_3290,N_1106);
and U8146 (N_8146,N_4172,N_1201);
or U8147 (N_8147,N_2208,N_3846);
nor U8148 (N_8148,N_2807,N_3223);
nand U8149 (N_8149,N_1624,N_3587);
xor U8150 (N_8150,N_2190,N_2837);
nand U8151 (N_8151,N_136,N_291);
and U8152 (N_8152,N_2837,N_973);
xnor U8153 (N_8153,N_767,N_2415);
or U8154 (N_8154,N_3790,N_1102);
and U8155 (N_8155,N_3126,N_904);
nand U8156 (N_8156,N_3494,N_764);
and U8157 (N_8157,N_4849,N_621);
nand U8158 (N_8158,N_744,N_4421);
or U8159 (N_8159,N_3877,N_2667);
and U8160 (N_8160,N_3178,N_1357);
or U8161 (N_8161,N_2632,N_3990);
or U8162 (N_8162,N_3728,N_951);
nor U8163 (N_8163,N_1873,N_4187);
or U8164 (N_8164,N_3881,N_4943);
nand U8165 (N_8165,N_4273,N_1382);
and U8166 (N_8166,N_3158,N_1517);
and U8167 (N_8167,N_4092,N_836);
nor U8168 (N_8168,N_1589,N_4204);
nor U8169 (N_8169,N_4112,N_1314);
or U8170 (N_8170,N_502,N_1400);
and U8171 (N_8171,N_3623,N_3519);
nor U8172 (N_8172,N_252,N_2396);
or U8173 (N_8173,N_3570,N_292);
or U8174 (N_8174,N_4230,N_598);
xor U8175 (N_8175,N_3056,N_4849);
or U8176 (N_8176,N_398,N_2413);
nor U8177 (N_8177,N_2299,N_2507);
nand U8178 (N_8178,N_3695,N_2453);
and U8179 (N_8179,N_1675,N_4529);
or U8180 (N_8180,N_2203,N_56);
or U8181 (N_8181,N_4072,N_329);
and U8182 (N_8182,N_1895,N_2235);
nand U8183 (N_8183,N_2049,N_3469);
nand U8184 (N_8184,N_3212,N_1808);
nor U8185 (N_8185,N_13,N_1518);
or U8186 (N_8186,N_2711,N_3027);
or U8187 (N_8187,N_4019,N_3191);
or U8188 (N_8188,N_4684,N_4723);
nand U8189 (N_8189,N_4403,N_244);
and U8190 (N_8190,N_1625,N_630);
nand U8191 (N_8191,N_1004,N_2760);
or U8192 (N_8192,N_2553,N_2379);
nand U8193 (N_8193,N_2517,N_758);
and U8194 (N_8194,N_769,N_2096);
and U8195 (N_8195,N_3879,N_4306);
or U8196 (N_8196,N_4783,N_723);
nand U8197 (N_8197,N_4807,N_1516);
nor U8198 (N_8198,N_2487,N_1379);
xor U8199 (N_8199,N_1423,N_3446);
nor U8200 (N_8200,N_1838,N_2732);
nor U8201 (N_8201,N_1560,N_707);
nand U8202 (N_8202,N_4210,N_4507);
or U8203 (N_8203,N_3091,N_625);
nor U8204 (N_8204,N_2075,N_189);
nor U8205 (N_8205,N_297,N_533);
nor U8206 (N_8206,N_1632,N_4614);
nand U8207 (N_8207,N_1644,N_134);
nand U8208 (N_8208,N_1135,N_689);
or U8209 (N_8209,N_4510,N_2925);
nand U8210 (N_8210,N_2939,N_273);
or U8211 (N_8211,N_1113,N_1736);
xnor U8212 (N_8212,N_1995,N_875);
and U8213 (N_8213,N_4693,N_1495);
xnor U8214 (N_8214,N_932,N_594);
xor U8215 (N_8215,N_4061,N_4808);
and U8216 (N_8216,N_3823,N_1392);
nand U8217 (N_8217,N_3120,N_4141);
nor U8218 (N_8218,N_1387,N_1041);
nand U8219 (N_8219,N_1279,N_523);
or U8220 (N_8220,N_4310,N_664);
xnor U8221 (N_8221,N_3584,N_265);
and U8222 (N_8222,N_3101,N_2590);
nand U8223 (N_8223,N_3665,N_3453);
or U8224 (N_8224,N_1034,N_835);
and U8225 (N_8225,N_3159,N_2920);
nand U8226 (N_8226,N_2786,N_4235);
or U8227 (N_8227,N_1089,N_2646);
nor U8228 (N_8228,N_2574,N_295);
nand U8229 (N_8229,N_918,N_2072);
xnor U8230 (N_8230,N_4222,N_3738);
and U8231 (N_8231,N_2362,N_3213);
xor U8232 (N_8232,N_1408,N_4912);
nor U8233 (N_8233,N_182,N_3373);
nand U8234 (N_8234,N_1157,N_23);
or U8235 (N_8235,N_1883,N_116);
nor U8236 (N_8236,N_87,N_67);
nand U8237 (N_8237,N_3000,N_2805);
or U8238 (N_8238,N_4887,N_3332);
or U8239 (N_8239,N_3564,N_306);
and U8240 (N_8240,N_2111,N_2016);
or U8241 (N_8241,N_96,N_2599);
or U8242 (N_8242,N_1390,N_3743);
or U8243 (N_8243,N_2855,N_3649);
and U8244 (N_8244,N_2023,N_3633);
and U8245 (N_8245,N_4594,N_3358);
nand U8246 (N_8246,N_2364,N_1373);
nor U8247 (N_8247,N_716,N_2997);
nand U8248 (N_8248,N_179,N_4100);
and U8249 (N_8249,N_932,N_1584);
and U8250 (N_8250,N_674,N_1411);
xor U8251 (N_8251,N_354,N_2649);
nand U8252 (N_8252,N_4073,N_1647);
nand U8253 (N_8253,N_2321,N_877);
xor U8254 (N_8254,N_4259,N_2550);
nor U8255 (N_8255,N_3319,N_4058);
nand U8256 (N_8256,N_3951,N_3701);
nor U8257 (N_8257,N_3131,N_4919);
nor U8258 (N_8258,N_1018,N_3621);
nor U8259 (N_8259,N_3806,N_456);
nor U8260 (N_8260,N_4783,N_4897);
nand U8261 (N_8261,N_943,N_3734);
xnor U8262 (N_8262,N_2688,N_2665);
nand U8263 (N_8263,N_944,N_263);
or U8264 (N_8264,N_513,N_3822);
nor U8265 (N_8265,N_1178,N_2026);
nand U8266 (N_8266,N_4560,N_4527);
nand U8267 (N_8267,N_2943,N_2168);
nor U8268 (N_8268,N_1978,N_3885);
nand U8269 (N_8269,N_4597,N_3330);
nor U8270 (N_8270,N_1049,N_4444);
and U8271 (N_8271,N_259,N_2544);
nor U8272 (N_8272,N_784,N_1651);
nand U8273 (N_8273,N_556,N_765);
nand U8274 (N_8274,N_73,N_3329);
and U8275 (N_8275,N_2685,N_4625);
nand U8276 (N_8276,N_3513,N_1437);
nand U8277 (N_8277,N_905,N_4621);
or U8278 (N_8278,N_4873,N_315);
nand U8279 (N_8279,N_679,N_1040);
nand U8280 (N_8280,N_2088,N_3763);
nand U8281 (N_8281,N_339,N_3454);
or U8282 (N_8282,N_4118,N_4111);
and U8283 (N_8283,N_3290,N_3254);
xor U8284 (N_8284,N_3091,N_261);
nor U8285 (N_8285,N_1336,N_4241);
nand U8286 (N_8286,N_3907,N_2359);
and U8287 (N_8287,N_3089,N_3206);
or U8288 (N_8288,N_3878,N_4345);
and U8289 (N_8289,N_3128,N_988);
or U8290 (N_8290,N_4564,N_2502);
and U8291 (N_8291,N_1709,N_3042);
nor U8292 (N_8292,N_2835,N_4184);
and U8293 (N_8293,N_944,N_336);
xor U8294 (N_8294,N_412,N_4147);
nor U8295 (N_8295,N_4463,N_2203);
or U8296 (N_8296,N_1364,N_3558);
xnor U8297 (N_8297,N_3012,N_2515);
nand U8298 (N_8298,N_3470,N_3133);
nand U8299 (N_8299,N_2529,N_1705);
and U8300 (N_8300,N_2036,N_3679);
or U8301 (N_8301,N_3556,N_130);
nor U8302 (N_8302,N_494,N_2832);
xnor U8303 (N_8303,N_900,N_4521);
nor U8304 (N_8304,N_644,N_1117);
and U8305 (N_8305,N_4850,N_3735);
or U8306 (N_8306,N_2721,N_3066);
or U8307 (N_8307,N_1157,N_1615);
or U8308 (N_8308,N_3643,N_1274);
nor U8309 (N_8309,N_2397,N_4651);
and U8310 (N_8310,N_4268,N_2587);
xor U8311 (N_8311,N_4829,N_2813);
xnor U8312 (N_8312,N_1929,N_151);
nand U8313 (N_8313,N_2437,N_3950);
and U8314 (N_8314,N_853,N_178);
or U8315 (N_8315,N_834,N_213);
nand U8316 (N_8316,N_2947,N_2225);
nor U8317 (N_8317,N_4784,N_3060);
nor U8318 (N_8318,N_3003,N_1588);
or U8319 (N_8319,N_1927,N_24);
nand U8320 (N_8320,N_3724,N_1019);
nor U8321 (N_8321,N_159,N_1301);
or U8322 (N_8322,N_1041,N_117);
or U8323 (N_8323,N_2668,N_668);
or U8324 (N_8324,N_4365,N_1570);
nor U8325 (N_8325,N_2192,N_466);
or U8326 (N_8326,N_1877,N_2438);
or U8327 (N_8327,N_4748,N_2154);
xnor U8328 (N_8328,N_2253,N_2483);
nor U8329 (N_8329,N_1466,N_4949);
or U8330 (N_8330,N_792,N_3991);
nand U8331 (N_8331,N_4429,N_2318);
nor U8332 (N_8332,N_1692,N_3381);
nand U8333 (N_8333,N_4908,N_2756);
nor U8334 (N_8334,N_2309,N_3097);
or U8335 (N_8335,N_3768,N_1581);
or U8336 (N_8336,N_2137,N_2245);
and U8337 (N_8337,N_961,N_122);
and U8338 (N_8338,N_3789,N_221);
and U8339 (N_8339,N_2955,N_2160);
or U8340 (N_8340,N_651,N_4751);
and U8341 (N_8341,N_3889,N_2537);
nor U8342 (N_8342,N_3790,N_3854);
or U8343 (N_8343,N_4637,N_4404);
nor U8344 (N_8344,N_3598,N_559);
nor U8345 (N_8345,N_4376,N_2538);
nand U8346 (N_8346,N_4752,N_288);
nand U8347 (N_8347,N_3337,N_4905);
nand U8348 (N_8348,N_2553,N_3967);
xor U8349 (N_8349,N_2145,N_2976);
nor U8350 (N_8350,N_3882,N_2425);
and U8351 (N_8351,N_3310,N_1979);
nor U8352 (N_8352,N_473,N_4657);
and U8353 (N_8353,N_1359,N_1157);
or U8354 (N_8354,N_4473,N_4174);
or U8355 (N_8355,N_4791,N_4102);
or U8356 (N_8356,N_1590,N_747);
nor U8357 (N_8357,N_57,N_3770);
and U8358 (N_8358,N_16,N_4180);
nor U8359 (N_8359,N_3268,N_2924);
or U8360 (N_8360,N_1892,N_3204);
and U8361 (N_8361,N_3102,N_3339);
and U8362 (N_8362,N_2252,N_79);
and U8363 (N_8363,N_4106,N_3040);
and U8364 (N_8364,N_2410,N_2025);
nand U8365 (N_8365,N_2044,N_1135);
nand U8366 (N_8366,N_4280,N_2334);
nor U8367 (N_8367,N_2006,N_3499);
or U8368 (N_8368,N_778,N_649);
or U8369 (N_8369,N_4189,N_2946);
and U8370 (N_8370,N_1077,N_250);
nor U8371 (N_8371,N_249,N_2298);
nor U8372 (N_8372,N_754,N_1624);
nand U8373 (N_8373,N_2932,N_3075);
xnor U8374 (N_8374,N_2079,N_3065);
nand U8375 (N_8375,N_1037,N_153);
or U8376 (N_8376,N_3256,N_3640);
and U8377 (N_8377,N_3394,N_93);
or U8378 (N_8378,N_3086,N_4117);
nor U8379 (N_8379,N_4305,N_1038);
nor U8380 (N_8380,N_2009,N_502);
xnor U8381 (N_8381,N_1317,N_2291);
or U8382 (N_8382,N_2837,N_2477);
xor U8383 (N_8383,N_93,N_2231);
and U8384 (N_8384,N_28,N_3972);
nand U8385 (N_8385,N_4747,N_947);
nand U8386 (N_8386,N_1561,N_4456);
xor U8387 (N_8387,N_4228,N_867);
or U8388 (N_8388,N_2385,N_2908);
xnor U8389 (N_8389,N_2553,N_2565);
nor U8390 (N_8390,N_1692,N_163);
nor U8391 (N_8391,N_1401,N_2577);
xor U8392 (N_8392,N_749,N_4699);
or U8393 (N_8393,N_3401,N_13);
nor U8394 (N_8394,N_943,N_1375);
nand U8395 (N_8395,N_4740,N_4104);
or U8396 (N_8396,N_2595,N_4519);
or U8397 (N_8397,N_4302,N_318);
and U8398 (N_8398,N_3637,N_810);
nor U8399 (N_8399,N_2454,N_3833);
nor U8400 (N_8400,N_1305,N_2287);
or U8401 (N_8401,N_4356,N_1241);
and U8402 (N_8402,N_3628,N_2606);
nand U8403 (N_8403,N_163,N_4044);
nor U8404 (N_8404,N_1952,N_4709);
nor U8405 (N_8405,N_3212,N_2189);
and U8406 (N_8406,N_1728,N_805);
nand U8407 (N_8407,N_2952,N_2280);
xnor U8408 (N_8408,N_1863,N_4763);
and U8409 (N_8409,N_2920,N_4521);
nand U8410 (N_8410,N_3994,N_701);
and U8411 (N_8411,N_269,N_4000);
nor U8412 (N_8412,N_163,N_3951);
nand U8413 (N_8413,N_598,N_4138);
nor U8414 (N_8414,N_1963,N_650);
or U8415 (N_8415,N_3048,N_2981);
or U8416 (N_8416,N_1708,N_1301);
or U8417 (N_8417,N_2738,N_1451);
nand U8418 (N_8418,N_4217,N_586);
and U8419 (N_8419,N_57,N_517);
nand U8420 (N_8420,N_1246,N_1577);
or U8421 (N_8421,N_1758,N_4033);
nor U8422 (N_8422,N_1618,N_1596);
or U8423 (N_8423,N_1102,N_210);
or U8424 (N_8424,N_3235,N_4942);
xnor U8425 (N_8425,N_4096,N_928);
nor U8426 (N_8426,N_4988,N_1558);
nor U8427 (N_8427,N_1636,N_1739);
and U8428 (N_8428,N_2718,N_3306);
nor U8429 (N_8429,N_1497,N_818);
or U8430 (N_8430,N_288,N_2627);
nand U8431 (N_8431,N_4175,N_3195);
or U8432 (N_8432,N_2982,N_3441);
nand U8433 (N_8433,N_241,N_1658);
nand U8434 (N_8434,N_2800,N_695);
nor U8435 (N_8435,N_4325,N_2240);
xnor U8436 (N_8436,N_1734,N_2490);
or U8437 (N_8437,N_4973,N_3579);
nor U8438 (N_8438,N_2124,N_2255);
or U8439 (N_8439,N_3765,N_728);
nand U8440 (N_8440,N_4481,N_1138);
and U8441 (N_8441,N_4169,N_1823);
nor U8442 (N_8442,N_1298,N_2519);
nand U8443 (N_8443,N_2289,N_1721);
and U8444 (N_8444,N_3180,N_4109);
or U8445 (N_8445,N_3744,N_3701);
xor U8446 (N_8446,N_1101,N_2949);
and U8447 (N_8447,N_1374,N_1598);
and U8448 (N_8448,N_3135,N_3885);
nand U8449 (N_8449,N_4862,N_2677);
or U8450 (N_8450,N_2182,N_4042);
xnor U8451 (N_8451,N_2888,N_382);
or U8452 (N_8452,N_4360,N_477);
and U8453 (N_8453,N_1348,N_3252);
or U8454 (N_8454,N_3513,N_3544);
nand U8455 (N_8455,N_3001,N_2760);
nor U8456 (N_8456,N_667,N_2957);
or U8457 (N_8457,N_310,N_4571);
xnor U8458 (N_8458,N_2788,N_4518);
nor U8459 (N_8459,N_2944,N_4067);
and U8460 (N_8460,N_2149,N_4384);
and U8461 (N_8461,N_2819,N_1438);
or U8462 (N_8462,N_1051,N_4361);
nand U8463 (N_8463,N_1255,N_35);
or U8464 (N_8464,N_1125,N_1674);
nand U8465 (N_8465,N_2362,N_3401);
and U8466 (N_8466,N_86,N_3833);
nor U8467 (N_8467,N_1692,N_1357);
or U8468 (N_8468,N_3945,N_3177);
or U8469 (N_8469,N_3985,N_3329);
xnor U8470 (N_8470,N_3614,N_2047);
nand U8471 (N_8471,N_1936,N_3522);
or U8472 (N_8472,N_4128,N_732);
and U8473 (N_8473,N_2365,N_2413);
nand U8474 (N_8474,N_1719,N_1037);
and U8475 (N_8475,N_1015,N_1400);
or U8476 (N_8476,N_4225,N_4065);
and U8477 (N_8477,N_1570,N_1088);
or U8478 (N_8478,N_1919,N_2823);
or U8479 (N_8479,N_1049,N_2869);
or U8480 (N_8480,N_519,N_1971);
nor U8481 (N_8481,N_4525,N_697);
nor U8482 (N_8482,N_1342,N_4811);
xor U8483 (N_8483,N_83,N_2191);
and U8484 (N_8484,N_2228,N_356);
and U8485 (N_8485,N_4772,N_2360);
nor U8486 (N_8486,N_1411,N_1850);
nand U8487 (N_8487,N_4185,N_1360);
nor U8488 (N_8488,N_800,N_4270);
and U8489 (N_8489,N_3683,N_2680);
and U8490 (N_8490,N_3203,N_404);
or U8491 (N_8491,N_2839,N_2782);
nor U8492 (N_8492,N_3059,N_289);
nor U8493 (N_8493,N_4157,N_1683);
nand U8494 (N_8494,N_3913,N_3816);
and U8495 (N_8495,N_3676,N_776);
nor U8496 (N_8496,N_2918,N_3763);
nor U8497 (N_8497,N_1554,N_2512);
nand U8498 (N_8498,N_4200,N_1959);
nor U8499 (N_8499,N_3402,N_481);
or U8500 (N_8500,N_3813,N_3120);
and U8501 (N_8501,N_4587,N_2756);
xnor U8502 (N_8502,N_1202,N_3852);
and U8503 (N_8503,N_2590,N_3406);
nor U8504 (N_8504,N_285,N_453);
nor U8505 (N_8505,N_4362,N_3680);
and U8506 (N_8506,N_1480,N_1926);
or U8507 (N_8507,N_3799,N_405);
and U8508 (N_8508,N_2212,N_1006);
xor U8509 (N_8509,N_3456,N_2520);
nor U8510 (N_8510,N_2892,N_737);
and U8511 (N_8511,N_3212,N_162);
nor U8512 (N_8512,N_4462,N_1704);
or U8513 (N_8513,N_1948,N_3202);
nand U8514 (N_8514,N_4094,N_819);
and U8515 (N_8515,N_2034,N_468);
or U8516 (N_8516,N_3033,N_4129);
xor U8517 (N_8517,N_734,N_4586);
or U8518 (N_8518,N_1640,N_2345);
and U8519 (N_8519,N_1832,N_3319);
or U8520 (N_8520,N_343,N_924);
nor U8521 (N_8521,N_1924,N_1893);
nand U8522 (N_8522,N_3159,N_4232);
or U8523 (N_8523,N_3471,N_2854);
or U8524 (N_8524,N_152,N_1146);
nor U8525 (N_8525,N_2856,N_4723);
xnor U8526 (N_8526,N_4601,N_2789);
or U8527 (N_8527,N_633,N_2229);
and U8528 (N_8528,N_3137,N_4391);
or U8529 (N_8529,N_4719,N_2576);
nand U8530 (N_8530,N_3928,N_1798);
or U8531 (N_8531,N_4854,N_907);
and U8532 (N_8532,N_1002,N_2950);
nor U8533 (N_8533,N_1987,N_3615);
and U8534 (N_8534,N_3112,N_3106);
or U8535 (N_8535,N_460,N_4152);
and U8536 (N_8536,N_1420,N_2895);
nand U8537 (N_8537,N_591,N_3238);
or U8538 (N_8538,N_2733,N_1796);
nand U8539 (N_8539,N_4841,N_2329);
nand U8540 (N_8540,N_3457,N_2794);
xnor U8541 (N_8541,N_4596,N_2407);
nand U8542 (N_8542,N_607,N_1494);
nand U8543 (N_8543,N_1530,N_2473);
nand U8544 (N_8544,N_4652,N_2097);
xor U8545 (N_8545,N_446,N_1304);
or U8546 (N_8546,N_4518,N_176);
nor U8547 (N_8547,N_4092,N_3788);
or U8548 (N_8548,N_1067,N_4837);
nor U8549 (N_8549,N_4548,N_611);
and U8550 (N_8550,N_521,N_1284);
or U8551 (N_8551,N_3560,N_3838);
or U8552 (N_8552,N_123,N_3743);
nor U8553 (N_8553,N_2489,N_2765);
nand U8554 (N_8554,N_4037,N_2898);
xnor U8555 (N_8555,N_3817,N_457);
nor U8556 (N_8556,N_38,N_3457);
and U8557 (N_8557,N_3341,N_4197);
or U8558 (N_8558,N_4575,N_1723);
or U8559 (N_8559,N_4795,N_63);
nor U8560 (N_8560,N_1766,N_3209);
and U8561 (N_8561,N_1428,N_4700);
and U8562 (N_8562,N_2812,N_2648);
nand U8563 (N_8563,N_1036,N_4212);
nand U8564 (N_8564,N_3430,N_4630);
nand U8565 (N_8565,N_4832,N_3392);
nor U8566 (N_8566,N_2943,N_2550);
nor U8567 (N_8567,N_82,N_4514);
nand U8568 (N_8568,N_4226,N_4710);
or U8569 (N_8569,N_1805,N_4788);
xor U8570 (N_8570,N_2381,N_4493);
xnor U8571 (N_8571,N_2475,N_4805);
nor U8572 (N_8572,N_6,N_8);
nand U8573 (N_8573,N_4417,N_77);
xnor U8574 (N_8574,N_1428,N_4914);
or U8575 (N_8575,N_4730,N_3672);
xnor U8576 (N_8576,N_1793,N_228);
nand U8577 (N_8577,N_2807,N_4862);
and U8578 (N_8578,N_1289,N_2858);
nor U8579 (N_8579,N_2198,N_3352);
nor U8580 (N_8580,N_1609,N_1457);
nor U8581 (N_8581,N_4644,N_3697);
nor U8582 (N_8582,N_2200,N_36);
or U8583 (N_8583,N_165,N_1008);
or U8584 (N_8584,N_1568,N_837);
or U8585 (N_8585,N_2572,N_886);
or U8586 (N_8586,N_4417,N_1571);
or U8587 (N_8587,N_240,N_3574);
nand U8588 (N_8588,N_1039,N_3586);
nand U8589 (N_8589,N_193,N_4249);
nor U8590 (N_8590,N_1416,N_2497);
and U8591 (N_8591,N_4703,N_515);
nand U8592 (N_8592,N_3527,N_1383);
or U8593 (N_8593,N_3261,N_1990);
nor U8594 (N_8594,N_4339,N_2339);
or U8595 (N_8595,N_4512,N_311);
nor U8596 (N_8596,N_3607,N_4345);
nor U8597 (N_8597,N_2539,N_193);
nand U8598 (N_8598,N_13,N_78);
or U8599 (N_8599,N_38,N_2431);
nor U8600 (N_8600,N_1561,N_3858);
nor U8601 (N_8601,N_2993,N_1246);
nor U8602 (N_8602,N_4198,N_4430);
or U8603 (N_8603,N_4997,N_4725);
and U8604 (N_8604,N_2973,N_4378);
xnor U8605 (N_8605,N_801,N_4124);
nand U8606 (N_8606,N_2872,N_2446);
or U8607 (N_8607,N_133,N_3178);
and U8608 (N_8608,N_578,N_2982);
nor U8609 (N_8609,N_3654,N_4804);
xor U8610 (N_8610,N_1117,N_1849);
nand U8611 (N_8611,N_2563,N_3886);
nor U8612 (N_8612,N_104,N_2161);
nand U8613 (N_8613,N_1481,N_23);
nand U8614 (N_8614,N_1644,N_781);
xor U8615 (N_8615,N_1674,N_2005);
and U8616 (N_8616,N_708,N_2247);
xor U8617 (N_8617,N_4129,N_261);
and U8618 (N_8618,N_1409,N_3175);
nand U8619 (N_8619,N_4486,N_2919);
and U8620 (N_8620,N_4553,N_397);
and U8621 (N_8621,N_2692,N_2257);
nor U8622 (N_8622,N_2615,N_107);
and U8623 (N_8623,N_3539,N_2741);
and U8624 (N_8624,N_1549,N_4900);
or U8625 (N_8625,N_3284,N_3716);
or U8626 (N_8626,N_905,N_1584);
nor U8627 (N_8627,N_1861,N_3114);
nor U8628 (N_8628,N_1268,N_4507);
or U8629 (N_8629,N_4658,N_110);
and U8630 (N_8630,N_4267,N_2965);
nand U8631 (N_8631,N_2801,N_3146);
and U8632 (N_8632,N_4876,N_3503);
and U8633 (N_8633,N_1950,N_1666);
nor U8634 (N_8634,N_1045,N_850);
nor U8635 (N_8635,N_4693,N_3441);
nor U8636 (N_8636,N_4699,N_1208);
or U8637 (N_8637,N_4948,N_756);
xnor U8638 (N_8638,N_3413,N_3730);
and U8639 (N_8639,N_3925,N_3924);
and U8640 (N_8640,N_970,N_3923);
nor U8641 (N_8641,N_161,N_2465);
or U8642 (N_8642,N_2730,N_2335);
and U8643 (N_8643,N_4438,N_2397);
nand U8644 (N_8644,N_4872,N_1433);
and U8645 (N_8645,N_2482,N_4237);
xnor U8646 (N_8646,N_616,N_1953);
or U8647 (N_8647,N_4564,N_2203);
or U8648 (N_8648,N_4366,N_4078);
or U8649 (N_8649,N_3915,N_2989);
xor U8650 (N_8650,N_2989,N_4675);
nand U8651 (N_8651,N_2702,N_818);
and U8652 (N_8652,N_2002,N_674);
and U8653 (N_8653,N_3217,N_3810);
xor U8654 (N_8654,N_2028,N_1167);
and U8655 (N_8655,N_2945,N_1223);
nor U8656 (N_8656,N_2746,N_4586);
or U8657 (N_8657,N_4338,N_2259);
nor U8658 (N_8658,N_4012,N_841);
nor U8659 (N_8659,N_1854,N_2193);
nor U8660 (N_8660,N_2902,N_2254);
and U8661 (N_8661,N_3818,N_476);
and U8662 (N_8662,N_3366,N_840);
nand U8663 (N_8663,N_1441,N_2241);
nor U8664 (N_8664,N_743,N_4586);
or U8665 (N_8665,N_3996,N_2242);
or U8666 (N_8666,N_1876,N_3560);
or U8667 (N_8667,N_2385,N_3267);
nor U8668 (N_8668,N_1168,N_520);
or U8669 (N_8669,N_3015,N_2502);
nand U8670 (N_8670,N_3249,N_4460);
nand U8671 (N_8671,N_148,N_1413);
nand U8672 (N_8672,N_3037,N_362);
nor U8673 (N_8673,N_3858,N_978);
and U8674 (N_8674,N_4832,N_3499);
nor U8675 (N_8675,N_249,N_732);
nor U8676 (N_8676,N_4102,N_4365);
nor U8677 (N_8677,N_2287,N_2692);
or U8678 (N_8678,N_4416,N_596);
nand U8679 (N_8679,N_4590,N_1482);
nand U8680 (N_8680,N_3558,N_1382);
xnor U8681 (N_8681,N_4924,N_3431);
nor U8682 (N_8682,N_2154,N_3844);
and U8683 (N_8683,N_4466,N_4017);
nand U8684 (N_8684,N_2055,N_2889);
nor U8685 (N_8685,N_3895,N_2142);
nor U8686 (N_8686,N_558,N_4484);
or U8687 (N_8687,N_3119,N_4035);
or U8688 (N_8688,N_536,N_1945);
xnor U8689 (N_8689,N_1556,N_1732);
nand U8690 (N_8690,N_2665,N_1403);
and U8691 (N_8691,N_92,N_2805);
or U8692 (N_8692,N_3873,N_968);
nor U8693 (N_8693,N_2290,N_3801);
or U8694 (N_8694,N_3147,N_2792);
xnor U8695 (N_8695,N_418,N_2027);
nand U8696 (N_8696,N_1794,N_3213);
nand U8697 (N_8697,N_1749,N_1679);
nor U8698 (N_8698,N_4156,N_3626);
and U8699 (N_8699,N_2448,N_313);
or U8700 (N_8700,N_3705,N_1637);
and U8701 (N_8701,N_3796,N_1088);
or U8702 (N_8702,N_1039,N_238);
xnor U8703 (N_8703,N_1142,N_3006);
or U8704 (N_8704,N_4938,N_3344);
or U8705 (N_8705,N_3508,N_892);
nor U8706 (N_8706,N_4191,N_1331);
nor U8707 (N_8707,N_1541,N_2974);
nand U8708 (N_8708,N_2709,N_4548);
or U8709 (N_8709,N_2943,N_277);
or U8710 (N_8710,N_686,N_3480);
nand U8711 (N_8711,N_186,N_4301);
nand U8712 (N_8712,N_3951,N_2540);
and U8713 (N_8713,N_4933,N_3176);
nor U8714 (N_8714,N_2588,N_1993);
nor U8715 (N_8715,N_1576,N_3181);
nor U8716 (N_8716,N_872,N_2765);
and U8717 (N_8717,N_3263,N_4617);
or U8718 (N_8718,N_3615,N_3352);
and U8719 (N_8719,N_4416,N_3161);
and U8720 (N_8720,N_4638,N_1458);
and U8721 (N_8721,N_997,N_2744);
nor U8722 (N_8722,N_4936,N_4498);
and U8723 (N_8723,N_2533,N_1241);
nor U8724 (N_8724,N_1512,N_4988);
and U8725 (N_8725,N_1415,N_1647);
or U8726 (N_8726,N_1969,N_1859);
nand U8727 (N_8727,N_4037,N_1742);
xnor U8728 (N_8728,N_4096,N_4682);
nor U8729 (N_8729,N_2186,N_4921);
and U8730 (N_8730,N_4324,N_2542);
nand U8731 (N_8731,N_1101,N_2368);
nor U8732 (N_8732,N_2347,N_1039);
nand U8733 (N_8733,N_1654,N_2865);
xnor U8734 (N_8734,N_3384,N_3396);
nor U8735 (N_8735,N_4199,N_4722);
nor U8736 (N_8736,N_3677,N_4254);
nand U8737 (N_8737,N_2457,N_4910);
or U8738 (N_8738,N_605,N_3433);
nor U8739 (N_8739,N_1584,N_2399);
nand U8740 (N_8740,N_3920,N_2013);
xor U8741 (N_8741,N_777,N_80);
nand U8742 (N_8742,N_4803,N_3611);
nand U8743 (N_8743,N_1746,N_4707);
xor U8744 (N_8744,N_2805,N_3548);
and U8745 (N_8745,N_3216,N_1380);
or U8746 (N_8746,N_3354,N_2475);
nand U8747 (N_8747,N_567,N_4430);
and U8748 (N_8748,N_492,N_1350);
and U8749 (N_8749,N_2076,N_469);
or U8750 (N_8750,N_4964,N_290);
and U8751 (N_8751,N_1899,N_3740);
nand U8752 (N_8752,N_4551,N_836);
and U8753 (N_8753,N_1666,N_1925);
nand U8754 (N_8754,N_3308,N_2911);
and U8755 (N_8755,N_2884,N_2221);
nand U8756 (N_8756,N_4069,N_503);
and U8757 (N_8757,N_2613,N_2135);
or U8758 (N_8758,N_3394,N_79);
and U8759 (N_8759,N_4879,N_4971);
and U8760 (N_8760,N_730,N_4971);
or U8761 (N_8761,N_3376,N_3591);
or U8762 (N_8762,N_1560,N_4160);
nor U8763 (N_8763,N_3867,N_154);
nor U8764 (N_8764,N_4289,N_1636);
and U8765 (N_8765,N_2699,N_2184);
nand U8766 (N_8766,N_1178,N_47);
and U8767 (N_8767,N_1632,N_8);
or U8768 (N_8768,N_3722,N_1063);
nor U8769 (N_8769,N_260,N_651);
nor U8770 (N_8770,N_4446,N_1417);
and U8771 (N_8771,N_667,N_2513);
and U8772 (N_8772,N_1650,N_2596);
nand U8773 (N_8773,N_1047,N_4139);
or U8774 (N_8774,N_2352,N_3770);
and U8775 (N_8775,N_4518,N_1857);
xnor U8776 (N_8776,N_1585,N_3670);
nand U8777 (N_8777,N_4642,N_4209);
and U8778 (N_8778,N_1730,N_3979);
and U8779 (N_8779,N_1198,N_4186);
xor U8780 (N_8780,N_3260,N_2332);
nand U8781 (N_8781,N_1812,N_2746);
or U8782 (N_8782,N_3620,N_2362);
or U8783 (N_8783,N_4897,N_3411);
xor U8784 (N_8784,N_671,N_207);
nor U8785 (N_8785,N_1219,N_3264);
and U8786 (N_8786,N_1978,N_3413);
nand U8787 (N_8787,N_3638,N_1838);
nand U8788 (N_8788,N_3139,N_3182);
nor U8789 (N_8789,N_4332,N_4253);
nor U8790 (N_8790,N_1446,N_3916);
or U8791 (N_8791,N_537,N_2450);
nand U8792 (N_8792,N_3750,N_3848);
nor U8793 (N_8793,N_3544,N_633);
and U8794 (N_8794,N_3199,N_1531);
nand U8795 (N_8795,N_3560,N_274);
xor U8796 (N_8796,N_1185,N_4043);
nand U8797 (N_8797,N_4282,N_1832);
nand U8798 (N_8798,N_1489,N_4456);
nand U8799 (N_8799,N_3353,N_460);
and U8800 (N_8800,N_4149,N_1192);
nand U8801 (N_8801,N_3932,N_552);
or U8802 (N_8802,N_2149,N_3728);
nor U8803 (N_8803,N_3612,N_4361);
nor U8804 (N_8804,N_4343,N_1561);
nand U8805 (N_8805,N_505,N_1903);
nor U8806 (N_8806,N_1012,N_801);
and U8807 (N_8807,N_1654,N_4445);
nor U8808 (N_8808,N_1547,N_2132);
and U8809 (N_8809,N_4078,N_4083);
nor U8810 (N_8810,N_3158,N_1890);
and U8811 (N_8811,N_2741,N_3211);
nand U8812 (N_8812,N_4223,N_4414);
nand U8813 (N_8813,N_2345,N_3066);
nor U8814 (N_8814,N_1187,N_924);
and U8815 (N_8815,N_1777,N_3650);
nand U8816 (N_8816,N_3349,N_4477);
nor U8817 (N_8817,N_4410,N_2029);
or U8818 (N_8818,N_3518,N_3432);
nor U8819 (N_8819,N_3767,N_1544);
nand U8820 (N_8820,N_1652,N_87);
nor U8821 (N_8821,N_1795,N_439);
nor U8822 (N_8822,N_511,N_999);
and U8823 (N_8823,N_3597,N_2860);
nor U8824 (N_8824,N_1559,N_2793);
nor U8825 (N_8825,N_1862,N_1465);
xor U8826 (N_8826,N_3320,N_4929);
or U8827 (N_8827,N_1196,N_3393);
xnor U8828 (N_8828,N_331,N_446);
and U8829 (N_8829,N_2456,N_3641);
or U8830 (N_8830,N_2953,N_4383);
and U8831 (N_8831,N_454,N_56);
nor U8832 (N_8832,N_112,N_1330);
nor U8833 (N_8833,N_2538,N_4568);
nor U8834 (N_8834,N_867,N_4741);
nor U8835 (N_8835,N_3369,N_2167);
or U8836 (N_8836,N_4411,N_773);
nand U8837 (N_8837,N_213,N_1998);
nor U8838 (N_8838,N_1320,N_1811);
xor U8839 (N_8839,N_4569,N_2954);
nand U8840 (N_8840,N_963,N_2238);
nor U8841 (N_8841,N_1498,N_2540);
nor U8842 (N_8842,N_2230,N_1502);
nor U8843 (N_8843,N_1564,N_1910);
nor U8844 (N_8844,N_3262,N_3717);
nand U8845 (N_8845,N_3161,N_4270);
and U8846 (N_8846,N_1679,N_2803);
nand U8847 (N_8847,N_1130,N_813);
nand U8848 (N_8848,N_217,N_2871);
nor U8849 (N_8849,N_3610,N_3360);
xor U8850 (N_8850,N_4510,N_2354);
nand U8851 (N_8851,N_4576,N_766);
nand U8852 (N_8852,N_4324,N_4255);
and U8853 (N_8853,N_2766,N_1701);
nor U8854 (N_8854,N_2927,N_2591);
and U8855 (N_8855,N_783,N_178);
or U8856 (N_8856,N_4635,N_636);
nor U8857 (N_8857,N_4688,N_1439);
and U8858 (N_8858,N_4230,N_2111);
and U8859 (N_8859,N_2744,N_2839);
nor U8860 (N_8860,N_1786,N_4486);
nand U8861 (N_8861,N_2863,N_1148);
or U8862 (N_8862,N_4916,N_1088);
nand U8863 (N_8863,N_4494,N_4397);
nand U8864 (N_8864,N_3578,N_4011);
nor U8865 (N_8865,N_1121,N_2956);
xnor U8866 (N_8866,N_3068,N_116);
and U8867 (N_8867,N_1080,N_3593);
nor U8868 (N_8868,N_2907,N_2087);
or U8869 (N_8869,N_4663,N_49);
and U8870 (N_8870,N_4779,N_3160);
nor U8871 (N_8871,N_2618,N_436);
nor U8872 (N_8872,N_3265,N_3128);
or U8873 (N_8873,N_1680,N_536);
nand U8874 (N_8874,N_2976,N_3940);
nor U8875 (N_8875,N_4967,N_730);
nor U8876 (N_8876,N_1829,N_305);
or U8877 (N_8877,N_2874,N_3341);
or U8878 (N_8878,N_3046,N_2002);
nor U8879 (N_8879,N_4745,N_1867);
nor U8880 (N_8880,N_645,N_2492);
xnor U8881 (N_8881,N_2197,N_1971);
or U8882 (N_8882,N_2467,N_4464);
nand U8883 (N_8883,N_270,N_2345);
and U8884 (N_8884,N_2542,N_2552);
nand U8885 (N_8885,N_263,N_1794);
nand U8886 (N_8886,N_1430,N_2412);
nand U8887 (N_8887,N_2219,N_3605);
nand U8888 (N_8888,N_3592,N_3059);
xnor U8889 (N_8889,N_1245,N_3841);
or U8890 (N_8890,N_3316,N_1851);
nand U8891 (N_8891,N_3711,N_555);
or U8892 (N_8892,N_1621,N_2818);
and U8893 (N_8893,N_1100,N_4106);
xnor U8894 (N_8894,N_2358,N_1025);
nand U8895 (N_8895,N_1849,N_2490);
nand U8896 (N_8896,N_3645,N_3623);
nor U8897 (N_8897,N_2472,N_3864);
or U8898 (N_8898,N_2078,N_4630);
nand U8899 (N_8899,N_2853,N_2401);
xnor U8900 (N_8900,N_4157,N_2715);
nand U8901 (N_8901,N_3565,N_1342);
or U8902 (N_8902,N_274,N_1948);
nor U8903 (N_8903,N_889,N_4165);
nand U8904 (N_8904,N_266,N_2082);
and U8905 (N_8905,N_274,N_4471);
or U8906 (N_8906,N_3978,N_3850);
nand U8907 (N_8907,N_529,N_4072);
or U8908 (N_8908,N_4677,N_2510);
nor U8909 (N_8909,N_1107,N_1029);
nand U8910 (N_8910,N_3820,N_631);
and U8911 (N_8911,N_2715,N_3481);
xnor U8912 (N_8912,N_484,N_3034);
and U8913 (N_8913,N_275,N_3414);
nor U8914 (N_8914,N_2491,N_3723);
nand U8915 (N_8915,N_1230,N_760);
or U8916 (N_8916,N_3119,N_2287);
nor U8917 (N_8917,N_2665,N_2078);
nand U8918 (N_8918,N_3886,N_1224);
nand U8919 (N_8919,N_2384,N_2420);
or U8920 (N_8920,N_3788,N_3102);
nor U8921 (N_8921,N_770,N_4445);
xnor U8922 (N_8922,N_3434,N_1104);
or U8923 (N_8923,N_4949,N_3630);
and U8924 (N_8924,N_2723,N_2278);
nand U8925 (N_8925,N_2491,N_3028);
nand U8926 (N_8926,N_4949,N_1739);
xor U8927 (N_8927,N_178,N_3487);
nor U8928 (N_8928,N_3303,N_2593);
xnor U8929 (N_8929,N_809,N_878);
and U8930 (N_8930,N_2352,N_4112);
or U8931 (N_8931,N_2878,N_4563);
nor U8932 (N_8932,N_4678,N_3678);
and U8933 (N_8933,N_1336,N_1202);
and U8934 (N_8934,N_2917,N_1040);
or U8935 (N_8935,N_2278,N_2689);
nor U8936 (N_8936,N_4904,N_651);
or U8937 (N_8937,N_934,N_3465);
or U8938 (N_8938,N_1088,N_4909);
xor U8939 (N_8939,N_4124,N_362);
and U8940 (N_8940,N_3368,N_253);
and U8941 (N_8941,N_3358,N_760);
nor U8942 (N_8942,N_1805,N_2783);
and U8943 (N_8943,N_4598,N_1082);
nor U8944 (N_8944,N_2106,N_2783);
and U8945 (N_8945,N_744,N_4282);
and U8946 (N_8946,N_6,N_1067);
nand U8947 (N_8947,N_2101,N_1672);
nand U8948 (N_8948,N_1160,N_2239);
xnor U8949 (N_8949,N_815,N_1621);
xor U8950 (N_8950,N_93,N_2800);
nor U8951 (N_8951,N_4500,N_2345);
nand U8952 (N_8952,N_3527,N_4333);
nand U8953 (N_8953,N_1236,N_4036);
and U8954 (N_8954,N_3545,N_2769);
nand U8955 (N_8955,N_4376,N_2904);
or U8956 (N_8956,N_1770,N_2970);
nand U8957 (N_8957,N_2198,N_3046);
xor U8958 (N_8958,N_3569,N_1667);
nor U8959 (N_8959,N_3260,N_3042);
xor U8960 (N_8960,N_3565,N_4018);
nand U8961 (N_8961,N_3282,N_3599);
nor U8962 (N_8962,N_4949,N_4426);
nand U8963 (N_8963,N_4220,N_203);
nor U8964 (N_8964,N_1864,N_1335);
nand U8965 (N_8965,N_1530,N_2861);
and U8966 (N_8966,N_1892,N_2168);
xor U8967 (N_8967,N_4338,N_503);
nor U8968 (N_8968,N_406,N_3671);
nor U8969 (N_8969,N_3907,N_3205);
or U8970 (N_8970,N_3040,N_3804);
nand U8971 (N_8971,N_2464,N_1565);
and U8972 (N_8972,N_1553,N_4371);
and U8973 (N_8973,N_3415,N_1701);
or U8974 (N_8974,N_2888,N_3101);
or U8975 (N_8975,N_11,N_2095);
nand U8976 (N_8976,N_4454,N_1982);
and U8977 (N_8977,N_3667,N_779);
and U8978 (N_8978,N_1597,N_2081);
and U8979 (N_8979,N_3427,N_1189);
nor U8980 (N_8980,N_3708,N_843);
and U8981 (N_8981,N_3286,N_1840);
and U8982 (N_8982,N_730,N_4876);
nand U8983 (N_8983,N_4800,N_1899);
nand U8984 (N_8984,N_4393,N_2317);
nand U8985 (N_8985,N_3189,N_3294);
or U8986 (N_8986,N_1654,N_454);
xnor U8987 (N_8987,N_92,N_2490);
nor U8988 (N_8988,N_4479,N_256);
or U8989 (N_8989,N_1199,N_3792);
nand U8990 (N_8990,N_2376,N_371);
nand U8991 (N_8991,N_1680,N_2589);
or U8992 (N_8992,N_3339,N_2423);
nand U8993 (N_8993,N_4019,N_2107);
xor U8994 (N_8994,N_3879,N_4193);
nor U8995 (N_8995,N_3357,N_4278);
or U8996 (N_8996,N_1261,N_4896);
nor U8997 (N_8997,N_4956,N_2229);
nand U8998 (N_8998,N_1660,N_3616);
xor U8999 (N_8999,N_472,N_1239);
nor U9000 (N_9000,N_2236,N_1011);
or U9001 (N_9001,N_3144,N_316);
nor U9002 (N_9002,N_1221,N_913);
and U9003 (N_9003,N_3084,N_1441);
and U9004 (N_9004,N_4230,N_3014);
nor U9005 (N_9005,N_1522,N_2451);
and U9006 (N_9006,N_3365,N_2604);
and U9007 (N_9007,N_1929,N_895);
nor U9008 (N_9008,N_757,N_2091);
xor U9009 (N_9009,N_907,N_4708);
nor U9010 (N_9010,N_0,N_1519);
and U9011 (N_9011,N_4103,N_1422);
xor U9012 (N_9012,N_2089,N_3513);
nand U9013 (N_9013,N_1867,N_1159);
or U9014 (N_9014,N_2163,N_212);
nor U9015 (N_9015,N_4471,N_1689);
xor U9016 (N_9016,N_527,N_1978);
nand U9017 (N_9017,N_3046,N_2245);
nand U9018 (N_9018,N_2266,N_1367);
and U9019 (N_9019,N_2298,N_2402);
or U9020 (N_9020,N_1221,N_2779);
or U9021 (N_9021,N_4989,N_3981);
xnor U9022 (N_9022,N_2004,N_517);
nor U9023 (N_9023,N_2531,N_4648);
or U9024 (N_9024,N_4765,N_693);
or U9025 (N_9025,N_3496,N_1193);
and U9026 (N_9026,N_89,N_3373);
nor U9027 (N_9027,N_4566,N_4191);
and U9028 (N_9028,N_3367,N_4587);
nor U9029 (N_9029,N_4214,N_1373);
nand U9030 (N_9030,N_3802,N_4763);
or U9031 (N_9031,N_586,N_3768);
nor U9032 (N_9032,N_1664,N_4642);
or U9033 (N_9033,N_4954,N_1430);
or U9034 (N_9034,N_1308,N_2132);
nor U9035 (N_9035,N_2947,N_2862);
nand U9036 (N_9036,N_3184,N_2408);
nor U9037 (N_9037,N_4544,N_2244);
nor U9038 (N_9038,N_4094,N_4546);
nand U9039 (N_9039,N_639,N_3244);
nor U9040 (N_9040,N_422,N_1170);
or U9041 (N_9041,N_3876,N_906);
or U9042 (N_9042,N_627,N_3225);
nand U9043 (N_9043,N_1037,N_575);
nand U9044 (N_9044,N_590,N_2453);
and U9045 (N_9045,N_2473,N_2416);
nand U9046 (N_9046,N_518,N_4653);
nand U9047 (N_9047,N_1087,N_4607);
xor U9048 (N_9048,N_969,N_1473);
xnor U9049 (N_9049,N_2591,N_1285);
and U9050 (N_9050,N_1583,N_1897);
nor U9051 (N_9051,N_1634,N_114);
and U9052 (N_9052,N_3176,N_1697);
nand U9053 (N_9053,N_1986,N_1504);
nor U9054 (N_9054,N_1312,N_3915);
or U9055 (N_9055,N_294,N_2975);
xor U9056 (N_9056,N_371,N_3636);
nor U9057 (N_9057,N_4894,N_4226);
nor U9058 (N_9058,N_3474,N_175);
nand U9059 (N_9059,N_3147,N_1734);
xnor U9060 (N_9060,N_929,N_286);
nor U9061 (N_9061,N_3538,N_3416);
nand U9062 (N_9062,N_475,N_2893);
or U9063 (N_9063,N_3994,N_2393);
xor U9064 (N_9064,N_4637,N_113);
nor U9065 (N_9065,N_463,N_3942);
nor U9066 (N_9066,N_4036,N_2124);
nand U9067 (N_9067,N_4001,N_3780);
or U9068 (N_9068,N_1551,N_2536);
nand U9069 (N_9069,N_1963,N_4746);
or U9070 (N_9070,N_1737,N_1329);
nand U9071 (N_9071,N_3636,N_1369);
and U9072 (N_9072,N_3174,N_1213);
nand U9073 (N_9073,N_4050,N_138);
nor U9074 (N_9074,N_2189,N_1259);
nand U9075 (N_9075,N_3985,N_3948);
nand U9076 (N_9076,N_2357,N_4795);
and U9077 (N_9077,N_1417,N_3112);
xnor U9078 (N_9078,N_1975,N_3184);
nand U9079 (N_9079,N_3267,N_3155);
nand U9080 (N_9080,N_2495,N_2399);
xnor U9081 (N_9081,N_3794,N_1604);
or U9082 (N_9082,N_2145,N_3951);
nand U9083 (N_9083,N_3307,N_4891);
nand U9084 (N_9084,N_3333,N_248);
nor U9085 (N_9085,N_1616,N_250);
and U9086 (N_9086,N_1572,N_2531);
xor U9087 (N_9087,N_1366,N_1985);
nand U9088 (N_9088,N_1785,N_2004);
and U9089 (N_9089,N_281,N_4736);
nand U9090 (N_9090,N_618,N_3744);
xor U9091 (N_9091,N_2575,N_2778);
nand U9092 (N_9092,N_4445,N_1931);
nand U9093 (N_9093,N_704,N_1757);
nor U9094 (N_9094,N_1048,N_1450);
nand U9095 (N_9095,N_527,N_3780);
nor U9096 (N_9096,N_3374,N_3895);
xor U9097 (N_9097,N_4657,N_3104);
nor U9098 (N_9098,N_648,N_3303);
nor U9099 (N_9099,N_2356,N_1861);
nor U9100 (N_9100,N_987,N_3581);
nand U9101 (N_9101,N_3766,N_1431);
nand U9102 (N_9102,N_3599,N_2489);
nor U9103 (N_9103,N_4013,N_4239);
or U9104 (N_9104,N_22,N_1711);
or U9105 (N_9105,N_379,N_3575);
nand U9106 (N_9106,N_2644,N_3354);
or U9107 (N_9107,N_1297,N_1199);
or U9108 (N_9108,N_4880,N_1561);
and U9109 (N_9109,N_4196,N_719);
nor U9110 (N_9110,N_4875,N_4221);
nand U9111 (N_9111,N_3090,N_2213);
and U9112 (N_9112,N_3303,N_1030);
nor U9113 (N_9113,N_4025,N_2449);
nand U9114 (N_9114,N_3103,N_2960);
and U9115 (N_9115,N_4100,N_2696);
nand U9116 (N_9116,N_465,N_782);
and U9117 (N_9117,N_1599,N_4260);
nor U9118 (N_9118,N_3630,N_1992);
and U9119 (N_9119,N_1495,N_3000);
or U9120 (N_9120,N_67,N_2225);
nor U9121 (N_9121,N_1650,N_4169);
nor U9122 (N_9122,N_383,N_2055);
nand U9123 (N_9123,N_4242,N_1788);
nand U9124 (N_9124,N_558,N_1105);
nand U9125 (N_9125,N_4126,N_4864);
or U9126 (N_9126,N_4593,N_2010);
and U9127 (N_9127,N_3452,N_4323);
nor U9128 (N_9128,N_3501,N_1942);
nand U9129 (N_9129,N_4503,N_4783);
xor U9130 (N_9130,N_3035,N_2880);
or U9131 (N_9131,N_4757,N_986);
or U9132 (N_9132,N_3017,N_3479);
nor U9133 (N_9133,N_610,N_1376);
nand U9134 (N_9134,N_4667,N_4878);
xor U9135 (N_9135,N_1781,N_3325);
or U9136 (N_9136,N_1090,N_2926);
nor U9137 (N_9137,N_4945,N_2639);
xor U9138 (N_9138,N_2155,N_788);
and U9139 (N_9139,N_1691,N_1259);
xor U9140 (N_9140,N_4660,N_2635);
xor U9141 (N_9141,N_15,N_4336);
nand U9142 (N_9142,N_3709,N_3427);
or U9143 (N_9143,N_1538,N_939);
nor U9144 (N_9144,N_1349,N_4961);
nand U9145 (N_9145,N_957,N_3986);
or U9146 (N_9146,N_943,N_726);
or U9147 (N_9147,N_1538,N_3622);
nand U9148 (N_9148,N_1035,N_3494);
and U9149 (N_9149,N_4093,N_4589);
or U9150 (N_9150,N_1519,N_1744);
nor U9151 (N_9151,N_3619,N_4577);
and U9152 (N_9152,N_4128,N_1815);
and U9153 (N_9153,N_2100,N_570);
or U9154 (N_9154,N_1094,N_4976);
nor U9155 (N_9155,N_4121,N_571);
nand U9156 (N_9156,N_423,N_3364);
nand U9157 (N_9157,N_4475,N_3280);
and U9158 (N_9158,N_1936,N_2905);
nor U9159 (N_9159,N_4004,N_1898);
xor U9160 (N_9160,N_532,N_3261);
xnor U9161 (N_9161,N_3198,N_2471);
nor U9162 (N_9162,N_1399,N_1346);
and U9163 (N_9163,N_429,N_2958);
nand U9164 (N_9164,N_4227,N_1818);
nor U9165 (N_9165,N_2196,N_4419);
or U9166 (N_9166,N_4936,N_2590);
or U9167 (N_9167,N_760,N_4100);
nand U9168 (N_9168,N_283,N_2159);
xor U9169 (N_9169,N_1045,N_3183);
nand U9170 (N_9170,N_4188,N_3267);
and U9171 (N_9171,N_733,N_287);
or U9172 (N_9172,N_2754,N_3516);
nand U9173 (N_9173,N_1956,N_3391);
xnor U9174 (N_9174,N_4269,N_2075);
nor U9175 (N_9175,N_2012,N_1226);
nand U9176 (N_9176,N_1239,N_2401);
nand U9177 (N_9177,N_3345,N_3417);
nor U9178 (N_9178,N_2086,N_1498);
and U9179 (N_9179,N_841,N_2620);
and U9180 (N_9180,N_1413,N_4418);
xnor U9181 (N_9181,N_4264,N_2465);
and U9182 (N_9182,N_3921,N_563);
and U9183 (N_9183,N_4124,N_4840);
or U9184 (N_9184,N_1631,N_2378);
nor U9185 (N_9185,N_1166,N_1117);
and U9186 (N_9186,N_2640,N_6);
nand U9187 (N_9187,N_4577,N_1957);
or U9188 (N_9188,N_2528,N_4219);
and U9189 (N_9189,N_1396,N_2709);
nand U9190 (N_9190,N_3360,N_1419);
nand U9191 (N_9191,N_1949,N_1055);
xnor U9192 (N_9192,N_3975,N_370);
and U9193 (N_9193,N_2283,N_1610);
or U9194 (N_9194,N_2256,N_4690);
nor U9195 (N_9195,N_1486,N_1653);
xnor U9196 (N_9196,N_1602,N_726);
and U9197 (N_9197,N_3481,N_893);
nor U9198 (N_9198,N_892,N_2783);
nand U9199 (N_9199,N_3271,N_220);
and U9200 (N_9200,N_251,N_2251);
nand U9201 (N_9201,N_445,N_2034);
xnor U9202 (N_9202,N_704,N_428);
nor U9203 (N_9203,N_2545,N_2725);
and U9204 (N_9204,N_3133,N_1984);
nor U9205 (N_9205,N_4969,N_2162);
and U9206 (N_9206,N_239,N_1610);
nand U9207 (N_9207,N_331,N_4888);
and U9208 (N_9208,N_3733,N_4214);
nand U9209 (N_9209,N_533,N_3552);
or U9210 (N_9210,N_647,N_4522);
and U9211 (N_9211,N_4575,N_2242);
nand U9212 (N_9212,N_3371,N_2239);
nand U9213 (N_9213,N_2804,N_775);
nand U9214 (N_9214,N_4477,N_849);
nor U9215 (N_9215,N_3790,N_3771);
nor U9216 (N_9216,N_1771,N_3229);
nor U9217 (N_9217,N_2608,N_1860);
nand U9218 (N_9218,N_918,N_1960);
or U9219 (N_9219,N_621,N_4410);
nand U9220 (N_9220,N_743,N_3426);
or U9221 (N_9221,N_2745,N_780);
nand U9222 (N_9222,N_286,N_385);
nand U9223 (N_9223,N_3736,N_1435);
nand U9224 (N_9224,N_2881,N_4553);
and U9225 (N_9225,N_284,N_2687);
and U9226 (N_9226,N_1066,N_2173);
or U9227 (N_9227,N_2249,N_2276);
nor U9228 (N_9228,N_1597,N_3871);
or U9229 (N_9229,N_2772,N_1334);
nand U9230 (N_9230,N_1979,N_1630);
or U9231 (N_9231,N_1582,N_4190);
or U9232 (N_9232,N_1742,N_1672);
nor U9233 (N_9233,N_2220,N_4537);
nor U9234 (N_9234,N_3775,N_4767);
nand U9235 (N_9235,N_4337,N_450);
nor U9236 (N_9236,N_4091,N_4614);
and U9237 (N_9237,N_585,N_2046);
nand U9238 (N_9238,N_601,N_4719);
and U9239 (N_9239,N_1994,N_4769);
xnor U9240 (N_9240,N_697,N_219);
and U9241 (N_9241,N_2250,N_2043);
and U9242 (N_9242,N_122,N_564);
nor U9243 (N_9243,N_4578,N_929);
nor U9244 (N_9244,N_2879,N_3611);
nor U9245 (N_9245,N_4363,N_537);
xnor U9246 (N_9246,N_121,N_4010);
xnor U9247 (N_9247,N_4963,N_1063);
or U9248 (N_9248,N_4106,N_4246);
and U9249 (N_9249,N_327,N_1048);
nand U9250 (N_9250,N_1829,N_2495);
and U9251 (N_9251,N_3882,N_2302);
or U9252 (N_9252,N_1981,N_4446);
nand U9253 (N_9253,N_2915,N_4187);
nor U9254 (N_9254,N_2398,N_1073);
or U9255 (N_9255,N_3954,N_835);
nand U9256 (N_9256,N_1139,N_3889);
nand U9257 (N_9257,N_4704,N_3425);
nor U9258 (N_9258,N_1419,N_1259);
or U9259 (N_9259,N_4269,N_2473);
and U9260 (N_9260,N_1029,N_1224);
nand U9261 (N_9261,N_3193,N_337);
or U9262 (N_9262,N_2994,N_3072);
and U9263 (N_9263,N_4146,N_2348);
and U9264 (N_9264,N_4925,N_2681);
nand U9265 (N_9265,N_2616,N_1672);
xnor U9266 (N_9266,N_2942,N_2507);
and U9267 (N_9267,N_3841,N_11);
nand U9268 (N_9268,N_1738,N_446);
xnor U9269 (N_9269,N_4038,N_2885);
xor U9270 (N_9270,N_1507,N_3374);
nor U9271 (N_9271,N_4919,N_507);
and U9272 (N_9272,N_4819,N_4146);
or U9273 (N_9273,N_1892,N_4709);
nand U9274 (N_9274,N_4361,N_3564);
nor U9275 (N_9275,N_2647,N_457);
nor U9276 (N_9276,N_4739,N_4620);
xnor U9277 (N_9277,N_968,N_35);
or U9278 (N_9278,N_2720,N_899);
nand U9279 (N_9279,N_787,N_1134);
and U9280 (N_9280,N_3876,N_2340);
and U9281 (N_9281,N_3631,N_997);
and U9282 (N_9282,N_4332,N_2850);
nand U9283 (N_9283,N_450,N_4907);
and U9284 (N_9284,N_2508,N_679);
nand U9285 (N_9285,N_647,N_1888);
or U9286 (N_9286,N_1232,N_4659);
or U9287 (N_9287,N_2963,N_4016);
or U9288 (N_9288,N_725,N_1450);
xor U9289 (N_9289,N_4632,N_2677);
nand U9290 (N_9290,N_3984,N_2054);
and U9291 (N_9291,N_3426,N_3834);
nor U9292 (N_9292,N_296,N_2879);
nand U9293 (N_9293,N_231,N_3931);
and U9294 (N_9294,N_381,N_3364);
nand U9295 (N_9295,N_1039,N_2435);
nand U9296 (N_9296,N_1802,N_4856);
and U9297 (N_9297,N_2165,N_3531);
and U9298 (N_9298,N_3505,N_2443);
nand U9299 (N_9299,N_1356,N_4660);
nand U9300 (N_9300,N_4809,N_813);
nand U9301 (N_9301,N_4836,N_4591);
and U9302 (N_9302,N_1390,N_3524);
and U9303 (N_9303,N_4256,N_1998);
nor U9304 (N_9304,N_1653,N_2936);
and U9305 (N_9305,N_4325,N_2948);
nor U9306 (N_9306,N_460,N_2553);
nand U9307 (N_9307,N_1085,N_2009);
or U9308 (N_9308,N_3721,N_546);
or U9309 (N_9309,N_2066,N_1117);
or U9310 (N_9310,N_3202,N_3174);
or U9311 (N_9311,N_2636,N_2585);
and U9312 (N_9312,N_590,N_1552);
and U9313 (N_9313,N_2911,N_4504);
nand U9314 (N_9314,N_2081,N_4850);
xnor U9315 (N_9315,N_3035,N_467);
or U9316 (N_9316,N_4313,N_4819);
or U9317 (N_9317,N_4596,N_3268);
nand U9318 (N_9318,N_2621,N_3317);
or U9319 (N_9319,N_2979,N_1057);
and U9320 (N_9320,N_2627,N_424);
or U9321 (N_9321,N_2026,N_3723);
xnor U9322 (N_9322,N_3124,N_2796);
nand U9323 (N_9323,N_3506,N_2059);
nand U9324 (N_9324,N_1426,N_3691);
or U9325 (N_9325,N_1335,N_4791);
or U9326 (N_9326,N_4618,N_4213);
nor U9327 (N_9327,N_3568,N_3259);
and U9328 (N_9328,N_2736,N_1644);
nand U9329 (N_9329,N_2627,N_3582);
nand U9330 (N_9330,N_4568,N_1199);
and U9331 (N_9331,N_3675,N_3879);
nor U9332 (N_9332,N_4088,N_2615);
nor U9333 (N_9333,N_375,N_2107);
or U9334 (N_9334,N_302,N_3561);
and U9335 (N_9335,N_1838,N_2259);
or U9336 (N_9336,N_1387,N_48);
or U9337 (N_9337,N_4918,N_1828);
nor U9338 (N_9338,N_1438,N_1180);
nand U9339 (N_9339,N_4669,N_2672);
xnor U9340 (N_9340,N_3058,N_1386);
and U9341 (N_9341,N_4600,N_858);
nor U9342 (N_9342,N_4645,N_4804);
xor U9343 (N_9343,N_620,N_1184);
nor U9344 (N_9344,N_661,N_2867);
nand U9345 (N_9345,N_3970,N_1286);
nor U9346 (N_9346,N_1119,N_1811);
nand U9347 (N_9347,N_2825,N_4423);
or U9348 (N_9348,N_2651,N_3832);
nand U9349 (N_9349,N_4044,N_3320);
nand U9350 (N_9350,N_1988,N_1912);
or U9351 (N_9351,N_1653,N_3974);
or U9352 (N_9352,N_1927,N_3336);
or U9353 (N_9353,N_3072,N_4151);
nand U9354 (N_9354,N_3192,N_2989);
or U9355 (N_9355,N_1007,N_1008);
nand U9356 (N_9356,N_3002,N_4960);
nor U9357 (N_9357,N_2592,N_1311);
xor U9358 (N_9358,N_3622,N_4283);
or U9359 (N_9359,N_743,N_2716);
and U9360 (N_9360,N_3302,N_4825);
nor U9361 (N_9361,N_3977,N_3532);
nor U9362 (N_9362,N_4690,N_3522);
or U9363 (N_9363,N_2287,N_939);
nor U9364 (N_9364,N_2008,N_3935);
nor U9365 (N_9365,N_1257,N_4231);
and U9366 (N_9366,N_4389,N_4928);
or U9367 (N_9367,N_154,N_3291);
nor U9368 (N_9368,N_3144,N_1016);
nor U9369 (N_9369,N_256,N_2536);
and U9370 (N_9370,N_1026,N_991);
nor U9371 (N_9371,N_4449,N_272);
nor U9372 (N_9372,N_3865,N_978);
or U9373 (N_9373,N_930,N_3358);
nor U9374 (N_9374,N_390,N_1998);
xnor U9375 (N_9375,N_37,N_3967);
and U9376 (N_9376,N_3874,N_3746);
or U9377 (N_9377,N_1799,N_152);
nor U9378 (N_9378,N_3526,N_1247);
xnor U9379 (N_9379,N_1280,N_107);
nand U9380 (N_9380,N_3773,N_723);
and U9381 (N_9381,N_4441,N_3578);
and U9382 (N_9382,N_1515,N_474);
nor U9383 (N_9383,N_3950,N_2611);
nor U9384 (N_9384,N_2947,N_3233);
and U9385 (N_9385,N_3186,N_3486);
nor U9386 (N_9386,N_3876,N_3023);
xor U9387 (N_9387,N_2753,N_3318);
nand U9388 (N_9388,N_732,N_4747);
nor U9389 (N_9389,N_4783,N_1527);
nor U9390 (N_9390,N_354,N_3563);
or U9391 (N_9391,N_3597,N_3929);
and U9392 (N_9392,N_3071,N_2435);
nand U9393 (N_9393,N_442,N_2918);
nand U9394 (N_9394,N_1901,N_1084);
nand U9395 (N_9395,N_2817,N_3708);
or U9396 (N_9396,N_4829,N_88);
and U9397 (N_9397,N_790,N_487);
nor U9398 (N_9398,N_1633,N_3524);
or U9399 (N_9399,N_3772,N_4722);
and U9400 (N_9400,N_4853,N_1469);
nor U9401 (N_9401,N_4108,N_3622);
and U9402 (N_9402,N_954,N_1348);
or U9403 (N_9403,N_3929,N_3085);
xnor U9404 (N_9404,N_3012,N_4594);
nor U9405 (N_9405,N_1414,N_434);
and U9406 (N_9406,N_4922,N_1065);
nand U9407 (N_9407,N_4446,N_580);
xor U9408 (N_9408,N_4620,N_3032);
and U9409 (N_9409,N_1415,N_3269);
nor U9410 (N_9410,N_4793,N_2761);
and U9411 (N_9411,N_1917,N_1432);
xnor U9412 (N_9412,N_1914,N_150);
nand U9413 (N_9413,N_2782,N_99);
or U9414 (N_9414,N_888,N_1713);
nand U9415 (N_9415,N_616,N_2195);
and U9416 (N_9416,N_1559,N_3603);
and U9417 (N_9417,N_2632,N_2118);
and U9418 (N_9418,N_820,N_3514);
and U9419 (N_9419,N_3198,N_3464);
and U9420 (N_9420,N_3552,N_4166);
or U9421 (N_9421,N_2766,N_2815);
nand U9422 (N_9422,N_1118,N_2786);
xnor U9423 (N_9423,N_3057,N_4839);
nor U9424 (N_9424,N_1045,N_1494);
and U9425 (N_9425,N_41,N_1824);
or U9426 (N_9426,N_1037,N_1746);
nor U9427 (N_9427,N_2603,N_3305);
nor U9428 (N_9428,N_4826,N_1018);
nor U9429 (N_9429,N_1698,N_409);
or U9430 (N_9430,N_436,N_1719);
and U9431 (N_9431,N_4950,N_261);
nor U9432 (N_9432,N_1017,N_2758);
nand U9433 (N_9433,N_4646,N_1410);
and U9434 (N_9434,N_860,N_3142);
nand U9435 (N_9435,N_4702,N_3730);
and U9436 (N_9436,N_4179,N_4232);
and U9437 (N_9437,N_1803,N_4981);
nand U9438 (N_9438,N_2889,N_1250);
nor U9439 (N_9439,N_898,N_2956);
nor U9440 (N_9440,N_741,N_4270);
nor U9441 (N_9441,N_2269,N_262);
or U9442 (N_9442,N_3395,N_4376);
nand U9443 (N_9443,N_4562,N_1371);
xor U9444 (N_9444,N_4484,N_2783);
nand U9445 (N_9445,N_2782,N_3992);
nand U9446 (N_9446,N_291,N_3790);
nor U9447 (N_9447,N_85,N_2826);
nor U9448 (N_9448,N_1125,N_2003);
or U9449 (N_9449,N_2527,N_88);
xor U9450 (N_9450,N_4441,N_105);
and U9451 (N_9451,N_1697,N_3525);
and U9452 (N_9452,N_4509,N_505);
xor U9453 (N_9453,N_4981,N_3586);
and U9454 (N_9454,N_782,N_2207);
xor U9455 (N_9455,N_1898,N_2531);
nand U9456 (N_9456,N_4953,N_1456);
nand U9457 (N_9457,N_586,N_2790);
and U9458 (N_9458,N_284,N_1995);
or U9459 (N_9459,N_3765,N_4517);
and U9460 (N_9460,N_1027,N_235);
and U9461 (N_9461,N_3078,N_1582);
or U9462 (N_9462,N_1492,N_3628);
or U9463 (N_9463,N_804,N_2792);
and U9464 (N_9464,N_551,N_785);
and U9465 (N_9465,N_3400,N_3443);
nor U9466 (N_9466,N_3958,N_502);
xor U9467 (N_9467,N_2410,N_562);
xnor U9468 (N_9468,N_4385,N_3585);
or U9469 (N_9469,N_3699,N_4356);
nor U9470 (N_9470,N_1972,N_347);
nor U9471 (N_9471,N_2616,N_3753);
or U9472 (N_9472,N_8,N_3684);
and U9473 (N_9473,N_3843,N_738);
nand U9474 (N_9474,N_3754,N_3647);
nor U9475 (N_9475,N_1645,N_1498);
and U9476 (N_9476,N_4646,N_3812);
nand U9477 (N_9477,N_4663,N_964);
and U9478 (N_9478,N_3863,N_200);
nor U9479 (N_9479,N_2806,N_2677);
nand U9480 (N_9480,N_4109,N_772);
nor U9481 (N_9481,N_4563,N_3572);
or U9482 (N_9482,N_4591,N_566);
nand U9483 (N_9483,N_4715,N_4811);
or U9484 (N_9484,N_4146,N_1323);
or U9485 (N_9485,N_4829,N_4218);
nor U9486 (N_9486,N_1691,N_1725);
nand U9487 (N_9487,N_2362,N_4108);
xnor U9488 (N_9488,N_4077,N_50);
xnor U9489 (N_9489,N_4825,N_3398);
nor U9490 (N_9490,N_4412,N_2715);
nand U9491 (N_9491,N_4939,N_4349);
nor U9492 (N_9492,N_2471,N_1040);
or U9493 (N_9493,N_3848,N_538);
nor U9494 (N_9494,N_4411,N_3423);
nand U9495 (N_9495,N_2418,N_494);
nand U9496 (N_9496,N_627,N_24);
nand U9497 (N_9497,N_4294,N_2630);
or U9498 (N_9498,N_759,N_219);
or U9499 (N_9499,N_3388,N_704);
nor U9500 (N_9500,N_3662,N_803);
nor U9501 (N_9501,N_3516,N_4174);
or U9502 (N_9502,N_2042,N_4878);
nor U9503 (N_9503,N_4970,N_828);
nor U9504 (N_9504,N_2655,N_2757);
or U9505 (N_9505,N_4223,N_2572);
nand U9506 (N_9506,N_576,N_1322);
nor U9507 (N_9507,N_2391,N_4274);
nand U9508 (N_9508,N_4763,N_1100);
nor U9509 (N_9509,N_2212,N_3937);
nor U9510 (N_9510,N_884,N_2278);
nor U9511 (N_9511,N_3764,N_4693);
xnor U9512 (N_9512,N_802,N_2062);
nand U9513 (N_9513,N_3520,N_3224);
nand U9514 (N_9514,N_1111,N_724);
and U9515 (N_9515,N_218,N_687);
and U9516 (N_9516,N_2954,N_2945);
or U9517 (N_9517,N_4019,N_2840);
and U9518 (N_9518,N_4005,N_136);
nand U9519 (N_9519,N_3882,N_2286);
and U9520 (N_9520,N_3362,N_4016);
nor U9521 (N_9521,N_4328,N_2454);
and U9522 (N_9522,N_2005,N_489);
and U9523 (N_9523,N_3626,N_3444);
nor U9524 (N_9524,N_3095,N_1246);
and U9525 (N_9525,N_4464,N_3545);
and U9526 (N_9526,N_3172,N_1500);
nand U9527 (N_9527,N_941,N_4981);
or U9528 (N_9528,N_3440,N_4814);
xnor U9529 (N_9529,N_4917,N_1391);
and U9530 (N_9530,N_4033,N_859);
or U9531 (N_9531,N_4784,N_267);
nor U9532 (N_9532,N_2417,N_292);
nand U9533 (N_9533,N_192,N_1405);
nand U9534 (N_9534,N_1931,N_2826);
nor U9535 (N_9535,N_2329,N_449);
and U9536 (N_9536,N_2164,N_2985);
nand U9537 (N_9537,N_3982,N_2615);
nor U9538 (N_9538,N_4489,N_91);
nor U9539 (N_9539,N_4169,N_1927);
and U9540 (N_9540,N_1955,N_4814);
or U9541 (N_9541,N_796,N_3406);
xor U9542 (N_9542,N_3282,N_1067);
nand U9543 (N_9543,N_2514,N_1564);
or U9544 (N_9544,N_1631,N_1072);
or U9545 (N_9545,N_2669,N_2835);
or U9546 (N_9546,N_4302,N_4746);
or U9547 (N_9547,N_436,N_4044);
nand U9548 (N_9548,N_2538,N_1215);
and U9549 (N_9549,N_949,N_4866);
or U9550 (N_9550,N_1933,N_4405);
nand U9551 (N_9551,N_2591,N_435);
or U9552 (N_9552,N_4969,N_3494);
nand U9553 (N_9553,N_3083,N_4833);
or U9554 (N_9554,N_1530,N_4331);
nand U9555 (N_9555,N_3362,N_3708);
nor U9556 (N_9556,N_97,N_1485);
nand U9557 (N_9557,N_1301,N_2933);
or U9558 (N_9558,N_2611,N_4223);
nand U9559 (N_9559,N_51,N_4454);
or U9560 (N_9560,N_4741,N_2911);
and U9561 (N_9561,N_955,N_4488);
nand U9562 (N_9562,N_4057,N_395);
and U9563 (N_9563,N_1752,N_4381);
nand U9564 (N_9564,N_581,N_3262);
nand U9565 (N_9565,N_770,N_738);
nor U9566 (N_9566,N_4869,N_2729);
nand U9567 (N_9567,N_4945,N_1526);
nand U9568 (N_9568,N_4146,N_1504);
nor U9569 (N_9569,N_1483,N_4088);
and U9570 (N_9570,N_3142,N_575);
nand U9571 (N_9571,N_2141,N_4994);
or U9572 (N_9572,N_196,N_2446);
nor U9573 (N_9573,N_3384,N_3930);
nand U9574 (N_9574,N_1216,N_4131);
nand U9575 (N_9575,N_3762,N_3665);
or U9576 (N_9576,N_3592,N_693);
nor U9577 (N_9577,N_4504,N_11);
xnor U9578 (N_9578,N_4126,N_3574);
or U9579 (N_9579,N_2088,N_1799);
or U9580 (N_9580,N_3158,N_306);
nor U9581 (N_9581,N_1793,N_2286);
and U9582 (N_9582,N_3835,N_3737);
xor U9583 (N_9583,N_419,N_4353);
nand U9584 (N_9584,N_3427,N_604);
nor U9585 (N_9585,N_3198,N_3779);
nand U9586 (N_9586,N_3390,N_3694);
or U9587 (N_9587,N_3600,N_694);
xor U9588 (N_9588,N_2518,N_1553);
xor U9589 (N_9589,N_717,N_1046);
nand U9590 (N_9590,N_2009,N_4080);
and U9591 (N_9591,N_933,N_4196);
and U9592 (N_9592,N_2056,N_960);
nor U9593 (N_9593,N_1851,N_4298);
and U9594 (N_9594,N_1795,N_777);
xnor U9595 (N_9595,N_4937,N_2020);
and U9596 (N_9596,N_1467,N_1077);
and U9597 (N_9597,N_2865,N_4262);
or U9598 (N_9598,N_1700,N_1644);
nand U9599 (N_9599,N_430,N_205);
nand U9600 (N_9600,N_1738,N_2616);
nor U9601 (N_9601,N_4543,N_2840);
or U9602 (N_9602,N_738,N_3725);
nor U9603 (N_9603,N_344,N_2605);
or U9604 (N_9604,N_757,N_2777);
or U9605 (N_9605,N_1945,N_4043);
nand U9606 (N_9606,N_3273,N_3018);
or U9607 (N_9607,N_1759,N_3892);
nor U9608 (N_9608,N_4893,N_3440);
nor U9609 (N_9609,N_4213,N_873);
nor U9610 (N_9610,N_3350,N_3731);
xor U9611 (N_9611,N_2773,N_2079);
nor U9612 (N_9612,N_3393,N_1005);
nand U9613 (N_9613,N_4671,N_811);
nor U9614 (N_9614,N_4784,N_1064);
xor U9615 (N_9615,N_2301,N_1850);
nor U9616 (N_9616,N_1131,N_4942);
nand U9617 (N_9617,N_2342,N_3169);
nor U9618 (N_9618,N_4151,N_2681);
and U9619 (N_9619,N_3196,N_1727);
and U9620 (N_9620,N_1862,N_2788);
and U9621 (N_9621,N_1355,N_2644);
or U9622 (N_9622,N_996,N_3211);
xnor U9623 (N_9623,N_2306,N_2591);
nand U9624 (N_9624,N_953,N_629);
nor U9625 (N_9625,N_3107,N_1872);
nand U9626 (N_9626,N_3941,N_678);
xor U9627 (N_9627,N_3366,N_2623);
nand U9628 (N_9628,N_1554,N_539);
and U9629 (N_9629,N_3925,N_3807);
nand U9630 (N_9630,N_1433,N_2695);
or U9631 (N_9631,N_4150,N_4872);
nor U9632 (N_9632,N_2306,N_4993);
and U9633 (N_9633,N_3413,N_358);
and U9634 (N_9634,N_1835,N_363);
nand U9635 (N_9635,N_1500,N_2929);
or U9636 (N_9636,N_4172,N_212);
or U9637 (N_9637,N_3076,N_4860);
nand U9638 (N_9638,N_1077,N_3292);
or U9639 (N_9639,N_1417,N_547);
or U9640 (N_9640,N_3614,N_211);
nand U9641 (N_9641,N_2252,N_4109);
and U9642 (N_9642,N_3711,N_4018);
and U9643 (N_9643,N_4945,N_3481);
or U9644 (N_9644,N_1094,N_3977);
and U9645 (N_9645,N_4857,N_2098);
or U9646 (N_9646,N_657,N_1819);
and U9647 (N_9647,N_1008,N_4345);
xnor U9648 (N_9648,N_4354,N_4789);
nor U9649 (N_9649,N_3496,N_2091);
nand U9650 (N_9650,N_3971,N_112);
or U9651 (N_9651,N_4514,N_4240);
nor U9652 (N_9652,N_2686,N_2243);
and U9653 (N_9653,N_1347,N_4277);
or U9654 (N_9654,N_3390,N_3822);
or U9655 (N_9655,N_1487,N_2764);
nand U9656 (N_9656,N_883,N_1383);
and U9657 (N_9657,N_4291,N_2886);
or U9658 (N_9658,N_4067,N_1203);
nor U9659 (N_9659,N_1142,N_4955);
xnor U9660 (N_9660,N_3720,N_3823);
nand U9661 (N_9661,N_2910,N_2375);
nor U9662 (N_9662,N_718,N_3283);
and U9663 (N_9663,N_3841,N_4734);
and U9664 (N_9664,N_53,N_2650);
or U9665 (N_9665,N_4445,N_737);
and U9666 (N_9666,N_4363,N_788);
or U9667 (N_9667,N_1965,N_3256);
nand U9668 (N_9668,N_1641,N_2842);
or U9669 (N_9669,N_93,N_4027);
and U9670 (N_9670,N_2305,N_364);
and U9671 (N_9671,N_2367,N_4286);
nor U9672 (N_9672,N_4107,N_422);
and U9673 (N_9673,N_4974,N_3640);
nor U9674 (N_9674,N_2585,N_3257);
nor U9675 (N_9675,N_227,N_346);
or U9676 (N_9676,N_1868,N_1849);
or U9677 (N_9677,N_4156,N_4143);
or U9678 (N_9678,N_970,N_390);
nand U9679 (N_9679,N_4943,N_3727);
nand U9680 (N_9680,N_2225,N_2480);
or U9681 (N_9681,N_3740,N_1007);
xnor U9682 (N_9682,N_1045,N_3833);
or U9683 (N_9683,N_4594,N_2640);
xnor U9684 (N_9684,N_513,N_3401);
nand U9685 (N_9685,N_738,N_3164);
nand U9686 (N_9686,N_3772,N_2395);
or U9687 (N_9687,N_3692,N_1530);
and U9688 (N_9688,N_106,N_2230);
or U9689 (N_9689,N_4275,N_2135);
nand U9690 (N_9690,N_2611,N_4427);
nor U9691 (N_9691,N_4811,N_457);
or U9692 (N_9692,N_764,N_1919);
or U9693 (N_9693,N_1323,N_2449);
nand U9694 (N_9694,N_2412,N_3355);
nand U9695 (N_9695,N_1733,N_1165);
nand U9696 (N_9696,N_1676,N_3255);
xnor U9697 (N_9697,N_3705,N_1816);
and U9698 (N_9698,N_2691,N_3809);
and U9699 (N_9699,N_3505,N_3139);
and U9700 (N_9700,N_4296,N_1230);
nand U9701 (N_9701,N_1624,N_4803);
xnor U9702 (N_9702,N_2283,N_1065);
nor U9703 (N_9703,N_2344,N_2947);
nand U9704 (N_9704,N_2107,N_2354);
nand U9705 (N_9705,N_1131,N_4199);
nor U9706 (N_9706,N_2874,N_1029);
and U9707 (N_9707,N_3064,N_2249);
or U9708 (N_9708,N_1100,N_4824);
and U9709 (N_9709,N_3340,N_1312);
nor U9710 (N_9710,N_731,N_2020);
nor U9711 (N_9711,N_2807,N_64);
nand U9712 (N_9712,N_2814,N_2551);
or U9713 (N_9713,N_4460,N_4332);
and U9714 (N_9714,N_3544,N_3985);
xnor U9715 (N_9715,N_2434,N_3987);
or U9716 (N_9716,N_2629,N_2876);
xnor U9717 (N_9717,N_3201,N_2735);
or U9718 (N_9718,N_1698,N_197);
or U9719 (N_9719,N_591,N_3491);
nor U9720 (N_9720,N_4440,N_1687);
nor U9721 (N_9721,N_469,N_4343);
nor U9722 (N_9722,N_3850,N_2167);
nand U9723 (N_9723,N_588,N_1452);
and U9724 (N_9724,N_1121,N_26);
nor U9725 (N_9725,N_1279,N_2079);
nand U9726 (N_9726,N_2807,N_2320);
nor U9727 (N_9727,N_4749,N_1393);
and U9728 (N_9728,N_3476,N_3266);
nand U9729 (N_9729,N_1844,N_699);
nand U9730 (N_9730,N_502,N_4498);
nand U9731 (N_9731,N_2182,N_4147);
and U9732 (N_9732,N_126,N_1889);
nor U9733 (N_9733,N_1825,N_259);
nand U9734 (N_9734,N_3693,N_1810);
xnor U9735 (N_9735,N_1546,N_2831);
xor U9736 (N_9736,N_3676,N_417);
nand U9737 (N_9737,N_1486,N_1890);
or U9738 (N_9738,N_471,N_1464);
nor U9739 (N_9739,N_4956,N_3223);
or U9740 (N_9740,N_3359,N_1692);
nor U9741 (N_9741,N_2262,N_277);
or U9742 (N_9742,N_4444,N_4620);
nor U9743 (N_9743,N_512,N_3702);
nand U9744 (N_9744,N_2210,N_2732);
nand U9745 (N_9745,N_878,N_3152);
nand U9746 (N_9746,N_3904,N_3149);
nand U9747 (N_9747,N_495,N_875);
nand U9748 (N_9748,N_4487,N_1351);
or U9749 (N_9749,N_2563,N_158);
and U9750 (N_9750,N_4114,N_3890);
and U9751 (N_9751,N_1115,N_2373);
xor U9752 (N_9752,N_4662,N_3862);
nand U9753 (N_9753,N_3141,N_3302);
nor U9754 (N_9754,N_4489,N_4003);
nand U9755 (N_9755,N_4561,N_314);
nand U9756 (N_9756,N_2417,N_3442);
or U9757 (N_9757,N_4200,N_658);
nor U9758 (N_9758,N_1908,N_3592);
and U9759 (N_9759,N_2897,N_2658);
and U9760 (N_9760,N_1592,N_4753);
or U9761 (N_9761,N_644,N_3788);
and U9762 (N_9762,N_1384,N_3860);
or U9763 (N_9763,N_2805,N_1056);
nor U9764 (N_9764,N_621,N_2184);
and U9765 (N_9765,N_4486,N_519);
nand U9766 (N_9766,N_1835,N_3167);
nor U9767 (N_9767,N_4839,N_4045);
or U9768 (N_9768,N_3149,N_3950);
xnor U9769 (N_9769,N_4006,N_4283);
and U9770 (N_9770,N_235,N_3592);
or U9771 (N_9771,N_707,N_2993);
and U9772 (N_9772,N_3213,N_3889);
and U9773 (N_9773,N_654,N_4516);
nand U9774 (N_9774,N_919,N_4263);
xnor U9775 (N_9775,N_3174,N_3710);
nor U9776 (N_9776,N_3683,N_415);
or U9777 (N_9777,N_3337,N_3254);
or U9778 (N_9778,N_1894,N_4909);
and U9779 (N_9779,N_267,N_735);
and U9780 (N_9780,N_1383,N_3988);
and U9781 (N_9781,N_1003,N_3233);
or U9782 (N_9782,N_69,N_2884);
nand U9783 (N_9783,N_665,N_2760);
and U9784 (N_9784,N_3858,N_2847);
or U9785 (N_9785,N_4381,N_690);
nor U9786 (N_9786,N_914,N_4953);
and U9787 (N_9787,N_4661,N_3634);
or U9788 (N_9788,N_3586,N_202);
or U9789 (N_9789,N_2562,N_1064);
or U9790 (N_9790,N_2345,N_4239);
nand U9791 (N_9791,N_2027,N_4859);
or U9792 (N_9792,N_72,N_2669);
and U9793 (N_9793,N_3008,N_3014);
and U9794 (N_9794,N_2734,N_2062);
nand U9795 (N_9795,N_3917,N_2220);
and U9796 (N_9796,N_3171,N_1501);
and U9797 (N_9797,N_488,N_4464);
nand U9798 (N_9798,N_2476,N_947);
and U9799 (N_9799,N_2874,N_3315);
or U9800 (N_9800,N_1576,N_1077);
nor U9801 (N_9801,N_404,N_2303);
or U9802 (N_9802,N_3580,N_1159);
nor U9803 (N_9803,N_81,N_2507);
nor U9804 (N_9804,N_1578,N_3996);
nor U9805 (N_9805,N_531,N_2743);
nor U9806 (N_9806,N_857,N_2768);
and U9807 (N_9807,N_2458,N_3524);
nand U9808 (N_9808,N_1059,N_939);
nand U9809 (N_9809,N_3682,N_2115);
and U9810 (N_9810,N_3048,N_2951);
nand U9811 (N_9811,N_4893,N_3852);
or U9812 (N_9812,N_191,N_2227);
nand U9813 (N_9813,N_1096,N_2981);
xor U9814 (N_9814,N_3833,N_3350);
nand U9815 (N_9815,N_2634,N_4681);
and U9816 (N_9816,N_1466,N_3234);
nor U9817 (N_9817,N_773,N_1418);
nand U9818 (N_9818,N_33,N_4640);
nand U9819 (N_9819,N_1043,N_1646);
nand U9820 (N_9820,N_1208,N_1489);
nor U9821 (N_9821,N_4820,N_3163);
or U9822 (N_9822,N_1644,N_3808);
or U9823 (N_9823,N_3119,N_42);
or U9824 (N_9824,N_4352,N_2321);
or U9825 (N_9825,N_1538,N_3917);
and U9826 (N_9826,N_1735,N_3747);
and U9827 (N_9827,N_4639,N_789);
nor U9828 (N_9828,N_4665,N_3875);
and U9829 (N_9829,N_4082,N_3883);
and U9830 (N_9830,N_647,N_4556);
and U9831 (N_9831,N_1786,N_4252);
and U9832 (N_9832,N_4082,N_2296);
or U9833 (N_9833,N_254,N_2704);
nand U9834 (N_9834,N_4372,N_511);
or U9835 (N_9835,N_1714,N_4555);
or U9836 (N_9836,N_16,N_760);
nand U9837 (N_9837,N_283,N_4659);
or U9838 (N_9838,N_4799,N_2524);
and U9839 (N_9839,N_1765,N_1798);
nor U9840 (N_9840,N_2500,N_3875);
and U9841 (N_9841,N_1176,N_1385);
or U9842 (N_9842,N_592,N_1496);
nor U9843 (N_9843,N_478,N_3635);
and U9844 (N_9844,N_869,N_783);
or U9845 (N_9845,N_4673,N_2382);
or U9846 (N_9846,N_1341,N_571);
xor U9847 (N_9847,N_4772,N_2465);
nor U9848 (N_9848,N_921,N_1777);
nor U9849 (N_9849,N_2084,N_3571);
or U9850 (N_9850,N_2183,N_110);
or U9851 (N_9851,N_4043,N_105);
nor U9852 (N_9852,N_3224,N_1959);
and U9853 (N_9853,N_4668,N_3798);
or U9854 (N_9854,N_2041,N_3236);
or U9855 (N_9855,N_5,N_3165);
nor U9856 (N_9856,N_2391,N_144);
and U9857 (N_9857,N_4163,N_538);
nor U9858 (N_9858,N_4967,N_4228);
xor U9859 (N_9859,N_1190,N_693);
and U9860 (N_9860,N_2616,N_3778);
nand U9861 (N_9861,N_4255,N_3742);
xnor U9862 (N_9862,N_297,N_3540);
or U9863 (N_9863,N_3586,N_2313);
nand U9864 (N_9864,N_4142,N_4010);
nor U9865 (N_9865,N_1958,N_662);
xnor U9866 (N_9866,N_1239,N_1244);
and U9867 (N_9867,N_933,N_261);
and U9868 (N_9868,N_2026,N_4354);
and U9869 (N_9869,N_2419,N_756);
and U9870 (N_9870,N_1107,N_3389);
nand U9871 (N_9871,N_1321,N_2302);
xor U9872 (N_9872,N_2503,N_224);
nand U9873 (N_9873,N_4638,N_3001);
nor U9874 (N_9874,N_1109,N_1301);
nand U9875 (N_9875,N_2943,N_1398);
nand U9876 (N_9876,N_375,N_902);
nand U9877 (N_9877,N_2355,N_269);
or U9878 (N_9878,N_2823,N_2652);
nand U9879 (N_9879,N_3024,N_3306);
nand U9880 (N_9880,N_2089,N_4044);
and U9881 (N_9881,N_2919,N_783);
nand U9882 (N_9882,N_4651,N_3842);
nor U9883 (N_9883,N_3219,N_244);
nor U9884 (N_9884,N_392,N_2499);
nor U9885 (N_9885,N_3901,N_4394);
nor U9886 (N_9886,N_3843,N_108);
nor U9887 (N_9887,N_215,N_4534);
nand U9888 (N_9888,N_1134,N_3936);
or U9889 (N_9889,N_1880,N_1534);
and U9890 (N_9890,N_3197,N_1102);
or U9891 (N_9891,N_4708,N_4569);
nor U9892 (N_9892,N_2462,N_4790);
nand U9893 (N_9893,N_179,N_2400);
and U9894 (N_9894,N_3020,N_3012);
nand U9895 (N_9895,N_4089,N_1551);
nand U9896 (N_9896,N_798,N_1620);
and U9897 (N_9897,N_3696,N_4702);
nand U9898 (N_9898,N_3113,N_4756);
xor U9899 (N_9899,N_2121,N_3934);
xnor U9900 (N_9900,N_3453,N_3493);
xnor U9901 (N_9901,N_1357,N_4311);
or U9902 (N_9902,N_684,N_4560);
nor U9903 (N_9903,N_153,N_3814);
nor U9904 (N_9904,N_2013,N_2029);
or U9905 (N_9905,N_1550,N_1414);
nor U9906 (N_9906,N_2785,N_1129);
xnor U9907 (N_9907,N_2412,N_987);
or U9908 (N_9908,N_4930,N_352);
and U9909 (N_9909,N_3233,N_1137);
or U9910 (N_9910,N_598,N_2764);
nor U9911 (N_9911,N_4292,N_4969);
and U9912 (N_9912,N_2268,N_262);
nor U9913 (N_9913,N_1897,N_4397);
nor U9914 (N_9914,N_4997,N_2631);
or U9915 (N_9915,N_3036,N_705);
and U9916 (N_9916,N_545,N_3281);
and U9917 (N_9917,N_1171,N_1733);
or U9918 (N_9918,N_1035,N_4352);
nor U9919 (N_9919,N_2907,N_1446);
nand U9920 (N_9920,N_614,N_2818);
nand U9921 (N_9921,N_2423,N_1432);
nor U9922 (N_9922,N_3643,N_776);
or U9923 (N_9923,N_828,N_1155);
and U9924 (N_9924,N_1488,N_764);
xnor U9925 (N_9925,N_1296,N_4309);
and U9926 (N_9926,N_4508,N_4107);
nor U9927 (N_9927,N_2666,N_70);
nand U9928 (N_9928,N_1639,N_3691);
or U9929 (N_9929,N_525,N_1161);
nand U9930 (N_9930,N_314,N_4147);
nand U9931 (N_9931,N_1133,N_1475);
nor U9932 (N_9932,N_442,N_130);
and U9933 (N_9933,N_2672,N_4382);
nor U9934 (N_9934,N_838,N_2216);
nor U9935 (N_9935,N_1116,N_2789);
and U9936 (N_9936,N_4540,N_2534);
nor U9937 (N_9937,N_3388,N_230);
and U9938 (N_9938,N_2292,N_934);
nand U9939 (N_9939,N_4054,N_3904);
xor U9940 (N_9940,N_4040,N_1405);
and U9941 (N_9941,N_1145,N_1940);
nand U9942 (N_9942,N_956,N_2352);
or U9943 (N_9943,N_4245,N_1152);
or U9944 (N_9944,N_1327,N_525);
nor U9945 (N_9945,N_3114,N_18);
nand U9946 (N_9946,N_3182,N_1679);
nor U9947 (N_9947,N_2399,N_3654);
or U9948 (N_9948,N_4421,N_216);
and U9949 (N_9949,N_2696,N_1432);
nand U9950 (N_9950,N_172,N_4007);
and U9951 (N_9951,N_3405,N_987);
nand U9952 (N_9952,N_1017,N_154);
and U9953 (N_9953,N_1402,N_1359);
or U9954 (N_9954,N_1972,N_809);
nor U9955 (N_9955,N_856,N_4258);
or U9956 (N_9956,N_718,N_4263);
and U9957 (N_9957,N_4296,N_1166);
or U9958 (N_9958,N_4469,N_1776);
and U9959 (N_9959,N_4788,N_4158);
nand U9960 (N_9960,N_1268,N_3143);
nor U9961 (N_9961,N_4653,N_1084);
nand U9962 (N_9962,N_365,N_1171);
or U9963 (N_9963,N_1409,N_1916);
nor U9964 (N_9964,N_1344,N_1955);
and U9965 (N_9965,N_1105,N_3913);
nand U9966 (N_9966,N_3715,N_328);
and U9967 (N_9967,N_832,N_3441);
nand U9968 (N_9968,N_1170,N_4780);
or U9969 (N_9969,N_3603,N_4313);
nand U9970 (N_9970,N_2103,N_53);
and U9971 (N_9971,N_4678,N_2451);
nor U9972 (N_9972,N_3993,N_53);
and U9973 (N_9973,N_2270,N_3121);
nor U9974 (N_9974,N_2804,N_4156);
or U9975 (N_9975,N_4388,N_1356);
nor U9976 (N_9976,N_3879,N_4742);
and U9977 (N_9977,N_1712,N_2618);
and U9978 (N_9978,N_4561,N_1974);
nand U9979 (N_9979,N_4759,N_4967);
xnor U9980 (N_9980,N_4630,N_4981);
nand U9981 (N_9981,N_3266,N_1905);
nand U9982 (N_9982,N_4402,N_4876);
or U9983 (N_9983,N_2452,N_3289);
and U9984 (N_9984,N_4625,N_1010);
nor U9985 (N_9985,N_1868,N_1493);
xnor U9986 (N_9986,N_2328,N_66);
nand U9987 (N_9987,N_4574,N_4362);
nor U9988 (N_9988,N_3833,N_4042);
xor U9989 (N_9989,N_4095,N_4289);
nand U9990 (N_9990,N_93,N_3052);
nor U9991 (N_9991,N_4318,N_4835);
or U9992 (N_9992,N_1886,N_4553);
nand U9993 (N_9993,N_4348,N_3332);
or U9994 (N_9994,N_2457,N_4052);
nand U9995 (N_9995,N_2398,N_2380);
nand U9996 (N_9996,N_1258,N_1285);
nand U9997 (N_9997,N_2689,N_2446);
nand U9998 (N_9998,N_2968,N_435);
nand U9999 (N_9999,N_4978,N_2);
xor U10000 (N_10000,N_6651,N_5673);
and U10001 (N_10001,N_5560,N_8871);
nand U10002 (N_10002,N_5979,N_7663);
nor U10003 (N_10003,N_7732,N_5398);
nand U10004 (N_10004,N_6203,N_5940);
and U10005 (N_10005,N_5162,N_5920);
nor U10006 (N_10006,N_7064,N_5137);
and U10007 (N_10007,N_8859,N_7394);
and U10008 (N_10008,N_5619,N_8266);
or U10009 (N_10009,N_8002,N_7504);
and U10010 (N_10010,N_7983,N_8431);
nor U10011 (N_10011,N_5810,N_8020);
nand U10012 (N_10012,N_7517,N_6570);
and U10013 (N_10013,N_8535,N_5428);
nand U10014 (N_10014,N_6787,N_8417);
nor U10015 (N_10015,N_9496,N_9128);
xnor U10016 (N_10016,N_6033,N_8425);
nand U10017 (N_10017,N_7414,N_8962);
or U10018 (N_10018,N_5842,N_9426);
and U10019 (N_10019,N_5366,N_6726);
xnor U10020 (N_10020,N_9117,N_8361);
nor U10021 (N_10021,N_5678,N_6015);
or U10022 (N_10022,N_6069,N_7440);
xor U10023 (N_10023,N_5070,N_7799);
and U10024 (N_10024,N_6409,N_8124);
nand U10025 (N_10025,N_6902,N_9202);
xor U10026 (N_10026,N_9382,N_8900);
and U10027 (N_10027,N_7933,N_7914);
and U10028 (N_10028,N_8059,N_8125);
xnor U10029 (N_10029,N_7744,N_5613);
and U10030 (N_10030,N_8147,N_5958);
nand U10031 (N_10031,N_8148,N_8809);
and U10032 (N_10032,N_6245,N_7409);
or U10033 (N_10033,N_5515,N_9990);
and U10034 (N_10034,N_8830,N_5983);
and U10035 (N_10035,N_7727,N_6893);
nand U10036 (N_10036,N_5306,N_6950);
nor U10037 (N_10037,N_6866,N_5074);
nand U10038 (N_10038,N_9639,N_8617);
nor U10039 (N_10039,N_6420,N_6675);
nand U10040 (N_10040,N_6102,N_8380);
and U10041 (N_10041,N_9361,N_8468);
nand U10042 (N_10042,N_7925,N_8267);
or U10043 (N_10043,N_9675,N_9800);
nand U10044 (N_10044,N_6290,N_6062);
nor U10045 (N_10045,N_6418,N_8390);
nor U10046 (N_10046,N_7157,N_9122);
nand U10047 (N_10047,N_9616,N_5537);
and U10048 (N_10048,N_9353,N_9478);
and U10049 (N_10049,N_9648,N_8221);
or U10050 (N_10050,N_5874,N_7619);
or U10051 (N_10051,N_9060,N_6775);
nor U10052 (N_10052,N_6309,N_6227);
nand U10053 (N_10053,N_5575,N_5125);
and U10054 (N_10054,N_8430,N_8365);
and U10055 (N_10055,N_9347,N_8190);
nor U10056 (N_10056,N_8415,N_7491);
nand U10057 (N_10057,N_5655,N_9785);
and U10058 (N_10058,N_8207,N_8941);
and U10059 (N_10059,N_8455,N_9723);
and U10060 (N_10060,N_5670,N_6984);
xnor U10061 (N_10061,N_6337,N_6006);
xnor U10062 (N_10062,N_8352,N_7588);
xnor U10063 (N_10063,N_9217,N_6987);
nor U10064 (N_10064,N_9106,N_5139);
nor U10065 (N_10065,N_9484,N_6286);
or U10066 (N_10066,N_8860,N_5669);
or U10067 (N_10067,N_7523,N_7314);
nor U10068 (N_10068,N_6876,N_7907);
xor U10069 (N_10069,N_6164,N_5975);
and U10070 (N_10070,N_5078,N_5486);
or U10071 (N_10071,N_9645,N_8853);
xnor U10072 (N_10072,N_7735,N_9579);
nand U10073 (N_10073,N_6345,N_7185);
or U10074 (N_10074,N_8399,N_5335);
or U10075 (N_10075,N_6129,N_9195);
nor U10076 (N_10076,N_8142,N_9190);
nand U10077 (N_10077,N_5760,N_5020);
or U10078 (N_10078,N_9621,N_7029);
nand U10079 (N_10079,N_8780,N_7250);
and U10080 (N_10080,N_5587,N_6177);
xnor U10081 (N_10081,N_8915,N_7834);
xor U10082 (N_10082,N_7980,N_7860);
nand U10083 (N_10083,N_8721,N_8533);
and U10084 (N_10084,N_6378,N_6222);
nand U10085 (N_10085,N_5511,N_8566);
nand U10086 (N_10086,N_6784,N_6603);
nor U10087 (N_10087,N_9370,N_9201);
nand U10088 (N_10088,N_8400,N_7711);
or U10089 (N_10089,N_5068,N_9010);
or U10090 (N_10090,N_6248,N_8748);
nor U10091 (N_10091,N_9330,N_8593);
nand U10092 (N_10092,N_5865,N_5329);
and U10093 (N_10093,N_7658,N_7515);
and U10094 (N_10094,N_9769,N_6920);
and U10095 (N_10095,N_6824,N_9524);
or U10096 (N_10096,N_7994,N_6528);
and U10097 (N_10097,N_9149,N_7263);
and U10098 (N_10098,N_9164,N_7003);
or U10099 (N_10099,N_9869,N_5939);
nand U10100 (N_10100,N_9047,N_5835);
or U10101 (N_10101,N_5437,N_7922);
nand U10102 (N_10102,N_6729,N_7345);
nand U10103 (N_10103,N_7981,N_6904);
nand U10104 (N_10104,N_8310,N_8713);
or U10105 (N_10105,N_7573,N_5585);
nand U10106 (N_10106,N_5463,N_5418);
or U10107 (N_10107,N_5941,N_9981);
or U10108 (N_10108,N_5572,N_5854);
xor U10109 (N_10109,N_6773,N_6441);
nand U10110 (N_10110,N_6398,N_6255);
or U10111 (N_10111,N_5396,N_7717);
xnor U10112 (N_10112,N_9389,N_8539);
or U10113 (N_10113,N_5342,N_7646);
or U10114 (N_10114,N_6184,N_8594);
or U10115 (N_10115,N_7698,N_9980);
nor U10116 (N_10116,N_8225,N_7818);
nand U10117 (N_10117,N_7264,N_5925);
or U10118 (N_10118,N_6009,N_6611);
and U10119 (N_10119,N_8543,N_9792);
and U10120 (N_10120,N_9181,N_6044);
and U10121 (N_10121,N_6746,N_7301);
and U10122 (N_10122,N_6445,N_9740);
nand U10123 (N_10123,N_8739,N_7328);
or U10124 (N_10124,N_9635,N_5741);
or U10125 (N_10125,N_5151,N_7316);
or U10126 (N_10126,N_6846,N_5974);
or U10127 (N_10127,N_7387,N_9861);
xor U10128 (N_10128,N_6148,N_7742);
nand U10129 (N_10129,N_8297,N_5972);
or U10130 (N_10130,N_5258,N_8832);
and U10131 (N_10131,N_9345,N_9231);
and U10132 (N_10132,N_8628,N_7303);
or U10133 (N_10133,N_8326,N_8169);
and U10134 (N_10134,N_7889,N_5318);
nor U10135 (N_10135,N_8796,N_5438);
nor U10136 (N_10136,N_8107,N_8498);
nor U10137 (N_10137,N_6186,N_9337);
and U10138 (N_10138,N_9246,N_8086);
and U10139 (N_10139,N_8677,N_8931);
and U10140 (N_10140,N_6406,N_6559);
nand U10141 (N_10141,N_5429,N_8171);
xor U10142 (N_10142,N_9995,N_7976);
xnor U10143 (N_10143,N_6656,N_7299);
and U10144 (N_10144,N_8000,N_6568);
or U10145 (N_10145,N_8482,N_6986);
nand U10146 (N_10146,N_6300,N_5028);
and U10147 (N_10147,N_5172,N_6483);
or U10148 (N_10148,N_5197,N_9743);
nand U10149 (N_10149,N_5032,N_9768);
nand U10150 (N_10150,N_9071,N_7516);
nor U10151 (N_10151,N_7298,N_5853);
and U10152 (N_10152,N_7965,N_6548);
xor U10153 (N_10153,N_7770,N_6356);
nand U10154 (N_10154,N_9433,N_8973);
and U10155 (N_10155,N_5589,N_6688);
nor U10156 (N_10156,N_6967,N_7974);
nor U10157 (N_10157,N_9462,N_9022);
nor U10158 (N_10158,N_7804,N_5959);
nor U10159 (N_10159,N_5998,N_5986);
nor U10160 (N_10160,N_6502,N_9958);
and U10161 (N_10161,N_9984,N_9797);
and U10162 (N_10162,N_6679,N_9256);
or U10163 (N_10163,N_5698,N_5803);
and U10164 (N_10164,N_6229,N_6217);
and U10165 (N_10165,N_6320,N_5757);
nor U10166 (N_10166,N_5790,N_6435);
nor U10167 (N_10167,N_7542,N_9511);
nand U10168 (N_10168,N_7119,N_5002);
or U10169 (N_10169,N_6993,N_6505);
nand U10170 (N_10170,N_7112,N_6175);
xnor U10171 (N_10171,N_9843,N_8131);
nor U10172 (N_10172,N_7026,N_9271);
and U10173 (N_10173,N_8737,N_5241);
nor U10174 (N_10174,N_8876,N_7603);
nor U10175 (N_10175,N_6094,N_7370);
xor U10176 (N_10176,N_5521,N_8693);
nand U10177 (N_10177,N_8986,N_9001);
or U10178 (N_10178,N_8090,N_5245);
nand U10179 (N_10179,N_7346,N_6192);
or U10180 (N_10180,N_5733,N_8626);
nor U10181 (N_10181,N_7247,N_7783);
or U10182 (N_10182,N_7478,N_5194);
and U10183 (N_10183,N_8551,N_5365);
or U10184 (N_10184,N_8449,N_7775);
and U10185 (N_10185,N_9957,N_5007);
nor U10186 (N_10186,N_8157,N_5155);
and U10187 (N_10187,N_7617,N_7940);
nand U10188 (N_10188,N_8492,N_9825);
or U10189 (N_10189,N_5409,N_9114);
or U10190 (N_10190,N_7463,N_5580);
nor U10191 (N_10191,N_5562,N_8298);
and U10192 (N_10192,N_8908,N_5203);
nand U10193 (N_10193,N_7023,N_7849);
nand U10194 (N_10194,N_9727,N_8133);
or U10195 (N_10195,N_9362,N_7715);
nand U10196 (N_10196,N_8862,N_6718);
and U10197 (N_10197,N_9120,N_8282);
or U10198 (N_10198,N_9220,N_8254);
and U10199 (N_10199,N_5136,N_6820);
nor U10200 (N_10200,N_9576,N_8681);
nand U10201 (N_10201,N_7237,N_6292);
and U10202 (N_10202,N_9987,N_6312);
or U10203 (N_10203,N_8103,N_5981);
or U10204 (N_10204,N_7363,N_9240);
or U10205 (N_10205,N_6975,N_8052);
nand U10206 (N_10206,N_7074,N_6293);
or U10207 (N_10207,N_6220,N_6176);
xor U10208 (N_10208,N_6779,N_8630);
or U10209 (N_10209,N_8706,N_7612);
nand U10210 (N_10210,N_5071,N_9365);
nor U10211 (N_10211,N_8443,N_9724);
nor U10212 (N_10212,N_7969,N_5937);
nor U10213 (N_10213,N_6317,N_8005);
nor U10214 (N_10214,N_7146,N_8318);
nor U10215 (N_10215,N_6683,N_9831);
nand U10216 (N_10216,N_8027,N_5262);
or U10217 (N_10217,N_6953,N_6349);
and U10218 (N_10218,N_7359,N_9399);
or U10219 (N_10219,N_5130,N_6289);
nor U10220 (N_10220,N_7281,N_6010);
nor U10221 (N_10221,N_6396,N_7168);
nand U10222 (N_10222,N_9857,N_6829);
nor U10223 (N_10223,N_7189,N_8026);
nor U10224 (N_10224,N_7641,N_5341);
nand U10225 (N_10225,N_8822,N_6952);
nand U10226 (N_10226,N_6689,N_5085);
nand U10227 (N_10227,N_7134,N_5378);
nand U10228 (N_10228,N_7145,N_8684);
or U10229 (N_10229,N_9998,N_5484);
or U10230 (N_10230,N_7309,N_6673);
nor U10231 (N_10231,N_6374,N_7561);
nor U10232 (N_10232,N_7737,N_9186);
and U10233 (N_10233,N_5199,N_5031);
nand U10234 (N_10234,N_7423,N_5173);
nor U10235 (N_10235,N_5561,N_9448);
nor U10236 (N_10236,N_6985,N_6257);
or U10237 (N_10237,N_6545,N_6926);
nor U10238 (N_10238,N_8374,N_7874);
or U10239 (N_10239,N_6209,N_9821);
nand U10240 (N_10240,N_5758,N_9782);
xnor U10241 (N_10241,N_9111,N_5891);
nand U10242 (N_10242,N_6159,N_8178);
or U10243 (N_10243,N_7798,N_6226);
nor U10244 (N_10244,N_6947,N_8401);
nor U10245 (N_10245,N_8159,N_7691);
nand U10246 (N_10246,N_8838,N_9539);
or U10247 (N_10247,N_9683,N_6024);
nand U10248 (N_10248,N_9127,N_6249);
or U10249 (N_10249,N_8306,N_8510);
and U10250 (N_10250,N_9809,N_8534);
and U10251 (N_10251,N_6230,N_8726);
nand U10252 (N_10252,N_8958,N_8666);
nor U10253 (N_10253,N_7405,N_8553);
or U10254 (N_10254,N_7792,N_9307);
nor U10255 (N_10255,N_9783,N_8152);
nand U10256 (N_10256,N_5022,N_8453);
nor U10257 (N_10257,N_7091,N_9679);
nor U10258 (N_10258,N_8343,N_8968);
and U10259 (N_10259,N_5610,N_8727);
and U10260 (N_10260,N_8951,N_7081);
nor U10261 (N_10261,N_7248,N_7623);
nand U10262 (N_10262,N_9214,N_7817);
nor U10263 (N_10263,N_5179,N_6654);
nand U10264 (N_10264,N_6500,N_8409);
or U10265 (N_10265,N_8228,N_8555);
nand U10266 (N_10266,N_6691,N_6650);
or U10267 (N_10267,N_9184,N_9508);
or U10268 (N_10268,N_9881,N_9044);
and U10269 (N_10269,N_7886,N_5174);
nor U10270 (N_10270,N_9827,N_5631);
and U10271 (N_10271,N_9529,N_5750);
nand U10272 (N_10272,N_8004,N_9932);
nor U10273 (N_10273,N_8237,N_5186);
nor U10274 (N_10274,N_7195,N_5475);
or U10275 (N_10275,N_6279,N_9767);
xor U10276 (N_10276,N_5200,N_7092);
nor U10277 (N_10277,N_8489,N_7225);
and U10278 (N_10278,N_7100,N_5767);
nor U10279 (N_10279,N_6138,N_8154);
nand U10280 (N_10280,N_5577,N_6327);
nor U10281 (N_10281,N_9025,N_5259);
nand U10282 (N_10282,N_7055,N_9589);
nand U10283 (N_10283,N_9215,N_9053);
xnor U10284 (N_10284,N_5065,N_8682);
xor U10285 (N_10285,N_9334,N_8299);
nand U10286 (N_10286,N_5873,N_5114);
nand U10287 (N_10287,N_8919,N_7272);
nor U10288 (N_10288,N_7764,N_7106);
nand U10289 (N_10289,N_9130,N_7004);
nor U10290 (N_10290,N_6633,N_9725);
nor U10291 (N_10291,N_8511,N_6273);
nand U10292 (N_10292,N_7174,N_5805);
and U10293 (N_10293,N_6411,N_9213);
and U10294 (N_10294,N_7318,N_6881);
nand U10295 (N_10295,N_5745,N_6328);
and U10296 (N_10296,N_8637,N_5158);
and U10297 (N_10297,N_6826,N_8045);
nor U10298 (N_10298,N_6897,N_8526);
nor U10299 (N_10299,N_6468,N_7388);
nor U10300 (N_10300,N_8011,N_8912);
or U10301 (N_10301,N_8802,N_7001);
or U10302 (N_10302,N_6088,N_9608);
or U10303 (N_10303,N_7321,N_5879);
or U10304 (N_10304,N_7752,N_8634);
xnor U10305 (N_10305,N_9855,N_8261);
nand U10306 (N_10306,N_5599,N_8913);
xor U10307 (N_10307,N_9832,N_8143);
and U10308 (N_10308,N_6520,N_7570);
or U10309 (N_10309,N_5381,N_7453);
and U10310 (N_10310,N_7203,N_7209);
xor U10311 (N_10311,N_7104,N_6607);
nor U10312 (N_10312,N_6433,N_9810);
xor U10313 (N_10313,N_6386,N_6901);
nand U10314 (N_10314,N_9077,N_9729);
nand U10315 (N_10315,N_6955,N_9878);
or U10316 (N_10316,N_6613,N_5037);
or U10317 (N_10317,N_9139,N_7011);
nor U10318 (N_10318,N_5944,N_6804);
or U10319 (N_10319,N_8121,N_6208);
nor U10320 (N_10320,N_5731,N_5243);
or U10321 (N_10321,N_7261,N_5233);
nand U10322 (N_10322,N_7945,N_6614);
or U10323 (N_10323,N_8692,N_5993);
or U10324 (N_10324,N_7111,N_5824);
or U10325 (N_10325,N_8928,N_7354);
xnor U10326 (N_10326,N_9983,N_5509);
and U10327 (N_10327,N_6032,N_9269);
xor U10328 (N_10328,N_5392,N_9449);
or U10329 (N_10329,N_8970,N_6862);
nand U10330 (N_10330,N_8377,N_8246);
nor U10331 (N_10331,N_5863,N_5569);
xnor U10332 (N_10332,N_7322,N_9336);
nor U10333 (N_10333,N_6686,N_7009);
and U10334 (N_10334,N_6809,N_6096);
nor U10335 (N_10335,N_8975,N_9419);
and U10336 (N_10336,N_7544,N_5749);
nor U10337 (N_10337,N_7957,N_6627);
xor U10338 (N_10338,N_9793,N_5473);
or U10339 (N_10339,N_6912,N_8477);
and U10340 (N_10340,N_6270,N_6593);
or U10341 (N_10341,N_6900,N_9302);
nand U10342 (N_10342,N_6153,N_9751);
nor U10343 (N_10343,N_7633,N_6670);
nor U10344 (N_10344,N_8939,N_9989);
nor U10345 (N_10345,N_7049,N_6456);
and U10346 (N_10346,N_7788,N_5650);
nor U10347 (N_10347,N_5798,N_5783);
and U10348 (N_10348,N_5080,N_5751);
or U10349 (N_10349,N_6000,N_8158);
and U10350 (N_10350,N_5132,N_7873);
nor U10351 (N_10351,N_9663,N_5956);
nor U10352 (N_10352,N_5701,N_8797);
nand U10353 (N_10353,N_6535,N_6158);
or U10354 (N_10354,N_8836,N_6080);
nand U10355 (N_10355,N_9016,N_6313);
nor U10356 (N_10356,N_9252,N_9844);
or U10357 (N_10357,N_9297,N_5311);
nor U10358 (N_10358,N_6195,N_7724);
xnor U10359 (N_10359,N_5642,N_6421);
and U10360 (N_10360,N_6664,N_6423);
and U10361 (N_10361,N_7996,N_5025);
or U10362 (N_10362,N_9379,N_5682);
or U10363 (N_10363,N_5355,N_6905);
nand U10364 (N_10364,N_9046,N_7319);
and U10365 (N_10365,N_9673,N_5044);
nand U10366 (N_10366,N_9943,N_9391);
or U10367 (N_10367,N_9378,N_7769);
and U10368 (N_10368,N_6348,N_7270);
nand U10369 (N_10369,N_6855,N_8742);
xnor U10370 (N_10370,N_9094,N_7707);
and U10371 (N_10371,N_8439,N_7459);
and U10372 (N_10372,N_5838,N_8683);
or U10373 (N_10373,N_7694,N_8123);
and U10374 (N_10374,N_8203,N_6049);
nor U10375 (N_10375,N_7396,N_8396);
nand U10376 (N_10376,N_7404,N_7142);
nand U10377 (N_10377,N_7509,N_8979);
nor U10378 (N_10378,N_9546,N_6547);
nand U10379 (N_10379,N_5076,N_7918);
or U10380 (N_10380,N_5296,N_5104);
or U10381 (N_10381,N_5960,N_7729);
or U10382 (N_10382,N_9210,N_7390);
nand U10383 (N_10383,N_9075,N_7946);
and U10384 (N_10384,N_8213,N_8955);
and U10385 (N_10385,N_7560,N_8173);
or U10386 (N_10386,N_5982,N_9002);
or U10387 (N_10387,N_7436,N_7128);
or U10388 (N_10388,N_6193,N_5964);
or U10389 (N_10389,N_9418,N_9474);
or U10390 (N_10390,N_6287,N_5639);
or U10391 (N_10391,N_6324,N_6853);
and U10392 (N_10392,N_9351,N_7073);
and U10393 (N_10393,N_9909,N_8281);
nand U10394 (N_10394,N_6163,N_8785);
or U10395 (N_10395,N_6916,N_9520);
and U10396 (N_10396,N_5553,N_5953);
or U10397 (N_10397,N_6600,N_7018);
nand U10398 (N_10398,N_7317,N_9410);
nand U10399 (N_10399,N_6026,N_5083);
nor U10400 (N_10400,N_5752,N_8812);
or U10401 (N_10401,N_7503,N_8226);
nand U10402 (N_10402,N_5229,N_6021);
nor U10403 (N_10403,N_6361,N_6243);
xnor U10404 (N_10404,N_8050,N_7094);
or U10405 (N_10405,N_6971,N_5544);
nor U10406 (N_10406,N_5344,N_7524);
nand U10407 (N_10407,N_8927,N_9574);
and U10408 (N_10408,N_9678,N_5985);
and U10409 (N_10409,N_9339,N_7852);
nor U10410 (N_10410,N_5322,N_8884);
nor U10411 (N_10411,N_8701,N_8337);
nand U10412 (N_10412,N_8088,N_5009);
nor U10413 (N_10413,N_9052,N_6860);
nand U10414 (N_10414,N_9865,N_6384);
nor U10415 (N_10415,N_5713,N_6206);
nand U10416 (N_10416,N_5176,N_9008);
nand U10417 (N_10417,N_5178,N_5019);
xnor U10418 (N_10418,N_5570,N_9477);
nor U10419 (N_10419,N_5620,N_7496);
nor U10420 (N_10420,N_5274,N_6127);
nand U10421 (N_10421,N_7728,N_6929);
and U10422 (N_10422,N_6045,N_7052);
or U10423 (N_10423,N_7098,N_9708);
xor U10424 (N_10424,N_9179,N_8700);
nor U10425 (N_10425,N_9328,N_5738);
nor U10426 (N_10426,N_6090,N_7276);
nand U10427 (N_10427,N_5555,N_7820);
nor U10428 (N_10428,N_9512,N_9386);
nor U10429 (N_10429,N_6427,N_6724);
nor U10430 (N_10430,N_9487,N_9985);
and U10431 (N_10431,N_5491,N_6076);
nand U10432 (N_10432,N_5282,N_6232);
xor U10433 (N_10433,N_6628,N_5578);
nor U10434 (N_10434,N_9384,N_5568);
xor U10435 (N_10435,N_5317,N_5916);
nor U10436 (N_10436,N_9828,N_9939);
xnor U10437 (N_10437,N_7267,N_5106);
or U10438 (N_10438,N_8994,N_5115);
and U10439 (N_10439,N_8814,N_6281);
and U10440 (N_10440,N_7625,N_5809);
nor U10441 (N_10441,N_5657,N_9820);
nor U10442 (N_10442,N_9867,N_9475);
and U10443 (N_10443,N_7725,N_7238);
and U10444 (N_10444,N_8869,N_9282);
or U10445 (N_10445,N_9890,N_6365);
nand U10446 (N_10446,N_5605,N_8771);
nor U10447 (N_10447,N_8252,N_8679);
nor U10448 (N_10448,N_5904,N_6643);
nor U10449 (N_10449,N_8105,N_7289);
or U10450 (N_10450,N_8301,N_5348);
nor U10451 (N_10451,N_9770,N_8640);
nor U10452 (N_10452,N_8215,N_9750);
nand U10453 (N_10453,N_7920,N_9198);
and U10454 (N_10454,N_9526,N_5460);
or U10455 (N_10455,N_6099,N_9509);
nor U10456 (N_10456,N_9559,N_6737);
nor U10457 (N_10457,N_7442,N_6624);
nand U10458 (N_10458,N_5036,N_8490);
and U10459 (N_10459,N_8272,N_7337);
and U10460 (N_10460,N_9722,N_9940);
and U10461 (N_10461,N_6119,N_9280);
nand U10462 (N_10462,N_5780,N_6595);
nand U10463 (N_10463,N_8744,N_6425);
nand U10464 (N_10464,N_8084,N_7068);
and U10465 (N_10465,N_8010,N_5770);
nand U10466 (N_10466,N_5247,N_8513);
or U10467 (N_10467,N_7466,N_5299);
nand U10468 (N_10468,N_8022,N_9401);
nand U10469 (N_10469,N_7230,N_7632);
and U10470 (N_10470,N_8804,N_5225);
nand U10471 (N_10471,N_7484,N_8294);
xor U10472 (N_10472,N_5600,N_8805);
xor U10473 (N_10473,N_8678,N_9930);
nor U10474 (N_10474,N_6666,N_9817);
and U10475 (N_10475,N_7749,N_8168);
nand U10476 (N_10476,N_9295,N_6513);
nor U10477 (N_10477,N_6939,N_9069);
nand U10478 (N_10478,N_7452,N_5908);
and U10479 (N_10479,N_7110,N_8393);
or U10480 (N_10480,N_5331,N_6711);
and U10481 (N_10481,N_8283,N_6850);
xnor U10482 (N_10482,N_8846,N_9306);
nor U10483 (N_10483,N_8504,N_6400);
xor U10484 (N_10484,N_7520,N_9625);
nand U10485 (N_10485,N_6295,N_7713);
nand U10486 (N_10486,N_9692,N_6354);
nand U10487 (N_10487,N_9176,N_5621);
and U10488 (N_10488,N_5629,N_6544);
xor U10489 (N_10489,N_7294,N_5107);
nand U10490 (N_10490,N_5327,N_7149);
nand U10491 (N_10491,N_8581,N_8977);
nor U10492 (N_10492,N_5470,N_5235);
or U10493 (N_10493,N_7762,N_5954);
nand U10494 (N_10494,N_9331,N_8575);
xor U10495 (N_10495,N_7857,N_6852);
or U10496 (N_10496,N_6360,N_5691);
nor U10497 (N_10497,N_7959,N_9795);
nor U10498 (N_10498,N_7639,N_6790);
xnor U10499 (N_10499,N_5143,N_9997);
or U10500 (N_10500,N_6821,N_9090);
or U10501 (N_10501,N_9588,N_7342);
nand U10502 (N_10502,N_7648,N_7652);
and U10503 (N_10503,N_7156,N_7313);
nand U10504 (N_10504,N_7446,N_7039);
or U10505 (N_10505,N_7386,N_9207);
and U10506 (N_10506,N_5559,N_8704);
nor U10507 (N_10507,N_7778,N_8360);
nand U10508 (N_10508,N_6491,N_5353);
or U10509 (N_10509,N_5441,N_8642);
nand U10510 (N_10510,N_7973,N_7721);
nand U10511 (N_10511,N_8503,N_8255);
or U10512 (N_10512,N_9922,N_7099);
or U10513 (N_10513,N_5607,N_8756);
nor U10514 (N_10514,N_5756,N_7896);
and U10515 (N_10515,N_5523,N_5851);
or U10516 (N_10516,N_9429,N_9834);
nand U10517 (N_10517,N_7494,N_9924);
nand U10518 (N_10518,N_9695,N_5945);
and U10519 (N_10519,N_5822,N_5324);
and U10520 (N_10520,N_6818,N_9092);
xor U10521 (N_10521,N_5995,N_8714);
xor U10522 (N_10522,N_7600,N_6878);
nor U10523 (N_10523,N_8825,N_5462);
xnor U10524 (N_10524,N_5914,N_9806);
nor U10525 (N_10525,N_6402,N_6518);
xor U10526 (N_10526,N_5430,N_8795);
or U10527 (N_10527,N_8211,N_8943);
nand U10528 (N_10528,N_6147,N_7988);
nand U10529 (N_10529,N_9360,N_5645);
nand U10530 (N_10530,N_9618,N_7836);
nor U10531 (N_10531,N_7305,N_7406);
nor U10532 (N_10532,N_6749,N_7143);
and U10533 (N_10533,N_7636,N_8627);
or U10534 (N_10534,N_8236,N_6692);
and U10535 (N_10535,N_7862,N_9966);
nor U10536 (N_10536,N_6036,N_6936);
xnor U10537 (N_10537,N_6087,N_5506);
nand U10538 (N_10538,N_5761,N_5426);
or U10539 (N_10539,N_6842,N_5526);
nor U10540 (N_10540,N_6834,N_8817);
nor U10541 (N_10541,N_6067,N_7371);
or U10542 (N_10542,N_5887,N_7082);
nor U10543 (N_10543,N_7883,N_8911);
or U10544 (N_10544,N_6029,N_6757);
or U10545 (N_10545,N_5911,N_9826);
nand U10546 (N_10546,N_6994,N_6648);
or U10547 (N_10547,N_5685,N_8312);
xnor U10548 (N_10548,N_9585,N_5831);
nand U10549 (N_10549,N_8388,N_6272);
nand U10550 (N_10550,N_6074,N_6296);
xnor U10551 (N_10551,N_6874,N_8878);
nor U10552 (N_10552,N_5948,N_9617);
nor U10553 (N_10553,N_7703,N_8163);
and U10554 (N_10554,N_9876,N_9312);
nor U10555 (N_10555,N_7779,N_9741);
and U10556 (N_10556,N_6370,N_5604);
xor U10557 (N_10557,N_6951,N_9013);
nand U10558 (N_10558,N_8330,N_8284);
nor U10559 (N_10559,N_5525,N_6918);
xor U10560 (N_10560,N_5189,N_8335);
nand U10561 (N_10561,N_6669,N_9182);
and U10562 (N_10562,N_9057,N_7982);
and U10563 (N_10563,N_6769,N_7433);
nor U10564 (N_10564,N_5397,N_5035);
nor U10565 (N_10565,N_8671,N_9761);
and U10566 (N_10566,N_8290,N_6007);
nor U10567 (N_10567,N_5679,N_7279);
and U10568 (N_10568,N_7816,N_9661);
or U10569 (N_10569,N_8387,N_6512);
or U10570 (N_10570,N_8491,N_8291);
nand U10571 (N_10571,N_5285,N_9003);
nor U10572 (N_10572,N_8728,N_5618);
or U10573 (N_10573,N_7577,N_8229);
or U10574 (N_10574,N_8950,N_9752);
or U10575 (N_10575,N_9454,N_6047);
or U10576 (N_10576,N_9934,N_6859);
and U10577 (N_10577,N_8636,N_7992);
and U10578 (N_10578,N_9322,N_5049);
and U10579 (N_10579,N_7731,N_9613);
nor U10580 (N_10580,N_7302,N_9253);
or U10581 (N_10581,N_9897,N_9759);
or U10582 (N_10582,N_9287,N_6304);
and U10583 (N_10583,N_8046,N_9728);
nand U10584 (N_10584,N_7269,N_7266);
nor U10585 (N_10585,N_7477,N_8669);
xnor U10586 (N_10586,N_9045,N_5968);
xnor U10587 (N_10587,N_9168,N_5016);
nand U10588 (N_10588,N_8725,N_8085);
and U10589 (N_10589,N_5204,N_5542);
nor U10590 (N_10590,N_9690,N_7163);
xnor U10591 (N_10591,N_6426,N_6747);
nand U10592 (N_10592,N_8777,N_5326);
or U10593 (N_10593,N_8153,N_7184);
nand U10594 (N_10594,N_8258,N_6672);
and U10595 (N_10595,N_8867,N_9407);
and U10596 (N_10596,N_8508,N_6213);
nand U10597 (N_10597,N_6125,N_6136);
nor U10598 (N_10598,N_9313,N_6139);
xnor U10599 (N_10599,N_9461,N_5417);
and U10600 (N_10600,N_6755,N_7175);
and U10601 (N_10601,N_6368,N_8589);
nand U10602 (N_10602,N_9514,N_6133);
nor U10603 (N_10603,N_8076,N_9737);
and U10604 (N_10604,N_5672,N_9584);
nor U10605 (N_10605,N_6828,N_7326);
nand U10606 (N_10606,N_6965,N_9640);
nor U10607 (N_10607,N_8749,N_8398);
and U10608 (N_10608,N_5684,N_8437);
nand U10609 (N_10609,N_5443,N_6961);
or U10610 (N_10610,N_6503,N_8907);
nand U10611 (N_10611,N_5739,N_8354);
xnor U10612 (N_10612,N_6599,N_5743);
or U10613 (N_10613,N_9275,N_5906);
xor U10614 (N_10614,N_8113,N_5160);
nor U10615 (N_10615,N_9630,N_9096);
and U10616 (N_10616,N_5784,N_7838);
or U10617 (N_10617,N_5432,N_9250);
nor U10618 (N_10618,N_9055,N_6644);
or U10619 (N_10619,N_6380,N_8806);
nand U10620 (N_10620,N_9747,N_9553);
xnor U10621 (N_10621,N_7872,N_9291);
nor U10622 (N_10622,N_8655,N_5583);
nor U10623 (N_10623,N_7187,N_6189);
nor U10624 (N_10624,N_6336,N_7684);
and U10625 (N_10625,N_5116,N_7554);
or U10626 (N_10626,N_6780,N_8095);
nor U10627 (N_10627,N_9024,N_6389);
nor U10628 (N_10628,N_7581,N_7840);
or U10629 (N_10629,N_9239,N_7627);
and U10630 (N_10630,N_5361,N_9814);
and U10631 (N_10631,N_6011,N_9856);
and U10632 (N_10632,N_7954,N_6130);
nor U10633 (N_10633,N_9333,N_5992);
or U10634 (N_10634,N_6362,N_9655);
and U10635 (N_10635,N_8077,N_9264);
nand U10636 (N_10636,N_9923,N_5099);
or U10637 (N_10637,N_9535,N_6478);
nor U10638 (N_10638,N_9975,N_8766);
nand U10639 (N_10639,N_6481,N_7960);
nand U10640 (N_10640,N_6075,N_6395);
or U10641 (N_10641,N_9501,N_5786);
or U10642 (N_10642,N_7575,N_6390);
and U10643 (N_10643,N_8736,N_8238);
and U10644 (N_10644,N_5888,N_8760);
nand U10645 (N_10645,N_7766,N_7399);
nand U10646 (N_10646,N_8324,N_5005);
or U10647 (N_10647,N_8106,N_7911);
or U10648 (N_10648,N_6563,N_8823);
nor U10649 (N_10649,N_6124,N_7010);
nor U10650 (N_10650,N_5765,N_6408);
nor U10651 (N_10651,N_5703,N_6632);
or U10652 (N_10652,N_5687,N_5617);
nor U10653 (N_10653,N_6363,N_7075);
xnor U10654 (N_10654,N_6943,N_5269);
and U10655 (N_10655,N_7897,N_5674);
and U10656 (N_10656,N_7800,N_5855);
or U10657 (N_10657,N_9387,N_8665);
nor U10658 (N_10658,N_5171,N_6188);
xor U10659 (N_10659,N_9356,N_5690);
or U10660 (N_10660,N_8614,N_7537);
or U10661 (N_10661,N_7031,N_6439);
or U10662 (N_10662,N_7998,N_6095);
or U10663 (N_10663,N_5689,N_8898);
or U10664 (N_10664,N_5693,N_8557);
nand U10665 (N_10665,N_5265,N_9102);
nand U10666 (N_10666,N_8793,N_6367);
or U10667 (N_10667,N_6638,N_8755);
xnor U10668 (N_10668,N_9595,N_5815);
or U10669 (N_10669,N_8835,N_8279);
or U10670 (N_10670,N_7125,N_7545);
and U10671 (N_10671,N_8916,N_5928);
and U10672 (N_10672,N_5812,N_5885);
nand U10673 (N_10673,N_6789,N_8036);
and U10674 (N_10674,N_8521,N_5157);
and U10675 (N_10675,N_5219,N_8322);
nand U10676 (N_10676,N_5183,N_8497);
nand U10677 (N_10677,N_6344,N_8662);
and U10678 (N_10678,N_7441,N_7890);
nor U10679 (N_10679,N_7415,N_7402);
or U10680 (N_10680,N_5952,N_5581);
and U10681 (N_10681,N_8942,N_9936);
nor U10682 (N_10682,N_7701,N_7153);
nor U10683 (N_10683,N_5279,N_5170);
nand U10684 (N_10684,N_6066,N_9363);
and U10685 (N_10685,N_8485,N_8081);
or U10686 (N_10686,N_9097,N_5175);
or U10687 (N_10687,N_9542,N_7162);
nor U10688 (N_10688,N_9845,N_7258);
nand U10689 (N_10689,N_5556,N_5943);
xor U10690 (N_10690,N_9979,N_8657);
or U10691 (N_10691,N_9951,N_7597);
nor U10692 (N_10692,N_5821,N_9972);
or U10693 (N_10693,N_6169,N_7232);
nand U10694 (N_10694,N_6432,N_5946);
and U10695 (N_10695,N_9430,N_8340);
and U10696 (N_10696,N_7593,N_9882);
or U10697 (N_10697,N_5781,N_9650);
nor U10698 (N_10698,N_6371,N_8947);
and U10699 (N_10699,N_5830,N_9919);
nor U10700 (N_10700,N_7380,N_7601);
or U10701 (N_10701,N_5500,N_8222);
nand U10702 (N_10702,N_5431,N_6849);
xor U10703 (N_10703,N_9394,N_7682);
or U10704 (N_10704,N_8198,N_9343);
nand U10705 (N_10705,N_9702,N_6671);
and U10706 (N_10706,N_5626,N_5133);
nand U10707 (N_10707,N_7366,N_7527);
xor U10708 (N_10708,N_8827,N_8759);
nor U10709 (N_10709,N_8419,N_5989);
nor U10710 (N_10710,N_7204,N_8092);
and U10711 (N_10711,N_9414,N_5064);
and U10712 (N_10712,N_6879,N_6140);
nand U10713 (N_10713,N_9308,N_6598);
or U10714 (N_10714,N_5419,N_7062);
nor U10715 (N_10715,N_7614,N_5901);
or U10716 (N_10716,N_7704,N_7487);
or U10717 (N_10717,N_5708,N_5263);
or U10718 (N_10718,N_6974,N_9541);
or U10719 (N_10719,N_6885,N_6097);
nand U10720 (N_10720,N_7330,N_8969);
nor U10721 (N_10721,N_9298,N_6494);
and U10722 (N_10722,N_8048,N_7041);
or U10723 (N_10723,N_5680,N_8949);
nand U10724 (N_10724,N_7024,N_6461);
xor U10725 (N_10725,N_6144,N_5434);
nor U10726 (N_10726,N_9523,N_6931);
nand U10727 (N_10727,N_7051,N_6429);
and U10728 (N_10728,N_7683,N_5563);
nand U10729 (N_10729,N_8242,N_9310);
nand U10730 (N_10730,N_7710,N_6743);
nor U10731 (N_10731,N_6800,N_6835);
nand U10732 (N_10732,N_7312,N_6155);
xor U10733 (N_10733,N_8887,N_5057);
and U10734 (N_10734,N_8260,N_7070);
and U10735 (N_10735,N_7284,N_5467);
or U10736 (N_10736,N_8194,N_8167);
xor U10737 (N_10737,N_6658,N_6730);
nor U10738 (N_10738,N_9175,N_5487);
xnor U10739 (N_10739,N_5303,N_7909);
and U10740 (N_10740,N_9875,N_7332);
and U10741 (N_10741,N_8460,N_6265);
or U10742 (N_10742,N_6172,N_9718);
or U10743 (N_10743,N_6107,N_5502);
nand U10744 (N_10744,N_8126,N_5671);
or U10745 (N_10745,N_9083,N_5535);
or U10746 (N_10746,N_8181,N_7224);
and U10747 (N_10747,N_8658,N_8128);
nor U10748 (N_10748,N_8003,N_7829);
nor U10749 (N_10749,N_7103,N_6736);
nor U10750 (N_10750,N_7333,N_6816);
or U10751 (N_10751,N_6250,N_5849);
nand U10752 (N_10752,N_6516,N_9942);
and U10753 (N_10753,N_5406,N_5492);
or U10754 (N_10754,N_5154,N_7558);
nand U10755 (N_10755,N_7121,N_9125);
and U10756 (N_10756,N_8988,N_8373);
and U10757 (N_10757,N_6892,N_9892);
nor U10758 (N_10758,N_7881,N_7864);
and U10759 (N_10759,N_5895,N_9816);
or U10760 (N_10760,N_5722,N_7336);
and U10761 (N_10761,N_5903,N_9007);
and U10762 (N_10762,N_7460,N_6700);
nand U10763 (N_10763,N_7286,N_5881);
or U10764 (N_10764,N_6412,N_7549);
and U10765 (N_10765,N_8654,N_7927);
and U10766 (N_10766,N_7349,N_9126);
or U10767 (N_10767,N_5079,N_7325);
nor U10768 (N_10768,N_8422,N_8139);
and U10769 (N_10769,N_9124,N_8009);
nand U10770 (N_10770,N_9232,N_6996);
nor U10771 (N_10771,N_7464,N_5740);
nor U10772 (N_10772,N_6428,N_5090);
xor U10773 (N_10773,N_7392,N_9590);
nor U10774 (N_10774,N_8894,N_7410);
nor U10775 (N_10775,N_6703,N_9713);
or U10776 (N_10776,N_9917,N_7767);
or U10777 (N_10777,N_8746,N_6655);
nand U10778 (N_10778,N_7686,N_9086);
nand U10779 (N_10779,N_9495,N_6781);
nand U10780 (N_10780,N_9054,N_9963);
nand U10781 (N_10781,N_8652,N_9392);
and U10782 (N_10782,N_6244,N_5403);
xor U10783 (N_10783,N_7970,N_5866);
and U10784 (N_10784,N_9355,N_6112);
nand U10785 (N_10785,N_5847,N_8741);
xnor U10786 (N_10786,N_5814,N_7822);
and U10787 (N_10787,N_5704,N_9779);
and U10788 (N_10788,N_8605,N_8549);
nor U10789 (N_10789,N_9148,N_8035);
or U10790 (N_10790,N_5497,N_6539);
and U10791 (N_10791,N_5421,N_5060);
nor U10792 (N_10792,N_8917,N_8565);
xor U10793 (N_10793,N_8414,N_9085);
or U10794 (N_10794,N_8807,N_5997);
nor U10795 (N_10795,N_7420,N_7118);
or U10796 (N_10796,N_9945,N_8454);
nand U10797 (N_10797,N_7879,N_7171);
nand U10798 (N_10798,N_9573,N_7587);
or U10799 (N_10799,N_9929,N_5640);
or U10800 (N_10800,N_8995,N_5454);
nand U10801 (N_10801,N_9627,N_9067);
nand U10802 (N_10802,N_8909,N_7458);
nor U10803 (N_10803,N_7942,N_9714);
and U10804 (N_10804,N_8021,N_8978);
and U10805 (N_10805,N_5261,N_6832);
and U10806 (N_10806,N_9516,N_5270);
nand U10807 (N_10807,N_7532,N_9815);
and U10808 (N_10808,N_6198,N_5638);
xnor U10809 (N_10809,N_6338,N_7277);
xnor U10810 (N_10810,N_9036,N_7054);
or U10811 (N_10811,N_9874,N_6896);
and U10812 (N_10812,N_5571,N_9432);
nor U10813 (N_10813,N_6665,N_5024);
nor U10814 (N_10814,N_8042,N_7985);
nor U10815 (N_10815,N_7397,N_7961);
nand U10816 (N_10816,N_5436,N_6622);
nand U10817 (N_10817,N_9311,N_5347);
nor U10818 (N_10818,N_9744,N_7253);
xor U10819 (N_10819,N_5357,N_7502);
nand U10820 (N_10820,N_8205,N_7594);
and U10821 (N_10821,N_7271,N_9236);
nand U10822 (N_10822,N_8475,N_9976);
and U10823 (N_10823,N_5455,N_9062);
nor U10824 (N_10824,N_5550,N_5977);
or U10825 (N_10825,N_8550,N_7474);
nand U10826 (N_10826,N_7531,N_6771);
nand U10827 (N_10827,N_8470,N_5734);
nand U10828 (N_10828,N_7972,N_7469);
nand U10829 (N_10829,N_8435,N_6562);
nand U10830 (N_10830,N_8858,N_9161);
or U10831 (N_10831,N_8758,N_5485);
and U10832 (N_10832,N_6870,N_7454);
or U10833 (N_10833,N_8345,N_8517);
nand U10834 (N_10834,N_6237,N_9381);
or U10835 (N_10835,N_5252,N_9911);
or U10836 (N_10836,N_9423,N_9234);
and U10837 (N_10837,N_9536,N_7891);
and U10838 (N_10838,N_6488,N_8329);
nor U10839 (N_10839,N_8685,N_9859);
nor U10840 (N_10840,N_9241,N_5328);
nor U10841 (N_10841,N_7559,N_6869);
and U10842 (N_10842,N_5483,N_8347);
and U10843 (N_10843,N_5246,N_9178);
nand U10844 (N_10844,N_9259,N_7368);
nor U10845 (N_10845,N_6204,N_7695);
nand U10846 (N_10846,N_9578,N_7109);
nand U10847 (N_10847,N_6282,N_6667);
nand U10848 (N_10848,N_6694,N_8429);
xor U10849 (N_10849,N_5963,N_7835);
and U10850 (N_10850,N_7708,N_5209);
or U10851 (N_10851,N_6844,N_5062);
or U10852 (N_10852,N_6134,N_6606);
xnor U10853 (N_10853,N_9158,N_9604);
and U10854 (N_10854,N_6280,N_9799);
and U10855 (N_10855,N_5254,N_6104);
or U10856 (N_10856,N_6661,N_9730);
and U10857 (N_10857,N_5826,N_7147);
nor U10858 (N_10858,N_6242,N_9140);
or U10859 (N_10859,N_9950,N_7438);
or U10860 (N_10860,N_9790,N_5666);
or U10861 (N_10861,N_7595,N_5272);
or U10862 (N_10862,N_8531,N_5350);
or U10863 (N_10863,N_6693,N_8484);
and U10864 (N_10864,N_6572,N_7280);
nand U10865 (N_10865,N_5880,N_7357);
nand U10866 (N_10866,N_5858,N_8044);
or U10867 (N_10867,N_8768,N_6224);
nand U10868 (N_10868,N_9513,N_8512);
nor U10869 (N_10869,N_5315,N_5969);
nor U10870 (N_10870,N_8323,N_5066);
nor U10871 (N_10871,N_9841,N_5469);
xnor U10872 (N_10872,N_9996,N_7066);
and U10873 (N_10873,N_9937,N_6895);
nor U10874 (N_10874,N_5852,N_5800);
nor U10875 (N_10875,N_7200,N_7219);
and U10876 (N_10876,N_6531,N_8561);
and U10877 (N_10877,N_7760,N_5833);
nand U10878 (N_10878,N_9499,N_8598);
and U10879 (N_10879,N_7198,N_7934);
nor U10880 (N_10880,N_5973,N_7757);
nor U10881 (N_10881,N_7939,N_9652);
or U10882 (N_10882,N_9305,N_6739);
and U10883 (N_10883,N_9349,N_7461);
xor U10884 (N_10884,N_6676,N_5222);
nor U10885 (N_10885,N_9375,N_5073);
nand U10886 (N_10886,N_8120,N_8089);
nor U10887 (N_10887,N_7854,N_5055);
or U10888 (N_10888,N_5924,N_8432);
or U10889 (N_10889,N_6316,N_7668);
or U10890 (N_10890,N_5420,N_5498);
nand U10891 (N_10891,N_6485,N_6238);
and U10892 (N_10892,N_9350,N_5255);
and U10893 (N_10893,N_9864,N_7931);
nand U10894 (N_10894,N_7352,N_9489);
or U10895 (N_10895,N_8892,N_8585);
nor U10896 (N_10896,N_8865,N_6476);
and U10897 (N_10897,N_7780,N_9113);
and U10898 (N_10898,N_6267,N_9780);
nor U10899 (N_10899,N_5495,N_6836);
and U10900 (N_10900,N_5439,N_9177);
and U10901 (N_10901,N_7930,N_5330);
nand U10902 (N_10902,N_5742,N_9973);
nor U10903 (N_10903,N_5721,N_9600);
nand U10904 (N_10904,N_8688,N_6116);
nor U10905 (N_10905,N_7120,N_8778);
and U10906 (N_10906,N_5442,N_5301);
xnor U10907 (N_10907,N_8162,N_7574);
and U10908 (N_10908,N_9956,N_5410);
nand U10909 (N_10909,N_8997,N_9031);
or U10910 (N_10910,N_7861,N_5496);
or U10911 (N_10911,N_6543,N_8160);
nor U10912 (N_10912,N_7069,N_8137);
and U10913 (N_10913,N_7678,N_7538);
nor U10914 (N_10914,N_8087,N_7493);
or U10915 (N_10915,N_7884,N_9606);
nand U10916 (N_10916,N_5705,N_5816);
and U10917 (N_10917,N_7885,N_8509);
or U10918 (N_10918,N_7306,N_6387);
and U10919 (N_10919,N_7007,N_7362);
and U10920 (N_10920,N_7814,N_7378);
nand U10921 (N_10921,N_7815,N_9257);
nor U10922 (N_10922,N_7685,N_9159);
or U10923 (N_10923,N_7900,N_9525);
or U10924 (N_10924,N_6605,N_5582);
nand U10925 (N_10925,N_6586,N_9591);
nor U10926 (N_10926,N_5287,N_8378);
and U10927 (N_10927,N_7944,N_8570);
nor U10928 (N_10928,N_5015,N_7071);
or U10929 (N_10929,N_6472,N_5351);
and U10930 (N_10930,N_9693,N_8328);
xnor U10931 (N_10931,N_5875,N_5603);
nor U10932 (N_10932,N_7917,N_8233);
xor U10933 (N_10933,N_8525,N_7689);
nand U10934 (N_10934,N_6152,N_5633);
xor U10935 (N_10935,N_9967,N_9470);
nand U10936 (N_10936,N_6825,N_6659);
and U10937 (N_10937,N_6609,N_8715);
nand U10938 (N_10938,N_8075,N_7553);
nor U10939 (N_10939,N_5046,N_8843);
nor U10940 (N_10940,N_9665,N_7888);
nand U10941 (N_10941,N_7654,N_6123);
nor U10942 (N_10942,N_5987,N_9026);
or U10943 (N_10943,N_9359,N_9715);
nor U10944 (N_10944,N_5994,N_6063);
or U10945 (N_10945,N_5889,N_5346);
or U10946 (N_10946,N_8944,N_7268);
and U10947 (N_10947,N_9657,N_8897);
nand U10948 (N_10948,N_7733,N_5988);
nand U10949 (N_10949,N_5653,N_6616);
nor U10950 (N_10950,N_6325,N_5148);
and U10951 (N_10951,N_5787,N_9441);
and U10952 (N_10952,N_9039,N_8775);
xor U10953 (N_10953,N_5198,N_7951);
or U10954 (N_10954,N_5932,N_7643);
and U10955 (N_10955,N_8038,N_5651);
nand U10956 (N_10956,N_6696,N_5163);
or U10957 (N_10957,N_8444,N_9033);
nand U10958 (N_10958,N_8334,N_5793);
nand U10959 (N_10959,N_8697,N_9528);
nor U10960 (N_10960,N_5823,N_6914);
nand U10961 (N_10961,N_6173,N_5239);
or U10962 (N_10962,N_9335,N_9505);
xnor U10963 (N_10963,N_7022,N_5513);
nor U10964 (N_10964,N_5829,N_5929);
or U10965 (N_10965,N_7486,N_5167);
xnor U10966 (N_10966,N_7256,N_7067);
or U10967 (N_10967,N_6653,N_7702);
nor U10968 (N_10968,N_8982,N_7843);
nor U10969 (N_10969,N_6311,N_5913);
or U10970 (N_10970,N_6319,N_9786);
or U10971 (N_10971,N_8538,N_5192);
nand U10972 (N_10972,N_7565,N_7519);
or U10973 (N_10973,N_5912,N_9836);
xnor U10974 (N_10974,N_9532,N_8607);
and U10975 (N_10975,N_7283,N_6487);
and U10976 (N_10976,N_8965,N_5481);
or U10977 (N_10977,N_7043,N_8461);
and U10978 (N_10978,N_8542,N_6333);
and U10979 (N_10979,N_9104,N_6777);
nor U10980 (N_10980,N_9283,N_5056);
or U10981 (N_10981,N_5113,N_6973);
or U10982 (N_10982,N_9689,N_7159);
xnor U10983 (N_10983,N_7199,N_9504);
and U10984 (N_10984,N_5412,N_6838);
xor U10985 (N_10985,N_6806,N_8174);
nor U10986 (N_10986,N_6962,N_8779);
and U10987 (N_10987,N_8007,N_5030);
nand U10988 (N_10988,N_7379,N_8116);
nand U10989 (N_10989,N_9209,N_6276);
and U10990 (N_10990,N_8619,N_8663);
nand U10991 (N_10991,N_9206,N_5516);
nor U10992 (N_10992,N_6471,N_5281);
and U10993 (N_10993,N_5202,N_7805);
nand U10994 (N_10994,N_6811,N_8954);
xnor U10995 (N_10995,N_5774,N_6031);
and U10996 (N_10996,N_8976,N_7919);
or U10997 (N_10997,N_9830,N_5744);
and U10998 (N_10998,N_9626,N_8695);
or U10999 (N_10999,N_8612,N_9108);
or U11000 (N_11000,N_9223,N_5314);
or U11001 (N_11001,N_6883,N_9671);
xor U11002 (N_11002,N_5688,N_9266);
nand U11003 (N_11003,N_5919,N_6604);
and U11004 (N_11004,N_6517,N_6793);
nand U11005 (N_11005,N_7046,N_8930);
or U11006 (N_11006,N_7365,N_6657);
and U11007 (N_11007,N_5659,N_8127);
nor U11008 (N_11008,N_6449,N_7936);
xnor U11009 (N_11009,N_7226,N_7090);
nor U11010 (N_11010,N_6783,N_7036);
or U11011 (N_11011,N_6201,N_8078);
or U11012 (N_11012,N_5042,N_8650);
nand U11013 (N_11013,N_7550,N_7430);
nand U11014 (N_11014,N_8244,N_7739);
and U11015 (N_11015,N_7826,N_6774);
nand U11016 (N_11016,N_7511,N_6910);
nor U11017 (N_11017,N_7991,N_9970);
nand U11018 (N_11018,N_7307,N_6592);
nand U11019 (N_11019,N_8729,N_6721);
nand U11020 (N_11020,N_6583,N_8478);
nand U11021 (N_11021,N_6715,N_7186);
and U11022 (N_11022,N_5976,N_8574);
xor U11023 (N_11023,N_5579,N_9572);
nand U11024 (N_11024,N_7726,N_6017);
nand U11025 (N_11025,N_8500,N_9163);
nor U11026 (N_11026,N_5092,N_5227);
nor U11027 (N_11027,N_9417,N_6680);
nor U11028 (N_11028,N_5861,N_5053);
or U11029 (N_11029,N_5293,N_9451);
or U11030 (N_11030,N_7803,N_8935);
nand U11031 (N_11031,N_5422,N_6262);
nor U11032 (N_11032,N_6857,N_7021);
nor U11033 (N_11033,N_6575,N_9155);
and U11034 (N_11034,N_5356,N_9051);
or U11035 (N_11035,N_6121,N_6071);
nand U11036 (N_11036,N_8559,N_9615);
xnor U11037 (N_11037,N_8356,N_9696);
nor U11038 (N_11038,N_6647,N_7655);
or U11039 (N_11039,N_8262,N_6863);
and U11040 (N_11040,N_9059,N_7657);
and U11041 (N_11041,N_8451,N_5716);
nand U11042 (N_11042,N_8249,N_5962);
nor U11043 (N_11043,N_8670,N_7913);
nor U11044 (N_11044,N_5295,N_6394);
or U11045 (N_11045,N_9160,N_8278);
nand U11046 (N_11046,N_7679,N_7647);
nor U11047 (N_11047,N_5190,N_8268);
nor U11048 (N_11048,N_7672,N_9154);
or U11049 (N_11049,N_9348,N_8302);
nand U11050 (N_11050,N_8548,N_9317);
or U11051 (N_11051,N_7177,N_6167);
or U11052 (N_11052,N_8351,N_5763);
and U11053 (N_11053,N_6536,N_5416);
xnor U11054 (N_11054,N_8093,N_7564);
nand U11055 (N_11055,N_9469,N_5440);
or U11056 (N_11056,N_6523,N_6567);
nor U11057 (N_11057,N_7669,N_9571);
nand U11058 (N_11058,N_7037,N_9607);
and U11059 (N_11059,N_6813,N_6709);
xnor U11060 (N_11060,N_5546,N_9138);
or U11061 (N_11061,N_6174,N_9258);
and U11062 (N_11062,N_7367,N_5292);
nor U11063 (N_11063,N_7154,N_7358);
and U11064 (N_11064,N_8344,N_7419);
xnor U11065 (N_11065,N_6385,N_8708);
and U11066 (N_11066,N_5768,N_7676);
or U11067 (N_11067,N_9200,N_9896);
or U11068 (N_11068,N_6180,N_9157);
or U11069 (N_11069,N_5714,N_9486);
nand U11070 (N_11070,N_7690,N_5567);
and U11071 (N_11071,N_8102,N_6573);
and U11072 (N_11072,N_5930,N_8686);
nand U11073 (N_11073,N_8336,N_5257);
nand U11074 (N_11074,N_8932,N_9144);
and U11075 (N_11075,N_5720,N_9151);
or U11076 (N_11076,N_5405,N_9073);
or U11077 (N_11077,N_9685,N_9545);
or U11078 (N_11078,N_9457,N_5773);
nor U11079 (N_11079,N_5637,N_7273);
or U11080 (N_11080,N_6183,N_9150);
nand U11081 (N_11081,N_7621,N_9270);
nand U11082 (N_11082,N_7242,N_7391);
or U11083 (N_11083,N_9745,N_9082);
nand U11084 (N_11084,N_6191,N_9368);
or U11085 (N_11085,N_7340,N_6264);
nand U11086 (N_11086,N_8855,N_5108);
nand U11087 (N_11087,N_9805,N_6034);
nor U11088 (N_11088,N_8989,N_7428);
and U11089 (N_11089,N_7456,N_5890);
nand U11090 (N_11090,N_6541,N_5082);
nand U11091 (N_11091,N_8296,N_8017);
nor U11092 (N_11092,N_9697,N_8495);
or U11093 (N_11093,N_7915,N_8192);
or U11094 (N_11094,N_6571,N_8953);
nor U11095 (N_11095,N_5297,N_6532);
nor U11096 (N_11096,N_7034,N_8056);
nand U11097 (N_11097,N_7451,N_8097);
nor U11098 (N_11098,N_6382,N_6915);
or U11099 (N_11099,N_8108,N_9840);
nor U11100 (N_11100,N_5043,N_6020);
nor U11101 (N_11101,N_5539,N_5185);
xnor U11102 (N_11102,N_9537,N_5517);
or U11103 (N_11103,N_5807,N_7839);
xor U11104 (N_11104,N_7999,N_9778);
nor U11105 (N_11105,N_7794,N_6438);
and U11106 (N_11106,N_7755,N_7645);
or U11107 (N_11107,N_6805,N_6663);
nor U11108 (N_11108,N_7591,N_8792);
or U11109 (N_11109,N_6982,N_8457);
nor U11110 (N_11110,N_6867,N_6960);
nand U11111 (N_11111,N_7955,N_8711);
nor U11112 (N_11112,N_5950,N_5466);
or U11113 (N_11113,N_6799,N_6275);
nor U11114 (N_11114,N_6877,N_7772);
or U11115 (N_11115,N_9404,N_7497);
xor U11116 (N_11116,N_7488,N_6802);
nor U11117 (N_11117,N_6796,N_6524);
or U11118 (N_11118,N_9872,N_9450);
nor U11119 (N_11119,N_7526,N_5862);
nand U11120 (N_11120,N_5902,N_8956);
and U11121 (N_11121,N_7522,N_8369);
and U11122 (N_11122,N_9656,N_5664);
nand U11123 (N_11123,N_8937,N_5834);
nand U11124 (N_11124,N_9261,N_8896);
nand U11125 (N_11125,N_7220,N_6268);
xnor U11126 (N_11126,N_9848,N_8752);
nor U11127 (N_11127,N_8803,N_7626);
nand U11128 (N_11128,N_5027,N_8155);
nand U11129 (N_11129,N_7201,N_8307);
nand U11130 (N_11130,N_7616,N_7122);
nor U11131 (N_11131,N_8140,N_7806);
or U11132 (N_11132,N_8135,N_9005);
nor U11133 (N_11133,N_9153,N_9344);
or U11134 (N_11134,N_5778,N_5859);
or U11135 (N_11135,N_7096,N_8463);
xor U11136 (N_11136,N_7080,N_7720);
nand U11137 (N_11137,N_5893,N_9798);
and U11138 (N_11138,N_5249,N_7002);
nand U11139 (N_11139,N_9593,N_5882);
nand U11140 (N_11140,N_9204,N_5766);
or U11141 (N_11141,N_7602,N_6837);
or U11142 (N_11142,N_5061,N_6972);
nor U11143 (N_11143,N_7260,N_9174);
nor U11144 (N_11144,N_6392,N_9409);
nor U11145 (N_11145,N_8243,N_8717);
and U11146 (N_11146,N_6415,N_6529);
nand U11147 (N_11147,N_6722,N_6417);
or U11148 (N_11148,N_9460,N_7030);
nor U11149 (N_11149,N_6591,N_7662);
nor U11150 (N_11150,N_9412,N_5712);
nor U11151 (N_11151,N_9229,N_6585);
and U11152 (N_11152,N_8371,N_8132);
or U11153 (N_11153,N_5574,N_9569);
and U11154 (N_11154,N_6128,N_9883);
or U11155 (N_11155,N_5586,N_8609);
or U11156 (N_11156,N_7763,N_5096);
and U11157 (N_11157,N_7369,N_6913);
nand U11158 (N_11158,N_9357,N_8273);
or U11159 (N_11159,N_6318,N_6113);
and U11160 (N_11160,N_5505,N_8524);
xor U11161 (N_11161,N_6713,N_8948);
or U11162 (N_11162,N_8280,N_7579);
or U11163 (N_11163,N_5414,N_5141);
nand U11164 (N_11164,N_7207,N_9129);
xor U11165 (N_11165,N_6864,N_8638);
and U11166 (N_11166,N_6719,N_6685);
nor U11167 (N_11167,N_8580,N_5214);
nor U11168 (N_11168,N_9304,N_7202);
and U11169 (N_11169,N_8456,N_7206);
xnor U11170 (N_11170,N_8819,N_6253);
or U11171 (N_11171,N_8201,N_6788);
or U11172 (N_11172,N_6004,N_5217);
and U11173 (N_11173,N_8514,N_7585);
and U11174 (N_11174,N_7376,N_8579);
nor U11175 (N_11175,N_9694,N_7697);
nor U11176 (N_11176,N_5728,N_9614);
nand U11177 (N_11177,N_9510,N_5508);
and U11178 (N_11178,N_7876,N_8060);
and U11179 (N_11179,N_5636,N_5210);
xnor U11180 (N_11180,N_9012,N_7117);
or U11181 (N_11181,N_7667,N_9916);
or U11182 (N_11182,N_7688,N_7751);
nor U11183 (N_11183,N_7310,N_7904);
and U11184 (N_11184,N_5843,N_5709);
nand U11185 (N_11185,N_5084,N_7285);
nand U11186 (N_11186,N_5717,N_8516);
nand U11187 (N_11187,N_8300,N_9920);
or U11188 (N_11188,N_5910,N_7027);
and U11189 (N_11189,N_9278,N_8418);
and U11190 (N_11190,N_6357,N_7304);
or U11191 (N_11191,N_9858,N_6728);
and U11192 (N_11192,N_7887,N_8633);
or U11193 (N_11193,N_8813,N_7827);
nor U11194 (N_11194,N_8129,N_6490);
nand U11195 (N_11195,N_7875,N_6241);
xor U11196 (N_11196,N_5536,N_8055);
xnor U11197 (N_11197,N_6690,N_9944);
or U11198 (N_11198,N_8150,N_9596);
nand U11199 (N_11199,N_5014,N_5841);
nor U11200 (N_11200,N_9443,N_8754);
and U11201 (N_11201,N_5769,N_6463);
and U11202 (N_11202,N_6170,N_5452);
and U11203 (N_11203,N_6521,N_5404);
or U11204 (N_11204,N_7194,N_5122);
nand U11205 (N_11205,N_7417,N_8620);
nand U11206 (N_11206,N_8476,N_9080);
nand U11207 (N_11207,N_8067,N_8138);
xor U11208 (N_11208,N_9156,N_7513);
nor U11209 (N_11209,N_7032,N_7364);
and U11210 (N_11210,N_6968,N_7631);
nor U11211 (N_11211,N_8286,N_8144);
and U11212 (N_11212,N_6246,N_6830);
and U11213 (N_11213,N_6093,N_5045);
nor U11214 (N_11214,N_8062,N_7033);
nor U11215 (N_11215,N_5832,N_8664);
nand U11216 (N_11216,N_6447,N_9852);
nor U11217 (N_11217,N_8573,N_5820);
nor U11218 (N_11218,N_6542,N_5736);
and U11219 (N_11219,N_6100,N_8868);
or U11220 (N_11220,N_8597,N_9262);
nand U11221 (N_11221,N_6738,N_7941);
nor U11222 (N_11222,N_9705,N_8791);
nor U11223 (N_11223,N_5312,N_8277);
xor U11224 (N_11224,N_8864,N_9133);
xnor U11225 (N_11225,N_9185,N_6618);
xor U11226 (N_11226,N_8926,N_5699);
nand U11227 (N_11227,N_9027,N_8383);
xor U11228 (N_11228,N_6988,N_9633);
nand U11229 (N_11229,N_8773,N_5119);
or U11230 (N_11230,N_5923,N_9777);
nor U11231 (N_11231,N_6785,N_8112);
and U11232 (N_11232,N_5248,N_9434);
nand U11233 (N_11233,N_9774,N_7086);
or U11234 (N_11234,N_8849,N_8488);
nand U11235 (N_11235,N_5597,N_6211);
nand U11236 (N_11236,N_7903,N_6436);
nand U11237 (N_11237,N_7393,N_7831);
and U11238 (N_11238,N_5808,N_8327);
and U11239 (N_11239,N_9143,N_9030);
nor U11240 (N_11240,N_8019,N_6640);
and U11241 (N_11241,N_7008,N_7056);
nand U11242 (N_11242,N_8407,N_5187);
or U11243 (N_11243,N_5354,N_9479);
xor U11244 (N_11244,N_7480,N_9691);
or U11245 (N_11245,N_8395,N_5126);
nand U11246 (N_11246,N_5611,N_5697);
xor U11247 (N_11247,N_6957,N_6919);
nor U11248 (N_11248,N_9084,N_7395);
xor U11249 (N_11249,N_8071,N_5339);
and U11250 (N_11250,N_5211,N_9203);
and U11251 (N_11251,N_7734,N_6083);
nand U11252 (N_11252,N_6310,N_8122);
or U11253 (N_11253,N_9684,N_6477);
or U11254 (N_11254,N_9522,N_7932);
xor U11255 (N_11255,N_5220,N_7790);
and U11256 (N_11256,N_7339,N_8961);
nor U11257 (N_11257,N_6149,N_7746);
nor U11258 (N_11258,N_5394,N_9732);
nor U11259 (N_11259,N_6118,N_6050);
nor U11260 (N_11260,N_9592,N_5683);
nor U11261 (N_11261,N_5086,N_8032);
or U11262 (N_11262,N_5182,N_9518);
nand U11263 (N_11263,N_6868,N_5146);
and U11264 (N_11264,N_7061,N_7275);
nor U11265 (N_11265,N_8338,N_8659);
xnor U11266 (N_11266,N_5615,N_9666);
and U11267 (N_11267,N_8733,N_7850);
or U11268 (N_11268,N_7221,N_5870);
nand U11269 (N_11269,N_8906,N_5686);
or U11270 (N_11270,N_8996,N_7530);
nor U11271 (N_11271,N_5276,N_8933);
nand U11272 (N_11272,N_6334,N_5727);
nand U11273 (N_11273,N_6239,N_6207);
xor U11274 (N_11274,N_6992,N_6617);
and U11275 (N_11275,N_9061,N_7618);
and U11276 (N_11276,N_9763,N_6373);
or U11277 (N_11277,N_7842,N_7938);
or U11278 (N_11278,N_9716,N_9134);
and U11279 (N_11279,N_5590,N_8528);
and U11280 (N_11280,N_8309,N_8922);
and U11281 (N_11281,N_8080,N_6462);
xnor U11282 (N_11282,N_8753,N_6258);
nor U11283 (N_11283,N_8187,N_8474);
or U11284 (N_11284,N_7435,N_5267);
nor U11285 (N_11285,N_7963,N_8905);
nor U11286 (N_11286,N_5180,N_9436);
and U11287 (N_11287,N_9813,N_8146);
nand U11288 (N_11288,N_8259,N_9629);
or U11289 (N_11289,N_5038,N_5236);
or U11290 (N_11290,N_8053,N_5153);
or U11291 (N_11291,N_6522,N_6637);
nor U11292 (N_11292,N_5490,N_8204);
or U11293 (N_11293,N_6898,N_8199);
nand U11294 (N_11294,N_7649,N_7015);
xnor U11295 (N_11295,N_6223,N_9803);
nand U11296 (N_11296,N_6215,N_9230);
nor U11297 (N_11297,N_5782,N_8645);
nor U11298 (N_11298,N_7290,N_8219);
and U11299 (N_11299,N_8452,N_8763);
xnor U11300 (N_11300,N_5003,N_7492);
and U11301 (N_11301,N_7747,N_9638);
nor U11302 (N_11302,N_8568,N_6060);
and U11303 (N_11303,N_9829,N_9928);
and U11304 (N_11304,N_6254,N_8991);
or U11305 (N_11305,N_6963,N_5644);
or U11306 (N_11306,N_7592,N_5134);
nor U11307 (N_11307,N_5547,N_7361);
or U11308 (N_11308,N_8065,N_9849);
nor U11309 (N_11309,N_5218,N_8735);
nor U11310 (N_11310,N_6452,N_5584);
and U11311 (N_11311,N_8635,N_6964);
nor U11312 (N_11312,N_7473,N_6210);
nand U11313 (N_11313,N_6634,N_9244);
nor U11314 (N_11314,N_9099,N_5169);
and U11315 (N_11315,N_6814,N_7562);
nand U11316 (N_11316,N_8992,N_5737);
nand U11317 (N_11317,N_6048,N_5488);
nor U11318 (N_11318,N_8202,N_7124);
nand U11319 (N_11319,N_9933,N_5795);
and U11320 (N_11320,N_8025,N_8596);
or U11321 (N_11321,N_8880,N_5905);
and U11322 (N_11322,N_6498,N_9734);
and U11323 (N_11323,N_9802,N_7088);
nor U11324 (N_11324,N_5892,N_7265);
or U11325 (N_11325,N_8772,N_9165);
and U11326 (N_11326,N_8938,N_7126);
or U11327 (N_11327,N_5242,N_8839);
or U11328 (N_11328,N_5724,N_9058);
or U11329 (N_11329,N_7514,N_6511);
or U11330 (N_11330,N_7389,N_5383);
and U11331 (N_11331,N_9017,N_8100);
nor U11332 (N_11332,N_9070,N_9644);
or U11333 (N_11333,N_9490,N_9788);
and U11334 (N_11334,N_6509,N_5336);
or U11335 (N_11335,N_5872,N_5196);
xnor U11336 (N_11336,N_9020,N_6765);
xor U11337 (N_11337,N_7784,N_9225);
nor U11338 (N_11338,N_5616,N_6168);
xor U11339 (N_11339,N_6506,N_6110);
or U11340 (N_11340,N_5271,N_5389);
or U11341 (N_11341,N_8902,N_8774);
xor U11342 (N_11342,N_7539,N_6068);
nor U11343 (N_11343,N_5545,N_5103);
nand U11344 (N_11344,N_7624,N_8210);
and U11345 (N_11345,N_5482,N_8857);
and U11346 (N_11346,N_5284,N_7536);
nor U11347 (N_11347,N_6073,N_6596);
nand U11348 (N_11348,N_5386,N_7190);
or U11349 (N_11349,N_5538,N_6303);
nor U11350 (N_11350,N_8410,N_5707);
or U11351 (N_11351,N_7426,N_6597);
and U11352 (N_11352,N_6923,N_5401);
nor U11353 (N_11353,N_7129,N_6103);
and U11354 (N_11354,N_7510,N_5732);
or U11355 (N_11355,N_6157,N_7495);
nand U11356 (N_11356,N_8304,N_5237);
nor U11357 (N_11357,N_5999,N_9581);
or U11358 (N_11358,N_9819,N_8428);
nor U11359 (N_11359,N_5402,N_5797);
and U11360 (N_11360,N_9491,N_5775);
nor U11361 (N_11361,N_7644,N_5321);
xor U11362 (N_11362,N_5075,N_6891);
nand U11363 (N_11363,N_6997,N_8537);
nor U11364 (N_11364,N_6980,N_7786);
nor U11365 (N_11365,N_5332,N_5131);
or U11366 (N_11366,N_9480,N_8434);
nor U11367 (N_11367,N_8381,N_6454);
xor U11368 (N_11368,N_6843,N_7439);
xnor U11369 (N_11369,N_8886,N_6678);
nand U11370 (N_11370,N_6833,N_7445);
and U11371 (N_11371,N_7334,N_5996);
or U11372 (N_11372,N_5836,N_6405);
nand U11373 (N_11373,N_5961,N_9248);
nor U11374 (N_11374,N_8441,N_8702);
nand U11375 (N_11375,N_9456,N_9719);
xnor U11376 (N_11376,N_8505,N_5520);
nor U11377 (N_11377,N_9035,N_8740);
nor U11378 (N_11378,N_5848,N_6732);
and U11379 (N_11379,N_5608,N_6762);
or U11380 (N_11380,N_9006,N_7089);
or U11381 (N_11381,N_9804,N_7630);
nor U11382 (N_11382,N_6530,N_6949);
nor U11383 (N_11383,N_7546,N_6917);
and U11384 (N_11384,N_6340,N_6958);
nand U11385 (N_11385,N_7508,N_9471);
or U11386 (N_11386,N_9534,N_9371);
nand U11387 (N_11387,N_5382,N_7953);
nor U11388 (N_11388,N_6459,N_9894);
and U11389 (N_11389,N_9323,N_7947);
nand U11390 (N_11390,N_8929,N_7964);
nand U11391 (N_11391,N_8041,N_8499);
and U11392 (N_11392,N_5779,N_6003);
xor U11393 (N_11393,N_5260,N_5658);
nor U11394 (N_11394,N_7935,N_9517);
nor U11395 (N_11395,N_7135,N_8186);
nor U11396 (N_11396,N_7580,N_9056);
and U11397 (N_11397,N_8651,N_5081);
and U11398 (N_11398,N_5896,N_5518);
or U11399 (N_11399,N_7596,N_9493);
and U11400 (N_11400,N_9421,N_7604);
and U11401 (N_11401,N_9681,N_8069);
xnor U11402 (N_11402,N_8600,N_6381);
nor U11403 (N_11403,N_5224,N_7877);
or U11404 (N_11404,N_5711,N_8788);
nand U11405 (N_11405,N_7866,N_6795);
nor U11406 (N_11406,N_7809,N_6496);
nor U11407 (N_11407,N_9823,N_5450);
xor U11408 (N_11408,N_9279,N_9506);
or U11409 (N_11409,N_8397,N_5240);
and U11410 (N_11410,N_5647,N_7984);
xnor U11411 (N_11411,N_8567,N_5156);
xnor U11412 (N_11412,N_7236,N_8987);
xnor U11413 (N_11413,N_5054,N_9971);
xor U11414 (N_11414,N_8523,N_5012);
xnor U11415 (N_11415,N_9994,N_8040);
and U11416 (N_11416,N_6778,N_7582);
nor U11417 (N_11417,N_7044,N_6040);
and U11418 (N_11418,N_6767,N_9807);
and U11419 (N_11419,N_6081,N_5652);
and U11420 (N_11420,N_9726,N_6019);
nand U11421 (N_11421,N_5216,N_7677);
or U11422 (N_11422,N_8013,N_9318);
nor U11423 (N_11423,N_6160,N_5138);
and U11424 (N_11424,N_8333,N_8616);
nand U11425 (N_11425,N_6937,N_5465);
nand U11426 (N_11426,N_6519,N_5828);
and U11427 (N_11427,N_5349,N_6839);
nand U11428 (N_11428,N_6827,N_9424);
or U11429 (N_11429,N_6016,N_6760);
nand U11430 (N_11430,N_7971,N_8507);
and U11431 (N_11431,N_9340,N_7178);
xnor U11432 (N_11432,N_6294,N_8096);
and U11433 (N_11433,N_6098,N_8486);
nor U11434 (N_11434,N_9801,N_9043);
nor U11435 (N_11435,N_5110,N_7101);
xnor U11436 (N_11436,N_6082,N_8603);
nand U11437 (N_11437,N_5856,N_5168);
nor U11438 (N_11438,N_8519,N_6735);
or U11439 (N_11439,N_9445,N_6493);
nor U11440 (N_11440,N_8732,N_9949);
and U11441 (N_11441,N_5230,N_6150);
or U11442 (N_11442,N_5696,N_8632);
or U11443 (N_11443,N_5623,N_8808);
nand U11444 (N_11444,N_9324,N_9623);
nand U11445 (N_11445,N_6492,N_6137);
and U11446 (N_11446,N_8818,N_8837);
or U11447 (N_11447,N_8547,N_6684);
nand U11448 (N_11448,N_8358,N_6701);
nand U11449 (N_11449,N_5018,N_7811);
and U11450 (N_11450,N_6331,N_9839);
xnor U11451 (N_11451,N_8572,N_5710);
or U11452 (N_11452,N_8185,N_6030);
nand U11453 (N_11453,N_5360,N_8265);
xor U11454 (N_11454,N_8391,N_8826);
nand U11455 (N_11455,N_6792,N_7151);
nand U11456 (N_11456,N_6526,N_8611);
nand U11457 (N_11457,N_6848,N_9903);
nor U11458 (N_11458,N_7855,N_6928);
nor U11459 (N_11459,N_9643,N_8209);
and U11460 (N_11460,N_5464,N_8918);
nor U11461 (N_11461,N_7848,N_5788);
or U11462 (N_11462,N_7659,N_8295);
or U11463 (N_11463,N_9895,N_8481);
nor U11464 (N_11464,N_9947,N_5289);
and U11465 (N_11465,N_5477,N_5565);
nor U11466 (N_11466,N_5530,N_7796);
xnor U11467 (N_11467,N_9796,N_8006);
nor U11468 (N_11468,N_5368,N_7856);
and U11469 (N_11469,N_5512,N_6179);
xor U11470 (N_11470,N_7057,N_8440);
nand U11471 (N_11471,N_7181,N_6305);
and U11472 (N_11472,N_5702,N_9712);
or U11473 (N_11473,N_6744,N_8016);
xor U11474 (N_11474,N_9873,N_6641);
xnor U11475 (N_11475,N_7908,N_7987);
nand U11476 (N_11476,N_5359,N_6092);
nand U11477 (N_11477,N_6540,N_8710);
nand U11478 (N_11478,N_6084,N_7482);
nor U11479 (N_11479,N_5371,N_9530);
or U11480 (N_11480,N_5433,N_6979);
nor U11481 (N_11481,N_9373,N_9521);
xor U11482 (N_11482,N_5540,N_6443);
nor U11483 (N_11483,N_6460,N_5676);
and U11484 (N_11484,N_7871,N_9960);
nor U11485 (N_11485,N_8285,N_6687);
nand U11486 (N_11486,N_8578,N_9527);
nand U11487 (N_11487,N_7005,N_6479);
or U11488 (N_11488,N_5663,N_9009);
nor U11489 (N_11489,N_8023,N_8083);
nor U11490 (N_11490,N_5451,N_6002);
and U11491 (N_11491,N_8844,N_5527);
or U11492 (N_11492,N_5307,N_8622);
nand U11493 (N_11493,N_7628,N_7476);
xnor U11494 (N_11494,N_6377,N_8584);
nand U11495 (N_11495,N_7411,N_7292);
xor U11496 (N_11496,N_8873,N_9977);
nor U11497 (N_11497,N_7196,N_5384);
or U11498 (N_11498,N_6269,N_8564);
and U11499 (N_11499,N_6431,N_6761);
or U11500 (N_11500,N_7810,N_6803);
nand U11501 (N_11501,N_8647,N_6577);
nor U11502 (N_11502,N_5184,N_9263);
or U11503 (N_11503,N_5668,N_9533);
nor U11504 (N_11504,N_5474,N_6772);
and U11505 (N_11505,N_7709,N_6888);
or U11506 (N_11506,N_8921,N_6484);
nor U11507 (N_11507,N_9428,N_6199);
nand U11508 (N_11508,N_7485,N_7506);
nand U11509 (N_11509,N_7164,N_8799);
nand U11510 (N_11510,N_7228,N_7605);
nor U11511 (N_11511,N_8175,N_7576);
and U11512 (N_11512,N_9637,N_9838);
xor U11513 (N_11513,N_7812,N_7087);
xnor U11514 (N_11514,N_9110,N_5965);
nor U11515 (N_11515,N_8250,N_9519);
nor U11516 (N_11516,N_5725,N_9758);
or U11517 (N_11517,N_8877,N_7385);
or U11518 (N_11518,N_9265,N_8245);
nor U11519 (N_11519,N_9676,N_8560);
nor U11520 (N_11520,N_9437,N_7350);
xnor U11521 (N_11521,N_8074,N_6284);
or U11522 (N_11522,N_7233,N_9773);
or U11523 (N_11523,N_9733,N_9227);
or U11524 (N_11524,N_6847,N_8368);
nand U11525 (N_11525,N_6038,N_6610);
xnor U11526 (N_11526,N_8119,N_7781);
or U11527 (N_11527,N_7642,N_9023);
nor U11528 (N_11528,N_5387,N_6464);
or U11529 (N_11529,N_8675,N_9888);
or U11530 (N_11530,N_9555,N_8389);
nor U11531 (N_11531,N_5900,N_6635);
xnor U11532 (N_11532,N_7730,N_6631);
or U11533 (N_11533,N_5291,N_9891);
nand U11534 (N_11534,N_5077,N_8851);
nor U11535 (N_11535,N_8527,N_9180);
nand U11536 (N_11536,N_7943,N_8522);
nand U11537 (N_11537,N_9254,N_6039);
or U11538 (N_11538,N_9364,N_9566);
and U11539 (N_11539,N_6710,N_5251);
xnor U11540 (N_11540,N_8136,N_5226);
nor U11541 (N_11541,N_5747,N_6455);
or U11542 (N_11542,N_5135,N_7795);
nand U11543 (N_11543,N_7997,N_9145);
and U11544 (N_11544,N_8672,N_7095);
and U11545 (N_11545,N_5423,N_6181);
or U11546 (N_11546,N_8402,N_9567);
nand U11547 (N_11547,N_7471,N_6424);
and U11548 (N_11548,N_6259,N_7830);
nand U11549 (N_11549,N_9274,N_7851);
or U11550 (N_11550,N_6819,N_8899);
nand U11551 (N_11551,N_9393,N_6812);
or U11552 (N_11552,N_9704,N_9753);
or U11553 (N_11553,N_7699,N_9415);
nor U11554 (N_11554,N_5777,N_6205);
nand U11555 (N_11555,N_6642,N_5050);
or U11556 (N_11556,N_8705,N_5124);
or U11557 (N_11557,N_6682,N_6978);
nand U11558 (N_11558,N_9870,N_7377);
nor U11559 (N_11559,N_8940,N_9251);
and U11560 (N_11560,N_9918,N_5510);
or U11561 (N_11561,N_8786,N_5091);
or U11562 (N_11562,N_5564,N_8099);
nor U11563 (N_11563,N_5921,N_9194);
nor U11564 (N_11564,N_6549,N_9216);
nor U11565 (N_11565,N_9847,N_9004);
nand U11566 (N_11566,N_7016,N_8957);
nand U11567 (N_11567,N_5771,N_6256);
or U11568 (N_11568,N_6970,N_7793);
or U11569 (N_11569,N_5059,N_7821);
and U11570 (N_11570,N_9946,N_8288);
nand U11571 (N_11571,N_6782,N_7152);
nor U11572 (N_11572,N_7670,N_5534);
nand U11573 (N_11573,N_5449,N_6146);
and U11574 (N_11574,N_6720,N_9492);
nand U11575 (N_11575,N_6861,N_5541);
nor U11576 (N_11576,N_6064,N_8466);
and U11577 (N_11577,N_5864,N_7692);
or U11578 (N_11578,N_6053,N_9889);
nand U11579 (N_11579,N_5118,N_6240);
nor U11580 (N_11580,N_8184,N_8276);
or U11581 (N_11581,N_9925,N_7472);
or U11582 (N_11582,N_7568,N_9411);
nor U11583 (N_11583,N_8648,N_9906);
nor U11584 (N_11584,N_9762,N_5715);
or U11585 (N_11585,N_7673,N_6465);
and U11586 (N_11586,N_8840,N_9601);
nand U11587 (N_11587,N_8321,N_9610);
and U11588 (N_11588,N_9228,N_9561);
xnor U11589 (N_11589,N_6807,N_8224);
nor U11590 (N_11590,N_7329,N_7450);
xnor U11591 (N_11591,N_7425,N_9221);
xor U11592 (N_11592,N_8494,N_7551);
nand U11593 (N_11593,N_6171,N_9938);
nand U11594 (N_11594,N_6442,N_7227);
or U11595 (N_11595,N_5238,N_5635);
nor U11596 (N_11596,N_9620,N_7311);
and U11597 (N_11597,N_5558,N_9115);
or U11598 (N_11598,N_7705,N_9982);
nor U11599 (N_11599,N_8392,N_7950);
or U11600 (N_11600,N_5661,N_9941);
xor U11601 (N_11601,N_6266,N_5614);
and U11602 (N_11602,N_8386,N_9398);
nor U11603 (N_11603,N_7218,N_6808);
xnor U11604 (N_11604,N_6236,N_8798);
or U11605 (N_11605,N_5458,N_8212);
nor U11606 (N_11606,N_8438,N_5660);
or U11607 (N_11607,N_9700,N_9299);
nor U11608 (N_11608,N_9147,N_6646);
nand U11609 (N_11609,N_9276,N_9116);
and U11610 (N_11610,N_9455,N_9811);
or U11611 (N_11611,N_9284,N_9586);
and U11612 (N_11612,N_8984,N_9735);
and U11613 (N_11613,N_5776,N_6037);
or U11614 (N_11614,N_6499,N_9000);
or U11615 (N_11615,N_8847,N_7167);
nand U11616 (N_11616,N_5933,N_6404);
and U11617 (N_11617,N_5641,N_6942);
or U11618 (N_11618,N_8613,N_6625);
xor U11619 (N_11619,N_5147,N_9377);
and U11620 (N_11620,N_8980,N_8687);
nor U11621 (N_11621,N_8592,N_5548);
and U11622 (N_11622,N_7687,N_7028);
or U11623 (N_11623,N_6822,N_9746);
nor U11624 (N_11624,N_5072,N_9749);
or U11625 (N_11625,N_5445,N_9273);
or U11626 (N_11626,N_7432,N_5529);
xnor U11627 (N_11627,N_9032,N_9435);
or U11628 (N_11628,N_7609,N_5325);
or U11629 (N_11629,N_5380,N_6594);
and U11630 (N_11630,N_6085,N_5320);
nor U11631 (N_11631,N_7801,N_6794);
xor U11632 (N_11632,N_5622,N_6576);
and U11633 (N_11633,N_9954,N_6225);
nor U11634 (N_11634,N_5627,N_8945);
or U11635 (N_11635,N_7241,N_8875);
nand U11636 (N_11636,N_9853,N_9500);
or U11637 (N_11637,N_5898,N_6587);
nor U11638 (N_11638,N_7183,N_5040);
nand U11639 (N_11639,N_7894,N_8057);
and U11640 (N_11640,N_9706,N_8404);
nand U11641 (N_11641,N_7895,N_7819);
and U11642 (N_11642,N_9907,N_8104);
nor U11643 (N_11643,N_9397,N_8998);
and U11644 (N_11644,N_8608,N_5144);
or U11645 (N_11645,N_9682,N_5806);
and U11646 (N_11646,N_8014,N_9912);
nor U11647 (N_11647,N_6875,N_8972);
nand U11648 (N_11648,N_9332,N_9105);
nand U11649 (N_11649,N_6142,N_7552);
nand U11650 (N_11650,N_5566,N_5273);
nand U11651 (N_11651,N_6321,N_7443);
nand U11652 (N_11652,N_5480,N_8251);
or U11653 (N_11653,N_8031,N_9467);
nor U11654 (N_11654,N_9654,N_9286);
or U11655 (N_11655,N_7215,N_7047);
nand U11656 (N_11656,N_7424,N_8767);
nand U11657 (N_11657,N_6948,N_7916);
or U11658 (N_11658,N_6922,N_9162);
and U11659 (N_11659,N_9598,N_6601);
nand U11660 (N_11660,N_8024,N_6660);
nor U11661 (N_11661,N_9562,N_5844);
and U11662 (N_11662,N_7076,N_9602);
and U11663 (N_11663,N_9898,N_8029);
and U11664 (N_11664,N_9739,N_8618);
and U11665 (N_11665,N_9789,N_6379);
nand U11666 (N_11666,N_7785,N_9862);
and U11667 (N_11667,N_9208,N_6554);
or U11668 (N_11668,N_7170,N_5646);
and U11669 (N_11669,N_8872,N_9886);
and U11670 (N_11670,N_8292,N_6602);
and U11671 (N_11671,N_6639,N_6197);
and U11672 (N_11672,N_6991,N_9969);
nand U11673 (N_11673,N_8990,N_8967);
or U11674 (N_11674,N_6351,N_7188);
xnor U11675 (N_11675,N_8180,N_6725);
nand U11676 (N_11676,N_6884,N_6615);
and U11677 (N_11677,N_7722,N_7634);
and U11678 (N_11678,N_5531,N_9452);
or U11679 (N_11679,N_8313,N_8384);
nand U11680 (N_11680,N_5748,N_6903);
xor U11681 (N_11681,N_7025,N_8064);
nand U11682 (N_11682,N_5753,N_9544);
and U11683 (N_11683,N_9570,N_6369);
and U11684 (N_11684,N_5364,N_7756);
or U11685 (N_11685,N_9112,N_5907);
or U11686 (N_11686,N_5886,N_9109);
or U11687 (N_11687,N_7789,N_8690);
and U11688 (N_11688,N_9959,N_8317);
nor U11689 (N_11689,N_9034,N_9952);
xnor U11690 (N_11690,N_7045,N_9551);
or U11691 (N_11691,N_9408,N_7620);
and U11692 (N_11692,N_7130,N_8049);
or U11693 (N_11693,N_6114,N_6945);
or U11694 (N_11694,N_7867,N_8134);
or U11695 (N_11695,N_8769,N_7977);
or U11696 (N_11696,N_5358,N_9854);
nor U11697 (N_11697,N_7608,N_8270);
and U11698 (N_11698,N_7431,N_6911);
nor U11699 (N_11699,N_8789,N_5145);
nor U11700 (N_11700,N_6315,N_6584);
nand U11701 (N_11701,N_8881,N_6716);
and U11702 (N_11702,N_7210,N_8601);
xnor U11703 (N_11703,N_8889,N_7754);
nand U11704 (N_11704,N_9447,N_5675);
and U11705 (N_11705,N_5628,N_5942);
and U11706 (N_11706,N_9063,N_7462);
or U11707 (N_11707,N_8070,N_7291);
nand U11708 (N_11708,N_9088,N_6043);
nand U11709 (N_11709,N_5883,N_7416);
nand U11710 (N_11710,N_5694,N_5094);
nor U11711 (N_11711,N_9309,N_6525);
or U11712 (N_11712,N_7097,N_9554);
nand U11713 (N_11713,N_7341,N_5109);
and U11714 (N_11714,N_9877,N_5250);
nand U11715 (N_11715,N_8413,N_7192);
or U11716 (N_11716,N_5021,N_8532);
and U11717 (N_11717,N_8483,N_8959);
or U11718 (N_11718,N_8079,N_9772);
nand U11719 (N_11719,N_8816,N_9699);
or U11720 (N_11720,N_6626,N_9123);
xnor U11721 (N_11721,N_6486,N_6025);
and U11722 (N_11722,N_7293,N_7155);
nor U11723 (N_11723,N_6028,N_6277);
nor U11724 (N_11724,N_7160,N_9619);
nand U11725 (N_11725,N_9908,N_7447);
and U11726 (N_11726,N_5323,N_7912);
and U11727 (N_11727,N_8842,N_8303);
or U11728 (N_11728,N_7297,N_7598);
xnor U11729 (N_11729,N_5316,N_9738);
or U11730 (N_11730,N_6768,N_9580);
nand U11731 (N_11731,N_5723,N_5052);
nand U11732 (N_11732,N_6797,N_6504);
nor U11733 (N_11733,N_6552,N_8588);
and U11734 (N_11734,N_7753,N_6550);
and U11735 (N_11735,N_5369,N_5957);
or U11736 (N_11736,N_8723,N_8411);
and U11737 (N_11737,N_9255,N_5223);
nand U11738 (N_11738,N_5471,N_9292);
or U11739 (N_11739,N_9885,N_9222);
nand U11740 (N_11740,N_7622,N_5552);
nand U11741 (N_11741,N_5472,N_7229);
nor U11742 (N_11742,N_9050,N_9531);
and U11743 (N_11743,N_6055,N_9582);
nand U11744 (N_11744,N_8653,N_7498);
nor U11745 (N_11745,N_5039,N_6899);
nand U11746 (N_11746,N_8595,N_6944);
xnor U11747 (N_11747,N_6823,N_8436);
nor U11748 (N_11748,N_8253,N_5507);
and U11749 (N_11749,N_7418,N_9402);
nor U11750 (N_11750,N_6298,N_5063);
and U11751 (N_11751,N_5304,N_5034);
nand U11752 (N_11752,N_6561,N_8033);
nor U11753 (N_11753,N_7042,N_5041);
nand U11754 (N_11754,N_9453,N_6629);
and U11755 (N_11755,N_8480,N_8239);
xor U11756 (N_11756,N_5922,N_6871);
nand U11757 (N_11757,N_7437,N_5533);
and U11758 (N_11758,N_7765,N_6165);
and U11759 (N_11759,N_9472,N_7578);
or U11760 (N_11760,N_5069,N_8063);
and U11761 (N_11761,N_7403,N_5305);
nor U11762 (N_11762,N_9342,N_6235);
or U11763 (N_11763,N_5000,N_6393);
and U11764 (N_11764,N_7905,N_9824);
nor U11765 (N_11765,N_8536,N_6966);
or U11766 (N_11766,N_8195,N_9029);
and U11767 (N_11767,N_8227,N_7693);
nor U11768 (N_11768,N_9603,N_9612);
nand U11769 (N_11769,N_9380,N_8794);
xnor U11770 (N_11770,N_6764,N_9515);
xor U11771 (N_11771,N_5221,N_8405);
nor U11772 (N_11772,N_8156,N_6352);
nand U11773 (N_11773,N_9242,N_9968);
or U11774 (N_11774,N_9594,N_6419);
xnor U11775 (N_11775,N_6880,N_9736);
nor U11776 (N_11776,N_5632,N_6776);
or U11777 (N_11777,N_6407,N_8230);
and U11778 (N_11778,N_5391,N_5503);
nand U11779 (N_11779,N_6283,N_6935);
nand U11780 (N_11780,N_8314,N_9851);
and U11781 (N_11781,N_5195,N_9465);
or U11782 (N_11782,N_5915,N_8464);
nor U11783 (N_11783,N_6453,N_7637);
nor U11784 (N_11784,N_8408,N_5008);
nand U11785 (N_11785,N_9587,N_6537);
nor U11786 (N_11786,N_9986,N_9757);
xnor U11787 (N_11787,N_8649,N_7231);
nand U11788 (N_11788,N_7059,N_9078);
nor U11789 (N_11789,N_5947,N_8985);
and U11790 (N_11790,N_6297,N_5105);
and U11791 (N_11791,N_9167,N_7723);
nor U11792 (N_11792,N_7541,N_6668);
nor U11793 (N_11793,N_7671,N_6959);
and U11794 (N_11794,N_7141,N_6151);
nor U11795 (N_11795,N_8934,N_8801);
nand U11796 (N_11796,N_5846,N_5448);
nor U11797 (N_11797,N_6981,N_6938);
nor U11798 (N_11798,N_5370,N_6745);
xnor U11799 (N_11799,N_6514,N_7127);
xnor U11800 (N_11800,N_9921,N_9717);
nor U11801 (N_11801,N_9483,N_7169);
nor U11802 (N_11802,N_7828,N_5811);
and U11803 (N_11803,N_6588,N_8660);
or U11804 (N_11804,N_5837,N_9926);
or U11805 (N_11805,N_8446,N_7222);
nor U11806 (N_11806,N_8357,N_7507);
or U11807 (N_11807,N_9550,N_6501);
nand U11808 (N_11808,N_8810,N_8487);
or U11809 (N_11809,N_9385,N_7296);
or U11810 (N_11810,N_6109,N_5244);
or U11811 (N_11811,N_9212,N_7743);
and U11812 (N_11812,N_5726,N_7761);
and U11813 (N_11813,N_9871,N_6763);
nand U11814 (N_11814,N_6758,N_9549);
nor U11815 (N_11815,N_6329,N_5719);
and U11816 (N_11816,N_6475,N_7212);
nand U11817 (N_11817,N_9927,N_5231);
nor U11818 (N_11818,N_6054,N_6212);
xnor U11819 (N_11819,N_7610,N_9765);
nor U11820 (N_11820,N_5444,N_9880);
nor U11821 (N_11821,N_6856,N_8751);
nor U11822 (N_11822,N_6508,N_9319);
or U11823 (N_11823,N_6791,N_7320);
and U11824 (N_11824,N_9974,N_8856);
nand U11825 (N_11825,N_7929,N_6196);
or U11826 (N_11826,N_6770,N_8091);
nor U11827 (N_11827,N_8114,N_8834);
nand U11828 (N_11828,N_9624,N_9219);
nand U11829 (N_11829,N_6946,N_8183);
nand U11830 (N_11830,N_8644,N_6335);
and U11831 (N_11831,N_6894,N_8315);
xor U11832 (N_11832,N_5256,N_7859);
and U11833 (N_11833,N_8068,N_8189);
xnor U11834 (N_11834,N_8496,N_8724);
xor U11835 (N_11835,N_9187,N_8641);
nand U11836 (N_11836,N_8072,N_7158);
and U11837 (N_11837,N_5232,N_5938);
xor U11838 (N_11838,N_7629,N_5177);
or U11839 (N_11839,N_6976,N_9646);
or U11840 (N_11840,N_8745,N_5362);
or U11841 (N_11841,N_6274,N_5294);
and U11842 (N_11842,N_8372,N_9425);
or U11843 (N_11843,N_7567,N_7434);
or U11844 (N_11844,N_9081,N_9277);
nand U11845 (N_11845,N_6089,N_7893);
and U11846 (N_11846,N_8750,N_5991);
nand U11847 (N_11847,N_8037,N_9900);
or U11848 (N_11848,N_9636,N_5048);
nand U11849 (N_11849,N_8467,N_6120);
and U11850 (N_11850,N_9038,N_9087);
or U11851 (N_11851,N_5193,N_9100);
nand U11852 (N_11852,N_5399,N_7521);
and U11853 (N_11853,N_7674,N_5909);
nor U11854 (N_11854,N_5268,N_8423);
nand U11855 (N_11855,N_9680,N_6401);
and U11856 (N_11856,N_9338,N_8546);
and U11857 (N_11857,N_8406,N_5010);
nor U11858 (N_11858,N_9642,N_6086);
nand U11859 (N_11859,N_7131,N_7398);
nand U11860 (N_11860,N_7006,N_8257);
and U11861 (N_11861,N_5425,N_6558);
nor U11862 (N_11862,N_8782,N_7501);
nor U11863 (N_11863,N_6018,N_8981);
nand U11864 (N_11864,N_7777,N_7638);
or U11865 (N_11865,N_7968,N_5338);
or U11866 (N_11866,N_9494,N_8058);
and U11867 (N_11867,N_5205,N_8232);
and U11868 (N_11868,N_6574,N_7664);
and U11869 (N_11869,N_6831,N_5334);
and U11870 (N_11870,N_8043,N_8850);
and U11871 (N_11871,N_8716,N_9658);
nor U11872 (N_11872,N_9224,N_5264);
and U11873 (N_11873,N_8993,N_5791);
nand U11874 (N_11874,N_9497,N_5926);
and U11875 (N_11875,N_5871,N_7651);
and U11876 (N_11876,N_6202,N_6515);
and U11877 (N_11877,N_6708,N_6061);
nor U11878 (N_11878,N_9709,N_5459);
nand U11879 (N_11879,N_9137,N_9503);
or U11880 (N_11880,N_5867,N_8458);
and U11881 (N_11881,N_9388,N_7844);
nor U11882 (N_11882,N_9988,N_6727);
or U11883 (N_11883,N_5677,N_8420);
xor U11884 (N_11884,N_6023,N_9366);
nor U11885 (N_11885,N_6677,N_9095);
and U11886 (N_11886,N_6751,N_5593);
and U11887 (N_11887,N_7077,N_7427);
or U11888 (N_11888,N_7448,N_6131);
xnor U11889 (N_11889,N_6260,N_5662);
or U11890 (N_11890,N_5612,N_5093);
nor U11891 (N_11891,N_5839,N_7543);
nor U11892 (N_11892,N_6990,N_7465);
nand U11893 (N_11893,N_5897,N_8518);
or U11894 (N_11894,N_8923,N_6873);
or U11895 (N_11895,N_8709,N_9662);
nor U11896 (N_11896,N_5917,N_5827);
nor U11897 (N_11897,N_8394,N_9327);
nor U11898 (N_11898,N_5379,N_6801);
nand U11899 (N_11899,N_9079,N_9152);
nor U11900 (N_11900,N_6434,N_9993);
or U11901 (N_11901,N_9556,N_9622);
nor U11902 (N_11902,N_7696,N_9444);
nor U11903 (N_11903,N_9632,N_8870);
nor U11904 (N_11904,N_9674,N_7381);
or U11905 (N_11905,N_8235,N_7989);
nand U11906 (N_11906,N_9731,N_7758);
or U11907 (N_11907,N_9463,N_7315);
nand U11908 (N_11908,N_9507,N_6482);
and U11909 (N_11909,N_5234,N_9383);
nor U11910 (N_11910,N_7114,N_7144);
and U11911 (N_11911,N_9014,N_7255);
and U11912 (N_11912,N_8289,N_8883);
xnor U11913 (N_11913,N_5966,N_5648);
or U11914 (N_11914,N_5206,N_9481);
and U11915 (N_11915,N_8473,N_9226);
or U11916 (N_11916,N_7058,N_8707);
and U11917 (N_11917,N_7179,N_8197);
or U11918 (N_11918,N_9822,N_9142);
nand U11919 (N_11919,N_8946,N_8625);
or U11920 (N_11920,N_6233,N_8193);
and U11921 (N_11921,N_7287,N_9427);
nor U11922 (N_11922,N_7085,N_9628);
xor U11923 (N_11923,N_7599,N_9396);
nor U11924 (N_11924,N_8639,N_8964);
or U11925 (N_11925,N_7586,N_6845);
nand U11926 (N_11926,N_6495,N_8269);
and U11927 (N_11927,N_8370,N_6187);
nor U11928 (N_11928,N_7180,N_8188);
or U11929 (N_11929,N_9564,N_6059);
or U11930 (N_11930,N_7353,N_7217);
xnor U11931 (N_11931,N_7123,N_5345);
nand U11932 (N_11932,N_6271,N_6263);
nand U11933 (N_11933,N_9121,N_9597);
nand U11934 (N_11934,N_7079,N_7774);
nand U11935 (N_11935,N_8054,N_9118);
and U11936 (N_11936,N_5309,N_5400);
and U11937 (N_11937,N_6457,N_6507);
nor U11938 (N_11938,N_9543,N_5067);
or U11939 (N_11939,N_5802,N_6851);
and U11940 (N_11940,N_6106,N_5191);
and U11941 (N_11941,N_8117,N_5029);
or U11942 (N_11942,N_9431,N_8828);
or U11943 (N_11943,N_9583,N_7666);
xor U11944 (N_11944,N_5980,N_6108);
or U11945 (N_11945,N_9440,N_6551);
nor U11946 (N_11946,N_8890,N_7373);
and U11947 (N_11947,N_5695,N_5123);
nor U11948 (N_11948,N_5188,N_5013);
nand U11949 (N_11949,N_5117,N_8217);
or U11950 (N_11950,N_6582,N_5087);
or U11951 (N_11951,N_8815,N_6467);
and U11952 (N_11952,N_5088,N_7102);
xnor U11953 (N_11953,N_7555,N_7590);
nand U11954 (N_11954,N_7993,N_7116);
and U11955 (N_11955,N_5280,N_8861);
and U11956 (N_11956,N_9019,N_5596);
or U11957 (N_11957,N_8540,N_5319);
xnor U11958 (N_11958,N_6889,N_9485);
or U11959 (N_11959,N_7050,N_7072);
nand U11960 (N_11960,N_8172,N_7375);
nor U11961 (N_11961,N_6301,N_9575);
or U11962 (N_11962,N_8971,N_5935);
xnor U11963 (N_11963,N_7140,N_8845);
nand U11964 (N_11964,N_9439,N_5643);
or U11965 (N_11965,N_8734,N_7825);
nor U11966 (N_11966,N_8501,N_5869);
and U11967 (N_11967,N_5978,N_8910);
nor U11968 (N_11968,N_9787,N_6698);
nor U11969 (N_11969,N_5290,N_8179);
or U11970 (N_11970,N_9064,N_5557);
nor U11971 (N_11971,N_8545,N_5288);
or U11972 (N_11972,N_7882,N_7356);
nor U11973 (N_11973,N_8621,N_9641);
nand U11974 (N_11974,N_9931,N_5528);
or U11975 (N_11975,N_8141,N_6983);
nand U11976 (N_11976,N_5051,N_8703);
xor U11977 (N_11977,N_9136,N_9904);
nand U11978 (N_11978,N_9538,N_8606);
and U11979 (N_11979,N_8576,N_6854);
nand U11980 (N_11980,N_8353,N_9183);
nand U11981 (N_11981,N_7211,N_6132);
or U11982 (N_11982,N_8610,N_8196);
xor U11983 (N_11983,N_6566,N_6841);
xnor U11984 (N_11984,N_6969,N_9141);
and U11985 (N_11985,N_8696,N_8375);
and U11986 (N_11986,N_6057,N_7845);
nand U11987 (N_11987,N_9631,N_6704);
and U11988 (N_11988,N_9420,N_8743);
nand U11989 (N_11989,N_8591,N_7257);
xor U11990 (N_11990,N_5667,N_8130);
nand U11991 (N_11991,N_5374,N_9074);
xor U11992 (N_11992,N_9953,N_7584);
or U11993 (N_11993,N_6145,N_7773);
nand U11994 (N_11994,N_7853,N_6052);
and U11995 (N_11995,N_9072,N_7656);
nor U11996 (N_11996,N_9955,N_6538);
nor U11997 (N_11997,N_7193,N_6752);
and U11998 (N_11998,N_5792,N_9540);
or U11999 (N_11999,N_7000,N_9329);
xnor U12000 (N_12000,N_7540,N_9459);
nor U12001 (N_12001,N_8355,N_9193);
and U12002 (N_12002,N_7833,N_8920);
or U12003 (N_12003,N_6569,N_8731);
nor U12004 (N_12004,N_9964,N_7748);
or U12005 (N_12005,N_9289,N_5283);
xnor U12006 (N_12006,N_7115,N_8403);
or U12007 (N_12007,N_7216,N_8200);
nor U12008 (N_12008,N_5097,N_8164);
or U12009 (N_12009,N_5789,N_7898);
and U12010 (N_12010,N_8151,N_8848);
nand U12011 (N_12011,N_9784,N_5984);
and U12012 (N_12012,N_6308,N_8082);
or U12013 (N_12013,N_9119,N_5971);
xnor U12014 (N_12014,N_9649,N_9833);
nor U12015 (N_12015,N_8308,N_9887);
or U12016 (N_12016,N_9498,N_9991);
nor U12017 (N_12017,N_8176,N_8385);
nor U12018 (N_12018,N_6251,N_9170);
xor U12019 (N_12019,N_6619,N_7782);
xor U12020 (N_12020,N_6934,N_9189);
nand U12021 (N_12021,N_6995,N_6886);
and U12022 (N_12022,N_9672,N_7583);
nor U12023 (N_12023,N_7967,N_7249);
xnor U12024 (N_12024,N_7278,N_5817);
nand U12025 (N_12025,N_7615,N_8960);
nor U12026 (N_12026,N_6154,N_5300);
nand U12027 (N_12027,N_6580,N_5001);
nand U12028 (N_12028,N_5624,N_5181);
and U12029 (N_12029,N_9367,N_8762);
or U12030 (N_12030,N_6399,N_5424);
xor U12031 (N_12031,N_7921,N_6630);
nand U12032 (N_12032,N_9300,N_7324);
nand U12033 (N_12033,N_5478,N_9611);
nand U12034 (N_12034,N_5149,N_8412);
xor U12035 (N_12035,N_6341,N_6383);
or U12036 (N_12036,N_5588,N_6214);
and U12037 (N_12037,N_6652,N_5479);
or U12038 (N_12038,N_8182,N_6141);
and U12039 (N_12039,N_8903,N_7475);
or U12040 (N_12040,N_7750,N_9281);
nor U12041 (N_12041,N_5700,N_7197);
or U12042 (N_12042,N_6810,N_9670);
nor U12043 (N_12043,N_7019,N_8166);
nor U12044 (N_12044,N_9899,N_6027);
and U12045 (N_12045,N_8966,N_6977);
and U12046 (N_12046,N_5333,N_8066);
xnor U12047 (N_12047,N_5735,N_6840);
nor U12048 (N_12048,N_7847,N_9653);
xnor U12049 (N_12049,N_6288,N_9893);
xnor U12050 (N_12050,N_7400,N_7360);
nand U12051 (N_12051,N_8359,N_7251);
or U12052 (N_12052,N_9406,N_8924);
nor U12053 (N_12053,N_5504,N_7880);
nor U12054 (N_12054,N_7525,N_8895);
nand U12055 (N_12055,N_9466,N_5730);
nand U12056 (N_12056,N_7768,N_5951);
nand U12057 (N_12057,N_5253,N_8824);
nor U12058 (N_12058,N_6347,N_7797);
nand U12059 (N_12059,N_9438,N_7467);
xor U12060 (N_12060,N_7589,N_5878);
or U12061 (N_12061,N_5681,N_7407);
nand U12062 (N_12062,N_5818,N_9935);
or U12063 (N_12063,N_9703,N_8667);
nand U12064 (N_12064,N_5201,N_6872);
nand U12065 (N_12065,N_6750,N_8448);
nand U12066 (N_12066,N_7680,N_7837);
nor U12067 (N_12067,N_5894,N_8008);
xor U12068 (N_12068,N_8936,N_7846);
nor U12069 (N_12069,N_5413,N_7787);
or U12070 (N_12070,N_6858,N_8223);
nand U12071 (N_12071,N_9290,N_9659);
and U12072 (N_12072,N_7736,N_8367);
nand U12073 (N_12073,N_8784,N_7449);
and U12074 (N_12074,N_6228,N_9374);
xnor U12075 (N_12075,N_9707,N_5522);
and U12076 (N_12076,N_6589,N_8661);
nor U12077 (N_12077,N_9488,N_5447);
xor U12078 (N_12078,N_6343,N_7949);
xor U12079 (N_12079,N_7083,N_8623);
or U12080 (N_12080,N_9781,N_9688);
nor U12081 (N_12081,N_7429,N_8469);
nor U12082 (N_12082,N_5706,N_9547);
nand U12083 (N_12083,N_8694,N_8234);
nor U12084 (N_12084,N_5047,N_5493);
nor U12085 (N_12085,N_5884,N_8342);
nor U12086 (N_12086,N_7813,N_7331);
and U12087 (N_12087,N_9914,N_8287);
xor U12088 (N_12088,N_5006,N_8698);
nand U12089 (N_12089,N_7878,N_7490);
nand U12090 (N_12090,N_8604,N_8018);
xor U12091 (N_12091,N_8841,N_5868);
nand U12092 (N_12092,N_7245,N_9131);
nor U12093 (N_12093,N_7133,N_6299);
nand U12094 (N_12094,N_9135,N_6740);
and U12095 (N_12095,N_5799,N_8866);
and U12096 (N_12096,N_6339,N_5427);
or U12097 (N_12097,N_5026,N_6815);
nor U12098 (N_12098,N_9369,N_9766);
nor U12099 (N_12099,N_8034,N_7234);
xnor U12100 (N_12100,N_9314,N_9764);
nand U12101 (N_12101,N_8506,N_6190);
and U12102 (N_12102,N_6998,N_7383);
or U12103 (N_12103,N_6989,N_8552);
or U12104 (N_12104,N_7776,N_5212);
nor U12105 (N_12105,N_7863,N_6448);
nand U12106 (N_12106,N_5625,N_5549);
nor U12107 (N_12107,N_9293,N_5476);
xnor U12108 (N_12108,N_8366,N_9021);
and U12109 (N_12109,N_5877,N_9320);
nor U12110 (N_12110,N_9235,N_7740);
nand U12111 (N_12111,N_7274,N_6346);
nor U12112 (N_12112,N_8047,N_7906);
nor U12113 (N_12113,N_9837,N_7150);
nor U12114 (N_12114,N_7235,N_6422);
and U12115 (N_12115,N_6590,N_9303);
nor U12116 (N_12116,N_6714,N_6358);
nor U12117 (N_12117,N_7899,N_8502);
nand U12118 (N_12118,N_6079,N_7505);
or U12119 (N_12119,N_6413,N_6451);
and U12120 (N_12120,N_6450,N_7191);
nor U12121 (N_12121,N_7344,N_7675);
or U12122 (N_12122,N_9669,N_6742);
nor U12123 (N_12123,N_5337,N_8530);
nor U12124 (N_12124,N_8833,N_9066);
and U12125 (N_12125,N_9860,N_7372);
nor U12126 (N_12126,N_9325,N_6219);
nor U12127 (N_12127,N_6391,N_7870);
and U12128 (N_12128,N_6252,N_8854);
nand U12129 (N_12129,N_6178,N_5532);
and U12130 (N_12130,N_5970,N_8362);
and U12131 (N_12131,N_8472,N_7557);
or U12132 (N_12132,N_8783,N_7107);
nor U12133 (N_12133,N_6489,N_6941);
or U12134 (N_12134,N_9093,N_5302);
or U12135 (N_12135,N_6907,N_7166);
and U12136 (N_12136,N_8051,N_5754);
or U12137 (N_12137,N_5729,N_6662);
nand U12138 (N_12138,N_7771,N_8718);
nor U12139 (N_12139,N_8811,N_7865);
or U12140 (N_12140,N_9294,N_8719);
and U12141 (N_12141,N_5102,N_8363);
and U12142 (N_12142,N_8901,N_5759);
or U12143 (N_12143,N_5489,N_9482);
nor U12144 (N_12144,N_6126,N_5543);
nand U12145 (N_12145,N_5159,N_6887);
nand U12146 (N_12146,N_9199,N_6166);
and U12147 (N_12147,N_8852,N_5949);
nor U12148 (N_12148,N_8339,N_6014);
nor U12149 (N_12149,N_5142,N_5967);
nand U12150 (N_12150,N_9560,N_8433);
and U12151 (N_12151,N_8558,N_9197);
or U12152 (N_12152,N_8757,N_9557);
or U12153 (N_12153,N_5772,N_8787);
or U12154 (N_12154,N_5918,N_5551);
or U12155 (N_12155,N_8445,N_9403);
or U12156 (N_12156,N_6314,N_7823);
nor U12157 (N_12157,N_7499,N_9913);
or U12158 (N_12158,N_7444,N_8293);
and U12159 (N_12159,N_8416,N_7868);
or U12160 (N_12160,N_6001,N_9321);
and U12161 (N_12161,N_8615,N_6332);
nor U12162 (N_12162,N_8214,N_5278);
and U12163 (N_12163,N_9132,N_6078);
nor U12164 (N_12164,N_8781,N_6388);
xnor U12165 (N_12165,N_9742,N_9565);
or U12166 (N_12166,N_8590,N_7563);
nand U12167 (N_12167,N_7979,N_5796);
or U12168 (N_12168,N_7975,N_9948);
and U12169 (N_12169,N_6416,N_7335);
and U12170 (N_12170,N_7408,N_5207);
nor U12171 (N_12171,N_8764,N_9211);
and U12172 (N_12172,N_7063,N_5372);
nor U12173 (N_12173,N_7137,N_8770);
or U12174 (N_12174,N_8274,N_7213);
or U12175 (N_12175,N_6105,N_8668);
and U12176 (N_12176,N_7832,N_9992);
or U12177 (N_12177,N_6403,N_5127);
and U12178 (N_12178,N_8349,N_7165);
xor U12179 (N_12179,N_8599,N_6906);
and U12180 (N_12180,N_7173,N_5415);
or U12181 (N_12181,N_7640,N_8098);
and U12182 (N_12182,N_5313,N_8271);
or U12183 (N_12183,N_6364,N_8577);
nand U12184 (N_12184,N_6497,N_7244);
xnor U12185 (N_12185,N_6470,N_6578);
nand U12186 (N_12186,N_8800,N_8712);
and U12187 (N_12187,N_7148,N_6022);
xor U12188 (N_12188,N_8145,N_7712);
or U12189 (N_12189,N_9863,N_7489);
or U12190 (N_12190,N_9042,N_6579);
or U12191 (N_12191,N_9091,N_5764);
nor U12192 (N_12192,N_8208,N_9846);
nor U12193 (N_12193,N_5554,N_7534);
or U12194 (N_12194,N_8264,N_6077);
or U12195 (N_12195,N_5801,N_7512);
and U12196 (N_12196,N_8556,N_5825);
nor U12197 (N_12197,N_5494,N_9233);
nand U12198 (N_12198,N_7413,N_5390);
and U12199 (N_12199,N_9400,N_8624);
nor U12200 (N_12200,N_9464,N_9458);
or U12201 (N_12201,N_9720,N_5017);
or U12202 (N_12202,N_9171,N_6999);
nand U12203 (N_12203,N_8831,N_9191);
nor U12204 (N_12204,N_9413,N_7481);
and U12205 (N_12205,N_9192,N_8765);
and U12206 (N_12206,N_5385,N_7569);
and U12207 (N_12207,N_5499,N_7572);
or U12208 (N_12208,N_7681,N_8462);
or U12209 (N_12209,N_6444,N_7665);
xnor U12210 (N_12210,N_5166,N_5634);
xor U12211 (N_12211,N_7300,N_7901);
or U12212 (N_12212,N_7053,N_9660);
and U12213 (N_12213,N_6925,N_8738);
xor U12214 (N_12214,N_6437,N_5602);
and U12215 (N_12215,N_6410,N_9285);
and U12216 (N_12216,N_5762,N_5411);
and U12217 (N_12217,N_7205,N_7338);
xor U12218 (N_12218,N_7650,N_8586);
nand U12219 (N_12219,N_6218,N_7548);
nor U12220 (N_12220,N_8379,N_8631);
and U12221 (N_12221,N_6285,N_5656);
nor U12222 (N_12222,N_8364,N_7468);
nor U12223 (N_12223,N_9687,N_5860);
nor U12224 (N_12224,N_6307,N_5033);
xor U12225 (N_12225,N_5011,N_5120);
or U12226 (N_12226,N_5213,N_5845);
nor U12227 (N_12227,N_8563,N_8426);
and U12228 (N_12228,N_9884,N_6956);
nor U12229 (N_12229,N_9599,N_5591);
or U12230 (N_12230,N_5461,N_7259);
or U12231 (N_12231,N_7254,N_6458);
nor U12232 (N_12232,N_5785,N_5286);
or U12233 (N_12233,N_5004,N_7132);
or U12234 (N_12234,N_6041,N_6723);
nor U12235 (N_12235,N_6924,N_9760);
or U12236 (N_12236,N_6712,N_5934);
nand U12237 (N_12237,N_6302,N_8562);
nand U12238 (N_12238,N_8094,N_8829);
or U12239 (N_12239,N_9568,N_7706);
and U12240 (N_12240,N_8073,N_5654);
and U12241 (N_12241,N_8015,N_8699);
and U12242 (N_12242,N_7012,N_7529);
or U12243 (N_12243,N_9755,N_6012);
xor U12244 (N_12244,N_7741,N_5393);
or U12245 (N_12245,N_6733,N_9999);
nand U12246 (N_12246,N_6291,N_9651);
nand U12247 (N_12247,N_5573,N_9315);
and U12248 (N_12248,N_6115,N_8030);
xnor U12249 (N_12249,N_6890,N_9103);
nand U12250 (N_12250,N_7611,N_6731);
or U12251 (N_12251,N_9272,N_8350);
and U12252 (N_12252,N_5755,N_9260);
nand U12253 (N_12253,N_6527,N_9354);
nor U12254 (N_12254,N_6143,N_5804);
or U12255 (N_12255,N_6940,N_5395);
nand U12256 (N_12256,N_7479,N_6908);
and U12257 (N_12257,N_8248,N_5813);
or U12258 (N_12258,N_6111,N_6534);
nor U12259 (N_12259,N_7176,N_9101);
and U12260 (N_12260,N_9107,N_9018);
and U12261 (N_12261,N_6697,N_7351);
nand U12262 (N_12262,N_7013,N_7014);
nor U12263 (N_12263,N_6326,N_9842);
nor U12264 (N_12264,N_9868,N_7613);
and U12265 (N_12265,N_9326,N_7384);
nand U12266 (N_12266,N_7035,N_5101);
or U12267 (N_12267,N_8820,N_6440);
nor U12268 (N_12268,N_7653,N_7902);
or U12269 (N_12269,N_5089,N_5388);
xnor U12270 (N_12270,N_8885,N_8730);
and U12271 (N_12271,N_9068,N_6759);
or U12272 (N_12272,N_8376,N_5023);
nor U12273 (N_12273,N_6533,N_8479);
or U12274 (N_12274,N_8325,N_7661);
nand U12275 (N_12275,N_8571,N_8220);
nand U12276 (N_12276,N_8316,N_7808);
and U12277 (N_12277,N_6786,N_6702);
or U12278 (N_12278,N_8247,N_8602);
nand U12279 (N_12279,N_6216,N_6546);
nor U12280 (N_12280,N_6070,N_8177);
xnor U12281 (N_12281,N_9698,N_6817);
and U12282 (N_12282,N_5501,N_5129);
or U12283 (N_12283,N_6756,N_5340);
and U12284 (N_12284,N_5595,N_5456);
or U12285 (N_12285,N_9268,N_6927);
nand U12286 (N_12286,N_6342,N_8001);
nand U12287 (N_12287,N_6051,N_7956);
or U12288 (N_12288,N_9098,N_8341);
xnor U12289 (N_12289,N_9901,N_6865);
nand U12290 (N_12290,N_9011,N_6182);
and U12291 (N_12291,N_5376,N_6221);
or U12292 (N_12292,N_6480,N_9686);
nand U12293 (N_12293,N_6008,N_8447);
and U12294 (N_12294,N_9609,N_6754);
nand U12295 (N_12295,N_8240,N_5794);
xor U12296 (N_12296,N_6091,N_9346);
or U12297 (N_12297,N_6882,N_9237);
and U12298 (N_12298,N_6323,N_7635);
or U12299 (N_12299,N_5111,N_8275);
nand U12300 (N_12300,N_5228,N_8231);
nand U12301 (N_12301,N_7308,N_7214);
nand U12302 (N_12302,N_8720,N_9502);
or U12303 (N_12303,N_7923,N_8863);
or U12304 (N_12304,N_7986,N_6366);
or U12305 (N_12305,N_9879,N_7084);
or U12306 (N_12306,N_9188,N_6101);
nand U12307 (N_12307,N_9301,N_6565);
or U12308 (N_12308,N_6200,N_7483);
and U12309 (N_12309,N_9395,N_7355);
and U12310 (N_12310,N_5876,N_5128);
nor U12311 (N_12311,N_8882,N_5100);
or U12312 (N_12312,N_5594,N_7374);
nor U12313 (N_12313,N_9711,N_9850);
xnor U12314 (N_12314,N_8544,N_7457);
or U12315 (N_12315,N_7060,N_8061);
or U12316 (N_12316,N_7807,N_7556);
nand U12317 (N_12317,N_7136,N_9422);
or U12318 (N_12318,N_9405,N_8643);
and U12319 (N_12319,N_7500,N_7910);
nand U12320 (N_12320,N_8427,N_5435);
or U12321 (N_12321,N_6707,N_7937);
xnor U12322 (N_12322,N_8111,N_5308);
nor U12323 (N_12323,N_6717,N_7718);
and U12324 (N_12324,N_9473,N_9605);
nor U12325 (N_12325,N_8891,N_9267);
nor U12326 (N_12326,N_7172,N_8331);
and U12327 (N_12327,N_8039,N_8332);
nand U12328 (N_12328,N_6556,N_5955);
nand U12329 (N_12329,N_8904,N_7105);
nor U12330 (N_12330,N_7223,N_6278);
or U12331 (N_12331,N_8582,N_8691);
or U12332 (N_12332,N_8471,N_5931);
xnor U12333 (N_12333,N_9548,N_6954);
nor U12334 (N_12334,N_5718,N_7978);
xor U12335 (N_12335,N_6734,N_8914);
and U12336 (N_12336,N_8999,N_9358);
or U12337 (N_12337,N_6446,N_7606);
xor U12338 (N_12338,N_5819,N_5408);
nand U12339 (N_12339,N_8149,N_6621);
or U12340 (N_12340,N_6042,N_9902);
and U12341 (N_12341,N_8241,N_7208);
or U12342 (N_12342,N_7252,N_8629);
nand U12343 (N_12343,N_6355,N_6705);
or U12344 (N_12344,N_7282,N_7528);
nor U12345 (N_12345,N_9243,N_6581);
nand U12346 (N_12346,N_7048,N_7841);
nor U12347 (N_12347,N_9416,N_5375);
and U12348 (N_12348,N_7571,N_9791);
nand U12349 (N_12349,N_5692,N_5524);
xnor U12350 (N_12350,N_9065,N_5277);
nand U12351 (N_12351,N_5592,N_6560);
xnor U12352 (N_12352,N_9771,N_8319);
nand U12353 (N_12353,N_6330,N_9668);
nor U12354 (N_12354,N_8311,N_6117);
nand U12355 (N_12355,N_6376,N_7719);
nand U12356 (N_12356,N_9965,N_7078);
nor U12357 (N_12357,N_9296,N_8680);
xnor U12358 (N_12358,N_8109,N_9667);
nor U12359 (N_12359,N_5152,N_9316);
nand U12360 (N_12360,N_9037,N_9756);
and U12361 (N_12361,N_5598,N_9710);
nor U12362 (N_12362,N_6065,N_8028);
or U12363 (N_12363,N_6261,N_8348);
nor U12364 (N_12364,N_6474,N_8722);
nand U12365 (N_12365,N_6674,N_9238);
or U12366 (N_12366,N_5899,N_8529);
and U12367 (N_12367,N_6013,N_5606);
and U12368 (N_12368,N_5161,N_8191);
nor U12369 (N_12369,N_6359,N_8424);
and U12370 (N_12370,N_7700,N_5310);
nand U12371 (N_12371,N_6234,N_6056);
and U12372 (N_12372,N_9245,N_6156);
and U12373 (N_12373,N_6557,N_5377);
or U12374 (N_12374,N_8110,N_7108);
and U12375 (N_12375,N_7240,N_7327);
xor U12376 (N_12376,N_6766,N_7607);
nand U12377 (N_12377,N_9146,N_9754);
nor U12378 (N_12378,N_5457,N_7139);
xnor U12379 (N_12379,N_7017,N_7295);
or U12380 (N_12380,N_7714,N_8170);
and U12381 (N_12381,N_6430,N_7745);
or U12382 (N_12382,N_7239,N_6072);
nand U12383 (N_12383,N_5150,N_8893);
and U12384 (N_12384,N_8450,N_7948);
or U12385 (N_12385,N_8674,N_9818);
and U12386 (N_12386,N_7243,N_8493);
nand U12387 (N_12387,N_9794,N_5840);
nor U12388 (N_12388,N_5367,N_9468);
or U12389 (N_12389,N_6473,N_7759);
nand U12390 (N_12390,N_5373,N_6553);
and U12391 (N_12391,N_6741,N_5601);
nand U12392 (N_12392,N_9835,N_9446);
nor U12393 (N_12393,N_5927,N_8165);
nor U12394 (N_12394,N_6414,N_8676);
nor U12395 (N_12395,N_9915,N_9962);
nand U12396 (N_12396,N_8216,N_6612);
or U12397 (N_12397,N_9775,N_6555);
nor U12398 (N_12398,N_5746,N_6921);
nand U12399 (N_12399,N_7138,N_7958);
or U12400 (N_12400,N_9978,N_5208);
and U12401 (N_12401,N_9577,N_8583);
and U12402 (N_12402,N_6636,N_9249);
or U12403 (N_12403,N_8925,N_9166);
xor U12404 (N_12404,N_7347,N_5519);
nand U12405 (N_12405,N_5266,N_5468);
or U12406 (N_12406,N_9372,N_8012);
nand U12407 (N_12407,N_8305,N_6930);
or U12408 (N_12408,N_7952,N_7348);
and U12409 (N_12409,N_8218,N_7382);
nor U12410 (N_12410,N_6005,N_6162);
xnor U12411 (N_12411,N_6058,N_5850);
nor U12412 (N_12412,N_7113,N_7995);
nand U12413 (N_12413,N_7738,N_8421);
or U12414 (N_12414,N_7892,N_7716);
or U12415 (N_12415,N_8888,N_9169);
nand U12416 (N_12416,N_7926,N_9808);
and U12417 (N_12417,N_7858,N_8587);
nor U12418 (N_12418,N_9563,N_9173);
nand U12419 (N_12419,N_7412,N_9552);
nor U12420 (N_12420,N_9089,N_8256);
xnor U12421 (N_12421,N_8161,N_9721);
and U12422 (N_12422,N_6353,N_9558);
and U12423 (N_12423,N_9634,N_7869);
nand U12424 (N_12424,N_5098,N_9812);
and U12425 (N_12425,N_7962,N_9748);
and U12426 (N_12426,N_6185,N_7093);
nand U12427 (N_12427,N_6706,N_9476);
xnor U12428 (N_12428,N_7038,N_7566);
nor U12429 (N_12429,N_7040,N_5936);
or U12430 (N_12430,N_8761,N_9341);
xnor U12431 (N_12431,N_9028,N_8541);
and U12432 (N_12432,N_7990,N_6231);
or U12433 (N_12433,N_6350,N_7020);
nor U12434 (N_12434,N_9196,N_9905);
xor U12435 (N_12435,N_7421,N_5215);
or U12436 (N_12436,N_8465,N_5095);
and U12437 (N_12437,N_9776,N_7288);
and U12438 (N_12438,N_9172,N_7161);
nor U12439 (N_12439,N_7262,N_5165);
nand U12440 (N_12440,N_7470,N_9866);
nor U12441 (N_12441,N_5112,N_6035);
nand U12442 (N_12442,N_8983,N_8963);
nand U12443 (N_12443,N_8101,N_6649);
nor U12444 (N_12444,N_5446,N_6510);
nand U12445 (N_12445,N_7533,N_8515);
nor U12446 (N_12446,N_8974,N_9049);
and U12447 (N_12447,N_8459,N_7791);
or U12448 (N_12448,N_5453,N_6608);
nor U12449 (N_12449,N_6695,N_7928);
nand U12450 (N_12450,N_6372,N_8952);
nor U12451 (N_12451,N_5990,N_6397);
xnor U12452 (N_12452,N_5352,N_7343);
nand U12453 (N_12453,N_7182,N_6699);
nor U12454 (N_12454,N_8689,N_8442);
xor U12455 (N_12455,N_6375,N_5275);
nor U12456 (N_12456,N_6564,N_6623);
nand U12457 (N_12457,N_9910,N_5665);
xnor U12458 (N_12458,N_8554,N_5649);
or U12459 (N_12459,N_6046,N_5576);
nand U12460 (N_12460,N_5630,N_6748);
nand U12461 (N_12461,N_9664,N_6135);
or U12462 (N_12462,N_7246,N_8790);
nor U12463 (N_12463,N_6620,N_9288);
nand U12464 (N_12464,N_9961,N_5407);
nor U12465 (N_12465,N_9390,N_6322);
or U12466 (N_12466,N_5363,N_5609);
and U12467 (N_12467,N_8118,N_9205);
and U12468 (N_12468,N_7518,N_5058);
or U12469 (N_12469,N_9442,N_9076);
and U12470 (N_12470,N_6247,N_7401);
and U12471 (N_12471,N_7966,N_8382);
nor U12472 (N_12472,N_7323,N_8115);
and U12473 (N_12473,N_6932,N_7547);
and U12474 (N_12474,N_8673,N_6161);
nand U12475 (N_12475,N_9247,N_9040);
xnor U12476 (N_12476,N_5121,N_8646);
or U12477 (N_12477,N_6933,N_7422);
or U12478 (N_12478,N_9647,N_8263);
nand U12479 (N_12479,N_8776,N_9015);
or U12480 (N_12480,N_6122,N_5857);
and U12481 (N_12481,N_7065,N_9041);
xor U12482 (N_12482,N_9701,N_8320);
xor U12483 (N_12483,N_8879,N_8569);
nor U12484 (N_12484,N_9048,N_8206);
nand U12485 (N_12485,N_6469,N_7535);
nor U12486 (N_12486,N_8656,N_7924);
nor U12487 (N_12487,N_5164,N_6306);
xor U12488 (N_12488,N_6753,N_9677);
nand U12489 (N_12489,N_8520,N_6909);
nand U12490 (N_12490,N_6466,N_5298);
and U12491 (N_12491,N_7824,N_6194);
xor U12492 (N_12492,N_9352,N_9376);
and U12493 (N_12493,N_6645,N_8874);
nand U12494 (N_12494,N_9218,N_7660);
xnor U12495 (N_12495,N_7802,N_5343);
nand U12496 (N_12496,N_8747,N_5514);
and U12497 (N_12497,N_8346,N_5140);
xnor U12498 (N_12498,N_7455,N_6681);
and U12499 (N_12499,N_8821,N_6798);
nand U12500 (N_12500,N_7237,N_6082);
or U12501 (N_12501,N_6390,N_6077);
and U12502 (N_12502,N_6730,N_6423);
or U12503 (N_12503,N_6553,N_8932);
nor U12504 (N_12504,N_6701,N_7053);
nand U12505 (N_12505,N_5326,N_6345);
or U12506 (N_12506,N_6976,N_9522);
and U12507 (N_12507,N_7254,N_7151);
nand U12508 (N_12508,N_6633,N_9750);
nor U12509 (N_12509,N_8438,N_7654);
nand U12510 (N_12510,N_8973,N_7671);
or U12511 (N_12511,N_9382,N_9549);
nand U12512 (N_12512,N_5280,N_8975);
and U12513 (N_12513,N_7696,N_9075);
and U12514 (N_12514,N_7906,N_7264);
nor U12515 (N_12515,N_9854,N_5609);
nand U12516 (N_12516,N_9009,N_7353);
and U12517 (N_12517,N_5535,N_9764);
nand U12518 (N_12518,N_5985,N_7010);
or U12519 (N_12519,N_5260,N_7633);
nor U12520 (N_12520,N_6402,N_5472);
and U12521 (N_12521,N_5078,N_6809);
nand U12522 (N_12522,N_8405,N_5337);
nand U12523 (N_12523,N_9680,N_5120);
nor U12524 (N_12524,N_9558,N_9228);
xor U12525 (N_12525,N_9807,N_8373);
or U12526 (N_12526,N_7403,N_7470);
and U12527 (N_12527,N_7276,N_5807);
xor U12528 (N_12528,N_8662,N_5297);
nand U12529 (N_12529,N_5871,N_6665);
or U12530 (N_12530,N_7358,N_6076);
nand U12531 (N_12531,N_8934,N_7892);
xor U12532 (N_12532,N_9018,N_6279);
nand U12533 (N_12533,N_6136,N_5297);
nor U12534 (N_12534,N_7703,N_8198);
or U12535 (N_12535,N_5897,N_8208);
nor U12536 (N_12536,N_6780,N_6752);
or U12537 (N_12537,N_7193,N_6581);
or U12538 (N_12538,N_9067,N_9642);
nor U12539 (N_12539,N_7904,N_5554);
xor U12540 (N_12540,N_7081,N_7566);
and U12541 (N_12541,N_5737,N_7739);
xnor U12542 (N_12542,N_7828,N_8278);
or U12543 (N_12543,N_9600,N_5415);
nor U12544 (N_12544,N_8462,N_6885);
nor U12545 (N_12545,N_5415,N_6266);
or U12546 (N_12546,N_6107,N_6017);
nor U12547 (N_12547,N_7912,N_9767);
nand U12548 (N_12548,N_9889,N_8985);
nor U12549 (N_12549,N_6930,N_8884);
nand U12550 (N_12550,N_5583,N_5218);
nand U12551 (N_12551,N_6771,N_5403);
and U12552 (N_12552,N_7548,N_8938);
or U12553 (N_12553,N_7766,N_5544);
nand U12554 (N_12554,N_8822,N_8672);
or U12555 (N_12555,N_7020,N_7656);
or U12556 (N_12556,N_6154,N_5772);
and U12557 (N_12557,N_7603,N_6691);
xnor U12558 (N_12558,N_6784,N_8073);
nor U12559 (N_12559,N_8825,N_5720);
and U12560 (N_12560,N_7574,N_8566);
or U12561 (N_12561,N_9808,N_7082);
or U12562 (N_12562,N_7380,N_5570);
or U12563 (N_12563,N_9060,N_8090);
nor U12564 (N_12564,N_5354,N_9453);
and U12565 (N_12565,N_9391,N_9364);
and U12566 (N_12566,N_5994,N_8849);
nand U12567 (N_12567,N_5977,N_5128);
xnor U12568 (N_12568,N_6917,N_7331);
nor U12569 (N_12569,N_8532,N_7979);
and U12570 (N_12570,N_6733,N_7497);
nor U12571 (N_12571,N_5112,N_5702);
and U12572 (N_12572,N_9042,N_9950);
xor U12573 (N_12573,N_9856,N_7409);
nand U12574 (N_12574,N_5909,N_6131);
and U12575 (N_12575,N_8733,N_5365);
or U12576 (N_12576,N_5306,N_7832);
and U12577 (N_12577,N_6973,N_5546);
or U12578 (N_12578,N_9763,N_9259);
nor U12579 (N_12579,N_6917,N_5981);
nor U12580 (N_12580,N_9578,N_9981);
nand U12581 (N_12581,N_8998,N_6568);
nor U12582 (N_12582,N_6622,N_9453);
nand U12583 (N_12583,N_5831,N_5474);
nor U12584 (N_12584,N_9836,N_9825);
xor U12585 (N_12585,N_8035,N_7565);
xnor U12586 (N_12586,N_7384,N_6209);
nand U12587 (N_12587,N_6656,N_6324);
nand U12588 (N_12588,N_5311,N_9299);
and U12589 (N_12589,N_5147,N_9623);
or U12590 (N_12590,N_6527,N_5962);
xnor U12591 (N_12591,N_7231,N_7521);
nand U12592 (N_12592,N_8252,N_6986);
or U12593 (N_12593,N_8238,N_5480);
nor U12594 (N_12594,N_7442,N_8741);
nor U12595 (N_12595,N_8337,N_9947);
nand U12596 (N_12596,N_6096,N_7555);
nand U12597 (N_12597,N_8218,N_9503);
nor U12598 (N_12598,N_6872,N_7972);
or U12599 (N_12599,N_8408,N_5943);
nor U12600 (N_12600,N_7216,N_6360);
or U12601 (N_12601,N_6583,N_5603);
xnor U12602 (N_12602,N_6611,N_9883);
and U12603 (N_12603,N_5096,N_7061);
and U12604 (N_12604,N_5707,N_5506);
or U12605 (N_12605,N_8850,N_6027);
nand U12606 (N_12606,N_6189,N_7902);
and U12607 (N_12607,N_9892,N_9574);
and U12608 (N_12608,N_7934,N_9458);
or U12609 (N_12609,N_9125,N_8775);
nand U12610 (N_12610,N_9954,N_5133);
and U12611 (N_12611,N_6786,N_8844);
nand U12612 (N_12612,N_5601,N_6321);
nand U12613 (N_12613,N_7586,N_5247);
nand U12614 (N_12614,N_6714,N_9748);
or U12615 (N_12615,N_9197,N_6990);
nor U12616 (N_12616,N_7317,N_8946);
nand U12617 (N_12617,N_9519,N_5335);
nand U12618 (N_12618,N_7075,N_7055);
xor U12619 (N_12619,N_8936,N_7014);
or U12620 (N_12620,N_7758,N_7645);
or U12621 (N_12621,N_7997,N_8736);
and U12622 (N_12622,N_9925,N_8343);
nand U12623 (N_12623,N_6722,N_5809);
or U12624 (N_12624,N_6319,N_6861);
nand U12625 (N_12625,N_8894,N_8289);
nand U12626 (N_12626,N_5070,N_7882);
nor U12627 (N_12627,N_7541,N_6146);
and U12628 (N_12628,N_7142,N_5930);
nor U12629 (N_12629,N_6603,N_6610);
and U12630 (N_12630,N_9260,N_9202);
and U12631 (N_12631,N_5683,N_6507);
or U12632 (N_12632,N_8827,N_8435);
or U12633 (N_12633,N_6704,N_5732);
nand U12634 (N_12634,N_9421,N_8663);
and U12635 (N_12635,N_5499,N_9985);
nor U12636 (N_12636,N_5547,N_5974);
nand U12637 (N_12637,N_9387,N_9033);
and U12638 (N_12638,N_6077,N_8850);
nor U12639 (N_12639,N_5814,N_5850);
and U12640 (N_12640,N_6072,N_7437);
and U12641 (N_12641,N_7161,N_8554);
and U12642 (N_12642,N_6631,N_9029);
xor U12643 (N_12643,N_7413,N_7314);
nand U12644 (N_12644,N_8672,N_6741);
xnor U12645 (N_12645,N_6484,N_5717);
and U12646 (N_12646,N_8057,N_7583);
or U12647 (N_12647,N_7418,N_8784);
or U12648 (N_12648,N_5141,N_6116);
xor U12649 (N_12649,N_5740,N_6730);
nand U12650 (N_12650,N_6653,N_5645);
nand U12651 (N_12651,N_6169,N_7624);
xnor U12652 (N_12652,N_5401,N_6175);
and U12653 (N_12653,N_7362,N_7739);
or U12654 (N_12654,N_9476,N_8068);
nor U12655 (N_12655,N_7606,N_9421);
and U12656 (N_12656,N_9637,N_7142);
and U12657 (N_12657,N_9984,N_9125);
nor U12658 (N_12658,N_5745,N_5289);
xnor U12659 (N_12659,N_6868,N_5695);
xor U12660 (N_12660,N_9806,N_6267);
xor U12661 (N_12661,N_8220,N_5244);
or U12662 (N_12662,N_9436,N_9022);
and U12663 (N_12663,N_8452,N_9819);
or U12664 (N_12664,N_7498,N_9516);
nand U12665 (N_12665,N_5703,N_7661);
nand U12666 (N_12666,N_5816,N_7052);
xor U12667 (N_12667,N_5957,N_8795);
nand U12668 (N_12668,N_9986,N_5056);
nand U12669 (N_12669,N_6624,N_7308);
xnor U12670 (N_12670,N_9556,N_7626);
nand U12671 (N_12671,N_8323,N_6316);
nor U12672 (N_12672,N_7295,N_5379);
nor U12673 (N_12673,N_7864,N_9045);
xnor U12674 (N_12674,N_5926,N_6545);
and U12675 (N_12675,N_5213,N_7723);
and U12676 (N_12676,N_8558,N_7954);
nand U12677 (N_12677,N_9540,N_8581);
nor U12678 (N_12678,N_5358,N_5361);
nor U12679 (N_12679,N_5618,N_7957);
or U12680 (N_12680,N_9739,N_5475);
nor U12681 (N_12681,N_6090,N_5022);
nand U12682 (N_12682,N_5161,N_8453);
xnor U12683 (N_12683,N_5578,N_8585);
xnor U12684 (N_12684,N_9153,N_8364);
nand U12685 (N_12685,N_7724,N_8027);
and U12686 (N_12686,N_5706,N_6200);
nor U12687 (N_12687,N_9474,N_7209);
nand U12688 (N_12688,N_8152,N_6524);
xnor U12689 (N_12689,N_9697,N_6840);
nor U12690 (N_12690,N_5779,N_8791);
nor U12691 (N_12691,N_8359,N_5996);
nor U12692 (N_12692,N_8862,N_5434);
nor U12693 (N_12693,N_9503,N_5520);
nand U12694 (N_12694,N_6003,N_8542);
and U12695 (N_12695,N_9371,N_5980);
nor U12696 (N_12696,N_7126,N_8928);
nor U12697 (N_12697,N_5468,N_6613);
or U12698 (N_12698,N_9947,N_9642);
and U12699 (N_12699,N_9237,N_8793);
nor U12700 (N_12700,N_7807,N_6384);
nand U12701 (N_12701,N_7578,N_7711);
nand U12702 (N_12702,N_7227,N_7601);
and U12703 (N_12703,N_7846,N_9115);
or U12704 (N_12704,N_8789,N_9412);
nor U12705 (N_12705,N_6853,N_8968);
nand U12706 (N_12706,N_7944,N_6056);
or U12707 (N_12707,N_8625,N_9552);
nand U12708 (N_12708,N_8398,N_5871);
or U12709 (N_12709,N_9803,N_6184);
or U12710 (N_12710,N_8747,N_7296);
and U12711 (N_12711,N_7129,N_7263);
and U12712 (N_12712,N_8693,N_5181);
and U12713 (N_12713,N_5096,N_9100);
and U12714 (N_12714,N_6986,N_5636);
nand U12715 (N_12715,N_9006,N_5236);
nor U12716 (N_12716,N_5938,N_7233);
nor U12717 (N_12717,N_9655,N_5805);
or U12718 (N_12718,N_6945,N_8601);
or U12719 (N_12719,N_8317,N_6742);
or U12720 (N_12720,N_9049,N_9282);
xor U12721 (N_12721,N_8410,N_9826);
nand U12722 (N_12722,N_7359,N_5928);
or U12723 (N_12723,N_9801,N_5608);
nor U12724 (N_12724,N_9082,N_6378);
xor U12725 (N_12725,N_5471,N_6728);
nor U12726 (N_12726,N_9576,N_7725);
or U12727 (N_12727,N_5634,N_9309);
and U12728 (N_12728,N_8329,N_7733);
xor U12729 (N_12729,N_7657,N_5121);
nor U12730 (N_12730,N_6883,N_8524);
and U12731 (N_12731,N_7733,N_9588);
xor U12732 (N_12732,N_7835,N_8133);
nor U12733 (N_12733,N_8305,N_7553);
and U12734 (N_12734,N_5530,N_8288);
xor U12735 (N_12735,N_5156,N_9236);
nor U12736 (N_12736,N_6578,N_9898);
or U12737 (N_12737,N_6262,N_8144);
xnor U12738 (N_12738,N_8110,N_6560);
nor U12739 (N_12739,N_9541,N_7423);
or U12740 (N_12740,N_8881,N_6775);
nor U12741 (N_12741,N_6373,N_7147);
nand U12742 (N_12742,N_8619,N_6310);
nor U12743 (N_12743,N_5240,N_7784);
or U12744 (N_12744,N_5613,N_7050);
nor U12745 (N_12745,N_6566,N_9023);
nand U12746 (N_12746,N_9033,N_6270);
nand U12747 (N_12747,N_6675,N_8259);
nand U12748 (N_12748,N_5483,N_5868);
nand U12749 (N_12749,N_9036,N_9601);
nor U12750 (N_12750,N_9121,N_6953);
or U12751 (N_12751,N_9438,N_5200);
nor U12752 (N_12752,N_6301,N_5626);
nand U12753 (N_12753,N_5877,N_9850);
or U12754 (N_12754,N_5626,N_5260);
xnor U12755 (N_12755,N_6179,N_5280);
nor U12756 (N_12756,N_9287,N_9264);
nand U12757 (N_12757,N_8639,N_6669);
nand U12758 (N_12758,N_5436,N_8289);
xnor U12759 (N_12759,N_9413,N_5193);
and U12760 (N_12760,N_8200,N_9011);
nand U12761 (N_12761,N_9343,N_7046);
or U12762 (N_12762,N_7511,N_7790);
or U12763 (N_12763,N_9827,N_6617);
xnor U12764 (N_12764,N_8900,N_7853);
or U12765 (N_12765,N_8644,N_9447);
nand U12766 (N_12766,N_7526,N_9351);
nor U12767 (N_12767,N_7020,N_6981);
nand U12768 (N_12768,N_9531,N_6216);
or U12769 (N_12769,N_5735,N_7100);
nor U12770 (N_12770,N_5485,N_9568);
nand U12771 (N_12771,N_9558,N_8836);
nand U12772 (N_12772,N_6870,N_9225);
or U12773 (N_12773,N_8075,N_6367);
nand U12774 (N_12774,N_5093,N_9220);
nand U12775 (N_12775,N_5586,N_6487);
or U12776 (N_12776,N_8860,N_8831);
and U12777 (N_12777,N_5170,N_6644);
nand U12778 (N_12778,N_5157,N_5260);
nand U12779 (N_12779,N_5009,N_7034);
xor U12780 (N_12780,N_7996,N_9564);
and U12781 (N_12781,N_8458,N_5662);
or U12782 (N_12782,N_5067,N_7079);
nor U12783 (N_12783,N_5149,N_8067);
and U12784 (N_12784,N_5148,N_9286);
and U12785 (N_12785,N_9461,N_6196);
or U12786 (N_12786,N_9315,N_7097);
xor U12787 (N_12787,N_5306,N_5212);
xnor U12788 (N_12788,N_8360,N_5155);
nand U12789 (N_12789,N_5612,N_9049);
xor U12790 (N_12790,N_8241,N_6030);
nand U12791 (N_12791,N_9079,N_6722);
nor U12792 (N_12792,N_7778,N_9985);
xor U12793 (N_12793,N_7270,N_6229);
or U12794 (N_12794,N_5371,N_8069);
xnor U12795 (N_12795,N_5459,N_9927);
and U12796 (N_12796,N_9427,N_6623);
and U12797 (N_12797,N_9972,N_5415);
nor U12798 (N_12798,N_5772,N_9051);
or U12799 (N_12799,N_7336,N_9797);
nor U12800 (N_12800,N_9227,N_5265);
nand U12801 (N_12801,N_8592,N_6925);
nor U12802 (N_12802,N_9234,N_8040);
nor U12803 (N_12803,N_9953,N_6780);
and U12804 (N_12804,N_6601,N_5695);
or U12805 (N_12805,N_6124,N_9272);
nand U12806 (N_12806,N_7817,N_5508);
or U12807 (N_12807,N_5233,N_5945);
xnor U12808 (N_12808,N_7392,N_9385);
and U12809 (N_12809,N_5402,N_6449);
xnor U12810 (N_12810,N_6858,N_7726);
nand U12811 (N_12811,N_7874,N_9640);
nand U12812 (N_12812,N_7013,N_8882);
nor U12813 (N_12813,N_7605,N_9105);
nand U12814 (N_12814,N_6497,N_8116);
or U12815 (N_12815,N_9605,N_7486);
or U12816 (N_12816,N_9260,N_6727);
nor U12817 (N_12817,N_5801,N_8308);
and U12818 (N_12818,N_7824,N_7755);
xor U12819 (N_12819,N_9178,N_6832);
nor U12820 (N_12820,N_5265,N_7295);
nand U12821 (N_12821,N_8496,N_5769);
nand U12822 (N_12822,N_6589,N_6967);
and U12823 (N_12823,N_8228,N_5351);
or U12824 (N_12824,N_9542,N_7437);
nand U12825 (N_12825,N_7699,N_7934);
and U12826 (N_12826,N_9940,N_7202);
xor U12827 (N_12827,N_7186,N_7657);
or U12828 (N_12828,N_5306,N_7715);
nor U12829 (N_12829,N_6898,N_9629);
and U12830 (N_12830,N_6590,N_6389);
xnor U12831 (N_12831,N_7532,N_8754);
or U12832 (N_12832,N_8563,N_9345);
nor U12833 (N_12833,N_7044,N_7421);
and U12834 (N_12834,N_7402,N_5633);
or U12835 (N_12835,N_5404,N_6856);
nand U12836 (N_12836,N_5725,N_6562);
nand U12837 (N_12837,N_9025,N_7878);
and U12838 (N_12838,N_7448,N_5851);
nor U12839 (N_12839,N_6055,N_8914);
and U12840 (N_12840,N_7434,N_8208);
nand U12841 (N_12841,N_5613,N_5219);
xor U12842 (N_12842,N_5458,N_9978);
or U12843 (N_12843,N_8765,N_6090);
and U12844 (N_12844,N_8623,N_5360);
and U12845 (N_12845,N_6809,N_9975);
and U12846 (N_12846,N_6111,N_7671);
or U12847 (N_12847,N_8014,N_7397);
nor U12848 (N_12848,N_6021,N_6011);
and U12849 (N_12849,N_8328,N_8687);
nand U12850 (N_12850,N_6282,N_8309);
nand U12851 (N_12851,N_6534,N_5078);
nor U12852 (N_12852,N_8121,N_6579);
and U12853 (N_12853,N_6212,N_6327);
and U12854 (N_12854,N_5713,N_8243);
and U12855 (N_12855,N_9921,N_9925);
or U12856 (N_12856,N_8276,N_5705);
nand U12857 (N_12857,N_9580,N_7156);
xnor U12858 (N_12858,N_5901,N_8745);
nor U12859 (N_12859,N_5486,N_7851);
or U12860 (N_12860,N_8707,N_6564);
nand U12861 (N_12861,N_8202,N_8394);
nor U12862 (N_12862,N_6488,N_8795);
nor U12863 (N_12863,N_6159,N_9387);
and U12864 (N_12864,N_8499,N_8922);
and U12865 (N_12865,N_7808,N_6357);
nand U12866 (N_12866,N_5511,N_5101);
and U12867 (N_12867,N_5681,N_9294);
nor U12868 (N_12868,N_8435,N_5874);
nor U12869 (N_12869,N_7428,N_6087);
nor U12870 (N_12870,N_5745,N_7485);
nand U12871 (N_12871,N_5440,N_5180);
nor U12872 (N_12872,N_5914,N_5666);
nor U12873 (N_12873,N_7637,N_8049);
xor U12874 (N_12874,N_6682,N_8106);
nor U12875 (N_12875,N_5440,N_8520);
or U12876 (N_12876,N_7212,N_7917);
nor U12877 (N_12877,N_9121,N_6907);
or U12878 (N_12878,N_6027,N_7214);
nand U12879 (N_12879,N_7121,N_6512);
nor U12880 (N_12880,N_9498,N_5006);
nand U12881 (N_12881,N_9516,N_7821);
nand U12882 (N_12882,N_7962,N_7689);
or U12883 (N_12883,N_7887,N_6136);
nor U12884 (N_12884,N_8244,N_5727);
nand U12885 (N_12885,N_7734,N_8462);
or U12886 (N_12886,N_7919,N_7382);
nand U12887 (N_12887,N_8203,N_8376);
nand U12888 (N_12888,N_9443,N_8835);
xor U12889 (N_12889,N_5230,N_8016);
nand U12890 (N_12890,N_9747,N_6646);
xor U12891 (N_12891,N_6410,N_5047);
and U12892 (N_12892,N_7976,N_6264);
or U12893 (N_12893,N_5439,N_8401);
xnor U12894 (N_12894,N_6736,N_7899);
and U12895 (N_12895,N_5368,N_5974);
nor U12896 (N_12896,N_9985,N_6089);
xor U12897 (N_12897,N_6689,N_8789);
nand U12898 (N_12898,N_8184,N_6123);
nand U12899 (N_12899,N_6231,N_8632);
nor U12900 (N_12900,N_6679,N_7902);
and U12901 (N_12901,N_9650,N_8564);
or U12902 (N_12902,N_9899,N_8770);
nor U12903 (N_12903,N_7670,N_6289);
or U12904 (N_12904,N_6930,N_5601);
nor U12905 (N_12905,N_5624,N_5880);
nor U12906 (N_12906,N_6119,N_5591);
nand U12907 (N_12907,N_7512,N_5321);
or U12908 (N_12908,N_9481,N_6104);
nor U12909 (N_12909,N_7590,N_5317);
nor U12910 (N_12910,N_7758,N_9653);
nand U12911 (N_12911,N_9186,N_7172);
or U12912 (N_12912,N_6016,N_5205);
or U12913 (N_12913,N_8570,N_8616);
or U12914 (N_12914,N_9346,N_6362);
nand U12915 (N_12915,N_6091,N_5105);
xor U12916 (N_12916,N_6984,N_9824);
nand U12917 (N_12917,N_6260,N_7783);
xor U12918 (N_12918,N_5267,N_6182);
nand U12919 (N_12919,N_5070,N_7860);
and U12920 (N_12920,N_5575,N_6100);
nor U12921 (N_12921,N_5764,N_5683);
and U12922 (N_12922,N_5599,N_8057);
nor U12923 (N_12923,N_7104,N_6543);
or U12924 (N_12924,N_8218,N_6008);
nand U12925 (N_12925,N_7367,N_5358);
nor U12926 (N_12926,N_6817,N_5093);
or U12927 (N_12927,N_6360,N_5278);
and U12928 (N_12928,N_5160,N_5532);
or U12929 (N_12929,N_5142,N_8840);
or U12930 (N_12930,N_9340,N_8086);
nor U12931 (N_12931,N_9355,N_8362);
nor U12932 (N_12932,N_9839,N_5095);
nor U12933 (N_12933,N_5200,N_9944);
nand U12934 (N_12934,N_9014,N_8177);
and U12935 (N_12935,N_9405,N_6905);
and U12936 (N_12936,N_9145,N_6311);
nor U12937 (N_12937,N_8233,N_7906);
or U12938 (N_12938,N_7388,N_9950);
nand U12939 (N_12939,N_8972,N_7838);
and U12940 (N_12940,N_7640,N_6945);
xnor U12941 (N_12941,N_8608,N_9428);
nand U12942 (N_12942,N_9125,N_5635);
and U12943 (N_12943,N_5556,N_6104);
nand U12944 (N_12944,N_6533,N_8961);
or U12945 (N_12945,N_8090,N_8137);
nor U12946 (N_12946,N_7081,N_8991);
and U12947 (N_12947,N_7416,N_9853);
and U12948 (N_12948,N_8927,N_7190);
or U12949 (N_12949,N_7929,N_9670);
xnor U12950 (N_12950,N_6961,N_5128);
nand U12951 (N_12951,N_5209,N_6278);
and U12952 (N_12952,N_9423,N_5620);
or U12953 (N_12953,N_8231,N_8488);
nand U12954 (N_12954,N_9667,N_8665);
or U12955 (N_12955,N_6754,N_7748);
or U12956 (N_12956,N_8381,N_9551);
nand U12957 (N_12957,N_7859,N_9481);
or U12958 (N_12958,N_6180,N_8006);
or U12959 (N_12959,N_5442,N_6903);
nand U12960 (N_12960,N_6604,N_6943);
or U12961 (N_12961,N_9895,N_5696);
nor U12962 (N_12962,N_9196,N_7537);
nor U12963 (N_12963,N_7386,N_5049);
and U12964 (N_12964,N_9302,N_9378);
nand U12965 (N_12965,N_7022,N_6452);
xor U12966 (N_12966,N_6214,N_6016);
or U12967 (N_12967,N_8317,N_5828);
and U12968 (N_12968,N_7050,N_6878);
nor U12969 (N_12969,N_7133,N_9541);
nand U12970 (N_12970,N_8328,N_7482);
xnor U12971 (N_12971,N_6831,N_5777);
nor U12972 (N_12972,N_8280,N_9700);
xnor U12973 (N_12973,N_5153,N_8564);
nand U12974 (N_12974,N_5220,N_8824);
and U12975 (N_12975,N_5996,N_7546);
nand U12976 (N_12976,N_6568,N_8914);
nor U12977 (N_12977,N_8820,N_7555);
xor U12978 (N_12978,N_6750,N_7932);
nor U12979 (N_12979,N_7753,N_8148);
or U12980 (N_12980,N_6255,N_9915);
xnor U12981 (N_12981,N_7173,N_9238);
nand U12982 (N_12982,N_8423,N_6157);
nor U12983 (N_12983,N_7087,N_8212);
or U12984 (N_12984,N_9912,N_8880);
or U12985 (N_12985,N_6597,N_9814);
and U12986 (N_12986,N_7738,N_6474);
xor U12987 (N_12987,N_5732,N_7415);
or U12988 (N_12988,N_5088,N_9207);
xnor U12989 (N_12989,N_6244,N_7984);
nand U12990 (N_12990,N_8321,N_5905);
nor U12991 (N_12991,N_5064,N_7268);
or U12992 (N_12992,N_5328,N_5299);
nor U12993 (N_12993,N_5201,N_5564);
and U12994 (N_12994,N_6890,N_7277);
and U12995 (N_12995,N_5955,N_7549);
xor U12996 (N_12996,N_6952,N_7228);
nor U12997 (N_12997,N_9751,N_7254);
nand U12998 (N_12998,N_6323,N_8887);
or U12999 (N_12999,N_5228,N_7526);
or U13000 (N_13000,N_7870,N_6891);
nor U13001 (N_13001,N_5752,N_9646);
and U13002 (N_13002,N_5327,N_6980);
xnor U13003 (N_13003,N_9277,N_9409);
and U13004 (N_13004,N_6363,N_5484);
nor U13005 (N_13005,N_5099,N_9552);
nor U13006 (N_13006,N_5088,N_5738);
or U13007 (N_13007,N_5039,N_8555);
or U13008 (N_13008,N_7969,N_5912);
xor U13009 (N_13009,N_8523,N_5497);
or U13010 (N_13010,N_9633,N_7089);
or U13011 (N_13011,N_7426,N_8408);
xnor U13012 (N_13012,N_8328,N_5513);
nand U13013 (N_13013,N_6118,N_5681);
nand U13014 (N_13014,N_7570,N_7162);
or U13015 (N_13015,N_7908,N_9725);
and U13016 (N_13016,N_9648,N_8853);
nand U13017 (N_13017,N_7790,N_8148);
or U13018 (N_13018,N_7939,N_9190);
and U13019 (N_13019,N_6864,N_9106);
and U13020 (N_13020,N_9766,N_5079);
nor U13021 (N_13021,N_5325,N_8114);
and U13022 (N_13022,N_8669,N_9808);
xnor U13023 (N_13023,N_7724,N_6703);
nor U13024 (N_13024,N_8473,N_6955);
and U13025 (N_13025,N_5184,N_5041);
nor U13026 (N_13026,N_6013,N_9302);
or U13027 (N_13027,N_6657,N_6001);
and U13028 (N_13028,N_7486,N_5385);
nor U13029 (N_13029,N_9685,N_6884);
nor U13030 (N_13030,N_6991,N_5806);
or U13031 (N_13031,N_9908,N_8293);
and U13032 (N_13032,N_6888,N_5829);
or U13033 (N_13033,N_7144,N_7387);
or U13034 (N_13034,N_8081,N_7003);
nand U13035 (N_13035,N_5843,N_7525);
and U13036 (N_13036,N_5349,N_8186);
nand U13037 (N_13037,N_9934,N_5116);
or U13038 (N_13038,N_9791,N_8827);
and U13039 (N_13039,N_6643,N_8365);
nor U13040 (N_13040,N_8150,N_9206);
nand U13041 (N_13041,N_7635,N_8674);
or U13042 (N_13042,N_6499,N_5447);
nor U13043 (N_13043,N_8366,N_6700);
nand U13044 (N_13044,N_9362,N_9496);
or U13045 (N_13045,N_5896,N_6274);
and U13046 (N_13046,N_7749,N_7027);
nand U13047 (N_13047,N_8808,N_6088);
nand U13048 (N_13048,N_8738,N_9038);
nor U13049 (N_13049,N_5326,N_6763);
and U13050 (N_13050,N_8620,N_9265);
nor U13051 (N_13051,N_9696,N_5100);
xor U13052 (N_13052,N_9184,N_9867);
nor U13053 (N_13053,N_7777,N_9228);
nand U13054 (N_13054,N_8113,N_8413);
nand U13055 (N_13055,N_8471,N_5220);
xor U13056 (N_13056,N_6571,N_7597);
nor U13057 (N_13057,N_5084,N_5547);
nor U13058 (N_13058,N_6097,N_6224);
nor U13059 (N_13059,N_8066,N_9747);
and U13060 (N_13060,N_9437,N_7401);
and U13061 (N_13061,N_8176,N_7879);
or U13062 (N_13062,N_7111,N_5441);
nor U13063 (N_13063,N_8090,N_7302);
xnor U13064 (N_13064,N_7195,N_6243);
nor U13065 (N_13065,N_7952,N_9497);
nand U13066 (N_13066,N_8207,N_6720);
nor U13067 (N_13067,N_7008,N_5839);
and U13068 (N_13068,N_7915,N_9570);
nor U13069 (N_13069,N_9217,N_6236);
or U13070 (N_13070,N_7535,N_6223);
or U13071 (N_13071,N_5128,N_5186);
nor U13072 (N_13072,N_7276,N_7345);
or U13073 (N_13073,N_6146,N_8387);
nor U13074 (N_13074,N_5692,N_7679);
or U13075 (N_13075,N_8847,N_6460);
xor U13076 (N_13076,N_9529,N_6268);
nand U13077 (N_13077,N_9342,N_6613);
or U13078 (N_13078,N_7926,N_5653);
or U13079 (N_13079,N_9997,N_8403);
and U13080 (N_13080,N_6856,N_5983);
nand U13081 (N_13081,N_8533,N_5837);
or U13082 (N_13082,N_7169,N_9568);
and U13083 (N_13083,N_5857,N_6906);
and U13084 (N_13084,N_9984,N_8795);
nor U13085 (N_13085,N_9719,N_5618);
nor U13086 (N_13086,N_7380,N_5324);
nor U13087 (N_13087,N_5040,N_9793);
nand U13088 (N_13088,N_7973,N_5905);
nor U13089 (N_13089,N_8160,N_9928);
or U13090 (N_13090,N_7835,N_6398);
and U13091 (N_13091,N_9746,N_8628);
nor U13092 (N_13092,N_9160,N_8382);
or U13093 (N_13093,N_6844,N_6403);
or U13094 (N_13094,N_5670,N_9819);
nand U13095 (N_13095,N_7419,N_5094);
xnor U13096 (N_13096,N_7293,N_7387);
nand U13097 (N_13097,N_7152,N_7244);
or U13098 (N_13098,N_9676,N_5782);
nor U13099 (N_13099,N_5874,N_5429);
nor U13100 (N_13100,N_8061,N_7104);
xor U13101 (N_13101,N_9292,N_9578);
nor U13102 (N_13102,N_5051,N_5201);
and U13103 (N_13103,N_8533,N_8063);
or U13104 (N_13104,N_5103,N_5993);
nand U13105 (N_13105,N_5026,N_9935);
and U13106 (N_13106,N_5774,N_7024);
nor U13107 (N_13107,N_6338,N_6506);
or U13108 (N_13108,N_6549,N_8076);
nor U13109 (N_13109,N_6685,N_6333);
xor U13110 (N_13110,N_6354,N_5552);
nand U13111 (N_13111,N_7443,N_8191);
nor U13112 (N_13112,N_8208,N_9380);
and U13113 (N_13113,N_6463,N_8243);
and U13114 (N_13114,N_8714,N_6409);
and U13115 (N_13115,N_9489,N_6185);
nor U13116 (N_13116,N_7412,N_7409);
and U13117 (N_13117,N_6326,N_8985);
and U13118 (N_13118,N_6546,N_7597);
or U13119 (N_13119,N_5835,N_5271);
nor U13120 (N_13120,N_7008,N_6670);
or U13121 (N_13121,N_6732,N_6324);
and U13122 (N_13122,N_6786,N_5134);
nor U13123 (N_13123,N_5719,N_5575);
or U13124 (N_13124,N_5802,N_7956);
nand U13125 (N_13125,N_8304,N_5988);
or U13126 (N_13126,N_8726,N_8647);
nor U13127 (N_13127,N_7335,N_9328);
nand U13128 (N_13128,N_9839,N_6962);
and U13129 (N_13129,N_5451,N_7488);
or U13130 (N_13130,N_9473,N_6742);
or U13131 (N_13131,N_7056,N_9353);
or U13132 (N_13132,N_9908,N_5804);
xnor U13133 (N_13133,N_6714,N_5086);
or U13134 (N_13134,N_7007,N_8512);
nor U13135 (N_13135,N_8511,N_7497);
and U13136 (N_13136,N_5558,N_6236);
nand U13137 (N_13137,N_7073,N_7014);
nor U13138 (N_13138,N_6995,N_8415);
nor U13139 (N_13139,N_5136,N_7537);
nand U13140 (N_13140,N_6043,N_7131);
or U13141 (N_13141,N_8372,N_5564);
nor U13142 (N_13142,N_8991,N_5203);
nor U13143 (N_13143,N_8145,N_5590);
xnor U13144 (N_13144,N_5709,N_9959);
and U13145 (N_13145,N_5927,N_9338);
or U13146 (N_13146,N_8606,N_8820);
or U13147 (N_13147,N_6777,N_7978);
or U13148 (N_13148,N_9689,N_9966);
nor U13149 (N_13149,N_6338,N_5735);
nor U13150 (N_13150,N_5356,N_7581);
and U13151 (N_13151,N_9459,N_9658);
and U13152 (N_13152,N_9795,N_8587);
nor U13153 (N_13153,N_8349,N_5342);
nor U13154 (N_13154,N_7878,N_8662);
xnor U13155 (N_13155,N_6251,N_6547);
xnor U13156 (N_13156,N_6840,N_8150);
nor U13157 (N_13157,N_5013,N_9772);
nor U13158 (N_13158,N_7255,N_6408);
and U13159 (N_13159,N_7163,N_7166);
and U13160 (N_13160,N_9615,N_5878);
nor U13161 (N_13161,N_5319,N_5874);
xor U13162 (N_13162,N_6734,N_8769);
xor U13163 (N_13163,N_5343,N_9047);
and U13164 (N_13164,N_6841,N_6139);
nand U13165 (N_13165,N_5028,N_5395);
nand U13166 (N_13166,N_8320,N_7276);
and U13167 (N_13167,N_7545,N_5470);
and U13168 (N_13168,N_8096,N_8170);
xor U13169 (N_13169,N_8543,N_6389);
nand U13170 (N_13170,N_6973,N_7594);
nand U13171 (N_13171,N_6292,N_7757);
and U13172 (N_13172,N_7002,N_7293);
xor U13173 (N_13173,N_9712,N_5791);
and U13174 (N_13174,N_8304,N_8288);
nand U13175 (N_13175,N_6426,N_7442);
and U13176 (N_13176,N_6702,N_6641);
nand U13177 (N_13177,N_5165,N_8885);
nand U13178 (N_13178,N_5636,N_7909);
or U13179 (N_13179,N_6316,N_5428);
nand U13180 (N_13180,N_9060,N_8104);
and U13181 (N_13181,N_6831,N_9651);
and U13182 (N_13182,N_8986,N_8579);
nand U13183 (N_13183,N_5850,N_6400);
and U13184 (N_13184,N_6493,N_6987);
or U13185 (N_13185,N_5630,N_5938);
nand U13186 (N_13186,N_9371,N_5567);
or U13187 (N_13187,N_6826,N_5764);
nand U13188 (N_13188,N_6857,N_7937);
or U13189 (N_13189,N_9350,N_5626);
nor U13190 (N_13190,N_8908,N_8007);
xnor U13191 (N_13191,N_8534,N_7791);
and U13192 (N_13192,N_7501,N_6733);
nand U13193 (N_13193,N_6029,N_8620);
or U13194 (N_13194,N_9563,N_5955);
or U13195 (N_13195,N_7318,N_9566);
or U13196 (N_13196,N_7443,N_5930);
nand U13197 (N_13197,N_7888,N_5378);
xor U13198 (N_13198,N_8125,N_6177);
nor U13199 (N_13199,N_6831,N_8594);
or U13200 (N_13200,N_8648,N_6182);
nand U13201 (N_13201,N_5913,N_9880);
nor U13202 (N_13202,N_7286,N_5229);
and U13203 (N_13203,N_5277,N_6056);
and U13204 (N_13204,N_7621,N_5018);
nand U13205 (N_13205,N_9523,N_5330);
nor U13206 (N_13206,N_5043,N_5963);
and U13207 (N_13207,N_7844,N_8880);
and U13208 (N_13208,N_9257,N_8290);
and U13209 (N_13209,N_6335,N_6643);
or U13210 (N_13210,N_7540,N_5990);
nor U13211 (N_13211,N_8867,N_6913);
nor U13212 (N_13212,N_5896,N_6987);
nand U13213 (N_13213,N_8283,N_9840);
nand U13214 (N_13214,N_7852,N_9294);
nand U13215 (N_13215,N_6860,N_5970);
and U13216 (N_13216,N_6225,N_5248);
nand U13217 (N_13217,N_8401,N_9409);
nor U13218 (N_13218,N_7186,N_9255);
or U13219 (N_13219,N_5931,N_8141);
nand U13220 (N_13220,N_6977,N_5499);
nor U13221 (N_13221,N_7730,N_7791);
nor U13222 (N_13222,N_7180,N_7205);
or U13223 (N_13223,N_5879,N_6902);
nand U13224 (N_13224,N_6872,N_5463);
or U13225 (N_13225,N_9626,N_7470);
or U13226 (N_13226,N_8880,N_6427);
nand U13227 (N_13227,N_7488,N_8808);
nand U13228 (N_13228,N_5161,N_6465);
and U13229 (N_13229,N_7770,N_5700);
and U13230 (N_13230,N_8110,N_7973);
or U13231 (N_13231,N_8084,N_7279);
nor U13232 (N_13232,N_6379,N_9510);
nand U13233 (N_13233,N_9875,N_8766);
or U13234 (N_13234,N_9919,N_9464);
or U13235 (N_13235,N_8591,N_8367);
nor U13236 (N_13236,N_9361,N_9443);
nor U13237 (N_13237,N_8804,N_6995);
nor U13238 (N_13238,N_9940,N_5018);
nand U13239 (N_13239,N_6918,N_6374);
and U13240 (N_13240,N_5456,N_7289);
nand U13241 (N_13241,N_8733,N_5843);
or U13242 (N_13242,N_7316,N_5385);
nor U13243 (N_13243,N_7069,N_6046);
or U13244 (N_13244,N_6329,N_6726);
nor U13245 (N_13245,N_5803,N_6072);
nand U13246 (N_13246,N_8835,N_5627);
and U13247 (N_13247,N_5663,N_8981);
nand U13248 (N_13248,N_5446,N_8632);
xnor U13249 (N_13249,N_5220,N_9317);
and U13250 (N_13250,N_9498,N_6497);
or U13251 (N_13251,N_6130,N_7142);
and U13252 (N_13252,N_5134,N_9507);
and U13253 (N_13253,N_8146,N_7848);
nor U13254 (N_13254,N_5370,N_6143);
or U13255 (N_13255,N_8757,N_6104);
xor U13256 (N_13256,N_8670,N_6444);
or U13257 (N_13257,N_9794,N_9576);
and U13258 (N_13258,N_6531,N_7899);
nand U13259 (N_13259,N_5503,N_6824);
nand U13260 (N_13260,N_5858,N_5852);
and U13261 (N_13261,N_7531,N_6461);
and U13262 (N_13262,N_9922,N_8570);
xnor U13263 (N_13263,N_9814,N_7312);
or U13264 (N_13264,N_8405,N_9350);
and U13265 (N_13265,N_9936,N_5357);
nor U13266 (N_13266,N_6410,N_6570);
and U13267 (N_13267,N_5696,N_6065);
nor U13268 (N_13268,N_6554,N_5524);
and U13269 (N_13269,N_6721,N_5719);
nor U13270 (N_13270,N_6401,N_6976);
and U13271 (N_13271,N_8826,N_9186);
and U13272 (N_13272,N_5854,N_7327);
or U13273 (N_13273,N_6991,N_6080);
or U13274 (N_13274,N_6825,N_7877);
or U13275 (N_13275,N_7741,N_7174);
xnor U13276 (N_13276,N_7219,N_9007);
or U13277 (N_13277,N_5600,N_8274);
xor U13278 (N_13278,N_5887,N_7287);
nand U13279 (N_13279,N_5477,N_7657);
nor U13280 (N_13280,N_5039,N_8587);
or U13281 (N_13281,N_7051,N_9685);
or U13282 (N_13282,N_6616,N_6998);
and U13283 (N_13283,N_5062,N_9903);
nand U13284 (N_13284,N_5356,N_9900);
nor U13285 (N_13285,N_7842,N_9667);
nand U13286 (N_13286,N_8312,N_9910);
and U13287 (N_13287,N_6628,N_7322);
and U13288 (N_13288,N_9784,N_7412);
nand U13289 (N_13289,N_9395,N_9729);
and U13290 (N_13290,N_8514,N_7276);
nor U13291 (N_13291,N_9137,N_8430);
or U13292 (N_13292,N_9374,N_5338);
or U13293 (N_13293,N_5967,N_8562);
or U13294 (N_13294,N_9365,N_9204);
and U13295 (N_13295,N_8777,N_7263);
nor U13296 (N_13296,N_8206,N_5422);
xnor U13297 (N_13297,N_5035,N_9412);
nor U13298 (N_13298,N_8913,N_5633);
xor U13299 (N_13299,N_9767,N_8405);
or U13300 (N_13300,N_5583,N_9003);
nor U13301 (N_13301,N_9889,N_8250);
or U13302 (N_13302,N_7587,N_8762);
nor U13303 (N_13303,N_6473,N_8017);
and U13304 (N_13304,N_6999,N_5058);
or U13305 (N_13305,N_7081,N_5548);
nor U13306 (N_13306,N_5845,N_9505);
nand U13307 (N_13307,N_9038,N_9664);
or U13308 (N_13308,N_7904,N_9582);
or U13309 (N_13309,N_5071,N_7714);
nor U13310 (N_13310,N_5803,N_5110);
and U13311 (N_13311,N_7111,N_6692);
nand U13312 (N_13312,N_8073,N_6421);
nor U13313 (N_13313,N_8983,N_9510);
or U13314 (N_13314,N_5383,N_8444);
xor U13315 (N_13315,N_7879,N_9950);
nor U13316 (N_13316,N_7351,N_5541);
nor U13317 (N_13317,N_6467,N_9782);
or U13318 (N_13318,N_6489,N_5782);
or U13319 (N_13319,N_6791,N_7436);
nor U13320 (N_13320,N_9663,N_7775);
or U13321 (N_13321,N_5952,N_5148);
nor U13322 (N_13322,N_7286,N_9052);
or U13323 (N_13323,N_5643,N_8089);
and U13324 (N_13324,N_7388,N_6203);
nand U13325 (N_13325,N_8767,N_5054);
and U13326 (N_13326,N_5761,N_9879);
nand U13327 (N_13327,N_6227,N_6790);
xor U13328 (N_13328,N_6199,N_7594);
or U13329 (N_13329,N_8163,N_8518);
nor U13330 (N_13330,N_8421,N_7070);
nand U13331 (N_13331,N_8324,N_6062);
xnor U13332 (N_13332,N_9074,N_5557);
nor U13333 (N_13333,N_8643,N_5023);
nor U13334 (N_13334,N_9592,N_5714);
nand U13335 (N_13335,N_5021,N_7803);
nand U13336 (N_13336,N_9588,N_8406);
or U13337 (N_13337,N_5012,N_8405);
nand U13338 (N_13338,N_8160,N_6438);
nand U13339 (N_13339,N_5188,N_7983);
nor U13340 (N_13340,N_8552,N_9424);
nand U13341 (N_13341,N_5116,N_5835);
xnor U13342 (N_13342,N_6348,N_9799);
nand U13343 (N_13343,N_8882,N_6455);
nor U13344 (N_13344,N_5698,N_5014);
or U13345 (N_13345,N_7822,N_8073);
or U13346 (N_13346,N_6756,N_5874);
nand U13347 (N_13347,N_8415,N_6518);
xnor U13348 (N_13348,N_6631,N_6326);
nand U13349 (N_13349,N_8160,N_6970);
nand U13350 (N_13350,N_6125,N_5997);
or U13351 (N_13351,N_5086,N_7018);
nor U13352 (N_13352,N_8236,N_6872);
or U13353 (N_13353,N_9087,N_5528);
or U13354 (N_13354,N_8413,N_7393);
nand U13355 (N_13355,N_6709,N_5918);
or U13356 (N_13356,N_6847,N_9226);
nand U13357 (N_13357,N_7211,N_6491);
nand U13358 (N_13358,N_5529,N_5875);
nand U13359 (N_13359,N_8146,N_5567);
or U13360 (N_13360,N_5576,N_8757);
xor U13361 (N_13361,N_5985,N_9788);
or U13362 (N_13362,N_6711,N_7391);
nor U13363 (N_13363,N_5001,N_7919);
or U13364 (N_13364,N_6033,N_8821);
and U13365 (N_13365,N_6803,N_6281);
nand U13366 (N_13366,N_7808,N_6125);
or U13367 (N_13367,N_9398,N_8197);
or U13368 (N_13368,N_8204,N_5272);
xor U13369 (N_13369,N_6068,N_6786);
xnor U13370 (N_13370,N_9615,N_6741);
and U13371 (N_13371,N_9757,N_8514);
nor U13372 (N_13372,N_6195,N_6626);
or U13373 (N_13373,N_9527,N_7439);
or U13374 (N_13374,N_5879,N_5956);
or U13375 (N_13375,N_5753,N_7596);
or U13376 (N_13376,N_5331,N_9374);
or U13377 (N_13377,N_6480,N_5340);
and U13378 (N_13378,N_7275,N_6406);
or U13379 (N_13379,N_7915,N_5524);
nor U13380 (N_13380,N_8970,N_5056);
and U13381 (N_13381,N_5438,N_6168);
nor U13382 (N_13382,N_8873,N_6819);
nand U13383 (N_13383,N_7030,N_7740);
or U13384 (N_13384,N_6906,N_6088);
nand U13385 (N_13385,N_8043,N_9893);
and U13386 (N_13386,N_8625,N_7509);
xnor U13387 (N_13387,N_6734,N_9365);
nor U13388 (N_13388,N_9391,N_6574);
or U13389 (N_13389,N_8449,N_5967);
nor U13390 (N_13390,N_8774,N_7068);
nand U13391 (N_13391,N_7722,N_9071);
nand U13392 (N_13392,N_9673,N_7237);
or U13393 (N_13393,N_7402,N_5423);
or U13394 (N_13394,N_7359,N_7779);
xor U13395 (N_13395,N_5136,N_5579);
nand U13396 (N_13396,N_8506,N_9940);
nor U13397 (N_13397,N_6455,N_5109);
and U13398 (N_13398,N_6635,N_7406);
and U13399 (N_13399,N_8149,N_9061);
nor U13400 (N_13400,N_7510,N_6562);
xnor U13401 (N_13401,N_7589,N_8972);
and U13402 (N_13402,N_6204,N_9627);
and U13403 (N_13403,N_7158,N_6033);
or U13404 (N_13404,N_8013,N_9636);
or U13405 (N_13405,N_7053,N_7034);
xor U13406 (N_13406,N_9281,N_8923);
or U13407 (N_13407,N_6739,N_8552);
or U13408 (N_13408,N_7853,N_9292);
nor U13409 (N_13409,N_8874,N_8665);
nand U13410 (N_13410,N_6587,N_6688);
nand U13411 (N_13411,N_9451,N_7928);
nor U13412 (N_13412,N_8442,N_9692);
nor U13413 (N_13413,N_9486,N_6124);
or U13414 (N_13414,N_8142,N_8599);
nor U13415 (N_13415,N_8396,N_9122);
or U13416 (N_13416,N_6538,N_8775);
nor U13417 (N_13417,N_8618,N_9614);
nand U13418 (N_13418,N_6203,N_9938);
and U13419 (N_13419,N_6559,N_8854);
or U13420 (N_13420,N_7257,N_5900);
or U13421 (N_13421,N_7255,N_7378);
and U13422 (N_13422,N_9157,N_5259);
nand U13423 (N_13423,N_8924,N_9657);
and U13424 (N_13424,N_6303,N_6897);
or U13425 (N_13425,N_6251,N_6066);
nor U13426 (N_13426,N_9412,N_7028);
and U13427 (N_13427,N_9277,N_9912);
and U13428 (N_13428,N_6021,N_7315);
and U13429 (N_13429,N_6367,N_9235);
nor U13430 (N_13430,N_8894,N_8585);
or U13431 (N_13431,N_8752,N_6540);
nor U13432 (N_13432,N_7551,N_5054);
and U13433 (N_13433,N_7203,N_5891);
nor U13434 (N_13434,N_8277,N_8246);
or U13435 (N_13435,N_7385,N_8673);
and U13436 (N_13436,N_5609,N_5962);
nand U13437 (N_13437,N_8377,N_9087);
nor U13438 (N_13438,N_9803,N_5661);
nand U13439 (N_13439,N_8332,N_6759);
or U13440 (N_13440,N_6816,N_8164);
nor U13441 (N_13441,N_7730,N_9128);
or U13442 (N_13442,N_6494,N_8571);
or U13443 (N_13443,N_5428,N_6659);
nand U13444 (N_13444,N_8486,N_9996);
nor U13445 (N_13445,N_6100,N_5571);
xor U13446 (N_13446,N_6196,N_7317);
nand U13447 (N_13447,N_9831,N_8173);
and U13448 (N_13448,N_6744,N_9206);
xnor U13449 (N_13449,N_6220,N_8068);
nor U13450 (N_13450,N_5236,N_8479);
or U13451 (N_13451,N_8055,N_7689);
xnor U13452 (N_13452,N_8434,N_9911);
nor U13453 (N_13453,N_8798,N_5549);
nand U13454 (N_13454,N_6717,N_9427);
or U13455 (N_13455,N_9809,N_9251);
or U13456 (N_13456,N_6257,N_6938);
xnor U13457 (N_13457,N_8849,N_8092);
nand U13458 (N_13458,N_5795,N_5895);
or U13459 (N_13459,N_7360,N_5943);
or U13460 (N_13460,N_6922,N_7378);
nand U13461 (N_13461,N_7158,N_9478);
nand U13462 (N_13462,N_8051,N_5452);
nor U13463 (N_13463,N_6298,N_7046);
nor U13464 (N_13464,N_9246,N_6561);
nor U13465 (N_13465,N_7299,N_9297);
nor U13466 (N_13466,N_7103,N_8292);
nand U13467 (N_13467,N_9605,N_7383);
or U13468 (N_13468,N_6327,N_5844);
and U13469 (N_13469,N_8232,N_5030);
nor U13470 (N_13470,N_9993,N_7074);
and U13471 (N_13471,N_5816,N_5564);
and U13472 (N_13472,N_8948,N_5944);
nor U13473 (N_13473,N_6267,N_6763);
nand U13474 (N_13474,N_9376,N_5268);
or U13475 (N_13475,N_7121,N_7325);
or U13476 (N_13476,N_6650,N_7384);
nor U13477 (N_13477,N_9345,N_5062);
and U13478 (N_13478,N_9198,N_6340);
nor U13479 (N_13479,N_9402,N_6172);
nand U13480 (N_13480,N_9206,N_7667);
or U13481 (N_13481,N_9781,N_6722);
nor U13482 (N_13482,N_8999,N_7934);
nor U13483 (N_13483,N_5487,N_8899);
nor U13484 (N_13484,N_7591,N_9504);
and U13485 (N_13485,N_9253,N_5266);
or U13486 (N_13486,N_7611,N_9915);
nor U13487 (N_13487,N_6407,N_9339);
xnor U13488 (N_13488,N_9777,N_9077);
or U13489 (N_13489,N_5111,N_6483);
and U13490 (N_13490,N_6801,N_9701);
nand U13491 (N_13491,N_6627,N_7302);
and U13492 (N_13492,N_6739,N_5824);
or U13493 (N_13493,N_5041,N_9651);
nand U13494 (N_13494,N_6738,N_8320);
nor U13495 (N_13495,N_9894,N_7206);
xor U13496 (N_13496,N_9746,N_7145);
nor U13497 (N_13497,N_7580,N_5607);
and U13498 (N_13498,N_9378,N_9707);
and U13499 (N_13499,N_8917,N_9517);
and U13500 (N_13500,N_8902,N_7398);
nor U13501 (N_13501,N_7414,N_8825);
nor U13502 (N_13502,N_8335,N_5675);
xnor U13503 (N_13503,N_7512,N_5771);
and U13504 (N_13504,N_9021,N_8717);
nand U13505 (N_13505,N_6360,N_9952);
and U13506 (N_13506,N_7394,N_5674);
and U13507 (N_13507,N_7620,N_5994);
nor U13508 (N_13508,N_7361,N_6975);
nand U13509 (N_13509,N_7031,N_9123);
or U13510 (N_13510,N_8790,N_7839);
xnor U13511 (N_13511,N_9804,N_5267);
nor U13512 (N_13512,N_5641,N_5526);
and U13513 (N_13513,N_9355,N_5210);
nand U13514 (N_13514,N_6552,N_9181);
xnor U13515 (N_13515,N_5877,N_5714);
nand U13516 (N_13516,N_9518,N_6905);
and U13517 (N_13517,N_9402,N_6240);
and U13518 (N_13518,N_6195,N_7008);
or U13519 (N_13519,N_8645,N_8887);
and U13520 (N_13520,N_7762,N_5620);
or U13521 (N_13521,N_7465,N_5578);
or U13522 (N_13522,N_7970,N_8658);
and U13523 (N_13523,N_9020,N_6673);
nor U13524 (N_13524,N_8750,N_9650);
nor U13525 (N_13525,N_9908,N_6857);
or U13526 (N_13526,N_8192,N_7648);
and U13527 (N_13527,N_5709,N_7803);
xnor U13528 (N_13528,N_5753,N_5779);
nand U13529 (N_13529,N_9490,N_9046);
and U13530 (N_13530,N_9267,N_9790);
nor U13531 (N_13531,N_6369,N_6044);
and U13532 (N_13532,N_6946,N_6055);
and U13533 (N_13533,N_5949,N_9961);
xor U13534 (N_13534,N_6358,N_7489);
or U13535 (N_13535,N_8235,N_9338);
or U13536 (N_13536,N_5956,N_7332);
or U13537 (N_13537,N_9671,N_5758);
and U13538 (N_13538,N_8201,N_5882);
nor U13539 (N_13539,N_5075,N_7933);
or U13540 (N_13540,N_8495,N_9923);
and U13541 (N_13541,N_6389,N_5936);
or U13542 (N_13542,N_6311,N_8964);
xor U13543 (N_13543,N_7246,N_7221);
nor U13544 (N_13544,N_7591,N_9187);
nor U13545 (N_13545,N_9850,N_6821);
or U13546 (N_13546,N_9086,N_7980);
and U13547 (N_13547,N_7964,N_6725);
nand U13548 (N_13548,N_5511,N_8430);
or U13549 (N_13549,N_6135,N_5650);
xnor U13550 (N_13550,N_7568,N_7942);
and U13551 (N_13551,N_9261,N_7031);
nand U13552 (N_13552,N_6505,N_7074);
or U13553 (N_13553,N_6988,N_9928);
xnor U13554 (N_13554,N_5708,N_9115);
nor U13555 (N_13555,N_7301,N_7369);
nor U13556 (N_13556,N_6589,N_6521);
nor U13557 (N_13557,N_6415,N_7797);
or U13558 (N_13558,N_9673,N_9186);
nor U13559 (N_13559,N_8117,N_6859);
nor U13560 (N_13560,N_7481,N_9721);
or U13561 (N_13561,N_9538,N_5803);
nor U13562 (N_13562,N_6272,N_5451);
nand U13563 (N_13563,N_5697,N_7876);
and U13564 (N_13564,N_6266,N_8304);
nand U13565 (N_13565,N_8469,N_7467);
nor U13566 (N_13566,N_9036,N_7068);
nor U13567 (N_13567,N_5634,N_7951);
and U13568 (N_13568,N_7472,N_8710);
and U13569 (N_13569,N_9460,N_7601);
and U13570 (N_13570,N_6698,N_7698);
xor U13571 (N_13571,N_9805,N_5559);
xnor U13572 (N_13572,N_6635,N_8309);
and U13573 (N_13573,N_6023,N_5959);
or U13574 (N_13574,N_9977,N_8171);
nor U13575 (N_13575,N_9575,N_7788);
xor U13576 (N_13576,N_6127,N_5827);
nand U13577 (N_13577,N_6644,N_5047);
nand U13578 (N_13578,N_6897,N_6667);
nand U13579 (N_13579,N_9783,N_7596);
and U13580 (N_13580,N_5688,N_7160);
and U13581 (N_13581,N_7556,N_7535);
xor U13582 (N_13582,N_9098,N_5782);
nand U13583 (N_13583,N_9132,N_8472);
nand U13584 (N_13584,N_6717,N_8411);
nand U13585 (N_13585,N_7592,N_5125);
nor U13586 (N_13586,N_5993,N_7546);
and U13587 (N_13587,N_5091,N_5785);
nand U13588 (N_13588,N_5344,N_7639);
nand U13589 (N_13589,N_7064,N_7305);
or U13590 (N_13590,N_6978,N_5505);
and U13591 (N_13591,N_6271,N_5712);
nand U13592 (N_13592,N_7979,N_5591);
or U13593 (N_13593,N_5694,N_9554);
and U13594 (N_13594,N_8371,N_5552);
nor U13595 (N_13595,N_8406,N_9476);
or U13596 (N_13596,N_8597,N_6888);
or U13597 (N_13597,N_8056,N_5698);
nand U13598 (N_13598,N_7087,N_6812);
or U13599 (N_13599,N_9431,N_8627);
and U13600 (N_13600,N_6316,N_8074);
nand U13601 (N_13601,N_8763,N_5157);
xor U13602 (N_13602,N_5902,N_8872);
or U13603 (N_13603,N_5016,N_7641);
and U13604 (N_13604,N_5593,N_6680);
and U13605 (N_13605,N_5734,N_8699);
or U13606 (N_13606,N_5018,N_8084);
xor U13607 (N_13607,N_5827,N_8860);
and U13608 (N_13608,N_9773,N_9037);
nand U13609 (N_13609,N_7029,N_9316);
nand U13610 (N_13610,N_9459,N_9225);
xor U13611 (N_13611,N_9530,N_8747);
and U13612 (N_13612,N_8535,N_5973);
or U13613 (N_13613,N_6521,N_9985);
or U13614 (N_13614,N_8715,N_8425);
nor U13615 (N_13615,N_6524,N_7135);
nor U13616 (N_13616,N_9993,N_9363);
and U13617 (N_13617,N_7053,N_6249);
xor U13618 (N_13618,N_5472,N_9672);
or U13619 (N_13619,N_7868,N_7835);
nand U13620 (N_13620,N_6275,N_9909);
nand U13621 (N_13621,N_5125,N_8617);
xor U13622 (N_13622,N_8427,N_6542);
nor U13623 (N_13623,N_5051,N_5002);
and U13624 (N_13624,N_5493,N_8922);
nand U13625 (N_13625,N_9656,N_5758);
nand U13626 (N_13626,N_6482,N_8847);
or U13627 (N_13627,N_6057,N_6226);
or U13628 (N_13628,N_7966,N_5301);
and U13629 (N_13629,N_5154,N_5469);
nor U13630 (N_13630,N_5438,N_7064);
or U13631 (N_13631,N_7620,N_6996);
and U13632 (N_13632,N_8051,N_9640);
or U13633 (N_13633,N_8595,N_9435);
xnor U13634 (N_13634,N_9591,N_6952);
and U13635 (N_13635,N_5468,N_6910);
nand U13636 (N_13636,N_5813,N_6931);
nor U13637 (N_13637,N_8345,N_9206);
nand U13638 (N_13638,N_5172,N_6790);
or U13639 (N_13639,N_8023,N_5466);
and U13640 (N_13640,N_5741,N_5848);
nor U13641 (N_13641,N_9039,N_9124);
or U13642 (N_13642,N_8817,N_9639);
or U13643 (N_13643,N_9368,N_6944);
and U13644 (N_13644,N_7579,N_5130);
and U13645 (N_13645,N_5191,N_9386);
and U13646 (N_13646,N_5816,N_6254);
xnor U13647 (N_13647,N_5733,N_6977);
xor U13648 (N_13648,N_8422,N_9981);
xor U13649 (N_13649,N_7028,N_8412);
or U13650 (N_13650,N_8133,N_7545);
nand U13651 (N_13651,N_9327,N_9985);
xor U13652 (N_13652,N_8766,N_9035);
and U13653 (N_13653,N_6358,N_8310);
nor U13654 (N_13654,N_8989,N_5187);
nor U13655 (N_13655,N_9289,N_8317);
and U13656 (N_13656,N_7426,N_9613);
nor U13657 (N_13657,N_9168,N_9062);
and U13658 (N_13658,N_9102,N_9883);
nor U13659 (N_13659,N_7541,N_6129);
nand U13660 (N_13660,N_5836,N_6093);
xor U13661 (N_13661,N_7488,N_7219);
nand U13662 (N_13662,N_6763,N_8618);
or U13663 (N_13663,N_8356,N_9002);
or U13664 (N_13664,N_6557,N_9847);
nor U13665 (N_13665,N_5918,N_9523);
or U13666 (N_13666,N_8172,N_8660);
or U13667 (N_13667,N_5203,N_8695);
nor U13668 (N_13668,N_7015,N_5201);
nor U13669 (N_13669,N_7655,N_6146);
or U13670 (N_13670,N_5676,N_9328);
nand U13671 (N_13671,N_5630,N_9901);
xnor U13672 (N_13672,N_9747,N_8104);
nor U13673 (N_13673,N_8830,N_7427);
and U13674 (N_13674,N_7256,N_5916);
or U13675 (N_13675,N_9031,N_5036);
and U13676 (N_13676,N_9511,N_9525);
nand U13677 (N_13677,N_7928,N_5266);
nand U13678 (N_13678,N_8292,N_9050);
and U13679 (N_13679,N_6876,N_5190);
and U13680 (N_13680,N_9666,N_9751);
nand U13681 (N_13681,N_5489,N_9501);
xnor U13682 (N_13682,N_9102,N_7638);
nand U13683 (N_13683,N_8892,N_6909);
or U13684 (N_13684,N_5581,N_5660);
nor U13685 (N_13685,N_8680,N_8659);
and U13686 (N_13686,N_6297,N_6276);
and U13687 (N_13687,N_7706,N_8370);
nand U13688 (N_13688,N_9633,N_5341);
nand U13689 (N_13689,N_7326,N_7640);
xnor U13690 (N_13690,N_5120,N_7325);
nor U13691 (N_13691,N_6080,N_8974);
nor U13692 (N_13692,N_6554,N_5253);
xnor U13693 (N_13693,N_9391,N_6850);
or U13694 (N_13694,N_7377,N_8812);
or U13695 (N_13695,N_7638,N_8890);
nor U13696 (N_13696,N_8534,N_7015);
and U13697 (N_13697,N_9939,N_7782);
or U13698 (N_13698,N_7182,N_5589);
or U13699 (N_13699,N_7664,N_9591);
nor U13700 (N_13700,N_7750,N_8534);
and U13701 (N_13701,N_8532,N_9623);
or U13702 (N_13702,N_7323,N_8779);
and U13703 (N_13703,N_6437,N_9144);
or U13704 (N_13704,N_8243,N_8208);
and U13705 (N_13705,N_9110,N_5012);
nor U13706 (N_13706,N_8364,N_6961);
and U13707 (N_13707,N_9809,N_6209);
or U13708 (N_13708,N_8875,N_8643);
or U13709 (N_13709,N_6941,N_6532);
nor U13710 (N_13710,N_9169,N_7054);
and U13711 (N_13711,N_9691,N_8839);
or U13712 (N_13712,N_8296,N_9719);
or U13713 (N_13713,N_9869,N_9452);
or U13714 (N_13714,N_5855,N_8926);
or U13715 (N_13715,N_8423,N_5894);
nor U13716 (N_13716,N_7761,N_7139);
and U13717 (N_13717,N_6853,N_5626);
or U13718 (N_13718,N_9352,N_8552);
and U13719 (N_13719,N_9820,N_9932);
nand U13720 (N_13720,N_5234,N_6899);
or U13721 (N_13721,N_8864,N_9672);
nand U13722 (N_13722,N_6589,N_9004);
or U13723 (N_13723,N_6878,N_7573);
nand U13724 (N_13724,N_7589,N_8625);
nor U13725 (N_13725,N_8565,N_6491);
and U13726 (N_13726,N_5192,N_6997);
or U13727 (N_13727,N_8675,N_9070);
nor U13728 (N_13728,N_7989,N_5383);
or U13729 (N_13729,N_5520,N_7564);
or U13730 (N_13730,N_9776,N_5256);
or U13731 (N_13731,N_6956,N_7856);
or U13732 (N_13732,N_5555,N_7716);
and U13733 (N_13733,N_8292,N_9606);
or U13734 (N_13734,N_7999,N_7172);
or U13735 (N_13735,N_5794,N_7523);
nand U13736 (N_13736,N_7244,N_9028);
nor U13737 (N_13737,N_8332,N_7679);
or U13738 (N_13738,N_7894,N_6369);
or U13739 (N_13739,N_9394,N_6501);
or U13740 (N_13740,N_6137,N_7197);
nor U13741 (N_13741,N_6780,N_9704);
xor U13742 (N_13742,N_5276,N_5034);
and U13743 (N_13743,N_6719,N_9432);
nor U13744 (N_13744,N_5057,N_9919);
or U13745 (N_13745,N_8706,N_6895);
nor U13746 (N_13746,N_7669,N_5426);
nor U13747 (N_13747,N_5144,N_8644);
xnor U13748 (N_13748,N_8109,N_9984);
and U13749 (N_13749,N_5939,N_6139);
nand U13750 (N_13750,N_5358,N_7906);
nor U13751 (N_13751,N_5586,N_5256);
xor U13752 (N_13752,N_5524,N_7871);
nor U13753 (N_13753,N_6023,N_5334);
nand U13754 (N_13754,N_8606,N_8819);
nor U13755 (N_13755,N_7352,N_7614);
or U13756 (N_13756,N_8373,N_7148);
and U13757 (N_13757,N_5068,N_6509);
or U13758 (N_13758,N_7507,N_5330);
nor U13759 (N_13759,N_9565,N_5291);
xnor U13760 (N_13760,N_5605,N_6755);
nand U13761 (N_13761,N_5901,N_9675);
or U13762 (N_13762,N_8013,N_5210);
nand U13763 (N_13763,N_8641,N_5906);
and U13764 (N_13764,N_9395,N_5355);
nor U13765 (N_13765,N_7512,N_8863);
and U13766 (N_13766,N_8796,N_5007);
nand U13767 (N_13767,N_5257,N_9482);
nor U13768 (N_13768,N_5884,N_6457);
and U13769 (N_13769,N_8463,N_8965);
or U13770 (N_13770,N_8553,N_6748);
and U13771 (N_13771,N_6445,N_9596);
nor U13772 (N_13772,N_7044,N_7227);
nor U13773 (N_13773,N_8149,N_6030);
nand U13774 (N_13774,N_6202,N_7971);
or U13775 (N_13775,N_9104,N_8818);
nor U13776 (N_13776,N_5372,N_7343);
and U13777 (N_13777,N_8490,N_6762);
or U13778 (N_13778,N_9265,N_7624);
nor U13779 (N_13779,N_8646,N_5749);
and U13780 (N_13780,N_5112,N_8986);
or U13781 (N_13781,N_8184,N_9975);
or U13782 (N_13782,N_9184,N_7069);
nor U13783 (N_13783,N_8437,N_8663);
or U13784 (N_13784,N_8262,N_9300);
xor U13785 (N_13785,N_6688,N_8693);
or U13786 (N_13786,N_5759,N_8748);
or U13787 (N_13787,N_8334,N_6893);
and U13788 (N_13788,N_8695,N_9879);
nand U13789 (N_13789,N_8708,N_6172);
or U13790 (N_13790,N_8812,N_8737);
xnor U13791 (N_13791,N_7380,N_9015);
nand U13792 (N_13792,N_5291,N_5025);
or U13793 (N_13793,N_9906,N_9430);
nand U13794 (N_13794,N_8892,N_9660);
nor U13795 (N_13795,N_6119,N_7419);
or U13796 (N_13796,N_7006,N_6947);
or U13797 (N_13797,N_9101,N_5053);
and U13798 (N_13798,N_8351,N_7207);
nand U13799 (N_13799,N_7728,N_7844);
and U13800 (N_13800,N_7912,N_7683);
or U13801 (N_13801,N_7401,N_8049);
nand U13802 (N_13802,N_6065,N_9754);
xor U13803 (N_13803,N_9515,N_7045);
nor U13804 (N_13804,N_5815,N_5826);
nor U13805 (N_13805,N_7134,N_9837);
nand U13806 (N_13806,N_8726,N_5413);
nor U13807 (N_13807,N_9691,N_8851);
and U13808 (N_13808,N_7721,N_7599);
nand U13809 (N_13809,N_7874,N_9567);
and U13810 (N_13810,N_5292,N_9435);
and U13811 (N_13811,N_6012,N_6927);
nor U13812 (N_13812,N_8074,N_5561);
nor U13813 (N_13813,N_7610,N_5931);
and U13814 (N_13814,N_5064,N_6310);
xor U13815 (N_13815,N_7292,N_5626);
and U13816 (N_13816,N_5486,N_6320);
nand U13817 (N_13817,N_9436,N_5168);
nor U13818 (N_13818,N_7390,N_7114);
and U13819 (N_13819,N_5771,N_5010);
and U13820 (N_13820,N_5213,N_8029);
and U13821 (N_13821,N_8997,N_5152);
and U13822 (N_13822,N_6400,N_6809);
or U13823 (N_13823,N_7955,N_6060);
xor U13824 (N_13824,N_6037,N_9553);
and U13825 (N_13825,N_7589,N_7907);
nand U13826 (N_13826,N_7374,N_7724);
nand U13827 (N_13827,N_6938,N_7935);
nor U13828 (N_13828,N_7499,N_7612);
and U13829 (N_13829,N_8227,N_9322);
and U13830 (N_13830,N_8714,N_8610);
xnor U13831 (N_13831,N_6981,N_9574);
nand U13832 (N_13832,N_9749,N_6904);
or U13833 (N_13833,N_8109,N_9791);
nor U13834 (N_13834,N_5596,N_9088);
nor U13835 (N_13835,N_5625,N_8986);
and U13836 (N_13836,N_8310,N_6538);
nor U13837 (N_13837,N_6156,N_6505);
and U13838 (N_13838,N_8472,N_9848);
nor U13839 (N_13839,N_9544,N_6952);
nand U13840 (N_13840,N_6216,N_5912);
xnor U13841 (N_13841,N_5439,N_7629);
nor U13842 (N_13842,N_5818,N_5382);
and U13843 (N_13843,N_9592,N_5925);
or U13844 (N_13844,N_7450,N_7075);
nor U13845 (N_13845,N_9723,N_5899);
and U13846 (N_13846,N_7238,N_5526);
nor U13847 (N_13847,N_8306,N_7806);
and U13848 (N_13848,N_6765,N_8177);
and U13849 (N_13849,N_6974,N_9109);
nor U13850 (N_13850,N_6442,N_6114);
xor U13851 (N_13851,N_6787,N_9325);
nor U13852 (N_13852,N_6480,N_7585);
nor U13853 (N_13853,N_9244,N_5831);
nor U13854 (N_13854,N_7465,N_7329);
and U13855 (N_13855,N_6455,N_9372);
or U13856 (N_13856,N_6163,N_6830);
or U13857 (N_13857,N_6579,N_7270);
or U13858 (N_13858,N_5751,N_6362);
and U13859 (N_13859,N_8941,N_6221);
or U13860 (N_13860,N_8559,N_8565);
xnor U13861 (N_13861,N_7354,N_5904);
nor U13862 (N_13862,N_6899,N_8468);
nor U13863 (N_13863,N_6448,N_8357);
and U13864 (N_13864,N_6581,N_6907);
nor U13865 (N_13865,N_8301,N_8193);
and U13866 (N_13866,N_8532,N_6044);
nand U13867 (N_13867,N_8431,N_8711);
and U13868 (N_13868,N_6148,N_6130);
nor U13869 (N_13869,N_8806,N_6337);
nor U13870 (N_13870,N_7359,N_8336);
and U13871 (N_13871,N_9842,N_7117);
xor U13872 (N_13872,N_5230,N_5121);
nor U13873 (N_13873,N_6377,N_9494);
nand U13874 (N_13874,N_5950,N_8493);
and U13875 (N_13875,N_6392,N_5616);
xor U13876 (N_13876,N_5455,N_6654);
and U13877 (N_13877,N_9235,N_8205);
nor U13878 (N_13878,N_9371,N_9440);
nand U13879 (N_13879,N_5540,N_8594);
xnor U13880 (N_13880,N_6774,N_5201);
xnor U13881 (N_13881,N_5721,N_7880);
and U13882 (N_13882,N_7837,N_6222);
nand U13883 (N_13883,N_9331,N_7979);
nor U13884 (N_13884,N_9800,N_5612);
nand U13885 (N_13885,N_8493,N_7405);
nand U13886 (N_13886,N_5603,N_9435);
nor U13887 (N_13887,N_6351,N_9760);
or U13888 (N_13888,N_5504,N_7239);
nor U13889 (N_13889,N_9117,N_7661);
and U13890 (N_13890,N_8792,N_9540);
and U13891 (N_13891,N_7934,N_9555);
nand U13892 (N_13892,N_5329,N_9635);
nand U13893 (N_13893,N_5516,N_7152);
nor U13894 (N_13894,N_5839,N_6481);
nand U13895 (N_13895,N_5294,N_9465);
nand U13896 (N_13896,N_7180,N_5563);
and U13897 (N_13897,N_6143,N_6482);
and U13898 (N_13898,N_7659,N_5916);
and U13899 (N_13899,N_5181,N_5567);
nor U13900 (N_13900,N_6065,N_9115);
or U13901 (N_13901,N_6679,N_9413);
nand U13902 (N_13902,N_7664,N_8069);
or U13903 (N_13903,N_7812,N_7412);
or U13904 (N_13904,N_6940,N_7412);
nand U13905 (N_13905,N_6785,N_9049);
and U13906 (N_13906,N_6435,N_7151);
nor U13907 (N_13907,N_6810,N_9408);
nor U13908 (N_13908,N_8935,N_8221);
or U13909 (N_13909,N_5804,N_8684);
nor U13910 (N_13910,N_7051,N_9609);
nand U13911 (N_13911,N_9217,N_5996);
or U13912 (N_13912,N_6091,N_5873);
or U13913 (N_13913,N_8746,N_9621);
or U13914 (N_13914,N_7753,N_6515);
nand U13915 (N_13915,N_6418,N_8685);
nand U13916 (N_13916,N_6763,N_8308);
or U13917 (N_13917,N_5874,N_6796);
xor U13918 (N_13918,N_7606,N_8597);
xnor U13919 (N_13919,N_6153,N_7014);
and U13920 (N_13920,N_7954,N_9645);
or U13921 (N_13921,N_6177,N_8873);
nand U13922 (N_13922,N_8775,N_8616);
nor U13923 (N_13923,N_9327,N_7126);
nor U13924 (N_13924,N_6739,N_7265);
and U13925 (N_13925,N_8873,N_6835);
and U13926 (N_13926,N_6602,N_9589);
or U13927 (N_13927,N_8627,N_9098);
nand U13928 (N_13928,N_9415,N_7733);
and U13929 (N_13929,N_8135,N_6143);
or U13930 (N_13930,N_7044,N_9330);
or U13931 (N_13931,N_7941,N_9113);
or U13932 (N_13932,N_6152,N_7158);
nor U13933 (N_13933,N_9659,N_7845);
or U13934 (N_13934,N_8305,N_9894);
and U13935 (N_13935,N_7818,N_5451);
nor U13936 (N_13936,N_6508,N_8035);
xor U13937 (N_13937,N_9595,N_6702);
nand U13938 (N_13938,N_9801,N_9404);
nor U13939 (N_13939,N_9853,N_7854);
and U13940 (N_13940,N_6560,N_5873);
and U13941 (N_13941,N_9738,N_9987);
nor U13942 (N_13942,N_9668,N_8842);
or U13943 (N_13943,N_6308,N_6170);
nand U13944 (N_13944,N_5468,N_5824);
or U13945 (N_13945,N_8195,N_5793);
nor U13946 (N_13946,N_5531,N_5363);
or U13947 (N_13947,N_6998,N_8867);
and U13948 (N_13948,N_5706,N_8967);
and U13949 (N_13949,N_7825,N_8634);
and U13950 (N_13950,N_9918,N_9032);
nand U13951 (N_13951,N_8075,N_6979);
or U13952 (N_13952,N_7647,N_7221);
and U13953 (N_13953,N_5368,N_7303);
nand U13954 (N_13954,N_8773,N_5282);
nor U13955 (N_13955,N_8711,N_8074);
and U13956 (N_13956,N_7882,N_5813);
xor U13957 (N_13957,N_5759,N_8728);
and U13958 (N_13958,N_6263,N_8002);
nand U13959 (N_13959,N_5344,N_7822);
nand U13960 (N_13960,N_5690,N_9264);
or U13961 (N_13961,N_9458,N_7482);
nor U13962 (N_13962,N_8631,N_5968);
nor U13963 (N_13963,N_6291,N_9420);
and U13964 (N_13964,N_7437,N_5619);
and U13965 (N_13965,N_5673,N_7982);
nand U13966 (N_13966,N_7573,N_9425);
nor U13967 (N_13967,N_7014,N_8418);
xnor U13968 (N_13968,N_7645,N_9510);
or U13969 (N_13969,N_7558,N_6087);
nor U13970 (N_13970,N_6645,N_5768);
nand U13971 (N_13971,N_7250,N_6542);
nand U13972 (N_13972,N_6170,N_8757);
nand U13973 (N_13973,N_6267,N_8560);
xnor U13974 (N_13974,N_8472,N_5078);
xor U13975 (N_13975,N_5922,N_7590);
nand U13976 (N_13976,N_8668,N_9062);
nor U13977 (N_13977,N_9672,N_8267);
and U13978 (N_13978,N_6509,N_5579);
and U13979 (N_13979,N_7549,N_6356);
xnor U13980 (N_13980,N_7414,N_5160);
or U13981 (N_13981,N_5987,N_9741);
and U13982 (N_13982,N_6646,N_6331);
and U13983 (N_13983,N_6495,N_6511);
nand U13984 (N_13984,N_6496,N_5314);
nor U13985 (N_13985,N_7110,N_5408);
and U13986 (N_13986,N_8956,N_7295);
or U13987 (N_13987,N_6758,N_8748);
xor U13988 (N_13988,N_6238,N_8452);
and U13989 (N_13989,N_8326,N_6504);
nor U13990 (N_13990,N_8723,N_8374);
nand U13991 (N_13991,N_8324,N_8167);
nor U13992 (N_13992,N_5085,N_6566);
and U13993 (N_13993,N_6973,N_6297);
nand U13994 (N_13994,N_5380,N_9020);
xor U13995 (N_13995,N_8204,N_8949);
or U13996 (N_13996,N_8104,N_8600);
or U13997 (N_13997,N_7150,N_5441);
and U13998 (N_13998,N_7654,N_6546);
or U13999 (N_13999,N_9924,N_7262);
and U14000 (N_14000,N_8380,N_6523);
or U14001 (N_14001,N_7493,N_6571);
nor U14002 (N_14002,N_9686,N_6598);
nor U14003 (N_14003,N_5149,N_9926);
and U14004 (N_14004,N_6293,N_7014);
nand U14005 (N_14005,N_9020,N_9629);
and U14006 (N_14006,N_5849,N_7086);
and U14007 (N_14007,N_6644,N_7108);
xnor U14008 (N_14008,N_7518,N_9355);
or U14009 (N_14009,N_7455,N_7229);
nor U14010 (N_14010,N_7292,N_8725);
and U14011 (N_14011,N_7314,N_8041);
nor U14012 (N_14012,N_5398,N_5748);
or U14013 (N_14013,N_9146,N_8830);
nor U14014 (N_14014,N_9413,N_6417);
and U14015 (N_14015,N_9850,N_8998);
nor U14016 (N_14016,N_5813,N_6120);
nand U14017 (N_14017,N_9119,N_9247);
nand U14018 (N_14018,N_6226,N_5627);
nand U14019 (N_14019,N_6038,N_7730);
and U14020 (N_14020,N_8903,N_6815);
or U14021 (N_14021,N_7334,N_8021);
nor U14022 (N_14022,N_8711,N_9134);
or U14023 (N_14023,N_5302,N_5370);
or U14024 (N_14024,N_5703,N_7277);
nor U14025 (N_14025,N_6869,N_7762);
nand U14026 (N_14026,N_6192,N_6029);
or U14027 (N_14027,N_5404,N_6402);
and U14028 (N_14028,N_5321,N_8958);
nor U14029 (N_14029,N_6961,N_6045);
and U14030 (N_14030,N_5417,N_7979);
nand U14031 (N_14031,N_7958,N_8530);
and U14032 (N_14032,N_6034,N_8964);
or U14033 (N_14033,N_7534,N_7256);
nand U14034 (N_14034,N_7463,N_6846);
xnor U14035 (N_14035,N_5285,N_5015);
nand U14036 (N_14036,N_6937,N_5836);
nand U14037 (N_14037,N_7198,N_9475);
and U14038 (N_14038,N_8271,N_5564);
nand U14039 (N_14039,N_7283,N_8747);
or U14040 (N_14040,N_7838,N_8150);
and U14041 (N_14041,N_6900,N_7044);
or U14042 (N_14042,N_5583,N_6542);
or U14043 (N_14043,N_5285,N_9200);
nor U14044 (N_14044,N_5201,N_7588);
nor U14045 (N_14045,N_9579,N_7806);
nand U14046 (N_14046,N_8501,N_7562);
or U14047 (N_14047,N_5880,N_6147);
and U14048 (N_14048,N_6157,N_8822);
or U14049 (N_14049,N_8347,N_7370);
or U14050 (N_14050,N_5817,N_8598);
nor U14051 (N_14051,N_8524,N_8540);
or U14052 (N_14052,N_6858,N_9585);
or U14053 (N_14053,N_6402,N_7022);
nor U14054 (N_14054,N_7998,N_6187);
or U14055 (N_14055,N_7128,N_9502);
or U14056 (N_14056,N_5039,N_5574);
or U14057 (N_14057,N_8264,N_9031);
nor U14058 (N_14058,N_6041,N_7789);
nand U14059 (N_14059,N_6143,N_6240);
xor U14060 (N_14060,N_9701,N_5083);
or U14061 (N_14061,N_7498,N_7199);
xnor U14062 (N_14062,N_5427,N_6044);
nand U14063 (N_14063,N_8693,N_9196);
or U14064 (N_14064,N_5776,N_6480);
or U14065 (N_14065,N_9334,N_6464);
nand U14066 (N_14066,N_9203,N_8962);
and U14067 (N_14067,N_5581,N_6954);
nand U14068 (N_14068,N_8258,N_8621);
nand U14069 (N_14069,N_5295,N_5595);
and U14070 (N_14070,N_8492,N_7795);
nor U14071 (N_14071,N_5940,N_9100);
or U14072 (N_14072,N_8202,N_8766);
nor U14073 (N_14073,N_9869,N_6584);
or U14074 (N_14074,N_9437,N_9245);
nand U14075 (N_14075,N_6804,N_9245);
nor U14076 (N_14076,N_6120,N_6491);
or U14077 (N_14077,N_6151,N_7206);
or U14078 (N_14078,N_8648,N_6032);
nor U14079 (N_14079,N_9162,N_5534);
nor U14080 (N_14080,N_7523,N_9434);
nor U14081 (N_14081,N_8262,N_7335);
and U14082 (N_14082,N_7235,N_5064);
or U14083 (N_14083,N_7711,N_7806);
nand U14084 (N_14084,N_5855,N_9695);
and U14085 (N_14085,N_6047,N_6186);
nand U14086 (N_14086,N_7113,N_9062);
nor U14087 (N_14087,N_7752,N_5458);
nor U14088 (N_14088,N_5940,N_9630);
xnor U14089 (N_14089,N_7121,N_7729);
and U14090 (N_14090,N_6396,N_9026);
or U14091 (N_14091,N_6850,N_6225);
nor U14092 (N_14092,N_7408,N_7883);
nor U14093 (N_14093,N_7614,N_5894);
nor U14094 (N_14094,N_7453,N_5409);
nand U14095 (N_14095,N_7945,N_8210);
nand U14096 (N_14096,N_5078,N_9428);
nand U14097 (N_14097,N_6364,N_8854);
nand U14098 (N_14098,N_8224,N_5429);
nor U14099 (N_14099,N_5906,N_8831);
and U14100 (N_14100,N_9259,N_5877);
nor U14101 (N_14101,N_6967,N_7358);
or U14102 (N_14102,N_9752,N_5486);
nand U14103 (N_14103,N_7395,N_8381);
or U14104 (N_14104,N_5924,N_8146);
or U14105 (N_14105,N_9562,N_8047);
or U14106 (N_14106,N_7381,N_5389);
or U14107 (N_14107,N_6496,N_9540);
or U14108 (N_14108,N_9329,N_5115);
nor U14109 (N_14109,N_5353,N_5024);
nor U14110 (N_14110,N_8884,N_6066);
nor U14111 (N_14111,N_7307,N_7119);
nor U14112 (N_14112,N_9374,N_8496);
and U14113 (N_14113,N_8572,N_6398);
nor U14114 (N_14114,N_9200,N_9182);
or U14115 (N_14115,N_6045,N_8699);
and U14116 (N_14116,N_8129,N_5636);
or U14117 (N_14117,N_9935,N_7717);
nor U14118 (N_14118,N_6552,N_6489);
and U14119 (N_14119,N_6032,N_9041);
nand U14120 (N_14120,N_5911,N_9475);
xnor U14121 (N_14121,N_7046,N_6397);
and U14122 (N_14122,N_5811,N_5661);
nand U14123 (N_14123,N_7074,N_6813);
nor U14124 (N_14124,N_5946,N_6284);
xnor U14125 (N_14125,N_7975,N_7378);
or U14126 (N_14126,N_8041,N_8256);
or U14127 (N_14127,N_7003,N_8485);
nand U14128 (N_14128,N_9643,N_6460);
or U14129 (N_14129,N_8139,N_6571);
nand U14130 (N_14130,N_9638,N_7905);
and U14131 (N_14131,N_8177,N_5503);
or U14132 (N_14132,N_9505,N_7221);
nor U14133 (N_14133,N_9060,N_9852);
xor U14134 (N_14134,N_7806,N_7953);
nand U14135 (N_14135,N_5544,N_9964);
and U14136 (N_14136,N_6456,N_9944);
nand U14137 (N_14137,N_7548,N_9027);
xor U14138 (N_14138,N_8308,N_6174);
nor U14139 (N_14139,N_8030,N_6960);
and U14140 (N_14140,N_6632,N_9311);
or U14141 (N_14141,N_9556,N_7235);
and U14142 (N_14142,N_7510,N_6906);
nand U14143 (N_14143,N_9948,N_8806);
nand U14144 (N_14144,N_8828,N_5366);
and U14145 (N_14145,N_8649,N_5844);
and U14146 (N_14146,N_9211,N_5468);
nand U14147 (N_14147,N_8547,N_8729);
nand U14148 (N_14148,N_9428,N_6721);
and U14149 (N_14149,N_8959,N_9502);
and U14150 (N_14150,N_8594,N_8769);
or U14151 (N_14151,N_5746,N_5974);
nor U14152 (N_14152,N_9162,N_6863);
xor U14153 (N_14153,N_7867,N_6629);
or U14154 (N_14154,N_6528,N_6135);
and U14155 (N_14155,N_5961,N_9291);
or U14156 (N_14156,N_6350,N_5065);
nand U14157 (N_14157,N_8426,N_9430);
nand U14158 (N_14158,N_6662,N_8274);
and U14159 (N_14159,N_9898,N_7041);
and U14160 (N_14160,N_5948,N_6253);
nand U14161 (N_14161,N_5170,N_5668);
nor U14162 (N_14162,N_9610,N_6954);
and U14163 (N_14163,N_6534,N_7608);
or U14164 (N_14164,N_5355,N_8725);
or U14165 (N_14165,N_7286,N_5458);
and U14166 (N_14166,N_9001,N_5916);
and U14167 (N_14167,N_8281,N_6563);
and U14168 (N_14168,N_6404,N_8975);
and U14169 (N_14169,N_8149,N_7239);
nand U14170 (N_14170,N_6527,N_8137);
or U14171 (N_14171,N_7186,N_8358);
and U14172 (N_14172,N_5020,N_9893);
and U14173 (N_14173,N_9707,N_6119);
nor U14174 (N_14174,N_9113,N_9651);
nor U14175 (N_14175,N_8867,N_5552);
nand U14176 (N_14176,N_5812,N_8994);
and U14177 (N_14177,N_5398,N_8247);
nor U14178 (N_14178,N_7116,N_7210);
nand U14179 (N_14179,N_8288,N_8950);
and U14180 (N_14180,N_8250,N_5440);
nand U14181 (N_14181,N_5204,N_7920);
nand U14182 (N_14182,N_5565,N_6601);
nand U14183 (N_14183,N_7244,N_9058);
and U14184 (N_14184,N_7479,N_7422);
or U14185 (N_14185,N_7734,N_6994);
nand U14186 (N_14186,N_7811,N_5984);
or U14187 (N_14187,N_6545,N_7456);
nor U14188 (N_14188,N_6716,N_9234);
or U14189 (N_14189,N_8395,N_8157);
and U14190 (N_14190,N_8300,N_5792);
nand U14191 (N_14191,N_5033,N_8119);
nor U14192 (N_14192,N_8352,N_7286);
or U14193 (N_14193,N_8912,N_6346);
xnor U14194 (N_14194,N_5347,N_7918);
nor U14195 (N_14195,N_5443,N_5002);
or U14196 (N_14196,N_5057,N_7125);
nand U14197 (N_14197,N_8237,N_7870);
nand U14198 (N_14198,N_5854,N_5699);
and U14199 (N_14199,N_9976,N_7942);
and U14200 (N_14200,N_8232,N_9115);
and U14201 (N_14201,N_6938,N_7442);
nand U14202 (N_14202,N_9019,N_9512);
or U14203 (N_14203,N_6220,N_7877);
or U14204 (N_14204,N_7287,N_7297);
nor U14205 (N_14205,N_6024,N_6218);
xnor U14206 (N_14206,N_5703,N_9059);
xor U14207 (N_14207,N_7130,N_6584);
or U14208 (N_14208,N_8952,N_7296);
or U14209 (N_14209,N_9956,N_5821);
nor U14210 (N_14210,N_7540,N_9639);
xor U14211 (N_14211,N_5196,N_7769);
nor U14212 (N_14212,N_5030,N_8840);
nor U14213 (N_14213,N_5194,N_8811);
or U14214 (N_14214,N_8360,N_7854);
and U14215 (N_14215,N_7412,N_7768);
nand U14216 (N_14216,N_5552,N_9826);
xnor U14217 (N_14217,N_7978,N_8666);
or U14218 (N_14218,N_5027,N_5182);
nand U14219 (N_14219,N_8341,N_7133);
nor U14220 (N_14220,N_6321,N_9738);
and U14221 (N_14221,N_8862,N_6816);
nand U14222 (N_14222,N_9973,N_6722);
and U14223 (N_14223,N_5620,N_5240);
xnor U14224 (N_14224,N_5433,N_7173);
nor U14225 (N_14225,N_6101,N_9655);
or U14226 (N_14226,N_7875,N_6542);
nor U14227 (N_14227,N_7833,N_6437);
and U14228 (N_14228,N_7195,N_5223);
nor U14229 (N_14229,N_7047,N_5506);
and U14230 (N_14230,N_7825,N_7522);
xor U14231 (N_14231,N_6270,N_6327);
nor U14232 (N_14232,N_6568,N_9617);
xnor U14233 (N_14233,N_9477,N_9564);
nand U14234 (N_14234,N_8117,N_8660);
nand U14235 (N_14235,N_8774,N_5254);
nand U14236 (N_14236,N_5268,N_5546);
or U14237 (N_14237,N_9798,N_7126);
and U14238 (N_14238,N_8932,N_8389);
nand U14239 (N_14239,N_7055,N_7488);
nand U14240 (N_14240,N_5277,N_9337);
nor U14241 (N_14241,N_9763,N_9771);
and U14242 (N_14242,N_9752,N_6461);
or U14243 (N_14243,N_8391,N_6175);
nor U14244 (N_14244,N_9170,N_8468);
nor U14245 (N_14245,N_8762,N_8695);
nand U14246 (N_14246,N_7940,N_9305);
and U14247 (N_14247,N_6802,N_6970);
xnor U14248 (N_14248,N_9277,N_5882);
nor U14249 (N_14249,N_7517,N_9593);
nor U14250 (N_14250,N_9196,N_9336);
and U14251 (N_14251,N_5305,N_8387);
and U14252 (N_14252,N_9354,N_6902);
xor U14253 (N_14253,N_7109,N_8768);
and U14254 (N_14254,N_7648,N_5583);
and U14255 (N_14255,N_9772,N_5670);
nor U14256 (N_14256,N_7542,N_5202);
nor U14257 (N_14257,N_9668,N_9568);
nand U14258 (N_14258,N_6145,N_6477);
and U14259 (N_14259,N_8169,N_8688);
and U14260 (N_14260,N_6551,N_7579);
or U14261 (N_14261,N_5194,N_5578);
and U14262 (N_14262,N_7002,N_5133);
or U14263 (N_14263,N_8382,N_8977);
nand U14264 (N_14264,N_7493,N_5680);
nor U14265 (N_14265,N_9080,N_6650);
nor U14266 (N_14266,N_8766,N_7879);
nand U14267 (N_14267,N_6064,N_6733);
nand U14268 (N_14268,N_6380,N_6105);
nor U14269 (N_14269,N_8274,N_5764);
nand U14270 (N_14270,N_9907,N_8588);
and U14271 (N_14271,N_5641,N_7695);
and U14272 (N_14272,N_8420,N_5522);
nand U14273 (N_14273,N_7482,N_5939);
nand U14274 (N_14274,N_8241,N_7178);
nor U14275 (N_14275,N_9843,N_6951);
and U14276 (N_14276,N_7075,N_7007);
or U14277 (N_14277,N_6967,N_8402);
nand U14278 (N_14278,N_5114,N_5468);
xor U14279 (N_14279,N_8240,N_5155);
or U14280 (N_14280,N_5238,N_7725);
nand U14281 (N_14281,N_6931,N_5493);
or U14282 (N_14282,N_9444,N_7341);
nand U14283 (N_14283,N_7964,N_9298);
and U14284 (N_14284,N_9412,N_5843);
nand U14285 (N_14285,N_7627,N_5600);
nand U14286 (N_14286,N_6234,N_8439);
nor U14287 (N_14287,N_9120,N_8570);
nand U14288 (N_14288,N_7357,N_7865);
nand U14289 (N_14289,N_8775,N_6810);
or U14290 (N_14290,N_8008,N_7870);
nand U14291 (N_14291,N_7649,N_7828);
xor U14292 (N_14292,N_6502,N_9959);
nor U14293 (N_14293,N_5363,N_6872);
nand U14294 (N_14294,N_7281,N_8718);
xnor U14295 (N_14295,N_5734,N_9041);
xor U14296 (N_14296,N_9236,N_5113);
and U14297 (N_14297,N_7389,N_5017);
nor U14298 (N_14298,N_9492,N_9883);
nor U14299 (N_14299,N_7674,N_8885);
nor U14300 (N_14300,N_7682,N_5049);
and U14301 (N_14301,N_9150,N_5944);
and U14302 (N_14302,N_8804,N_7441);
xor U14303 (N_14303,N_6064,N_6391);
or U14304 (N_14304,N_7079,N_9049);
nand U14305 (N_14305,N_5156,N_8365);
xnor U14306 (N_14306,N_6659,N_5836);
and U14307 (N_14307,N_8773,N_5012);
xnor U14308 (N_14308,N_6214,N_6769);
and U14309 (N_14309,N_5967,N_8488);
nand U14310 (N_14310,N_9259,N_5868);
or U14311 (N_14311,N_9877,N_5958);
nand U14312 (N_14312,N_5620,N_9323);
or U14313 (N_14313,N_6065,N_6775);
or U14314 (N_14314,N_5281,N_8951);
xor U14315 (N_14315,N_8313,N_9075);
nand U14316 (N_14316,N_8791,N_8469);
and U14317 (N_14317,N_9010,N_9556);
nor U14318 (N_14318,N_6760,N_8133);
nand U14319 (N_14319,N_5224,N_9982);
nor U14320 (N_14320,N_6050,N_9802);
nor U14321 (N_14321,N_9212,N_8740);
nand U14322 (N_14322,N_5878,N_6554);
or U14323 (N_14323,N_8542,N_7112);
and U14324 (N_14324,N_6950,N_9137);
nor U14325 (N_14325,N_8916,N_5306);
nand U14326 (N_14326,N_7102,N_8881);
nor U14327 (N_14327,N_6985,N_5573);
and U14328 (N_14328,N_9922,N_8770);
and U14329 (N_14329,N_8010,N_7303);
or U14330 (N_14330,N_5994,N_5655);
or U14331 (N_14331,N_7876,N_6788);
nor U14332 (N_14332,N_7615,N_5692);
and U14333 (N_14333,N_6252,N_5048);
and U14334 (N_14334,N_9292,N_8612);
nand U14335 (N_14335,N_8913,N_7135);
and U14336 (N_14336,N_8743,N_8173);
nor U14337 (N_14337,N_9060,N_7574);
nor U14338 (N_14338,N_8528,N_8414);
and U14339 (N_14339,N_9197,N_8025);
and U14340 (N_14340,N_9800,N_5023);
or U14341 (N_14341,N_9355,N_6319);
and U14342 (N_14342,N_6488,N_7765);
nor U14343 (N_14343,N_7918,N_5627);
nand U14344 (N_14344,N_8892,N_9307);
nand U14345 (N_14345,N_5733,N_5155);
xnor U14346 (N_14346,N_5726,N_9202);
or U14347 (N_14347,N_8399,N_9428);
nand U14348 (N_14348,N_6014,N_7896);
nor U14349 (N_14349,N_7837,N_6743);
nand U14350 (N_14350,N_8166,N_6072);
and U14351 (N_14351,N_8057,N_7187);
nor U14352 (N_14352,N_5263,N_6485);
nor U14353 (N_14353,N_9146,N_8067);
xor U14354 (N_14354,N_8789,N_7266);
nand U14355 (N_14355,N_9330,N_8680);
nor U14356 (N_14356,N_8841,N_5042);
nand U14357 (N_14357,N_9486,N_5512);
nor U14358 (N_14358,N_8187,N_8217);
and U14359 (N_14359,N_7192,N_5458);
nor U14360 (N_14360,N_5958,N_6838);
nand U14361 (N_14361,N_9559,N_8656);
nand U14362 (N_14362,N_9807,N_6080);
and U14363 (N_14363,N_5627,N_8379);
or U14364 (N_14364,N_6399,N_7807);
xnor U14365 (N_14365,N_8389,N_5686);
nor U14366 (N_14366,N_6256,N_6436);
nand U14367 (N_14367,N_7042,N_6969);
and U14368 (N_14368,N_5477,N_9795);
nor U14369 (N_14369,N_5079,N_8714);
nor U14370 (N_14370,N_5465,N_7837);
nand U14371 (N_14371,N_5499,N_9599);
nand U14372 (N_14372,N_5333,N_9389);
or U14373 (N_14373,N_9620,N_7024);
and U14374 (N_14374,N_5260,N_9772);
xor U14375 (N_14375,N_9668,N_8151);
and U14376 (N_14376,N_6436,N_5572);
and U14377 (N_14377,N_7277,N_7849);
nor U14378 (N_14378,N_8704,N_7239);
nor U14379 (N_14379,N_6999,N_5165);
or U14380 (N_14380,N_8830,N_9122);
and U14381 (N_14381,N_8542,N_8189);
and U14382 (N_14382,N_7000,N_9180);
nor U14383 (N_14383,N_6611,N_8329);
or U14384 (N_14384,N_7868,N_6176);
nand U14385 (N_14385,N_6534,N_9234);
nor U14386 (N_14386,N_5216,N_6423);
and U14387 (N_14387,N_5303,N_9834);
and U14388 (N_14388,N_8766,N_8564);
or U14389 (N_14389,N_7213,N_7394);
nor U14390 (N_14390,N_6831,N_6010);
xnor U14391 (N_14391,N_6717,N_7686);
nand U14392 (N_14392,N_6852,N_5552);
and U14393 (N_14393,N_7481,N_6269);
or U14394 (N_14394,N_6920,N_8612);
nand U14395 (N_14395,N_7457,N_5420);
or U14396 (N_14396,N_5974,N_7664);
or U14397 (N_14397,N_5278,N_8431);
xnor U14398 (N_14398,N_7702,N_5577);
nor U14399 (N_14399,N_7551,N_7863);
or U14400 (N_14400,N_8843,N_7423);
xor U14401 (N_14401,N_6950,N_6765);
or U14402 (N_14402,N_5080,N_5683);
xnor U14403 (N_14403,N_7449,N_5282);
nor U14404 (N_14404,N_8812,N_6946);
or U14405 (N_14405,N_8028,N_5735);
and U14406 (N_14406,N_7440,N_6581);
and U14407 (N_14407,N_8726,N_7394);
and U14408 (N_14408,N_8736,N_9042);
and U14409 (N_14409,N_9926,N_9788);
or U14410 (N_14410,N_8232,N_5770);
or U14411 (N_14411,N_6707,N_8140);
and U14412 (N_14412,N_6392,N_7313);
or U14413 (N_14413,N_6884,N_5677);
nand U14414 (N_14414,N_9756,N_9483);
nor U14415 (N_14415,N_5292,N_8987);
nor U14416 (N_14416,N_7552,N_7225);
nand U14417 (N_14417,N_8848,N_5606);
nand U14418 (N_14418,N_9724,N_7516);
xnor U14419 (N_14419,N_6747,N_6464);
and U14420 (N_14420,N_8569,N_9980);
nand U14421 (N_14421,N_8083,N_6885);
or U14422 (N_14422,N_9435,N_8611);
nand U14423 (N_14423,N_9335,N_9606);
or U14424 (N_14424,N_7243,N_8303);
nor U14425 (N_14425,N_6762,N_6657);
nand U14426 (N_14426,N_7204,N_7358);
or U14427 (N_14427,N_9512,N_6151);
nand U14428 (N_14428,N_5060,N_8364);
nor U14429 (N_14429,N_6938,N_9741);
or U14430 (N_14430,N_7577,N_9935);
nand U14431 (N_14431,N_6018,N_8475);
and U14432 (N_14432,N_7890,N_7766);
or U14433 (N_14433,N_7402,N_7048);
nand U14434 (N_14434,N_8631,N_8268);
xor U14435 (N_14435,N_9879,N_6668);
nand U14436 (N_14436,N_6304,N_7595);
nor U14437 (N_14437,N_7758,N_8184);
nand U14438 (N_14438,N_8937,N_8455);
nor U14439 (N_14439,N_8291,N_6607);
nor U14440 (N_14440,N_9736,N_8038);
nor U14441 (N_14441,N_7279,N_7339);
nor U14442 (N_14442,N_9143,N_9917);
and U14443 (N_14443,N_5125,N_7101);
nor U14444 (N_14444,N_7186,N_8829);
and U14445 (N_14445,N_5751,N_7707);
or U14446 (N_14446,N_6249,N_7796);
and U14447 (N_14447,N_7654,N_7457);
xnor U14448 (N_14448,N_5767,N_5952);
or U14449 (N_14449,N_6297,N_9080);
nand U14450 (N_14450,N_7235,N_9751);
or U14451 (N_14451,N_9112,N_7216);
xnor U14452 (N_14452,N_8909,N_9684);
or U14453 (N_14453,N_5248,N_5466);
and U14454 (N_14454,N_8767,N_9817);
nand U14455 (N_14455,N_8625,N_7511);
and U14456 (N_14456,N_7722,N_9340);
nor U14457 (N_14457,N_6219,N_5384);
nor U14458 (N_14458,N_7280,N_7578);
or U14459 (N_14459,N_8957,N_8606);
and U14460 (N_14460,N_7104,N_6194);
or U14461 (N_14461,N_7667,N_5397);
or U14462 (N_14462,N_8753,N_6921);
nor U14463 (N_14463,N_5417,N_7678);
nand U14464 (N_14464,N_8440,N_7556);
nor U14465 (N_14465,N_6750,N_8876);
or U14466 (N_14466,N_5677,N_6205);
nand U14467 (N_14467,N_9347,N_8195);
and U14468 (N_14468,N_7067,N_6522);
or U14469 (N_14469,N_5439,N_7399);
nand U14470 (N_14470,N_8283,N_7480);
and U14471 (N_14471,N_8994,N_9127);
or U14472 (N_14472,N_5940,N_8621);
nand U14473 (N_14473,N_7718,N_5707);
nor U14474 (N_14474,N_8488,N_9494);
and U14475 (N_14475,N_9670,N_8141);
and U14476 (N_14476,N_7447,N_7674);
or U14477 (N_14477,N_6759,N_9562);
nor U14478 (N_14478,N_8073,N_6596);
xnor U14479 (N_14479,N_7983,N_8057);
nor U14480 (N_14480,N_5611,N_6145);
or U14481 (N_14481,N_6893,N_5529);
xor U14482 (N_14482,N_6341,N_7284);
nand U14483 (N_14483,N_5171,N_8868);
or U14484 (N_14484,N_8163,N_9941);
xor U14485 (N_14485,N_9583,N_9772);
or U14486 (N_14486,N_6202,N_6751);
or U14487 (N_14487,N_8023,N_8492);
or U14488 (N_14488,N_9981,N_9945);
xnor U14489 (N_14489,N_5625,N_7898);
nor U14490 (N_14490,N_9345,N_9887);
nor U14491 (N_14491,N_8114,N_6034);
nor U14492 (N_14492,N_6951,N_7577);
or U14493 (N_14493,N_6512,N_5266);
nand U14494 (N_14494,N_6858,N_9726);
nor U14495 (N_14495,N_6313,N_7593);
and U14496 (N_14496,N_9227,N_5915);
nand U14497 (N_14497,N_9088,N_6967);
nand U14498 (N_14498,N_6896,N_5736);
nor U14499 (N_14499,N_7499,N_8545);
and U14500 (N_14500,N_9789,N_8041);
and U14501 (N_14501,N_6470,N_9987);
nor U14502 (N_14502,N_6803,N_9975);
nor U14503 (N_14503,N_6777,N_6260);
nor U14504 (N_14504,N_6138,N_5182);
nor U14505 (N_14505,N_8210,N_7508);
or U14506 (N_14506,N_7124,N_5436);
or U14507 (N_14507,N_8322,N_5046);
nand U14508 (N_14508,N_5454,N_7146);
xnor U14509 (N_14509,N_5866,N_8184);
and U14510 (N_14510,N_7017,N_9029);
nor U14511 (N_14511,N_9611,N_7051);
or U14512 (N_14512,N_9344,N_9455);
xor U14513 (N_14513,N_6133,N_7681);
nor U14514 (N_14514,N_5352,N_6806);
or U14515 (N_14515,N_5483,N_6289);
or U14516 (N_14516,N_6843,N_7515);
nor U14517 (N_14517,N_6510,N_6290);
or U14518 (N_14518,N_9385,N_6116);
nand U14519 (N_14519,N_6255,N_9232);
or U14520 (N_14520,N_8118,N_5478);
or U14521 (N_14521,N_7176,N_8650);
and U14522 (N_14522,N_7957,N_6906);
and U14523 (N_14523,N_8044,N_8941);
nand U14524 (N_14524,N_9928,N_6034);
and U14525 (N_14525,N_8723,N_8343);
nor U14526 (N_14526,N_9549,N_9286);
nand U14527 (N_14527,N_6570,N_9456);
xor U14528 (N_14528,N_5430,N_7262);
and U14529 (N_14529,N_6502,N_8364);
or U14530 (N_14530,N_6434,N_7552);
and U14531 (N_14531,N_9931,N_6147);
or U14532 (N_14532,N_8541,N_8202);
nand U14533 (N_14533,N_8856,N_8528);
xnor U14534 (N_14534,N_7756,N_9910);
nor U14535 (N_14535,N_8678,N_5173);
or U14536 (N_14536,N_7967,N_8081);
xor U14537 (N_14537,N_8614,N_6565);
or U14538 (N_14538,N_8108,N_9603);
nor U14539 (N_14539,N_8669,N_5295);
nor U14540 (N_14540,N_5054,N_9685);
nand U14541 (N_14541,N_8014,N_8380);
or U14542 (N_14542,N_7616,N_6382);
nand U14543 (N_14543,N_9354,N_7070);
nand U14544 (N_14544,N_8999,N_5201);
nor U14545 (N_14545,N_6925,N_8712);
nor U14546 (N_14546,N_9196,N_8482);
nand U14547 (N_14547,N_8323,N_6497);
and U14548 (N_14548,N_5201,N_5187);
or U14549 (N_14549,N_5801,N_7702);
nand U14550 (N_14550,N_9740,N_7101);
nor U14551 (N_14551,N_7964,N_7260);
nor U14552 (N_14552,N_5229,N_7694);
or U14553 (N_14553,N_8190,N_5178);
and U14554 (N_14554,N_5975,N_9768);
nand U14555 (N_14555,N_7917,N_9448);
nor U14556 (N_14556,N_5337,N_8563);
nand U14557 (N_14557,N_9407,N_7808);
nor U14558 (N_14558,N_7556,N_5867);
xnor U14559 (N_14559,N_8691,N_7375);
xor U14560 (N_14560,N_6316,N_8039);
nand U14561 (N_14561,N_9859,N_5396);
nand U14562 (N_14562,N_9076,N_8894);
nor U14563 (N_14563,N_9225,N_5378);
xor U14564 (N_14564,N_5044,N_6893);
nand U14565 (N_14565,N_5360,N_9925);
or U14566 (N_14566,N_6108,N_8068);
nor U14567 (N_14567,N_6861,N_9081);
nand U14568 (N_14568,N_8250,N_8113);
nor U14569 (N_14569,N_7168,N_9341);
and U14570 (N_14570,N_5894,N_9979);
nand U14571 (N_14571,N_7437,N_8746);
nor U14572 (N_14572,N_8665,N_8274);
nor U14573 (N_14573,N_8810,N_9398);
and U14574 (N_14574,N_5825,N_6935);
or U14575 (N_14575,N_6105,N_6214);
and U14576 (N_14576,N_7750,N_6355);
nand U14577 (N_14577,N_6548,N_5065);
nand U14578 (N_14578,N_8789,N_6622);
nor U14579 (N_14579,N_8491,N_7119);
or U14580 (N_14580,N_8863,N_9467);
nor U14581 (N_14581,N_8562,N_9311);
nor U14582 (N_14582,N_5411,N_5705);
nand U14583 (N_14583,N_9984,N_7041);
or U14584 (N_14584,N_6154,N_8072);
and U14585 (N_14585,N_7317,N_5138);
or U14586 (N_14586,N_7986,N_5127);
nor U14587 (N_14587,N_9143,N_5266);
nand U14588 (N_14588,N_5677,N_8058);
xor U14589 (N_14589,N_7485,N_7974);
nand U14590 (N_14590,N_8966,N_9017);
or U14591 (N_14591,N_9987,N_9198);
nand U14592 (N_14592,N_9088,N_8819);
and U14593 (N_14593,N_6791,N_7561);
and U14594 (N_14594,N_5914,N_5388);
nand U14595 (N_14595,N_9758,N_9964);
or U14596 (N_14596,N_5631,N_9362);
xnor U14597 (N_14597,N_5015,N_5155);
xnor U14598 (N_14598,N_6602,N_9818);
or U14599 (N_14599,N_8729,N_8375);
or U14600 (N_14600,N_7103,N_6024);
and U14601 (N_14601,N_5426,N_5644);
and U14602 (N_14602,N_5064,N_5103);
and U14603 (N_14603,N_5329,N_9091);
xor U14604 (N_14604,N_8991,N_6308);
or U14605 (N_14605,N_8347,N_5908);
or U14606 (N_14606,N_6286,N_7049);
nor U14607 (N_14607,N_6698,N_7878);
nor U14608 (N_14608,N_5419,N_7703);
or U14609 (N_14609,N_7575,N_6923);
and U14610 (N_14610,N_8558,N_8864);
and U14611 (N_14611,N_7341,N_7889);
nand U14612 (N_14612,N_9641,N_8125);
nor U14613 (N_14613,N_7303,N_8489);
nand U14614 (N_14614,N_5792,N_9698);
nand U14615 (N_14615,N_9355,N_9121);
or U14616 (N_14616,N_8362,N_6905);
or U14617 (N_14617,N_7524,N_5825);
nor U14618 (N_14618,N_9183,N_6365);
and U14619 (N_14619,N_9372,N_5589);
nor U14620 (N_14620,N_7757,N_6494);
or U14621 (N_14621,N_6669,N_5009);
nand U14622 (N_14622,N_8804,N_9690);
xnor U14623 (N_14623,N_7430,N_7871);
or U14624 (N_14624,N_7796,N_8902);
or U14625 (N_14625,N_6362,N_7349);
or U14626 (N_14626,N_6513,N_8667);
or U14627 (N_14627,N_7743,N_9206);
or U14628 (N_14628,N_6364,N_7649);
nand U14629 (N_14629,N_5806,N_8037);
or U14630 (N_14630,N_8195,N_9394);
and U14631 (N_14631,N_6227,N_6079);
nand U14632 (N_14632,N_9904,N_8471);
and U14633 (N_14633,N_7535,N_9337);
nor U14634 (N_14634,N_6067,N_8725);
and U14635 (N_14635,N_8355,N_6018);
nand U14636 (N_14636,N_5379,N_9584);
nor U14637 (N_14637,N_9783,N_7032);
nor U14638 (N_14638,N_9445,N_6072);
or U14639 (N_14639,N_8458,N_9368);
xnor U14640 (N_14640,N_7904,N_8906);
or U14641 (N_14641,N_7228,N_8482);
nand U14642 (N_14642,N_8000,N_6514);
nor U14643 (N_14643,N_8314,N_5536);
or U14644 (N_14644,N_9529,N_5003);
and U14645 (N_14645,N_5427,N_8711);
nor U14646 (N_14646,N_7702,N_7992);
nor U14647 (N_14647,N_9333,N_6395);
and U14648 (N_14648,N_7050,N_6560);
or U14649 (N_14649,N_6037,N_6204);
or U14650 (N_14650,N_7320,N_9655);
or U14651 (N_14651,N_8176,N_9331);
xor U14652 (N_14652,N_8042,N_9474);
nor U14653 (N_14653,N_5329,N_8230);
nand U14654 (N_14654,N_6412,N_5163);
nand U14655 (N_14655,N_6543,N_5108);
nand U14656 (N_14656,N_7204,N_8987);
or U14657 (N_14657,N_5460,N_7197);
nand U14658 (N_14658,N_8106,N_5816);
and U14659 (N_14659,N_5538,N_6414);
nor U14660 (N_14660,N_9496,N_5672);
and U14661 (N_14661,N_8744,N_6570);
or U14662 (N_14662,N_8141,N_6870);
nor U14663 (N_14663,N_9355,N_7900);
xor U14664 (N_14664,N_9525,N_7342);
nor U14665 (N_14665,N_7187,N_7891);
or U14666 (N_14666,N_8657,N_6700);
xnor U14667 (N_14667,N_5580,N_9439);
xor U14668 (N_14668,N_9504,N_5718);
nand U14669 (N_14669,N_9159,N_8970);
nand U14670 (N_14670,N_5059,N_5119);
nor U14671 (N_14671,N_6458,N_7017);
nor U14672 (N_14672,N_5127,N_7069);
nor U14673 (N_14673,N_7562,N_8483);
or U14674 (N_14674,N_8044,N_7975);
and U14675 (N_14675,N_5662,N_6738);
nand U14676 (N_14676,N_9675,N_7787);
and U14677 (N_14677,N_7482,N_9878);
xnor U14678 (N_14678,N_7160,N_5087);
nand U14679 (N_14679,N_8976,N_7117);
or U14680 (N_14680,N_7870,N_8409);
nor U14681 (N_14681,N_9394,N_6894);
xnor U14682 (N_14682,N_7050,N_7848);
xor U14683 (N_14683,N_5821,N_9015);
nand U14684 (N_14684,N_7608,N_7875);
nand U14685 (N_14685,N_8593,N_8081);
nand U14686 (N_14686,N_9477,N_5700);
nand U14687 (N_14687,N_8873,N_9700);
or U14688 (N_14688,N_5500,N_6521);
or U14689 (N_14689,N_7414,N_6189);
nand U14690 (N_14690,N_8407,N_5358);
xnor U14691 (N_14691,N_8475,N_9335);
xor U14692 (N_14692,N_7386,N_9779);
nand U14693 (N_14693,N_7020,N_9590);
or U14694 (N_14694,N_8626,N_5604);
or U14695 (N_14695,N_8680,N_8937);
nand U14696 (N_14696,N_7453,N_7365);
or U14697 (N_14697,N_7965,N_7572);
nand U14698 (N_14698,N_5968,N_8577);
nor U14699 (N_14699,N_8804,N_6439);
or U14700 (N_14700,N_6744,N_6313);
nor U14701 (N_14701,N_9855,N_9882);
and U14702 (N_14702,N_6306,N_8221);
nand U14703 (N_14703,N_5932,N_8960);
nor U14704 (N_14704,N_5817,N_9334);
or U14705 (N_14705,N_5755,N_5691);
or U14706 (N_14706,N_8209,N_7063);
and U14707 (N_14707,N_8542,N_9236);
nand U14708 (N_14708,N_8555,N_8786);
nor U14709 (N_14709,N_6980,N_9774);
or U14710 (N_14710,N_7472,N_7195);
nor U14711 (N_14711,N_9671,N_5052);
nand U14712 (N_14712,N_7971,N_5441);
or U14713 (N_14713,N_5793,N_7952);
nor U14714 (N_14714,N_7757,N_6974);
and U14715 (N_14715,N_9329,N_8179);
nand U14716 (N_14716,N_6499,N_8648);
nor U14717 (N_14717,N_8784,N_6955);
nand U14718 (N_14718,N_7714,N_8261);
xor U14719 (N_14719,N_8093,N_5886);
nand U14720 (N_14720,N_7042,N_6648);
and U14721 (N_14721,N_6939,N_8926);
or U14722 (N_14722,N_7305,N_6529);
or U14723 (N_14723,N_9583,N_6800);
nor U14724 (N_14724,N_6938,N_9011);
xnor U14725 (N_14725,N_5749,N_9624);
nor U14726 (N_14726,N_9449,N_7483);
and U14727 (N_14727,N_9450,N_6023);
nand U14728 (N_14728,N_6461,N_5498);
or U14729 (N_14729,N_6867,N_5079);
and U14730 (N_14730,N_7741,N_7116);
nor U14731 (N_14731,N_5900,N_8417);
nand U14732 (N_14732,N_6138,N_8303);
nor U14733 (N_14733,N_6395,N_5230);
and U14734 (N_14734,N_6301,N_7109);
nor U14735 (N_14735,N_5815,N_6690);
nand U14736 (N_14736,N_5555,N_7791);
nand U14737 (N_14737,N_8387,N_7236);
xnor U14738 (N_14738,N_5118,N_9544);
and U14739 (N_14739,N_9920,N_6915);
nand U14740 (N_14740,N_7996,N_6150);
nand U14741 (N_14741,N_6718,N_5809);
nand U14742 (N_14742,N_7803,N_5971);
and U14743 (N_14743,N_6604,N_6148);
or U14744 (N_14744,N_8756,N_7363);
nand U14745 (N_14745,N_9430,N_6223);
and U14746 (N_14746,N_8518,N_9883);
or U14747 (N_14747,N_8186,N_5127);
and U14748 (N_14748,N_9329,N_9543);
xor U14749 (N_14749,N_9634,N_8027);
nand U14750 (N_14750,N_7957,N_5930);
nand U14751 (N_14751,N_8766,N_9724);
and U14752 (N_14752,N_5211,N_9425);
nand U14753 (N_14753,N_9293,N_5869);
nand U14754 (N_14754,N_9094,N_6972);
xnor U14755 (N_14755,N_6543,N_5492);
nand U14756 (N_14756,N_8729,N_8321);
nor U14757 (N_14757,N_7425,N_7486);
nand U14758 (N_14758,N_5698,N_6519);
xnor U14759 (N_14759,N_8300,N_9128);
nor U14760 (N_14760,N_9435,N_9243);
and U14761 (N_14761,N_5548,N_8339);
or U14762 (N_14762,N_5223,N_8700);
nand U14763 (N_14763,N_7278,N_7223);
nor U14764 (N_14764,N_8418,N_7470);
xnor U14765 (N_14765,N_8711,N_9855);
and U14766 (N_14766,N_9498,N_5302);
and U14767 (N_14767,N_5800,N_6510);
nand U14768 (N_14768,N_9693,N_9848);
or U14769 (N_14769,N_9382,N_7001);
xnor U14770 (N_14770,N_9206,N_6604);
nand U14771 (N_14771,N_7688,N_5590);
or U14772 (N_14772,N_8306,N_7091);
nand U14773 (N_14773,N_5007,N_5615);
nand U14774 (N_14774,N_7122,N_6634);
or U14775 (N_14775,N_6117,N_5396);
or U14776 (N_14776,N_9043,N_7488);
nor U14777 (N_14777,N_7529,N_6723);
and U14778 (N_14778,N_9890,N_9183);
xor U14779 (N_14779,N_7360,N_9306);
nor U14780 (N_14780,N_8451,N_6530);
and U14781 (N_14781,N_8439,N_9935);
or U14782 (N_14782,N_9064,N_9391);
and U14783 (N_14783,N_5554,N_8261);
xnor U14784 (N_14784,N_7121,N_9469);
and U14785 (N_14785,N_8596,N_6787);
nand U14786 (N_14786,N_8539,N_9576);
or U14787 (N_14787,N_9196,N_6720);
and U14788 (N_14788,N_5565,N_5647);
xor U14789 (N_14789,N_8458,N_8478);
or U14790 (N_14790,N_8088,N_6415);
nor U14791 (N_14791,N_6393,N_9223);
or U14792 (N_14792,N_6343,N_6701);
nand U14793 (N_14793,N_9024,N_7001);
and U14794 (N_14794,N_9086,N_7075);
nand U14795 (N_14795,N_5399,N_8604);
nor U14796 (N_14796,N_7067,N_8551);
nand U14797 (N_14797,N_5999,N_9229);
and U14798 (N_14798,N_9789,N_6669);
xor U14799 (N_14799,N_6270,N_8321);
nand U14800 (N_14800,N_9692,N_7255);
or U14801 (N_14801,N_7566,N_8069);
or U14802 (N_14802,N_7777,N_5620);
or U14803 (N_14803,N_7632,N_8123);
or U14804 (N_14804,N_9391,N_9431);
nor U14805 (N_14805,N_5721,N_5007);
and U14806 (N_14806,N_7030,N_6356);
nor U14807 (N_14807,N_9864,N_7922);
and U14808 (N_14808,N_7183,N_6363);
or U14809 (N_14809,N_8463,N_9387);
xor U14810 (N_14810,N_9858,N_7059);
or U14811 (N_14811,N_6752,N_5085);
or U14812 (N_14812,N_7089,N_8850);
nand U14813 (N_14813,N_6551,N_8509);
and U14814 (N_14814,N_7968,N_6690);
nand U14815 (N_14815,N_7675,N_5850);
or U14816 (N_14816,N_8266,N_8160);
and U14817 (N_14817,N_9336,N_9939);
nand U14818 (N_14818,N_5404,N_9152);
or U14819 (N_14819,N_7731,N_9606);
and U14820 (N_14820,N_9768,N_5983);
nand U14821 (N_14821,N_9540,N_7951);
nand U14822 (N_14822,N_8607,N_6317);
or U14823 (N_14823,N_6522,N_5602);
and U14824 (N_14824,N_8868,N_9673);
or U14825 (N_14825,N_7614,N_7161);
nand U14826 (N_14826,N_6490,N_5283);
and U14827 (N_14827,N_6597,N_9907);
xnor U14828 (N_14828,N_6341,N_7208);
or U14829 (N_14829,N_7970,N_5735);
nor U14830 (N_14830,N_5245,N_7094);
nand U14831 (N_14831,N_5263,N_9383);
nand U14832 (N_14832,N_8153,N_9965);
nand U14833 (N_14833,N_8798,N_5387);
nand U14834 (N_14834,N_8326,N_6351);
and U14835 (N_14835,N_7299,N_5074);
and U14836 (N_14836,N_5392,N_8925);
xnor U14837 (N_14837,N_5401,N_7397);
nor U14838 (N_14838,N_5073,N_8920);
and U14839 (N_14839,N_8912,N_5756);
nor U14840 (N_14840,N_6310,N_8203);
nand U14841 (N_14841,N_5639,N_7715);
and U14842 (N_14842,N_5551,N_5176);
nand U14843 (N_14843,N_6662,N_6729);
nor U14844 (N_14844,N_9750,N_8432);
nor U14845 (N_14845,N_9857,N_5837);
xnor U14846 (N_14846,N_8245,N_9493);
xor U14847 (N_14847,N_8912,N_6794);
nor U14848 (N_14848,N_8429,N_8252);
nand U14849 (N_14849,N_5378,N_8830);
nor U14850 (N_14850,N_9777,N_9360);
and U14851 (N_14851,N_5041,N_9817);
nand U14852 (N_14852,N_7441,N_5896);
nor U14853 (N_14853,N_5166,N_9797);
nor U14854 (N_14854,N_5452,N_8507);
or U14855 (N_14855,N_5391,N_9019);
nand U14856 (N_14856,N_8951,N_6521);
nor U14857 (N_14857,N_6299,N_9250);
nand U14858 (N_14858,N_8803,N_5708);
nor U14859 (N_14859,N_5901,N_9742);
or U14860 (N_14860,N_7685,N_6573);
xnor U14861 (N_14861,N_7081,N_7366);
and U14862 (N_14862,N_8194,N_9243);
xnor U14863 (N_14863,N_8829,N_5226);
and U14864 (N_14864,N_6663,N_5387);
and U14865 (N_14865,N_9278,N_9185);
xnor U14866 (N_14866,N_7716,N_5373);
nand U14867 (N_14867,N_8899,N_9849);
and U14868 (N_14868,N_8371,N_8082);
nand U14869 (N_14869,N_6587,N_9445);
or U14870 (N_14870,N_9657,N_7384);
xor U14871 (N_14871,N_7926,N_8350);
xnor U14872 (N_14872,N_7708,N_7493);
nand U14873 (N_14873,N_5491,N_7157);
xor U14874 (N_14874,N_6119,N_5522);
and U14875 (N_14875,N_8578,N_9658);
and U14876 (N_14876,N_8424,N_6392);
or U14877 (N_14877,N_6146,N_8446);
nand U14878 (N_14878,N_5939,N_9892);
or U14879 (N_14879,N_5297,N_6413);
or U14880 (N_14880,N_6484,N_6629);
nand U14881 (N_14881,N_6967,N_9966);
and U14882 (N_14882,N_7602,N_7721);
or U14883 (N_14883,N_6070,N_8426);
xnor U14884 (N_14884,N_5223,N_8502);
nand U14885 (N_14885,N_9203,N_9089);
nor U14886 (N_14886,N_5183,N_6165);
nor U14887 (N_14887,N_6222,N_5630);
or U14888 (N_14888,N_5526,N_8522);
nor U14889 (N_14889,N_7976,N_6348);
nor U14890 (N_14890,N_5718,N_5915);
nand U14891 (N_14891,N_7175,N_8270);
or U14892 (N_14892,N_8754,N_8583);
or U14893 (N_14893,N_6354,N_6286);
nor U14894 (N_14894,N_8084,N_6055);
nor U14895 (N_14895,N_8270,N_9659);
and U14896 (N_14896,N_7737,N_7770);
nand U14897 (N_14897,N_9582,N_6248);
nand U14898 (N_14898,N_8986,N_7128);
nor U14899 (N_14899,N_7278,N_9117);
and U14900 (N_14900,N_5097,N_5201);
and U14901 (N_14901,N_7896,N_5868);
and U14902 (N_14902,N_6093,N_9082);
or U14903 (N_14903,N_8319,N_6666);
and U14904 (N_14904,N_8562,N_7656);
nor U14905 (N_14905,N_7678,N_8572);
or U14906 (N_14906,N_5132,N_8188);
and U14907 (N_14907,N_5011,N_6241);
nand U14908 (N_14908,N_9185,N_8850);
nand U14909 (N_14909,N_9827,N_5837);
or U14910 (N_14910,N_6114,N_5704);
and U14911 (N_14911,N_7014,N_9345);
nand U14912 (N_14912,N_8765,N_8062);
nor U14913 (N_14913,N_5070,N_5495);
and U14914 (N_14914,N_9348,N_6060);
nand U14915 (N_14915,N_9719,N_6354);
and U14916 (N_14916,N_7169,N_5896);
and U14917 (N_14917,N_7542,N_6768);
nand U14918 (N_14918,N_6990,N_8688);
or U14919 (N_14919,N_8900,N_8943);
nor U14920 (N_14920,N_6069,N_6414);
and U14921 (N_14921,N_7259,N_8850);
nor U14922 (N_14922,N_5643,N_7079);
or U14923 (N_14923,N_6076,N_5331);
or U14924 (N_14924,N_6622,N_8970);
nand U14925 (N_14925,N_9965,N_8964);
xnor U14926 (N_14926,N_9064,N_9177);
and U14927 (N_14927,N_6056,N_9212);
and U14928 (N_14928,N_6999,N_5147);
nor U14929 (N_14929,N_9644,N_8360);
nand U14930 (N_14930,N_8221,N_7205);
and U14931 (N_14931,N_5124,N_6041);
nor U14932 (N_14932,N_6694,N_8363);
xor U14933 (N_14933,N_5165,N_8890);
nor U14934 (N_14934,N_5201,N_6688);
nand U14935 (N_14935,N_5861,N_8287);
nand U14936 (N_14936,N_7274,N_6184);
nand U14937 (N_14937,N_8546,N_7459);
or U14938 (N_14938,N_8149,N_5798);
or U14939 (N_14939,N_8227,N_6807);
and U14940 (N_14940,N_8515,N_8351);
nand U14941 (N_14941,N_5578,N_6030);
xor U14942 (N_14942,N_9568,N_5149);
and U14943 (N_14943,N_8122,N_8022);
or U14944 (N_14944,N_8206,N_8124);
or U14945 (N_14945,N_9563,N_8392);
or U14946 (N_14946,N_8923,N_7991);
nor U14947 (N_14947,N_9630,N_7480);
nor U14948 (N_14948,N_9034,N_9629);
nand U14949 (N_14949,N_9455,N_5223);
and U14950 (N_14950,N_6140,N_5921);
xnor U14951 (N_14951,N_8169,N_5671);
or U14952 (N_14952,N_6172,N_7608);
nand U14953 (N_14953,N_8283,N_7137);
xnor U14954 (N_14954,N_5866,N_7144);
nand U14955 (N_14955,N_5786,N_9220);
nand U14956 (N_14956,N_8887,N_8728);
or U14957 (N_14957,N_6694,N_5915);
nand U14958 (N_14958,N_6433,N_9395);
and U14959 (N_14959,N_7512,N_6264);
nor U14960 (N_14960,N_7963,N_6521);
and U14961 (N_14961,N_6296,N_8952);
nand U14962 (N_14962,N_5107,N_8455);
and U14963 (N_14963,N_5917,N_9233);
or U14964 (N_14964,N_8299,N_5394);
xnor U14965 (N_14965,N_6486,N_5207);
nor U14966 (N_14966,N_8832,N_7010);
or U14967 (N_14967,N_6991,N_6234);
or U14968 (N_14968,N_6732,N_6784);
xnor U14969 (N_14969,N_6205,N_9677);
and U14970 (N_14970,N_7206,N_8195);
and U14971 (N_14971,N_8379,N_6532);
or U14972 (N_14972,N_7217,N_7130);
nand U14973 (N_14973,N_6652,N_7578);
nand U14974 (N_14974,N_5055,N_7705);
and U14975 (N_14975,N_8247,N_8846);
nor U14976 (N_14976,N_9270,N_8409);
and U14977 (N_14977,N_6557,N_7017);
nor U14978 (N_14978,N_6983,N_7267);
nand U14979 (N_14979,N_5227,N_7977);
and U14980 (N_14980,N_7288,N_6525);
and U14981 (N_14981,N_9291,N_7160);
and U14982 (N_14982,N_5427,N_9010);
or U14983 (N_14983,N_5407,N_5585);
nor U14984 (N_14984,N_8366,N_5998);
nor U14985 (N_14985,N_8270,N_5560);
nand U14986 (N_14986,N_9761,N_8685);
and U14987 (N_14987,N_8536,N_8343);
nand U14988 (N_14988,N_9124,N_8464);
and U14989 (N_14989,N_8292,N_7815);
and U14990 (N_14990,N_7867,N_8570);
and U14991 (N_14991,N_6862,N_7704);
nor U14992 (N_14992,N_9330,N_8149);
and U14993 (N_14993,N_6268,N_9026);
nor U14994 (N_14994,N_9355,N_5533);
nor U14995 (N_14995,N_7941,N_5047);
xor U14996 (N_14996,N_8656,N_6250);
nand U14997 (N_14997,N_9507,N_7218);
or U14998 (N_14998,N_9219,N_6374);
nor U14999 (N_14999,N_7026,N_5446);
xor UO_0 (O_0,N_12519,N_14206);
nand UO_1 (O_1,N_11805,N_11741);
and UO_2 (O_2,N_12080,N_13611);
xnor UO_3 (O_3,N_10428,N_14867);
nor UO_4 (O_4,N_14574,N_12283);
nor UO_5 (O_5,N_11573,N_11197);
or UO_6 (O_6,N_10998,N_12290);
nor UO_7 (O_7,N_12030,N_13376);
nor UO_8 (O_8,N_14579,N_12661);
and UO_9 (O_9,N_12565,N_14092);
or UO_10 (O_10,N_10129,N_11541);
and UO_11 (O_11,N_12880,N_12557);
or UO_12 (O_12,N_11790,N_14042);
nor UO_13 (O_13,N_10850,N_12141);
xor UO_14 (O_14,N_11222,N_11376);
or UO_15 (O_15,N_12922,N_11331);
or UO_16 (O_16,N_14685,N_13014);
or UO_17 (O_17,N_14837,N_10705);
and UO_18 (O_18,N_14032,N_10501);
nand UO_19 (O_19,N_10945,N_11780);
and UO_20 (O_20,N_10314,N_12125);
nand UO_21 (O_21,N_14910,N_13832);
or UO_22 (O_22,N_14664,N_14834);
nand UO_23 (O_23,N_10874,N_14791);
nor UO_24 (O_24,N_13406,N_11430);
nor UO_25 (O_25,N_10577,N_14940);
and UO_26 (O_26,N_12464,N_14635);
and UO_27 (O_27,N_13175,N_14045);
or UO_28 (O_28,N_10287,N_10980);
or UO_29 (O_29,N_14737,N_11891);
nor UO_30 (O_30,N_13689,N_12605);
nand UO_31 (O_31,N_10585,N_13395);
or UO_32 (O_32,N_10591,N_13384);
nor UO_33 (O_33,N_14824,N_13531);
and UO_34 (O_34,N_11545,N_11426);
or UO_35 (O_35,N_12157,N_13559);
and UO_36 (O_36,N_14238,N_12222);
nand UO_37 (O_37,N_14479,N_11909);
and UO_38 (O_38,N_12311,N_11188);
and UO_39 (O_39,N_13577,N_13150);
nor UO_40 (O_40,N_10515,N_14217);
nor UO_41 (O_41,N_12475,N_14708);
xor UO_42 (O_42,N_13479,N_12753);
nand UO_43 (O_43,N_14854,N_14457);
nand UO_44 (O_44,N_13124,N_10159);
and UO_45 (O_45,N_12574,N_10711);
nor UO_46 (O_46,N_14922,N_10059);
nor UO_47 (O_47,N_10066,N_10824);
nor UO_48 (O_48,N_13498,N_11184);
nand UO_49 (O_49,N_13623,N_13226);
xor UO_50 (O_50,N_14117,N_13591);
or UO_51 (O_51,N_14591,N_11735);
xnor UO_52 (O_52,N_14857,N_14973);
and UO_53 (O_53,N_14272,N_13888);
nor UO_54 (O_54,N_13523,N_14802);
nand UO_55 (O_55,N_11215,N_10975);
nand UO_56 (O_56,N_12213,N_14723);
or UO_57 (O_57,N_12429,N_14220);
or UO_58 (O_58,N_14616,N_14356);
or UO_59 (O_59,N_14269,N_14843);
nor UO_60 (O_60,N_10497,N_12214);
or UO_61 (O_61,N_11610,N_14602);
and UO_62 (O_62,N_14765,N_12749);
nand UO_63 (O_63,N_13590,N_11076);
and UO_64 (O_64,N_14986,N_11913);
nand UO_65 (O_65,N_13461,N_13847);
nor UO_66 (O_66,N_12722,N_14548);
or UO_67 (O_67,N_11239,N_14582);
nand UO_68 (O_68,N_12850,N_10897);
and UO_69 (O_69,N_12020,N_14241);
or UO_70 (O_70,N_10036,N_12910);
nor UO_71 (O_71,N_10598,N_13836);
and UO_72 (O_72,N_12669,N_11703);
nor UO_73 (O_73,N_11737,N_13251);
and UO_74 (O_74,N_12066,N_10098);
nand UO_75 (O_75,N_12160,N_12510);
and UO_76 (O_76,N_12422,N_13002);
nand UO_77 (O_77,N_10388,N_13549);
xor UO_78 (O_78,N_10793,N_10871);
or UO_79 (O_79,N_13660,N_12024);
or UO_80 (O_80,N_10640,N_11846);
nor UO_81 (O_81,N_13131,N_11067);
nor UO_82 (O_82,N_13451,N_14360);
nand UO_83 (O_83,N_10589,N_13919);
nor UO_84 (O_84,N_14514,N_12779);
or UO_85 (O_85,N_11186,N_12412);
nor UO_86 (O_86,N_14482,N_14641);
or UO_87 (O_87,N_13053,N_13626);
nor UO_88 (O_88,N_12645,N_11098);
and UO_89 (O_89,N_14619,N_11924);
xor UO_90 (O_90,N_10986,N_14778);
nand UO_91 (O_91,N_10113,N_12360);
or UO_92 (O_92,N_14759,N_14415);
or UO_93 (O_93,N_12576,N_13264);
nor UO_94 (O_94,N_14433,N_10649);
or UO_95 (O_95,N_11662,N_13991);
or UO_96 (O_96,N_10639,N_12727);
nand UO_97 (O_97,N_13229,N_11264);
and UO_98 (O_98,N_12294,N_14148);
xnor UO_99 (O_99,N_14449,N_11890);
or UO_100 (O_100,N_10456,N_10333);
xnor UO_101 (O_101,N_12695,N_11212);
or UO_102 (O_102,N_12385,N_11588);
nor UO_103 (O_103,N_14210,N_12054);
nand UO_104 (O_104,N_12707,N_14028);
or UO_105 (O_105,N_11893,N_13690);
nor UO_106 (O_106,N_13650,N_14448);
or UO_107 (O_107,N_13501,N_12419);
and UO_108 (O_108,N_10034,N_12365);
nor UO_109 (O_109,N_10226,N_14104);
and UO_110 (O_110,N_11260,N_14462);
nor UO_111 (O_111,N_10909,N_12920);
and UO_112 (O_112,N_13331,N_11606);
nand UO_113 (O_113,N_10527,N_13496);
or UO_114 (O_114,N_12699,N_11395);
and UO_115 (O_115,N_13894,N_14311);
nor UO_116 (O_116,N_14048,N_14819);
xor UO_117 (O_117,N_13716,N_11285);
nand UO_118 (O_118,N_13587,N_14652);
or UO_119 (O_119,N_11847,N_11629);
nand UO_120 (O_120,N_11486,N_13058);
nor UO_121 (O_121,N_14866,N_10142);
nand UO_122 (O_122,N_13080,N_13973);
nand UO_123 (O_123,N_12937,N_14534);
or UO_124 (O_124,N_12599,N_10804);
nor UO_125 (O_125,N_11991,N_11992);
nor UO_126 (O_126,N_12352,N_11295);
nor UO_127 (O_127,N_10387,N_12562);
nor UO_128 (O_128,N_10817,N_12447);
nand UO_129 (O_129,N_13333,N_14649);
nand UO_130 (O_130,N_12381,N_11999);
and UO_131 (O_131,N_10115,N_12697);
nor UO_132 (O_132,N_12162,N_10016);
xnor UO_133 (O_133,N_10475,N_13319);
or UO_134 (O_134,N_11088,N_13774);
nand UO_135 (O_135,N_12050,N_14670);
and UO_136 (O_136,N_11551,N_14453);
or UO_137 (O_137,N_10143,N_13318);
nor UO_138 (O_138,N_14851,N_12477);
or UO_139 (O_139,N_14389,N_10813);
nand UO_140 (O_140,N_14103,N_14036);
and UO_141 (O_141,N_13492,N_10123);
or UO_142 (O_142,N_11613,N_14746);
nand UO_143 (O_143,N_13624,N_13541);
nor UO_144 (O_144,N_12793,N_13134);
nor UO_145 (O_145,N_11571,N_12698);
and UO_146 (O_146,N_10770,N_14056);
nand UO_147 (O_147,N_14853,N_10434);
nor UO_148 (O_148,N_12855,N_14501);
and UO_149 (O_149,N_11500,N_10555);
or UO_150 (O_150,N_13108,N_11174);
and UO_151 (O_151,N_12396,N_10575);
and UO_152 (O_152,N_14455,N_14595);
nor UO_153 (O_153,N_14142,N_11172);
nand UO_154 (O_154,N_12487,N_12692);
or UO_155 (O_155,N_13816,N_13109);
nand UO_156 (O_156,N_11785,N_12232);
and UO_157 (O_157,N_14067,N_14143);
or UO_158 (O_158,N_12187,N_14964);
nor UO_159 (O_159,N_14275,N_10661);
nand UO_160 (O_160,N_14307,N_11346);
or UO_161 (O_161,N_14370,N_14601);
nand UO_162 (O_162,N_13420,N_13332);
and UO_163 (O_163,N_14733,N_13462);
nor UO_164 (O_164,N_14088,N_11363);
and UO_165 (O_165,N_10329,N_10199);
nand UO_166 (O_166,N_13314,N_11866);
or UO_167 (O_167,N_14810,N_14406);
and UO_168 (O_168,N_11114,N_11825);
xnor UO_169 (O_169,N_10603,N_12279);
nor UO_170 (O_170,N_10863,N_14956);
and UO_171 (O_171,N_11634,N_14618);
nor UO_172 (O_172,N_12632,N_11600);
nand UO_173 (O_173,N_10091,N_10438);
nand UO_174 (O_174,N_13830,N_10706);
xor UO_175 (O_175,N_14700,N_11727);
nand UO_176 (O_176,N_10315,N_10522);
xor UO_177 (O_177,N_12830,N_14299);
or UO_178 (O_178,N_10245,N_11607);
nand UO_179 (O_179,N_12949,N_11468);
nor UO_180 (O_180,N_14296,N_13633);
or UO_181 (O_181,N_10297,N_10222);
or UO_182 (O_182,N_14913,N_13557);
nand UO_183 (O_183,N_11210,N_11747);
or UO_184 (O_184,N_12056,N_14876);
nor UO_185 (O_185,N_10203,N_10959);
nor UO_186 (O_186,N_13714,N_12603);
nand UO_187 (O_187,N_14536,N_10030);
or UO_188 (O_188,N_14014,N_12478);
nand UO_189 (O_189,N_14914,N_13979);
and UO_190 (O_190,N_11681,N_10787);
or UO_191 (O_191,N_12837,N_13750);
xor UO_192 (O_192,N_12355,N_11489);
or UO_193 (O_193,N_13011,N_13293);
and UO_194 (O_194,N_12517,N_12821);
nor UO_195 (O_195,N_11935,N_11522);
nor UO_196 (O_196,N_13339,N_12264);
or UO_197 (O_197,N_10043,N_11742);
or UO_198 (O_198,N_14147,N_13683);
nand UO_199 (O_199,N_14283,N_10925);
and UO_200 (O_200,N_10865,N_10570);
or UO_201 (O_201,N_12914,N_11147);
or UO_202 (O_202,N_12458,N_14306);
nand UO_203 (O_203,N_10478,N_14197);
nor UO_204 (O_204,N_10678,N_11560);
or UO_205 (O_205,N_12975,N_11989);
xor UO_206 (O_206,N_10077,N_14101);
nor UO_207 (O_207,N_14471,N_14425);
nand UO_208 (O_208,N_10581,N_11388);
and UO_209 (O_209,N_13940,N_14183);
nand UO_210 (O_210,N_14812,N_10557);
or UO_211 (O_211,N_11936,N_12220);
nor UO_212 (O_212,N_10085,N_13394);
nand UO_213 (O_213,N_12659,N_13146);
nor UO_214 (O_214,N_12223,N_10768);
and UO_215 (O_215,N_10718,N_13405);
and UO_216 (O_216,N_12567,N_12465);
xnor UO_217 (O_217,N_13929,N_11862);
nand UO_218 (O_218,N_11422,N_13110);
and UO_219 (O_219,N_12463,N_10453);
nand UO_220 (O_220,N_12498,N_13643);
nand UO_221 (O_221,N_12641,N_11765);
xor UO_222 (O_222,N_14452,N_11365);
nand UO_223 (O_223,N_12990,N_10331);
and UO_224 (O_224,N_10141,N_12179);
and UO_225 (O_225,N_14862,N_10647);
or UO_226 (O_226,N_13439,N_14312);
and UO_227 (O_227,N_14571,N_14083);
and UO_228 (O_228,N_10014,N_10671);
or UO_229 (O_229,N_13342,N_13117);
or UO_230 (O_230,N_12849,N_14015);
and UO_231 (O_231,N_10134,N_14253);
nand UO_232 (O_232,N_12243,N_11589);
and UO_233 (O_233,N_12732,N_11550);
xor UO_234 (O_234,N_14458,N_13598);
nor UO_235 (O_235,N_11865,N_12008);
xor UO_236 (O_236,N_10426,N_10336);
nor UO_237 (O_237,N_12958,N_11046);
and UO_238 (O_238,N_11763,N_14764);
nand UO_239 (O_239,N_14881,N_12560);
nor UO_240 (O_240,N_13572,N_13355);
nor UO_241 (O_241,N_11996,N_14889);
and UO_242 (O_242,N_14123,N_10357);
nor UO_243 (O_243,N_12048,N_11964);
nand UO_244 (O_244,N_11042,N_14232);
or UO_245 (O_245,N_12773,N_11837);
and UO_246 (O_246,N_10324,N_12272);
and UO_247 (O_247,N_10551,N_13688);
and UO_248 (O_248,N_14125,N_12114);
and UO_249 (O_249,N_10814,N_10481);
nor UO_250 (O_250,N_12600,N_13540);
or UO_251 (O_251,N_11575,N_12948);
nand UO_252 (O_252,N_13675,N_12065);
nand UO_253 (O_253,N_12173,N_14599);
nand UO_254 (O_254,N_12897,N_12282);
xnor UO_255 (O_255,N_14727,N_13207);
xor UO_256 (O_256,N_12084,N_10025);
nand UO_257 (O_257,N_13198,N_13310);
nand UO_258 (O_258,N_13133,N_14419);
nor UO_259 (O_259,N_13760,N_13773);
xor UO_260 (O_260,N_10547,N_14520);
or UO_261 (O_261,N_14613,N_13844);
nand UO_262 (O_262,N_13083,N_14392);
or UO_263 (O_263,N_11353,N_13087);
xnor UO_264 (O_264,N_11436,N_10473);
and UO_265 (O_265,N_11157,N_12312);
and UO_266 (O_266,N_11040,N_13842);
nand UO_267 (O_267,N_12268,N_10356);
xor UO_268 (O_268,N_14758,N_10617);
and UO_269 (O_269,N_12684,N_10961);
or UO_270 (O_270,N_10274,N_13041);
and UO_271 (O_271,N_11033,N_12266);
or UO_272 (O_272,N_10485,N_12893);
nor UO_273 (O_273,N_11087,N_11848);
and UO_274 (O_274,N_12186,N_12941);
nor UO_275 (O_275,N_10634,N_14258);
and UO_276 (O_276,N_12476,N_14276);
nor UO_277 (O_277,N_13486,N_14584);
nor UO_278 (O_278,N_12806,N_11107);
or UO_279 (O_279,N_14378,N_10566);
nand UO_280 (O_280,N_13596,N_10916);
and UO_281 (O_281,N_14545,N_14355);
xnor UO_282 (O_282,N_13446,N_14978);
and UO_283 (O_283,N_12170,N_11746);
and UO_284 (O_284,N_11757,N_13050);
nand UO_285 (O_285,N_11858,N_11685);
nand UO_286 (O_286,N_14712,N_14081);
xor UO_287 (O_287,N_11798,N_12159);
nor UO_288 (O_288,N_12131,N_10496);
nor UO_289 (O_289,N_14608,N_10687);
or UO_290 (O_290,N_11927,N_13694);
nand UO_291 (O_291,N_12852,N_14057);
or UO_292 (O_292,N_13076,N_10120);
or UO_293 (O_293,N_12354,N_10796);
or UO_294 (O_294,N_11292,N_11901);
nand UO_295 (O_295,N_13222,N_11962);
xnor UO_296 (O_296,N_13582,N_11656);
nand UO_297 (O_297,N_10312,N_10751);
xnor UO_298 (O_298,N_11884,N_10786);
and UO_299 (O_299,N_12053,N_13506);
nand UO_300 (O_300,N_14351,N_11908);
nand UO_301 (O_301,N_11017,N_12956);
and UO_302 (O_302,N_11438,N_10472);
or UO_303 (O_303,N_10450,N_14397);
and UO_304 (O_304,N_13491,N_11041);
nand UO_305 (O_305,N_11649,N_10499);
nand UO_306 (O_306,N_11066,N_11739);
or UO_307 (O_307,N_12531,N_10645);
nor UO_308 (O_308,N_13114,N_14215);
xor UO_309 (O_309,N_14776,N_14063);
nand UO_310 (O_310,N_14807,N_14456);
xor UO_311 (O_311,N_11193,N_10258);
or UO_312 (O_312,N_11048,N_12198);
and UO_313 (O_313,N_10266,N_11849);
nor UO_314 (O_314,N_11441,N_11294);
and UO_315 (O_315,N_11071,N_10346);
or UO_316 (O_316,N_12110,N_14991);
or UO_317 (O_317,N_10212,N_14981);
nand UO_318 (O_318,N_11064,N_11319);
or UO_319 (O_319,N_11933,N_12529);
nand UO_320 (O_320,N_11444,N_13959);
and UO_321 (O_321,N_14633,N_13353);
or UO_322 (O_322,N_12480,N_12960);
nand UO_323 (O_323,N_14838,N_14836);
nand UO_324 (O_324,N_10549,N_10702);
or UO_325 (O_325,N_12548,N_12321);
or UO_326 (O_326,N_14491,N_12143);
and UO_327 (O_327,N_10621,N_14129);
nor UO_328 (O_328,N_13885,N_10064);
nor UO_329 (O_329,N_10174,N_13920);
nor UO_330 (O_330,N_12535,N_14346);
nor UO_331 (O_331,N_12763,N_12289);
xor UO_332 (O_332,N_12474,N_13326);
or UO_333 (O_333,N_13543,N_14199);
or UO_334 (O_334,N_12023,N_11715);
nor UO_335 (O_335,N_14974,N_13911);
nand UO_336 (O_336,N_13519,N_14407);
xnor UO_337 (O_337,N_12402,N_12655);
xnor UO_338 (O_338,N_13008,N_11281);
nand UO_339 (O_339,N_11756,N_10592);
xnor UO_340 (O_340,N_14839,N_13316);
and UO_341 (O_341,N_11667,N_13909);
and UO_342 (O_342,N_11868,N_12998);
and UO_343 (O_343,N_10761,N_10410);
nand UO_344 (O_344,N_13240,N_11330);
nor UO_345 (O_345,N_13980,N_12930);
nor UO_346 (O_346,N_14598,N_14752);
nand UO_347 (O_347,N_10765,N_14200);
or UO_348 (O_348,N_10139,N_13669);
xnor UO_349 (O_349,N_14895,N_13585);
nor UO_350 (O_350,N_11787,N_14177);
and UO_351 (O_351,N_13465,N_13672);
nor UO_352 (O_352,N_13667,N_13530);
xor UO_353 (O_353,N_10891,N_13195);
and UO_354 (O_354,N_12060,N_11855);
nor UO_355 (O_355,N_12137,N_14451);
or UO_356 (O_356,N_13105,N_12524);
nand UO_357 (O_357,N_13219,N_14364);
xor UO_358 (O_358,N_14716,N_10658);
xor UO_359 (O_359,N_11897,N_12123);
or UO_360 (O_360,N_11484,N_13184);
and UO_361 (O_361,N_11795,N_11100);
nand UO_362 (O_362,N_11604,N_14628);
nor UO_363 (O_363,N_12401,N_11085);
nor UO_364 (O_364,N_14093,N_10225);
nand UO_365 (O_365,N_10738,N_14988);
or UO_366 (O_366,N_10444,N_11978);
nor UO_367 (O_367,N_10597,N_13261);
or UO_368 (O_368,N_12586,N_10827);
nor UO_369 (O_369,N_11204,N_14025);
nand UO_370 (O_370,N_10483,N_11333);
nor UO_371 (O_371,N_10951,N_13796);
nor UO_372 (O_372,N_12261,N_10146);
and UO_373 (O_373,N_12759,N_12151);
nor UO_374 (O_374,N_12967,N_13655);
xor UO_375 (O_375,N_13098,N_10633);
or UO_376 (O_376,N_10525,N_13101);
or UO_377 (O_377,N_14636,N_11410);
or UO_378 (O_378,N_12391,N_10966);
nor UO_379 (O_379,N_13415,N_13306);
nor UO_380 (O_380,N_12484,N_13256);
xnor UO_381 (O_381,N_10180,N_10970);
or UO_382 (O_382,N_11515,N_11934);
and UO_383 (O_383,N_11128,N_13234);
or UO_384 (O_384,N_11655,N_11099);
and UO_385 (O_385,N_13097,N_12751);
and UO_386 (O_386,N_13554,N_14698);
nor UO_387 (O_387,N_12523,N_14787);
and UO_388 (O_388,N_14040,N_11517);
nand UO_389 (O_389,N_12057,N_10112);
nor UO_390 (O_390,N_14745,N_12974);
and UO_391 (O_391,N_12424,N_14750);
nor UO_392 (O_392,N_14905,N_11002);
nor UO_393 (O_393,N_14097,N_13983);
nand UO_394 (O_394,N_12052,N_14322);
nor UO_395 (O_395,N_14376,N_13410);
nand UO_396 (O_396,N_13283,N_10283);
and UO_397 (O_397,N_12456,N_12988);
nor UO_398 (O_398,N_13346,N_10624);
nand UO_399 (O_399,N_10904,N_10715);
and UO_400 (O_400,N_14717,N_12711);
or UO_401 (O_401,N_10936,N_13879);
nand UO_402 (O_402,N_13236,N_11643);
nand UO_403 (O_403,N_12296,N_10248);
nand UO_404 (O_404,N_14893,N_11697);
or UO_405 (O_405,N_11078,N_13154);
nor UO_406 (O_406,N_14151,N_10477);
and UO_407 (O_407,N_12269,N_12769);
or UO_408 (O_408,N_14185,N_13200);
and UO_409 (O_409,N_13536,N_14263);
or UO_410 (O_410,N_14417,N_10504);
nor UO_411 (O_411,N_13452,N_14180);
or UO_412 (O_412,N_11421,N_11888);
nor UO_413 (O_413,N_10806,N_11531);
and UO_414 (O_414,N_13791,N_12746);
or UO_415 (O_415,N_12251,N_12202);
nand UO_416 (O_416,N_12657,N_14512);
nor UO_417 (O_417,N_13875,N_11902);
or UO_418 (O_418,N_13471,N_10582);
or UO_419 (O_419,N_11984,N_12395);
nand UO_420 (O_420,N_11959,N_13330);
nor UO_421 (O_421,N_14943,N_12128);
or UO_422 (O_422,N_10632,N_13814);
nand UO_423 (O_423,N_13642,N_11428);
nor UO_424 (O_424,N_11781,N_12446);
or UO_425 (O_425,N_10535,N_14509);
or UO_426 (O_426,N_11401,N_12511);
and UO_427 (O_427,N_12549,N_13381);
nor UO_428 (O_428,N_13629,N_11635);
or UO_429 (O_429,N_14367,N_13951);
and UO_430 (O_430,N_13317,N_11065);
or UO_431 (O_431,N_12227,N_11458);
xnor UO_432 (O_432,N_12579,N_11886);
nor UO_433 (O_433,N_10458,N_14437);
nor UO_434 (O_434,N_12298,N_10474);
nor UO_435 (O_435,N_12813,N_10752);
or UO_436 (O_436,N_14987,N_14577);
or UO_437 (O_437,N_14050,N_10107);
nor UO_438 (O_438,N_11730,N_13102);
nor UO_439 (O_439,N_11030,N_14314);
or UO_440 (O_440,N_13499,N_14373);
and UO_441 (O_441,N_10612,N_12278);
xnor UO_442 (O_442,N_10580,N_10693);
xor UO_443 (O_443,N_12415,N_11835);
or UO_444 (O_444,N_11381,N_10003);
nor UO_445 (O_445,N_10486,N_12113);
nand UO_446 (O_446,N_11247,N_11833);
nor UO_447 (O_447,N_13432,N_13328);
nor UO_448 (O_448,N_12775,N_10719);
nand UO_449 (O_449,N_13977,N_12546);
nand UO_450 (O_450,N_10057,N_11325);
and UO_451 (O_451,N_11615,N_12715);
and UO_452 (O_452,N_11993,N_11297);
nand UO_453 (O_453,N_10267,N_11016);
or UO_454 (O_454,N_13387,N_12488);
or UO_455 (O_455,N_13091,N_14879);
and UO_456 (O_456,N_12393,N_10625);
and UO_457 (O_457,N_12106,N_10399);
and UO_458 (O_458,N_10655,N_10000);
or UO_459 (O_459,N_12903,N_12687);
nor UO_460 (O_460,N_10783,N_10701);
nand UO_461 (O_461,N_11267,N_14580);
and UO_462 (O_462,N_13854,N_14609);
and UO_463 (O_463,N_13607,N_13368);
or UO_464 (O_464,N_12260,N_11856);
nand UO_465 (O_465,N_13696,N_13848);
nor UO_466 (O_466,N_10048,N_14494);
xnor UO_467 (O_467,N_11622,N_11268);
nor UO_468 (O_468,N_14975,N_11774);
nor UO_469 (O_469,N_11692,N_12445);
nand UO_470 (O_470,N_13925,N_14607);
or UO_471 (O_471,N_13225,N_14855);
nor UO_472 (O_472,N_11973,N_11129);
or UO_473 (O_473,N_14679,N_12330);
nor UO_474 (O_474,N_13803,N_11125);
nor UO_475 (O_475,N_10099,N_12189);
and UO_476 (O_476,N_14701,N_12224);
nor UO_477 (O_477,N_11338,N_14153);
nand UO_478 (O_478,N_12758,N_14310);
and UO_479 (O_479,N_14684,N_10389);
and UO_480 (O_480,N_11861,N_12558);
nor UO_481 (O_481,N_13952,N_13600);
and UO_482 (O_482,N_11802,N_13282);
nor UO_483 (O_483,N_11312,N_14768);
nor UO_484 (O_484,N_12590,N_12399);
nand UO_485 (O_485,N_11488,N_10564);
nand UO_486 (O_486,N_10449,N_10455);
or UO_487 (O_487,N_11412,N_11561);
xor UO_488 (O_488,N_10251,N_12537);
nand UO_489 (O_489,N_11683,N_10548);
nand UO_490 (O_490,N_13833,N_13341);
nand UO_491 (O_491,N_13826,N_11369);
nand UO_492 (O_492,N_10332,N_14037);
xor UO_493 (O_493,N_14486,N_13456);
xor UO_494 (O_494,N_13678,N_10921);
or UO_495 (O_495,N_10166,N_12468);
and UO_496 (O_496,N_14247,N_13325);
nor UO_497 (O_497,N_11714,N_10619);
nand UO_498 (O_498,N_11710,N_13377);
nand UO_499 (O_499,N_13687,N_14444);
nand UO_500 (O_500,N_14076,N_13403);
nor UO_501 (O_501,N_14762,N_11340);
and UO_502 (O_502,N_10923,N_14557);
nor UO_503 (O_503,N_11439,N_13950);
and UO_504 (O_504,N_12622,N_10821);
nand UO_505 (O_505,N_12504,N_11852);
nand UO_506 (O_506,N_11648,N_11138);
and UO_507 (O_507,N_10208,N_12146);
xor UO_508 (O_508,N_12000,N_14096);
nor UO_509 (O_509,N_10561,N_11496);
and UO_510 (O_510,N_14693,N_13637);
and UO_511 (O_511,N_12863,N_14469);
and UO_512 (O_512,N_12947,N_14632);
or UO_513 (O_513,N_13015,N_14046);
or UO_514 (O_514,N_14049,N_14022);
xor UO_515 (O_515,N_10156,N_14979);
nor UO_516 (O_516,N_12373,N_13709);
nand UO_517 (O_517,N_12884,N_14128);
nand UO_518 (O_518,N_11497,N_12273);
nand UO_519 (O_519,N_12101,N_10102);
or UO_520 (O_520,N_11905,N_10150);
nand UO_521 (O_521,N_10650,N_14436);
xor UO_522 (O_522,N_12790,N_14647);
or UO_523 (O_523,N_11972,N_14902);
xor UO_524 (O_524,N_12262,N_12240);
nor UO_525 (O_525,N_10100,N_12072);
and UO_526 (O_526,N_11969,N_12149);
nor UO_527 (O_527,N_13770,N_13776);
nor UO_528 (O_528,N_10778,N_12877);
nand UO_529 (O_529,N_14588,N_13740);
nand UO_530 (O_530,N_12772,N_13211);
nor UO_531 (O_531,N_12428,N_10311);
and UO_532 (O_532,N_13505,N_14439);
and UO_533 (O_533,N_12492,N_12069);
or UO_534 (O_534,N_14506,N_13388);
nor UO_535 (O_535,N_12230,N_11045);
nor UO_536 (O_536,N_12843,N_11269);
xor UO_537 (O_537,N_14427,N_13069);
nand UO_538 (O_538,N_14401,N_14657);
and UO_539 (O_539,N_12677,N_10464);
or UO_540 (O_540,N_13663,N_11022);
and UO_541 (O_541,N_14773,N_13923);
or UO_542 (O_542,N_14581,N_14907);
nor UO_543 (O_543,N_13955,N_12915);
nor UO_544 (O_544,N_14541,N_11451);
nand UO_545 (O_545,N_14138,N_12135);
and UO_546 (O_546,N_13168,N_10378);
nand UO_547 (O_547,N_13065,N_14721);
xnor UO_548 (O_548,N_14655,N_14438);
nand UO_549 (O_549,N_14250,N_11413);
nor UO_550 (O_550,N_12566,N_10668);
or UO_551 (O_551,N_10939,N_13547);
xnor UO_552 (O_552,N_10031,N_10913);
nand UO_553 (O_553,N_13799,N_11366);
or UO_554 (O_554,N_12862,N_14236);
nor UO_555 (O_555,N_14511,N_12994);
or UO_556 (O_556,N_12380,N_10361);
nand UO_557 (O_557,N_12770,N_12502);
nor UO_558 (O_558,N_12314,N_13527);
and UO_559 (O_559,N_10869,N_13907);
and UO_560 (O_560,N_14174,N_13370);
or UO_561 (O_561,N_10732,N_12658);
nor UO_562 (O_562,N_11359,N_10067);
and UO_563 (O_563,N_13526,N_11361);
nand UO_564 (O_564,N_13253,N_13771);
nor UO_565 (O_565,N_13174,N_12723);
nand UO_566 (O_566,N_10771,N_13797);
and UO_567 (O_567,N_10177,N_14445);
and UO_568 (O_568,N_13427,N_13731);
nor UO_569 (O_569,N_12271,N_11102);
and UO_570 (O_570,N_10151,N_12774);
and UO_571 (O_571,N_11814,N_10739);
and UO_572 (O_572,N_10119,N_12088);
nor UO_573 (O_573,N_12095,N_11068);
and UO_574 (O_574,N_10679,N_14399);
xor UO_575 (O_575,N_12129,N_14001);
xor UO_576 (O_576,N_12670,N_13373);
nand UO_577 (O_577,N_10853,N_10197);
or UO_578 (O_578,N_10981,N_13137);
nor UO_579 (O_579,N_11457,N_11404);
and UO_580 (O_580,N_14969,N_12741);
or UO_581 (O_581,N_10073,N_10153);
or UO_582 (O_582,N_14245,N_13654);
nor UO_583 (O_583,N_11548,N_12085);
nor UO_584 (O_584,N_10819,N_14784);
nor UO_585 (O_585,N_12828,N_10988);
xor UO_586 (O_586,N_10345,N_12865);
or UO_587 (O_587,N_10341,N_12582);
nor UO_588 (O_588,N_10364,N_10321);
nand UO_589 (O_589,N_14919,N_13963);
or UO_590 (O_590,N_12700,N_11841);
nor UO_591 (O_591,N_12580,N_13913);
nand UO_592 (O_592,N_10089,N_14996);
nor UO_593 (O_593,N_11974,N_11539);
xor UO_594 (O_594,N_12545,N_10875);
and UO_595 (O_595,N_14980,N_10012);
or UO_596 (O_596,N_13473,N_11305);
nand UO_597 (O_597,N_14167,N_12568);
xnor UO_598 (O_598,N_13412,N_12924);
nand UO_599 (O_599,N_13735,N_11673);
xnor UO_600 (O_600,N_12018,N_10210);
nor UO_601 (O_601,N_11598,N_12652);
nand UO_602 (O_602,N_13827,N_12842);
nor UO_603 (O_603,N_10293,N_14216);
nor UO_604 (O_604,N_10131,N_11318);
nor UO_605 (O_605,N_14198,N_13685);
and UO_606 (O_606,N_14377,N_13573);
nor UO_607 (O_607,N_10673,N_10529);
and UO_608 (O_608,N_11465,N_12839);
nor UO_609 (O_609,N_14883,N_14144);
nor UO_610 (O_610,N_14626,N_11680);
nand UO_611 (O_611,N_10035,N_10278);
or UO_612 (O_612,N_11243,N_10187);
or UO_613 (O_613,N_11750,N_14549);
or UO_614 (O_614,N_11518,N_12191);
and UO_615 (O_615,N_11083,N_11047);
and UO_616 (O_616,N_13005,N_10638);
and UO_617 (O_617,N_10855,N_10382);
nand UO_618 (O_618,N_10753,N_14603);
or UO_619 (O_619,N_10613,N_11585);
or UO_620 (O_620,N_13246,N_14877);
nor UO_621 (O_621,N_10275,N_14977);
and UO_622 (O_622,N_14179,N_13389);
or UO_623 (O_623,N_13233,N_14428);
nor UO_624 (O_624,N_13202,N_11594);
nor UO_625 (O_625,N_11552,N_12804);
nor UO_626 (O_626,N_12226,N_13761);
nand UO_627 (O_627,N_10710,N_13495);
nor UO_628 (O_628,N_11981,N_10838);
nand UO_629 (O_629,N_14463,N_14966);
xor UO_630 (O_630,N_11475,N_11175);
and UO_631 (O_631,N_10263,N_14869);
nor UO_632 (O_632,N_10993,N_13841);
or UO_633 (O_633,N_13104,N_12001);
or UO_634 (O_634,N_13484,N_13764);
or UO_635 (O_635,N_14669,N_12680);
and UO_636 (O_636,N_12740,N_10046);
nor UO_637 (O_637,N_11171,N_10637);
and UO_638 (O_638,N_12696,N_13897);
and UO_639 (O_639,N_14753,N_10895);
or UO_640 (O_640,N_12210,N_12507);
nor UO_641 (O_641,N_13088,N_13166);
xnor UO_642 (O_642,N_14543,N_11836);
nor UO_643 (O_643,N_10670,N_13135);
and UO_644 (O_644,N_14324,N_10754);
nand UO_645 (O_645,N_12121,N_14694);
or UO_646 (O_646,N_11554,N_13859);
nand UO_647 (O_647,N_12503,N_11156);
and UO_648 (O_648,N_10465,N_12148);
or UO_649 (O_649,N_14208,N_12506);
nor UO_650 (O_650,N_12882,N_13932);
and UO_651 (O_651,N_10708,N_14064);
nor UO_652 (O_652,N_14523,N_12551);
or UO_653 (O_653,N_13784,N_12055);
nand UO_654 (O_654,N_14010,N_10491);
nand UO_655 (O_655,N_10976,N_11699);
xnor UO_656 (O_656,N_12666,N_13849);
or UO_657 (O_657,N_12336,N_14783);
or UO_658 (O_658,N_14842,N_12703);
xor UO_659 (O_659,N_10096,N_10365);
xnor UO_660 (O_660,N_11160,N_11568);
xnor UO_661 (O_661,N_10833,N_14754);
and UO_662 (O_662,N_14440,N_10894);
or UO_663 (O_663,N_12377,N_14012);
xnor UO_664 (O_664,N_11957,N_14017);
and UO_665 (O_665,N_13197,N_10353);
nand UO_666 (O_666,N_11482,N_14478);
nand UO_667 (O_667,N_10234,N_11657);
nor UO_668 (O_668,N_12342,N_14219);
xnor UO_669 (O_669,N_11944,N_13752);
xor UO_670 (O_670,N_11339,N_11379);
and UO_671 (O_671,N_14505,N_14435);
and UO_672 (O_672,N_13812,N_13865);
and UO_673 (O_673,N_10513,N_14375);
and UO_674 (O_674,N_12649,N_14426);
nand UO_675 (O_675,N_10273,N_12120);
nor UO_676 (O_676,N_12397,N_12177);
or UO_677 (O_677,N_11131,N_11664);
nor UO_678 (O_678,N_12891,N_12675);
or UO_679 (O_679,N_12901,N_13901);
and UO_680 (O_680,N_13220,N_13867);
or UO_681 (O_681,N_14942,N_14186);
nand UO_682 (O_682,N_11010,N_10126);
or UO_683 (O_683,N_11504,N_11498);
xnor UO_684 (O_684,N_11940,N_11954);
nand UO_685 (O_685,N_10733,N_11581);
nor UO_686 (O_686,N_11789,N_14099);
or UO_687 (O_687,N_13575,N_14795);
and UO_688 (O_688,N_11006,N_12313);
xor UO_689 (O_689,N_10683,N_13986);
or UO_690 (O_690,N_11840,N_10795);
or UO_691 (O_691,N_14170,N_10163);
or UO_692 (O_692,N_12338,N_13721);
nor UO_693 (O_693,N_12204,N_11450);
or UO_694 (O_694,N_11303,N_12229);
and UO_695 (O_695,N_13445,N_11931);
xnor UO_696 (O_696,N_12686,N_10192);
nand UO_697 (O_697,N_14909,N_12408);
nand UO_698 (O_698,N_10133,N_14848);
or UO_699 (O_699,N_11392,N_14303);
nand UO_700 (O_700,N_11152,N_13546);
nor UO_701 (O_701,N_14132,N_14596);
or UO_702 (O_702,N_10729,N_11229);
and UO_703 (O_703,N_14352,N_14422);
xnor UO_704 (O_704,N_11462,N_13537);
nand UO_705 (O_705,N_10911,N_14567);
or UO_706 (O_706,N_14423,N_13601);
or UO_707 (O_707,N_11638,N_10610);
and UO_708 (O_708,N_12826,N_12859);
nor UO_709 (O_709,N_14755,N_13302);
or UO_710 (O_710,N_12145,N_10442);
or UO_711 (O_711,N_13271,N_10760);
nand UO_712 (O_712,N_12521,N_12794);
or UO_713 (O_713,N_14850,N_13082);
and UO_714 (O_714,N_10652,N_12616);
nor UO_715 (O_715,N_14658,N_13255);
nand UO_716 (O_716,N_12571,N_12216);
or UO_717 (O_717,N_14817,N_13329);
and UO_718 (O_718,N_14280,N_13372);
nand UO_719 (O_719,N_12203,N_14234);
or UO_720 (O_720,N_11053,N_13493);
or UO_721 (O_721,N_14072,N_14121);
and UO_722 (O_722,N_10461,N_11644);
or UO_723 (O_723,N_14349,N_11481);
or UO_724 (O_724,N_13989,N_12678);
nand UO_725 (O_725,N_12021,N_11503);
nand UO_726 (O_726,N_10330,N_14885);
or UO_727 (O_727,N_13210,N_12375);
and UO_728 (O_728,N_10605,N_13638);
xnor UO_729 (O_729,N_10949,N_12376);
nand UO_730 (O_730,N_11870,N_11587);
and UO_731 (O_731,N_10304,N_10759);
and UO_732 (O_732,N_10953,N_11231);
xnor UO_733 (O_733,N_12987,N_13350);
nand UO_734 (O_734,N_10588,N_13340);
nand UO_735 (O_735,N_10902,N_10253);
nand UO_736 (O_736,N_13829,N_12780);
xnor UO_737 (O_737,N_11226,N_12505);
or UO_738 (O_738,N_13309,N_10642);
nor UO_739 (O_739,N_14725,N_11873);
or UO_740 (O_740,N_12514,N_13659);
or UO_741 (O_741,N_14927,N_14544);
and UO_742 (O_742,N_13156,N_13453);
and UO_743 (O_743,N_11745,N_12154);
or UO_744 (O_744,N_13217,N_10747);
and UO_745 (O_745,N_12388,N_11527);
nor UO_746 (O_746,N_11270,N_14267);
nor UO_747 (O_747,N_11717,N_12993);
or UO_748 (O_748,N_10924,N_11577);
nor UO_749 (O_749,N_11327,N_13935);
or UO_750 (O_750,N_14627,N_10766);
and UO_751 (O_751,N_13480,N_13242);
nor UO_752 (O_752,N_10938,N_11402);
or UO_753 (O_753,N_14686,N_10480);
nor UO_754 (O_754,N_11425,N_11650);
nor UO_755 (O_755,N_14041,N_12872);
nand UO_756 (O_756,N_11997,N_13161);
or UO_757 (O_757,N_11723,N_13631);
nand UO_758 (O_758,N_13027,N_10422);
nand UO_759 (O_759,N_12899,N_10905);
and UO_760 (O_760,N_13583,N_12333);
or UO_761 (O_761,N_13576,N_14481);
and UO_762 (O_762,N_13708,N_11120);
and UO_763 (O_763,N_14396,N_12152);
and UO_764 (O_764,N_11032,N_14374);
nor UO_765 (O_765,N_13769,N_11364);
nor UO_766 (O_766,N_12489,N_10144);
nor UO_767 (O_767,N_10717,N_12423);
nand UO_768 (O_768,N_11180,N_10294);
nor UO_769 (O_769,N_11744,N_10825);
nor UO_770 (O_770,N_10415,N_11372);
or UO_771 (O_771,N_10492,N_10362);
or UO_772 (O_772,N_11896,N_11612);
and UO_773 (O_773,N_13855,N_12980);
and UO_774 (O_774,N_13459,N_10509);
and UO_775 (O_775,N_12386,N_12874);
nor UO_776 (O_776,N_12522,N_14568);
or UO_777 (O_777,N_13745,N_12046);
nor UO_778 (O_778,N_12628,N_14903);
or UO_779 (O_779,N_12366,N_13227);
nor UO_780 (O_780,N_13818,N_13170);
and UO_781 (O_781,N_14366,N_11800);
and UO_782 (O_782,N_13119,N_10276);
nor UO_783 (O_783,N_10616,N_10183);
and UO_784 (O_784,N_12032,N_10172);
and UO_785 (O_785,N_12392,N_14052);
nand UO_786 (O_786,N_14865,N_14516);
nor UO_787 (O_787,N_11233,N_13142);
nand UO_788 (O_788,N_11182,N_13470);
and UO_789 (O_789,N_11135,N_12633);
or UO_790 (O_790,N_11813,N_13386);
nor UO_791 (O_791,N_14731,N_11158);
nand UO_792 (O_792,N_11059,N_10926);
or UO_793 (O_793,N_14835,N_11698);
nand UO_794 (O_794,N_14722,N_12982);
nand UO_795 (O_795,N_14929,N_11446);
nand UO_796 (O_796,N_14944,N_13775);
or UO_797 (O_797,N_13178,N_11704);
nor UO_798 (O_798,N_12432,N_13525);
nand UO_799 (O_799,N_12117,N_12783);
nand UO_800 (O_800,N_13632,N_14274);
or UO_801 (O_801,N_12630,N_10235);
nor UO_802 (O_802,N_14313,N_13960);
nand UO_803 (O_803,N_12720,N_11477);
nand UO_804 (O_804,N_11803,N_11090);
nand UO_805 (O_805,N_14024,N_10950);
or UO_806 (O_806,N_12414,N_11828);
or UO_807 (O_807,N_11596,N_11777);
xnor UO_808 (O_808,N_13478,N_12542);
nand UO_809 (O_809,N_12267,N_12265);
nand UO_810 (O_810,N_14499,N_13241);
nand UO_811 (O_811,N_12411,N_12033);
or UO_812 (O_812,N_13698,N_12971);
nand UO_813 (O_813,N_11572,N_11883);
nand UO_814 (O_814,N_14689,N_13880);
or UO_815 (O_815,N_11845,N_12784);
or UO_816 (O_816,N_14085,N_14493);
nor UO_817 (O_817,N_13617,N_12672);
and UO_818 (O_818,N_10006,N_12440);
or UO_819 (O_819,N_13171,N_12346);
nand UO_820 (O_820,N_14338,N_13221);
or UO_821 (O_821,N_13819,N_10774);
nor UO_822 (O_822,N_10574,N_11265);
nand UO_823 (O_823,N_10623,N_11910);
nand UO_824 (O_824,N_12789,N_12344);
nor UO_825 (O_825,N_14204,N_10578);
nand UO_826 (O_826,N_12892,N_13428);
or UO_827 (O_827,N_14212,N_10092);
nand UO_828 (O_828,N_12583,N_11218);
and UO_829 (O_829,N_13485,N_12725);
nor UO_830 (O_830,N_12788,N_12416);
and UO_831 (O_831,N_12096,N_10342);
and UO_832 (O_832,N_10508,N_12185);
and UO_833 (O_833,N_10032,N_14223);
or UO_834 (O_834,N_11618,N_10256);
xnor UO_835 (O_835,N_14748,N_11702);
nand UO_836 (O_836,N_10743,N_11044);
and UO_837 (O_837,N_12916,N_13999);
and UO_838 (O_838,N_12933,N_12885);
nand UO_839 (O_839,N_10413,N_14008);
and UO_840 (O_840,N_10433,N_11977);
or UO_841 (O_841,N_12064,N_14408);
nor UO_842 (O_842,N_12339,N_11015);
or UO_843 (O_843,N_12076,N_12184);
and UO_844 (O_844,N_14289,N_10797);
or UO_845 (O_845,N_10493,N_11543);
xnor UO_846 (O_846,N_11652,N_13123);
nand UO_847 (O_847,N_13300,N_12835);
nor UO_848 (O_848,N_10065,N_10217);
nor UO_849 (O_849,N_11400,N_10929);
and UO_850 (O_850,N_13817,N_12051);
nor UO_851 (O_851,N_11393,N_12439);
or UO_852 (O_852,N_10595,N_14741);
or UO_853 (O_853,N_11074,N_11139);
or UO_854 (O_854,N_14656,N_13658);
or UO_855 (O_855,N_11509,N_13474);
and UO_856 (O_856,N_12581,N_10780);
nand UO_857 (O_857,N_12322,N_11433);
or UO_858 (O_858,N_11232,N_12760);
or UO_859 (O_859,N_11706,N_11164);
or UO_860 (O_860,N_10108,N_13021);
nand UO_861 (O_861,N_11885,N_14517);
and UO_862 (O_862,N_12923,N_12167);
or UO_863 (O_863,N_12361,N_12969);
or UO_864 (O_864,N_10423,N_11035);
or UO_865 (O_865,N_11329,N_13265);
and UO_866 (O_866,N_10009,N_12832);
nand UO_867 (O_867,N_13628,N_10756);
and UO_868 (O_868,N_12809,N_14467);
nand UO_869 (O_869,N_10918,N_14724);
or UO_870 (O_870,N_10809,N_14803);
and UO_871 (O_871,N_12035,N_11278);
nand UO_872 (O_872,N_10946,N_14359);
nor UO_873 (O_873,N_12683,N_10694);
nand UO_874 (O_874,N_13177,N_14029);
nor UO_875 (O_875,N_12374,N_12104);
nor UO_876 (O_876,N_13748,N_13567);
or UO_877 (O_877,N_14772,N_10082);
and UO_878 (O_878,N_11279,N_10443);
and UO_879 (O_879,N_12690,N_11110);
nor UO_880 (O_880,N_11494,N_13535);
nand UO_881 (O_881,N_13754,N_10818);
nand UO_882 (O_882,N_10999,N_11614);
and UO_883 (O_883,N_14989,N_10220);
nor UO_884 (O_884,N_11206,N_11322);
xor UO_885 (O_885,N_11728,N_13231);
nor UO_886 (O_886,N_12134,N_11118);
nor UO_887 (O_887,N_13085,N_12400);
nor UO_888 (O_888,N_12010,N_11342);
nand UO_889 (O_889,N_13604,N_10152);
and UO_890 (O_890,N_10811,N_11389);
nor UO_891 (O_891,N_12124,N_14720);
and UO_892 (O_892,N_13692,N_13931);
and UO_893 (O_893,N_14239,N_12111);
and UO_894 (O_894,N_11592,N_10121);
xnor UO_895 (O_895,N_12682,N_11762);
or UO_896 (O_896,N_12379,N_11192);
xor UO_897 (O_897,N_14470,N_10677);
nor UO_898 (O_898,N_13281,N_11257);
nand UO_899 (O_899,N_10927,N_12483);
xor UO_900 (O_900,N_14344,N_13578);
and UO_901 (O_901,N_14362,N_11190);
nor UO_902 (O_902,N_10726,N_11660);
nor UO_903 (O_903,N_11812,N_10054);
or UO_904 (O_904,N_12620,N_11209);
and UO_905 (O_905,N_14080,N_14354);
nand UO_906 (O_906,N_11918,N_10609);
nand UO_907 (O_907,N_12708,N_11682);
and UO_908 (O_908,N_10887,N_11166);
xnor UO_909 (O_909,N_13710,N_14925);
and UO_910 (O_910,N_11850,N_12554);
nand UO_911 (O_911,N_10542,N_13247);
and UO_912 (O_912,N_11466,N_12195);
or UO_913 (O_913,N_14528,N_12823);
or UO_914 (O_914,N_13294,N_10596);
or UO_915 (O_915,N_13866,N_12803);
xnor UO_916 (O_916,N_14954,N_14697);
or UO_917 (O_917,N_12662,N_10854);
nand UO_918 (O_918,N_14797,N_13785);
or UO_919 (O_919,N_10334,N_10405);
nand UO_920 (O_920,N_12771,N_11245);
and UO_921 (O_921,N_13668,N_13730);
and UO_922 (O_922,N_11467,N_10132);
and UO_923 (O_923,N_13136,N_13997);
and UO_924 (O_924,N_14124,N_10236);
nor UO_925 (O_925,N_11797,N_12245);
nor UO_926 (O_926,N_13401,N_14140);
or UO_927 (O_927,N_14062,N_13365);
nor UO_928 (O_928,N_13469,N_11408);
or UO_929 (O_929,N_12748,N_12257);
nand UO_930 (O_930,N_13676,N_14915);
nand UO_931 (O_931,N_11191,N_13656);
nand UO_932 (O_932,N_11377,N_14071);
and UO_933 (O_933,N_11470,N_13176);
and UO_934 (O_934,N_12378,N_13367);
and UO_935 (O_935,N_14751,N_13444);
nand UO_936 (O_936,N_14894,N_10841);
xor UO_937 (O_937,N_11854,N_14259);
nand UO_938 (O_938,N_14027,N_11371);
xnor UO_939 (O_939,N_11932,N_11472);
nor UO_940 (O_940,N_11159,N_10420);
nand UO_941 (O_941,N_10285,N_11987);
nand UO_942 (O_942,N_11601,N_12970);
nor UO_943 (O_943,N_14106,N_13392);
or UO_944 (O_944,N_13853,N_13640);
or UO_945 (O_945,N_14270,N_10403);
nand UO_946 (O_946,N_14668,N_12973);
xor UO_947 (O_947,N_11397,N_11437);
and UO_948 (O_948,N_10604,N_10892);
and UO_949 (O_949,N_10688,N_12800);
and UO_950 (O_950,N_13279,N_11448);
nor UO_951 (O_951,N_13216,N_13804);
and UO_952 (O_952,N_14757,N_10611);
nand UO_953 (O_953,N_11262,N_10375);
xor UO_954 (O_954,N_13440,N_12426);
nor UO_955 (O_955,N_10764,N_14286);
nand UO_956 (O_956,N_11290,N_10742);
nor UO_957 (O_957,N_14141,N_11326);
and UO_958 (O_958,N_12370,N_14639);
nand UO_959 (O_959,N_12287,N_14524);
and UO_960 (O_960,N_14683,N_13034);
nor UO_961 (O_961,N_14157,N_10857);
nand UO_962 (O_962,N_12520,N_12791);
nor UO_963 (O_963,N_14692,N_12329);
or UO_964 (O_964,N_12449,N_13772);
or UO_965 (O_965,N_10459,N_12592);
and UO_966 (O_966,N_10391,N_10886);
or UO_967 (O_967,N_10482,N_10019);
nand UO_968 (O_968,N_10079,N_14805);
xor UO_969 (O_969,N_14680,N_12140);
nand UO_970 (O_970,N_14146,N_13421);
xnor UO_971 (O_971,N_10883,N_10318);
and UO_972 (O_972,N_13597,N_12639);
or UO_973 (O_973,N_12997,N_14203);
nor UO_974 (O_974,N_14908,N_14711);
and UO_975 (O_975,N_12097,N_13417);
or UO_976 (O_976,N_13023,N_11094);
nor UO_977 (O_977,N_10648,N_10406);
or UO_978 (O_978,N_14137,N_10730);
or UO_979 (O_979,N_11878,N_13621);
or UO_980 (O_980,N_14340,N_13379);
nand UO_981 (O_981,N_12040,N_14983);
nor UO_982 (O_982,N_13364,N_11900);
and UO_983 (O_983,N_14139,N_12082);
or UO_984 (O_984,N_14550,N_12836);
and UO_985 (O_985,N_11738,N_13982);
xnor UO_986 (O_986,N_11356,N_11630);
or UO_987 (O_987,N_10201,N_14331);
nand UO_988 (O_988,N_13719,N_12796);
or UO_989 (O_989,N_13048,N_12618);
nand UO_990 (O_990,N_12873,N_11559);
nor UO_991 (O_991,N_10973,N_10470);
nand UO_992 (O_992,N_13971,N_11700);
and UO_993 (O_993,N_10181,N_10862);
nor UO_994 (O_994,N_13511,N_11725);
xor UO_995 (O_995,N_12673,N_12840);
nand UO_996 (O_996,N_14454,N_12734);
nand UO_997 (O_997,N_14587,N_12918);
and UO_998 (O_998,N_12944,N_11775);
nand UO_999 (O_999,N_13933,N_11134);
nand UO_1000 (O_1000,N_13081,N_12200);
or UO_1001 (O_1001,N_13442,N_14785);
nand UO_1002 (O_1002,N_11718,N_14059);
and UO_1003 (O_1003,N_13352,N_12197);
nor UO_1004 (O_1004,N_13237,N_14369);
or UO_1005 (O_1005,N_13565,N_13052);
or UO_1006 (O_1006,N_14998,N_11037);
nor UO_1007 (O_1007,N_10531,N_14166);
nand UO_1008 (O_1008,N_13046,N_13066);
nor UO_1009 (O_1009,N_14094,N_12610);
or UO_1010 (O_1010,N_14190,N_14194);
nand UO_1011 (O_1011,N_14476,N_12888);
nor UO_1012 (O_1012,N_13805,N_14033);
nand UO_1013 (O_1013,N_12246,N_13794);
nor UO_1014 (O_1014,N_12192,N_14213);
and UO_1015 (O_1015,N_12274,N_11922);
or UO_1016 (O_1016,N_14007,N_11375);
or UO_1017 (O_1017,N_12303,N_12671);
nand UO_1018 (O_1018,N_12728,N_11453);
nor UO_1019 (O_1019,N_10316,N_12025);
nor UO_1020 (O_1020,N_11335,N_14530);
and UO_1021 (O_1021,N_10495,N_14039);
nor UO_1022 (O_1022,N_13561,N_13682);
or UO_1023 (O_1023,N_11637,N_11310);
or UO_1024 (O_1024,N_14918,N_11505);
or UO_1025 (O_1025,N_14713,N_14777);
or UO_1026 (O_1026,N_14405,N_11007);
xnor UO_1027 (O_1027,N_11028,N_11224);
nor UO_1028 (O_1028,N_10042,N_11411);
or UO_1029 (O_1029,N_11432,N_10922);
nand UO_1030 (O_1030,N_11001,N_10137);
or UO_1031 (O_1031,N_13756,N_11653);
and UO_1032 (O_1032,N_11244,N_14341);
nor UO_1033 (O_1033,N_14933,N_12550);
nor UO_1034 (O_1034,N_10657,N_12270);
and UO_1035 (O_1035,N_13564,N_10063);
xor UO_1036 (O_1036,N_13193,N_14442);
nor UO_1037 (O_1037,N_13863,N_13095);
or UO_1038 (O_1038,N_10600,N_12898);
or UO_1039 (O_1039,N_11769,N_10441);
and UO_1040 (O_1040,N_13252,N_13348);
or UO_1041 (O_1041,N_12454,N_11670);
nor UO_1042 (O_1042,N_10978,N_13323);
xor UO_1043 (O_1043,N_12242,N_14898);
or UO_1044 (O_1044,N_14960,N_11101);
and UO_1045 (O_1045,N_10635,N_10045);
and UO_1046 (O_1046,N_11949,N_10462);
and UO_1047 (O_1047,N_12591,N_11946);
or UO_1048 (O_1048,N_14483,N_13551);
or UO_1049 (O_1049,N_13297,N_13861);
or UO_1050 (O_1050,N_13019,N_11799);
and UO_1051 (O_1051,N_12022,N_10667);
nand UO_1052 (O_1052,N_13418,N_12028);
and UO_1053 (O_1053,N_10681,N_13899);
nand UO_1054 (O_1054,N_12883,N_12218);
xnor UO_1055 (O_1055,N_11130,N_13003);
and UO_1056 (O_1056,N_10118,N_14446);
nand UO_1057 (O_1057,N_14696,N_14688);
nor UO_1058 (O_1058,N_11011,N_14262);
and UO_1059 (O_1059,N_13187,N_11619);
nand UO_1060 (O_1060,N_11565,N_12561);
or UO_1061 (O_1061,N_11501,N_10127);
or UO_1062 (O_1062,N_11442,N_13100);
nand UO_1063 (O_1063,N_13113,N_14823);
and UO_1064 (O_1064,N_11832,N_14226);
or UO_1065 (O_1065,N_13949,N_10007);
or UO_1066 (O_1066,N_10347,N_11547);
nor UO_1067 (O_1067,N_13128,N_14521);
nand UO_1068 (O_1068,N_12629,N_13099);
and UO_1069 (O_1069,N_11349,N_13215);
and UO_1070 (O_1070,N_11020,N_13695);
or UO_1071 (O_1071,N_12927,N_10563);
or UO_1072 (O_1072,N_12533,N_13324);
nor UO_1073 (O_1073,N_14533,N_11106);
or UO_1074 (O_1074,N_10041,N_14009);
xnor UO_1075 (O_1075,N_10071,N_12304);
and UO_1076 (O_1076,N_12631,N_13000);
xnor UO_1077 (O_1077,N_10390,N_10565);
xnor UO_1078 (O_1078,N_14240,N_13071);
and UO_1079 (O_1079,N_14818,N_14266);
nor UO_1080 (O_1080,N_13928,N_11755);
xnor UO_1081 (O_1081,N_10842,N_12710);
and UO_1082 (O_1082,N_10984,N_10545);
and UO_1083 (O_1083,N_13747,N_12705);
nor UO_1084 (O_1084,N_13802,N_12867);
and UO_1085 (O_1085,N_14004,N_10029);
and UO_1086 (O_1086,N_14820,N_14886);
nand UO_1087 (O_1087,N_11863,N_13850);
or UO_1088 (O_1088,N_14705,N_11490);
xnor UO_1089 (O_1089,N_13793,N_13751);
nor UO_1090 (O_1090,N_13998,N_13315);
nor UO_1091 (O_1091,N_10877,N_11391);
and UO_1092 (O_1092,N_13768,N_11880);
or UO_1093 (O_1093,N_13434,N_10644);
or UO_1094 (O_1094,N_12845,N_11760);
nor UO_1095 (O_1095,N_14970,N_12068);
and UO_1096 (O_1096,N_11579,N_13077);
and UO_1097 (O_1097,N_10662,N_12019);
and UO_1098 (O_1098,N_14254,N_10601);
and UO_1099 (O_1099,N_12706,N_14794);
and UO_1100 (O_1100,N_14087,N_12441);
and UO_1101 (O_1101,N_10994,N_14443);
and UO_1102 (O_1102,N_13425,N_14380);
nand UO_1103 (O_1103,N_12909,N_13762);
xor UO_1104 (O_1104,N_11690,N_13996);
nor UO_1105 (O_1105,N_14079,N_14475);
or UO_1106 (O_1106,N_14682,N_14875);
nor UO_1107 (O_1107,N_12989,N_13508);
nor UO_1108 (O_1108,N_12238,N_11716);
or UO_1109 (O_1109,N_10335,N_13520);
nor UO_1110 (O_1110,N_11530,N_11645);
xnor UO_1111 (O_1111,N_14896,N_10431);
and UO_1112 (O_1112,N_10543,N_14000);
nand UO_1113 (O_1113,N_14304,N_10653);
nand UO_1114 (O_1114,N_10056,N_14880);
and UO_1115 (O_1115,N_14985,N_14961);
or UO_1116 (O_1116,N_13732,N_12664);
xnor UO_1117 (O_1117,N_10977,N_14726);
nor UO_1118 (O_1118,N_11132,N_10076);
nand UO_1119 (O_1119,N_14845,N_13301);
nor UO_1120 (O_1120,N_11343,N_14921);
and UO_1121 (O_1121,N_11676,N_14555);
or UO_1122 (O_1122,N_14844,N_12083);
nor UO_1123 (O_1123,N_12778,N_14760);
and UO_1124 (O_1124,N_12436,N_12405);
xor UO_1125 (O_1125,N_13800,N_11420);
nand UO_1126 (O_1126,N_14502,N_13032);
and UO_1127 (O_1127,N_12327,N_13677);
and UO_1128 (O_1128,N_12012,N_10521);
nor UO_1129 (O_1129,N_13266,N_13514);
and UO_1130 (O_1130,N_12491,N_12818);
and UO_1131 (O_1131,N_12921,N_12570);
nor UO_1132 (O_1132,N_12857,N_14832);
nand UO_1133 (O_1133,N_14152,N_13739);
and UO_1134 (O_1134,N_10363,N_11898);
and UO_1135 (O_1135,N_14623,N_13017);
xor UO_1136 (O_1136,N_13889,N_12717);
or UO_1137 (O_1137,N_13815,N_12105);
xnor UO_1138 (O_1138,N_12390,N_14761);
nand UO_1139 (O_1139,N_14675,N_12061);
or UO_1140 (O_1140,N_13699,N_11154);
nand UO_1141 (O_1141,N_10282,N_13887);
and UO_1142 (O_1142,N_10286,N_11616);
nor UO_1143 (O_1143,N_14257,N_12004);
nor UO_1144 (O_1144,N_14578,N_14821);
nor UO_1145 (O_1145,N_13679,N_12443);
nand UO_1146 (O_1146,N_12199,N_13260);
nand UO_1147 (O_1147,N_13810,N_11113);
or UO_1148 (O_1148,N_12089,N_11195);
and UO_1149 (O_1149,N_13693,N_12943);
or UO_1150 (O_1150,N_11537,N_12328);
nand UO_1151 (O_1151,N_13299,N_12563);
xnor UO_1152 (O_1152,N_13864,N_14111);
and UO_1153 (O_1153,N_12078,N_10317);
and UO_1154 (O_1154,N_13943,N_12573);
and UO_1155 (O_1155,N_13634,N_10556);
nand UO_1156 (O_1156,N_13334,N_13224);
nor UO_1157 (O_1157,N_14606,N_14164);
nand UO_1158 (O_1158,N_14188,N_10861);
nor UO_1159 (O_1159,N_14546,N_14931);
nor UO_1160 (O_1160,N_11487,N_10024);
nand UO_1161 (O_1161,N_12276,N_13595);
and UO_1162 (O_1162,N_14882,N_11567);
or UO_1163 (O_1163,N_11023,N_13666);
and UO_1164 (O_1164,N_12331,N_13262);
nand UO_1165 (O_1165,N_13482,N_11165);
or UO_1166 (O_1166,N_13056,N_12394);
nand UO_1167 (O_1167,N_11533,N_12847);
nor UO_1168 (O_1168,N_11235,N_10147);
nand UO_1169 (O_1169,N_11569,N_13026);
nor UO_1170 (O_1170,N_11299,N_12718);
or UO_1171 (O_1171,N_12733,N_11384);
nand UO_1172 (O_1172,N_10337,N_12607);
nand UO_1173 (O_1173,N_14339,N_12674);
or UO_1174 (O_1174,N_12777,N_12335);
nor UO_1175 (O_1175,N_10835,N_14330);
nand UO_1176 (O_1176,N_10404,N_12147);
nand UO_1177 (O_1177,N_12249,N_12834);
or UO_1178 (O_1178,N_11502,N_11764);
nor UO_1179 (O_1179,N_13605,N_11695);
xnor UO_1180 (O_1180,N_13393,N_13347);
nand UO_1181 (O_1181,N_10271,N_13004);
and UO_1182 (O_1182,N_14743,N_12183);
nand UO_1183 (O_1183,N_11256,N_10075);
nor UO_1184 (O_1184,N_11693,N_10265);
and UO_1185 (O_1185,N_14774,N_10175);
or UO_1186 (O_1186,N_13054,N_12015);
nor UO_1187 (O_1187,N_12310,N_13016);
nor UO_1188 (O_1188,N_11452,N_10259);
nor UO_1189 (O_1189,N_10494,N_14172);
or UO_1190 (O_1190,N_14847,N_14384);
xnor UO_1191 (O_1191,N_12547,N_13378);
nor UO_1192 (O_1192,N_13107,N_14614);
and UO_1193 (O_1193,N_10689,N_13416);
and UO_1194 (O_1194,N_12601,N_14831);
nor UO_1195 (O_1195,N_13132,N_14119);
and UO_1196 (O_1196,N_12985,N_13269);
xnor UO_1197 (O_1197,N_12820,N_11665);
or UO_1198 (O_1198,N_10878,N_14939);
nand UO_1199 (O_1199,N_11027,N_10956);
xor UO_1200 (O_1200,N_10238,N_13001);
xor UO_1201 (O_1201,N_12013,N_14327);
or UO_1202 (O_1202,N_13086,N_12917);
nand UO_1203 (O_1203,N_11398,N_12851);
nor UO_1204 (O_1204,N_14265,N_10243);
or UO_1205 (O_1205,N_13780,N_14207);
or UO_1206 (O_1206,N_11148,N_13292);
nor UO_1207 (O_1207,N_13515,N_11507);
and UO_1208 (O_1208,N_10896,N_11228);
nor UO_1209 (O_1209,N_12900,N_14872);
nand UO_1210 (O_1210,N_13129,N_11348);
nand UO_1211 (O_1211,N_14120,N_10844);
or UO_1212 (O_1212,N_11168,N_12595);
nand UO_1213 (O_1213,N_14061,N_10170);
nand UO_1214 (O_1214,N_14082,N_13837);
nor UO_1215 (O_1215,N_13201,N_14434);
and UO_1216 (O_1216,N_14098,N_14371);
nand UO_1217 (O_1217,N_11178,N_11916);
or UO_1218 (O_1218,N_13424,N_13588);
and UO_1219 (O_1219,N_14002,N_10026);
or UO_1220 (O_1220,N_11879,N_12315);
nor UO_1221 (O_1221,N_12325,N_12744);
and UO_1222 (O_1222,N_10849,N_11791);
or UO_1223 (O_1223,N_10627,N_11817);
nand UO_1224 (O_1224,N_11394,N_11624);
and UO_1225 (O_1225,N_11492,N_12626);
and UO_1226 (O_1226,N_11323,N_11669);
or UO_1227 (O_1227,N_12324,N_10379);
nor UO_1228 (O_1228,N_14118,N_14075);
nor UO_1229 (O_1229,N_10308,N_10991);
xor UO_1230 (O_1230,N_13189,N_12174);
or UO_1231 (O_1231,N_14735,N_12337);
and UO_1232 (O_1232,N_14766,N_10920);
nor UO_1233 (O_1233,N_11221,N_10840);
or UO_1234 (O_1234,N_13916,N_13006);
nor UO_1235 (O_1235,N_13158,N_14100);
and UO_1236 (O_1236,N_12555,N_14237);
and UO_1237 (O_1237,N_11983,N_13268);
or UO_1238 (O_1238,N_12005,N_11555);
and UO_1239 (O_1239,N_14804,N_11641);
and UO_1240 (O_1240,N_13455,N_12992);
nand UO_1241 (O_1241,N_12797,N_12263);
xnor UO_1242 (O_1242,N_13622,N_10369);
and UO_1243 (O_1243,N_11043,N_10325);
and UO_1244 (O_1244,N_10209,N_10964);
nor UO_1245 (O_1245,N_12188,N_14329);
nand UO_1246 (O_1246,N_10148,N_14830);
xnor UO_1247 (O_1247,N_11779,N_12404);
xor UO_1248 (O_1248,N_13970,N_11719);
and UO_1249 (O_1249,N_14251,N_11145);
nor UO_1250 (O_1250,N_14500,N_10554);
or UO_1251 (O_1251,N_11198,N_10010);
nand UO_1252 (O_1252,N_10023,N_10193);
nor UO_1253 (O_1253,N_11506,N_14403);
nand UO_1254 (O_1254,N_10829,N_13181);
nand UO_1255 (O_1255,N_10884,N_12070);
or UO_1256 (O_1256,N_11449,N_10430);
xnor UO_1257 (O_1257,N_11478,N_11627);
nand UO_1258 (O_1258,N_10327,N_14221);
or UO_1259 (O_1259,N_13044,N_11079);
and UO_1260 (O_1260,N_12512,N_12724);
or UO_1261 (O_1261,N_11358,N_10223);
xnor UO_1262 (O_1262,N_10130,N_14068);
or UO_1263 (O_1263,N_14945,N_11734);
nor UO_1264 (O_1264,N_11990,N_10866);
nor UO_1265 (O_1265,N_11536,N_14852);
nor UO_1266 (O_1266,N_12356,N_13712);
nor UO_1267 (O_1267,N_12306,N_11283);
xor UO_1268 (O_1268,N_13702,N_14168);
and UO_1269 (O_1269,N_14155,N_12833);
nor UO_1270 (O_1270,N_12651,N_10104);
xnor UO_1271 (O_1271,N_11097,N_11766);
and UO_1272 (O_1272,N_12090,N_11701);
xnor UO_1273 (O_1273,N_11768,N_13212);
nor UO_1274 (O_1274,N_11464,N_10602);
xnor UO_1275 (O_1275,N_13454,N_12357);
or UO_1276 (O_1276,N_11170,N_13152);
nand UO_1277 (O_1277,N_10425,N_14358);
nand UO_1278 (O_1278,N_14295,N_13787);
and UO_1279 (O_1279,N_11050,N_13981);
nand UO_1280 (O_1280,N_14849,N_11194);
and UO_1281 (O_1281,N_13433,N_12978);
xnor UO_1282 (O_1282,N_10864,N_12319);
and UO_1283 (O_1283,N_12116,N_11570);
or UO_1284 (O_1284,N_12621,N_13169);
or UO_1285 (O_1285,N_11396,N_13968);
nand UO_1286 (O_1286,N_14288,N_14801);
nand UO_1287 (O_1287,N_11246,N_14868);
nor UO_1288 (O_1288,N_10558,N_10445);
nand UO_1289 (O_1289,N_11320,N_10526);
xor UO_1290 (O_1290,N_13125,N_10249);
nor UO_1291 (O_1291,N_11018,N_13993);
nand UO_1292 (O_1292,N_12490,N_13160);
and UO_1293 (O_1293,N_12792,N_11771);
xor UO_1294 (O_1294,N_12950,N_11882);
nand UO_1295 (O_1295,N_12905,N_10820);
nor UO_1296 (O_1296,N_13969,N_10520);
xnor UO_1297 (O_1297,N_14911,N_11711);
or UO_1298 (O_1298,N_10777,N_11374);
and UO_1299 (O_1299,N_11677,N_13976);
and UO_1300 (O_1300,N_14992,N_14073);
and UO_1301 (O_1301,N_10359,N_12525);
xor UO_1302 (O_1302,N_10669,N_12413);
nor UO_1303 (O_1303,N_11611,N_12627);
and UO_1304 (O_1304,N_10607,N_10101);
and UO_1305 (O_1305,N_11523,N_13892);
nor UO_1306 (O_1306,N_14681,N_12876);
nor UO_1307 (O_1307,N_13930,N_11185);
nor UO_1308 (O_1308,N_13603,N_13020);
or UO_1309 (O_1309,N_14976,N_14863);
nand UO_1310 (O_1310,N_10784,N_11907);
or UO_1311 (O_1311,N_12059,N_10698);
nor UO_1312 (O_1312,N_13937,N_12611);
xnor UO_1313 (O_1313,N_11623,N_10583);
nand UO_1314 (O_1314,N_12913,N_13296);
xnor UO_1315 (O_1315,N_10229,N_12762);
and UO_1316 (O_1316,N_10503,N_12193);
or UO_1317 (O_1317,N_11911,N_10055);
nand UO_1318 (O_1318,N_14323,N_12665);
nand UO_1319 (O_1319,N_14089,N_10967);
xnor UO_1320 (O_1320,N_10636,N_12928);
nor UO_1321 (O_1321,N_14337,N_11642);
or UO_1322 (O_1322,N_11816,N_12795);
or UO_1323 (O_1323,N_11105,N_13580);
nand UO_1324 (O_1324,N_12172,N_12878);
nor UO_1325 (O_1325,N_14189,N_14273);
nor UO_1326 (O_1326,N_12709,N_12372);
nor UO_1327 (O_1327,N_14242,N_10974);
and UO_1328 (O_1328,N_12689,N_12881);
nand UO_1329 (O_1329,N_14055,N_12540);
nor UO_1330 (O_1330,N_12300,N_11005);
and UO_1331 (O_1331,N_14348,N_11149);
nor UO_1332 (O_1332,N_10125,N_13064);
nand UO_1333 (O_1333,N_14127,N_14756);
and UO_1334 (O_1334,N_10870,N_10872);
and UO_1335 (O_1335,N_10344,N_11137);
or UO_1336 (O_1336,N_12308,N_14890);
nand UO_1337 (O_1337,N_14150,N_12829);
nand UO_1338 (O_1338,N_14317,N_11674);
and UO_1339 (O_1339,N_12250,N_11955);
or UO_1340 (O_1340,N_14126,N_12255);
nand UO_1341 (O_1341,N_12486,N_13230);
or UO_1342 (O_1342,N_10963,N_10725);
nor UO_1343 (O_1343,N_12122,N_10646);
and UO_1344 (O_1344,N_10419,N_13090);
and UO_1345 (O_1345,N_14593,N_11080);
xor UO_1346 (O_1346,N_12455,N_14538);
and UO_1347 (O_1347,N_11853,N_14654);
and UO_1348 (O_1348,N_11761,N_13562);
and UO_1349 (O_1349,N_13040,N_14955);
and UO_1350 (O_1350,N_10103,N_10087);
nand UO_1351 (O_1351,N_10714,N_11000);
xnor UO_1352 (O_1352,N_13338,N_11514);
nand UO_1353 (O_1353,N_12624,N_13612);
and UO_1354 (O_1354,N_11124,N_13390);
xor UO_1355 (O_1355,N_10837,N_12473);
xnor UO_1356 (O_1356,N_12808,N_14884);
nand UO_1357 (O_1357,N_10933,N_14659);
nand UO_1358 (O_1358,N_14729,N_12515);
nand UO_1359 (O_1359,N_14814,N_10262);
and UO_1360 (O_1360,N_14006,N_13533);
nand UO_1361 (O_1361,N_14244,N_12640);
and UO_1362 (O_1362,N_14799,N_13906);
and UO_1363 (O_1363,N_12074,N_14813);
nand UO_1364 (O_1364,N_14589,N_13312);
or UO_1365 (O_1365,N_12434,N_11183);
nand UO_1366 (O_1366,N_10519,N_10140);
and UO_1367 (O_1367,N_10506,N_13890);
nor UO_1368 (O_1368,N_12115,N_11122);
or UO_1369 (O_1369,N_12911,N_11491);
and UO_1370 (O_1370,N_13431,N_12194);
nand UO_1371 (O_1371,N_10001,N_10427);
or UO_1372 (O_1372,N_12609,N_11306);
or UO_1373 (O_1373,N_13286,N_11036);
and UO_1374 (O_1374,N_11621,N_12049);
and UO_1375 (O_1375,N_13371,N_13407);
nor UO_1376 (O_1376,N_14594,N_10280);
nor UO_1377 (O_1377,N_14160,N_11471);
nor UO_1378 (O_1378,N_10206,N_12351);
nor UO_1379 (O_1379,N_14154,N_14811);
and UO_1380 (O_1380,N_11463,N_13116);
or UO_1381 (O_1381,N_14229,N_10227);
nor UO_1382 (O_1382,N_13448,N_13254);
nand UO_1383 (O_1383,N_10618,N_14488);
nor UO_1384 (O_1384,N_11708,N_11963);
and UO_1385 (O_1385,N_14342,N_13860);
nor UO_1386 (O_1386,N_12858,N_11970);
and UO_1387 (O_1387,N_13555,N_11199);
or UO_1388 (O_1388,N_13964,N_12026);
and UO_1389 (O_1389,N_10376,N_11461);
nor UO_1390 (O_1390,N_11678,N_14013);
nand UO_1391 (O_1391,N_12205,N_10358);
nand UO_1392 (O_1392,N_14965,N_13635);
nor UO_1393 (O_1393,N_10721,N_10020);
nor UO_1394 (O_1394,N_10576,N_13059);
nand UO_1395 (O_1395,N_13902,N_11925);
xor UO_1396 (O_1396,N_13782,N_10791);
nand UO_1397 (O_1397,N_11956,N_11271);
and UO_1398 (O_1398,N_10788,N_10196);
or UO_1399 (O_1399,N_13674,N_11988);
nor UO_1400 (O_1400,N_13354,N_12634);
xor UO_1401 (O_1401,N_12093,N_10906);
or UO_1402 (O_1402,N_14926,N_14518);
xnor UO_1403 (O_1403,N_10744,N_13942);
nand UO_1404 (O_1404,N_13966,N_10207);
nand UO_1405 (O_1405,N_10374,N_13423);
xnor UO_1406 (O_1406,N_14044,N_13013);
nand UO_1407 (O_1407,N_10264,N_10799);
and UO_1408 (O_1408,N_10254,N_12169);
and UO_1409 (O_1409,N_12954,N_11273);
and UO_1410 (O_1410,N_14249,N_13138);
and UO_1411 (O_1411,N_14430,N_11407);
or UO_1412 (O_1412,N_13738,N_10269);
or UO_1413 (O_1413,N_10322,N_10631);
xor UO_1414 (O_1414,N_11593,N_10416);
and UO_1415 (O_1415,N_12043,N_14637);
or UO_1416 (O_1416,N_12241,N_12092);
or UO_1417 (O_1417,N_11284,N_12860);
or UO_1418 (O_1418,N_14815,N_14334);
and UO_1419 (O_1419,N_10882,N_11557);
nor UO_1420 (O_1420,N_14498,N_13548);
or UO_1421 (O_1421,N_12011,N_13733);
nand UO_1422 (O_1422,N_10674,N_14390);
nand UO_1423 (O_1423,N_12934,N_14287);
nor UO_1424 (O_1424,N_10432,N_11640);
nand UO_1425 (O_1425,N_13647,N_13345);
or UO_1426 (O_1426,N_13957,N_11726);
or UO_1427 (O_1427,N_14474,N_11431);
nand UO_1428 (O_1428,N_11483,N_13664);
nand UO_1429 (O_1429,N_13939,N_10058);
xnor UO_1430 (O_1430,N_14856,N_13718);
nand UO_1431 (O_1431,N_13068,N_14990);
nand UO_1432 (O_1432,N_10901,N_10541);
xor UO_1433 (O_1433,N_11237,N_11899);
or UO_1434 (O_1434,N_12743,N_11729);
nor UO_1435 (O_1435,N_13681,N_11823);
nand UO_1436 (O_1436,N_13707,N_11004);
nand UO_1437 (O_1437,N_14559,N_12237);
or UO_1438 (O_1438,N_10451,N_14450);
nand UO_1439 (O_1439,N_14497,N_11843);
and UO_1440 (O_1440,N_11857,N_14948);
nand UO_1441 (O_1441,N_12207,N_13518);
or UO_1442 (O_1442,N_13363,N_10246);
nand UO_1443 (O_1443,N_10394,N_14414);
or UO_1444 (O_1444,N_14539,N_12130);
or UO_1445 (O_1445,N_13343,N_11923);
nor UO_1446 (O_1446,N_11819,N_14644);
nand UO_1447 (O_1447,N_10195,N_11146);
nand UO_1448 (O_1448,N_13697,N_10138);
and UO_1449 (O_1449,N_14492,N_10095);
and UO_1450 (O_1450,N_12757,N_12347);
nand UO_1451 (O_1451,N_11309,N_13529);
nor UO_1452 (O_1452,N_11196,N_11445);
nor UO_1453 (O_1453,N_13627,N_10932);
or UO_1454 (O_1454,N_13509,N_14135);
nor UO_1455 (O_1455,N_12389,N_13411);
xnor UO_1456 (O_1456,N_12736,N_11039);
or UO_1457 (O_1457,N_14095,N_14345);
and UO_1458 (O_1458,N_10758,N_11332);
nand UO_1459 (O_1459,N_13419,N_11671);
nor UO_1460 (O_1460,N_10934,N_10122);
and UO_1461 (O_1461,N_10960,N_13449);
or UO_1462 (O_1462,N_11679,N_12729);
or UO_1463 (O_1463,N_14400,N_10037);
and UO_1464 (O_1464,N_10173,N_13488);
or UO_1465 (O_1465,N_13593,N_14826);
or UO_1466 (O_1466,N_14368,N_14592);
and UO_1467 (O_1467,N_11620,N_13728);
or UO_1468 (O_1468,N_12869,N_12693);
or UO_1469 (O_1469,N_11367,N_14084);
or UO_1470 (O_1470,N_12027,N_12940);
nor UO_1471 (O_1471,N_10062,N_11301);
and UO_1472 (O_1472,N_12215,N_11108);
nand UO_1473 (O_1473,N_13349,N_14928);
nor UO_1474 (O_1474,N_10408,N_13397);
and UO_1475 (O_1475,N_10762,N_11227);
and UO_1476 (O_1476,N_13404,N_13248);
and UO_1477 (O_1477,N_10622,N_12608);
xnor UO_1478 (O_1478,N_13893,N_13196);
xnor UO_1479 (O_1479,N_11903,N_11535);
nand UO_1480 (O_1480,N_11941,N_12063);
nand UO_1481 (O_1481,N_14490,N_12042);
xor UO_1482 (O_1482,N_13545,N_13037);
nand UO_1483 (O_1483,N_14736,N_11069);
nand UO_1484 (O_1484,N_10720,N_11994);
nand UO_1485 (O_1485,N_12964,N_11296);
nand UO_1486 (O_1486,N_13502,N_13806);
xnor UO_1487 (O_1487,N_10114,N_12318);
or UO_1488 (O_1488,N_14110,N_13789);
xor UO_1489 (O_1489,N_12038,N_12470);
nor UO_1490 (O_1490,N_10186,N_12209);
and UO_1491 (O_1491,N_10340,N_13584);
nor UO_1492 (O_1492,N_10889,N_13385);
nand UO_1493 (O_1493,N_14321,N_10083);
xnor UO_1494 (O_1494,N_11203,N_13120);
nand UO_1495 (O_1495,N_12150,N_14026);
or UO_1496 (O_1496,N_13759,N_10831);
nor UO_1497 (O_1497,N_13162,N_14293);
nand UO_1498 (O_1498,N_12039,N_11872);
nand UO_1499 (O_1499,N_11082,N_12825);
nand UO_1500 (O_1500,N_10040,N_12668);
nand UO_1501 (O_1501,N_10510,N_13033);
or UO_1502 (O_1502,N_13620,N_11272);
nand UO_1503 (O_1503,N_14388,N_13277);
nor UO_1504 (O_1504,N_14537,N_11058);
nand UO_1505 (O_1505,N_13028,N_11792);
or UO_1506 (O_1506,N_10213,N_13270);
or UO_1507 (O_1507,N_11651,N_13307);
and UO_1508 (O_1508,N_13185,N_12301);
xor UO_1509 (O_1509,N_11985,N_11315);
and UO_1510 (O_1510,N_14357,N_13457);
and UO_1511 (O_1511,N_11801,N_10446);
or UO_1512 (O_1512,N_13438,N_14038);
nor UO_1513 (O_1513,N_11205,N_14290);
or UO_1514 (O_1514,N_10169,N_14281);
nor UO_1515 (O_1515,N_13873,N_11476);
nand UO_1516 (O_1516,N_11562,N_10782);
nand UO_1517 (O_1517,N_13475,N_12047);
xnor UO_1518 (O_1518,N_12870,N_12838);
and UO_1519 (O_1519,N_10022,N_13163);
or UO_1520 (O_1520,N_12142,N_11055);
xor UO_1521 (O_1521,N_12323,N_11696);
xnor UO_1522 (O_1522,N_11003,N_12448);
nor UO_1523 (O_1523,N_10489,N_14196);
nand UO_1524 (O_1524,N_13521,N_13613);
nand UO_1525 (O_1525,N_10145,N_13031);
and UO_1526 (O_1526,N_14461,N_13029);
xnor UO_1527 (O_1527,N_13995,N_13194);
nor UO_1528 (O_1528,N_10680,N_12701);
nand UO_1529 (O_1529,N_10952,N_13822);
xor UO_1530 (O_1530,N_11838,N_14432);
or UO_1531 (O_1531,N_12156,N_13512);
and UO_1532 (O_1532,N_12348,N_14058);
nand UO_1533 (O_1533,N_10155,N_14298);
nand UO_1534 (O_1534,N_13538,N_12383);
xor UO_1535 (O_1535,N_14264,N_11072);
nand UO_1536 (O_1536,N_10880,N_10448);
or UO_1537 (O_1537,N_10355,N_13070);
and UO_1538 (O_1538,N_12500,N_13736);
or UO_1539 (O_1539,N_13835,N_13910);
nor UO_1540 (O_1540,N_14796,N_12691);
nor UO_1541 (O_1541,N_14995,N_13792);
nand UO_1542 (O_1542,N_14090,N_12799);
nand UO_1543 (O_1543,N_14507,N_13568);
and UO_1544 (O_1544,N_10690,N_13924);
nor UO_1545 (O_1545,N_11289,N_10407);
or UO_1546 (O_1546,N_13917,N_11151);
and UO_1547 (O_1547,N_11625,N_14665);
nand UO_1548 (O_1548,N_12190,N_13074);
nand UO_1549 (O_1549,N_12451,N_10051);
xnor UO_1550 (O_1550,N_12648,N_10785);
or UO_1551 (O_1551,N_13904,N_11248);
or UO_1552 (O_1552,N_14112,N_13857);
or UO_1553 (O_1553,N_13927,N_10218);
nor UO_1554 (O_1554,N_10157,N_14677);
nand UO_1555 (O_1555,N_12073,N_10672);
nor UO_1556 (O_1556,N_11025,N_14704);
nor UO_1557 (O_1557,N_12737,N_12827);
nor UO_1558 (O_1558,N_14065,N_11542);
and UO_1559 (O_1559,N_12457,N_10997);
nand UO_1560 (O_1560,N_14629,N_13276);
nand UO_1561 (O_1561,N_13303,N_10439);
or UO_1562 (O_1562,N_14468,N_13662);
nor UO_1563 (O_1563,N_13945,N_13703);
nand UO_1564 (O_1564,N_10695,N_12819);
and UO_1565 (O_1565,N_12472,N_10296);
and UO_1566 (O_1566,N_13589,N_13895);
nor UO_1567 (O_1567,N_13954,N_11093);
xor UO_1568 (O_1568,N_14691,N_13619);
nand UO_1569 (O_1569,N_14612,N_11217);
nand UO_1570 (O_1570,N_14291,N_13922);
nor UO_1571 (O_1571,N_11906,N_13402);
nor UO_1572 (O_1572,N_11119,N_13118);
and UO_1573 (O_1573,N_12951,N_11796);
xor UO_1574 (O_1574,N_11721,N_13437);
and UO_1575 (O_1575,N_13552,N_14165);
or UO_1576 (O_1576,N_12935,N_10769);
nor UO_1577 (O_1577,N_10685,N_10851);
nand UO_1578 (O_1578,N_12409,N_10216);
nand UO_1579 (O_1579,N_12817,N_13741);
and UO_1580 (O_1580,N_10178,N_10381);
nor UO_1581 (O_1581,N_10002,N_13467);
nand UO_1582 (O_1582,N_11876,N_13809);
xor UO_1583 (O_1583,N_11772,N_13157);
nor UO_1584 (O_1584,N_13823,N_11549);
nor UO_1585 (O_1585,N_12588,N_11141);
nand UO_1586 (O_1586,N_12981,N_14702);
or UO_1587 (O_1587,N_10873,N_13965);
nand UO_1588 (O_1588,N_13610,N_14923);
nand UO_1589 (O_1589,N_13400,N_11919);
xor UO_1590 (O_1590,N_10323,N_10893);
nor UO_1591 (O_1591,N_10524,N_14460);
or UO_1592 (O_1592,N_11544,N_10982);
nand UO_1593 (O_1593,N_10808,N_13208);
or UO_1594 (O_1594,N_14391,N_12719);
nand UO_1595 (O_1595,N_12597,N_11282);
and UO_1596 (O_1596,N_13737,N_12444);
nand UO_1597 (O_1597,N_13357,N_14182);
nand UO_1598 (O_1598,N_13359,N_11707);
nand UO_1599 (O_1599,N_14542,N_14687);
and UO_1600 (O_1600,N_10969,N_12029);
nand UO_1601 (O_1601,N_11778,N_13093);
nand UO_1602 (O_1602,N_10839,N_10728);
xor UO_1603 (O_1603,N_12235,N_11347);
or UO_1604 (O_1604,N_13025,N_11864);
nand UO_1605 (O_1605,N_12275,N_11052);
nor UO_1606 (O_1606,N_10221,N_10398);
nor UO_1607 (O_1607,N_10313,N_11112);
nor UO_1608 (O_1608,N_13947,N_10930);
nand UO_1609 (O_1609,N_10663,N_10244);
nor UO_1610 (O_1610,N_12866,N_14997);
and UO_1611 (O_1611,N_13084,N_10985);
or UO_1612 (O_1612,N_11479,N_11167);
nor UO_1613 (O_1613,N_14513,N_13494);
and UO_1614 (O_1614,N_13691,N_12045);
nand UO_1615 (O_1615,N_12126,N_14786);
and UO_1616 (O_1616,N_11350,N_14640);
xnor UO_1617 (O_1617,N_13250,N_14781);
nor UO_1618 (O_1618,N_10990,N_13651);
nand UO_1619 (O_1619,N_12598,N_10149);
or UO_1620 (O_1620,N_13886,N_14864);
or UO_1621 (O_1621,N_14690,N_14651);
and UO_1622 (O_1622,N_12564,N_14676);
and UO_1623 (O_1623,N_10081,N_14113);
or UO_1624 (O_1624,N_13036,N_10412);
nor UO_1625 (O_1625,N_14284,N_11749);
and UO_1626 (O_1626,N_10704,N_14671);
or UO_1627 (O_1627,N_12844,N_12578);
nor UO_1628 (O_1628,N_11869,N_11063);
xor UO_1629 (O_1629,N_10165,N_13010);
xnor UO_1630 (O_1630,N_14699,N_13700);
or UO_1631 (O_1631,N_12442,N_10979);
xnor UO_1632 (O_1632,N_14211,N_12925);
nand UO_1633 (O_1633,N_10660,N_14561);
nand UO_1634 (O_1634,N_13126,N_11743);
and UO_1635 (O_1635,N_14030,N_10628);
or UO_1636 (O_1636,N_12003,N_13592);
nand UO_1637 (O_1637,N_10792,N_12438);
nand UO_1638 (O_1638,N_12368,N_14573);
or UO_1639 (O_1639,N_13188,N_13921);
nand UO_1640 (O_1640,N_12965,N_10928);
and UO_1641 (O_1641,N_10736,N_11783);
and UO_1642 (O_1642,N_11526,N_14968);
xnor UO_1643 (O_1643,N_10053,N_14402);
and UO_1644 (O_1644,N_14487,N_12433);
xnor UO_1645 (O_1645,N_12919,N_11029);
or UO_1646 (O_1646,N_10471,N_10447);
nor UO_1647 (O_1647,N_10307,N_12752);
or UO_1648 (O_1648,N_13838,N_14953);
or UO_1649 (O_1649,N_14672,N_13022);
and UO_1650 (O_1650,N_12868,N_10500);
nor UO_1651 (O_1651,N_10552,N_14728);
xor UO_1652 (O_1652,N_13443,N_10182);
nand UO_1653 (O_1653,N_13831,N_10536);
nor UO_1654 (O_1654,N_10463,N_12007);
and UO_1655 (O_1655,N_13720,N_11773);
or UO_1656 (O_1656,N_12178,N_11525);
and UO_1657 (O_1657,N_12326,N_14846);
nand UO_1658 (O_1658,N_11370,N_14496);
nor UO_1659 (O_1659,N_12747,N_10836);
nor UO_1660 (O_1660,N_11121,N_13149);
nor UO_1661 (O_1661,N_14315,N_14564);
and UO_1662 (O_1662,N_14554,N_11820);
and UO_1663 (O_1663,N_14381,N_12754);
nand UO_1664 (O_1664,N_10154,N_10958);
xor UO_1665 (O_1665,N_12353,N_11499);
and UO_1666 (O_1666,N_10800,N_11485);
and UO_1667 (O_1667,N_11512,N_12619);
nand UO_1668 (O_1668,N_13205,N_11307);
nor UO_1669 (O_1669,N_14930,N_14576);
nand UO_1670 (O_1670,N_12461,N_11511);
nor UO_1671 (O_1671,N_12807,N_10211);
and UO_1672 (O_1672,N_14011,N_12107);
nand UO_1673 (O_1673,N_10676,N_12031);
nor UO_1674 (O_1674,N_12459,N_12569);
nor UO_1675 (O_1675,N_10230,N_13045);
nand UO_1676 (O_1676,N_14532,N_14335);
or UO_1677 (O_1677,N_14972,N_14034);
and UO_1678 (O_1678,N_12702,N_14993);
nand UO_1679 (O_1679,N_14770,N_11440);
nand UO_1680 (O_1680,N_14703,N_11578);
or UO_1681 (O_1681,N_14268,N_13570);
nor UO_1682 (O_1682,N_14480,N_12731);
nor UO_1683 (O_1683,N_10807,N_12864);
nor UO_1684 (O_1684,N_12735,N_14891);
xor UO_1685 (O_1685,N_14719,N_12653);
xor UO_1686 (O_1686,N_10380,N_14878);
nand UO_1687 (O_1687,N_13788,N_11242);
nand UO_1688 (O_1688,N_11945,N_12364);
xnor UO_1689 (O_1689,N_13192,N_11950);
xor UO_1690 (O_1690,N_10571,N_13558);
and UO_1691 (O_1691,N_12577,N_13487);
nand UO_1692 (O_1692,N_11694,N_12100);
or UO_1693 (O_1693,N_14935,N_12155);
nor UO_1694 (O_1694,N_13985,N_12764);
and UO_1695 (O_1695,N_11753,N_10171);
or UO_1696 (O_1696,N_14967,N_10261);
or UO_1697 (O_1697,N_13974,N_14108);
nand UO_1698 (O_1698,N_10523,N_10803);
nor UO_1699 (O_1699,N_11839,N_11563);
and UO_1700 (O_1700,N_11049,N_13436);
xnor UO_1701 (O_1701,N_11240,N_13608);
or UO_1702 (O_1702,N_11142,N_11926);
nand UO_1703 (O_1703,N_13661,N_13362);
or UO_1704 (O_1704,N_11423,N_14934);
xnor UO_1705 (O_1705,N_12704,N_10250);
nor UO_1706 (O_1706,N_12730,N_10436);
nor UO_1707 (O_1707,N_14792,N_13542);
nor UO_1708 (O_1708,N_14202,N_11254);
and UO_1709 (O_1709,N_12138,N_12602);
nand UO_1710 (O_1710,N_14870,N_13869);
or UO_1711 (O_1711,N_10198,N_14504);
xor UO_1712 (O_1712,N_14102,N_14763);
xnor UO_1713 (O_1713,N_10659,N_11286);
nand UO_1714 (O_1714,N_10740,N_13153);
or UO_1715 (O_1715,N_11976,N_11751);
nand UO_1716 (O_1716,N_12305,N_14904);
and UO_1717 (O_1717,N_11793,N_12786);
nand UO_1718 (O_1718,N_12081,N_13553);
nand UO_1719 (O_1719,N_10931,N_10989);
nor UO_1720 (O_1720,N_12316,N_13513);
xor UO_1721 (O_1721,N_10802,N_14404);
nand UO_1722 (O_1722,N_14643,N_14181);
or UO_1723 (O_1723,N_10039,N_13096);
or UO_1724 (O_1724,N_11874,N_11236);
nor UO_1725 (O_1725,N_10528,N_14806);
nor UO_1726 (O_1726,N_12382,N_11824);
or UO_1727 (O_1727,N_13030,N_12168);
and UO_1728 (O_1728,N_14793,N_10569);
or UO_1729 (O_1729,N_10033,N_12848);
or UO_1730 (O_1730,N_12345,N_14133);
and UO_1731 (O_1731,N_12952,N_14744);
or UO_1732 (O_1732,N_10763,N_12962);
and UO_1733 (O_1733,N_11385,N_11686);
nor UO_1734 (O_1734,N_10767,N_10060);
xor UO_1735 (O_1735,N_13285,N_10630);
nand UO_1736 (O_1736,N_14175,N_11434);
or UO_1737 (O_1737,N_13884,N_12494);
nand UO_1738 (O_1738,N_13900,N_11894);
nor UO_1739 (O_1739,N_14645,N_10005);
or UO_1740 (O_1740,N_10502,N_11636);
and UO_1741 (O_1741,N_11912,N_13115);
or UO_1742 (O_1742,N_13765,N_14947);
and UO_1743 (O_1743,N_10017,N_11732);
nor UO_1744 (O_1744,N_11216,N_14860);
or UO_1745 (O_1745,N_13757,N_13503);
nand UO_1746 (O_1746,N_13218,N_10955);
nand UO_1747 (O_1747,N_14214,N_12824);
nor UO_1748 (O_1748,N_11416,N_11092);
and UO_1749 (O_1749,N_10339,N_14617);
and UO_1750 (O_1750,N_13422,N_10722);
nand UO_1751 (O_1751,N_12165,N_13891);
nand UO_1752 (O_1752,N_14252,N_10699);
and UO_1753 (O_1753,N_10879,N_11060);
or UO_1754 (O_1754,N_13344,N_12782);
or UO_1755 (O_1755,N_11070,N_13089);
nand UO_1756 (O_1756,N_14255,N_13821);
nor UO_1757 (O_1757,N_11163,N_13361);
nor UO_1758 (O_1758,N_13182,N_13790);
or UO_1759 (O_1759,N_11443,N_10038);
and UO_1760 (O_1760,N_10466,N_12118);
nor UO_1761 (O_1761,N_14472,N_11583);
nor UO_1762 (O_1762,N_12497,N_10069);
nor UO_1763 (O_1763,N_11508,N_13191);
and UO_1764 (O_1764,N_10231,N_14418);
or UO_1765 (O_1765,N_13594,N_13984);
or UO_1766 (O_1766,N_12846,N_14398);
and UO_1767 (O_1767,N_10011,N_11127);
nor UO_1768 (O_1768,N_11373,N_12534);
or UO_1769 (O_1769,N_12637,N_10377);
and UO_1770 (O_1770,N_13938,N_14674);
nand UO_1771 (O_1771,N_13289,N_13305);
and UO_1772 (O_1772,N_13539,N_10161);
nand UO_1773 (O_1773,N_11556,N_13704);
and UO_1774 (O_1774,N_12946,N_14387);
nor UO_1775 (O_1775,N_12341,N_13881);
nand UO_1776 (O_1776,N_10418,N_13483);
nand UO_1777 (O_1777,N_12805,N_11705);
or UO_1778 (O_1778,N_12996,N_13948);
or UO_1779 (O_1779,N_13287,N_11460);
nand UO_1780 (O_1780,N_10185,N_14562);
and UO_1781 (O_1781,N_14459,N_13896);
nor UO_1782 (O_1782,N_12513,N_13426);
or UO_1783 (O_1783,N_12798,N_14767);
or UO_1784 (O_1784,N_11086,N_13199);
or UO_1785 (O_1785,N_14230,N_14191);
nand UO_1786 (O_1786,N_13121,N_14771);
and UO_1787 (O_1787,N_12879,N_13946);
and UO_1788 (O_1788,N_13204,N_12103);
nand UO_1789 (O_1789,N_14447,N_12889);
xnor UO_1790 (O_1790,N_14091,N_10397);
xor UO_1791 (O_1791,N_12572,N_13409);
nand UO_1792 (O_1792,N_13489,N_11162);
or UO_1793 (O_1793,N_11591,N_12208);
or UO_1794 (O_1794,N_14624,N_10584);
or UO_1795 (O_1795,N_12217,N_14525);
or UO_1796 (O_1796,N_13978,N_14621);
or UO_1797 (O_1797,N_10559,N_14416);
or UO_1798 (O_1798,N_11546,N_14585);
nor UO_1799 (O_1799,N_12528,N_12164);
and UO_1800 (O_1800,N_14888,N_12077);
nor UO_1801 (O_1801,N_10479,N_14325);
nor UO_1802 (O_1802,N_11929,N_12181);
and UO_1803 (O_1803,N_12350,N_14808);
xnor UO_1804 (O_1804,N_10319,N_11626);
and UO_1805 (O_1805,N_12087,N_11513);
and UO_1806 (O_1806,N_10992,N_10507);
or UO_1807 (O_1807,N_10550,N_11516);
and UO_1808 (O_1808,N_11953,N_12643);
and UO_1809 (O_1809,N_13263,N_11590);
and UO_1810 (O_1810,N_11979,N_14347);
and UO_1811 (O_1811,N_10779,N_11818);
and UO_1812 (O_1812,N_11980,N_10260);
nand UO_1813 (O_1813,N_12929,N_11684);
or UO_1814 (O_1814,N_14663,N_12712);
and UO_1815 (O_1815,N_10072,N_10414);
or UO_1816 (O_1816,N_14424,N_10572);
or UO_1817 (O_1817,N_11298,N_13257);
nand UO_1818 (O_1818,N_11917,N_14420);
nand UO_1819 (O_1819,N_13007,N_10781);
and UO_1820 (O_1820,N_12861,N_10716);
nand UO_1821 (O_1821,N_10912,N_12766);
nor UO_1822 (O_1822,N_14316,N_11181);
nand UO_1823 (O_1823,N_11051,N_10579);
or UO_1824 (O_1824,N_14873,N_10094);
nand UO_1825 (O_1825,N_11258,N_10917);
or UO_1826 (O_1826,N_13926,N_13843);
nand UO_1827 (O_1827,N_13295,N_10947);
nor UO_1828 (O_1828,N_14650,N_11387);
xnor UO_1829 (O_1829,N_13245,N_13375);
nor UO_1830 (O_1830,N_14569,N_14714);
or UO_1831 (O_1831,N_11291,N_12508);
and UO_1832 (O_1832,N_10417,N_11275);
xnor UO_1833 (O_1833,N_12942,N_12654);
nor UO_1834 (O_1834,N_10666,N_14828);
nand UO_1835 (O_1835,N_14282,N_10191);
and UO_1836 (O_1836,N_10110,N_10828);
and UO_1837 (O_1837,N_14515,N_11859);
nand UO_1838 (O_1838,N_11302,N_10070);
nand UO_1839 (O_1839,N_11153,N_12410);
and UO_1840 (O_1840,N_10401,N_10712);
nor UO_1841 (O_1841,N_14074,N_14566);
and UO_1842 (O_1842,N_10810,N_13705);
or UO_1843 (O_1843,N_10888,N_12098);
and UO_1844 (O_1844,N_13463,N_13606);
or UO_1845 (O_1845,N_13615,N_11019);
nor UO_1846 (O_1846,N_11595,N_10691);
nor UO_1847 (O_1847,N_11031,N_11646);
and UO_1848 (O_1848,N_10074,N_13078);
nand UO_1849 (O_1849,N_13744,N_13652);
nor UO_1850 (O_1850,N_13898,N_14529);
nor UO_1851 (O_1851,N_10898,N_12667);
nor UO_1852 (O_1852,N_11599,N_13060);
nand UO_1853 (O_1853,N_11077,N_13358);
and UO_1854 (O_1854,N_14661,N_14134);
nand UO_1855 (O_1855,N_13840,N_12094);
nand UO_1856 (O_1856,N_10890,N_14158);
or UO_1857 (O_1857,N_14858,N_10517);
and UO_1858 (O_1858,N_11061,N_13308);
or UO_1859 (O_1859,N_13846,N_13155);
xnor UO_1860 (O_1860,N_14277,N_13644);
nor UO_1861 (O_1861,N_10750,N_11429);
nand UO_1862 (O_1862,N_11672,N_13724);
and UO_1863 (O_1863,N_10257,N_10219);
or UO_1864 (O_1864,N_13962,N_11211);
xor UO_1865 (O_1865,N_14477,N_13290);
and UO_1866 (O_1866,N_10116,N_13779);
nor UO_1867 (O_1867,N_14231,N_13646);
or UO_1868 (O_1868,N_13213,N_13024);
xor UO_1869 (O_1869,N_11263,N_13073);
nand UO_1870 (O_1870,N_10830,N_11073);
and UO_1871 (O_1871,N_11034,N_13369);
nand UO_1872 (O_1872,N_10822,N_12291);
nand UO_1873 (O_1873,N_11176,N_14353);
xor UO_1874 (O_1874,N_14653,N_14558);
nand UO_1875 (O_1875,N_10900,N_10538);
nand UO_1876 (O_1876,N_10745,N_10395);
or UO_1877 (O_1877,N_11860,N_12453);
nor UO_1878 (O_1878,N_12119,N_12359);
and UO_1879 (O_1879,N_12656,N_14292);
or UO_1880 (O_1880,N_12302,N_11566);
xor UO_1881 (O_1881,N_12280,N_12635);
nand UO_1882 (O_1882,N_14385,N_11608);
xor UO_1883 (O_1883,N_10846,N_14920);
and UO_1884 (O_1884,N_14302,N_13232);
and UO_1885 (O_1885,N_13267,N_14318);
nand UO_1886 (O_1886,N_10731,N_13510);
nor UO_1887 (O_1887,N_12938,N_10457);
and UO_1888 (O_1888,N_11584,N_13734);
and UO_1889 (O_1889,N_12362,N_12075);
nor UO_1890 (O_1890,N_12894,N_14551);
and UO_1891 (O_1891,N_11214,N_10452);
and UO_1892 (O_1892,N_11794,N_12986);
or UO_1893 (O_1893,N_10511,N_13472);
nor UO_1894 (O_1894,N_12469,N_13180);
nand UO_1895 (O_1895,N_14201,N_11455);
or UO_1896 (O_1896,N_11351,N_10656);
or UO_1897 (O_1897,N_10540,N_10168);
or UO_1898 (O_1898,N_12681,N_11807);
nor UO_1899 (O_1899,N_13322,N_10303);
or UO_1900 (O_1900,N_11647,N_13238);
and UO_1901 (O_1901,N_12334,N_10845);
or UO_1902 (O_1902,N_10620,N_11921);
xnor UO_1903 (O_1903,N_10848,N_12180);
and UO_1904 (O_1904,N_11995,N_10868);
or UO_1905 (O_1905,N_12612,N_13713);
or UO_1906 (O_1906,N_14874,N_13179);
and UO_1907 (O_1907,N_11406,N_11510);
and UO_1908 (O_1908,N_10467,N_14531);
xor UO_1909 (O_1909,N_10158,N_12112);
nand UO_1910 (O_1910,N_12556,N_11480);
or UO_1911 (O_1911,N_12485,N_10856);
nor UO_1912 (O_1912,N_13868,N_13140);
nor UO_1913 (O_1913,N_12358,N_12516);
and UO_1914 (O_1914,N_11961,N_10957);
nor UO_1915 (O_1915,N_12435,N_11754);
or UO_1916 (O_1916,N_11300,N_11261);
or UO_1917 (O_1917,N_10086,N_10626);
and UO_1918 (O_1918,N_13490,N_10826);
or UO_1919 (O_1919,N_10440,N_11380);
nor UO_1920 (O_1920,N_12196,N_13072);
nor UO_1921 (O_1921,N_10593,N_10776);
nand UO_1922 (O_1922,N_11143,N_11574);
nand UO_1923 (O_1923,N_13657,N_14769);
nor UO_1924 (O_1924,N_11308,N_12526);
nor UO_1925 (O_1925,N_11117,N_12420);
nor UO_1926 (O_1926,N_13571,N_14294);
nand UO_1927 (O_1927,N_13450,N_14951);
nor UO_1928 (O_1928,N_10176,N_12136);
nor UO_1929 (O_1929,N_12236,N_13723);
or UO_1930 (O_1930,N_11109,N_12761);
nand UO_1931 (O_1931,N_13825,N_11712);
nand UO_1932 (O_1932,N_14070,N_13476);
and UO_1933 (O_1933,N_12253,N_11495);
nor UO_1934 (O_1934,N_12166,N_11255);
or UO_1935 (O_1935,N_12908,N_10544);
nand UO_1936 (O_1936,N_14363,N_14825);
and UO_1937 (O_1937,N_12745,N_10429);
nand UO_1938 (O_1938,N_13953,N_12206);
or UO_1939 (O_1939,N_13206,N_13481);
and UO_1940 (O_1940,N_10349,N_10281);
xnor UO_1941 (O_1941,N_11782,N_10326);
and UO_1942 (O_1942,N_10983,N_10775);
or UO_1943 (O_1943,N_13665,N_10692);
or UO_1944 (O_1944,N_11892,N_12071);
or UO_1945 (O_1945,N_10996,N_14678);
and UO_1946 (O_1946,N_13586,N_11915);
nor UO_1947 (O_1947,N_13994,N_11553);
nor UO_1948 (O_1948,N_13972,N_10078);
nand UO_1949 (O_1949,N_13043,N_12467);
xnor UO_1950 (O_1950,N_12403,N_10755);
and UO_1951 (O_1951,N_10697,N_12427);
nor UO_1952 (O_1952,N_13321,N_14195);
xor UO_1953 (O_1953,N_11971,N_12587);
nand UO_1954 (O_1954,N_14361,N_13139);
xor UO_1955 (O_1955,N_12421,N_14994);
nor UO_1956 (O_1956,N_13244,N_10968);
and UO_1957 (O_1957,N_12685,N_13039);
or UO_1958 (O_1958,N_12099,N_13507);
nand UO_1959 (O_1959,N_12259,N_14431);
nor UO_1960 (O_1960,N_14209,N_10899);
nand UO_1961 (O_1961,N_11456,N_12939);
or UO_1962 (O_1962,N_11405,N_10241);
and UO_1963 (O_1963,N_10194,N_14957);
nand UO_1964 (O_1964,N_13872,N_10741);
nand UO_1965 (O_1965,N_14178,N_13067);
and UO_1966 (O_1966,N_13845,N_13684);
nor UO_1967 (O_1967,N_10987,N_14328);
and UO_1968 (O_1968,N_14590,N_14169);
xnor UO_1969 (O_1969,N_14053,N_11150);
nor UO_1970 (O_1970,N_10832,N_13172);
nand UO_1971 (O_1971,N_12527,N_13524);
and UO_1972 (O_1972,N_12481,N_11021);
nor UO_1973 (O_1973,N_14642,N_14709);
nor UO_1974 (O_1974,N_11177,N_12153);
nor UO_1975 (O_1975,N_13778,N_13856);
and UO_1976 (O_1976,N_10940,N_11920);
or UO_1977 (O_1977,N_12349,N_13956);
nand UO_1978 (O_1978,N_10713,N_13609);
or UO_1979 (O_1979,N_12371,N_13645);
or UO_1980 (O_1980,N_12387,N_10309);
nand UO_1981 (O_1981,N_13035,N_11223);
nor UO_1982 (O_1982,N_10396,N_10435);
nand UO_1983 (O_1983,N_10328,N_12139);
and UO_1984 (O_1984,N_13468,N_10105);
and UO_1985 (O_1985,N_12613,N_14662);
xnor UO_1986 (O_1986,N_11829,N_14841);
and UO_1987 (O_1987,N_14822,N_14109);
nand UO_1988 (O_1988,N_14740,N_10696);
or UO_1989 (O_1989,N_10008,N_13183);
and UO_1990 (O_1990,N_13725,N_13441);
xor UO_1991 (O_1991,N_14634,N_14950);
nand UO_1992 (O_1992,N_11534,N_12536);
and UO_1993 (O_1993,N_14519,N_10773);
xnor UO_1994 (O_1994,N_13275,N_10643);
or UO_1995 (O_1995,N_14583,N_13106);
or UO_1996 (O_1996,N_14412,N_12650);
xnor UO_1997 (O_1997,N_12642,N_13798);
nand UO_1998 (O_1998,N_13062,N_11414);
nand UO_1999 (O_1999,N_10301,N_13711);
endmodule