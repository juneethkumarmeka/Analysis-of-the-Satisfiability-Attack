module basic_1500_15000_2000_100_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_32,In_126);
or U1 (N_1,In_288,In_1181);
xor U2 (N_2,In_1383,In_563);
xor U3 (N_3,In_624,In_103);
nand U4 (N_4,In_138,In_1173);
or U5 (N_5,In_53,In_130);
xnor U6 (N_6,In_210,In_300);
nor U7 (N_7,In_964,In_823);
or U8 (N_8,In_1315,In_856);
or U9 (N_9,In_749,In_482);
nor U10 (N_10,In_453,In_144);
nand U11 (N_11,In_294,In_943);
and U12 (N_12,In_717,In_618);
and U13 (N_13,In_1276,In_744);
or U14 (N_14,In_109,In_837);
nand U15 (N_15,In_814,In_617);
and U16 (N_16,In_1443,In_861);
nand U17 (N_17,In_44,In_1079);
and U18 (N_18,In_1297,In_683);
nor U19 (N_19,In_90,In_1103);
xnor U20 (N_20,In_1037,In_732);
nor U21 (N_21,In_451,In_1038);
nand U22 (N_22,In_894,In_438);
nor U23 (N_23,In_1180,In_656);
nand U24 (N_24,In_984,In_1040);
and U25 (N_25,In_1302,In_1339);
or U26 (N_26,In_1005,In_1417);
or U27 (N_27,In_1430,In_501);
xnor U28 (N_28,In_755,In_63);
nand U29 (N_29,In_860,In_1406);
and U30 (N_30,In_918,In_845);
and U31 (N_31,In_958,In_157);
or U32 (N_32,In_784,In_672);
nor U33 (N_33,In_296,In_1027);
and U34 (N_34,In_1404,In_605);
xnor U35 (N_35,In_1244,In_390);
nand U36 (N_36,In_1022,In_415);
xor U37 (N_37,In_594,In_123);
and U38 (N_38,In_1481,In_599);
and U39 (N_39,In_416,In_88);
or U40 (N_40,In_245,In_951);
or U41 (N_41,In_893,In_1014);
xor U42 (N_42,In_1301,In_1015);
xnor U43 (N_43,In_364,In_566);
nand U44 (N_44,In_1168,In_848);
xnor U45 (N_45,In_237,In_897);
xor U46 (N_46,In_378,In_332);
xnor U47 (N_47,In_1496,In_1405);
and U48 (N_48,In_214,In_1092);
and U49 (N_49,In_602,In_1444);
or U50 (N_50,In_831,In_1207);
or U51 (N_51,In_1255,In_388);
and U52 (N_52,In_734,In_906);
nand U53 (N_53,In_968,In_211);
nor U54 (N_54,In_525,In_61);
or U55 (N_55,In_440,In_112);
xor U56 (N_56,In_302,In_1165);
nand U57 (N_57,In_1157,In_1493);
and U58 (N_58,In_878,In_881);
nor U59 (N_59,In_649,In_79);
xor U60 (N_60,In_354,In_763);
nor U61 (N_61,In_785,In_1139);
and U62 (N_62,In_1019,In_1296);
xnor U63 (N_63,In_1273,In_475);
xor U64 (N_64,In_1119,In_1312);
and U65 (N_65,In_427,In_338);
nor U66 (N_66,In_236,In_1064);
nand U67 (N_67,In_853,In_570);
and U68 (N_68,In_373,In_932);
nand U69 (N_69,In_419,In_244);
or U70 (N_70,In_804,In_162);
or U71 (N_71,In_1003,In_585);
nand U72 (N_72,In_205,In_1412);
xor U73 (N_73,In_69,In_486);
nand U74 (N_74,In_1020,In_1024);
and U75 (N_75,In_885,In_838);
nand U76 (N_76,In_177,In_406);
and U77 (N_77,In_640,In_658);
nor U78 (N_78,In_587,In_43);
nor U79 (N_79,In_39,In_231);
nor U80 (N_80,In_1182,In_912);
or U81 (N_81,In_914,In_521);
or U82 (N_82,In_456,In_1216);
nand U83 (N_83,In_1466,In_1378);
nand U84 (N_84,In_13,In_1099);
nand U85 (N_85,In_1490,In_619);
xnor U86 (N_86,In_20,In_926);
xnor U87 (N_87,In_645,In_1475);
or U88 (N_88,In_414,In_197);
or U89 (N_89,In_8,In_956);
nor U90 (N_90,In_1470,In_361);
or U91 (N_91,In_212,In_1056);
nor U92 (N_92,In_1042,In_1329);
nand U93 (N_93,In_1460,In_1367);
or U94 (N_94,In_1425,In_407);
xnor U95 (N_95,In_685,In_310);
nor U96 (N_96,In_439,In_864);
nand U97 (N_97,In_994,In_622);
and U98 (N_98,In_1049,In_91);
xnor U99 (N_99,In_304,In_1034);
nor U100 (N_100,In_815,In_1159);
nor U101 (N_101,In_124,In_345);
or U102 (N_102,In_1243,In_792);
and U103 (N_103,In_224,In_835);
nand U104 (N_104,In_836,In_1130);
xnor U105 (N_105,In_616,In_1433);
or U106 (N_106,In_1375,In_106);
and U107 (N_107,In_1438,In_1007);
and U108 (N_108,In_735,In_972);
and U109 (N_109,In_319,In_134);
and U110 (N_110,In_1010,In_148);
and U111 (N_111,In_1121,In_1374);
xnor U112 (N_112,In_242,In_195);
and U113 (N_113,In_203,In_676);
xnor U114 (N_114,In_494,In_1437);
nand U115 (N_115,In_27,In_1285);
xor U116 (N_116,In_1091,In_1381);
xnor U117 (N_117,In_1318,In_1472);
xnor U118 (N_118,In_983,In_557);
or U119 (N_119,In_297,In_28);
and U120 (N_120,In_259,In_510);
or U121 (N_121,In_396,In_1222);
nor U122 (N_122,In_322,In_1150);
or U123 (N_123,In_1424,In_1449);
or U124 (N_124,In_905,In_1248);
or U125 (N_125,In_324,In_398);
or U126 (N_126,In_1123,In_1429);
xnor U127 (N_127,In_712,In_953);
nor U128 (N_128,In_255,In_1242);
nand U129 (N_129,In_1464,In_1175);
and U130 (N_130,In_272,In_603);
and U131 (N_131,In_1454,In_583);
xnor U132 (N_132,In_800,In_397);
xor U133 (N_133,In_668,In_198);
or U134 (N_134,In_466,In_1304);
nand U135 (N_135,In_329,In_1346);
or U136 (N_136,In_1484,In_961);
nand U137 (N_137,In_1125,In_331);
or U138 (N_138,In_169,In_522);
nand U139 (N_139,In_1084,In_1256);
xor U140 (N_140,In_1253,In_1356);
xor U141 (N_141,In_209,In_377);
xnor U142 (N_142,In_1317,In_42);
and U143 (N_143,In_761,In_651);
nand U144 (N_144,In_988,In_796);
nor U145 (N_145,In_1044,In_1131);
nand U146 (N_146,In_110,In_751);
xor U147 (N_147,In_457,In_292);
xor U148 (N_148,In_430,In_1167);
nor U149 (N_149,In_908,In_1118);
nand U150 (N_150,In_748,In_21);
and U151 (N_151,N_110,In_479);
and U152 (N_152,In_524,In_62);
nor U153 (N_153,N_65,In_1314);
xnor U154 (N_154,In_353,In_37);
xnor U155 (N_155,In_253,N_2);
nand U156 (N_156,N_5,In_520);
nand U157 (N_157,In_218,In_386);
and U158 (N_158,In_1432,In_379);
or U159 (N_159,In_978,In_334);
and U160 (N_160,In_318,In_340);
or U161 (N_161,In_1266,In_1178);
or U162 (N_162,In_715,In_516);
or U163 (N_163,In_172,In_426);
and U164 (N_164,In_807,In_706);
and U165 (N_165,In_802,In_1499);
and U166 (N_166,In_1,In_995);
xnor U167 (N_167,In_1476,In_1197);
or U168 (N_168,In_560,In_281);
nor U169 (N_169,In_10,In_987);
xnor U170 (N_170,In_896,In_703);
and U171 (N_171,In_963,In_847);
nor U172 (N_172,In_190,In_1219);
nor U173 (N_173,In_1498,In_938);
and U174 (N_174,In_597,In_179);
and U175 (N_175,In_278,In_1043);
nand U176 (N_176,In_1284,In_1202);
xor U177 (N_177,In_173,In_1280);
nor U178 (N_178,In_258,In_1174);
xnor U179 (N_179,In_871,In_113);
nor U180 (N_180,In_684,N_116);
xnor U181 (N_181,In_1110,In_194);
or U182 (N_182,In_70,In_1000);
nand U183 (N_183,In_1289,In_1148);
or U184 (N_184,In_97,In_316);
nand U185 (N_185,In_277,In_757);
xnor U186 (N_186,In_370,In_1458);
nor U187 (N_187,In_700,In_1013);
nor U188 (N_188,In_863,N_62);
or U189 (N_189,In_1385,In_1361);
and U190 (N_190,In_18,In_1436);
nor U191 (N_191,In_980,In_875);
xor U192 (N_192,In_1259,In_1446);
and U193 (N_193,In_753,In_382);
nor U194 (N_194,In_1495,In_1392);
xor U195 (N_195,In_1387,In_787);
nor U196 (N_196,In_727,In_678);
xnor U197 (N_197,In_1188,In_852);
nor U198 (N_198,N_32,In_682);
and U199 (N_199,In_16,In_652);
nand U200 (N_200,In_770,In_311);
xor U201 (N_201,In_901,N_106);
and U202 (N_202,In_844,In_608);
or U203 (N_203,In_1221,N_122);
nor U204 (N_204,In_38,In_1163);
xor U205 (N_205,In_1154,In_478);
and U206 (N_206,N_102,N_142);
or U207 (N_207,In_1100,N_20);
nand U208 (N_208,In_745,In_517);
nand U209 (N_209,In_1334,In_546);
xnor U210 (N_210,In_632,In_363);
or U211 (N_211,In_202,In_946);
nor U212 (N_212,In_1113,In_58);
nor U213 (N_213,In_985,In_1347);
nor U214 (N_214,In_95,In_638);
xnor U215 (N_215,In_170,In_692);
nor U216 (N_216,In_154,In_1400);
xnor U217 (N_217,In_1184,In_455);
nand U218 (N_218,In_1105,In_358);
nand U219 (N_219,N_145,In_444);
or U220 (N_220,In_167,In_333);
xor U221 (N_221,In_1087,N_94);
nand U222 (N_222,In_40,In_343);
xnor U223 (N_223,In_376,In_1349);
or U224 (N_224,In_1135,In_428);
nor U225 (N_225,In_1360,In_164);
nor U226 (N_226,In_445,In_459);
xor U227 (N_227,N_22,In_1275);
and U228 (N_228,In_1068,In_1074);
or U229 (N_229,In_351,In_718);
nor U230 (N_230,In_556,In_1332);
nand U231 (N_231,In_1176,In_999);
xnor U232 (N_232,In_1377,In_653);
xor U233 (N_233,N_71,In_350);
or U234 (N_234,In_733,In_677);
nand U235 (N_235,In_1016,In_1048);
nor U236 (N_236,In_1257,In_634);
nor U237 (N_237,In_772,In_1127);
and U238 (N_238,In_403,N_45);
nor U239 (N_239,In_799,In_261);
or U240 (N_240,In_737,N_146);
xor U241 (N_241,In_35,In_1166);
nand U242 (N_242,In_232,In_468);
nor U243 (N_243,In_222,N_33);
nor U244 (N_244,In_591,In_1223);
or U245 (N_245,In_476,In_731);
or U246 (N_246,In_12,In_662);
xor U247 (N_247,In_1235,In_1201);
nor U248 (N_248,In_118,In_401);
and U249 (N_249,In_865,In_747);
and U250 (N_250,In_481,In_824);
or U251 (N_251,In_663,In_1316);
and U252 (N_252,In_565,In_492);
or U253 (N_253,N_128,In_1114);
or U254 (N_254,In_705,In_1250);
and U255 (N_255,In_564,N_53);
nor U256 (N_256,In_559,In_60);
nand U257 (N_257,N_126,In_1035);
xor U258 (N_258,In_1088,In_221);
xnor U259 (N_259,In_268,In_821);
or U260 (N_260,N_92,In_117);
or U261 (N_261,In_695,In_710);
and U262 (N_262,In_266,In_1463);
or U263 (N_263,N_86,In_1116);
or U264 (N_264,In_467,In_339);
and U265 (N_265,In_1149,In_1441);
nor U266 (N_266,In_1299,In_947);
or U267 (N_267,In_809,In_880);
and U268 (N_268,In_696,In_1109);
xor U269 (N_269,In_270,In_1211);
or U270 (N_270,In_1012,In_686);
and U271 (N_271,N_100,In_588);
nand U272 (N_272,In_1234,In_579);
nand U273 (N_273,In_568,In_1497);
or U274 (N_274,In_631,In_1155);
nand U275 (N_275,In_410,In_360);
nand U276 (N_276,In_889,In_85);
xnor U277 (N_277,In_1220,In_786);
or U278 (N_278,In_31,In_886);
and U279 (N_279,In_1473,In_771);
nor U280 (N_280,In_1058,In_129);
or U281 (N_281,In_1335,N_46);
or U282 (N_282,In_541,In_229);
nand U283 (N_283,In_491,In_1073);
and U284 (N_284,In_1342,N_105);
nand U285 (N_285,In_643,In_473);
xor U286 (N_286,In_1485,In_781);
or U287 (N_287,In_1214,In_1455);
and U288 (N_288,In_916,In_762);
or U289 (N_289,In_271,In_151);
and U290 (N_290,In_1144,In_470);
xor U291 (N_291,In_675,In_610);
or U292 (N_292,In_827,N_25);
or U293 (N_293,In_248,N_95);
nand U294 (N_294,In_741,In_709);
xnor U295 (N_295,In_829,In_1075);
nand U296 (N_296,In_1229,In_23);
nor U297 (N_297,In_82,In_1008);
or U298 (N_298,In_183,N_85);
nor U299 (N_299,In_295,In_573);
xnor U300 (N_300,In_145,In_1351);
or U301 (N_301,In_1295,In_93);
nand U302 (N_302,In_1230,In_65);
nor U303 (N_303,In_503,N_252);
nand U304 (N_304,N_236,In_1254);
nor U305 (N_305,In_56,In_1206);
and U306 (N_306,In_740,In_404);
nor U307 (N_307,N_83,In_1004);
xor U308 (N_308,In_1290,In_623);
nand U309 (N_309,N_179,In_1338);
xnor U310 (N_310,In_34,N_253);
nand U311 (N_311,In_1467,In_1002);
xnor U312 (N_312,N_123,In_974);
nor U313 (N_313,In_1423,In_891);
and U314 (N_314,In_1142,In_758);
or U315 (N_315,N_42,In_704);
nand U316 (N_316,In_1252,In_969);
or U317 (N_317,In_801,In_1479);
nor U318 (N_318,In_725,In_887);
nor U319 (N_319,In_1408,In_1122);
nand U320 (N_320,In_1399,In_738);
and U321 (N_321,In_511,In_857);
nor U322 (N_322,In_730,N_24);
or U323 (N_323,In_443,In_598);
and U324 (N_324,N_9,N_168);
and U325 (N_325,In_284,In_746);
and U326 (N_326,In_1245,In_869);
or U327 (N_327,N_220,In_321);
xor U328 (N_328,In_460,In_679);
nor U329 (N_329,In_1061,In_485);
nor U330 (N_330,In_1439,In_970);
xor U331 (N_331,N_255,In_776);
and U332 (N_332,In_674,In_250);
or U333 (N_333,In_646,In_55);
nor U334 (N_334,In_866,In_1205);
and U335 (N_335,In_447,In_25);
nor U336 (N_336,N_283,In_199);
nor U337 (N_337,In_1489,In_233);
and U338 (N_338,In_1369,In_760);
nor U339 (N_339,In_768,N_99);
nand U340 (N_340,In_842,In_508);
nor U341 (N_341,N_177,In_1321);
nand U342 (N_342,In_193,In_285);
and U343 (N_343,N_248,In_1161);
or U344 (N_344,In_904,N_166);
nor U345 (N_345,N_199,In_830);
nand U346 (N_346,In_323,In_775);
nand U347 (N_347,In_971,In_805);
and U348 (N_348,In_359,In_317);
nor U349 (N_349,In_1054,In_1162);
nand U350 (N_350,In_693,In_773);
and U351 (N_351,In_1066,In_385);
nor U352 (N_352,In_538,In_895);
nor U353 (N_353,In_1104,N_90);
xnor U354 (N_354,N_29,In_888);
nand U355 (N_355,N_133,In_660);
or U356 (N_356,In_965,In_1160);
and U357 (N_357,In_1031,In_1151);
xnor U358 (N_358,N_41,In_346);
nor U359 (N_359,In_287,In_1419);
nor U360 (N_360,N_262,N_91);
and U361 (N_361,In_514,In_581);
xor U362 (N_362,In_701,In_265);
nand U363 (N_363,In_1281,N_205);
or U364 (N_364,In_92,In_1390);
nor U365 (N_365,In_589,In_1070);
nand U366 (N_366,N_55,In_1396);
nor U367 (N_367,In_5,In_264);
xor U368 (N_368,N_185,In_902);
nand U369 (N_369,In_1124,N_31);
xnor U370 (N_370,N_160,N_290);
xor U371 (N_371,In_1210,In_882);
and U372 (N_372,In_697,In_647);
or U373 (N_373,N_233,In_384);
or U374 (N_374,In_1236,In_1358);
or U375 (N_375,N_72,In_979);
or U376 (N_376,In_924,In_724);
nor U377 (N_377,N_161,In_1021);
or U378 (N_378,In_14,N_15);
or U379 (N_379,In_555,N_230);
nand U380 (N_380,In_303,In_483);
xnor U381 (N_381,In_982,N_222);
xor U382 (N_382,In_158,In_873);
nand U383 (N_383,In_105,In_917);
nor U384 (N_384,In_267,N_203);
or U385 (N_385,In_862,In_1308);
nand U386 (N_386,N_190,N_260);
nor U387 (N_387,N_143,In_241);
or U388 (N_388,In_957,In_11);
nand U389 (N_389,In_436,N_132);
and U390 (N_390,N_70,N_98);
nand U391 (N_391,In_783,In_1364);
nor U392 (N_392,In_659,N_57);
or U393 (N_393,N_89,In_1132);
nor U394 (N_394,In_816,In_81);
and U395 (N_395,N_76,In_833);
nand U396 (N_396,In_68,In_1370);
or U397 (N_397,In_1327,In_1030);
and U398 (N_398,In_1409,In_506);
or U399 (N_399,In_17,In_1384);
and U400 (N_400,In_143,N_13);
nand U401 (N_401,In_1386,In_417);
nor U402 (N_402,N_1,In_1055);
nand U403 (N_403,In_174,In_490);
nand U404 (N_404,In_1143,In_1183);
nor U405 (N_405,In_422,In_642);
nand U406 (N_406,In_269,In_1133);
and U407 (N_407,In_1120,In_394);
nor U408 (N_408,In_368,In_235);
and U409 (N_409,N_279,In_477);
or U410 (N_410,In_448,In_769);
xor U411 (N_411,N_176,In_293);
or U412 (N_412,In_182,In_611);
nand U413 (N_413,In_919,In_797);
nand U414 (N_414,N_3,In_1486);
and U415 (N_415,N_271,In_1359);
or U416 (N_416,In_57,In_371);
nand U417 (N_417,N_266,In_1238);
and U418 (N_418,In_1270,N_104);
nand U419 (N_419,In_383,In_423);
and U420 (N_420,In_121,In_26);
and U421 (N_421,In_1146,N_112);
or U422 (N_422,N_239,N_23);
nor U423 (N_423,In_47,In_7);
or U424 (N_424,In_1213,In_99);
xor U425 (N_425,In_641,N_156);
and U426 (N_426,In_569,In_1089);
and U427 (N_427,N_163,In_185);
nand U428 (N_428,In_246,In_1106);
and U429 (N_429,In_1108,N_64);
nand U430 (N_430,In_462,In_180);
nand U431 (N_431,In_140,In_1413);
nand U432 (N_432,N_291,In_102);
xor U433 (N_433,N_6,In_22);
nor U434 (N_434,In_135,In_186);
nand U435 (N_435,In_960,N_294);
nand U436 (N_436,N_11,N_36);
and U437 (N_437,In_935,In_509);
and U438 (N_438,In_1366,In_89);
nand U439 (N_439,In_941,N_189);
and U440 (N_440,N_280,In_273);
nand U441 (N_441,In_247,In_561);
or U442 (N_442,In_975,In_1373);
and U443 (N_443,In_567,In_1264);
nor U444 (N_444,In_137,In_50);
nand U445 (N_445,In_592,N_38);
nand U446 (N_446,In_469,N_149);
nand U447 (N_447,In_290,In_874);
nor U448 (N_448,In_45,In_257);
nand U449 (N_449,In_1465,In_83);
and U450 (N_450,In_791,In_997);
nand U451 (N_451,N_16,N_296);
xor U452 (N_452,In_1185,N_394);
nor U453 (N_453,N_117,N_347);
xnor U454 (N_454,In_119,In_621);
nand U455 (N_455,N_272,In_480);
or U456 (N_456,In_513,In_149);
or U457 (N_457,N_427,In_849);
xor U458 (N_458,In_547,In_1028);
and U459 (N_459,N_162,In_615);
xnor U460 (N_460,In_774,In_1450);
and U461 (N_461,N_63,N_369);
or U462 (N_462,N_130,N_422);
nor U463 (N_463,In_6,N_115);
nand U464 (N_464,N_226,N_229);
xor U465 (N_465,In_936,In_533);
or U466 (N_466,In_1260,N_338);
nand U467 (N_467,In_155,In_1487);
xor U468 (N_468,N_224,In_1410);
nand U469 (N_469,In_1052,N_408);
xor U470 (N_470,In_165,In_530);
xnor U471 (N_471,N_155,In_29);
nor U472 (N_472,In_115,In_1324);
or U473 (N_473,In_713,In_1128);
nand U474 (N_474,In_1225,In_630);
or U475 (N_475,N_442,N_381);
nor U476 (N_476,In_1097,N_350);
nor U477 (N_477,In_1320,N_432);
or U478 (N_478,In_458,N_385);
nand U479 (N_479,In_519,In_518);
and U480 (N_480,N_147,In_1492);
or U481 (N_481,In_1363,In_661);
xnor U482 (N_482,N_259,In_367);
nor U483 (N_483,In_927,N_405);
nand U484 (N_484,In_408,In_851);
or U485 (N_485,N_274,In_1212);
nand U486 (N_486,In_806,N_169);
nand U487 (N_487,In_1083,N_12);
or U488 (N_488,N_52,In_1249);
nor U489 (N_489,N_180,In_314);
and U490 (N_490,In_1474,In_1469);
xor U491 (N_491,N_406,N_416);
nand U492 (N_492,In_798,In_959);
nand U493 (N_493,In_178,In_648);
nor U494 (N_494,In_254,In_381);
or U495 (N_495,In_215,N_302);
or U496 (N_496,In_1241,N_344);
nand U497 (N_497,N_412,In_702);
and U498 (N_498,In_1187,N_225);
xor U499 (N_499,N_358,In_1480);
nand U500 (N_500,In_545,In_217);
and U501 (N_501,N_299,N_66);
xor U502 (N_502,In_449,In_765);
or U503 (N_503,In_739,In_432);
or U504 (N_504,N_144,In_1102);
and U505 (N_505,In_1398,In_161);
xor U506 (N_506,N_295,N_251);
or U507 (N_507,In_1081,N_209);
and U508 (N_508,N_269,In_1305);
and U509 (N_509,In_1452,N_43);
and U510 (N_510,In_402,In_1397);
nand U511 (N_511,In_1426,N_327);
or U512 (N_512,In_107,In_282);
nand U513 (N_513,N_364,In_818);
nand U514 (N_514,In_418,In_542);
and U515 (N_515,N_325,N_215);
and U516 (N_516,In_1352,N_423);
nand U517 (N_517,In_962,N_127);
nor U518 (N_518,N_372,In_1263);
and U519 (N_519,In_1246,In_1231);
or U520 (N_520,N_228,In_1372);
xor U521 (N_521,In_750,In_471);
nand U522 (N_522,In_1388,In_41);
nand U523 (N_523,N_310,N_232);
nor U524 (N_524,N_240,In_990);
xnor U525 (N_525,In_301,In_613);
nor U526 (N_526,In_1494,N_390);
xor U527 (N_527,N_437,In_858);
or U528 (N_528,In_101,In_812);
nand U529 (N_529,N_194,N_159);
nand U530 (N_530,In_76,In_71);
and U531 (N_531,In_393,In_1448);
and U532 (N_532,N_19,In_527);
nand U533 (N_533,N_324,N_7);
or U534 (N_534,N_433,In_944);
nand U535 (N_535,In_1138,N_170);
or U536 (N_536,In_832,N_108);
nand U537 (N_537,N_289,In_1033);
nand U538 (N_538,N_332,In_1310);
nand U539 (N_539,In_1411,In_694);
and U540 (N_540,In_335,N_241);
nor U541 (N_541,In_132,In_1224);
or U542 (N_542,In_991,In_817);
nand U543 (N_543,In_1189,N_107);
and U544 (N_544,N_88,In_900);
nand U545 (N_545,In_722,N_387);
xor U546 (N_546,In_1483,N_111);
xnor U547 (N_547,In_276,N_319);
nand U548 (N_548,In_689,N_443);
or U549 (N_549,In_843,N_244);
nand U550 (N_550,In_488,In_1233);
nand U551 (N_551,In_1306,In_855);
nand U552 (N_552,N_403,In_450);
nor U553 (N_553,In_1442,In_1403);
nand U554 (N_554,N_449,In_1422);
and U555 (N_555,N_335,In_586);
nand U556 (N_556,In_1071,In_779);
and U557 (N_557,In_1247,In_411);
or U558 (N_558,In_434,N_311);
and U559 (N_559,In_472,In_220);
nand U560 (N_560,In_1440,In_374);
nor U561 (N_561,N_349,In_1001);
nor U562 (N_562,N_277,In_505);
xor U563 (N_563,In_1090,In_601);
or U564 (N_564,In_391,N_197);
nand U565 (N_565,In_1076,In_1357);
and U566 (N_566,In_726,N_309);
or U567 (N_567,In_620,In_1313);
and U568 (N_568,In_780,N_401);
and U569 (N_569,N_300,N_368);
or U570 (N_570,N_447,In_915);
xnor U571 (N_571,In_1158,In_910);
and U572 (N_572,In_307,In_854);
and U573 (N_573,N_188,In_120);
nand U574 (N_574,In_1190,In_299);
or U575 (N_575,In_1156,In_206);
xnor U576 (N_576,In_352,In_1177);
and U577 (N_577,N_0,N_125);
nand U578 (N_578,In_949,In_551);
nand U579 (N_579,N_264,In_24);
nand U580 (N_580,In_1186,In_1268);
nand U581 (N_581,In_841,N_249);
xor U582 (N_582,N_201,In_1298);
nand U583 (N_583,In_1191,N_17);
nand U584 (N_584,In_1307,N_184);
or U585 (N_585,In_1343,In_921);
and U586 (N_586,N_389,In_1111);
nand U587 (N_587,In_1291,In_1060);
or U588 (N_588,In_998,In_1193);
xnor U589 (N_589,N_56,In_948);
or U590 (N_590,N_247,In_1488);
or U591 (N_591,In_1228,In_934);
nand U592 (N_592,N_352,N_420);
and U593 (N_593,In_548,In_1407);
and U594 (N_594,In_312,In_64);
and U595 (N_595,In_196,N_448);
nand U596 (N_596,In_654,In_614);
nor U597 (N_597,In_899,In_30);
nor U598 (N_598,In_104,In_1326);
or U599 (N_599,In_507,N_114);
or U600 (N_600,In_1451,N_515);
nand U601 (N_601,N_87,In_937);
and U602 (N_602,In_1428,N_285);
xnor U603 (N_603,In_252,N_207);
nand U604 (N_604,In_1353,N_541);
and U605 (N_605,In_657,N_577);
nor U606 (N_606,N_59,In_719);
xor U607 (N_607,In_399,In_1368);
or U608 (N_608,In_515,N_131);
xnor U609 (N_609,In_156,In_441);
nand U610 (N_610,In_1414,In_680);
xor U611 (N_611,N_273,In_256);
nor U612 (N_612,In_540,N_139);
nand U613 (N_613,N_418,In_989);
nor U614 (N_614,N_370,In_1094);
xor U615 (N_615,N_383,In_1269);
nor U616 (N_616,N_113,N_424);
xnor U617 (N_617,In_208,In_766);
or U618 (N_618,N_473,N_526);
nand U619 (N_619,In_1379,N_554);
nor U620 (N_620,In_1331,N_235);
xnor U621 (N_621,In_1420,In_1072);
nand U622 (N_622,In_493,N_597);
and U623 (N_623,In_1086,N_44);
or U624 (N_624,In_1267,In_707);
nand U625 (N_625,In_1278,N_466);
nand U626 (N_626,In_133,In_72);
xor U627 (N_627,N_275,In_1457);
and U628 (N_628,N_297,In_239);
or U629 (N_629,In_1288,In_309);
and U630 (N_630,N_355,In_49);
nand U631 (N_631,N_246,N_79);
and U632 (N_632,In_1251,N_480);
xor U633 (N_633,N_292,N_154);
or U634 (N_634,N_588,N_396);
nand U635 (N_635,N_483,In_128);
and U636 (N_636,In_575,In_1279);
or U637 (N_637,N_21,In_337);
or U638 (N_638,N_238,In_859);
and U639 (N_639,N_216,In_52);
nor U640 (N_640,In_159,N_305);
xnor U641 (N_641,In_633,In_576);
xnor U642 (N_642,N_258,N_413);
and U643 (N_643,In_1355,N_500);
nand U644 (N_644,N_343,N_58);
and U645 (N_645,In_286,In_380);
and U646 (N_646,In_1401,N_376);
nor U647 (N_647,In_819,In_1371);
xnor U648 (N_648,In_1053,N_278);
nand U649 (N_649,In_187,In_2);
nand U650 (N_650,N_505,In_1340);
nand U651 (N_651,In_1200,N_587);
nor U652 (N_652,In_846,N_578);
or U653 (N_653,In_531,In_789);
nand U654 (N_654,In_298,N_499);
nand U655 (N_655,N_550,In_890);
xnor U656 (N_656,N_589,N_97);
or U657 (N_657,N_562,N_333);
nor U658 (N_658,In_1274,In_1478);
or U659 (N_659,In_839,N_470);
nor U660 (N_660,N_461,N_594);
or U661 (N_661,N_35,In_1218);
nor U662 (N_662,In_1491,In_986);
nor U663 (N_663,In_655,N_135);
xor U664 (N_664,N_479,In_803);
nand U665 (N_665,In_552,In_225);
xnor U666 (N_666,In_108,N_460);
nor U667 (N_667,N_459,In_1107);
xor U668 (N_668,N_212,N_213);
nor U669 (N_669,N_40,In_1322);
nand U670 (N_670,In_826,N_186);
and U671 (N_671,In_671,In_1018);
nor U672 (N_672,N_75,N_378);
and U673 (N_673,In_1431,In_1261);
xor U674 (N_674,N_164,In_1258);
nor U675 (N_675,In_498,N_231);
nand U676 (N_676,In_1101,N_60);
or U677 (N_677,N_458,In_1112);
nand U678 (N_678,In_142,N_476);
xnor U679 (N_679,In_1421,N_227);
nor U680 (N_680,In_176,N_439);
nor U681 (N_681,In_201,In_1391);
or U682 (N_682,In_238,N_129);
nor U683 (N_683,In_537,In_688);
xor U684 (N_684,In_356,In_1077);
and U685 (N_685,N_234,In_544);
xnor U686 (N_686,N_450,N_10);
nor U687 (N_687,In_928,In_141);
xor U688 (N_688,In_721,N_481);
nor U689 (N_689,N_267,N_535);
or U690 (N_690,N_357,In_365);
or U691 (N_691,In_504,N_560);
and U692 (N_692,In_499,In_283);
nor U693 (N_693,N_118,In_512);
nand U694 (N_694,In_536,N_573);
nand U695 (N_695,N_514,In_1325);
and U696 (N_696,In_67,N_263);
nand U697 (N_697,In_336,In_429);
xor U698 (N_698,N_322,In_1434);
nor U699 (N_699,In_868,N_429);
xor U700 (N_700,N_518,In_349);
or U701 (N_701,In_728,In_80);
nor U702 (N_702,N_441,N_493);
nor U703 (N_703,N_137,In_729);
or U704 (N_704,N_539,In_279);
nor U705 (N_705,In_1393,N_328);
or U706 (N_706,N_321,N_81);
xor U707 (N_707,In_474,In_595);
or U708 (N_708,N_377,N_326);
xnor U709 (N_709,N_542,In_1435);
and U710 (N_710,In_870,In_306);
nor U711 (N_711,In_1153,N_276);
nor U712 (N_712,N_482,N_206);
nor U713 (N_713,In_1286,In_670);
or U714 (N_714,In_1292,N_417);
nor U715 (N_715,N_286,In_1147);
or U716 (N_716,N_445,In_1382);
nand U717 (N_717,In_635,In_795);
xor U718 (N_718,N_152,N_566);
nand U719 (N_719,In_788,In_553);
or U720 (N_720,N_8,In_73);
nand U721 (N_721,In_903,In_883);
nor U722 (N_722,N_436,N_546);
and U723 (N_723,In_147,In_1350);
nor U724 (N_724,N_39,N_318);
nor U725 (N_725,In_1172,In_1416);
xor U726 (N_726,In_820,In_228);
or U727 (N_727,In_1395,In_572);
or U728 (N_728,In_940,In_1402);
nand U729 (N_729,N_313,N_457);
and U730 (N_730,In_1045,In_1262);
and U731 (N_731,In_627,N_580);
nand U732 (N_732,In_487,In_98);
nor U733 (N_733,N_477,In_681);
or U734 (N_734,In_146,In_395);
or U735 (N_735,In_528,N_84);
xnor U736 (N_736,N_487,In_362);
or U737 (N_737,N_517,N_153);
and U738 (N_738,In_939,In_240);
and U739 (N_739,In_1287,N_172);
nand U740 (N_740,N_558,N_419);
nor U741 (N_741,N_591,N_565);
nand U742 (N_742,In_1336,N_210);
and U743 (N_743,In_879,N_440);
nor U744 (N_744,N_485,In_1134);
nor U745 (N_745,In_234,In_86);
nor U746 (N_746,N_599,In_629);
and U747 (N_747,In_877,N_528);
nand U748 (N_748,In_1232,N_250);
xor U749 (N_749,N_221,In_66);
nor U750 (N_750,N_124,N_508);
and U751 (N_751,N_636,In_464);
xnor U752 (N_752,N_330,In_181);
nor U753 (N_753,N_261,In_184);
nor U754 (N_754,In_313,In_1080);
or U755 (N_755,N_93,N_467);
and U756 (N_756,N_682,N_486);
and U757 (N_757,N_362,N_576);
xnor U758 (N_758,In_1057,N_181);
nand U759 (N_759,In_420,N_421);
or U760 (N_760,In_1069,In_96);
xor U761 (N_761,N_724,In_759);
nand U762 (N_762,N_590,In_1098);
and U763 (N_763,N_635,N_30);
or U764 (N_764,N_4,In_1445);
nand U765 (N_765,In_163,In_644);
xnor U766 (N_766,In_171,In_810);
nor U767 (N_767,N_471,In_526);
or U768 (N_768,In_966,In_892);
or U769 (N_769,N_141,In_1380);
or U770 (N_770,In_1145,N_650);
and U771 (N_771,In_500,N_625);
and U772 (N_772,In_577,In_571);
nand U773 (N_773,N_684,In_19);
or U774 (N_774,N_603,In_973);
nor U775 (N_775,N_80,N_585);
xor U776 (N_776,In_263,N_749);
and U777 (N_777,N_384,N_699);
and U778 (N_778,N_257,N_121);
and U779 (N_779,N_495,N_654);
and U780 (N_780,In_558,N_444);
or U781 (N_781,In_767,N_497);
nand U782 (N_782,N_631,N_288);
xnor U783 (N_783,In_168,In_1239);
and U784 (N_784,In_192,N_637);
nor U785 (N_785,N_345,N_621);
or U786 (N_786,N_614,In_327);
nand U787 (N_787,In_930,N_407);
and U788 (N_788,N_672,In_922);
nor U789 (N_789,N_688,N_686);
xor U790 (N_790,In_1323,N_138);
nor U791 (N_791,N_346,In_280);
or U792 (N_792,N_592,In_850);
or U793 (N_793,In_976,N_559);
and U794 (N_794,N_506,In_125);
xnor U795 (N_795,In_1195,N_741);
nand U796 (N_796,N_678,N_191);
xor U797 (N_797,N_315,In_523);
nand U798 (N_798,In_945,In_1009);
and U799 (N_799,N_455,N_502);
xor U800 (N_800,N_37,In_1126);
and U801 (N_801,N_600,N_74);
nor U802 (N_802,N_648,In_46);
nand U803 (N_803,In_590,N_543);
or U804 (N_804,In_580,N_409);
nor U805 (N_805,N_312,In_687);
xnor U806 (N_806,N_134,N_520);
or U807 (N_807,N_217,In_977);
or U808 (N_808,N_464,N_398);
xnor U809 (N_809,In_1354,In_1215);
xnor U810 (N_810,In_36,N_469);
or U811 (N_811,N_649,In_1461);
and U812 (N_812,N_709,N_721);
and U813 (N_813,N_265,In_1217);
nand U814 (N_814,N_569,N_446);
xor U815 (N_815,N_610,N_54);
nand U816 (N_816,N_304,In_1011);
xnor U817 (N_817,In_549,In_778);
nor U818 (N_818,N_157,N_316);
nand U819 (N_819,In_75,N_193);
nand U820 (N_820,N_521,N_507);
xnor U821 (N_821,N_538,N_268);
nand U822 (N_822,N_659,In_1209);
nor U823 (N_823,In_1237,In_484);
nor U824 (N_824,N_703,N_737);
xnor U825 (N_825,N_681,In_325);
or U826 (N_826,In_754,N_548);
xnor U827 (N_827,N_651,N_697);
or U828 (N_828,In_1226,N_34);
xnor U829 (N_829,In_1169,N_687);
and U830 (N_830,N_339,N_732);
nor U831 (N_831,N_662,N_627);
and U832 (N_832,N_314,N_490);
xnor U833 (N_833,N_165,N_711);
nor U834 (N_834,In_328,N_671);
nor U835 (N_835,In_1047,N_622);
nand U836 (N_836,N_745,N_725);
nand U837 (N_837,N_611,N_642);
nand U838 (N_838,N_638,N_478);
or U839 (N_839,In_1137,N_151);
or U840 (N_840,In_1300,N_287);
or U841 (N_841,N_363,In_782);
nor U842 (N_842,N_204,N_103);
and U843 (N_843,N_382,In_1365);
or U844 (N_844,N_340,N_730);
or U845 (N_845,In_100,N_341);
or U846 (N_846,N_73,N_531);
xor U847 (N_847,In_1032,In_808);
nor U848 (N_848,N_632,N_698);
xor U849 (N_849,N_109,In_48);
and U850 (N_850,N_524,In_1362);
and U851 (N_851,In_1456,In_909);
nand U852 (N_852,N_451,In_1477);
nand U853 (N_853,In_550,N_402);
nand U854 (N_854,N_256,N_532);
and U855 (N_855,In_326,N_463);
nor U856 (N_856,In_87,In_454);
nor U857 (N_857,N_136,In_424);
nand U858 (N_858,N_685,N_359);
nor U859 (N_859,N_96,N_465);
or U860 (N_860,In_400,In_667);
nor U861 (N_861,In_664,N_348);
xnor U862 (N_862,N_308,N_705);
and U863 (N_863,N_509,N_472);
nand U864 (N_864,In_1023,In_489);
nand U865 (N_865,In_1394,In_1418);
nor U866 (N_866,In_639,N_150);
nor U867 (N_867,N_523,N_544);
or U868 (N_868,N_679,In_84);
or U869 (N_869,N_746,In_274);
xnor U870 (N_870,In_425,N_414);
and U871 (N_871,In_913,In_714);
xnor U872 (N_872,N_431,N_556);
xnor U873 (N_873,In_954,N_545);
xor U874 (N_874,N_488,N_522);
xor U875 (N_875,In_813,N_634);
nor U876 (N_876,N_691,N_657);
or U877 (N_877,In_227,In_1348);
and U878 (N_878,N_101,N_707);
or U879 (N_879,N_462,In_1482);
or U880 (N_880,N_723,N_484);
nor U881 (N_881,N_474,N_192);
and U882 (N_882,In_1095,N_623);
nand U883 (N_883,In_1294,N_607);
xor U884 (N_884,In_502,In_251);
nand U885 (N_885,N_742,N_533);
nand U886 (N_886,N_729,N_242);
nor U887 (N_887,N_710,In_495);
xor U888 (N_888,N_572,In_952);
and U889 (N_889,In_1141,In_1093);
nor U890 (N_890,N_198,N_669);
nand U891 (N_891,In_532,N_388);
xor U892 (N_892,In_1309,In_1078);
nor U893 (N_893,In_1085,N_624);
or U894 (N_894,N_586,In_207);
nand U895 (N_895,In_166,N_670);
nor U896 (N_896,In_465,N_14);
and U897 (N_897,N_561,In_925);
nand U898 (N_898,In_413,N_18);
nor U899 (N_899,In_539,N_158);
nand U900 (N_900,N_48,In_131);
nor U901 (N_901,In_699,In_923);
and U902 (N_902,In_562,In_920);
nand U903 (N_903,N_876,N_356);
nand U904 (N_904,In_612,N_491);
nor U905 (N_905,N_804,N_601);
nor U906 (N_906,N_49,N_187);
nand U907 (N_907,N_704,N_817);
nand U908 (N_908,N_765,N_619);
and U909 (N_909,N_674,N_763);
or U910 (N_910,N_391,N_837);
and U911 (N_911,In_992,N_715);
and U912 (N_912,N_689,N_881);
xnor U913 (N_913,In_1240,In_94);
nor U914 (N_914,In_1025,N_468);
xnor U915 (N_915,N_629,N_173);
nand U916 (N_916,N_816,N_595);
nand U917 (N_917,N_776,N_214);
nor U918 (N_918,In_1129,N_700);
nand U919 (N_919,In_907,N_307);
and U920 (N_920,In_691,N_510);
nand U921 (N_921,N_761,N_501);
and U922 (N_922,In_54,N_802);
or U923 (N_923,N_498,In_574);
nor U924 (N_924,In_1029,N_563);
xor U925 (N_925,In_219,N_148);
nand U926 (N_926,In_33,N_511);
nor U927 (N_927,In_1293,N_281);
and U928 (N_928,In_175,In_1059);
or U929 (N_929,N_284,N_854);
nand U930 (N_930,In_1136,N_867);
nor U931 (N_931,N_692,N_489);
or U932 (N_932,N_751,N_647);
or U933 (N_933,In_355,In_375);
and U934 (N_934,N_655,N_779);
xor U935 (N_935,In_1152,N_604);
and U936 (N_936,N_784,N_536);
xnor U937 (N_937,N_400,N_519);
or U938 (N_938,N_609,N_537);
xnor U939 (N_939,N_853,In_1171);
nand U940 (N_940,N_847,N_331);
xor U941 (N_941,N_26,In_1389);
and U942 (N_942,In_777,In_1471);
and U943 (N_943,In_347,In_275);
xor U944 (N_944,N_120,In_357);
and U945 (N_945,N_875,In_1337);
nor U946 (N_946,In_230,N_824);
nor U947 (N_947,In_793,In_1227);
xor U948 (N_948,In_1062,N_738);
xor U949 (N_949,N_598,N_800);
and U950 (N_950,N_646,N_877);
or U951 (N_951,N_371,N_883);
xnor U952 (N_952,In_636,N_895);
nand U953 (N_953,In_1194,N_628);
xor U954 (N_954,In_1345,N_380);
or U955 (N_955,N_795,N_616);
or U956 (N_956,In_1333,N_731);
or U957 (N_957,In_191,In_604);
nand U958 (N_958,In_223,In_405);
xnor U959 (N_959,N_208,N_584);
and U960 (N_960,N_61,N_805);
nand U961 (N_961,N_852,N_411);
or U962 (N_962,In_596,N_270);
nand U963 (N_963,N_834,N_719);
xnor U964 (N_964,In_996,N_683);
nand U965 (N_965,N_848,N_833);
xnor U966 (N_966,N_182,N_454);
nor U967 (N_967,N_397,N_894);
xor U968 (N_968,In_1192,N_809);
xor U969 (N_969,N_254,N_720);
nand U970 (N_970,N_568,N_799);
and U971 (N_971,In_1271,In_1041);
xor U972 (N_972,N_379,N_175);
and U973 (N_973,In_811,N_78);
nor U974 (N_974,In_1051,In_262);
nand U975 (N_975,N_838,In_1376);
and U976 (N_976,N_762,N_830);
nor U977 (N_977,N_617,In_993);
xnor U978 (N_978,N_819,N_718);
or U979 (N_979,In_1319,In_1283);
nand U980 (N_980,N_119,N_174);
nand U981 (N_981,In_315,N_211);
and U982 (N_982,N_862,N_808);
xnor U983 (N_983,In_669,In_51);
and U984 (N_984,N_845,N_716);
or U985 (N_985,N_760,In_1006);
or U986 (N_986,N_567,In_4);
nand U987 (N_987,N_366,N_825);
nor U988 (N_988,N_889,In_431);
xor U989 (N_989,N_726,N_870);
nand U990 (N_990,N_768,N_806);
nand U991 (N_991,N_866,N_897);
or U992 (N_992,N_525,In_1115);
xnor U993 (N_993,N_773,In_794);
nand U994 (N_994,In_1265,N_772);
and U995 (N_995,In_1415,N_167);
xor U996 (N_996,N_712,N_336);
xor U997 (N_997,N_878,N_639);
xor U998 (N_998,N_832,N_219);
nand U999 (N_999,N_606,In_226);
nor U1000 (N_1000,N_303,In_330);
nand U1001 (N_1001,In_756,N_552);
nand U1002 (N_1002,N_886,In_15);
or U1003 (N_1003,In_1017,N_529);
nand U1004 (N_1004,N_581,In_344);
xnor U1005 (N_1005,N_766,In_188);
nor U1006 (N_1006,In_637,In_626);
and U1007 (N_1007,In_1462,N_815);
nor U1008 (N_1008,In_204,N_298);
nand U1009 (N_1009,In_690,N_615);
nor U1010 (N_1010,In_933,In_160);
or U1011 (N_1011,N_818,N_666);
nor U1012 (N_1012,In_1277,N_633);
nor U1013 (N_1013,N_841,N_717);
nand U1014 (N_1014,N_869,N_223);
or U1015 (N_1015,In_716,N_823);
and U1016 (N_1016,N_652,N_596);
xnor U1017 (N_1017,In_825,In_666);
and U1018 (N_1018,In_260,In_584);
or U1019 (N_1019,In_74,N_504);
or U1020 (N_1020,N_813,In_898);
nor U1021 (N_1021,In_1330,N_667);
and U1022 (N_1022,In_867,In_1272);
nand U1023 (N_1023,N_415,In_828);
xor U1024 (N_1024,In_446,N_829);
nand U1025 (N_1025,N_677,N_337);
nand U1026 (N_1026,N_794,In_150);
or U1027 (N_1027,N_82,N_774);
and U1028 (N_1028,N_787,N_855);
or U1029 (N_1029,N_812,N_828);
or U1030 (N_1030,N_790,In_369);
xor U1031 (N_1031,N_722,In_78);
or U1032 (N_1032,In_139,N_301);
nand U1033 (N_1033,In_1204,N_899);
nor U1034 (N_1034,N_740,N_874);
nor U1035 (N_1035,N_668,In_1427);
and U1036 (N_1036,In_1282,N_822);
nand U1037 (N_1037,N_200,N_891);
or U1038 (N_1038,In_392,In_213);
nor U1039 (N_1039,N_475,In_1459);
nand U1040 (N_1040,N_827,N_218);
nand U1041 (N_1041,N_430,In_1117);
xnor U1042 (N_1042,N_492,In_955);
nor U1043 (N_1043,N_399,N_673);
xnor U1044 (N_1044,In_606,N_582);
or U1045 (N_1045,N_553,N_612);
nor U1046 (N_1046,In_931,N_512);
nor U1047 (N_1047,N_361,In_1164);
and U1048 (N_1048,N_675,In_435);
nand U1049 (N_1049,N_775,N_410);
xor U1050 (N_1050,N_963,N_1030);
nand U1051 (N_1051,N_937,N_503);
nand U1052 (N_1052,In_981,N_968);
xor U1053 (N_1053,N_367,In_421);
nor U1054 (N_1054,In_389,N_789);
or U1055 (N_1055,N_656,N_896);
and U1056 (N_1056,N_706,N_941);
or U1057 (N_1057,N_872,N_171);
or U1058 (N_1058,N_916,N_453);
xnor U1059 (N_1059,In_243,N_951);
nor U1060 (N_1060,N_1014,N_915);
or U1061 (N_1061,N_864,N_513);
or U1062 (N_1062,In_607,N_334);
nand U1063 (N_1063,N_982,In_1039);
and U1064 (N_1064,N_555,N_178);
xor U1065 (N_1065,N_351,N_1042);
or U1066 (N_1066,N_534,N_237);
xor U1067 (N_1067,In_736,N_826);
or U1068 (N_1068,N_1007,N_1025);
xor U1069 (N_1069,In_437,N_796);
nor U1070 (N_1070,In_628,N_922);
xnor U1071 (N_1071,N_734,N_969);
xnor U1072 (N_1072,N_898,N_395);
or U1073 (N_1073,N_927,In_348);
nand U1074 (N_1074,N_964,N_786);
nor U1075 (N_1075,N_924,N_859);
or U1076 (N_1076,N_945,In_1046);
nor U1077 (N_1077,N_831,N_890);
nand U1078 (N_1078,In_1050,In_3);
nand U1079 (N_1079,N_1031,In_720);
nand U1080 (N_1080,N_392,N_810);
nor U1081 (N_1081,N_990,In_1203);
nor U1082 (N_1082,N_970,N_975);
xor U1083 (N_1083,In_743,N_540);
xor U1084 (N_1084,In_122,N_680);
and U1085 (N_1085,N_991,N_1029);
xnor U1086 (N_1086,N_835,N_1002);
xnor U1087 (N_1087,In_578,N_428);
nand U1088 (N_1088,In_463,In_625);
or U1089 (N_1089,In_1170,N_1043);
nor U1090 (N_1090,In_114,In_200);
and U1091 (N_1091,N_613,N_747);
or U1092 (N_1092,N_739,N_69);
nand U1093 (N_1093,In_1208,In_0);
and U1094 (N_1094,In_967,In_291);
or U1095 (N_1095,N_714,N_353);
or U1096 (N_1096,N_386,N_844);
xor U1097 (N_1097,N_1023,N_955);
and U1098 (N_1098,N_1012,N_1027);
nand U1099 (N_1099,N_1018,In_127);
xnor U1100 (N_1100,N_342,In_534);
and U1101 (N_1101,N_931,In_320);
nand U1102 (N_1102,N_202,N_676);
nand U1103 (N_1103,N_494,N_928);
nand U1104 (N_1104,N_778,N_641);
or U1105 (N_1105,N_1015,N_695);
nand U1106 (N_1106,In_665,N_921);
and U1107 (N_1107,N_954,N_1040);
or U1108 (N_1108,N_981,N_860);
nor U1109 (N_1109,N_630,In_342);
nand U1110 (N_1110,N_373,N_195);
and U1111 (N_1111,N_914,N_839);
xnor U1112 (N_1112,N_933,In_582);
nor U1113 (N_1113,N_995,N_902);
xnor U1114 (N_1114,In_822,N_901);
nand U1115 (N_1115,N_51,N_736);
and U1116 (N_1116,N_557,N_583);
xor U1117 (N_1117,N_780,N_868);
xor U1118 (N_1118,N_767,N_1028);
nor U1119 (N_1119,N_575,N_811);
nor U1120 (N_1120,N_28,N_661);
nand U1121 (N_1121,N_243,N_910);
or U1122 (N_1122,N_858,N_653);
or U1123 (N_1123,N_727,N_551);
and U1124 (N_1124,N_1017,In_1468);
and U1125 (N_1125,N_1009,N_976);
or U1126 (N_1126,N_961,N_913);
nand U1127 (N_1127,N_984,N_985);
nor U1128 (N_1128,N_626,N_983);
nand U1129 (N_1129,N_888,N_950);
xnor U1130 (N_1130,In_433,N_842);
xor U1131 (N_1131,N_797,In_554);
nand U1132 (N_1132,In_77,N_998);
nor U1133 (N_1133,N_987,N_807);
nand U1134 (N_1134,In_216,N_856);
or U1135 (N_1135,In_189,In_305);
or U1136 (N_1136,In_711,In_1096);
and U1137 (N_1137,N_907,N_903);
nor U1138 (N_1138,In_1063,N_354);
nor U1139 (N_1139,N_527,N_404);
nand U1140 (N_1140,In_708,N_665);
nand U1141 (N_1141,N_840,N_571);
nand U1142 (N_1142,In_1198,N_947);
xnor U1143 (N_1143,N_926,N_994);
and U1144 (N_1144,In_609,N_375);
and U1145 (N_1145,N_863,In_911);
and U1146 (N_1146,N_923,N_803);
nor U1147 (N_1147,N_884,N_759);
and U1148 (N_1148,N_47,N_959);
and U1149 (N_1149,N_640,In_840);
nor U1150 (N_1150,In_116,N_67);
nand U1151 (N_1151,N_183,N_997);
xnor U1152 (N_1152,N_908,N_752);
and U1153 (N_1153,In_111,N_791);
nand U1154 (N_1154,In_764,N_836);
xor U1155 (N_1155,In_723,In_387);
or U1156 (N_1156,N_365,N_50);
and U1157 (N_1157,N_435,N_1008);
and U1158 (N_1158,N_857,N_1001);
nand U1159 (N_1159,In_593,N_793);
and U1160 (N_1160,N_936,In_412);
xor U1161 (N_1161,N_934,N_999);
nor U1162 (N_1162,N_880,N_393);
or U1163 (N_1163,N_694,N_756);
nand U1164 (N_1164,In_673,N_892);
nor U1165 (N_1165,N_282,N_939);
nor U1166 (N_1166,N_1044,N_977);
or U1167 (N_1167,N_664,N_530);
nor U1168 (N_1168,N_360,N_917);
nand U1169 (N_1169,N_769,N_755);
nand U1170 (N_1170,N_785,N_1004);
nand U1171 (N_1171,N_434,In_535);
nand U1172 (N_1172,N_851,N_801);
xor U1173 (N_1173,In_790,In_409);
and U1174 (N_1174,In_1341,In_153);
nand U1175 (N_1175,N_693,N_906);
xnor U1176 (N_1176,N_962,In_59);
or U1177 (N_1177,N_701,N_965);
nor U1178 (N_1178,N_958,N_938);
or U1179 (N_1179,N_948,N_702);
xor U1180 (N_1180,In_1140,N_733);
xnor U1181 (N_1181,N_549,N_893);
or U1182 (N_1182,N_873,N_1046);
or U1183 (N_1183,N_564,N_618);
or U1184 (N_1184,N_574,N_871);
nor U1185 (N_1185,N_861,N_912);
or U1186 (N_1186,In_289,In_752);
and U1187 (N_1187,N_925,N_949);
xor U1188 (N_1188,N_992,N_935);
xnor U1189 (N_1189,N_764,N_1021);
xnor U1190 (N_1190,N_957,N_1034);
and U1191 (N_1191,N_770,N_1022);
or U1192 (N_1192,In_1303,N_986);
nor U1193 (N_1193,N_1020,N_77);
xnor U1194 (N_1194,N_885,N_658);
or U1195 (N_1195,In_496,N_909);
nor U1196 (N_1196,N_974,N_245);
nor U1197 (N_1197,N_1048,N_516);
nand U1198 (N_1198,N_753,In_249);
nor U1199 (N_1199,N_973,In_136);
xor U1200 (N_1200,N_1105,N_1193);
xnor U1201 (N_1201,N_1153,N_1155);
or U1202 (N_1202,N_754,N_1111);
nand U1203 (N_1203,In_1026,N_1185);
xor U1204 (N_1204,N_750,N_1135);
nor U1205 (N_1205,N_1055,N_1162);
and U1206 (N_1206,N_918,N_798);
xnor U1207 (N_1207,N_1133,N_1108);
nor U1208 (N_1208,N_905,N_1016);
xnor U1209 (N_1209,N_1033,N_1013);
or U1210 (N_1210,N_1176,N_1130);
nor U1211 (N_1211,N_1122,N_1107);
xnor U1212 (N_1212,N_1114,N_1102);
nor U1213 (N_1213,N_1106,In_1199);
nor U1214 (N_1214,N_1082,N_1060);
and U1215 (N_1215,N_1041,N_1050);
nor U1216 (N_1216,N_1113,N_932);
nor U1217 (N_1217,N_1120,In_452);
xnor U1218 (N_1218,N_744,N_1104);
nor U1219 (N_1219,N_1138,N_1199);
nand U1220 (N_1220,N_788,N_1061);
nor U1221 (N_1221,In_152,N_1024);
or U1222 (N_1222,N_1149,N_1112);
nor U1223 (N_1223,N_887,In_1311);
nand U1224 (N_1224,N_1184,N_1195);
and U1225 (N_1225,N_1098,N_771);
nor U1226 (N_1226,N_953,N_919);
xnor U1227 (N_1227,N_1100,N_68);
xor U1228 (N_1228,N_1072,N_900);
xor U1229 (N_1229,N_820,N_644);
or U1230 (N_1230,N_1157,N_849);
or U1231 (N_1231,N_1189,In_1179);
or U1232 (N_1232,N_1158,N_1163);
or U1233 (N_1233,N_1070,N_608);
nand U1234 (N_1234,In_884,N_1110);
nor U1235 (N_1235,N_317,N_814);
xor U1236 (N_1236,N_960,N_456);
and U1237 (N_1237,N_988,N_850);
or U1238 (N_1238,N_944,N_777);
nor U1239 (N_1239,N_846,N_1091);
nand U1240 (N_1240,N_1064,N_547);
or U1241 (N_1241,N_1181,N_956);
nand U1242 (N_1242,In_366,N_1121);
nand U1243 (N_1243,In_1065,N_329);
or U1244 (N_1244,N_942,N_1069);
xor U1245 (N_1245,N_728,N_1154);
nand U1246 (N_1246,N_1140,N_882);
nor U1247 (N_1247,N_1179,N_972);
or U1248 (N_1248,In_497,N_1159);
nand U1249 (N_1249,N_1103,In_372);
or U1250 (N_1250,N_1035,N_1094);
nor U1251 (N_1251,N_1132,N_1167);
or U1252 (N_1252,N_1180,N_1150);
nand U1253 (N_1253,N_1006,In_872);
and U1254 (N_1254,N_1057,N_1000);
xor U1255 (N_1255,N_1003,N_425);
xor U1256 (N_1256,N_1188,N_1169);
nand U1257 (N_1257,N_1178,N_27);
nor U1258 (N_1258,In_1196,In_1328);
nand U1259 (N_1259,N_1062,N_1151);
and U1260 (N_1260,N_1143,N_743);
xnor U1261 (N_1261,N_940,In_834);
or U1262 (N_1262,N_570,In_876);
nand U1263 (N_1263,N_1177,N_1129);
or U1264 (N_1264,N_1010,N_1192);
nor U1265 (N_1265,N_1174,N_1124);
and U1266 (N_1266,N_971,N_1058);
xor U1267 (N_1267,N_978,N_1109);
nand U1268 (N_1268,N_1170,N_1141);
or U1269 (N_1269,N_1148,N_1099);
nor U1270 (N_1270,N_660,N_1085);
xor U1271 (N_1271,N_979,N_1054);
nor U1272 (N_1272,N_865,In_1082);
nor U1273 (N_1273,N_1011,N_1197);
nor U1274 (N_1274,N_426,N_1084);
xnor U1275 (N_1275,N_1191,N_1160);
or U1276 (N_1276,N_758,N_1045);
nor U1277 (N_1277,N_996,N_1093);
or U1278 (N_1278,In_9,N_1047);
or U1279 (N_1279,N_1139,N_1053);
nand U1280 (N_1280,N_1036,N_1076);
or U1281 (N_1281,N_1063,N_930);
or U1282 (N_1282,N_1096,N_748);
xor U1283 (N_1283,N_821,In_600);
nor U1284 (N_1284,N_690,N_1051);
nor U1285 (N_1285,N_1026,In_341);
nor U1286 (N_1286,N_1134,N_920);
or U1287 (N_1287,N_1081,N_579);
nand U1288 (N_1288,N_140,N_904);
xor U1289 (N_1289,N_1087,N_1083);
or U1290 (N_1290,N_911,In_698);
nor U1291 (N_1291,N_452,N_1131);
and U1292 (N_1292,N_783,N_989);
and U1293 (N_1293,N_1115,N_1075);
xor U1294 (N_1294,N_1090,N_1144);
or U1295 (N_1295,N_1183,In_1036);
xnor U1296 (N_1296,N_1066,In_950);
nor U1297 (N_1297,N_593,N_196);
nand U1298 (N_1298,N_1056,N_374);
xor U1299 (N_1299,N_293,N_1146);
xor U1300 (N_1300,N_1156,N_1123);
nor U1301 (N_1301,N_1068,N_929);
nand U1302 (N_1302,N_966,N_620);
nor U1303 (N_1303,N_1171,N_1071);
xnor U1304 (N_1304,N_1079,In_308);
nand U1305 (N_1305,N_943,N_1152);
and U1306 (N_1306,N_1136,In_1447);
nand U1307 (N_1307,N_1166,N_1065);
nor U1308 (N_1308,N_1101,N_1059);
and U1309 (N_1309,N_1182,N_663);
or U1310 (N_1310,N_1074,N_1164);
xor U1311 (N_1311,N_1190,N_1080);
nor U1312 (N_1312,N_1032,In_742);
and U1313 (N_1313,N_1117,N_1145);
nor U1314 (N_1314,In_1453,N_696);
or U1315 (N_1315,N_1165,N_735);
xnor U1316 (N_1316,N_1198,N_1147);
nor U1317 (N_1317,N_1142,N_602);
and U1318 (N_1318,N_1089,N_879);
or U1319 (N_1319,N_713,In_529);
and U1320 (N_1320,N_1175,In_1344);
or U1321 (N_1321,N_1092,N_1118);
xor U1322 (N_1322,N_967,N_757);
and U1323 (N_1323,N_1186,N_1161);
and U1324 (N_1324,N_1005,In_929);
and U1325 (N_1325,In_461,N_843);
or U1326 (N_1326,N_792,N_1116);
and U1327 (N_1327,In_650,N_1086);
and U1328 (N_1328,N_1194,In_1067);
nand U1329 (N_1329,N_1077,N_1095);
nor U1330 (N_1330,N_781,N_306);
nor U1331 (N_1331,N_1019,N_1038);
xnor U1332 (N_1332,N_1088,N_1196);
or U1333 (N_1333,N_1067,N_993);
and U1334 (N_1334,N_320,N_1127);
and U1335 (N_1335,N_438,N_605);
nand U1336 (N_1336,In_543,N_1049);
or U1337 (N_1337,N_1119,N_1168);
or U1338 (N_1338,N_1173,N_1137);
and U1339 (N_1339,N_782,N_1097);
nor U1340 (N_1340,N_1172,N_1187);
and U1341 (N_1341,N_1073,In_442);
and U1342 (N_1342,N_980,N_708);
nor U1343 (N_1343,N_323,N_952);
and U1344 (N_1344,N_1125,N_1126);
and U1345 (N_1345,In_942,N_643);
or U1346 (N_1346,N_1078,N_496);
nand U1347 (N_1347,N_1128,N_645);
or U1348 (N_1348,N_1039,N_1052);
nor U1349 (N_1349,N_946,N_1037);
xor U1350 (N_1350,N_1212,N_1216);
or U1351 (N_1351,N_1309,N_1349);
xor U1352 (N_1352,N_1269,N_1335);
and U1353 (N_1353,N_1291,N_1287);
or U1354 (N_1354,N_1319,N_1222);
or U1355 (N_1355,N_1228,N_1272);
nor U1356 (N_1356,N_1311,N_1277);
or U1357 (N_1357,N_1203,N_1262);
nor U1358 (N_1358,N_1226,N_1221);
or U1359 (N_1359,N_1202,N_1204);
and U1360 (N_1360,N_1298,N_1331);
nor U1361 (N_1361,N_1288,N_1206);
or U1362 (N_1362,N_1292,N_1253);
or U1363 (N_1363,N_1310,N_1315);
nand U1364 (N_1364,N_1205,N_1241);
or U1365 (N_1365,N_1313,N_1305);
xnor U1366 (N_1366,N_1254,N_1209);
nand U1367 (N_1367,N_1250,N_1289);
nor U1368 (N_1368,N_1236,N_1321);
and U1369 (N_1369,N_1265,N_1294);
or U1370 (N_1370,N_1258,N_1296);
and U1371 (N_1371,N_1246,N_1245);
xor U1372 (N_1372,N_1295,N_1260);
or U1373 (N_1373,N_1306,N_1279);
xnor U1374 (N_1374,N_1225,N_1213);
nand U1375 (N_1375,N_1318,N_1333);
xor U1376 (N_1376,N_1268,N_1345);
nand U1377 (N_1377,N_1242,N_1303);
nor U1378 (N_1378,N_1334,N_1290);
or U1379 (N_1379,N_1261,N_1264);
or U1380 (N_1380,N_1229,N_1324);
nor U1381 (N_1381,N_1314,N_1344);
xnor U1382 (N_1382,N_1256,N_1238);
xor U1383 (N_1383,N_1200,N_1281);
and U1384 (N_1384,N_1259,N_1342);
nor U1385 (N_1385,N_1224,N_1234);
nor U1386 (N_1386,N_1208,N_1348);
xor U1387 (N_1387,N_1337,N_1227);
and U1388 (N_1388,N_1270,N_1274);
xnor U1389 (N_1389,N_1230,N_1302);
and U1390 (N_1390,N_1341,N_1329);
or U1391 (N_1391,N_1220,N_1263);
nand U1392 (N_1392,N_1215,N_1330);
nand U1393 (N_1393,N_1340,N_1284);
nor U1394 (N_1394,N_1276,N_1223);
and U1395 (N_1395,N_1299,N_1332);
and U1396 (N_1396,N_1239,N_1231);
and U1397 (N_1397,N_1286,N_1325);
nor U1398 (N_1398,N_1338,N_1308);
or U1399 (N_1399,N_1322,N_1271);
nand U1400 (N_1400,N_1326,N_1243);
nand U1401 (N_1401,N_1343,N_1211);
xor U1402 (N_1402,N_1217,N_1249);
or U1403 (N_1403,N_1307,N_1237);
xor U1404 (N_1404,N_1339,N_1248);
xor U1405 (N_1405,N_1275,N_1328);
and U1406 (N_1406,N_1317,N_1293);
or U1407 (N_1407,N_1244,N_1219);
or U1408 (N_1408,N_1301,N_1235);
or U1409 (N_1409,N_1266,N_1267);
and U1410 (N_1410,N_1297,N_1280);
or U1411 (N_1411,N_1201,N_1255);
nand U1412 (N_1412,N_1232,N_1233);
nand U1413 (N_1413,N_1207,N_1285);
nor U1414 (N_1414,N_1300,N_1312);
nand U1415 (N_1415,N_1327,N_1282);
nor U1416 (N_1416,N_1251,N_1210);
or U1417 (N_1417,N_1214,N_1320);
nor U1418 (N_1418,N_1304,N_1347);
nor U1419 (N_1419,N_1240,N_1323);
nand U1420 (N_1420,N_1252,N_1316);
xor U1421 (N_1421,N_1283,N_1346);
xnor U1422 (N_1422,N_1257,N_1247);
xor U1423 (N_1423,N_1336,N_1278);
and U1424 (N_1424,N_1218,N_1273);
nor U1425 (N_1425,N_1291,N_1301);
or U1426 (N_1426,N_1258,N_1215);
nand U1427 (N_1427,N_1263,N_1325);
and U1428 (N_1428,N_1241,N_1246);
xor U1429 (N_1429,N_1277,N_1281);
xnor U1430 (N_1430,N_1210,N_1236);
nor U1431 (N_1431,N_1330,N_1348);
and U1432 (N_1432,N_1238,N_1208);
xor U1433 (N_1433,N_1313,N_1348);
nand U1434 (N_1434,N_1322,N_1325);
nand U1435 (N_1435,N_1325,N_1248);
or U1436 (N_1436,N_1307,N_1330);
xnor U1437 (N_1437,N_1310,N_1294);
xnor U1438 (N_1438,N_1276,N_1278);
and U1439 (N_1439,N_1295,N_1277);
xnor U1440 (N_1440,N_1250,N_1274);
xor U1441 (N_1441,N_1204,N_1326);
or U1442 (N_1442,N_1274,N_1331);
or U1443 (N_1443,N_1345,N_1321);
xor U1444 (N_1444,N_1239,N_1202);
nand U1445 (N_1445,N_1205,N_1319);
nor U1446 (N_1446,N_1267,N_1290);
xnor U1447 (N_1447,N_1288,N_1224);
nor U1448 (N_1448,N_1273,N_1249);
or U1449 (N_1449,N_1298,N_1282);
nand U1450 (N_1450,N_1222,N_1290);
or U1451 (N_1451,N_1259,N_1294);
xnor U1452 (N_1452,N_1225,N_1224);
nand U1453 (N_1453,N_1266,N_1342);
xnor U1454 (N_1454,N_1340,N_1288);
nand U1455 (N_1455,N_1283,N_1210);
xor U1456 (N_1456,N_1280,N_1287);
or U1457 (N_1457,N_1345,N_1203);
or U1458 (N_1458,N_1308,N_1312);
and U1459 (N_1459,N_1295,N_1283);
or U1460 (N_1460,N_1303,N_1232);
and U1461 (N_1461,N_1264,N_1200);
or U1462 (N_1462,N_1227,N_1258);
nand U1463 (N_1463,N_1279,N_1218);
xnor U1464 (N_1464,N_1264,N_1328);
nor U1465 (N_1465,N_1218,N_1342);
or U1466 (N_1466,N_1289,N_1279);
or U1467 (N_1467,N_1274,N_1313);
or U1468 (N_1468,N_1317,N_1224);
and U1469 (N_1469,N_1276,N_1236);
and U1470 (N_1470,N_1292,N_1250);
or U1471 (N_1471,N_1257,N_1320);
nand U1472 (N_1472,N_1332,N_1315);
and U1473 (N_1473,N_1249,N_1335);
or U1474 (N_1474,N_1241,N_1349);
xnor U1475 (N_1475,N_1334,N_1306);
or U1476 (N_1476,N_1200,N_1290);
or U1477 (N_1477,N_1338,N_1270);
and U1478 (N_1478,N_1209,N_1252);
nand U1479 (N_1479,N_1318,N_1252);
nor U1480 (N_1480,N_1203,N_1286);
xor U1481 (N_1481,N_1347,N_1339);
or U1482 (N_1482,N_1334,N_1265);
xor U1483 (N_1483,N_1279,N_1307);
nor U1484 (N_1484,N_1345,N_1219);
nand U1485 (N_1485,N_1249,N_1207);
or U1486 (N_1486,N_1271,N_1291);
xor U1487 (N_1487,N_1209,N_1346);
and U1488 (N_1488,N_1256,N_1344);
nor U1489 (N_1489,N_1217,N_1315);
xnor U1490 (N_1490,N_1290,N_1241);
xnor U1491 (N_1491,N_1244,N_1255);
nand U1492 (N_1492,N_1329,N_1304);
and U1493 (N_1493,N_1210,N_1293);
nor U1494 (N_1494,N_1270,N_1335);
nand U1495 (N_1495,N_1237,N_1309);
and U1496 (N_1496,N_1346,N_1219);
xor U1497 (N_1497,N_1278,N_1295);
and U1498 (N_1498,N_1303,N_1246);
or U1499 (N_1499,N_1314,N_1290);
or U1500 (N_1500,N_1470,N_1471);
nand U1501 (N_1501,N_1436,N_1487);
or U1502 (N_1502,N_1449,N_1386);
nand U1503 (N_1503,N_1454,N_1411);
nor U1504 (N_1504,N_1372,N_1481);
and U1505 (N_1505,N_1421,N_1445);
and U1506 (N_1506,N_1479,N_1416);
and U1507 (N_1507,N_1488,N_1477);
or U1508 (N_1508,N_1413,N_1398);
or U1509 (N_1509,N_1495,N_1485);
xnor U1510 (N_1510,N_1425,N_1426);
xor U1511 (N_1511,N_1406,N_1392);
and U1512 (N_1512,N_1382,N_1460);
and U1513 (N_1513,N_1461,N_1443);
or U1514 (N_1514,N_1351,N_1389);
and U1515 (N_1515,N_1394,N_1453);
nor U1516 (N_1516,N_1475,N_1467);
and U1517 (N_1517,N_1391,N_1415);
nand U1518 (N_1518,N_1383,N_1486);
nand U1519 (N_1519,N_1385,N_1466);
or U1520 (N_1520,N_1465,N_1494);
nand U1521 (N_1521,N_1366,N_1472);
nor U1522 (N_1522,N_1423,N_1356);
xnor U1523 (N_1523,N_1464,N_1367);
nand U1524 (N_1524,N_1387,N_1354);
xnor U1525 (N_1525,N_1408,N_1399);
nand U1526 (N_1526,N_1499,N_1404);
nand U1527 (N_1527,N_1388,N_1358);
or U1528 (N_1528,N_1396,N_1381);
or U1529 (N_1529,N_1492,N_1395);
or U1530 (N_1530,N_1473,N_1375);
or U1531 (N_1531,N_1365,N_1498);
or U1532 (N_1532,N_1462,N_1405);
nor U1533 (N_1533,N_1397,N_1352);
or U1534 (N_1534,N_1419,N_1360);
nand U1535 (N_1535,N_1402,N_1403);
nor U1536 (N_1536,N_1442,N_1418);
xor U1537 (N_1537,N_1378,N_1489);
nor U1538 (N_1538,N_1371,N_1446);
nand U1539 (N_1539,N_1409,N_1407);
or U1540 (N_1540,N_1448,N_1379);
or U1541 (N_1541,N_1417,N_1420);
or U1542 (N_1542,N_1390,N_1361);
xnor U1543 (N_1543,N_1490,N_1459);
xnor U1544 (N_1544,N_1455,N_1384);
and U1545 (N_1545,N_1496,N_1377);
xnor U1546 (N_1546,N_1373,N_1437);
nand U1547 (N_1547,N_1478,N_1374);
and U1548 (N_1548,N_1363,N_1410);
nor U1549 (N_1549,N_1456,N_1447);
xor U1550 (N_1550,N_1376,N_1439);
xnor U1551 (N_1551,N_1441,N_1457);
nand U1552 (N_1552,N_1440,N_1428);
xor U1553 (N_1553,N_1427,N_1483);
nor U1554 (N_1554,N_1435,N_1433);
xnor U1555 (N_1555,N_1359,N_1431);
nand U1556 (N_1556,N_1400,N_1434);
xor U1557 (N_1557,N_1480,N_1369);
nand U1558 (N_1558,N_1468,N_1355);
nor U1559 (N_1559,N_1497,N_1350);
or U1560 (N_1560,N_1414,N_1364);
nor U1561 (N_1561,N_1438,N_1422);
nor U1562 (N_1562,N_1429,N_1493);
nor U1563 (N_1563,N_1484,N_1491);
nand U1564 (N_1564,N_1469,N_1368);
or U1565 (N_1565,N_1458,N_1476);
and U1566 (N_1566,N_1474,N_1452);
or U1567 (N_1567,N_1424,N_1430);
nand U1568 (N_1568,N_1401,N_1482);
and U1569 (N_1569,N_1380,N_1432);
or U1570 (N_1570,N_1353,N_1450);
or U1571 (N_1571,N_1357,N_1463);
and U1572 (N_1572,N_1362,N_1444);
xor U1573 (N_1573,N_1451,N_1370);
nor U1574 (N_1574,N_1393,N_1412);
nand U1575 (N_1575,N_1394,N_1351);
and U1576 (N_1576,N_1375,N_1486);
or U1577 (N_1577,N_1475,N_1394);
or U1578 (N_1578,N_1371,N_1411);
nand U1579 (N_1579,N_1384,N_1423);
nand U1580 (N_1580,N_1440,N_1393);
or U1581 (N_1581,N_1398,N_1480);
nor U1582 (N_1582,N_1409,N_1362);
nor U1583 (N_1583,N_1392,N_1490);
or U1584 (N_1584,N_1389,N_1376);
nor U1585 (N_1585,N_1388,N_1481);
nor U1586 (N_1586,N_1472,N_1394);
or U1587 (N_1587,N_1474,N_1352);
nor U1588 (N_1588,N_1415,N_1382);
or U1589 (N_1589,N_1353,N_1409);
nand U1590 (N_1590,N_1408,N_1356);
nand U1591 (N_1591,N_1468,N_1435);
xnor U1592 (N_1592,N_1439,N_1453);
nand U1593 (N_1593,N_1457,N_1410);
nor U1594 (N_1594,N_1454,N_1398);
nor U1595 (N_1595,N_1453,N_1387);
nor U1596 (N_1596,N_1353,N_1437);
nor U1597 (N_1597,N_1499,N_1496);
or U1598 (N_1598,N_1415,N_1458);
nor U1599 (N_1599,N_1386,N_1472);
and U1600 (N_1600,N_1384,N_1482);
nor U1601 (N_1601,N_1461,N_1384);
or U1602 (N_1602,N_1407,N_1459);
and U1603 (N_1603,N_1367,N_1351);
nor U1604 (N_1604,N_1408,N_1455);
and U1605 (N_1605,N_1402,N_1412);
xnor U1606 (N_1606,N_1498,N_1380);
and U1607 (N_1607,N_1467,N_1394);
and U1608 (N_1608,N_1388,N_1432);
and U1609 (N_1609,N_1433,N_1425);
xnor U1610 (N_1610,N_1484,N_1379);
or U1611 (N_1611,N_1405,N_1400);
nor U1612 (N_1612,N_1351,N_1441);
or U1613 (N_1613,N_1351,N_1459);
and U1614 (N_1614,N_1467,N_1495);
xnor U1615 (N_1615,N_1419,N_1388);
or U1616 (N_1616,N_1460,N_1441);
or U1617 (N_1617,N_1472,N_1446);
nand U1618 (N_1618,N_1388,N_1483);
nor U1619 (N_1619,N_1397,N_1408);
xnor U1620 (N_1620,N_1416,N_1443);
or U1621 (N_1621,N_1426,N_1417);
and U1622 (N_1622,N_1380,N_1453);
and U1623 (N_1623,N_1460,N_1490);
and U1624 (N_1624,N_1357,N_1422);
or U1625 (N_1625,N_1499,N_1498);
nor U1626 (N_1626,N_1406,N_1431);
nand U1627 (N_1627,N_1438,N_1384);
or U1628 (N_1628,N_1425,N_1469);
or U1629 (N_1629,N_1486,N_1403);
nor U1630 (N_1630,N_1403,N_1465);
or U1631 (N_1631,N_1385,N_1493);
and U1632 (N_1632,N_1473,N_1361);
or U1633 (N_1633,N_1388,N_1498);
nand U1634 (N_1634,N_1435,N_1466);
nand U1635 (N_1635,N_1396,N_1395);
nand U1636 (N_1636,N_1443,N_1404);
nor U1637 (N_1637,N_1416,N_1430);
xnor U1638 (N_1638,N_1382,N_1447);
or U1639 (N_1639,N_1443,N_1455);
or U1640 (N_1640,N_1361,N_1472);
xnor U1641 (N_1641,N_1353,N_1456);
and U1642 (N_1642,N_1496,N_1434);
nand U1643 (N_1643,N_1485,N_1482);
or U1644 (N_1644,N_1488,N_1467);
nor U1645 (N_1645,N_1425,N_1419);
nand U1646 (N_1646,N_1449,N_1440);
xnor U1647 (N_1647,N_1416,N_1369);
xor U1648 (N_1648,N_1376,N_1413);
nand U1649 (N_1649,N_1421,N_1382);
nand U1650 (N_1650,N_1583,N_1598);
nor U1651 (N_1651,N_1547,N_1519);
nand U1652 (N_1652,N_1524,N_1614);
or U1653 (N_1653,N_1511,N_1588);
xor U1654 (N_1654,N_1516,N_1626);
and U1655 (N_1655,N_1646,N_1526);
nor U1656 (N_1656,N_1551,N_1538);
nand U1657 (N_1657,N_1591,N_1567);
and U1658 (N_1658,N_1550,N_1522);
and U1659 (N_1659,N_1618,N_1609);
nand U1660 (N_1660,N_1611,N_1571);
nand U1661 (N_1661,N_1521,N_1514);
xnor U1662 (N_1662,N_1507,N_1616);
or U1663 (N_1663,N_1564,N_1549);
nand U1664 (N_1664,N_1527,N_1530);
nand U1665 (N_1665,N_1606,N_1575);
nor U1666 (N_1666,N_1523,N_1561);
or U1667 (N_1667,N_1622,N_1587);
nor U1668 (N_1668,N_1607,N_1625);
and U1669 (N_1669,N_1581,N_1644);
xnor U1670 (N_1670,N_1534,N_1532);
nand U1671 (N_1671,N_1560,N_1544);
and U1672 (N_1672,N_1510,N_1518);
nor U1673 (N_1673,N_1610,N_1505);
xnor U1674 (N_1674,N_1556,N_1506);
xnor U1675 (N_1675,N_1565,N_1555);
nor U1676 (N_1676,N_1502,N_1623);
nor U1677 (N_1677,N_1536,N_1615);
xnor U1678 (N_1678,N_1582,N_1600);
or U1679 (N_1679,N_1554,N_1640);
and U1680 (N_1680,N_1585,N_1537);
nor U1681 (N_1681,N_1603,N_1533);
and U1682 (N_1682,N_1568,N_1621);
xnor U1683 (N_1683,N_1541,N_1608);
xnor U1684 (N_1684,N_1500,N_1590);
nor U1685 (N_1685,N_1508,N_1579);
xnor U1686 (N_1686,N_1636,N_1525);
or U1687 (N_1687,N_1557,N_1548);
nor U1688 (N_1688,N_1515,N_1617);
nor U1689 (N_1689,N_1627,N_1503);
xnor U1690 (N_1690,N_1535,N_1605);
or U1691 (N_1691,N_1577,N_1504);
nor U1692 (N_1692,N_1593,N_1631);
or U1693 (N_1693,N_1592,N_1558);
or U1694 (N_1694,N_1632,N_1566);
nor U1695 (N_1695,N_1562,N_1584);
or U1696 (N_1696,N_1572,N_1641);
or U1697 (N_1697,N_1559,N_1628);
and U1698 (N_1698,N_1634,N_1520);
or U1699 (N_1699,N_1546,N_1647);
and U1700 (N_1700,N_1529,N_1574);
nor U1701 (N_1701,N_1576,N_1619);
and U1702 (N_1702,N_1624,N_1596);
and U1703 (N_1703,N_1630,N_1589);
xor U1704 (N_1704,N_1542,N_1513);
nand U1705 (N_1705,N_1620,N_1509);
nand U1706 (N_1706,N_1642,N_1543);
xor U1707 (N_1707,N_1553,N_1633);
nor U1708 (N_1708,N_1638,N_1612);
nor U1709 (N_1709,N_1539,N_1629);
nand U1710 (N_1710,N_1649,N_1643);
nand U1711 (N_1711,N_1586,N_1639);
or U1712 (N_1712,N_1501,N_1517);
and U1713 (N_1713,N_1552,N_1635);
nand U1714 (N_1714,N_1569,N_1531);
xor U1715 (N_1715,N_1599,N_1648);
and U1716 (N_1716,N_1597,N_1563);
xnor U1717 (N_1717,N_1512,N_1540);
nand U1718 (N_1718,N_1595,N_1594);
xor U1719 (N_1719,N_1580,N_1637);
or U1720 (N_1720,N_1578,N_1604);
or U1721 (N_1721,N_1601,N_1528);
and U1722 (N_1722,N_1602,N_1613);
xnor U1723 (N_1723,N_1645,N_1545);
nand U1724 (N_1724,N_1570,N_1573);
nor U1725 (N_1725,N_1585,N_1584);
nor U1726 (N_1726,N_1507,N_1579);
and U1727 (N_1727,N_1592,N_1594);
nor U1728 (N_1728,N_1552,N_1544);
nor U1729 (N_1729,N_1639,N_1557);
or U1730 (N_1730,N_1575,N_1544);
or U1731 (N_1731,N_1587,N_1581);
and U1732 (N_1732,N_1525,N_1500);
and U1733 (N_1733,N_1614,N_1517);
xnor U1734 (N_1734,N_1576,N_1588);
nor U1735 (N_1735,N_1556,N_1640);
nor U1736 (N_1736,N_1619,N_1533);
nor U1737 (N_1737,N_1628,N_1567);
xnor U1738 (N_1738,N_1620,N_1529);
and U1739 (N_1739,N_1511,N_1625);
and U1740 (N_1740,N_1562,N_1622);
or U1741 (N_1741,N_1570,N_1512);
nor U1742 (N_1742,N_1538,N_1616);
nand U1743 (N_1743,N_1609,N_1619);
or U1744 (N_1744,N_1500,N_1508);
xnor U1745 (N_1745,N_1646,N_1528);
xor U1746 (N_1746,N_1510,N_1569);
nor U1747 (N_1747,N_1522,N_1582);
and U1748 (N_1748,N_1645,N_1624);
nor U1749 (N_1749,N_1610,N_1590);
nand U1750 (N_1750,N_1636,N_1564);
nand U1751 (N_1751,N_1571,N_1524);
or U1752 (N_1752,N_1538,N_1592);
nand U1753 (N_1753,N_1605,N_1520);
and U1754 (N_1754,N_1546,N_1580);
nand U1755 (N_1755,N_1552,N_1547);
and U1756 (N_1756,N_1518,N_1539);
xnor U1757 (N_1757,N_1507,N_1618);
or U1758 (N_1758,N_1558,N_1522);
nand U1759 (N_1759,N_1532,N_1602);
or U1760 (N_1760,N_1546,N_1627);
or U1761 (N_1761,N_1648,N_1610);
nand U1762 (N_1762,N_1596,N_1525);
and U1763 (N_1763,N_1613,N_1536);
nor U1764 (N_1764,N_1547,N_1598);
or U1765 (N_1765,N_1628,N_1516);
nand U1766 (N_1766,N_1649,N_1519);
xnor U1767 (N_1767,N_1626,N_1604);
nor U1768 (N_1768,N_1598,N_1580);
or U1769 (N_1769,N_1615,N_1620);
nor U1770 (N_1770,N_1635,N_1545);
xor U1771 (N_1771,N_1586,N_1597);
or U1772 (N_1772,N_1607,N_1623);
nand U1773 (N_1773,N_1600,N_1605);
or U1774 (N_1774,N_1504,N_1612);
or U1775 (N_1775,N_1547,N_1577);
and U1776 (N_1776,N_1632,N_1571);
nor U1777 (N_1777,N_1569,N_1541);
nor U1778 (N_1778,N_1522,N_1531);
nand U1779 (N_1779,N_1611,N_1591);
nor U1780 (N_1780,N_1624,N_1647);
nor U1781 (N_1781,N_1508,N_1641);
or U1782 (N_1782,N_1523,N_1518);
nor U1783 (N_1783,N_1618,N_1611);
nor U1784 (N_1784,N_1558,N_1510);
or U1785 (N_1785,N_1508,N_1578);
and U1786 (N_1786,N_1609,N_1640);
nor U1787 (N_1787,N_1585,N_1597);
nor U1788 (N_1788,N_1616,N_1646);
nand U1789 (N_1789,N_1501,N_1563);
and U1790 (N_1790,N_1617,N_1525);
nor U1791 (N_1791,N_1511,N_1547);
and U1792 (N_1792,N_1576,N_1608);
nand U1793 (N_1793,N_1637,N_1618);
nand U1794 (N_1794,N_1563,N_1618);
nand U1795 (N_1795,N_1609,N_1603);
xnor U1796 (N_1796,N_1598,N_1593);
nand U1797 (N_1797,N_1602,N_1621);
xnor U1798 (N_1798,N_1520,N_1531);
nor U1799 (N_1799,N_1617,N_1646);
and U1800 (N_1800,N_1709,N_1661);
and U1801 (N_1801,N_1714,N_1719);
and U1802 (N_1802,N_1653,N_1768);
and U1803 (N_1803,N_1671,N_1695);
and U1804 (N_1804,N_1741,N_1710);
xnor U1805 (N_1805,N_1788,N_1729);
and U1806 (N_1806,N_1692,N_1651);
or U1807 (N_1807,N_1789,N_1795);
and U1808 (N_1808,N_1670,N_1703);
and U1809 (N_1809,N_1732,N_1791);
and U1810 (N_1810,N_1799,N_1777);
or U1811 (N_1811,N_1718,N_1739);
and U1812 (N_1812,N_1750,N_1776);
xnor U1813 (N_1813,N_1775,N_1769);
nor U1814 (N_1814,N_1700,N_1765);
nand U1815 (N_1815,N_1756,N_1664);
or U1816 (N_1816,N_1697,N_1683);
and U1817 (N_1817,N_1781,N_1760);
nand U1818 (N_1818,N_1764,N_1684);
nor U1819 (N_1819,N_1736,N_1650);
and U1820 (N_1820,N_1699,N_1669);
and U1821 (N_1821,N_1672,N_1767);
or U1822 (N_1822,N_1704,N_1657);
nor U1823 (N_1823,N_1798,N_1783);
and U1824 (N_1824,N_1792,N_1687);
nor U1825 (N_1825,N_1786,N_1723);
nor U1826 (N_1826,N_1770,N_1762);
xor U1827 (N_1827,N_1678,N_1663);
xor U1828 (N_1828,N_1787,N_1757);
nand U1829 (N_1829,N_1754,N_1713);
or U1830 (N_1830,N_1674,N_1680);
nor U1831 (N_1831,N_1655,N_1705);
nor U1832 (N_1832,N_1726,N_1694);
or U1833 (N_1833,N_1766,N_1746);
and U1834 (N_1834,N_1759,N_1711);
nand U1835 (N_1835,N_1772,N_1779);
and U1836 (N_1836,N_1696,N_1763);
nor U1837 (N_1837,N_1720,N_1717);
and U1838 (N_1838,N_1780,N_1690);
nor U1839 (N_1839,N_1784,N_1676);
nor U1840 (N_1840,N_1706,N_1725);
nand U1841 (N_1841,N_1667,N_1708);
and U1842 (N_1842,N_1686,N_1737);
nor U1843 (N_1843,N_1749,N_1693);
or U1844 (N_1844,N_1773,N_1743);
nand U1845 (N_1845,N_1698,N_1796);
or U1846 (N_1846,N_1659,N_1730);
xnor U1847 (N_1847,N_1747,N_1734);
nor U1848 (N_1848,N_1738,N_1712);
and U1849 (N_1849,N_1652,N_1724);
xor U1850 (N_1850,N_1681,N_1656);
xor U1851 (N_1851,N_1771,N_1660);
xor U1852 (N_1852,N_1735,N_1761);
nand U1853 (N_1853,N_1665,N_1733);
nand U1854 (N_1854,N_1782,N_1673);
nand U1855 (N_1855,N_1797,N_1658);
xnor U1856 (N_1856,N_1745,N_1685);
xor U1857 (N_1857,N_1666,N_1662);
nor U1858 (N_1858,N_1755,N_1731);
and U1859 (N_1859,N_1785,N_1716);
xor U1860 (N_1860,N_1727,N_1778);
and U1861 (N_1861,N_1679,N_1675);
nand U1862 (N_1862,N_1691,N_1689);
and U1863 (N_1863,N_1707,N_1758);
or U1864 (N_1864,N_1774,N_1790);
and U1865 (N_1865,N_1702,N_1654);
and U1866 (N_1866,N_1742,N_1751);
and U1867 (N_1867,N_1748,N_1721);
xnor U1868 (N_1868,N_1701,N_1728);
or U1869 (N_1869,N_1740,N_1793);
nand U1870 (N_1870,N_1677,N_1715);
nand U1871 (N_1871,N_1744,N_1722);
nor U1872 (N_1872,N_1794,N_1668);
and U1873 (N_1873,N_1752,N_1753);
nand U1874 (N_1874,N_1688,N_1682);
and U1875 (N_1875,N_1744,N_1693);
nand U1876 (N_1876,N_1729,N_1779);
or U1877 (N_1877,N_1681,N_1785);
or U1878 (N_1878,N_1714,N_1667);
xnor U1879 (N_1879,N_1678,N_1672);
nor U1880 (N_1880,N_1677,N_1692);
and U1881 (N_1881,N_1747,N_1758);
xnor U1882 (N_1882,N_1776,N_1792);
xor U1883 (N_1883,N_1791,N_1727);
nand U1884 (N_1884,N_1782,N_1702);
xnor U1885 (N_1885,N_1669,N_1666);
nand U1886 (N_1886,N_1724,N_1745);
nor U1887 (N_1887,N_1782,N_1704);
nand U1888 (N_1888,N_1652,N_1788);
or U1889 (N_1889,N_1738,N_1713);
nand U1890 (N_1890,N_1761,N_1791);
nand U1891 (N_1891,N_1769,N_1773);
xor U1892 (N_1892,N_1672,N_1696);
or U1893 (N_1893,N_1748,N_1727);
nand U1894 (N_1894,N_1772,N_1686);
xor U1895 (N_1895,N_1781,N_1723);
and U1896 (N_1896,N_1687,N_1763);
nor U1897 (N_1897,N_1711,N_1689);
nand U1898 (N_1898,N_1670,N_1694);
xor U1899 (N_1899,N_1725,N_1699);
or U1900 (N_1900,N_1654,N_1710);
or U1901 (N_1901,N_1671,N_1741);
xor U1902 (N_1902,N_1740,N_1754);
xor U1903 (N_1903,N_1667,N_1723);
nand U1904 (N_1904,N_1739,N_1743);
nand U1905 (N_1905,N_1726,N_1703);
nor U1906 (N_1906,N_1658,N_1735);
and U1907 (N_1907,N_1782,N_1654);
nand U1908 (N_1908,N_1775,N_1677);
or U1909 (N_1909,N_1656,N_1746);
nand U1910 (N_1910,N_1722,N_1747);
xnor U1911 (N_1911,N_1784,N_1658);
nand U1912 (N_1912,N_1681,N_1799);
or U1913 (N_1913,N_1650,N_1758);
and U1914 (N_1914,N_1740,N_1775);
xor U1915 (N_1915,N_1686,N_1702);
or U1916 (N_1916,N_1795,N_1696);
or U1917 (N_1917,N_1778,N_1673);
nor U1918 (N_1918,N_1713,N_1741);
or U1919 (N_1919,N_1653,N_1733);
nand U1920 (N_1920,N_1795,N_1721);
or U1921 (N_1921,N_1750,N_1718);
xor U1922 (N_1922,N_1743,N_1678);
nand U1923 (N_1923,N_1696,N_1762);
nand U1924 (N_1924,N_1707,N_1775);
and U1925 (N_1925,N_1725,N_1653);
nand U1926 (N_1926,N_1686,N_1656);
nor U1927 (N_1927,N_1743,N_1776);
nor U1928 (N_1928,N_1758,N_1779);
nor U1929 (N_1929,N_1679,N_1698);
and U1930 (N_1930,N_1767,N_1651);
or U1931 (N_1931,N_1719,N_1677);
nand U1932 (N_1932,N_1777,N_1662);
and U1933 (N_1933,N_1707,N_1688);
nor U1934 (N_1934,N_1685,N_1736);
nor U1935 (N_1935,N_1778,N_1722);
and U1936 (N_1936,N_1699,N_1754);
and U1937 (N_1937,N_1697,N_1780);
or U1938 (N_1938,N_1703,N_1678);
nor U1939 (N_1939,N_1721,N_1728);
nand U1940 (N_1940,N_1682,N_1782);
and U1941 (N_1941,N_1729,N_1651);
nor U1942 (N_1942,N_1669,N_1773);
nor U1943 (N_1943,N_1704,N_1774);
or U1944 (N_1944,N_1763,N_1684);
or U1945 (N_1945,N_1663,N_1691);
and U1946 (N_1946,N_1712,N_1679);
nand U1947 (N_1947,N_1662,N_1698);
and U1948 (N_1948,N_1743,N_1687);
or U1949 (N_1949,N_1701,N_1772);
xor U1950 (N_1950,N_1845,N_1883);
nand U1951 (N_1951,N_1829,N_1899);
or U1952 (N_1952,N_1801,N_1949);
nand U1953 (N_1953,N_1930,N_1810);
xor U1954 (N_1954,N_1900,N_1922);
nand U1955 (N_1955,N_1889,N_1885);
and U1956 (N_1956,N_1827,N_1907);
and U1957 (N_1957,N_1923,N_1929);
nor U1958 (N_1958,N_1882,N_1800);
nand U1959 (N_1959,N_1818,N_1913);
nand U1960 (N_1960,N_1861,N_1833);
or U1961 (N_1961,N_1870,N_1921);
nand U1962 (N_1962,N_1931,N_1817);
xor U1963 (N_1963,N_1840,N_1808);
and U1964 (N_1964,N_1920,N_1828);
or U1965 (N_1965,N_1902,N_1830);
and U1966 (N_1966,N_1914,N_1877);
and U1967 (N_1967,N_1822,N_1925);
xor U1968 (N_1968,N_1935,N_1847);
and U1969 (N_1969,N_1897,N_1891);
or U1970 (N_1970,N_1881,N_1919);
nor U1971 (N_1971,N_1887,N_1896);
and U1972 (N_1972,N_1886,N_1823);
xor U1973 (N_1973,N_1836,N_1943);
nand U1974 (N_1974,N_1814,N_1936);
nor U1975 (N_1975,N_1873,N_1806);
or U1976 (N_1976,N_1893,N_1928);
nand U1977 (N_1977,N_1838,N_1851);
nand U1978 (N_1978,N_1831,N_1917);
or U1979 (N_1979,N_1804,N_1862);
and U1980 (N_1980,N_1908,N_1938);
and U1981 (N_1981,N_1942,N_1821);
or U1982 (N_1982,N_1909,N_1884);
nand U1983 (N_1983,N_1802,N_1812);
nor U1984 (N_1984,N_1820,N_1876);
and U1985 (N_1985,N_1859,N_1946);
or U1986 (N_1986,N_1941,N_1807);
nand U1987 (N_1987,N_1871,N_1932);
nand U1988 (N_1988,N_1865,N_1894);
and U1989 (N_1989,N_1854,N_1848);
xnor U1990 (N_1990,N_1846,N_1937);
or U1991 (N_1991,N_1944,N_1874);
xnor U1992 (N_1992,N_1903,N_1835);
and U1993 (N_1993,N_1869,N_1850);
xor U1994 (N_1994,N_1834,N_1849);
and U1995 (N_1995,N_1813,N_1905);
or U1996 (N_1996,N_1927,N_1853);
nand U1997 (N_1997,N_1888,N_1912);
and U1998 (N_1998,N_1890,N_1826);
nand U1999 (N_1999,N_1803,N_1841);
and U2000 (N_2000,N_1910,N_1839);
nor U2001 (N_2001,N_1857,N_1916);
or U2002 (N_2002,N_1948,N_1880);
or U2003 (N_2003,N_1867,N_1906);
and U2004 (N_2004,N_1918,N_1947);
xor U2005 (N_2005,N_1924,N_1911);
nor U2006 (N_2006,N_1852,N_1856);
nor U2007 (N_2007,N_1855,N_1878);
nand U2008 (N_2008,N_1868,N_1816);
or U2009 (N_2009,N_1805,N_1864);
nor U2010 (N_2010,N_1844,N_1939);
and U2011 (N_2011,N_1819,N_1940);
nand U2012 (N_2012,N_1915,N_1863);
or U2013 (N_2013,N_1934,N_1843);
xnor U2014 (N_2014,N_1811,N_1860);
xnor U2015 (N_2015,N_1872,N_1824);
nand U2016 (N_2016,N_1837,N_1933);
and U2017 (N_2017,N_1879,N_1825);
and U2018 (N_2018,N_1892,N_1875);
and U2019 (N_2019,N_1945,N_1832);
nand U2020 (N_2020,N_1815,N_1858);
and U2021 (N_2021,N_1866,N_1926);
nand U2022 (N_2022,N_1895,N_1901);
nand U2023 (N_2023,N_1809,N_1898);
and U2024 (N_2024,N_1842,N_1904);
nor U2025 (N_2025,N_1899,N_1817);
xnor U2026 (N_2026,N_1839,N_1918);
nor U2027 (N_2027,N_1855,N_1807);
or U2028 (N_2028,N_1931,N_1802);
nor U2029 (N_2029,N_1808,N_1905);
nor U2030 (N_2030,N_1849,N_1940);
or U2031 (N_2031,N_1809,N_1854);
or U2032 (N_2032,N_1935,N_1809);
or U2033 (N_2033,N_1838,N_1873);
and U2034 (N_2034,N_1819,N_1910);
xor U2035 (N_2035,N_1901,N_1876);
or U2036 (N_2036,N_1868,N_1914);
and U2037 (N_2037,N_1935,N_1944);
nor U2038 (N_2038,N_1807,N_1932);
xor U2039 (N_2039,N_1832,N_1858);
xnor U2040 (N_2040,N_1847,N_1906);
or U2041 (N_2041,N_1826,N_1895);
xnor U2042 (N_2042,N_1839,N_1836);
nand U2043 (N_2043,N_1907,N_1807);
or U2044 (N_2044,N_1935,N_1841);
nand U2045 (N_2045,N_1942,N_1891);
nor U2046 (N_2046,N_1898,N_1819);
nand U2047 (N_2047,N_1809,N_1848);
or U2048 (N_2048,N_1860,N_1943);
nand U2049 (N_2049,N_1821,N_1828);
xor U2050 (N_2050,N_1859,N_1894);
nand U2051 (N_2051,N_1904,N_1920);
and U2052 (N_2052,N_1900,N_1887);
or U2053 (N_2053,N_1844,N_1818);
or U2054 (N_2054,N_1918,N_1917);
nand U2055 (N_2055,N_1876,N_1828);
nor U2056 (N_2056,N_1876,N_1816);
nor U2057 (N_2057,N_1949,N_1824);
or U2058 (N_2058,N_1910,N_1915);
nor U2059 (N_2059,N_1854,N_1818);
nor U2060 (N_2060,N_1818,N_1851);
xnor U2061 (N_2061,N_1889,N_1894);
or U2062 (N_2062,N_1826,N_1914);
nand U2063 (N_2063,N_1946,N_1878);
nor U2064 (N_2064,N_1942,N_1896);
and U2065 (N_2065,N_1887,N_1825);
nor U2066 (N_2066,N_1830,N_1848);
nand U2067 (N_2067,N_1830,N_1824);
nor U2068 (N_2068,N_1844,N_1833);
and U2069 (N_2069,N_1817,N_1914);
and U2070 (N_2070,N_1944,N_1804);
xor U2071 (N_2071,N_1934,N_1901);
and U2072 (N_2072,N_1935,N_1832);
nor U2073 (N_2073,N_1866,N_1844);
nor U2074 (N_2074,N_1846,N_1862);
and U2075 (N_2075,N_1895,N_1839);
and U2076 (N_2076,N_1897,N_1840);
nor U2077 (N_2077,N_1900,N_1924);
and U2078 (N_2078,N_1817,N_1888);
xor U2079 (N_2079,N_1874,N_1942);
nor U2080 (N_2080,N_1855,N_1940);
and U2081 (N_2081,N_1831,N_1821);
and U2082 (N_2082,N_1832,N_1842);
nor U2083 (N_2083,N_1850,N_1944);
nor U2084 (N_2084,N_1808,N_1847);
and U2085 (N_2085,N_1802,N_1843);
and U2086 (N_2086,N_1861,N_1832);
or U2087 (N_2087,N_1889,N_1817);
and U2088 (N_2088,N_1854,N_1810);
or U2089 (N_2089,N_1919,N_1800);
nor U2090 (N_2090,N_1931,N_1896);
or U2091 (N_2091,N_1870,N_1873);
or U2092 (N_2092,N_1831,N_1942);
and U2093 (N_2093,N_1867,N_1822);
nor U2094 (N_2094,N_1941,N_1827);
xnor U2095 (N_2095,N_1920,N_1837);
xnor U2096 (N_2096,N_1949,N_1871);
and U2097 (N_2097,N_1876,N_1939);
xnor U2098 (N_2098,N_1856,N_1808);
or U2099 (N_2099,N_1873,N_1859);
xnor U2100 (N_2100,N_2078,N_2096);
nor U2101 (N_2101,N_2022,N_2032);
xnor U2102 (N_2102,N_2010,N_1950);
nor U2103 (N_2103,N_2057,N_1980);
nor U2104 (N_2104,N_2088,N_1981);
or U2105 (N_2105,N_2074,N_1961);
and U2106 (N_2106,N_2049,N_2089);
nand U2107 (N_2107,N_2060,N_2021);
xor U2108 (N_2108,N_2084,N_2018);
and U2109 (N_2109,N_1966,N_1973);
nor U2110 (N_2110,N_2005,N_2056);
nor U2111 (N_2111,N_2086,N_1968);
xnor U2112 (N_2112,N_1986,N_2027);
and U2113 (N_2113,N_2079,N_2071);
and U2114 (N_2114,N_1985,N_2004);
nand U2115 (N_2115,N_1974,N_2045);
nand U2116 (N_2116,N_2009,N_2034);
nor U2117 (N_2117,N_2041,N_2043);
nand U2118 (N_2118,N_2001,N_2047);
and U2119 (N_2119,N_2091,N_2007);
and U2120 (N_2120,N_2037,N_2092);
nor U2121 (N_2121,N_2019,N_2082);
xnor U2122 (N_2122,N_2099,N_2023);
and U2123 (N_2123,N_1953,N_1997);
and U2124 (N_2124,N_2024,N_2076);
nor U2125 (N_2125,N_2058,N_1963);
xnor U2126 (N_2126,N_2000,N_1951);
and U2127 (N_2127,N_2085,N_1960);
nor U2128 (N_2128,N_2053,N_1954);
and U2129 (N_2129,N_1958,N_2063);
nand U2130 (N_2130,N_2069,N_1990);
xnor U2131 (N_2131,N_2042,N_1994);
nand U2132 (N_2132,N_2039,N_2012);
xnor U2133 (N_2133,N_2097,N_2038);
nor U2134 (N_2134,N_2051,N_2017);
and U2135 (N_2135,N_2093,N_1955);
and U2136 (N_2136,N_2064,N_2026);
nand U2137 (N_2137,N_2025,N_2059);
and U2138 (N_2138,N_2080,N_2052);
nand U2139 (N_2139,N_1987,N_1962);
nand U2140 (N_2140,N_2048,N_2016);
xor U2141 (N_2141,N_1957,N_2072);
and U2142 (N_2142,N_1959,N_1952);
xor U2143 (N_2143,N_2095,N_2081);
xor U2144 (N_2144,N_1967,N_1969);
nand U2145 (N_2145,N_2062,N_2046);
xnor U2146 (N_2146,N_1998,N_2030);
nand U2147 (N_2147,N_2044,N_2066);
nor U2148 (N_2148,N_2029,N_1989);
and U2149 (N_2149,N_2008,N_2031);
and U2150 (N_2150,N_1956,N_1965);
and U2151 (N_2151,N_1988,N_2073);
nor U2152 (N_2152,N_2054,N_1978);
or U2153 (N_2153,N_1996,N_2055);
nor U2154 (N_2154,N_2061,N_2011);
or U2155 (N_2155,N_2033,N_1993);
nor U2156 (N_2156,N_1984,N_2075);
and U2157 (N_2157,N_1976,N_2098);
and U2158 (N_2158,N_1995,N_1975);
and U2159 (N_2159,N_1977,N_2087);
nand U2160 (N_2160,N_1999,N_2050);
and U2161 (N_2161,N_1964,N_1972);
nand U2162 (N_2162,N_2077,N_2014);
and U2163 (N_2163,N_1979,N_1983);
or U2164 (N_2164,N_1970,N_2013);
nor U2165 (N_2165,N_2015,N_2083);
nand U2166 (N_2166,N_1992,N_1971);
or U2167 (N_2167,N_2006,N_2002);
and U2168 (N_2168,N_2065,N_2090);
xnor U2169 (N_2169,N_1991,N_2040);
nor U2170 (N_2170,N_2028,N_2094);
xor U2171 (N_2171,N_2020,N_2068);
xnor U2172 (N_2172,N_2003,N_1982);
xor U2173 (N_2173,N_2035,N_2067);
and U2174 (N_2174,N_2036,N_2070);
and U2175 (N_2175,N_2093,N_2016);
and U2176 (N_2176,N_2027,N_2032);
and U2177 (N_2177,N_2092,N_2022);
nor U2178 (N_2178,N_2071,N_2032);
and U2179 (N_2179,N_2092,N_2096);
nand U2180 (N_2180,N_2053,N_1951);
or U2181 (N_2181,N_2030,N_1968);
nor U2182 (N_2182,N_2074,N_2073);
and U2183 (N_2183,N_2054,N_1972);
xnor U2184 (N_2184,N_1996,N_2039);
nor U2185 (N_2185,N_1952,N_1983);
nand U2186 (N_2186,N_1966,N_2024);
nand U2187 (N_2187,N_2087,N_1954);
nor U2188 (N_2188,N_2091,N_1964);
nand U2189 (N_2189,N_2036,N_2082);
nor U2190 (N_2190,N_2005,N_2014);
xnor U2191 (N_2191,N_1980,N_2045);
and U2192 (N_2192,N_2043,N_2019);
nor U2193 (N_2193,N_2052,N_2021);
or U2194 (N_2194,N_2024,N_1961);
nand U2195 (N_2195,N_1967,N_2047);
and U2196 (N_2196,N_1996,N_2051);
or U2197 (N_2197,N_2017,N_2058);
xor U2198 (N_2198,N_2034,N_2054);
nand U2199 (N_2199,N_1951,N_2036);
xnor U2200 (N_2200,N_1991,N_1968);
xor U2201 (N_2201,N_2062,N_2024);
or U2202 (N_2202,N_2075,N_1968);
or U2203 (N_2203,N_1964,N_2027);
nand U2204 (N_2204,N_2082,N_1969);
xnor U2205 (N_2205,N_1965,N_2081);
nand U2206 (N_2206,N_2019,N_2083);
and U2207 (N_2207,N_1980,N_2041);
nand U2208 (N_2208,N_2064,N_1993);
xnor U2209 (N_2209,N_2078,N_2052);
or U2210 (N_2210,N_2032,N_2063);
and U2211 (N_2211,N_2029,N_2093);
nor U2212 (N_2212,N_1956,N_2024);
and U2213 (N_2213,N_1966,N_1984);
and U2214 (N_2214,N_2029,N_2054);
or U2215 (N_2215,N_1986,N_2065);
nand U2216 (N_2216,N_2083,N_1959);
or U2217 (N_2217,N_2066,N_2061);
nand U2218 (N_2218,N_2088,N_2016);
or U2219 (N_2219,N_2072,N_2068);
or U2220 (N_2220,N_2079,N_2049);
and U2221 (N_2221,N_2020,N_2006);
nand U2222 (N_2222,N_2026,N_2036);
and U2223 (N_2223,N_2013,N_2082);
or U2224 (N_2224,N_1960,N_2046);
nand U2225 (N_2225,N_1953,N_1998);
or U2226 (N_2226,N_2028,N_2034);
xnor U2227 (N_2227,N_1950,N_1998);
nor U2228 (N_2228,N_2046,N_2003);
or U2229 (N_2229,N_2069,N_1957);
and U2230 (N_2230,N_2033,N_2050);
nand U2231 (N_2231,N_2037,N_1993);
nor U2232 (N_2232,N_2025,N_2056);
or U2233 (N_2233,N_2074,N_2086);
or U2234 (N_2234,N_1983,N_1989);
xnor U2235 (N_2235,N_1991,N_2043);
nor U2236 (N_2236,N_2063,N_2011);
nand U2237 (N_2237,N_2033,N_2091);
and U2238 (N_2238,N_2072,N_2022);
nand U2239 (N_2239,N_2001,N_1950);
or U2240 (N_2240,N_2041,N_2082);
xor U2241 (N_2241,N_1992,N_2004);
or U2242 (N_2242,N_1957,N_1958);
nor U2243 (N_2243,N_2032,N_2086);
and U2244 (N_2244,N_2096,N_1974);
and U2245 (N_2245,N_2066,N_2004);
nor U2246 (N_2246,N_2008,N_1969);
nor U2247 (N_2247,N_2070,N_2011);
nor U2248 (N_2248,N_1959,N_2082);
xnor U2249 (N_2249,N_1988,N_1950);
nand U2250 (N_2250,N_2224,N_2232);
nor U2251 (N_2251,N_2170,N_2102);
and U2252 (N_2252,N_2248,N_2128);
nor U2253 (N_2253,N_2180,N_2187);
nor U2254 (N_2254,N_2209,N_2111);
xor U2255 (N_2255,N_2117,N_2199);
nor U2256 (N_2256,N_2140,N_2197);
nand U2257 (N_2257,N_2127,N_2139);
and U2258 (N_2258,N_2191,N_2115);
or U2259 (N_2259,N_2112,N_2129);
nor U2260 (N_2260,N_2107,N_2132);
nand U2261 (N_2261,N_2223,N_2233);
xor U2262 (N_2262,N_2175,N_2100);
or U2263 (N_2263,N_2242,N_2103);
xor U2264 (N_2264,N_2169,N_2122);
xnor U2265 (N_2265,N_2196,N_2167);
nor U2266 (N_2266,N_2229,N_2190);
nand U2267 (N_2267,N_2125,N_2130);
and U2268 (N_2268,N_2154,N_2245);
and U2269 (N_2269,N_2135,N_2227);
xor U2270 (N_2270,N_2240,N_2219);
xor U2271 (N_2271,N_2136,N_2104);
and U2272 (N_2272,N_2145,N_2124);
or U2273 (N_2273,N_2147,N_2247);
and U2274 (N_2274,N_2174,N_2106);
nand U2275 (N_2275,N_2237,N_2194);
nor U2276 (N_2276,N_2173,N_2118);
xor U2277 (N_2277,N_2214,N_2109);
or U2278 (N_2278,N_2121,N_2171);
and U2279 (N_2279,N_2211,N_2220);
and U2280 (N_2280,N_2243,N_2179);
xnor U2281 (N_2281,N_2105,N_2207);
and U2282 (N_2282,N_2108,N_2119);
and U2283 (N_2283,N_2114,N_2182);
or U2284 (N_2284,N_2120,N_2158);
and U2285 (N_2285,N_2164,N_2153);
nand U2286 (N_2286,N_2210,N_2188);
nor U2287 (N_2287,N_2146,N_2244);
nand U2288 (N_2288,N_2217,N_2215);
nand U2289 (N_2289,N_2181,N_2131);
and U2290 (N_2290,N_2177,N_2221);
nor U2291 (N_2291,N_2116,N_2249);
xor U2292 (N_2292,N_2138,N_2226);
or U2293 (N_2293,N_2208,N_2113);
nand U2294 (N_2294,N_2151,N_2212);
nor U2295 (N_2295,N_2141,N_2205);
xnor U2296 (N_2296,N_2178,N_2168);
and U2297 (N_2297,N_2234,N_2101);
and U2298 (N_2298,N_2241,N_2201);
or U2299 (N_2299,N_2239,N_2192);
nand U2300 (N_2300,N_2200,N_2189);
and U2301 (N_2301,N_2184,N_2213);
nand U2302 (N_2302,N_2163,N_2159);
and U2303 (N_2303,N_2246,N_2142);
or U2304 (N_2304,N_2155,N_2123);
nand U2305 (N_2305,N_2149,N_2231);
nor U2306 (N_2306,N_2236,N_2193);
nor U2307 (N_2307,N_2156,N_2218);
and U2308 (N_2308,N_2204,N_2216);
or U2309 (N_2309,N_2152,N_2143);
and U2310 (N_2310,N_2161,N_2186);
nor U2311 (N_2311,N_2133,N_2150);
and U2312 (N_2312,N_2165,N_2203);
xor U2313 (N_2313,N_2235,N_2206);
nand U2314 (N_2314,N_2172,N_2225);
or U2315 (N_2315,N_2198,N_2157);
or U2316 (N_2316,N_2195,N_2230);
nand U2317 (N_2317,N_2183,N_2144);
xnor U2318 (N_2318,N_2222,N_2137);
or U2319 (N_2319,N_2126,N_2160);
nor U2320 (N_2320,N_2176,N_2185);
nand U2321 (N_2321,N_2238,N_2110);
or U2322 (N_2322,N_2228,N_2166);
or U2323 (N_2323,N_2148,N_2134);
nand U2324 (N_2324,N_2202,N_2162);
and U2325 (N_2325,N_2222,N_2239);
xnor U2326 (N_2326,N_2145,N_2130);
and U2327 (N_2327,N_2236,N_2179);
xnor U2328 (N_2328,N_2100,N_2248);
xor U2329 (N_2329,N_2120,N_2144);
nor U2330 (N_2330,N_2132,N_2204);
or U2331 (N_2331,N_2109,N_2225);
and U2332 (N_2332,N_2223,N_2234);
nor U2333 (N_2333,N_2184,N_2166);
or U2334 (N_2334,N_2178,N_2165);
nand U2335 (N_2335,N_2153,N_2158);
nand U2336 (N_2336,N_2143,N_2232);
nor U2337 (N_2337,N_2118,N_2116);
or U2338 (N_2338,N_2186,N_2165);
nor U2339 (N_2339,N_2232,N_2171);
nor U2340 (N_2340,N_2119,N_2144);
nor U2341 (N_2341,N_2120,N_2197);
or U2342 (N_2342,N_2231,N_2103);
or U2343 (N_2343,N_2108,N_2193);
or U2344 (N_2344,N_2241,N_2149);
xnor U2345 (N_2345,N_2231,N_2185);
or U2346 (N_2346,N_2233,N_2202);
or U2347 (N_2347,N_2194,N_2145);
xor U2348 (N_2348,N_2185,N_2244);
xnor U2349 (N_2349,N_2226,N_2123);
nand U2350 (N_2350,N_2135,N_2205);
xnor U2351 (N_2351,N_2190,N_2242);
xnor U2352 (N_2352,N_2123,N_2177);
xor U2353 (N_2353,N_2143,N_2185);
xor U2354 (N_2354,N_2127,N_2192);
or U2355 (N_2355,N_2186,N_2108);
xnor U2356 (N_2356,N_2157,N_2142);
nor U2357 (N_2357,N_2229,N_2169);
xor U2358 (N_2358,N_2144,N_2216);
nand U2359 (N_2359,N_2230,N_2192);
nor U2360 (N_2360,N_2125,N_2210);
or U2361 (N_2361,N_2105,N_2158);
and U2362 (N_2362,N_2159,N_2174);
nand U2363 (N_2363,N_2115,N_2106);
or U2364 (N_2364,N_2195,N_2236);
nor U2365 (N_2365,N_2110,N_2209);
nand U2366 (N_2366,N_2173,N_2130);
nand U2367 (N_2367,N_2109,N_2106);
or U2368 (N_2368,N_2145,N_2222);
and U2369 (N_2369,N_2223,N_2220);
or U2370 (N_2370,N_2144,N_2191);
or U2371 (N_2371,N_2124,N_2246);
nand U2372 (N_2372,N_2198,N_2100);
nor U2373 (N_2373,N_2107,N_2133);
or U2374 (N_2374,N_2188,N_2172);
and U2375 (N_2375,N_2128,N_2122);
and U2376 (N_2376,N_2154,N_2107);
and U2377 (N_2377,N_2117,N_2165);
nand U2378 (N_2378,N_2155,N_2208);
or U2379 (N_2379,N_2193,N_2169);
or U2380 (N_2380,N_2211,N_2167);
or U2381 (N_2381,N_2171,N_2175);
xnor U2382 (N_2382,N_2140,N_2178);
or U2383 (N_2383,N_2178,N_2139);
or U2384 (N_2384,N_2224,N_2196);
xor U2385 (N_2385,N_2230,N_2209);
xor U2386 (N_2386,N_2196,N_2150);
nor U2387 (N_2387,N_2154,N_2151);
xnor U2388 (N_2388,N_2101,N_2214);
or U2389 (N_2389,N_2100,N_2206);
nand U2390 (N_2390,N_2193,N_2229);
nor U2391 (N_2391,N_2225,N_2244);
or U2392 (N_2392,N_2212,N_2190);
xnor U2393 (N_2393,N_2208,N_2188);
and U2394 (N_2394,N_2190,N_2214);
nor U2395 (N_2395,N_2242,N_2182);
nand U2396 (N_2396,N_2174,N_2136);
or U2397 (N_2397,N_2160,N_2184);
or U2398 (N_2398,N_2240,N_2221);
xor U2399 (N_2399,N_2130,N_2178);
or U2400 (N_2400,N_2310,N_2258);
nand U2401 (N_2401,N_2357,N_2380);
or U2402 (N_2402,N_2277,N_2397);
xor U2403 (N_2403,N_2286,N_2331);
and U2404 (N_2404,N_2349,N_2253);
nand U2405 (N_2405,N_2392,N_2342);
or U2406 (N_2406,N_2263,N_2291);
or U2407 (N_2407,N_2303,N_2276);
nand U2408 (N_2408,N_2382,N_2289);
or U2409 (N_2409,N_2371,N_2295);
nor U2410 (N_2410,N_2312,N_2294);
nand U2411 (N_2411,N_2290,N_2302);
nor U2412 (N_2412,N_2255,N_2320);
nand U2413 (N_2413,N_2254,N_2298);
nand U2414 (N_2414,N_2370,N_2348);
or U2415 (N_2415,N_2364,N_2259);
nor U2416 (N_2416,N_2285,N_2318);
or U2417 (N_2417,N_2306,N_2372);
and U2418 (N_2418,N_2360,N_2262);
and U2419 (N_2419,N_2361,N_2338);
nor U2420 (N_2420,N_2250,N_2278);
and U2421 (N_2421,N_2282,N_2251);
xnor U2422 (N_2422,N_2396,N_2313);
nand U2423 (N_2423,N_2288,N_2319);
and U2424 (N_2424,N_2346,N_2381);
and U2425 (N_2425,N_2390,N_2307);
xor U2426 (N_2426,N_2356,N_2261);
nor U2427 (N_2427,N_2374,N_2353);
xor U2428 (N_2428,N_2293,N_2299);
nand U2429 (N_2429,N_2367,N_2332);
or U2430 (N_2430,N_2350,N_2383);
or U2431 (N_2431,N_2369,N_2373);
xnor U2432 (N_2432,N_2340,N_2337);
and U2433 (N_2433,N_2354,N_2375);
or U2434 (N_2434,N_2399,N_2386);
nand U2435 (N_2435,N_2268,N_2351);
and U2436 (N_2436,N_2335,N_2292);
nor U2437 (N_2437,N_2398,N_2344);
nand U2438 (N_2438,N_2378,N_2347);
or U2439 (N_2439,N_2265,N_2385);
nand U2440 (N_2440,N_2273,N_2274);
nand U2441 (N_2441,N_2287,N_2300);
or U2442 (N_2442,N_2322,N_2297);
xnor U2443 (N_2443,N_2366,N_2264);
nand U2444 (N_2444,N_2256,N_2393);
and U2445 (N_2445,N_2363,N_2267);
nor U2446 (N_2446,N_2391,N_2341);
nor U2447 (N_2447,N_2362,N_2368);
nor U2448 (N_2448,N_2394,N_2326);
xor U2449 (N_2449,N_2389,N_2321);
nand U2450 (N_2450,N_2266,N_2305);
or U2451 (N_2451,N_2325,N_2333);
and U2452 (N_2452,N_2352,N_2309);
and U2453 (N_2453,N_2315,N_2275);
or U2454 (N_2454,N_2296,N_2324);
nand U2455 (N_2455,N_2272,N_2387);
nand U2456 (N_2456,N_2334,N_2304);
nor U2457 (N_2457,N_2327,N_2388);
or U2458 (N_2458,N_2365,N_2345);
xor U2459 (N_2459,N_2270,N_2280);
or U2460 (N_2460,N_2252,N_2311);
xnor U2461 (N_2461,N_2316,N_2269);
or U2462 (N_2462,N_2358,N_2359);
nor U2463 (N_2463,N_2279,N_2377);
nor U2464 (N_2464,N_2260,N_2379);
nor U2465 (N_2465,N_2283,N_2330);
xnor U2466 (N_2466,N_2301,N_2308);
nand U2467 (N_2467,N_2257,N_2395);
nor U2468 (N_2468,N_2336,N_2339);
and U2469 (N_2469,N_2284,N_2355);
and U2470 (N_2470,N_2281,N_2376);
and U2471 (N_2471,N_2314,N_2317);
xnor U2472 (N_2472,N_2271,N_2328);
nor U2473 (N_2473,N_2329,N_2343);
and U2474 (N_2474,N_2323,N_2384);
nand U2475 (N_2475,N_2381,N_2312);
and U2476 (N_2476,N_2287,N_2272);
nor U2477 (N_2477,N_2322,N_2290);
nor U2478 (N_2478,N_2360,N_2396);
nand U2479 (N_2479,N_2294,N_2320);
nor U2480 (N_2480,N_2274,N_2293);
nor U2481 (N_2481,N_2395,N_2384);
xnor U2482 (N_2482,N_2387,N_2338);
and U2483 (N_2483,N_2383,N_2299);
and U2484 (N_2484,N_2300,N_2282);
nor U2485 (N_2485,N_2399,N_2306);
and U2486 (N_2486,N_2320,N_2295);
and U2487 (N_2487,N_2314,N_2367);
nor U2488 (N_2488,N_2285,N_2354);
and U2489 (N_2489,N_2390,N_2263);
and U2490 (N_2490,N_2297,N_2382);
nor U2491 (N_2491,N_2364,N_2282);
xor U2492 (N_2492,N_2329,N_2301);
nor U2493 (N_2493,N_2304,N_2368);
nand U2494 (N_2494,N_2291,N_2390);
nand U2495 (N_2495,N_2255,N_2372);
nand U2496 (N_2496,N_2258,N_2349);
nand U2497 (N_2497,N_2287,N_2286);
xor U2498 (N_2498,N_2393,N_2394);
nor U2499 (N_2499,N_2363,N_2316);
nand U2500 (N_2500,N_2312,N_2290);
and U2501 (N_2501,N_2274,N_2278);
or U2502 (N_2502,N_2350,N_2381);
nand U2503 (N_2503,N_2287,N_2390);
or U2504 (N_2504,N_2294,N_2282);
nand U2505 (N_2505,N_2369,N_2340);
nand U2506 (N_2506,N_2266,N_2388);
or U2507 (N_2507,N_2307,N_2361);
nand U2508 (N_2508,N_2327,N_2329);
nor U2509 (N_2509,N_2344,N_2290);
or U2510 (N_2510,N_2274,N_2252);
xor U2511 (N_2511,N_2348,N_2394);
nor U2512 (N_2512,N_2306,N_2351);
and U2513 (N_2513,N_2348,N_2287);
nand U2514 (N_2514,N_2305,N_2320);
nor U2515 (N_2515,N_2318,N_2292);
or U2516 (N_2516,N_2354,N_2368);
nand U2517 (N_2517,N_2266,N_2394);
and U2518 (N_2518,N_2381,N_2326);
or U2519 (N_2519,N_2378,N_2390);
and U2520 (N_2520,N_2300,N_2393);
or U2521 (N_2521,N_2261,N_2335);
or U2522 (N_2522,N_2335,N_2390);
nand U2523 (N_2523,N_2253,N_2323);
nor U2524 (N_2524,N_2305,N_2370);
and U2525 (N_2525,N_2366,N_2313);
or U2526 (N_2526,N_2356,N_2277);
xnor U2527 (N_2527,N_2310,N_2378);
nand U2528 (N_2528,N_2336,N_2381);
nand U2529 (N_2529,N_2252,N_2262);
or U2530 (N_2530,N_2387,N_2291);
xnor U2531 (N_2531,N_2296,N_2339);
or U2532 (N_2532,N_2308,N_2376);
xnor U2533 (N_2533,N_2398,N_2277);
and U2534 (N_2534,N_2359,N_2264);
and U2535 (N_2535,N_2349,N_2336);
nand U2536 (N_2536,N_2310,N_2329);
and U2537 (N_2537,N_2295,N_2251);
or U2538 (N_2538,N_2354,N_2270);
and U2539 (N_2539,N_2304,N_2391);
or U2540 (N_2540,N_2397,N_2267);
and U2541 (N_2541,N_2384,N_2271);
xor U2542 (N_2542,N_2384,N_2262);
nand U2543 (N_2543,N_2323,N_2258);
nor U2544 (N_2544,N_2281,N_2270);
xnor U2545 (N_2545,N_2276,N_2374);
nand U2546 (N_2546,N_2349,N_2366);
nand U2547 (N_2547,N_2356,N_2373);
or U2548 (N_2548,N_2337,N_2391);
and U2549 (N_2549,N_2357,N_2290);
nand U2550 (N_2550,N_2443,N_2512);
nand U2551 (N_2551,N_2472,N_2471);
nand U2552 (N_2552,N_2425,N_2493);
nor U2553 (N_2553,N_2439,N_2505);
or U2554 (N_2554,N_2547,N_2477);
nor U2555 (N_2555,N_2401,N_2453);
nand U2556 (N_2556,N_2460,N_2458);
xnor U2557 (N_2557,N_2464,N_2468);
xor U2558 (N_2558,N_2499,N_2543);
xnor U2559 (N_2559,N_2402,N_2495);
and U2560 (N_2560,N_2422,N_2545);
nor U2561 (N_2561,N_2410,N_2414);
nand U2562 (N_2562,N_2544,N_2549);
nor U2563 (N_2563,N_2409,N_2527);
xor U2564 (N_2564,N_2548,N_2537);
nand U2565 (N_2565,N_2481,N_2430);
xor U2566 (N_2566,N_2514,N_2429);
nor U2567 (N_2567,N_2497,N_2488);
or U2568 (N_2568,N_2475,N_2489);
nand U2569 (N_2569,N_2442,N_2516);
nor U2570 (N_2570,N_2513,N_2435);
nor U2571 (N_2571,N_2419,N_2426);
nand U2572 (N_2572,N_2522,N_2541);
xor U2573 (N_2573,N_2529,N_2519);
and U2574 (N_2574,N_2517,N_2530);
or U2575 (N_2575,N_2539,N_2417);
and U2576 (N_2576,N_2504,N_2482);
and U2577 (N_2577,N_2445,N_2463);
or U2578 (N_2578,N_2540,N_2491);
or U2579 (N_2579,N_2487,N_2474);
nand U2580 (N_2580,N_2492,N_2415);
nor U2581 (N_2581,N_2452,N_2420);
nor U2582 (N_2582,N_2434,N_2501);
or U2583 (N_2583,N_2534,N_2450);
xnor U2584 (N_2584,N_2418,N_2427);
nand U2585 (N_2585,N_2479,N_2500);
nand U2586 (N_2586,N_2538,N_2400);
or U2587 (N_2587,N_2525,N_2428);
xor U2588 (N_2588,N_2432,N_2451);
nand U2589 (N_2589,N_2531,N_2456);
xnor U2590 (N_2590,N_2421,N_2476);
and U2591 (N_2591,N_2508,N_2467);
and U2592 (N_2592,N_2405,N_2502);
xnor U2593 (N_2593,N_2457,N_2511);
and U2594 (N_2594,N_2473,N_2510);
or U2595 (N_2595,N_2446,N_2403);
xor U2596 (N_2596,N_2546,N_2536);
or U2597 (N_2597,N_2424,N_2532);
and U2598 (N_2598,N_2515,N_2485);
and U2599 (N_2599,N_2483,N_2521);
nor U2600 (N_2600,N_2447,N_2412);
nor U2601 (N_2601,N_2518,N_2433);
nand U2602 (N_2602,N_2454,N_2486);
and U2603 (N_2603,N_2509,N_2484);
nand U2604 (N_2604,N_2407,N_2503);
xor U2605 (N_2605,N_2423,N_2413);
xnor U2606 (N_2606,N_2438,N_2526);
and U2607 (N_2607,N_2478,N_2480);
nand U2608 (N_2608,N_2455,N_2524);
xnor U2609 (N_2609,N_2449,N_2440);
nand U2610 (N_2610,N_2461,N_2462);
nor U2611 (N_2611,N_2465,N_2404);
nor U2612 (N_2612,N_2528,N_2411);
or U2613 (N_2613,N_2490,N_2469);
xnor U2614 (N_2614,N_2496,N_2408);
xnor U2615 (N_2615,N_2441,N_2444);
nor U2616 (N_2616,N_2448,N_2535);
and U2617 (N_2617,N_2520,N_2436);
xor U2618 (N_2618,N_2466,N_2431);
or U2619 (N_2619,N_2498,N_2506);
nor U2620 (N_2620,N_2437,N_2459);
or U2621 (N_2621,N_2533,N_2406);
or U2622 (N_2622,N_2494,N_2470);
and U2623 (N_2623,N_2542,N_2416);
or U2624 (N_2624,N_2523,N_2507);
or U2625 (N_2625,N_2501,N_2400);
nor U2626 (N_2626,N_2507,N_2511);
nand U2627 (N_2627,N_2502,N_2431);
nor U2628 (N_2628,N_2430,N_2418);
xnor U2629 (N_2629,N_2405,N_2474);
nand U2630 (N_2630,N_2430,N_2419);
nand U2631 (N_2631,N_2427,N_2494);
nand U2632 (N_2632,N_2511,N_2470);
xnor U2633 (N_2633,N_2467,N_2517);
or U2634 (N_2634,N_2465,N_2477);
xnor U2635 (N_2635,N_2479,N_2480);
nor U2636 (N_2636,N_2447,N_2401);
nand U2637 (N_2637,N_2450,N_2467);
nor U2638 (N_2638,N_2479,N_2521);
and U2639 (N_2639,N_2440,N_2468);
nor U2640 (N_2640,N_2539,N_2542);
and U2641 (N_2641,N_2504,N_2457);
xnor U2642 (N_2642,N_2498,N_2410);
nand U2643 (N_2643,N_2425,N_2409);
xnor U2644 (N_2644,N_2533,N_2409);
nand U2645 (N_2645,N_2461,N_2401);
nor U2646 (N_2646,N_2505,N_2509);
nand U2647 (N_2647,N_2442,N_2444);
nor U2648 (N_2648,N_2548,N_2422);
and U2649 (N_2649,N_2528,N_2462);
and U2650 (N_2650,N_2480,N_2438);
or U2651 (N_2651,N_2426,N_2400);
and U2652 (N_2652,N_2522,N_2523);
nand U2653 (N_2653,N_2541,N_2444);
nand U2654 (N_2654,N_2451,N_2428);
xor U2655 (N_2655,N_2422,N_2499);
xnor U2656 (N_2656,N_2491,N_2500);
and U2657 (N_2657,N_2476,N_2497);
xnor U2658 (N_2658,N_2433,N_2526);
and U2659 (N_2659,N_2499,N_2500);
nor U2660 (N_2660,N_2433,N_2419);
xor U2661 (N_2661,N_2544,N_2451);
nand U2662 (N_2662,N_2459,N_2421);
nor U2663 (N_2663,N_2549,N_2487);
nand U2664 (N_2664,N_2492,N_2491);
or U2665 (N_2665,N_2500,N_2428);
and U2666 (N_2666,N_2536,N_2496);
and U2667 (N_2667,N_2510,N_2439);
and U2668 (N_2668,N_2426,N_2464);
xnor U2669 (N_2669,N_2487,N_2452);
and U2670 (N_2670,N_2540,N_2421);
and U2671 (N_2671,N_2411,N_2454);
xor U2672 (N_2672,N_2498,N_2497);
nor U2673 (N_2673,N_2453,N_2457);
and U2674 (N_2674,N_2537,N_2436);
or U2675 (N_2675,N_2462,N_2548);
nand U2676 (N_2676,N_2533,N_2544);
nor U2677 (N_2677,N_2525,N_2401);
and U2678 (N_2678,N_2423,N_2407);
nor U2679 (N_2679,N_2428,N_2493);
nand U2680 (N_2680,N_2463,N_2466);
nor U2681 (N_2681,N_2458,N_2464);
xor U2682 (N_2682,N_2503,N_2478);
or U2683 (N_2683,N_2520,N_2519);
or U2684 (N_2684,N_2436,N_2432);
xnor U2685 (N_2685,N_2508,N_2472);
and U2686 (N_2686,N_2464,N_2461);
or U2687 (N_2687,N_2549,N_2476);
nor U2688 (N_2688,N_2404,N_2476);
nor U2689 (N_2689,N_2444,N_2546);
and U2690 (N_2690,N_2411,N_2462);
nand U2691 (N_2691,N_2452,N_2524);
nor U2692 (N_2692,N_2450,N_2536);
xor U2693 (N_2693,N_2470,N_2477);
nor U2694 (N_2694,N_2439,N_2482);
nand U2695 (N_2695,N_2485,N_2486);
and U2696 (N_2696,N_2455,N_2431);
and U2697 (N_2697,N_2528,N_2492);
and U2698 (N_2698,N_2519,N_2491);
and U2699 (N_2699,N_2506,N_2502);
nor U2700 (N_2700,N_2641,N_2619);
or U2701 (N_2701,N_2614,N_2596);
nand U2702 (N_2702,N_2676,N_2670);
or U2703 (N_2703,N_2625,N_2660);
or U2704 (N_2704,N_2561,N_2569);
or U2705 (N_2705,N_2607,N_2620);
nor U2706 (N_2706,N_2680,N_2603);
xor U2707 (N_2707,N_2568,N_2677);
or U2708 (N_2708,N_2610,N_2593);
or U2709 (N_2709,N_2658,N_2585);
nand U2710 (N_2710,N_2692,N_2691);
or U2711 (N_2711,N_2693,N_2640);
nor U2712 (N_2712,N_2679,N_2590);
nor U2713 (N_2713,N_2555,N_2639);
and U2714 (N_2714,N_2674,N_2695);
and U2715 (N_2715,N_2635,N_2579);
xnor U2716 (N_2716,N_2652,N_2575);
nor U2717 (N_2717,N_2646,N_2554);
xor U2718 (N_2718,N_2591,N_2602);
xnor U2719 (N_2719,N_2638,N_2589);
nand U2720 (N_2720,N_2577,N_2557);
or U2721 (N_2721,N_2553,N_2664);
nand U2722 (N_2722,N_2694,N_2687);
xnor U2723 (N_2723,N_2583,N_2566);
and U2724 (N_2724,N_2690,N_2696);
nor U2725 (N_2725,N_2618,N_2653);
nand U2726 (N_2726,N_2616,N_2644);
and U2727 (N_2727,N_2651,N_2571);
nand U2728 (N_2728,N_2612,N_2661);
nand U2729 (N_2729,N_2552,N_2678);
nand U2730 (N_2730,N_2672,N_2592);
nor U2731 (N_2731,N_2605,N_2656);
xnor U2732 (N_2732,N_2580,N_2564);
xnor U2733 (N_2733,N_2617,N_2570);
xnor U2734 (N_2734,N_2645,N_2623);
xnor U2735 (N_2735,N_2599,N_2666);
or U2736 (N_2736,N_2634,N_2565);
xnor U2737 (N_2737,N_2560,N_2567);
nand U2738 (N_2738,N_2667,N_2576);
and U2739 (N_2739,N_2633,N_2584);
nand U2740 (N_2740,N_2626,N_2659);
nand U2741 (N_2741,N_2671,N_2594);
nand U2742 (N_2742,N_2588,N_2621);
nand U2743 (N_2743,N_2582,N_2628);
and U2744 (N_2744,N_2682,N_2647);
and U2745 (N_2745,N_2601,N_2636);
nand U2746 (N_2746,N_2632,N_2622);
nand U2747 (N_2747,N_2563,N_2688);
and U2748 (N_2748,N_2606,N_2663);
and U2749 (N_2749,N_2698,N_2574);
or U2750 (N_2750,N_2609,N_2551);
or U2751 (N_2751,N_2662,N_2699);
and U2752 (N_2752,N_2642,N_2598);
xor U2753 (N_2753,N_2572,N_2657);
nor U2754 (N_2754,N_2654,N_2686);
xnor U2755 (N_2755,N_2649,N_2665);
xor U2756 (N_2756,N_2558,N_2681);
or U2757 (N_2757,N_2556,N_2586);
or U2758 (N_2758,N_2629,N_2587);
xor U2759 (N_2759,N_2627,N_2615);
nor U2760 (N_2760,N_2600,N_2697);
nand U2761 (N_2761,N_2631,N_2595);
xor U2762 (N_2762,N_2648,N_2669);
xnor U2763 (N_2763,N_2578,N_2624);
and U2764 (N_2764,N_2573,N_2689);
nand U2765 (N_2765,N_2581,N_2630);
and U2766 (N_2766,N_2559,N_2675);
and U2767 (N_2767,N_2637,N_2604);
nand U2768 (N_2768,N_2562,N_2643);
xor U2769 (N_2769,N_2608,N_2668);
or U2770 (N_2770,N_2611,N_2597);
nor U2771 (N_2771,N_2655,N_2550);
nor U2772 (N_2772,N_2683,N_2650);
and U2773 (N_2773,N_2685,N_2684);
xnor U2774 (N_2774,N_2613,N_2673);
xor U2775 (N_2775,N_2644,N_2566);
nand U2776 (N_2776,N_2697,N_2625);
xor U2777 (N_2777,N_2617,N_2675);
and U2778 (N_2778,N_2599,N_2596);
nand U2779 (N_2779,N_2615,N_2575);
nand U2780 (N_2780,N_2638,N_2675);
or U2781 (N_2781,N_2586,N_2630);
or U2782 (N_2782,N_2554,N_2689);
and U2783 (N_2783,N_2565,N_2699);
xor U2784 (N_2784,N_2670,N_2585);
xnor U2785 (N_2785,N_2655,N_2631);
nor U2786 (N_2786,N_2644,N_2575);
nor U2787 (N_2787,N_2677,N_2576);
or U2788 (N_2788,N_2582,N_2622);
nor U2789 (N_2789,N_2613,N_2664);
and U2790 (N_2790,N_2582,N_2619);
and U2791 (N_2791,N_2644,N_2678);
xor U2792 (N_2792,N_2615,N_2691);
nand U2793 (N_2793,N_2551,N_2621);
and U2794 (N_2794,N_2683,N_2657);
nand U2795 (N_2795,N_2644,N_2675);
xnor U2796 (N_2796,N_2612,N_2692);
and U2797 (N_2797,N_2567,N_2600);
or U2798 (N_2798,N_2637,N_2614);
nand U2799 (N_2799,N_2633,N_2646);
nor U2800 (N_2800,N_2596,N_2686);
or U2801 (N_2801,N_2685,N_2630);
and U2802 (N_2802,N_2609,N_2680);
and U2803 (N_2803,N_2625,N_2571);
nand U2804 (N_2804,N_2554,N_2550);
or U2805 (N_2805,N_2689,N_2641);
or U2806 (N_2806,N_2552,N_2613);
xnor U2807 (N_2807,N_2679,N_2586);
nor U2808 (N_2808,N_2580,N_2666);
xor U2809 (N_2809,N_2629,N_2610);
and U2810 (N_2810,N_2637,N_2699);
nor U2811 (N_2811,N_2632,N_2606);
nor U2812 (N_2812,N_2570,N_2624);
and U2813 (N_2813,N_2688,N_2696);
or U2814 (N_2814,N_2609,N_2599);
nor U2815 (N_2815,N_2630,N_2614);
nor U2816 (N_2816,N_2688,N_2609);
xor U2817 (N_2817,N_2605,N_2697);
and U2818 (N_2818,N_2576,N_2663);
nor U2819 (N_2819,N_2673,N_2589);
and U2820 (N_2820,N_2617,N_2686);
nor U2821 (N_2821,N_2563,N_2576);
xor U2822 (N_2822,N_2586,N_2687);
nand U2823 (N_2823,N_2585,N_2615);
and U2824 (N_2824,N_2686,N_2607);
or U2825 (N_2825,N_2621,N_2630);
and U2826 (N_2826,N_2609,N_2607);
xor U2827 (N_2827,N_2570,N_2582);
xor U2828 (N_2828,N_2650,N_2657);
nand U2829 (N_2829,N_2640,N_2637);
xor U2830 (N_2830,N_2609,N_2588);
and U2831 (N_2831,N_2634,N_2583);
nor U2832 (N_2832,N_2551,N_2630);
nor U2833 (N_2833,N_2639,N_2592);
or U2834 (N_2834,N_2699,N_2550);
nand U2835 (N_2835,N_2627,N_2595);
xor U2836 (N_2836,N_2669,N_2658);
xnor U2837 (N_2837,N_2652,N_2667);
xor U2838 (N_2838,N_2615,N_2666);
nor U2839 (N_2839,N_2690,N_2667);
or U2840 (N_2840,N_2647,N_2688);
nor U2841 (N_2841,N_2667,N_2698);
nand U2842 (N_2842,N_2564,N_2587);
nor U2843 (N_2843,N_2636,N_2627);
or U2844 (N_2844,N_2646,N_2571);
and U2845 (N_2845,N_2567,N_2555);
or U2846 (N_2846,N_2635,N_2634);
xor U2847 (N_2847,N_2669,N_2551);
and U2848 (N_2848,N_2623,N_2559);
or U2849 (N_2849,N_2698,N_2583);
xor U2850 (N_2850,N_2823,N_2714);
nor U2851 (N_2851,N_2799,N_2710);
and U2852 (N_2852,N_2773,N_2786);
nor U2853 (N_2853,N_2723,N_2752);
nand U2854 (N_2854,N_2754,N_2804);
nand U2855 (N_2855,N_2836,N_2758);
nand U2856 (N_2856,N_2701,N_2821);
nor U2857 (N_2857,N_2757,N_2835);
nand U2858 (N_2858,N_2777,N_2817);
or U2859 (N_2859,N_2741,N_2713);
and U2860 (N_2860,N_2812,N_2730);
and U2861 (N_2861,N_2783,N_2768);
or U2862 (N_2862,N_2785,N_2769);
or U2863 (N_2863,N_2706,N_2822);
or U2864 (N_2864,N_2803,N_2738);
xnor U2865 (N_2865,N_2829,N_2734);
nor U2866 (N_2866,N_2815,N_2819);
and U2867 (N_2867,N_2728,N_2778);
and U2868 (N_2868,N_2750,N_2797);
or U2869 (N_2869,N_2762,N_2816);
and U2870 (N_2870,N_2833,N_2740);
and U2871 (N_2871,N_2761,N_2747);
and U2872 (N_2872,N_2790,N_2736);
and U2873 (N_2873,N_2726,N_2831);
nor U2874 (N_2874,N_2788,N_2746);
or U2875 (N_2875,N_2841,N_2832);
xor U2876 (N_2876,N_2789,N_2813);
or U2877 (N_2877,N_2733,N_2782);
nand U2878 (N_2878,N_2707,N_2784);
xnor U2879 (N_2879,N_2765,N_2827);
nor U2880 (N_2880,N_2742,N_2840);
or U2881 (N_2881,N_2828,N_2712);
and U2882 (N_2882,N_2808,N_2807);
nand U2883 (N_2883,N_2842,N_2763);
nor U2884 (N_2884,N_2766,N_2729);
or U2885 (N_2885,N_2796,N_2764);
nor U2886 (N_2886,N_2805,N_2751);
nand U2887 (N_2887,N_2849,N_2774);
or U2888 (N_2888,N_2770,N_2826);
and U2889 (N_2889,N_2834,N_2837);
and U2890 (N_2890,N_2737,N_2787);
and U2891 (N_2891,N_2776,N_2715);
nor U2892 (N_2892,N_2839,N_2814);
or U2893 (N_2893,N_2755,N_2838);
xnor U2894 (N_2894,N_2846,N_2779);
and U2895 (N_2895,N_2753,N_2731);
xnor U2896 (N_2896,N_2711,N_2749);
or U2897 (N_2897,N_2727,N_2847);
xnor U2898 (N_2898,N_2775,N_2767);
xnor U2899 (N_2899,N_2781,N_2818);
nand U2900 (N_2900,N_2709,N_2801);
xnor U2901 (N_2901,N_2795,N_2809);
nor U2902 (N_2902,N_2825,N_2700);
and U2903 (N_2903,N_2845,N_2719);
nor U2904 (N_2904,N_2708,N_2759);
xnor U2905 (N_2905,N_2725,N_2844);
xor U2906 (N_2906,N_2793,N_2802);
nand U2907 (N_2907,N_2848,N_2745);
and U2908 (N_2908,N_2744,N_2748);
xor U2909 (N_2909,N_2792,N_2800);
nor U2910 (N_2910,N_2705,N_2716);
or U2911 (N_2911,N_2717,N_2743);
nand U2912 (N_2912,N_2772,N_2721);
nor U2913 (N_2913,N_2820,N_2810);
or U2914 (N_2914,N_2718,N_2702);
nor U2915 (N_2915,N_2735,N_2806);
or U2916 (N_2916,N_2703,N_2724);
and U2917 (N_2917,N_2811,N_2732);
xnor U2918 (N_2918,N_2739,N_2704);
nor U2919 (N_2919,N_2791,N_2756);
xor U2920 (N_2920,N_2722,N_2798);
and U2921 (N_2921,N_2830,N_2843);
nor U2922 (N_2922,N_2780,N_2760);
and U2923 (N_2923,N_2794,N_2771);
nand U2924 (N_2924,N_2824,N_2720);
xor U2925 (N_2925,N_2711,N_2810);
nand U2926 (N_2926,N_2752,N_2787);
nor U2927 (N_2927,N_2727,N_2750);
xor U2928 (N_2928,N_2751,N_2795);
and U2929 (N_2929,N_2773,N_2750);
nor U2930 (N_2930,N_2832,N_2822);
nand U2931 (N_2931,N_2707,N_2843);
nand U2932 (N_2932,N_2741,N_2722);
and U2933 (N_2933,N_2767,N_2834);
nand U2934 (N_2934,N_2803,N_2714);
or U2935 (N_2935,N_2840,N_2829);
xor U2936 (N_2936,N_2801,N_2796);
nor U2937 (N_2937,N_2817,N_2822);
and U2938 (N_2938,N_2846,N_2773);
and U2939 (N_2939,N_2712,N_2793);
xor U2940 (N_2940,N_2817,N_2782);
or U2941 (N_2941,N_2842,N_2802);
or U2942 (N_2942,N_2811,N_2770);
xnor U2943 (N_2943,N_2707,N_2778);
and U2944 (N_2944,N_2736,N_2766);
or U2945 (N_2945,N_2732,N_2781);
xor U2946 (N_2946,N_2724,N_2780);
xor U2947 (N_2947,N_2801,N_2805);
xnor U2948 (N_2948,N_2788,N_2781);
xnor U2949 (N_2949,N_2772,N_2820);
nand U2950 (N_2950,N_2824,N_2764);
and U2951 (N_2951,N_2843,N_2806);
and U2952 (N_2952,N_2846,N_2791);
nor U2953 (N_2953,N_2742,N_2827);
nand U2954 (N_2954,N_2833,N_2806);
and U2955 (N_2955,N_2803,N_2711);
and U2956 (N_2956,N_2785,N_2728);
or U2957 (N_2957,N_2710,N_2717);
nand U2958 (N_2958,N_2719,N_2712);
nand U2959 (N_2959,N_2761,N_2816);
nand U2960 (N_2960,N_2712,N_2762);
and U2961 (N_2961,N_2802,N_2815);
or U2962 (N_2962,N_2750,N_2841);
and U2963 (N_2963,N_2738,N_2726);
nand U2964 (N_2964,N_2808,N_2794);
nand U2965 (N_2965,N_2840,N_2846);
nand U2966 (N_2966,N_2705,N_2718);
or U2967 (N_2967,N_2759,N_2792);
or U2968 (N_2968,N_2742,N_2767);
xor U2969 (N_2969,N_2727,N_2818);
nand U2970 (N_2970,N_2703,N_2721);
xor U2971 (N_2971,N_2716,N_2797);
xor U2972 (N_2972,N_2720,N_2840);
or U2973 (N_2973,N_2799,N_2739);
or U2974 (N_2974,N_2728,N_2841);
or U2975 (N_2975,N_2741,N_2832);
or U2976 (N_2976,N_2747,N_2750);
nand U2977 (N_2977,N_2799,N_2749);
nor U2978 (N_2978,N_2834,N_2725);
nor U2979 (N_2979,N_2805,N_2800);
and U2980 (N_2980,N_2758,N_2732);
nor U2981 (N_2981,N_2809,N_2747);
or U2982 (N_2982,N_2700,N_2795);
nor U2983 (N_2983,N_2847,N_2787);
or U2984 (N_2984,N_2745,N_2775);
xor U2985 (N_2985,N_2816,N_2837);
nand U2986 (N_2986,N_2753,N_2778);
xnor U2987 (N_2987,N_2752,N_2762);
xor U2988 (N_2988,N_2717,N_2754);
and U2989 (N_2989,N_2822,N_2840);
nor U2990 (N_2990,N_2769,N_2760);
nor U2991 (N_2991,N_2772,N_2814);
nand U2992 (N_2992,N_2815,N_2781);
or U2993 (N_2993,N_2750,N_2811);
xor U2994 (N_2994,N_2773,N_2789);
and U2995 (N_2995,N_2717,N_2832);
nor U2996 (N_2996,N_2845,N_2732);
xnor U2997 (N_2997,N_2832,N_2768);
nor U2998 (N_2998,N_2799,N_2792);
nand U2999 (N_2999,N_2719,N_2702);
nand U3000 (N_3000,N_2955,N_2933);
nand U3001 (N_3001,N_2935,N_2989);
and U3002 (N_3002,N_2873,N_2992);
nor U3003 (N_3003,N_2894,N_2887);
or U3004 (N_3004,N_2975,N_2931);
nand U3005 (N_3005,N_2890,N_2857);
nor U3006 (N_3006,N_2860,N_2971);
nor U3007 (N_3007,N_2994,N_2932);
or U3008 (N_3008,N_2930,N_2905);
or U3009 (N_3009,N_2962,N_2987);
or U3010 (N_3010,N_2973,N_2944);
nor U3011 (N_3011,N_2946,N_2924);
nor U3012 (N_3012,N_2895,N_2900);
nand U3013 (N_3013,N_2912,N_2880);
nor U3014 (N_3014,N_2999,N_2988);
nor U3015 (N_3015,N_2974,N_2993);
and U3016 (N_3016,N_2953,N_2885);
nand U3017 (N_3017,N_2956,N_2983);
or U3018 (N_3018,N_2906,N_2864);
xnor U3019 (N_3019,N_2856,N_2915);
nand U3020 (N_3020,N_2898,N_2875);
or U3021 (N_3021,N_2911,N_2929);
nand U3022 (N_3022,N_2865,N_2928);
nand U3023 (N_3023,N_2985,N_2909);
xnor U3024 (N_3024,N_2982,N_2964);
nor U3025 (N_3025,N_2899,N_2939);
and U3026 (N_3026,N_2959,N_2984);
nor U3027 (N_3027,N_2901,N_2947);
or U3028 (N_3028,N_2893,N_2876);
and U3029 (N_3029,N_2986,N_2854);
nor U3030 (N_3030,N_2936,N_2995);
or U3031 (N_3031,N_2997,N_2920);
nor U3032 (N_3032,N_2957,N_2980);
and U3033 (N_3033,N_2850,N_2948);
and U3034 (N_3034,N_2918,N_2938);
or U3035 (N_3035,N_2967,N_2877);
nand U3036 (N_3036,N_2851,N_2870);
nor U3037 (N_3037,N_2937,N_2934);
xor U3038 (N_3038,N_2969,N_2950);
nor U3039 (N_3039,N_2863,N_2917);
xnor U3040 (N_3040,N_2892,N_2926);
nor U3041 (N_3041,N_2963,N_2852);
or U3042 (N_3042,N_2861,N_2889);
nor U3043 (N_3043,N_2965,N_2881);
nor U3044 (N_3044,N_2859,N_2978);
and U3045 (N_3045,N_2990,N_2869);
or U3046 (N_3046,N_2991,N_2927);
nor U3047 (N_3047,N_2884,N_2872);
nor U3048 (N_3048,N_2976,N_2897);
or U3049 (N_3049,N_2960,N_2923);
xor U3050 (N_3050,N_2968,N_2882);
and U3051 (N_3051,N_2868,N_2855);
nor U3052 (N_3052,N_2943,N_2903);
nand U3053 (N_3053,N_2961,N_2871);
nand U3054 (N_3054,N_2874,N_2858);
nand U3055 (N_3055,N_2879,N_2891);
nor U3056 (N_3056,N_2981,N_2966);
nand U3057 (N_3057,N_2910,N_2945);
or U3058 (N_3058,N_2913,N_2896);
and U3059 (N_3059,N_2862,N_2904);
nor U3060 (N_3060,N_2941,N_2853);
xnor U3061 (N_3061,N_2952,N_2907);
or U3062 (N_3062,N_2922,N_2949);
nor U3063 (N_3063,N_2867,N_2886);
and U3064 (N_3064,N_2942,N_2914);
nor U3065 (N_3065,N_2921,N_2972);
xor U3066 (N_3066,N_2954,N_2977);
nand U3067 (N_3067,N_2925,N_2908);
xnor U3068 (N_3068,N_2979,N_2902);
or U3069 (N_3069,N_2998,N_2916);
or U3070 (N_3070,N_2919,N_2996);
nor U3071 (N_3071,N_2866,N_2883);
xor U3072 (N_3072,N_2958,N_2878);
or U3073 (N_3073,N_2940,N_2970);
xor U3074 (N_3074,N_2951,N_2888);
and U3075 (N_3075,N_2965,N_2905);
and U3076 (N_3076,N_2985,N_2893);
nor U3077 (N_3077,N_2964,N_2973);
or U3078 (N_3078,N_2908,N_2983);
or U3079 (N_3079,N_2906,N_2918);
xor U3080 (N_3080,N_2971,N_2937);
and U3081 (N_3081,N_2904,N_2922);
and U3082 (N_3082,N_2941,N_2869);
nand U3083 (N_3083,N_2911,N_2879);
nor U3084 (N_3084,N_2981,N_2878);
or U3085 (N_3085,N_2931,N_2985);
and U3086 (N_3086,N_2914,N_2972);
nand U3087 (N_3087,N_2881,N_2946);
and U3088 (N_3088,N_2969,N_2988);
or U3089 (N_3089,N_2866,N_2861);
nand U3090 (N_3090,N_2940,N_2993);
or U3091 (N_3091,N_2890,N_2881);
nor U3092 (N_3092,N_2917,N_2971);
and U3093 (N_3093,N_2874,N_2887);
and U3094 (N_3094,N_2937,N_2920);
and U3095 (N_3095,N_2851,N_2957);
or U3096 (N_3096,N_2915,N_2876);
xor U3097 (N_3097,N_2960,N_2871);
xor U3098 (N_3098,N_2917,N_2924);
and U3099 (N_3099,N_2909,N_2926);
or U3100 (N_3100,N_2948,N_2946);
and U3101 (N_3101,N_2936,N_2899);
nand U3102 (N_3102,N_2984,N_2901);
nor U3103 (N_3103,N_2986,N_2906);
xor U3104 (N_3104,N_2859,N_2954);
nor U3105 (N_3105,N_2929,N_2957);
and U3106 (N_3106,N_2909,N_2973);
or U3107 (N_3107,N_2911,N_2891);
or U3108 (N_3108,N_2999,N_2876);
nand U3109 (N_3109,N_2934,N_2857);
and U3110 (N_3110,N_2998,N_2874);
xnor U3111 (N_3111,N_2922,N_2965);
nor U3112 (N_3112,N_2990,N_2961);
and U3113 (N_3113,N_2952,N_2923);
xnor U3114 (N_3114,N_2888,N_2860);
nor U3115 (N_3115,N_2889,N_2853);
nand U3116 (N_3116,N_2870,N_2977);
nor U3117 (N_3117,N_2925,N_2885);
xor U3118 (N_3118,N_2992,N_2943);
xnor U3119 (N_3119,N_2973,N_2915);
xnor U3120 (N_3120,N_2891,N_2983);
nor U3121 (N_3121,N_2962,N_2912);
and U3122 (N_3122,N_2891,N_2851);
or U3123 (N_3123,N_2882,N_2955);
nor U3124 (N_3124,N_2925,N_2894);
xnor U3125 (N_3125,N_2859,N_2914);
nand U3126 (N_3126,N_2928,N_2910);
or U3127 (N_3127,N_2922,N_2875);
nand U3128 (N_3128,N_2947,N_2995);
and U3129 (N_3129,N_2958,N_2868);
nor U3130 (N_3130,N_2905,N_2866);
nor U3131 (N_3131,N_2971,N_2923);
xor U3132 (N_3132,N_2906,N_2960);
or U3133 (N_3133,N_2850,N_2908);
and U3134 (N_3134,N_2925,N_2867);
and U3135 (N_3135,N_2936,N_2935);
nand U3136 (N_3136,N_2922,N_2856);
and U3137 (N_3137,N_2910,N_2987);
nor U3138 (N_3138,N_2879,N_2857);
nand U3139 (N_3139,N_2943,N_2969);
nand U3140 (N_3140,N_2948,N_2892);
and U3141 (N_3141,N_2851,N_2875);
and U3142 (N_3142,N_2867,N_2923);
nor U3143 (N_3143,N_2984,N_2875);
nand U3144 (N_3144,N_2868,N_2944);
or U3145 (N_3145,N_2944,N_2929);
or U3146 (N_3146,N_2888,N_2850);
or U3147 (N_3147,N_2905,N_2924);
nor U3148 (N_3148,N_2991,N_2907);
xnor U3149 (N_3149,N_2965,N_2880);
or U3150 (N_3150,N_3130,N_3033);
or U3151 (N_3151,N_3149,N_3097);
nand U3152 (N_3152,N_3069,N_3023);
nand U3153 (N_3153,N_3073,N_3012);
nor U3154 (N_3154,N_3013,N_3057);
and U3155 (N_3155,N_3040,N_3122);
nand U3156 (N_3156,N_3030,N_3045);
xnor U3157 (N_3157,N_3135,N_3031);
or U3158 (N_3158,N_3016,N_3140);
nand U3159 (N_3159,N_3141,N_3022);
nand U3160 (N_3160,N_3017,N_3129);
or U3161 (N_3161,N_3037,N_3029);
xor U3162 (N_3162,N_3078,N_3131);
and U3163 (N_3163,N_3065,N_3103);
or U3164 (N_3164,N_3049,N_3002);
nand U3165 (N_3165,N_3063,N_3100);
nor U3166 (N_3166,N_3068,N_3041);
xnor U3167 (N_3167,N_3095,N_3005);
or U3168 (N_3168,N_3145,N_3123);
and U3169 (N_3169,N_3136,N_3044);
nand U3170 (N_3170,N_3094,N_3118);
and U3171 (N_3171,N_3116,N_3021);
nand U3172 (N_3172,N_3074,N_3142);
nor U3173 (N_3173,N_3056,N_3096);
nand U3174 (N_3174,N_3008,N_3088);
and U3175 (N_3175,N_3083,N_3082);
xor U3176 (N_3176,N_3015,N_3062);
nand U3177 (N_3177,N_3092,N_3014);
xor U3178 (N_3178,N_3038,N_3020);
nand U3179 (N_3179,N_3090,N_3007);
or U3180 (N_3180,N_3019,N_3146);
xnor U3181 (N_3181,N_3053,N_3138);
nor U3182 (N_3182,N_3132,N_3035);
and U3183 (N_3183,N_3050,N_3047);
xnor U3184 (N_3184,N_3107,N_3024);
nand U3185 (N_3185,N_3051,N_3032);
nor U3186 (N_3186,N_3076,N_3115);
xnor U3187 (N_3187,N_3060,N_3072);
xnor U3188 (N_3188,N_3148,N_3093);
and U3189 (N_3189,N_3067,N_3119);
and U3190 (N_3190,N_3025,N_3085);
nor U3191 (N_3191,N_3101,N_3006);
xor U3192 (N_3192,N_3059,N_3113);
and U3193 (N_3193,N_3018,N_3048);
or U3194 (N_3194,N_3043,N_3064);
nor U3195 (N_3195,N_3003,N_3147);
and U3196 (N_3196,N_3027,N_3066);
nand U3197 (N_3197,N_3106,N_3098);
nor U3198 (N_3198,N_3117,N_3128);
and U3199 (N_3199,N_3054,N_3061);
xnor U3200 (N_3200,N_3009,N_3111);
or U3201 (N_3201,N_3026,N_3144);
nor U3202 (N_3202,N_3124,N_3086);
nand U3203 (N_3203,N_3114,N_3070);
xor U3204 (N_3204,N_3084,N_3089);
nor U3205 (N_3205,N_3001,N_3112);
nand U3206 (N_3206,N_3105,N_3102);
or U3207 (N_3207,N_3104,N_3055);
xnor U3208 (N_3208,N_3139,N_3099);
nand U3209 (N_3209,N_3046,N_3036);
xnor U3210 (N_3210,N_3110,N_3081);
nor U3211 (N_3211,N_3087,N_3127);
nor U3212 (N_3212,N_3108,N_3039);
xor U3213 (N_3213,N_3133,N_3010);
xnor U3214 (N_3214,N_3126,N_3077);
or U3215 (N_3215,N_3071,N_3004);
xnor U3216 (N_3216,N_3120,N_3079);
nor U3217 (N_3217,N_3121,N_3125);
xnor U3218 (N_3218,N_3137,N_3143);
xor U3219 (N_3219,N_3000,N_3091);
nand U3220 (N_3220,N_3052,N_3109);
or U3221 (N_3221,N_3028,N_3011);
nand U3222 (N_3222,N_3075,N_3134);
nand U3223 (N_3223,N_3034,N_3042);
nor U3224 (N_3224,N_3058,N_3080);
nor U3225 (N_3225,N_3094,N_3020);
nand U3226 (N_3226,N_3104,N_3119);
nor U3227 (N_3227,N_3067,N_3003);
and U3228 (N_3228,N_3125,N_3128);
nor U3229 (N_3229,N_3022,N_3074);
nor U3230 (N_3230,N_3007,N_3126);
and U3231 (N_3231,N_3020,N_3085);
nand U3232 (N_3232,N_3044,N_3037);
nor U3233 (N_3233,N_3107,N_3021);
nand U3234 (N_3234,N_3046,N_3103);
nand U3235 (N_3235,N_3124,N_3012);
and U3236 (N_3236,N_3087,N_3077);
nand U3237 (N_3237,N_3054,N_3029);
xor U3238 (N_3238,N_3064,N_3084);
nand U3239 (N_3239,N_3126,N_3048);
nand U3240 (N_3240,N_3109,N_3016);
xor U3241 (N_3241,N_3147,N_3148);
nand U3242 (N_3242,N_3049,N_3147);
and U3243 (N_3243,N_3110,N_3104);
xnor U3244 (N_3244,N_3057,N_3133);
nor U3245 (N_3245,N_3120,N_3107);
or U3246 (N_3246,N_3052,N_3006);
or U3247 (N_3247,N_3125,N_3079);
nor U3248 (N_3248,N_3005,N_3069);
nor U3249 (N_3249,N_3036,N_3092);
or U3250 (N_3250,N_3092,N_3033);
nor U3251 (N_3251,N_3115,N_3144);
nor U3252 (N_3252,N_3046,N_3000);
nand U3253 (N_3253,N_3103,N_3074);
and U3254 (N_3254,N_3121,N_3070);
nand U3255 (N_3255,N_3089,N_3100);
or U3256 (N_3256,N_3110,N_3098);
or U3257 (N_3257,N_3015,N_3134);
nand U3258 (N_3258,N_3115,N_3100);
nor U3259 (N_3259,N_3102,N_3114);
and U3260 (N_3260,N_3132,N_3062);
nor U3261 (N_3261,N_3046,N_3049);
xnor U3262 (N_3262,N_3081,N_3134);
and U3263 (N_3263,N_3012,N_3103);
xor U3264 (N_3264,N_3119,N_3124);
nand U3265 (N_3265,N_3105,N_3087);
xnor U3266 (N_3266,N_3135,N_3028);
xnor U3267 (N_3267,N_3141,N_3129);
xor U3268 (N_3268,N_3070,N_3012);
nor U3269 (N_3269,N_3033,N_3036);
nand U3270 (N_3270,N_3009,N_3031);
or U3271 (N_3271,N_3043,N_3109);
or U3272 (N_3272,N_3134,N_3110);
or U3273 (N_3273,N_3136,N_3046);
or U3274 (N_3274,N_3063,N_3012);
nand U3275 (N_3275,N_3064,N_3018);
or U3276 (N_3276,N_3066,N_3141);
nand U3277 (N_3277,N_3132,N_3079);
and U3278 (N_3278,N_3103,N_3097);
nand U3279 (N_3279,N_3108,N_3139);
nand U3280 (N_3280,N_3121,N_3062);
and U3281 (N_3281,N_3119,N_3036);
and U3282 (N_3282,N_3082,N_3025);
or U3283 (N_3283,N_3079,N_3003);
and U3284 (N_3284,N_3052,N_3092);
nand U3285 (N_3285,N_3114,N_3050);
or U3286 (N_3286,N_3009,N_3134);
and U3287 (N_3287,N_3149,N_3024);
nor U3288 (N_3288,N_3013,N_3079);
nor U3289 (N_3289,N_3025,N_3141);
nor U3290 (N_3290,N_3107,N_3063);
xnor U3291 (N_3291,N_3118,N_3129);
xnor U3292 (N_3292,N_3076,N_3016);
or U3293 (N_3293,N_3098,N_3001);
or U3294 (N_3294,N_3082,N_3031);
nor U3295 (N_3295,N_3055,N_3029);
and U3296 (N_3296,N_3038,N_3032);
nor U3297 (N_3297,N_3000,N_3149);
xnor U3298 (N_3298,N_3114,N_3033);
or U3299 (N_3299,N_3035,N_3140);
nor U3300 (N_3300,N_3235,N_3278);
nor U3301 (N_3301,N_3284,N_3260);
xor U3302 (N_3302,N_3220,N_3207);
or U3303 (N_3303,N_3189,N_3266);
or U3304 (N_3304,N_3184,N_3162);
xor U3305 (N_3305,N_3229,N_3177);
nand U3306 (N_3306,N_3274,N_3298);
or U3307 (N_3307,N_3192,N_3227);
nor U3308 (N_3308,N_3290,N_3233);
xnor U3309 (N_3309,N_3152,N_3167);
or U3310 (N_3310,N_3232,N_3283);
xnor U3311 (N_3311,N_3244,N_3238);
or U3312 (N_3312,N_3247,N_3156);
nand U3313 (N_3313,N_3161,N_3191);
and U3314 (N_3314,N_3277,N_3288);
xor U3315 (N_3315,N_3195,N_3246);
and U3316 (N_3316,N_3250,N_3296);
xnor U3317 (N_3317,N_3263,N_3292);
or U3318 (N_3318,N_3255,N_3293);
and U3319 (N_3319,N_3159,N_3231);
nor U3320 (N_3320,N_3219,N_3271);
nand U3321 (N_3321,N_3200,N_3190);
xor U3322 (N_3322,N_3257,N_3234);
nor U3323 (N_3323,N_3272,N_3160);
nor U3324 (N_3324,N_3225,N_3222);
or U3325 (N_3325,N_3254,N_3201);
and U3326 (N_3326,N_3249,N_3258);
and U3327 (N_3327,N_3181,N_3275);
and U3328 (N_3328,N_3215,N_3178);
or U3329 (N_3329,N_3248,N_3173);
or U3330 (N_3330,N_3281,N_3228);
nor U3331 (N_3331,N_3256,N_3268);
or U3332 (N_3332,N_3174,N_3157);
xor U3333 (N_3333,N_3253,N_3150);
nor U3334 (N_3334,N_3203,N_3209);
nor U3335 (N_3335,N_3210,N_3230);
nand U3336 (N_3336,N_3205,N_3179);
xnor U3337 (N_3337,N_3226,N_3170);
or U3338 (N_3338,N_3198,N_3270);
xnor U3339 (N_3339,N_3180,N_3297);
or U3340 (N_3340,N_3267,N_3251);
or U3341 (N_3341,N_3237,N_3155);
and U3342 (N_3342,N_3199,N_3193);
and U3343 (N_3343,N_3213,N_3224);
and U3344 (N_3344,N_3216,N_3212);
nand U3345 (N_3345,N_3211,N_3289);
and U3346 (N_3346,N_3295,N_3279);
xnor U3347 (N_3347,N_3282,N_3204);
nand U3348 (N_3348,N_3208,N_3239);
xor U3349 (N_3349,N_3166,N_3245);
or U3350 (N_3350,N_3176,N_3165);
xor U3351 (N_3351,N_3168,N_3287);
xor U3352 (N_3352,N_3171,N_3158);
or U3353 (N_3353,N_3186,N_3196);
nor U3354 (N_3354,N_3291,N_3280);
and U3355 (N_3355,N_3241,N_3299);
or U3356 (N_3356,N_3172,N_3259);
nand U3357 (N_3357,N_3236,N_3182);
xnor U3358 (N_3358,N_3197,N_3214);
xnor U3359 (N_3359,N_3252,N_3151);
and U3360 (N_3360,N_3242,N_3285);
nor U3361 (N_3361,N_3240,N_3183);
nand U3362 (N_3362,N_3217,N_3218);
nor U3363 (N_3363,N_3273,N_3185);
or U3364 (N_3364,N_3276,N_3269);
and U3365 (N_3365,N_3261,N_3265);
nand U3366 (N_3366,N_3194,N_3188);
nor U3367 (N_3367,N_3164,N_3262);
nand U3368 (N_3368,N_3163,N_3175);
xor U3369 (N_3369,N_3223,N_3187);
xnor U3370 (N_3370,N_3286,N_3294);
and U3371 (N_3371,N_3202,N_3153);
or U3372 (N_3372,N_3243,N_3264);
or U3373 (N_3373,N_3221,N_3206);
or U3374 (N_3374,N_3154,N_3169);
xor U3375 (N_3375,N_3291,N_3160);
xnor U3376 (N_3376,N_3210,N_3224);
and U3377 (N_3377,N_3163,N_3260);
nor U3378 (N_3378,N_3260,N_3162);
nor U3379 (N_3379,N_3296,N_3264);
or U3380 (N_3380,N_3162,N_3263);
nor U3381 (N_3381,N_3173,N_3261);
nand U3382 (N_3382,N_3203,N_3287);
nand U3383 (N_3383,N_3268,N_3226);
xor U3384 (N_3384,N_3224,N_3179);
nor U3385 (N_3385,N_3251,N_3277);
and U3386 (N_3386,N_3222,N_3293);
nor U3387 (N_3387,N_3232,N_3208);
nand U3388 (N_3388,N_3245,N_3298);
and U3389 (N_3389,N_3186,N_3218);
nor U3390 (N_3390,N_3180,N_3161);
and U3391 (N_3391,N_3180,N_3230);
nor U3392 (N_3392,N_3179,N_3167);
nor U3393 (N_3393,N_3212,N_3184);
or U3394 (N_3394,N_3297,N_3205);
nor U3395 (N_3395,N_3158,N_3214);
xor U3396 (N_3396,N_3171,N_3240);
xnor U3397 (N_3397,N_3290,N_3225);
nand U3398 (N_3398,N_3293,N_3153);
xor U3399 (N_3399,N_3256,N_3197);
and U3400 (N_3400,N_3150,N_3187);
nor U3401 (N_3401,N_3274,N_3205);
and U3402 (N_3402,N_3269,N_3253);
nor U3403 (N_3403,N_3217,N_3213);
xnor U3404 (N_3404,N_3289,N_3165);
nand U3405 (N_3405,N_3207,N_3176);
or U3406 (N_3406,N_3205,N_3166);
and U3407 (N_3407,N_3200,N_3274);
or U3408 (N_3408,N_3165,N_3209);
xnor U3409 (N_3409,N_3162,N_3256);
or U3410 (N_3410,N_3230,N_3273);
nor U3411 (N_3411,N_3233,N_3219);
xor U3412 (N_3412,N_3231,N_3179);
nand U3413 (N_3413,N_3272,N_3291);
nor U3414 (N_3414,N_3235,N_3288);
or U3415 (N_3415,N_3246,N_3270);
and U3416 (N_3416,N_3279,N_3253);
xnor U3417 (N_3417,N_3277,N_3198);
xor U3418 (N_3418,N_3299,N_3291);
nand U3419 (N_3419,N_3227,N_3164);
and U3420 (N_3420,N_3287,N_3234);
nand U3421 (N_3421,N_3245,N_3274);
or U3422 (N_3422,N_3255,N_3179);
nor U3423 (N_3423,N_3223,N_3157);
and U3424 (N_3424,N_3182,N_3161);
nor U3425 (N_3425,N_3153,N_3225);
nand U3426 (N_3426,N_3163,N_3255);
nor U3427 (N_3427,N_3250,N_3178);
and U3428 (N_3428,N_3293,N_3263);
and U3429 (N_3429,N_3264,N_3270);
nor U3430 (N_3430,N_3164,N_3237);
nor U3431 (N_3431,N_3250,N_3210);
xor U3432 (N_3432,N_3235,N_3150);
and U3433 (N_3433,N_3204,N_3299);
nand U3434 (N_3434,N_3209,N_3184);
and U3435 (N_3435,N_3169,N_3268);
nand U3436 (N_3436,N_3295,N_3163);
nor U3437 (N_3437,N_3245,N_3189);
nor U3438 (N_3438,N_3277,N_3194);
and U3439 (N_3439,N_3209,N_3198);
nor U3440 (N_3440,N_3190,N_3167);
or U3441 (N_3441,N_3182,N_3252);
xor U3442 (N_3442,N_3179,N_3199);
and U3443 (N_3443,N_3239,N_3199);
nor U3444 (N_3444,N_3220,N_3268);
nor U3445 (N_3445,N_3278,N_3220);
nor U3446 (N_3446,N_3276,N_3185);
and U3447 (N_3447,N_3187,N_3181);
or U3448 (N_3448,N_3251,N_3289);
nor U3449 (N_3449,N_3242,N_3174);
or U3450 (N_3450,N_3415,N_3365);
or U3451 (N_3451,N_3342,N_3431);
or U3452 (N_3452,N_3407,N_3441);
nor U3453 (N_3453,N_3448,N_3438);
nor U3454 (N_3454,N_3339,N_3393);
nor U3455 (N_3455,N_3389,N_3440);
and U3456 (N_3456,N_3447,N_3306);
or U3457 (N_3457,N_3334,N_3400);
and U3458 (N_3458,N_3432,N_3316);
nand U3459 (N_3459,N_3344,N_3366);
nand U3460 (N_3460,N_3322,N_3378);
nand U3461 (N_3461,N_3370,N_3421);
xor U3462 (N_3462,N_3445,N_3330);
and U3463 (N_3463,N_3359,N_3398);
or U3464 (N_3464,N_3302,N_3315);
xnor U3465 (N_3465,N_3426,N_3435);
nor U3466 (N_3466,N_3368,N_3308);
nand U3467 (N_3467,N_3301,N_3351);
xnor U3468 (N_3468,N_3364,N_3312);
nor U3469 (N_3469,N_3347,N_3444);
nor U3470 (N_3470,N_3386,N_3382);
or U3471 (N_3471,N_3425,N_3323);
and U3472 (N_3472,N_3419,N_3317);
nor U3473 (N_3473,N_3420,N_3310);
or U3474 (N_3474,N_3380,N_3318);
nor U3475 (N_3475,N_3383,N_3385);
nor U3476 (N_3476,N_3362,N_3410);
xnor U3477 (N_3477,N_3436,N_3353);
nand U3478 (N_3478,N_3372,N_3417);
or U3479 (N_3479,N_3309,N_3409);
or U3480 (N_3480,N_3427,N_3331);
and U3481 (N_3481,N_3369,N_3337);
xor U3482 (N_3482,N_3329,N_3326);
nor U3483 (N_3483,N_3423,N_3402);
xnor U3484 (N_3484,N_3404,N_3406);
nand U3485 (N_3485,N_3416,N_3333);
or U3486 (N_3486,N_3336,N_3395);
nor U3487 (N_3487,N_3327,N_3300);
nand U3488 (N_3488,N_3422,N_3379);
nand U3489 (N_3489,N_3373,N_3341);
xnor U3490 (N_3490,N_3408,N_3411);
and U3491 (N_3491,N_3413,N_3412);
nor U3492 (N_3492,N_3350,N_3387);
nand U3493 (N_3493,N_3376,N_3443);
and U3494 (N_3494,N_3335,N_3303);
nor U3495 (N_3495,N_3401,N_3439);
nand U3496 (N_3496,N_3433,N_3442);
nor U3497 (N_3497,N_3345,N_3429);
nor U3498 (N_3498,N_3320,N_3394);
or U3499 (N_3499,N_3340,N_3360);
or U3500 (N_3500,N_3356,N_3346);
nand U3501 (N_3501,N_3313,N_3354);
or U3502 (N_3502,N_3338,N_3314);
and U3503 (N_3503,N_3374,N_3392);
xor U3504 (N_3504,N_3405,N_3397);
nand U3505 (N_3505,N_3352,N_3434);
xnor U3506 (N_3506,N_3377,N_3414);
nand U3507 (N_3507,N_3367,N_3399);
nand U3508 (N_3508,N_3446,N_3348);
xor U3509 (N_3509,N_3361,N_3403);
nor U3510 (N_3510,N_3449,N_3349);
and U3511 (N_3511,N_3325,N_3358);
nand U3512 (N_3512,N_3390,N_3428);
nor U3513 (N_3513,N_3391,N_3396);
and U3514 (N_3514,N_3304,N_3357);
nor U3515 (N_3515,N_3371,N_3321);
xnor U3516 (N_3516,N_3307,N_3305);
nand U3517 (N_3517,N_3388,N_3311);
xor U3518 (N_3518,N_3384,N_3355);
nand U3519 (N_3519,N_3343,N_3363);
nand U3520 (N_3520,N_3381,N_3324);
or U3521 (N_3521,N_3375,N_3332);
and U3522 (N_3522,N_3424,N_3430);
nor U3523 (N_3523,N_3319,N_3328);
nand U3524 (N_3524,N_3437,N_3418);
xnor U3525 (N_3525,N_3335,N_3361);
nor U3526 (N_3526,N_3378,N_3386);
nor U3527 (N_3527,N_3342,N_3369);
or U3528 (N_3528,N_3341,N_3420);
and U3529 (N_3529,N_3387,N_3332);
xnor U3530 (N_3530,N_3383,N_3334);
xor U3531 (N_3531,N_3374,N_3407);
and U3532 (N_3532,N_3398,N_3363);
nand U3533 (N_3533,N_3394,N_3339);
or U3534 (N_3534,N_3438,N_3392);
and U3535 (N_3535,N_3387,N_3365);
nand U3536 (N_3536,N_3367,N_3354);
and U3537 (N_3537,N_3410,N_3395);
or U3538 (N_3538,N_3300,N_3330);
and U3539 (N_3539,N_3310,N_3326);
and U3540 (N_3540,N_3425,N_3443);
xor U3541 (N_3541,N_3432,N_3357);
and U3542 (N_3542,N_3422,N_3366);
nor U3543 (N_3543,N_3375,N_3358);
nand U3544 (N_3544,N_3326,N_3448);
nor U3545 (N_3545,N_3354,N_3324);
nor U3546 (N_3546,N_3432,N_3360);
or U3547 (N_3547,N_3330,N_3449);
nor U3548 (N_3548,N_3310,N_3306);
nand U3549 (N_3549,N_3416,N_3414);
and U3550 (N_3550,N_3448,N_3316);
nor U3551 (N_3551,N_3394,N_3402);
or U3552 (N_3552,N_3388,N_3310);
nor U3553 (N_3553,N_3316,N_3320);
or U3554 (N_3554,N_3447,N_3319);
or U3555 (N_3555,N_3351,N_3375);
nand U3556 (N_3556,N_3424,N_3425);
xor U3557 (N_3557,N_3419,N_3359);
and U3558 (N_3558,N_3401,N_3312);
xor U3559 (N_3559,N_3367,N_3391);
or U3560 (N_3560,N_3403,N_3316);
nor U3561 (N_3561,N_3349,N_3324);
xor U3562 (N_3562,N_3449,N_3412);
or U3563 (N_3563,N_3399,N_3427);
and U3564 (N_3564,N_3373,N_3413);
nor U3565 (N_3565,N_3350,N_3420);
and U3566 (N_3566,N_3347,N_3301);
and U3567 (N_3567,N_3382,N_3427);
nand U3568 (N_3568,N_3332,N_3392);
nor U3569 (N_3569,N_3420,N_3349);
and U3570 (N_3570,N_3358,N_3405);
nor U3571 (N_3571,N_3395,N_3390);
nand U3572 (N_3572,N_3381,N_3394);
or U3573 (N_3573,N_3440,N_3419);
xor U3574 (N_3574,N_3360,N_3377);
nand U3575 (N_3575,N_3412,N_3372);
nor U3576 (N_3576,N_3344,N_3318);
and U3577 (N_3577,N_3324,N_3448);
or U3578 (N_3578,N_3330,N_3406);
xor U3579 (N_3579,N_3420,N_3362);
and U3580 (N_3580,N_3323,N_3438);
or U3581 (N_3581,N_3394,N_3414);
nor U3582 (N_3582,N_3380,N_3376);
and U3583 (N_3583,N_3383,N_3390);
xnor U3584 (N_3584,N_3384,N_3423);
nand U3585 (N_3585,N_3408,N_3412);
nand U3586 (N_3586,N_3374,N_3449);
nor U3587 (N_3587,N_3346,N_3399);
nor U3588 (N_3588,N_3360,N_3428);
and U3589 (N_3589,N_3385,N_3362);
or U3590 (N_3590,N_3441,N_3375);
and U3591 (N_3591,N_3407,N_3373);
xnor U3592 (N_3592,N_3315,N_3441);
and U3593 (N_3593,N_3428,N_3351);
or U3594 (N_3594,N_3397,N_3431);
xnor U3595 (N_3595,N_3435,N_3351);
or U3596 (N_3596,N_3435,N_3374);
nor U3597 (N_3597,N_3432,N_3386);
xor U3598 (N_3598,N_3315,N_3387);
nor U3599 (N_3599,N_3311,N_3423);
or U3600 (N_3600,N_3450,N_3491);
xnor U3601 (N_3601,N_3502,N_3527);
and U3602 (N_3602,N_3496,N_3472);
or U3603 (N_3603,N_3563,N_3560);
or U3604 (N_3604,N_3546,N_3485);
or U3605 (N_3605,N_3564,N_3545);
and U3606 (N_3606,N_3469,N_3483);
or U3607 (N_3607,N_3575,N_3598);
nor U3608 (N_3608,N_3479,N_3590);
xnor U3609 (N_3609,N_3520,N_3473);
nor U3610 (N_3610,N_3519,N_3461);
xnor U3611 (N_3611,N_3552,N_3530);
nand U3612 (N_3612,N_3467,N_3513);
nor U3613 (N_3613,N_3522,N_3567);
and U3614 (N_3614,N_3556,N_3458);
or U3615 (N_3615,N_3588,N_3532);
and U3616 (N_3616,N_3529,N_3537);
or U3617 (N_3617,N_3501,N_3538);
or U3618 (N_3618,N_3511,N_3454);
nand U3619 (N_3619,N_3570,N_3559);
nand U3620 (N_3620,N_3523,N_3474);
or U3621 (N_3621,N_3490,N_3548);
and U3622 (N_3622,N_3536,N_3494);
nand U3623 (N_3623,N_3573,N_3587);
xnor U3624 (N_3624,N_3478,N_3549);
nor U3625 (N_3625,N_3586,N_3475);
xor U3626 (N_3626,N_3488,N_3593);
nand U3627 (N_3627,N_3463,N_3540);
and U3628 (N_3628,N_3480,N_3464);
nand U3629 (N_3629,N_3525,N_3508);
or U3630 (N_3630,N_3535,N_3551);
or U3631 (N_3631,N_3471,N_3460);
and U3632 (N_3632,N_3515,N_3509);
nor U3633 (N_3633,N_3539,N_3544);
nor U3634 (N_3634,N_3569,N_3452);
nand U3635 (N_3635,N_3476,N_3486);
nor U3636 (N_3636,N_3571,N_3470);
or U3637 (N_3637,N_3459,N_3468);
and U3638 (N_3638,N_3578,N_3503);
nor U3639 (N_3639,N_3568,N_3497);
xor U3640 (N_3640,N_3561,N_3574);
xor U3641 (N_3641,N_3500,N_3555);
or U3642 (N_3642,N_3498,N_3594);
and U3643 (N_3643,N_3592,N_3596);
xnor U3644 (N_3644,N_3582,N_3521);
nand U3645 (N_3645,N_3453,N_3581);
nand U3646 (N_3646,N_3576,N_3566);
and U3647 (N_3647,N_3465,N_3565);
or U3648 (N_3648,N_3585,N_3462);
and U3649 (N_3649,N_3451,N_3487);
and U3650 (N_3650,N_3583,N_3492);
xnor U3651 (N_3651,N_3495,N_3499);
or U3652 (N_3652,N_3526,N_3482);
and U3653 (N_3653,N_3455,N_3518);
nor U3654 (N_3654,N_3512,N_3557);
nor U3655 (N_3655,N_3493,N_3584);
and U3656 (N_3656,N_3504,N_3481);
or U3657 (N_3657,N_3517,N_3554);
or U3658 (N_3658,N_3542,N_3599);
xnor U3659 (N_3659,N_3595,N_3456);
or U3660 (N_3660,N_3572,N_3489);
xor U3661 (N_3661,N_3533,N_3550);
xnor U3662 (N_3662,N_3531,N_3516);
nor U3663 (N_3663,N_3597,N_3562);
or U3664 (N_3664,N_3510,N_3457);
nor U3665 (N_3665,N_3484,N_3534);
or U3666 (N_3666,N_3589,N_3558);
nor U3667 (N_3667,N_3466,N_3514);
and U3668 (N_3668,N_3477,N_3541);
and U3669 (N_3669,N_3507,N_3553);
nand U3670 (N_3670,N_3524,N_3591);
nor U3671 (N_3671,N_3506,N_3579);
or U3672 (N_3672,N_3580,N_3577);
and U3673 (N_3673,N_3543,N_3528);
nor U3674 (N_3674,N_3547,N_3505);
xor U3675 (N_3675,N_3493,N_3516);
nor U3676 (N_3676,N_3599,N_3463);
xnor U3677 (N_3677,N_3562,N_3586);
or U3678 (N_3678,N_3518,N_3461);
nand U3679 (N_3679,N_3551,N_3559);
nor U3680 (N_3680,N_3529,N_3491);
xor U3681 (N_3681,N_3568,N_3460);
and U3682 (N_3682,N_3549,N_3486);
nand U3683 (N_3683,N_3476,N_3558);
or U3684 (N_3684,N_3595,N_3599);
nor U3685 (N_3685,N_3575,N_3583);
xor U3686 (N_3686,N_3518,N_3598);
and U3687 (N_3687,N_3494,N_3595);
and U3688 (N_3688,N_3507,N_3514);
or U3689 (N_3689,N_3542,N_3521);
xnor U3690 (N_3690,N_3566,N_3568);
and U3691 (N_3691,N_3572,N_3573);
and U3692 (N_3692,N_3593,N_3565);
xnor U3693 (N_3693,N_3473,N_3532);
nand U3694 (N_3694,N_3584,N_3547);
and U3695 (N_3695,N_3479,N_3503);
nor U3696 (N_3696,N_3520,N_3478);
xor U3697 (N_3697,N_3555,N_3521);
or U3698 (N_3698,N_3451,N_3486);
nor U3699 (N_3699,N_3529,N_3484);
and U3700 (N_3700,N_3453,N_3537);
or U3701 (N_3701,N_3467,N_3528);
or U3702 (N_3702,N_3491,N_3516);
or U3703 (N_3703,N_3559,N_3558);
xor U3704 (N_3704,N_3499,N_3589);
nor U3705 (N_3705,N_3547,N_3503);
nand U3706 (N_3706,N_3574,N_3598);
and U3707 (N_3707,N_3481,N_3453);
and U3708 (N_3708,N_3484,N_3521);
and U3709 (N_3709,N_3498,N_3530);
nor U3710 (N_3710,N_3530,N_3464);
nor U3711 (N_3711,N_3577,N_3543);
xnor U3712 (N_3712,N_3512,N_3472);
or U3713 (N_3713,N_3507,N_3511);
xnor U3714 (N_3714,N_3563,N_3464);
nor U3715 (N_3715,N_3455,N_3509);
nor U3716 (N_3716,N_3496,N_3499);
nor U3717 (N_3717,N_3545,N_3494);
or U3718 (N_3718,N_3473,N_3476);
nor U3719 (N_3719,N_3497,N_3551);
nor U3720 (N_3720,N_3460,N_3582);
nor U3721 (N_3721,N_3569,N_3558);
and U3722 (N_3722,N_3539,N_3488);
or U3723 (N_3723,N_3545,N_3579);
xnor U3724 (N_3724,N_3507,N_3500);
xnor U3725 (N_3725,N_3477,N_3591);
nor U3726 (N_3726,N_3535,N_3523);
or U3727 (N_3727,N_3540,N_3596);
or U3728 (N_3728,N_3528,N_3511);
and U3729 (N_3729,N_3596,N_3508);
xnor U3730 (N_3730,N_3532,N_3512);
or U3731 (N_3731,N_3457,N_3592);
nand U3732 (N_3732,N_3458,N_3543);
nor U3733 (N_3733,N_3522,N_3491);
or U3734 (N_3734,N_3465,N_3535);
nand U3735 (N_3735,N_3507,N_3540);
or U3736 (N_3736,N_3568,N_3550);
and U3737 (N_3737,N_3459,N_3583);
and U3738 (N_3738,N_3542,N_3595);
and U3739 (N_3739,N_3539,N_3589);
and U3740 (N_3740,N_3540,N_3575);
nand U3741 (N_3741,N_3522,N_3529);
nor U3742 (N_3742,N_3554,N_3523);
nand U3743 (N_3743,N_3590,N_3526);
nand U3744 (N_3744,N_3528,N_3560);
and U3745 (N_3745,N_3524,N_3587);
nand U3746 (N_3746,N_3480,N_3476);
xor U3747 (N_3747,N_3500,N_3564);
or U3748 (N_3748,N_3503,N_3560);
or U3749 (N_3749,N_3550,N_3546);
or U3750 (N_3750,N_3725,N_3604);
nor U3751 (N_3751,N_3668,N_3615);
xnor U3752 (N_3752,N_3632,N_3648);
nand U3753 (N_3753,N_3706,N_3697);
xnor U3754 (N_3754,N_3740,N_3652);
and U3755 (N_3755,N_3721,N_3636);
and U3756 (N_3756,N_3677,N_3620);
xor U3757 (N_3757,N_3645,N_3613);
nor U3758 (N_3758,N_3689,N_3618);
nor U3759 (N_3759,N_3609,N_3670);
xor U3760 (N_3760,N_3621,N_3674);
xnor U3761 (N_3761,N_3650,N_3711);
nor U3762 (N_3762,N_3681,N_3707);
or U3763 (N_3763,N_3710,N_3699);
and U3764 (N_3764,N_3608,N_3747);
nor U3765 (N_3765,N_3684,N_3654);
and U3766 (N_3766,N_3732,N_3735);
or U3767 (N_3767,N_3729,N_3746);
xnor U3768 (N_3768,N_3666,N_3682);
nor U3769 (N_3769,N_3683,N_3686);
or U3770 (N_3770,N_3687,N_3653);
xor U3771 (N_3771,N_3641,N_3680);
nand U3772 (N_3772,N_3694,N_3742);
xor U3773 (N_3773,N_3665,N_3663);
nand U3774 (N_3774,N_3626,N_3701);
nand U3775 (N_3775,N_3638,N_3605);
xnor U3776 (N_3776,N_3690,N_3606);
nor U3777 (N_3777,N_3679,N_3667);
and U3778 (N_3778,N_3612,N_3637);
nor U3779 (N_3779,N_3669,N_3722);
xor U3780 (N_3780,N_3745,N_3704);
nand U3781 (N_3781,N_3716,N_3622);
or U3782 (N_3782,N_3713,N_3741);
nand U3783 (N_3783,N_3610,N_3619);
or U3784 (N_3784,N_3696,N_3727);
nand U3785 (N_3785,N_3705,N_3734);
or U3786 (N_3786,N_3625,N_3691);
xor U3787 (N_3787,N_3749,N_3676);
nor U3788 (N_3788,N_3603,N_3644);
and U3789 (N_3789,N_3714,N_3744);
xnor U3790 (N_3790,N_3700,N_3703);
or U3791 (N_3791,N_3649,N_3731);
or U3792 (N_3792,N_3717,N_3600);
and U3793 (N_3793,N_3712,N_3658);
and U3794 (N_3794,N_3642,N_3631);
nand U3795 (N_3795,N_3662,N_3630);
and U3796 (N_3796,N_3624,N_3623);
nor U3797 (N_3797,N_3651,N_3616);
xnor U3798 (N_3798,N_3656,N_3660);
nor U3799 (N_3799,N_3692,N_3673);
xnor U3800 (N_3800,N_3672,N_3633);
nor U3801 (N_3801,N_3702,N_3678);
xor U3802 (N_3802,N_3743,N_3635);
and U3803 (N_3803,N_3655,N_3661);
nand U3804 (N_3804,N_3675,N_3646);
and U3805 (N_3805,N_3634,N_3693);
nor U3806 (N_3806,N_3739,N_3733);
nand U3807 (N_3807,N_3723,N_3728);
nand U3808 (N_3808,N_3708,N_3659);
xor U3809 (N_3809,N_3628,N_3685);
or U3810 (N_3810,N_3726,N_3688);
nand U3811 (N_3811,N_3720,N_3709);
or U3812 (N_3812,N_3602,N_3601);
and U3813 (N_3813,N_3736,N_3614);
nand U3814 (N_3814,N_3718,N_3695);
and U3815 (N_3815,N_3738,N_3748);
and U3816 (N_3816,N_3611,N_3640);
xor U3817 (N_3817,N_3627,N_3719);
xnor U3818 (N_3818,N_3715,N_3647);
xnor U3819 (N_3819,N_3639,N_3664);
nor U3820 (N_3820,N_3643,N_3737);
nand U3821 (N_3821,N_3724,N_3698);
and U3822 (N_3822,N_3607,N_3629);
nand U3823 (N_3823,N_3671,N_3657);
or U3824 (N_3824,N_3730,N_3617);
nor U3825 (N_3825,N_3605,N_3690);
or U3826 (N_3826,N_3744,N_3692);
xor U3827 (N_3827,N_3745,N_3743);
nand U3828 (N_3828,N_3714,N_3718);
and U3829 (N_3829,N_3608,N_3632);
nand U3830 (N_3830,N_3746,N_3682);
nand U3831 (N_3831,N_3725,N_3693);
or U3832 (N_3832,N_3657,N_3686);
and U3833 (N_3833,N_3646,N_3667);
nor U3834 (N_3834,N_3740,N_3730);
nand U3835 (N_3835,N_3613,N_3632);
or U3836 (N_3836,N_3749,N_3600);
nor U3837 (N_3837,N_3648,N_3643);
or U3838 (N_3838,N_3643,N_3728);
or U3839 (N_3839,N_3729,N_3624);
and U3840 (N_3840,N_3703,N_3602);
nor U3841 (N_3841,N_3669,N_3745);
nor U3842 (N_3842,N_3740,N_3627);
and U3843 (N_3843,N_3664,N_3681);
or U3844 (N_3844,N_3602,N_3659);
xor U3845 (N_3845,N_3628,N_3606);
or U3846 (N_3846,N_3659,N_3679);
xor U3847 (N_3847,N_3684,N_3602);
nand U3848 (N_3848,N_3640,N_3711);
nand U3849 (N_3849,N_3746,N_3657);
or U3850 (N_3850,N_3701,N_3646);
and U3851 (N_3851,N_3721,N_3627);
xnor U3852 (N_3852,N_3607,N_3612);
xor U3853 (N_3853,N_3727,N_3707);
nand U3854 (N_3854,N_3624,N_3617);
nor U3855 (N_3855,N_3687,N_3684);
nand U3856 (N_3856,N_3621,N_3652);
nor U3857 (N_3857,N_3717,N_3724);
and U3858 (N_3858,N_3706,N_3718);
and U3859 (N_3859,N_3635,N_3645);
and U3860 (N_3860,N_3658,N_3688);
nand U3861 (N_3861,N_3655,N_3701);
nor U3862 (N_3862,N_3684,N_3743);
nor U3863 (N_3863,N_3732,N_3743);
xnor U3864 (N_3864,N_3650,N_3730);
or U3865 (N_3865,N_3612,N_3736);
nor U3866 (N_3866,N_3696,N_3738);
nor U3867 (N_3867,N_3639,N_3621);
or U3868 (N_3868,N_3720,N_3723);
and U3869 (N_3869,N_3739,N_3629);
or U3870 (N_3870,N_3717,N_3623);
and U3871 (N_3871,N_3710,N_3647);
or U3872 (N_3872,N_3728,N_3677);
nand U3873 (N_3873,N_3667,N_3685);
nor U3874 (N_3874,N_3726,N_3639);
xnor U3875 (N_3875,N_3647,N_3702);
nand U3876 (N_3876,N_3662,N_3608);
nand U3877 (N_3877,N_3682,N_3693);
or U3878 (N_3878,N_3747,N_3685);
and U3879 (N_3879,N_3706,N_3629);
xnor U3880 (N_3880,N_3650,N_3637);
nand U3881 (N_3881,N_3736,N_3683);
and U3882 (N_3882,N_3673,N_3747);
or U3883 (N_3883,N_3724,N_3718);
and U3884 (N_3884,N_3700,N_3645);
nand U3885 (N_3885,N_3656,N_3722);
and U3886 (N_3886,N_3667,N_3630);
nor U3887 (N_3887,N_3735,N_3628);
or U3888 (N_3888,N_3707,N_3729);
xnor U3889 (N_3889,N_3649,N_3642);
nor U3890 (N_3890,N_3612,N_3651);
xor U3891 (N_3891,N_3662,N_3612);
nor U3892 (N_3892,N_3673,N_3733);
and U3893 (N_3893,N_3747,N_3655);
and U3894 (N_3894,N_3748,N_3660);
nand U3895 (N_3895,N_3730,N_3601);
xnor U3896 (N_3896,N_3665,N_3697);
xor U3897 (N_3897,N_3722,N_3725);
nand U3898 (N_3898,N_3606,N_3688);
and U3899 (N_3899,N_3709,N_3692);
nand U3900 (N_3900,N_3856,N_3774);
or U3901 (N_3901,N_3870,N_3886);
or U3902 (N_3902,N_3849,N_3865);
nand U3903 (N_3903,N_3755,N_3759);
nand U3904 (N_3904,N_3791,N_3787);
and U3905 (N_3905,N_3864,N_3779);
xnor U3906 (N_3906,N_3764,N_3862);
nor U3907 (N_3907,N_3883,N_3826);
nand U3908 (N_3908,N_3860,N_3793);
nand U3909 (N_3909,N_3812,N_3832);
or U3910 (N_3910,N_3808,N_3775);
nand U3911 (N_3911,N_3873,N_3859);
xnor U3912 (N_3912,N_3877,N_3843);
nand U3913 (N_3913,N_3811,N_3846);
or U3914 (N_3914,N_3762,N_3879);
and U3915 (N_3915,N_3894,N_3790);
or U3916 (N_3916,N_3829,N_3786);
xor U3917 (N_3917,N_3842,N_3890);
xor U3918 (N_3918,N_3854,N_3785);
xnor U3919 (N_3919,N_3835,N_3752);
or U3920 (N_3920,N_3821,N_3828);
nand U3921 (N_3921,N_3853,N_3781);
xnor U3922 (N_3922,N_3767,N_3803);
and U3923 (N_3923,N_3769,N_3796);
and U3924 (N_3924,N_3848,N_3872);
nand U3925 (N_3925,N_3758,N_3874);
or U3926 (N_3926,N_3822,N_3867);
or U3927 (N_3927,N_3809,N_3772);
nor U3928 (N_3928,N_3795,N_3851);
nor U3929 (N_3929,N_3757,N_3827);
nor U3930 (N_3930,N_3878,N_3751);
xnor U3931 (N_3931,N_3761,N_3852);
xor U3932 (N_3932,N_3783,N_3899);
and U3933 (N_3933,N_3869,N_3778);
xnor U3934 (N_3934,N_3861,N_3776);
xnor U3935 (N_3935,N_3845,N_3897);
xnor U3936 (N_3936,N_3750,N_3830);
or U3937 (N_3937,N_3804,N_3805);
and U3938 (N_3938,N_3875,N_3792);
nand U3939 (N_3939,N_3800,N_3798);
and U3940 (N_3940,N_3847,N_3754);
and U3941 (N_3941,N_3885,N_3893);
nand U3942 (N_3942,N_3797,N_3815);
nor U3943 (N_3943,N_3763,N_3844);
xnor U3944 (N_3944,N_3802,N_3756);
xor U3945 (N_3945,N_3863,N_3892);
or U3946 (N_3946,N_3810,N_3770);
nor U3947 (N_3947,N_3784,N_3868);
xor U3948 (N_3948,N_3888,N_3896);
xor U3949 (N_3949,N_3876,N_3880);
or U3950 (N_3950,N_3816,N_3801);
nor U3951 (N_3951,N_3833,N_3858);
nor U3952 (N_3952,N_3855,N_3794);
and U3953 (N_3953,N_3766,N_3838);
or U3954 (N_3954,N_3773,N_3825);
nand U3955 (N_3955,N_3771,N_3889);
xnor U3956 (N_3956,N_3850,N_3820);
nor U3957 (N_3957,N_3891,N_3768);
xor U3958 (N_3958,N_3807,N_3871);
nand U3959 (N_3959,N_3857,N_3814);
nor U3960 (N_3960,N_3765,N_3834);
xor U3961 (N_3961,N_3882,N_3823);
xnor U3962 (N_3962,N_3887,N_3898);
and U3963 (N_3963,N_3806,N_3895);
and U3964 (N_3964,N_3777,N_3837);
xnor U3965 (N_3965,N_3881,N_3841);
and U3966 (N_3966,N_3818,N_3866);
nand U3967 (N_3967,N_3788,N_3760);
nand U3968 (N_3968,N_3884,N_3780);
and U3969 (N_3969,N_3839,N_3813);
nor U3970 (N_3970,N_3819,N_3831);
nor U3971 (N_3971,N_3753,N_3817);
or U3972 (N_3972,N_3824,N_3782);
nand U3973 (N_3973,N_3840,N_3789);
or U3974 (N_3974,N_3836,N_3799);
xnor U3975 (N_3975,N_3881,N_3861);
or U3976 (N_3976,N_3886,N_3812);
or U3977 (N_3977,N_3760,N_3810);
xor U3978 (N_3978,N_3890,N_3790);
or U3979 (N_3979,N_3810,N_3855);
or U3980 (N_3980,N_3755,N_3884);
and U3981 (N_3981,N_3798,N_3795);
or U3982 (N_3982,N_3890,N_3774);
or U3983 (N_3983,N_3829,N_3868);
and U3984 (N_3984,N_3820,N_3766);
or U3985 (N_3985,N_3813,N_3833);
nand U3986 (N_3986,N_3818,N_3885);
and U3987 (N_3987,N_3808,N_3830);
nand U3988 (N_3988,N_3888,N_3841);
xnor U3989 (N_3989,N_3809,N_3787);
or U3990 (N_3990,N_3752,N_3807);
and U3991 (N_3991,N_3800,N_3795);
nand U3992 (N_3992,N_3807,N_3760);
or U3993 (N_3993,N_3834,N_3899);
nand U3994 (N_3994,N_3785,N_3776);
or U3995 (N_3995,N_3865,N_3879);
nor U3996 (N_3996,N_3843,N_3849);
or U3997 (N_3997,N_3784,N_3780);
xnor U3998 (N_3998,N_3817,N_3856);
and U3999 (N_3999,N_3850,N_3795);
xnor U4000 (N_4000,N_3784,N_3798);
nand U4001 (N_4001,N_3758,N_3772);
or U4002 (N_4002,N_3840,N_3889);
and U4003 (N_4003,N_3891,N_3803);
xor U4004 (N_4004,N_3765,N_3844);
nor U4005 (N_4005,N_3761,N_3765);
xor U4006 (N_4006,N_3766,N_3762);
or U4007 (N_4007,N_3788,N_3797);
xnor U4008 (N_4008,N_3873,N_3856);
or U4009 (N_4009,N_3894,N_3801);
nand U4010 (N_4010,N_3870,N_3777);
or U4011 (N_4011,N_3780,N_3758);
and U4012 (N_4012,N_3884,N_3794);
nand U4013 (N_4013,N_3820,N_3835);
or U4014 (N_4014,N_3898,N_3884);
nor U4015 (N_4015,N_3759,N_3817);
xor U4016 (N_4016,N_3817,N_3792);
nor U4017 (N_4017,N_3851,N_3882);
nor U4018 (N_4018,N_3889,N_3776);
xnor U4019 (N_4019,N_3862,N_3783);
or U4020 (N_4020,N_3850,N_3765);
nor U4021 (N_4021,N_3896,N_3872);
nor U4022 (N_4022,N_3892,N_3814);
nor U4023 (N_4023,N_3781,N_3879);
and U4024 (N_4024,N_3863,N_3822);
nor U4025 (N_4025,N_3827,N_3899);
or U4026 (N_4026,N_3890,N_3802);
nand U4027 (N_4027,N_3790,N_3854);
nor U4028 (N_4028,N_3751,N_3781);
nor U4029 (N_4029,N_3783,N_3823);
xnor U4030 (N_4030,N_3845,N_3851);
nor U4031 (N_4031,N_3774,N_3810);
nand U4032 (N_4032,N_3751,N_3774);
nor U4033 (N_4033,N_3845,N_3758);
xnor U4034 (N_4034,N_3886,N_3807);
nand U4035 (N_4035,N_3797,N_3870);
nor U4036 (N_4036,N_3829,N_3816);
xnor U4037 (N_4037,N_3844,N_3818);
nand U4038 (N_4038,N_3812,N_3861);
nor U4039 (N_4039,N_3835,N_3766);
nor U4040 (N_4040,N_3775,N_3781);
xor U4041 (N_4041,N_3805,N_3858);
xor U4042 (N_4042,N_3844,N_3823);
or U4043 (N_4043,N_3852,N_3850);
xnor U4044 (N_4044,N_3831,N_3760);
or U4045 (N_4045,N_3819,N_3829);
or U4046 (N_4046,N_3867,N_3836);
or U4047 (N_4047,N_3755,N_3814);
and U4048 (N_4048,N_3897,N_3788);
or U4049 (N_4049,N_3837,N_3854);
nor U4050 (N_4050,N_3965,N_3956);
xnor U4051 (N_4051,N_4006,N_3919);
xor U4052 (N_4052,N_3980,N_3997);
nand U4053 (N_4053,N_3959,N_3926);
or U4054 (N_4054,N_4043,N_3920);
xor U4055 (N_4055,N_4002,N_4005);
xnor U4056 (N_4056,N_3942,N_3989);
xnor U4057 (N_4057,N_3937,N_4041);
nor U4058 (N_4058,N_4025,N_4039);
or U4059 (N_4059,N_3978,N_3916);
nor U4060 (N_4060,N_3909,N_4042);
nor U4061 (N_4061,N_4016,N_3985);
and U4062 (N_4062,N_3975,N_3933);
and U4063 (N_4063,N_4020,N_3990);
or U4064 (N_4064,N_3960,N_4045);
and U4065 (N_4065,N_3945,N_4018);
xor U4066 (N_4066,N_4012,N_3973);
and U4067 (N_4067,N_4015,N_3939);
nand U4068 (N_4068,N_3952,N_3962);
or U4069 (N_4069,N_4032,N_3984);
nand U4070 (N_4070,N_3929,N_3904);
and U4071 (N_4071,N_3982,N_3955);
or U4072 (N_4072,N_3905,N_3961);
nor U4073 (N_4073,N_3999,N_3972);
and U4074 (N_4074,N_3967,N_3996);
xnor U4075 (N_4075,N_3950,N_4017);
and U4076 (N_4076,N_3979,N_3922);
and U4077 (N_4077,N_3969,N_4034);
nor U4078 (N_4078,N_3928,N_4029);
nor U4079 (N_4079,N_3991,N_3940);
and U4080 (N_4080,N_3949,N_3995);
xnor U4081 (N_4081,N_3968,N_3948);
and U4082 (N_4082,N_4009,N_4047);
and U4083 (N_4083,N_3914,N_3958);
and U4084 (N_4084,N_3908,N_3900);
and U4085 (N_4085,N_3983,N_4004);
and U4086 (N_4086,N_3966,N_3970);
nor U4087 (N_4087,N_4038,N_3935);
nor U4088 (N_4088,N_3981,N_3988);
and U4089 (N_4089,N_3925,N_3902);
nor U4090 (N_4090,N_4008,N_3906);
nand U4091 (N_4091,N_3934,N_3917);
nand U4092 (N_4092,N_3943,N_3946);
and U4093 (N_4093,N_4036,N_3915);
and U4094 (N_4094,N_4014,N_4044);
or U4095 (N_4095,N_3930,N_4037);
and U4096 (N_4096,N_3913,N_3907);
and U4097 (N_4097,N_4033,N_3901);
nand U4098 (N_4098,N_3957,N_3927);
nor U4099 (N_4099,N_3931,N_4010);
nand U4100 (N_4100,N_4027,N_3910);
nand U4101 (N_4101,N_3936,N_3971);
nor U4102 (N_4102,N_4011,N_4028);
nor U4103 (N_4103,N_4049,N_4046);
xnor U4104 (N_4104,N_4001,N_4031);
or U4105 (N_4105,N_4013,N_3992);
xor U4106 (N_4106,N_4023,N_4022);
or U4107 (N_4107,N_3986,N_4024);
nor U4108 (N_4108,N_4035,N_3944);
nand U4109 (N_4109,N_3964,N_3954);
nand U4110 (N_4110,N_3976,N_3993);
and U4111 (N_4111,N_4007,N_4000);
nor U4112 (N_4112,N_3938,N_4040);
xor U4113 (N_4113,N_3911,N_4030);
or U4114 (N_4114,N_3923,N_4048);
xnor U4115 (N_4115,N_3998,N_3941);
xnor U4116 (N_4116,N_4026,N_3947);
or U4117 (N_4117,N_3963,N_3918);
or U4118 (N_4118,N_3977,N_3912);
nor U4119 (N_4119,N_3921,N_3974);
nand U4120 (N_4120,N_3903,N_4003);
and U4121 (N_4121,N_3953,N_3994);
or U4122 (N_4122,N_3932,N_3924);
xnor U4123 (N_4123,N_3951,N_4019);
nand U4124 (N_4124,N_3987,N_4021);
and U4125 (N_4125,N_3970,N_3990);
xnor U4126 (N_4126,N_3927,N_3932);
xor U4127 (N_4127,N_3970,N_4038);
nor U4128 (N_4128,N_3950,N_4040);
and U4129 (N_4129,N_4034,N_4003);
nor U4130 (N_4130,N_3977,N_4047);
and U4131 (N_4131,N_4038,N_3930);
nor U4132 (N_4132,N_4020,N_4006);
xnor U4133 (N_4133,N_4031,N_4014);
and U4134 (N_4134,N_3933,N_4044);
and U4135 (N_4135,N_4009,N_4008);
or U4136 (N_4136,N_3966,N_4028);
nand U4137 (N_4137,N_3973,N_3999);
or U4138 (N_4138,N_3927,N_4044);
or U4139 (N_4139,N_3930,N_4005);
nand U4140 (N_4140,N_4037,N_3931);
or U4141 (N_4141,N_4046,N_4023);
or U4142 (N_4142,N_4041,N_3958);
and U4143 (N_4143,N_4035,N_3981);
and U4144 (N_4144,N_3917,N_3974);
or U4145 (N_4145,N_3996,N_3935);
or U4146 (N_4146,N_3917,N_3953);
nor U4147 (N_4147,N_3954,N_3946);
nand U4148 (N_4148,N_3900,N_4022);
or U4149 (N_4149,N_4025,N_3939);
nor U4150 (N_4150,N_3968,N_4024);
and U4151 (N_4151,N_4030,N_3959);
or U4152 (N_4152,N_3986,N_3996);
and U4153 (N_4153,N_4007,N_4018);
nand U4154 (N_4154,N_3995,N_3989);
and U4155 (N_4155,N_3945,N_3976);
or U4156 (N_4156,N_3913,N_3987);
and U4157 (N_4157,N_3963,N_3982);
or U4158 (N_4158,N_3990,N_3950);
and U4159 (N_4159,N_3984,N_4006);
xor U4160 (N_4160,N_4002,N_4015);
or U4161 (N_4161,N_3974,N_3960);
or U4162 (N_4162,N_3960,N_3906);
nand U4163 (N_4163,N_4040,N_4022);
and U4164 (N_4164,N_3963,N_4047);
xor U4165 (N_4165,N_3936,N_4026);
xnor U4166 (N_4166,N_3995,N_4029);
or U4167 (N_4167,N_3902,N_3954);
or U4168 (N_4168,N_3930,N_4008);
xnor U4169 (N_4169,N_3957,N_3960);
or U4170 (N_4170,N_3919,N_3947);
xnor U4171 (N_4171,N_4015,N_4013);
or U4172 (N_4172,N_4032,N_3907);
nand U4173 (N_4173,N_3940,N_3965);
xor U4174 (N_4174,N_3971,N_3934);
or U4175 (N_4175,N_3924,N_4029);
or U4176 (N_4176,N_3909,N_3959);
xnor U4177 (N_4177,N_4030,N_3991);
nand U4178 (N_4178,N_4033,N_3902);
and U4179 (N_4179,N_3954,N_3909);
and U4180 (N_4180,N_3930,N_4021);
or U4181 (N_4181,N_3978,N_3999);
nand U4182 (N_4182,N_3914,N_3909);
nand U4183 (N_4183,N_3989,N_4019);
nand U4184 (N_4184,N_3925,N_4016);
or U4185 (N_4185,N_4038,N_3955);
or U4186 (N_4186,N_3988,N_4022);
or U4187 (N_4187,N_3989,N_3968);
nor U4188 (N_4188,N_4034,N_3982);
nand U4189 (N_4189,N_3998,N_3918);
or U4190 (N_4190,N_3989,N_3911);
and U4191 (N_4191,N_3944,N_4037);
nand U4192 (N_4192,N_4014,N_4040);
or U4193 (N_4193,N_3934,N_3979);
and U4194 (N_4194,N_3931,N_3955);
nor U4195 (N_4195,N_4033,N_3965);
nor U4196 (N_4196,N_4049,N_3918);
or U4197 (N_4197,N_4049,N_4000);
or U4198 (N_4198,N_3987,N_4002);
nand U4199 (N_4199,N_3955,N_3994);
nand U4200 (N_4200,N_4055,N_4082);
nand U4201 (N_4201,N_4175,N_4177);
xor U4202 (N_4202,N_4072,N_4089);
and U4203 (N_4203,N_4108,N_4060);
and U4204 (N_4204,N_4078,N_4166);
nand U4205 (N_4205,N_4113,N_4173);
xor U4206 (N_4206,N_4097,N_4120);
xnor U4207 (N_4207,N_4121,N_4189);
and U4208 (N_4208,N_4056,N_4066);
and U4209 (N_4209,N_4172,N_4086);
nand U4210 (N_4210,N_4084,N_4099);
nor U4211 (N_4211,N_4143,N_4092);
nand U4212 (N_4212,N_4079,N_4083);
xor U4213 (N_4213,N_4116,N_4186);
xor U4214 (N_4214,N_4162,N_4180);
nand U4215 (N_4215,N_4137,N_4106);
nor U4216 (N_4216,N_4080,N_4102);
nor U4217 (N_4217,N_4155,N_4051);
xnor U4218 (N_4218,N_4168,N_4095);
nand U4219 (N_4219,N_4159,N_4067);
or U4220 (N_4220,N_4178,N_4076);
or U4221 (N_4221,N_4194,N_4052);
and U4222 (N_4222,N_4134,N_4088);
xor U4223 (N_4223,N_4061,N_4187);
nor U4224 (N_4224,N_4112,N_4125);
xor U4225 (N_4225,N_4109,N_4058);
xor U4226 (N_4226,N_4195,N_4114);
nor U4227 (N_4227,N_4149,N_4105);
xnor U4228 (N_4228,N_4179,N_4167);
nor U4229 (N_4229,N_4142,N_4190);
nor U4230 (N_4230,N_4164,N_4151);
and U4231 (N_4231,N_4132,N_4062);
or U4232 (N_4232,N_4170,N_4160);
and U4233 (N_4233,N_4139,N_4100);
or U4234 (N_4234,N_4050,N_4153);
and U4235 (N_4235,N_4127,N_4059);
nor U4236 (N_4236,N_4115,N_4140);
or U4237 (N_4237,N_4183,N_4117);
xnor U4238 (N_4238,N_4057,N_4145);
xor U4239 (N_4239,N_4182,N_4193);
nand U4240 (N_4240,N_4101,N_4133);
nor U4241 (N_4241,N_4053,N_4081);
or U4242 (N_4242,N_4104,N_4073);
xnor U4243 (N_4243,N_4070,N_4138);
and U4244 (N_4244,N_4161,N_4069);
or U4245 (N_4245,N_4157,N_4129);
or U4246 (N_4246,N_4174,N_4064);
and U4247 (N_4247,N_4093,N_4103);
and U4248 (N_4248,N_4146,N_4181);
nor U4249 (N_4249,N_4135,N_4148);
and U4250 (N_4250,N_4094,N_4128);
nand U4251 (N_4251,N_4123,N_4131);
and U4252 (N_4252,N_4163,N_4147);
nand U4253 (N_4253,N_4171,N_4185);
xnor U4254 (N_4254,N_4154,N_4199);
nand U4255 (N_4255,N_4150,N_4165);
and U4256 (N_4256,N_4107,N_4191);
xor U4257 (N_4257,N_4098,N_4071);
nor U4258 (N_4258,N_4111,N_4158);
nor U4259 (N_4259,N_4118,N_4090);
nand U4260 (N_4260,N_4119,N_4184);
nand U4261 (N_4261,N_4136,N_4091);
xnor U4262 (N_4262,N_4122,N_4192);
and U4263 (N_4263,N_4110,N_4152);
nor U4264 (N_4264,N_4054,N_4077);
nor U4265 (N_4265,N_4063,N_4198);
or U4266 (N_4266,N_4176,N_4141);
nor U4267 (N_4267,N_4156,N_4085);
nand U4268 (N_4268,N_4188,N_4197);
and U4269 (N_4269,N_4196,N_4096);
nor U4270 (N_4270,N_4126,N_4074);
or U4271 (N_4271,N_4065,N_4124);
or U4272 (N_4272,N_4169,N_4075);
and U4273 (N_4273,N_4144,N_4068);
nand U4274 (N_4274,N_4130,N_4087);
or U4275 (N_4275,N_4157,N_4193);
nand U4276 (N_4276,N_4094,N_4054);
or U4277 (N_4277,N_4071,N_4076);
and U4278 (N_4278,N_4072,N_4159);
nand U4279 (N_4279,N_4082,N_4139);
nand U4280 (N_4280,N_4097,N_4050);
nor U4281 (N_4281,N_4153,N_4077);
nor U4282 (N_4282,N_4070,N_4123);
nand U4283 (N_4283,N_4102,N_4186);
or U4284 (N_4284,N_4104,N_4164);
xor U4285 (N_4285,N_4117,N_4195);
and U4286 (N_4286,N_4142,N_4185);
and U4287 (N_4287,N_4149,N_4134);
xor U4288 (N_4288,N_4168,N_4177);
nand U4289 (N_4289,N_4073,N_4179);
or U4290 (N_4290,N_4099,N_4054);
nor U4291 (N_4291,N_4078,N_4054);
xnor U4292 (N_4292,N_4074,N_4153);
xnor U4293 (N_4293,N_4140,N_4154);
nand U4294 (N_4294,N_4172,N_4122);
xor U4295 (N_4295,N_4065,N_4115);
nor U4296 (N_4296,N_4132,N_4176);
xnor U4297 (N_4297,N_4090,N_4074);
or U4298 (N_4298,N_4110,N_4137);
and U4299 (N_4299,N_4054,N_4068);
nand U4300 (N_4300,N_4142,N_4133);
nor U4301 (N_4301,N_4061,N_4121);
nor U4302 (N_4302,N_4150,N_4199);
or U4303 (N_4303,N_4094,N_4066);
or U4304 (N_4304,N_4147,N_4159);
nand U4305 (N_4305,N_4197,N_4130);
nand U4306 (N_4306,N_4067,N_4122);
nor U4307 (N_4307,N_4107,N_4116);
xor U4308 (N_4308,N_4077,N_4057);
nand U4309 (N_4309,N_4066,N_4149);
and U4310 (N_4310,N_4181,N_4178);
or U4311 (N_4311,N_4113,N_4121);
or U4312 (N_4312,N_4063,N_4056);
nand U4313 (N_4313,N_4145,N_4066);
and U4314 (N_4314,N_4145,N_4172);
nor U4315 (N_4315,N_4137,N_4123);
nor U4316 (N_4316,N_4119,N_4062);
or U4317 (N_4317,N_4176,N_4105);
xor U4318 (N_4318,N_4119,N_4135);
or U4319 (N_4319,N_4116,N_4087);
nand U4320 (N_4320,N_4158,N_4105);
nand U4321 (N_4321,N_4164,N_4115);
or U4322 (N_4322,N_4112,N_4168);
nand U4323 (N_4323,N_4156,N_4084);
and U4324 (N_4324,N_4100,N_4109);
or U4325 (N_4325,N_4154,N_4134);
nand U4326 (N_4326,N_4195,N_4050);
and U4327 (N_4327,N_4078,N_4058);
nand U4328 (N_4328,N_4198,N_4073);
and U4329 (N_4329,N_4168,N_4169);
and U4330 (N_4330,N_4150,N_4164);
and U4331 (N_4331,N_4070,N_4061);
or U4332 (N_4332,N_4146,N_4067);
or U4333 (N_4333,N_4100,N_4156);
nor U4334 (N_4334,N_4050,N_4073);
nor U4335 (N_4335,N_4140,N_4108);
nor U4336 (N_4336,N_4074,N_4121);
nand U4337 (N_4337,N_4085,N_4124);
xnor U4338 (N_4338,N_4135,N_4187);
xor U4339 (N_4339,N_4078,N_4070);
and U4340 (N_4340,N_4122,N_4170);
nand U4341 (N_4341,N_4109,N_4082);
or U4342 (N_4342,N_4157,N_4174);
or U4343 (N_4343,N_4103,N_4184);
nand U4344 (N_4344,N_4165,N_4103);
and U4345 (N_4345,N_4118,N_4135);
or U4346 (N_4346,N_4159,N_4155);
and U4347 (N_4347,N_4122,N_4159);
nand U4348 (N_4348,N_4066,N_4098);
nor U4349 (N_4349,N_4105,N_4065);
nand U4350 (N_4350,N_4320,N_4213);
and U4351 (N_4351,N_4240,N_4277);
nand U4352 (N_4352,N_4235,N_4338);
and U4353 (N_4353,N_4255,N_4200);
or U4354 (N_4354,N_4348,N_4204);
and U4355 (N_4355,N_4268,N_4206);
nand U4356 (N_4356,N_4284,N_4209);
xor U4357 (N_4357,N_4290,N_4260);
and U4358 (N_4358,N_4286,N_4304);
xnor U4359 (N_4359,N_4230,N_4251);
xnor U4360 (N_4360,N_4258,N_4214);
nor U4361 (N_4361,N_4327,N_4229);
nand U4362 (N_4362,N_4246,N_4274);
and U4363 (N_4363,N_4281,N_4318);
nor U4364 (N_4364,N_4310,N_4216);
xnor U4365 (N_4365,N_4324,N_4344);
nor U4366 (N_4366,N_4237,N_4263);
nor U4367 (N_4367,N_4280,N_4288);
or U4368 (N_4368,N_4341,N_4339);
nor U4369 (N_4369,N_4331,N_4221);
or U4370 (N_4370,N_4308,N_4241);
nand U4371 (N_4371,N_4224,N_4223);
nand U4372 (N_4372,N_4326,N_4262);
or U4373 (N_4373,N_4231,N_4215);
nand U4374 (N_4374,N_4249,N_4259);
nand U4375 (N_4375,N_4265,N_4301);
and U4376 (N_4376,N_4305,N_4342);
nand U4377 (N_4377,N_4220,N_4325);
or U4378 (N_4378,N_4222,N_4210);
or U4379 (N_4379,N_4269,N_4317);
nand U4380 (N_4380,N_4270,N_4332);
and U4381 (N_4381,N_4303,N_4302);
and U4382 (N_4382,N_4296,N_4217);
and U4383 (N_4383,N_4218,N_4212);
nand U4384 (N_4384,N_4208,N_4349);
nand U4385 (N_4385,N_4239,N_4245);
nand U4386 (N_4386,N_4252,N_4337);
nand U4387 (N_4387,N_4219,N_4232);
nor U4388 (N_4388,N_4244,N_4287);
and U4389 (N_4389,N_4335,N_4295);
or U4390 (N_4390,N_4329,N_4247);
or U4391 (N_4391,N_4264,N_4340);
nand U4392 (N_4392,N_4333,N_4307);
nor U4393 (N_4393,N_4309,N_4312);
nand U4394 (N_4394,N_4273,N_4289);
nor U4395 (N_4395,N_4336,N_4306);
or U4396 (N_4396,N_4202,N_4347);
nand U4397 (N_4397,N_4233,N_4248);
nand U4398 (N_4398,N_4300,N_4238);
xnor U4399 (N_4399,N_4314,N_4285);
xor U4400 (N_4400,N_4279,N_4322);
or U4401 (N_4401,N_4294,N_4227);
or U4402 (N_4402,N_4315,N_4253);
nand U4403 (N_4403,N_4275,N_4323);
nand U4404 (N_4404,N_4278,N_4254);
nor U4405 (N_4405,N_4243,N_4313);
nor U4406 (N_4406,N_4234,N_4228);
and U4407 (N_4407,N_4226,N_4250);
nand U4408 (N_4408,N_4211,N_4321);
nor U4409 (N_4409,N_4345,N_4261);
or U4410 (N_4410,N_4319,N_4266);
nor U4411 (N_4411,N_4297,N_4225);
nand U4412 (N_4412,N_4256,N_4205);
nor U4413 (N_4413,N_4298,N_4299);
or U4414 (N_4414,N_4291,N_4201);
xnor U4415 (N_4415,N_4282,N_4316);
and U4416 (N_4416,N_4334,N_4328);
nand U4417 (N_4417,N_4293,N_4330);
nand U4418 (N_4418,N_4283,N_4346);
nand U4419 (N_4419,N_4311,N_4257);
xnor U4420 (N_4420,N_4292,N_4207);
nand U4421 (N_4421,N_4203,N_4343);
xor U4422 (N_4422,N_4242,N_4271);
nand U4423 (N_4423,N_4236,N_4272);
nand U4424 (N_4424,N_4276,N_4267);
nand U4425 (N_4425,N_4299,N_4273);
xor U4426 (N_4426,N_4283,N_4223);
nor U4427 (N_4427,N_4313,N_4273);
xor U4428 (N_4428,N_4294,N_4345);
and U4429 (N_4429,N_4301,N_4309);
and U4430 (N_4430,N_4254,N_4228);
xor U4431 (N_4431,N_4233,N_4264);
nor U4432 (N_4432,N_4287,N_4213);
or U4433 (N_4433,N_4252,N_4343);
nand U4434 (N_4434,N_4225,N_4230);
nor U4435 (N_4435,N_4246,N_4329);
and U4436 (N_4436,N_4309,N_4248);
nand U4437 (N_4437,N_4296,N_4299);
or U4438 (N_4438,N_4211,N_4318);
xor U4439 (N_4439,N_4273,N_4344);
or U4440 (N_4440,N_4333,N_4275);
nand U4441 (N_4441,N_4217,N_4290);
nand U4442 (N_4442,N_4285,N_4313);
or U4443 (N_4443,N_4316,N_4315);
nor U4444 (N_4444,N_4284,N_4328);
nand U4445 (N_4445,N_4293,N_4272);
xnor U4446 (N_4446,N_4227,N_4238);
nand U4447 (N_4447,N_4348,N_4328);
nand U4448 (N_4448,N_4286,N_4315);
nor U4449 (N_4449,N_4303,N_4222);
and U4450 (N_4450,N_4320,N_4227);
or U4451 (N_4451,N_4331,N_4218);
and U4452 (N_4452,N_4206,N_4263);
nand U4453 (N_4453,N_4208,N_4282);
and U4454 (N_4454,N_4205,N_4331);
or U4455 (N_4455,N_4241,N_4277);
and U4456 (N_4456,N_4274,N_4259);
xnor U4457 (N_4457,N_4290,N_4270);
nor U4458 (N_4458,N_4316,N_4321);
and U4459 (N_4459,N_4285,N_4251);
nor U4460 (N_4460,N_4306,N_4349);
and U4461 (N_4461,N_4213,N_4242);
nand U4462 (N_4462,N_4278,N_4234);
xor U4463 (N_4463,N_4219,N_4323);
nand U4464 (N_4464,N_4266,N_4223);
xnor U4465 (N_4465,N_4324,N_4275);
nor U4466 (N_4466,N_4292,N_4252);
and U4467 (N_4467,N_4261,N_4284);
xor U4468 (N_4468,N_4286,N_4252);
nor U4469 (N_4469,N_4207,N_4327);
nor U4470 (N_4470,N_4321,N_4270);
nand U4471 (N_4471,N_4233,N_4251);
xor U4472 (N_4472,N_4305,N_4257);
nand U4473 (N_4473,N_4314,N_4206);
or U4474 (N_4474,N_4267,N_4242);
or U4475 (N_4475,N_4271,N_4251);
xor U4476 (N_4476,N_4222,N_4347);
and U4477 (N_4477,N_4277,N_4267);
xor U4478 (N_4478,N_4335,N_4258);
nand U4479 (N_4479,N_4319,N_4307);
or U4480 (N_4480,N_4274,N_4227);
nand U4481 (N_4481,N_4289,N_4340);
and U4482 (N_4482,N_4236,N_4275);
or U4483 (N_4483,N_4226,N_4263);
xor U4484 (N_4484,N_4306,N_4262);
xnor U4485 (N_4485,N_4203,N_4253);
and U4486 (N_4486,N_4238,N_4280);
and U4487 (N_4487,N_4335,N_4251);
and U4488 (N_4488,N_4302,N_4254);
xor U4489 (N_4489,N_4256,N_4245);
or U4490 (N_4490,N_4316,N_4230);
and U4491 (N_4491,N_4258,N_4337);
xor U4492 (N_4492,N_4309,N_4205);
nor U4493 (N_4493,N_4247,N_4340);
xor U4494 (N_4494,N_4252,N_4321);
xor U4495 (N_4495,N_4348,N_4261);
nand U4496 (N_4496,N_4273,N_4308);
xor U4497 (N_4497,N_4243,N_4319);
xor U4498 (N_4498,N_4315,N_4234);
nor U4499 (N_4499,N_4289,N_4266);
nor U4500 (N_4500,N_4413,N_4434);
nor U4501 (N_4501,N_4438,N_4495);
xor U4502 (N_4502,N_4461,N_4424);
nand U4503 (N_4503,N_4457,N_4402);
nand U4504 (N_4504,N_4427,N_4436);
nor U4505 (N_4505,N_4359,N_4445);
or U4506 (N_4506,N_4405,N_4395);
or U4507 (N_4507,N_4426,N_4365);
or U4508 (N_4508,N_4475,N_4455);
xnor U4509 (N_4509,N_4448,N_4433);
nand U4510 (N_4510,N_4493,N_4383);
nand U4511 (N_4511,N_4488,N_4393);
and U4512 (N_4512,N_4418,N_4372);
and U4513 (N_4513,N_4358,N_4420);
or U4514 (N_4514,N_4469,N_4381);
nand U4515 (N_4515,N_4494,N_4463);
or U4516 (N_4516,N_4350,N_4437);
nand U4517 (N_4517,N_4392,N_4378);
xor U4518 (N_4518,N_4407,N_4484);
nand U4519 (N_4519,N_4357,N_4384);
nand U4520 (N_4520,N_4367,N_4412);
xor U4521 (N_4521,N_4399,N_4361);
nand U4522 (N_4522,N_4375,N_4444);
xnor U4523 (N_4523,N_4492,N_4496);
nor U4524 (N_4524,N_4397,N_4389);
nand U4525 (N_4525,N_4388,N_4429);
nor U4526 (N_4526,N_4370,N_4440);
nand U4527 (N_4527,N_4422,N_4451);
and U4528 (N_4528,N_4369,N_4385);
nor U4529 (N_4529,N_4462,N_4483);
nand U4530 (N_4530,N_4453,N_4362);
xnor U4531 (N_4531,N_4368,N_4481);
xor U4532 (N_4532,N_4460,N_4442);
nor U4533 (N_4533,N_4360,N_4421);
nor U4534 (N_4534,N_4431,N_4439);
nor U4535 (N_4535,N_4394,N_4473);
or U4536 (N_4536,N_4364,N_4497);
xor U4537 (N_4537,N_4356,N_4428);
xor U4538 (N_4538,N_4482,N_4472);
nand U4539 (N_4539,N_4355,N_4477);
xnor U4540 (N_4540,N_4404,N_4478);
nand U4541 (N_4541,N_4471,N_4386);
nand U4542 (N_4542,N_4470,N_4398);
nor U4543 (N_4543,N_4400,N_4425);
xor U4544 (N_4544,N_4474,N_4417);
nor U4545 (N_4545,N_4464,N_4351);
xnor U4546 (N_4546,N_4485,N_4486);
and U4547 (N_4547,N_4371,N_4387);
nor U4548 (N_4548,N_4353,N_4377);
xor U4549 (N_4549,N_4467,N_4376);
xnor U4550 (N_4550,N_4458,N_4466);
xor U4551 (N_4551,N_4373,N_4459);
and U4552 (N_4552,N_4415,N_4430);
xor U4553 (N_4553,N_4366,N_4499);
and U4554 (N_4554,N_4380,N_4450);
and U4555 (N_4555,N_4409,N_4490);
nand U4556 (N_4556,N_4476,N_4454);
nand U4557 (N_4557,N_4363,N_4396);
nor U4558 (N_4558,N_4449,N_4452);
and U4559 (N_4559,N_4408,N_4406);
or U4560 (N_4560,N_4411,N_4435);
and U4561 (N_4561,N_4391,N_4468);
and U4562 (N_4562,N_4456,N_4401);
and U4563 (N_4563,N_4465,N_4447);
nand U4564 (N_4564,N_4374,N_4479);
nor U4565 (N_4565,N_4487,N_4352);
nor U4566 (N_4566,N_4382,N_4498);
and U4567 (N_4567,N_4441,N_4414);
and U4568 (N_4568,N_4443,N_4403);
and U4569 (N_4569,N_4390,N_4423);
or U4570 (N_4570,N_4416,N_4354);
xor U4571 (N_4571,N_4446,N_4480);
xor U4572 (N_4572,N_4491,N_4410);
or U4573 (N_4573,N_4379,N_4419);
or U4574 (N_4574,N_4489,N_4432);
xor U4575 (N_4575,N_4478,N_4497);
or U4576 (N_4576,N_4361,N_4424);
nand U4577 (N_4577,N_4442,N_4419);
nor U4578 (N_4578,N_4377,N_4358);
nand U4579 (N_4579,N_4473,N_4358);
or U4580 (N_4580,N_4416,N_4439);
xor U4581 (N_4581,N_4470,N_4419);
and U4582 (N_4582,N_4459,N_4447);
and U4583 (N_4583,N_4360,N_4432);
or U4584 (N_4584,N_4454,N_4485);
xor U4585 (N_4585,N_4357,N_4374);
nand U4586 (N_4586,N_4497,N_4460);
xnor U4587 (N_4587,N_4451,N_4376);
xnor U4588 (N_4588,N_4488,N_4363);
or U4589 (N_4589,N_4405,N_4458);
or U4590 (N_4590,N_4381,N_4473);
xnor U4591 (N_4591,N_4444,N_4385);
and U4592 (N_4592,N_4364,N_4412);
and U4593 (N_4593,N_4353,N_4384);
and U4594 (N_4594,N_4427,N_4388);
nor U4595 (N_4595,N_4424,N_4366);
xnor U4596 (N_4596,N_4432,N_4380);
nor U4597 (N_4597,N_4414,N_4363);
or U4598 (N_4598,N_4424,N_4363);
nor U4599 (N_4599,N_4453,N_4378);
or U4600 (N_4600,N_4385,N_4367);
nand U4601 (N_4601,N_4366,N_4382);
nand U4602 (N_4602,N_4460,N_4368);
or U4603 (N_4603,N_4382,N_4467);
or U4604 (N_4604,N_4373,N_4417);
or U4605 (N_4605,N_4409,N_4426);
and U4606 (N_4606,N_4484,N_4370);
nor U4607 (N_4607,N_4378,N_4416);
nor U4608 (N_4608,N_4373,N_4353);
and U4609 (N_4609,N_4389,N_4432);
nor U4610 (N_4610,N_4437,N_4395);
xnor U4611 (N_4611,N_4359,N_4457);
and U4612 (N_4612,N_4438,N_4390);
nor U4613 (N_4613,N_4351,N_4434);
and U4614 (N_4614,N_4472,N_4457);
and U4615 (N_4615,N_4489,N_4415);
xor U4616 (N_4616,N_4393,N_4494);
nor U4617 (N_4617,N_4367,N_4428);
xor U4618 (N_4618,N_4381,N_4428);
or U4619 (N_4619,N_4481,N_4426);
nand U4620 (N_4620,N_4370,N_4433);
or U4621 (N_4621,N_4420,N_4389);
and U4622 (N_4622,N_4485,N_4478);
xnor U4623 (N_4623,N_4371,N_4392);
or U4624 (N_4624,N_4392,N_4434);
nand U4625 (N_4625,N_4396,N_4420);
or U4626 (N_4626,N_4465,N_4415);
nand U4627 (N_4627,N_4499,N_4421);
nand U4628 (N_4628,N_4374,N_4392);
nand U4629 (N_4629,N_4436,N_4430);
or U4630 (N_4630,N_4448,N_4481);
nor U4631 (N_4631,N_4357,N_4448);
nor U4632 (N_4632,N_4445,N_4363);
nand U4633 (N_4633,N_4455,N_4416);
xor U4634 (N_4634,N_4400,N_4358);
nor U4635 (N_4635,N_4420,N_4386);
or U4636 (N_4636,N_4409,N_4372);
or U4637 (N_4637,N_4393,N_4361);
nand U4638 (N_4638,N_4397,N_4406);
nor U4639 (N_4639,N_4443,N_4484);
nor U4640 (N_4640,N_4475,N_4473);
and U4641 (N_4641,N_4413,N_4363);
nor U4642 (N_4642,N_4368,N_4394);
nor U4643 (N_4643,N_4380,N_4477);
nand U4644 (N_4644,N_4448,N_4370);
or U4645 (N_4645,N_4478,N_4447);
xor U4646 (N_4646,N_4391,N_4412);
nand U4647 (N_4647,N_4469,N_4427);
or U4648 (N_4648,N_4414,N_4452);
and U4649 (N_4649,N_4472,N_4498);
and U4650 (N_4650,N_4602,N_4579);
and U4651 (N_4651,N_4548,N_4608);
nor U4652 (N_4652,N_4636,N_4582);
nand U4653 (N_4653,N_4613,N_4624);
and U4654 (N_4654,N_4633,N_4571);
nand U4655 (N_4655,N_4518,N_4589);
and U4656 (N_4656,N_4563,N_4632);
xor U4657 (N_4657,N_4533,N_4527);
xnor U4658 (N_4658,N_4596,N_4567);
nor U4659 (N_4659,N_4616,N_4587);
xnor U4660 (N_4660,N_4551,N_4509);
nor U4661 (N_4661,N_4619,N_4542);
nand U4662 (N_4662,N_4520,N_4645);
nand U4663 (N_4663,N_4559,N_4530);
and U4664 (N_4664,N_4510,N_4560);
nor U4665 (N_4665,N_4647,N_4588);
xnor U4666 (N_4666,N_4597,N_4547);
nor U4667 (N_4667,N_4543,N_4550);
xnor U4668 (N_4668,N_4515,N_4594);
xnor U4669 (N_4669,N_4521,N_4607);
nor U4670 (N_4670,N_4600,N_4611);
nand U4671 (N_4671,N_4536,N_4505);
and U4672 (N_4672,N_4554,N_4625);
and U4673 (N_4673,N_4541,N_4546);
nor U4674 (N_4674,N_4627,N_4524);
nand U4675 (N_4675,N_4584,N_4561);
nand U4676 (N_4676,N_4612,N_4593);
and U4677 (N_4677,N_4644,N_4605);
xnor U4678 (N_4678,N_4540,N_4620);
or U4679 (N_4679,N_4557,N_4523);
nand U4680 (N_4680,N_4519,N_4618);
or U4681 (N_4681,N_4570,N_4648);
nor U4682 (N_4682,N_4630,N_4506);
or U4683 (N_4683,N_4532,N_4553);
nand U4684 (N_4684,N_4501,N_4634);
or U4685 (N_4685,N_4535,N_4511);
or U4686 (N_4686,N_4604,N_4614);
nand U4687 (N_4687,N_4628,N_4512);
xnor U4688 (N_4688,N_4640,N_4615);
nand U4689 (N_4689,N_4569,N_4599);
nor U4690 (N_4690,N_4649,N_4573);
or U4691 (N_4691,N_4646,N_4622);
nand U4692 (N_4692,N_4603,N_4502);
xor U4693 (N_4693,N_4639,N_4525);
xor U4694 (N_4694,N_4508,N_4552);
and U4695 (N_4695,N_4631,N_4568);
nor U4696 (N_4696,N_4601,N_4606);
nand U4697 (N_4697,N_4516,N_4591);
xor U4698 (N_4698,N_4609,N_4642);
nor U4699 (N_4699,N_4580,N_4595);
and U4700 (N_4700,N_4590,N_4572);
xor U4701 (N_4701,N_4555,N_4514);
and U4702 (N_4702,N_4534,N_4507);
nand U4703 (N_4703,N_4577,N_4539);
and U4704 (N_4704,N_4643,N_4575);
or U4705 (N_4705,N_4621,N_4623);
nand U4706 (N_4706,N_4556,N_4637);
nand U4707 (N_4707,N_4517,N_4562);
nor U4708 (N_4708,N_4549,N_4522);
or U4709 (N_4709,N_4578,N_4629);
nand U4710 (N_4710,N_4526,N_4610);
and U4711 (N_4711,N_4531,N_4592);
xnor U4712 (N_4712,N_4617,N_4544);
nand U4713 (N_4713,N_4583,N_4564);
and U4714 (N_4714,N_4513,N_4529);
nor U4715 (N_4715,N_4566,N_4598);
xor U4716 (N_4716,N_4574,N_4638);
nor U4717 (N_4717,N_4545,N_4635);
nand U4718 (N_4718,N_4581,N_4503);
xor U4719 (N_4719,N_4537,N_4500);
and U4720 (N_4720,N_4565,N_4626);
or U4721 (N_4721,N_4504,N_4586);
nor U4722 (N_4722,N_4558,N_4641);
nand U4723 (N_4723,N_4528,N_4585);
or U4724 (N_4724,N_4538,N_4576);
nand U4725 (N_4725,N_4512,N_4537);
nand U4726 (N_4726,N_4527,N_4621);
xor U4727 (N_4727,N_4618,N_4641);
nor U4728 (N_4728,N_4637,N_4602);
or U4729 (N_4729,N_4507,N_4629);
or U4730 (N_4730,N_4629,N_4534);
nand U4731 (N_4731,N_4580,N_4576);
nand U4732 (N_4732,N_4571,N_4520);
xor U4733 (N_4733,N_4548,N_4544);
nand U4734 (N_4734,N_4626,N_4637);
or U4735 (N_4735,N_4500,N_4637);
or U4736 (N_4736,N_4588,N_4609);
and U4737 (N_4737,N_4531,N_4516);
or U4738 (N_4738,N_4590,N_4608);
nor U4739 (N_4739,N_4576,N_4579);
xnor U4740 (N_4740,N_4537,N_4637);
nor U4741 (N_4741,N_4561,N_4501);
nand U4742 (N_4742,N_4523,N_4579);
nor U4743 (N_4743,N_4594,N_4514);
or U4744 (N_4744,N_4558,N_4528);
or U4745 (N_4745,N_4622,N_4528);
xor U4746 (N_4746,N_4516,N_4618);
nand U4747 (N_4747,N_4568,N_4541);
and U4748 (N_4748,N_4614,N_4636);
xnor U4749 (N_4749,N_4501,N_4649);
nor U4750 (N_4750,N_4578,N_4622);
nor U4751 (N_4751,N_4630,N_4546);
xnor U4752 (N_4752,N_4538,N_4528);
nor U4753 (N_4753,N_4593,N_4507);
xnor U4754 (N_4754,N_4613,N_4577);
nand U4755 (N_4755,N_4628,N_4585);
and U4756 (N_4756,N_4636,N_4591);
or U4757 (N_4757,N_4583,N_4524);
nand U4758 (N_4758,N_4645,N_4540);
nand U4759 (N_4759,N_4613,N_4643);
nand U4760 (N_4760,N_4522,N_4632);
or U4761 (N_4761,N_4543,N_4625);
nand U4762 (N_4762,N_4504,N_4607);
or U4763 (N_4763,N_4604,N_4533);
or U4764 (N_4764,N_4604,N_4621);
xor U4765 (N_4765,N_4515,N_4581);
and U4766 (N_4766,N_4520,N_4542);
nand U4767 (N_4767,N_4560,N_4554);
nor U4768 (N_4768,N_4584,N_4602);
or U4769 (N_4769,N_4628,N_4611);
and U4770 (N_4770,N_4644,N_4538);
nor U4771 (N_4771,N_4503,N_4627);
or U4772 (N_4772,N_4591,N_4500);
and U4773 (N_4773,N_4648,N_4582);
or U4774 (N_4774,N_4548,N_4602);
nor U4775 (N_4775,N_4582,N_4600);
or U4776 (N_4776,N_4609,N_4648);
xnor U4777 (N_4777,N_4641,N_4556);
nor U4778 (N_4778,N_4580,N_4515);
xnor U4779 (N_4779,N_4505,N_4563);
or U4780 (N_4780,N_4514,N_4586);
or U4781 (N_4781,N_4580,N_4601);
and U4782 (N_4782,N_4510,N_4580);
and U4783 (N_4783,N_4619,N_4567);
or U4784 (N_4784,N_4632,N_4609);
or U4785 (N_4785,N_4647,N_4631);
or U4786 (N_4786,N_4572,N_4616);
xnor U4787 (N_4787,N_4633,N_4606);
or U4788 (N_4788,N_4522,N_4533);
nor U4789 (N_4789,N_4546,N_4574);
or U4790 (N_4790,N_4512,N_4538);
or U4791 (N_4791,N_4532,N_4580);
and U4792 (N_4792,N_4582,N_4605);
nand U4793 (N_4793,N_4616,N_4573);
xnor U4794 (N_4794,N_4615,N_4514);
and U4795 (N_4795,N_4607,N_4568);
xnor U4796 (N_4796,N_4610,N_4507);
xor U4797 (N_4797,N_4602,N_4610);
and U4798 (N_4798,N_4558,N_4531);
and U4799 (N_4799,N_4545,N_4596);
nand U4800 (N_4800,N_4689,N_4702);
and U4801 (N_4801,N_4701,N_4749);
xor U4802 (N_4802,N_4756,N_4695);
and U4803 (N_4803,N_4653,N_4725);
or U4804 (N_4804,N_4747,N_4736);
and U4805 (N_4805,N_4742,N_4762);
nor U4806 (N_4806,N_4670,N_4658);
or U4807 (N_4807,N_4730,N_4799);
xnor U4808 (N_4808,N_4726,N_4729);
and U4809 (N_4809,N_4697,N_4748);
or U4810 (N_4810,N_4751,N_4798);
xor U4811 (N_4811,N_4700,N_4755);
nor U4812 (N_4812,N_4754,N_4757);
or U4813 (N_4813,N_4792,N_4667);
or U4814 (N_4814,N_4680,N_4685);
nor U4815 (N_4815,N_4699,N_4777);
nor U4816 (N_4816,N_4740,N_4719);
xor U4817 (N_4817,N_4716,N_4674);
nand U4818 (N_4818,N_4779,N_4704);
nor U4819 (N_4819,N_4795,N_4760);
nand U4820 (N_4820,N_4723,N_4659);
nand U4821 (N_4821,N_4772,N_4678);
nor U4822 (N_4822,N_4744,N_4666);
nand U4823 (N_4823,N_4711,N_4710);
xor U4824 (N_4824,N_4722,N_4721);
or U4825 (N_4825,N_4652,N_4693);
xnor U4826 (N_4826,N_4684,N_4768);
or U4827 (N_4827,N_4797,N_4787);
and U4828 (N_4828,N_4793,N_4767);
or U4829 (N_4829,N_4675,N_4679);
nor U4830 (N_4830,N_4731,N_4746);
and U4831 (N_4831,N_4750,N_4681);
xor U4832 (N_4832,N_4656,N_4738);
and U4833 (N_4833,N_4717,N_4770);
xnor U4834 (N_4834,N_4790,N_4705);
nand U4835 (N_4835,N_4664,N_4739);
nand U4836 (N_4836,N_4724,N_4673);
nor U4837 (N_4837,N_4769,N_4708);
and U4838 (N_4838,N_4782,N_4672);
and U4839 (N_4839,N_4655,N_4669);
nor U4840 (N_4840,N_4773,N_4683);
or U4841 (N_4841,N_4758,N_4654);
nand U4842 (N_4842,N_4650,N_4663);
or U4843 (N_4843,N_4691,N_4706);
xor U4844 (N_4844,N_4774,N_4682);
nand U4845 (N_4845,N_4692,N_4671);
xor U4846 (N_4846,N_4686,N_4784);
nor U4847 (N_4847,N_4698,N_4665);
or U4848 (N_4848,N_4776,N_4752);
nand U4849 (N_4849,N_4660,N_4789);
nand U4850 (N_4850,N_4761,N_4796);
xnor U4851 (N_4851,N_4712,N_4728);
nand U4852 (N_4852,N_4668,N_4662);
nor U4853 (N_4853,N_4696,N_4709);
and U4854 (N_4854,N_4735,N_4713);
or U4855 (N_4855,N_4775,N_4661);
nand U4856 (N_4856,N_4786,N_4764);
nor U4857 (N_4857,N_4732,N_4765);
nor U4858 (N_4858,N_4657,N_4720);
or U4859 (N_4859,N_4785,N_4766);
xor U4860 (N_4860,N_4707,N_4788);
xor U4861 (N_4861,N_4727,N_4677);
xnor U4862 (N_4862,N_4781,N_4741);
xor U4863 (N_4863,N_4743,N_4794);
or U4864 (N_4864,N_4783,N_4753);
xnor U4865 (N_4865,N_4676,N_4737);
or U4866 (N_4866,N_4714,N_4703);
nand U4867 (N_4867,N_4694,N_4687);
nor U4868 (N_4868,N_4745,N_4718);
xnor U4869 (N_4869,N_4759,N_4733);
nor U4870 (N_4870,N_4778,N_4734);
nor U4871 (N_4871,N_4763,N_4780);
or U4872 (N_4872,N_4771,N_4690);
xnor U4873 (N_4873,N_4791,N_4688);
nor U4874 (N_4874,N_4651,N_4715);
or U4875 (N_4875,N_4742,N_4664);
or U4876 (N_4876,N_4749,N_4728);
or U4877 (N_4877,N_4791,N_4709);
xor U4878 (N_4878,N_4741,N_4753);
and U4879 (N_4879,N_4724,N_4695);
or U4880 (N_4880,N_4785,N_4790);
and U4881 (N_4881,N_4660,N_4776);
nand U4882 (N_4882,N_4693,N_4691);
and U4883 (N_4883,N_4748,N_4678);
xnor U4884 (N_4884,N_4663,N_4692);
nand U4885 (N_4885,N_4720,N_4686);
nor U4886 (N_4886,N_4688,N_4798);
nand U4887 (N_4887,N_4667,N_4758);
xor U4888 (N_4888,N_4685,N_4775);
or U4889 (N_4889,N_4799,N_4687);
nand U4890 (N_4890,N_4751,N_4790);
nor U4891 (N_4891,N_4754,N_4746);
nand U4892 (N_4892,N_4672,N_4661);
or U4893 (N_4893,N_4650,N_4681);
or U4894 (N_4894,N_4743,N_4775);
xor U4895 (N_4895,N_4798,N_4772);
nand U4896 (N_4896,N_4747,N_4688);
or U4897 (N_4897,N_4739,N_4758);
xnor U4898 (N_4898,N_4675,N_4748);
and U4899 (N_4899,N_4676,N_4734);
nor U4900 (N_4900,N_4667,N_4665);
nor U4901 (N_4901,N_4766,N_4762);
or U4902 (N_4902,N_4659,N_4711);
and U4903 (N_4903,N_4697,N_4735);
and U4904 (N_4904,N_4669,N_4771);
and U4905 (N_4905,N_4722,N_4673);
nand U4906 (N_4906,N_4759,N_4763);
or U4907 (N_4907,N_4685,N_4707);
xor U4908 (N_4908,N_4656,N_4686);
nor U4909 (N_4909,N_4715,N_4747);
xor U4910 (N_4910,N_4753,N_4797);
and U4911 (N_4911,N_4798,N_4789);
and U4912 (N_4912,N_4780,N_4752);
xor U4913 (N_4913,N_4704,N_4756);
nand U4914 (N_4914,N_4684,N_4769);
or U4915 (N_4915,N_4799,N_4710);
nor U4916 (N_4916,N_4718,N_4794);
nor U4917 (N_4917,N_4774,N_4759);
nand U4918 (N_4918,N_4728,N_4676);
or U4919 (N_4919,N_4721,N_4798);
or U4920 (N_4920,N_4651,N_4709);
xnor U4921 (N_4921,N_4770,N_4695);
or U4922 (N_4922,N_4672,N_4758);
and U4923 (N_4923,N_4670,N_4685);
nand U4924 (N_4924,N_4717,N_4765);
nor U4925 (N_4925,N_4712,N_4710);
nor U4926 (N_4926,N_4718,N_4652);
nand U4927 (N_4927,N_4778,N_4762);
xor U4928 (N_4928,N_4651,N_4670);
and U4929 (N_4929,N_4775,N_4732);
or U4930 (N_4930,N_4655,N_4726);
nand U4931 (N_4931,N_4667,N_4722);
or U4932 (N_4932,N_4685,N_4692);
xnor U4933 (N_4933,N_4705,N_4760);
and U4934 (N_4934,N_4680,N_4790);
nor U4935 (N_4935,N_4746,N_4795);
or U4936 (N_4936,N_4705,N_4672);
xor U4937 (N_4937,N_4775,N_4653);
nor U4938 (N_4938,N_4700,N_4662);
and U4939 (N_4939,N_4784,N_4787);
nor U4940 (N_4940,N_4764,N_4771);
nand U4941 (N_4941,N_4651,N_4736);
or U4942 (N_4942,N_4720,N_4703);
and U4943 (N_4943,N_4739,N_4771);
nand U4944 (N_4944,N_4650,N_4686);
nor U4945 (N_4945,N_4771,N_4782);
and U4946 (N_4946,N_4798,N_4658);
and U4947 (N_4947,N_4722,N_4654);
or U4948 (N_4948,N_4756,N_4672);
or U4949 (N_4949,N_4795,N_4790);
nand U4950 (N_4950,N_4856,N_4928);
nor U4951 (N_4951,N_4801,N_4811);
or U4952 (N_4952,N_4879,N_4855);
nor U4953 (N_4953,N_4890,N_4825);
nand U4954 (N_4954,N_4866,N_4867);
xnor U4955 (N_4955,N_4892,N_4816);
or U4956 (N_4956,N_4819,N_4891);
and U4957 (N_4957,N_4836,N_4909);
nand U4958 (N_4958,N_4925,N_4818);
xnor U4959 (N_4959,N_4804,N_4846);
or U4960 (N_4960,N_4913,N_4812);
nor U4961 (N_4961,N_4832,N_4884);
or U4962 (N_4962,N_4908,N_4802);
nand U4963 (N_4963,N_4937,N_4901);
nand U4964 (N_4964,N_4865,N_4841);
nor U4965 (N_4965,N_4949,N_4868);
and U4966 (N_4966,N_4839,N_4848);
and U4967 (N_4967,N_4806,N_4876);
or U4968 (N_4968,N_4851,N_4934);
xnor U4969 (N_4969,N_4916,N_4822);
or U4970 (N_4970,N_4809,N_4906);
nor U4971 (N_4971,N_4922,N_4911);
nor U4972 (N_4972,N_4942,N_4894);
and U4973 (N_4973,N_4902,N_4852);
nand U4974 (N_4974,N_4864,N_4877);
nand U4975 (N_4975,N_4920,N_4803);
and U4976 (N_4976,N_4943,N_4895);
or U4977 (N_4977,N_4835,N_4826);
or U4978 (N_4978,N_4938,N_4853);
nor U4979 (N_4979,N_4907,N_4815);
xor U4980 (N_4980,N_4861,N_4845);
or U4981 (N_4981,N_4823,N_4843);
xor U4982 (N_4982,N_4842,N_4810);
nand U4983 (N_4983,N_4946,N_4905);
nand U4984 (N_4984,N_4824,N_4880);
nor U4985 (N_4985,N_4927,N_4808);
and U4986 (N_4986,N_4947,N_4899);
nand U4987 (N_4987,N_4833,N_4838);
nor U4988 (N_4988,N_4917,N_4933);
xnor U4989 (N_4989,N_4805,N_4870);
nor U4990 (N_4990,N_4896,N_4932);
xor U4991 (N_4991,N_4923,N_4872);
and U4992 (N_4992,N_4807,N_4948);
nor U4993 (N_4993,N_4926,N_4915);
and U4994 (N_4994,N_4924,N_4886);
xnor U4995 (N_4995,N_4830,N_4914);
and U4996 (N_4996,N_4887,N_4847);
xnor U4997 (N_4997,N_4827,N_4945);
nand U4998 (N_4998,N_4828,N_4912);
or U4999 (N_4999,N_4854,N_4903);
nor U5000 (N_5000,N_4800,N_4820);
or U5001 (N_5001,N_4939,N_4871);
or U5002 (N_5002,N_4910,N_4834);
nand U5003 (N_5003,N_4936,N_4859);
xor U5004 (N_5004,N_4878,N_4889);
xnor U5005 (N_5005,N_4900,N_4849);
nor U5006 (N_5006,N_4875,N_4857);
or U5007 (N_5007,N_4940,N_4850);
nor U5008 (N_5008,N_4930,N_4941);
or U5009 (N_5009,N_4919,N_4874);
and U5010 (N_5010,N_4931,N_4893);
or U5011 (N_5011,N_4882,N_4829);
xnor U5012 (N_5012,N_4935,N_4904);
and U5013 (N_5013,N_4821,N_4898);
xnor U5014 (N_5014,N_4831,N_4814);
nand U5015 (N_5015,N_4862,N_4929);
and U5016 (N_5016,N_4837,N_4944);
nand U5017 (N_5017,N_4918,N_4897);
nor U5018 (N_5018,N_4817,N_4885);
and U5019 (N_5019,N_4863,N_4921);
xnor U5020 (N_5020,N_4860,N_4888);
xor U5021 (N_5021,N_4858,N_4881);
or U5022 (N_5022,N_4873,N_4844);
or U5023 (N_5023,N_4813,N_4840);
or U5024 (N_5024,N_4869,N_4883);
nor U5025 (N_5025,N_4889,N_4860);
nor U5026 (N_5026,N_4811,N_4828);
xor U5027 (N_5027,N_4800,N_4847);
and U5028 (N_5028,N_4840,N_4876);
nor U5029 (N_5029,N_4892,N_4801);
nand U5030 (N_5030,N_4888,N_4917);
or U5031 (N_5031,N_4835,N_4814);
nor U5032 (N_5032,N_4895,N_4870);
nand U5033 (N_5033,N_4840,N_4890);
nor U5034 (N_5034,N_4856,N_4946);
or U5035 (N_5035,N_4833,N_4824);
nor U5036 (N_5036,N_4886,N_4881);
nand U5037 (N_5037,N_4909,N_4888);
and U5038 (N_5038,N_4805,N_4827);
xnor U5039 (N_5039,N_4911,N_4801);
and U5040 (N_5040,N_4942,N_4860);
xor U5041 (N_5041,N_4909,N_4819);
nand U5042 (N_5042,N_4866,N_4850);
nor U5043 (N_5043,N_4876,N_4800);
and U5044 (N_5044,N_4846,N_4819);
nand U5045 (N_5045,N_4936,N_4916);
xnor U5046 (N_5046,N_4824,N_4832);
and U5047 (N_5047,N_4932,N_4803);
nand U5048 (N_5048,N_4843,N_4947);
or U5049 (N_5049,N_4855,N_4915);
and U5050 (N_5050,N_4831,N_4806);
nand U5051 (N_5051,N_4843,N_4902);
nor U5052 (N_5052,N_4829,N_4923);
xor U5053 (N_5053,N_4874,N_4903);
and U5054 (N_5054,N_4931,N_4867);
nor U5055 (N_5055,N_4922,N_4910);
nand U5056 (N_5056,N_4935,N_4808);
and U5057 (N_5057,N_4887,N_4802);
xor U5058 (N_5058,N_4867,N_4923);
nand U5059 (N_5059,N_4850,N_4878);
and U5060 (N_5060,N_4861,N_4827);
nor U5061 (N_5061,N_4864,N_4930);
xor U5062 (N_5062,N_4823,N_4880);
xor U5063 (N_5063,N_4930,N_4870);
and U5064 (N_5064,N_4926,N_4878);
nand U5065 (N_5065,N_4941,N_4846);
or U5066 (N_5066,N_4907,N_4900);
and U5067 (N_5067,N_4828,N_4829);
and U5068 (N_5068,N_4844,N_4917);
and U5069 (N_5069,N_4802,N_4807);
and U5070 (N_5070,N_4877,N_4806);
nor U5071 (N_5071,N_4827,N_4902);
nor U5072 (N_5072,N_4937,N_4823);
xnor U5073 (N_5073,N_4829,N_4821);
nor U5074 (N_5074,N_4867,N_4821);
nand U5075 (N_5075,N_4946,N_4911);
or U5076 (N_5076,N_4834,N_4866);
or U5077 (N_5077,N_4848,N_4878);
nand U5078 (N_5078,N_4888,N_4889);
or U5079 (N_5079,N_4857,N_4841);
nand U5080 (N_5080,N_4871,N_4899);
nand U5081 (N_5081,N_4926,N_4881);
nand U5082 (N_5082,N_4911,N_4818);
nand U5083 (N_5083,N_4916,N_4805);
nor U5084 (N_5084,N_4868,N_4885);
nor U5085 (N_5085,N_4944,N_4926);
nand U5086 (N_5086,N_4827,N_4877);
and U5087 (N_5087,N_4800,N_4865);
or U5088 (N_5088,N_4908,N_4846);
or U5089 (N_5089,N_4916,N_4918);
xor U5090 (N_5090,N_4941,N_4898);
and U5091 (N_5091,N_4827,N_4925);
nor U5092 (N_5092,N_4890,N_4888);
and U5093 (N_5093,N_4907,N_4924);
xor U5094 (N_5094,N_4881,N_4872);
and U5095 (N_5095,N_4903,N_4922);
xnor U5096 (N_5096,N_4940,N_4885);
nor U5097 (N_5097,N_4870,N_4857);
and U5098 (N_5098,N_4860,N_4920);
xor U5099 (N_5099,N_4847,N_4811);
nor U5100 (N_5100,N_5057,N_5086);
xnor U5101 (N_5101,N_4956,N_5073);
nor U5102 (N_5102,N_5046,N_5031);
xnor U5103 (N_5103,N_5095,N_5002);
or U5104 (N_5104,N_5028,N_5085);
or U5105 (N_5105,N_5033,N_5014);
or U5106 (N_5106,N_4991,N_4980);
or U5107 (N_5107,N_5022,N_5065);
and U5108 (N_5108,N_4986,N_5000);
and U5109 (N_5109,N_5071,N_5048);
xnor U5110 (N_5110,N_5015,N_5008);
nand U5111 (N_5111,N_5062,N_5081);
nand U5112 (N_5112,N_4978,N_5012);
nor U5113 (N_5113,N_4969,N_5027);
xnor U5114 (N_5114,N_5091,N_5013);
xnor U5115 (N_5115,N_4985,N_5049);
and U5116 (N_5116,N_4981,N_5068);
nand U5117 (N_5117,N_5041,N_5037);
and U5118 (N_5118,N_4995,N_4998);
nand U5119 (N_5119,N_5026,N_5098);
nor U5120 (N_5120,N_4999,N_4962);
xnor U5121 (N_5121,N_4987,N_5070);
nor U5122 (N_5122,N_5058,N_4990);
xnor U5123 (N_5123,N_4957,N_5003);
nand U5124 (N_5124,N_5030,N_5069);
xnor U5125 (N_5125,N_5010,N_4958);
or U5126 (N_5126,N_5061,N_5084);
or U5127 (N_5127,N_4963,N_5004);
xnor U5128 (N_5128,N_5052,N_4970);
nand U5129 (N_5129,N_5076,N_5089);
and U5130 (N_5130,N_4952,N_5087);
and U5131 (N_5131,N_5017,N_5016);
nand U5132 (N_5132,N_5066,N_5045);
xnor U5133 (N_5133,N_5019,N_5042);
or U5134 (N_5134,N_5064,N_4984);
nand U5135 (N_5135,N_4951,N_4993);
and U5136 (N_5136,N_5001,N_5036);
nor U5137 (N_5137,N_5054,N_5078);
xor U5138 (N_5138,N_5043,N_5025);
nand U5139 (N_5139,N_4977,N_4953);
nor U5140 (N_5140,N_5051,N_5032);
nor U5141 (N_5141,N_5063,N_5093);
xnor U5142 (N_5142,N_5006,N_5082);
xnor U5143 (N_5143,N_5074,N_5092);
nor U5144 (N_5144,N_5040,N_5060);
or U5145 (N_5145,N_4996,N_5007);
and U5146 (N_5146,N_4997,N_5088);
or U5147 (N_5147,N_5009,N_4973);
or U5148 (N_5148,N_4988,N_4975);
and U5149 (N_5149,N_5023,N_5035);
nand U5150 (N_5150,N_5056,N_4964);
or U5151 (N_5151,N_5096,N_4971);
nand U5152 (N_5152,N_4960,N_4966);
or U5153 (N_5153,N_5021,N_5047);
xnor U5154 (N_5154,N_5038,N_5083);
nand U5155 (N_5155,N_4965,N_4982);
nor U5156 (N_5156,N_5050,N_4954);
nor U5157 (N_5157,N_5055,N_4979);
and U5158 (N_5158,N_5079,N_4992);
xnor U5159 (N_5159,N_5097,N_5080);
and U5160 (N_5160,N_4983,N_5029);
nand U5161 (N_5161,N_4989,N_4994);
and U5162 (N_5162,N_5053,N_4974);
nor U5163 (N_5163,N_5075,N_5072);
xnor U5164 (N_5164,N_4961,N_5077);
or U5165 (N_5165,N_5024,N_5059);
or U5166 (N_5166,N_5005,N_5090);
or U5167 (N_5167,N_4976,N_4967);
xor U5168 (N_5168,N_5034,N_4972);
nor U5169 (N_5169,N_5018,N_5011);
nor U5170 (N_5170,N_5067,N_5094);
or U5171 (N_5171,N_4950,N_5099);
and U5172 (N_5172,N_5044,N_5039);
xor U5173 (N_5173,N_4968,N_4959);
or U5174 (N_5174,N_4955,N_5020);
nand U5175 (N_5175,N_4996,N_5097);
nand U5176 (N_5176,N_4982,N_5062);
nand U5177 (N_5177,N_5016,N_4977);
and U5178 (N_5178,N_4989,N_5049);
xor U5179 (N_5179,N_4987,N_5018);
xor U5180 (N_5180,N_4996,N_5038);
or U5181 (N_5181,N_4961,N_4983);
xor U5182 (N_5182,N_5048,N_5051);
and U5183 (N_5183,N_5072,N_5004);
nand U5184 (N_5184,N_4993,N_4952);
xor U5185 (N_5185,N_5046,N_4952);
or U5186 (N_5186,N_5049,N_4972);
and U5187 (N_5187,N_5000,N_5032);
xor U5188 (N_5188,N_5093,N_5091);
nand U5189 (N_5189,N_4979,N_4964);
or U5190 (N_5190,N_5036,N_4994);
and U5191 (N_5191,N_4970,N_5027);
or U5192 (N_5192,N_5075,N_4989);
nor U5193 (N_5193,N_5026,N_5083);
nand U5194 (N_5194,N_5003,N_5079);
nand U5195 (N_5195,N_5013,N_5089);
xnor U5196 (N_5196,N_5063,N_4984);
xnor U5197 (N_5197,N_5057,N_5076);
nand U5198 (N_5198,N_4980,N_4990);
nor U5199 (N_5199,N_4956,N_4982);
or U5200 (N_5200,N_5014,N_5023);
nand U5201 (N_5201,N_4993,N_4956);
nand U5202 (N_5202,N_4956,N_4978);
nor U5203 (N_5203,N_5031,N_4967);
xor U5204 (N_5204,N_5050,N_5094);
and U5205 (N_5205,N_4974,N_5050);
nor U5206 (N_5206,N_5048,N_5099);
or U5207 (N_5207,N_4972,N_4983);
xor U5208 (N_5208,N_5082,N_5051);
nor U5209 (N_5209,N_4981,N_5057);
nand U5210 (N_5210,N_4955,N_5025);
nor U5211 (N_5211,N_5070,N_5026);
nor U5212 (N_5212,N_4993,N_4990);
nand U5213 (N_5213,N_5039,N_5001);
nand U5214 (N_5214,N_5095,N_5077);
xnor U5215 (N_5215,N_5093,N_4977);
nor U5216 (N_5216,N_4985,N_5072);
or U5217 (N_5217,N_5008,N_4985);
nor U5218 (N_5218,N_5015,N_5007);
and U5219 (N_5219,N_5050,N_5079);
nand U5220 (N_5220,N_5032,N_4993);
xor U5221 (N_5221,N_5053,N_5045);
nor U5222 (N_5222,N_4994,N_5050);
nor U5223 (N_5223,N_4986,N_4994);
xor U5224 (N_5224,N_4996,N_4954);
or U5225 (N_5225,N_5022,N_4978);
nand U5226 (N_5226,N_5065,N_5066);
or U5227 (N_5227,N_4971,N_5064);
xor U5228 (N_5228,N_5063,N_4983);
xor U5229 (N_5229,N_5003,N_5045);
nand U5230 (N_5230,N_4988,N_5035);
and U5231 (N_5231,N_5053,N_4953);
nor U5232 (N_5232,N_5088,N_4952);
and U5233 (N_5233,N_5033,N_5032);
or U5234 (N_5234,N_5017,N_5066);
and U5235 (N_5235,N_5030,N_5005);
or U5236 (N_5236,N_4958,N_5086);
nor U5237 (N_5237,N_4995,N_5009);
nor U5238 (N_5238,N_5088,N_5095);
nor U5239 (N_5239,N_5084,N_5034);
xnor U5240 (N_5240,N_5093,N_5066);
nand U5241 (N_5241,N_4953,N_5096);
or U5242 (N_5242,N_5044,N_5005);
nor U5243 (N_5243,N_4963,N_5013);
nor U5244 (N_5244,N_5075,N_5042);
xor U5245 (N_5245,N_4969,N_4991);
nor U5246 (N_5246,N_5032,N_5063);
or U5247 (N_5247,N_5016,N_5004);
or U5248 (N_5248,N_5095,N_4987);
and U5249 (N_5249,N_5081,N_5072);
xor U5250 (N_5250,N_5212,N_5124);
nor U5251 (N_5251,N_5171,N_5128);
or U5252 (N_5252,N_5168,N_5110);
or U5253 (N_5253,N_5177,N_5213);
or U5254 (N_5254,N_5162,N_5237);
and U5255 (N_5255,N_5132,N_5148);
and U5256 (N_5256,N_5192,N_5102);
xnor U5257 (N_5257,N_5127,N_5143);
nor U5258 (N_5258,N_5231,N_5101);
xnor U5259 (N_5259,N_5178,N_5214);
nor U5260 (N_5260,N_5129,N_5244);
xnor U5261 (N_5261,N_5205,N_5123);
nand U5262 (N_5262,N_5133,N_5156);
nor U5263 (N_5263,N_5183,N_5152);
nor U5264 (N_5264,N_5140,N_5235);
and U5265 (N_5265,N_5160,N_5202);
nor U5266 (N_5266,N_5200,N_5158);
or U5267 (N_5267,N_5193,N_5220);
and U5268 (N_5268,N_5245,N_5209);
xnor U5269 (N_5269,N_5240,N_5204);
xnor U5270 (N_5270,N_5180,N_5189);
nor U5271 (N_5271,N_5163,N_5232);
nand U5272 (N_5272,N_5243,N_5219);
or U5273 (N_5273,N_5223,N_5185);
and U5274 (N_5274,N_5149,N_5221);
xnor U5275 (N_5275,N_5225,N_5198);
xnor U5276 (N_5276,N_5138,N_5142);
and U5277 (N_5277,N_5109,N_5119);
nor U5278 (N_5278,N_5179,N_5181);
nor U5279 (N_5279,N_5236,N_5208);
nor U5280 (N_5280,N_5117,N_5186);
nand U5281 (N_5281,N_5106,N_5233);
xor U5282 (N_5282,N_5136,N_5118);
or U5283 (N_5283,N_5157,N_5218);
or U5284 (N_5284,N_5104,N_5206);
or U5285 (N_5285,N_5176,N_5141);
or U5286 (N_5286,N_5131,N_5216);
or U5287 (N_5287,N_5125,N_5215);
xnor U5288 (N_5288,N_5120,N_5190);
and U5289 (N_5289,N_5210,N_5151);
or U5290 (N_5290,N_5108,N_5172);
xnor U5291 (N_5291,N_5197,N_5153);
nand U5292 (N_5292,N_5130,N_5227);
xor U5293 (N_5293,N_5241,N_5154);
nand U5294 (N_5294,N_5234,N_5196);
and U5295 (N_5295,N_5173,N_5112);
xor U5296 (N_5296,N_5116,N_5126);
nand U5297 (N_5297,N_5147,N_5228);
nor U5298 (N_5298,N_5195,N_5246);
nor U5299 (N_5299,N_5159,N_5230);
nand U5300 (N_5300,N_5155,N_5242);
xor U5301 (N_5301,N_5207,N_5164);
or U5302 (N_5302,N_5199,N_5201);
xor U5303 (N_5303,N_5146,N_5134);
nand U5304 (N_5304,N_5174,N_5184);
or U5305 (N_5305,N_5239,N_5107);
nor U5306 (N_5306,N_5248,N_5139);
nor U5307 (N_5307,N_5222,N_5111);
xnor U5308 (N_5308,N_5144,N_5249);
xnor U5309 (N_5309,N_5166,N_5114);
xor U5310 (N_5310,N_5238,N_5145);
or U5311 (N_5311,N_5150,N_5105);
xor U5312 (N_5312,N_5113,N_5100);
nor U5313 (N_5313,N_5175,N_5224);
xnor U5314 (N_5314,N_5135,N_5122);
or U5315 (N_5315,N_5188,N_5121);
nand U5316 (N_5316,N_5229,N_5226);
xnor U5317 (N_5317,N_5194,N_5217);
and U5318 (N_5318,N_5103,N_5167);
xnor U5319 (N_5319,N_5191,N_5203);
xnor U5320 (N_5320,N_5247,N_5170);
and U5321 (N_5321,N_5169,N_5182);
and U5322 (N_5322,N_5211,N_5165);
nor U5323 (N_5323,N_5137,N_5187);
nand U5324 (N_5324,N_5161,N_5115);
nor U5325 (N_5325,N_5101,N_5141);
and U5326 (N_5326,N_5108,N_5170);
nor U5327 (N_5327,N_5226,N_5194);
nand U5328 (N_5328,N_5217,N_5116);
and U5329 (N_5329,N_5161,N_5204);
xnor U5330 (N_5330,N_5119,N_5175);
and U5331 (N_5331,N_5141,N_5218);
nand U5332 (N_5332,N_5178,N_5174);
nor U5333 (N_5333,N_5107,N_5180);
or U5334 (N_5334,N_5124,N_5205);
or U5335 (N_5335,N_5177,N_5236);
xor U5336 (N_5336,N_5228,N_5166);
xor U5337 (N_5337,N_5152,N_5121);
nand U5338 (N_5338,N_5233,N_5100);
and U5339 (N_5339,N_5145,N_5101);
and U5340 (N_5340,N_5157,N_5168);
or U5341 (N_5341,N_5200,N_5234);
nor U5342 (N_5342,N_5211,N_5238);
nand U5343 (N_5343,N_5210,N_5248);
or U5344 (N_5344,N_5180,N_5235);
and U5345 (N_5345,N_5222,N_5188);
nand U5346 (N_5346,N_5224,N_5117);
nand U5347 (N_5347,N_5140,N_5110);
nor U5348 (N_5348,N_5102,N_5148);
xor U5349 (N_5349,N_5241,N_5120);
and U5350 (N_5350,N_5217,N_5165);
and U5351 (N_5351,N_5103,N_5119);
and U5352 (N_5352,N_5243,N_5111);
nor U5353 (N_5353,N_5212,N_5116);
nor U5354 (N_5354,N_5139,N_5132);
or U5355 (N_5355,N_5215,N_5247);
xnor U5356 (N_5356,N_5238,N_5248);
or U5357 (N_5357,N_5198,N_5197);
nand U5358 (N_5358,N_5156,N_5130);
xnor U5359 (N_5359,N_5200,N_5173);
nand U5360 (N_5360,N_5134,N_5109);
xor U5361 (N_5361,N_5248,N_5224);
and U5362 (N_5362,N_5142,N_5131);
or U5363 (N_5363,N_5129,N_5109);
nor U5364 (N_5364,N_5198,N_5247);
and U5365 (N_5365,N_5174,N_5239);
nor U5366 (N_5366,N_5175,N_5187);
nand U5367 (N_5367,N_5128,N_5131);
nand U5368 (N_5368,N_5124,N_5155);
xnor U5369 (N_5369,N_5185,N_5199);
nand U5370 (N_5370,N_5134,N_5181);
or U5371 (N_5371,N_5148,N_5209);
xor U5372 (N_5372,N_5231,N_5202);
nor U5373 (N_5373,N_5132,N_5202);
and U5374 (N_5374,N_5148,N_5115);
and U5375 (N_5375,N_5200,N_5122);
and U5376 (N_5376,N_5205,N_5189);
nor U5377 (N_5377,N_5128,N_5210);
nor U5378 (N_5378,N_5153,N_5135);
nor U5379 (N_5379,N_5242,N_5141);
or U5380 (N_5380,N_5183,N_5232);
nor U5381 (N_5381,N_5217,N_5189);
and U5382 (N_5382,N_5215,N_5101);
nand U5383 (N_5383,N_5123,N_5140);
xnor U5384 (N_5384,N_5240,N_5156);
nor U5385 (N_5385,N_5158,N_5214);
xnor U5386 (N_5386,N_5222,N_5226);
xor U5387 (N_5387,N_5185,N_5135);
nor U5388 (N_5388,N_5190,N_5155);
xnor U5389 (N_5389,N_5164,N_5212);
or U5390 (N_5390,N_5241,N_5150);
nand U5391 (N_5391,N_5195,N_5211);
nand U5392 (N_5392,N_5104,N_5189);
and U5393 (N_5393,N_5111,N_5152);
xnor U5394 (N_5394,N_5139,N_5142);
xnor U5395 (N_5395,N_5232,N_5119);
xor U5396 (N_5396,N_5110,N_5177);
nand U5397 (N_5397,N_5118,N_5230);
and U5398 (N_5398,N_5249,N_5216);
and U5399 (N_5399,N_5236,N_5187);
nand U5400 (N_5400,N_5360,N_5277);
and U5401 (N_5401,N_5280,N_5347);
nor U5402 (N_5402,N_5257,N_5274);
nor U5403 (N_5403,N_5252,N_5379);
nand U5404 (N_5404,N_5363,N_5265);
xnor U5405 (N_5405,N_5342,N_5326);
nor U5406 (N_5406,N_5377,N_5325);
nand U5407 (N_5407,N_5275,N_5298);
or U5408 (N_5408,N_5368,N_5260);
or U5409 (N_5409,N_5317,N_5345);
nand U5410 (N_5410,N_5375,N_5307);
and U5411 (N_5411,N_5319,N_5308);
or U5412 (N_5412,N_5392,N_5315);
xnor U5413 (N_5413,N_5362,N_5352);
and U5414 (N_5414,N_5271,N_5267);
xor U5415 (N_5415,N_5297,N_5369);
and U5416 (N_5416,N_5339,N_5365);
nor U5417 (N_5417,N_5374,N_5370);
nand U5418 (N_5418,N_5394,N_5385);
nand U5419 (N_5419,N_5367,N_5301);
nand U5420 (N_5420,N_5259,N_5349);
xor U5421 (N_5421,N_5321,N_5388);
nor U5422 (N_5422,N_5398,N_5263);
nand U5423 (N_5423,N_5284,N_5333);
nand U5424 (N_5424,N_5337,N_5296);
nor U5425 (N_5425,N_5285,N_5390);
or U5426 (N_5426,N_5381,N_5350);
nor U5427 (N_5427,N_5380,N_5310);
xor U5428 (N_5428,N_5251,N_5387);
and U5429 (N_5429,N_5292,N_5395);
and U5430 (N_5430,N_5279,N_5356);
and U5431 (N_5431,N_5290,N_5331);
xnor U5432 (N_5432,N_5357,N_5261);
or U5433 (N_5433,N_5266,N_5338);
nor U5434 (N_5434,N_5348,N_5295);
xor U5435 (N_5435,N_5322,N_5364);
nand U5436 (N_5436,N_5320,N_5330);
nand U5437 (N_5437,N_5335,N_5313);
nor U5438 (N_5438,N_5391,N_5373);
xnor U5439 (N_5439,N_5312,N_5359);
xor U5440 (N_5440,N_5316,N_5300);
nand U5441 (N_5441,N_5268,N_5289);
xnor U5442 (N_5442,N_5383,N_5272);
xnor U5443 (N_5443,N_5288,N_5334);
and U5444 (N_5444,N_5306,N_5318);
or U5445 (N_5445,N_5353,N_5329);
nor U5446 (N_5446,N_5305,N_5376);
nor U5447 (N_5447,N_5361,N_5250);
nor U5448 (N_5448,N_5314,N_5324);
nand U5449 (N_5449,N_5256,N_5327);
xor U5450 (N_5450,N_5382,N_5371);
xor U5451 (N_5451,N_5340,N_5293);
and U5452 (N_5452,N_5283,N_5343);
nor U5453 (N_5453,N_5273,N_5378);
and U5454 (N_5454,N_5386,N_5281);
xnor U5455 (N_5455,N_5393,N_5354);
xnor U5456 (N_5456,N_5355,N_5264);
and U5457 (N_5457,N_5346,N_5332);
xor U5458 (N_5458,N_5287,N_5328);
or U5459 (N_5459,N_5269,N_5384);
or U5460 (N_5460,N_5358,N_5309);
nor U5461 (N_5461,N_5372,N_5302);
nor U5462 (N_5462,N_5258,N_5304);
and U5463 (N_5463,N_5270,N_5299);
or U5464 (N_5464,N_5396,N_5303);
and U5465 (N_5465,N_5397,N_5351);
or U5466 (N_5466,N_5399,N_5253);
nand U5467 (N_5467,N_5389,N_5366);
and U5468 (N_5468,N_5341,N_5311);
nor U5469 (N_5469,N_5323,N_5254);
or U5470 (N_5470,N_5262,N_5294);
xnor U5471 (N_5471,N_5291,N_5344);
nand U5472 (N_5472,N_5255,N_5278);
nor U5473 (N_5473,N_5276,N_5286);
nor U5474 (N_5474,N_5336,N_5282);
nand U5475 (N_5475,N_5330,N_5322);
xnor U5476 (N_5476,N_5326,N_5334);
nor U5477 (N_5477,N_5302,N_5397);
or U5478 (N_5478,N_5329,N_5313);
and U5479 (N_5479,N_5283,N_5274);
nand U5480 (N_5480,N_5303,N_5275);
and U5481 (N_5481,N_5335,N_5348);
nand U5482 (N_5482,N_5271,N_5280);
xnor U5483 (N_5483,N_5384,N_5307);
or U5484 (N_5484,N_5321,N_5390);
nand U5485 (N_5485,N_5347,N_5313);
and U5486 (N_5486,N_5334,N_5317);
xor U5487 (N_5487,N_5250,N_5309);
xor U5488 (N_5488,N_5376,N_5382);
nand U5489 (N_5489,N_5330,N_5310);
xnor U5490 (N_5490,N_5314,N_5391);
nor U5491 (N_5491,N_5374,N_5303);
nand U5492 (N_5492,N_5359,N_5309);
nor U5493 (N_5493,N_5310,N_5268);
and U5494 (N_5494,N_5329,N_5310);
xor U5495 (N_5495,N_5383,N_5362);
and U5496 (N_5496,N_5277,N_5303);
xnor U5497 (N_5497,N_5284,N_5363);
nand U5498 (N_5498,N_5327,N_5322);
and U5499 (N_5499,N_5351,N_5307);
xor U5500 (N_5500,N_5276,N_5275);
and U5501 (N_5501,N_5297,N_5393);
xnor U5502 (N_5502,N_5347,N_5373);
or U5503 (N_5503,N_5332,N_5329);
and U5504 (N_5504,N_5334,N_5384);
and U5505 (N_5505,N_5279,N_5341);
nor U5506 (N_5506,N_5262,N_5355);
and U5507 (N_5507,N_5381,N_5364);
nand U5508 (N_5508,N_5291,N_5267);
nor U5509 (N_5509,N_5281,N_5371);
nor U5510 (N_5510,N_5356,N_5329);
nand U5511 (N_5511,N_5312,N_5295);
and U5512 (N_5512,N_5258,N_5331);
nand U5513 (N_5513,N_5356,N_5286);
nor U5514 (N_5514,N_5358,N_5366);
xnor U5515 (N_5515,N_5287,N_5329);
and U5516 (N_5516,N_5381,N_5292);
and U5517 (N_5517,N_5255,N_5285);
xor U5518 (N_5518,N_5384,N_5296);
and U5519 (N_5519,N_5324,N_5398);
xnor U5520 (N_5520,N_5263,N_5316);
nor U5521 (N_5521,N_5394,N_5291);
nand U5522 (N_5522,N_5311,N_5384);
nand U5523 (N_5523,N_5282,N_5314);
or U5524 (N_5524,N_5253,N_5347);
or U5525 (N_5525,N_5346,N_5308);
nor U5526 (N_5526,N_5399,N_5355);
xnor U5527 (N_5527,N_5375,N_5381);
nor U5528 (N_5528,N_5341,N_5355);
nand U5529 (N_5529,N_5277,N_5334);
nor U5530 (N_5530,N_5308,N_5379);
xnor U5531 (N_5531,N_5363,N_5256);
xnor U5532 (N_5532,N_5395,N_5282);
xor U5533 (N_5533,N_5345,N_5292);
nor U5534 (N_5534,N_5355,N_5256);
xor U5535 (N_5535,N_5335,N_5365);
and U5536 (N_5536,N_5301,N_5309);
or U5537 (N_5537,N_5311,N_5294);
xnor U5538 (N_5538,N_5386,N_5374);
nor U5539 (N_5539,N_5305,N_5337);
nand U5540 (N_5540,N_5327,N_5354);
or U5541 (N_5541,N_5386,N_5262);
and U5542 (N_5542,N_5339,N_5337);
nor U5543 (N_5543,N_5362,N_5283);
and U5544 (N_5544,N_5273,N_5262);
and U5545 (N_5545,N_5321,N_5359);
and U5546 (N_5546,N_5312,N_5315);
or U5547 (N_5547,N_5305,N_5385);
nand U5548 (N_5548,N_5389,N_5378);
or U5549 (N_5549,N_5279,N_5314);
nor U5550 (N_5550,N_5437,N_5466);
and U5551 (N_5551,N_5473,N_5538);
xnor U5552 (N_5552,N_5463,N_5404);
or U5553 (N_5553,N_5488,N_5403);
and U5554 (N_5554,N_5533,N_5494);
nand U5555 (N_5555,N_5441,N_5534);
and U5556 (N_5556,N_5448,N_5483);
or U5557 (N_5557,N_5467,N_5496);
nor U5558 (N_5558,N_5450,N_5407);
nor U5559 (N_5559,N_5435,N_5423);
xnor U5560 (N_5560,N_5472,N_5515);
or U5561 (N_5561,N_5523,N_5478);
xor U5562 (N_5562,N_5491,N_5481);
nor U5563 (N_5563,N_5546,N_5456);
nor U5564 (N_5564,N_5465,N_5477);
xnor U5565 (N_5565,N_5532,N_5504);
and U5566 (N_5566,N_5421,N_5508);
nand U5567 (N_5567,N_5531,N_5486);
or U5568 (N_5568,N_5543,N_5503);
xor U5569 (N_5569,N_5417,N_5425);
nand U5570 (N_5570,N_5443,N_5544);
nor U5571 (N_5571,N_5479,N_5433);
nand U5572 (N_5572,N_5452,N_5459);
or U5573 (N_5573,N_5514,N_5402);
and U5574 (N_5574,N_5414,N_5436);
nand U5575 (N_5575,N_5492,N_5445);
nand U5576 (N_5576,N_5470,N_5411);
and U5577 (N_5577,N_5429,N_5424);
nand U5578 (N_5578,N_5545,N_5539);
xor U5579 (N_5579,N_5455,N_5548);
or U5580 (N_5580,N_5406,N_5462);
xor U5581 (N_5581,N_5487,N_5529);
nand U5582 (N_5582,N_5474,N_5446);
and U5583 (N_5583,N_5464,N_5528);
nor U5584 (N_5584,N_5426,N_5519);
nand U5585 (N_5585,N_5507,N_5428);
nor U5586 (N_5586,N_5536,N_5432);
and U5587 (N_5587,N_5499,N_5449);
nor U5588 (N_5588,N_5468,N_5542);
and U5589 (N_5589,N_5495,N_5430);
or U5590 (N_5590,N_5439,N_5442);
xnor U5591 (N_5591,N_5475,N_5454);
or U5592 (N_5592,N_5530,N_5410);
and U5593 (N_5593,N_5513,N_5458);
or U5594 (N_5594,N_5505,N_5438);
xnor U5595 (N_5595,N_5447,N_5490);
nor U5596 (N_5596,N_5549,N_5511);
xnor U5597 (N_5597,N_5489,N_5516);
and U5598 (N_5598,N_5512,N_5498);
xnor U5599 (N_5599,N_5484,N_5510);
nor U5600 (N_5600,N_5521,N_5501);
or U5601 (N_5601,N_5418,N_5416);
nand U5602 (N_5602,N_5485,N_5413);
nor U5603 (N_5603,N_5527,N_5440);
nand U5604 (N_5604,N_5405,N_5453);
or U5605 (N_5605,N_5524,N_5427);
nand U5606 (N_5606,N_5420,N_5412);
xor U5607 (N_5607,N_5408,N_5517);
xor U5608 (N_5608,N_5506,N_5422);
and U5609 (N_5609,N_5482,N_5415);
xnor U5610 (N_5610,N_5526,N_5502);
xor U5611 (N_5611,N_5500,N_5457);
and U5612 (N_5612,N_5431,N_5535);
xor U5613 (N_5613,N_5541,N_5419);
or U5614 (N_5614,N_5497,N_5522);
nor U5615 (N_5615,N_5476,N_5537);
xnor U5616 (N_5616,N_5461,N_5520);
xor U5617 (N_5617,N_5434,N_5471);
xor U5618 (N_5618,N_5480,N_5401);
or U5619 (N_5619,N_5493,N_5509);
and U5620 (N_5620,N_5525,N_5547);
nand U5621 (N_5621,N_5444,N_5451);
nor U5622 (N_5622,N_5518,N_5409);
or U5623 (N_5623,N_5540,N_5400);
xor U5624 (N_5624,N_5460,N_5469);
nor U5625 (N_5625,N_5489,N_5453);
nor U5626 (N_5626,N_5493,N_5534);
nand U5627 (N_5627,N_5431,N_5450);
nand U5628 (N_5628,N_5482,N_5525);
nor U5629 (N_5629,N_5453,N_5488);
nor U5630 (N_5630,N_5523,N_5423);
nor U5631 (N_5631,N_5501,N_5405);
or U5632 (N_5632,N_5418,N_5536);
or U5633 (N_5633,N_5525,N_5533);
xnor U5634 (N_5634,N_5428,N_5452);
nor U5635 (N_5635,N_5529,N_5419);
nor U5636 (N_5636,N_5402,N_5422);
xnor U5637 (N_5637,N_5438,N_5428);
or U5638 (N_5638,N_5420,N_5531);
and U5639 (N_5639,N_5479,N_5432);
xor U5640 (N_5640,N_5426,N_5548);
or U5641 (N_5641,N_5491,N_5409);
and U5642 (N_5642,N_5510,N_5453);
or U5643 (N_5643,N_5400,N_5476);
or U5644 (N_5644,N_5460,N_5498);
or U5645 (N_5645,N_5489,N_5519);
nand U5646 (N_5646,N_5518,N_5525);
nor U5647 (N_5647,N_5450,N_5457);
xnor U5648 (N_5648,N_5517,N_5412);
nand U5649 (N_5649,N_5416,N_5521);
xnor U5650 (N_5650,N_5516,N_5496);
and U5651 (N_5651,N_5457,N_5405);
and U5652 (N_5652,N_5496,N_5450);
and U5653 (N_5653,N_5494,N_5479);
or U5654 (N_5654,N_5489,N_5529);
nor U5655 (N_5655,N_5455,N_5494);
nor U5656 (N_5656,N_5456,N_5504);
or U5657 (N_5657,N_5494,N_5521);
or U5658 (N_5658,N_5482,N_5497);
nor U5659 (N_5659,N_5457,N_5432);
or U5660 (N_5660,N_5447,N_5403);
or U5661 (N_5661,N_5528,N_5439);
or U5662 (N_5662,N_5426,N_5503);
or U5663 (N_5663,N_5523,N_5437);
xnor U5664 (N_5664,N_5442,N_5487);
nor U5665 (N_5665,N_5484,N_5409);
nand U5666 (N_5666,N_5533,N_5429);
nand U5667 (N_5667,N_5486,N_5538);
nand U5668 (N_5668,N_5435,N_5496);
xnor U5669 (N_5669,N_5546,N_5537);
and U5670 (N_5670,N_5478,N_5504);
nor U5671 (N_5671,N_5500,N_5474);
xor U5672 (N_5672,N_5526,N_5491);
xnor U5673 (N_5673,N_5444,N_5463);
nand U5674 (N_5674,N_5457,N_5442);
nand U5675 (N_5675,N_5537,N_5512);
or U5676 (N_5676,N_5479,N_5482);
and U5677 (N_5677,N_5535,N_5428);
xor U5678 (N_5678,N_5467,N_5481);
xnor U5679 (N_5679,N_5402,N_5470);
and U5680 (N_5680,N_5416,N_5469);
or U5681 (N_5681,N_5469,N_5453);
or U5682 (N_5682,N_5429,N_5410);
nand U5683 (N_5683,N_5448,N_5415);
or U5684 (N_5684,N_5547,N_5414);
and U5685 (N_5685,N_5547,N_5458);
and U5686 (N_5686,N_5539,N_5497);
or U5687 (N_5687,N_5466,N_5443);
and U5688 (N_5688,N_5434,N_5451);
nand U5689 (N_5689,N_5450,N_5508);
xor U5690 (N_5690,N_5445,N_5436);
nand U5691 (N_5691,N_5518,N_5453);
nand U5692 (N_5692,N_5488,N_5497);
xnor U5693 (N_5693,N_5403,N_5542);
nand U5694 (N_5694,N_5446,N_5403);
or U5695 (N_5695,N_5417,N_5401);
nand U5696 (N_5696,N_5518,N_5490);
xnor U5697 (N_5697,N_5433,N_5473);
and U5698 (N_5698,N_5414,N_5543);
nand U5699 (N_5699,N_5464,N_5489);
and U5700 (N_5700,N_5578,N_5555);
or U5701 (N_5701,N_5554,N_5677);
xnor U5702 (N_5702,N_5600,N_5646);
or U5703 (N_5703,N_5568,N_5579);
and U5704 (N_5704,N_5607,N_5552);
nand U5705 (N_5705,N_5662,N_5585);
and U5706 (N_5706,N_5630,N_5699);
or U5707 (N_5707,N_5593,N_5691);
or U5708 (N_5708,N_5692,N_5594);
or U5709 (N_5709,N_5671,N_5654);
xnor U5710 (N_5710,N_5611,N_5694);
and U5711 (N_5711,N_5620,N_5678);
nor U5712 (N_5712,N_5584,N_5696);
nor U5713 (N_5713,N_5642,N_5637);
xor U5714 (N_5714,N_5697,N_5682);
nor U5715 (N_5715,N_5582,N_5626);
and U5716 (N_5716,N_5603,N_5580);
or U5717 (N_5717,N_5689,N_5641);
nor U5718 (N_5718,N_5669,N_5596);
xor U5719 (N_5719,N_5681,N_5668);
and U5720 (N_5720,N_5569,N_5665);
nor U5721 (N_5721,N_5683,N_5590);
nor U5722 (N_5722,N_5564,N_5638);
or U5723 (N_5723,N_5635,N_5602);
or U5724 (N_5724,N_5631,N_5676);
xor U5725 (N_5725,N_5623,N_5560);
nand U5726 (N_5726,N_5618,N_5670);
xnor U5727 (N_5727,N_5595,N_5601);
and U5728 (N_5728,N_5655,N_5667);
nor U5729 (N_5729,N_5647,N_5586);
nand U5730 (N_5730,N_5605,N_5556);
nand U5731 (N_5731,N_5653,N_5643);
nand U5732 (N_5732,N_5688,N_5656);
nand U5733 (N_5733,N_5616,N_5649);
xor U5734 (N_5734,N_5612,N_5551);
xor U5735 (N_5735,N_5587,N_5563);
or U5736 (N_5736,N_5561,N_5562);
and U5737 (N_5737,N_5648,N_5591);
nand U5738 (N_5738,N_5686,N_5621);
nor U5739 (N_5739,N_5666,N_5664);
nor U5740 (N_5740,N_5687,N_5644);
or U5741 (N_5741,N_5583,N_5599);
and U5742 (N_5742,N_5650,N_5588);
and U5743 (N_5743,N_5559,N_5627);
and U5744 (N_5744,N_5572,N_5615);
nand U5745 (N_5745,N_5619,N_5639);
and U5746 (N_5746,N_5625,N_5571);
nand U5747 (N_5747,N_5632,N_5592);
or U5748 (N_5748,N_5698,N_5633);
and U5749 (N_5749,N_5680,N_5660);
or U5750 (N_5750,N_5613,N_5684);
and U5751 (N_5751,N_5622,N_5659);
and U5752 (N_5752,N_5575,N_5617);
or U5753 (N_5753,N_5557,N_5679);
or U5754 (N_5754,N_5629,N_5651);
nor U5755 (N_5755,N_5652,N_5565);
nand U5756 (N_5756,N_5614,N_5553);
or U5757 (N_5757,N_5598,N_5674);
or U5758 (N_5758,N_5574,N_5550);
or U5759 (N_5759,N_5645,N_5695);
xor U5760 (N_5760,N_5690,N_5604);
xor U5761 (N_5761,N_5663,N_5581);
nor U5762 (N_5762,N_5606,N_5566);
or U5763 (N_5763,N_5577,N_5685);
and U5764 (N_5764,N_5610,N_5636);
xor U5765 (N_5765,N_5576,N_5570);
or U5766 (N_5766,N_5672,N_5634);
or U5767 (N_5767,N_5673,N_5567);
and U5768 (N_5768,N_5597,N_5628);
nor U5769 (N_5769,N_5608,N_5573);
nand U5770 (N_5770,N_5589,N_5640);
xnor U5771 (N_5771,N_5675,N_5658);
xnor U5772 (N_5772,N_5609,N_5558);
nand U5773 (N_5773,N_5657,N_5693);
xor U5774 (N_5774,N_5624,N_5661);
or U5775 (N_5775,N_5665,N_5597);
nand U5776 (N_5776,N_5645,N_5605);
xnor U5777 (N_5777,N_5625,N_5672);
and U5778 (N_5778,N_5614,N_5595);
xor U5779 (N_5779,N_5681,N_5655);
nor U5780 (N_5780,N_5654,N_5589);
xor U5781 (N_5781,N_5592,N_5583);
and U5782 (N_5782,N_5556,N_5581);
or U5783 (N_5783,N_5644,N_5573);
xor U5784 (N_5784,N_5614,N_5668);
nand U5785 (N_5785,N_5675,N_5649);
xor U5786 (N_5786,N_5688,N_5683);
or U5787 (N_5787,N_5590,N_5562);
nand U5788 (N_5788,N_5633,N_5686);
nand U5789 (N_5789,N_5586,N_5599);
nor U5790 (N_5790,N_5694,N_5691);
or U5791 (N_5791,N_5652,N_5646);
or U5792 (N_5792,N_5576,N_5670);
or U5793 (N_5793,N_5640,N_5592);
nand U5794 (N_5794,N_5553,N_5629);
or U5795 (N_5795,N_5605,N_5656);
nand U5796 (N_5796,N_5687,N_5610);
nor U5797 (N_5797,N_5649,N_5634);
nor U5798 (N_5798,N_5671,N_5678);
and U5799 (N_5799,N_5627,N_5578);
nor U5800 (N_5800,N_5658,N_5618);
and U5801 (N_5801,N_5625,N_5553);
nor U5802 (N_5802,N_5652,N_5580);
nand U5803 (N_5803,N_5649,N_5579);
or U5804 (N_5804,N_5585,N_5633);
and U5805 (N_5805,N_5662,N_5617);
nand U5806 (N_5806,N_5591,N_5564);
or U5807 (N_5807,N_5610,N_5657);
or U5808 (N_5808,N_5608,N_5621);
or U5809 (N_5809,N_5566,N_5587);
nor U5810 (N_5810,N_5594,N_5571);
and U5811 (N_5811,N_5677,N_5681);
nor U5812 (N_5812,N_5635,N_5594);
or U5813 (N_5813,N_5589,N_5645);
and U5814 (N_5814,N_5653,N_5582);
and U5815 (N_5815,N_5697,N_5665);
or U5816 (N_5816,N_5655,N_5603);
and U5817 (N_5817,N_5651,N_5640);
nor U5818 (N_5818,N_5668,N_5628);
xor U5819 (N_5819,N_5693,N_5556);
and U5820 (N_5820,N_5590,N_5607);
xor U5821 (N_5821,N_5683,N_5693);
xnor U5822 (N_5822,N_5582,N_5678);
nand U5823 (N_5823,N_5694,N_5680);
nor U5824 (N_5824,N_5673,N_5688);
xnor U5825 (N_5825,N_5674,N_5651);
and U5826 (N_5826,N_5683,N_5694);
or U5827 (N_5827,N_5650,N_5680);
or U5828 (N_5828,N_5595,N_5621);
xor U5829 (N_5829,N_5585,N_5657);
xor U5830 (N_5830,N_5692,N_5599);
and U5831 (N_5831,N_5623,N_5586);
nand U5832 (N_5832,N_5633,N_5693);
and U5833 (N_5833,N_5657,N_5639);
nor U5834 (N_5834,N_5691,N_5685);
or U5835 (N_5835,N_5591,N_5592);
nor U5836 (N_5836,N_5683,N_5580);
nand U5837 (N_5837,N_5579,N_5667);
xor U5838 (N_5838,N_5647,N_5640);
nand U5839 (N_5839,N_5560,N_5589);
or U5840 (N_5840,N_5667,N_5551);
nand U5841 (N_5841,N_5621,N_5618);
nand U5842 (N_5842,N_5695,N_5550);
and U5843 (N_5843,N_5595,N_5650);
or U5844 (N_5844,N_5674,N_5583);
or U5845 (N_5845,N_5676,N_5606);
or U5846 (N_5846,N_5596,N_5670);
nor U5847 (N_5847,N_5617,N_5606);
nor U5848 (N_5848,N_5685,N_5553);
and U5849 (N_5849,N_5622,N_5663);
or U5850 (N_5850,N_5791,N_5712);
nor U5851 (N_5851,N_5825,N_5711);
xnor U5852 (N_5852,N_5740,N_5783);
nor U5853 (N_5853,N_5835,N_5796);
nor U5854 (N_5854,N_5819,N_5846);
xor U5855 (N_5855,N_5839,N_5832);
or U5856 (N_5856,N_5763,N_5743);
nor U5857 (N_5857,N_5773,N_5709);
or U5858 (N_5858,N_5821,N_5826);
and U5859 (N_5859,N_5784,N_5751);
and U5860 (N_5860,N_5706,N_5787);
nand U5861 (N_5861,N_5812,N_5744);
and U5862 (N_5862,N_5775,N_5845);
xnor U5863 (N_5863,N_5716,N_5800);
nand U5864 (N_5864,N_5766,N_5785);
or U5865 (N_5865,N_5734,N_5713);
xor U5866 (N_5866,N_5736,N_5781);
nand U5867 (N_5867,N_5776,N_5718);
or U5868 (N_5868,N_5707,N_5842);
xnor U5869 (N_5869,N_5760,N_5808);
nor U5870 (N_5870,N_5822,N_5770);
nand U5871 (N_5871,N_5813,N_5721);
xnor U5872 (N_5872,N_5789,N_5757);
nor U5873 (N_5873,N_5729,N_5714);
and U5874 (N_5874,N_5725,N_5829);
nand U5875 (N_5875,N_5764,N_5798);
xor U5876 (N_5876,N_5782,N_5802);
or U5877 (N_5877,N_5752,N_5737);
and U5878 (N_5878,N_5779,N_5804);
and U5879 (N_5879,N_5806,N_5815);
or U5880 (N_5880,N_5818,N_5755);
nor U5881 (N_5881,N_5768,N_5727);
nor U5882 (N_5882,N_5717,N_5723);
xnor U5883 (N_5883,N_5724,N_5807);
nand U5884 (N_5884,N_5728,N_5774);
and U5885 (N_5885,N_5843,N_5816);
nand U5886 (N_5886,N_5747,N_5742);
nor U5887 (N_5887,N_5705,N_5795);
nand U5888 (N_5888,N_5769,N_5739);
xnor U5889 (N_5889,N_5735,N_5704);
xor U5890 (N_5890,N_5827,N_5814);
xnor U5891 (N_5891,N_5820,N_5817);
nor U5892 (N_5892,N_5792,N_5756);
nor U5893 (N_5893,N_5754,N_5794);
and U5894 (N_5894,N_5749,N_5838);
nor U5895 (N_5895,N_5710,N_5703);
and U5896 (N_5896,N_5748,N_5823);
and U5897 (N_5897,N_5700,N_5702);
and U5898 (N_5898,N_5730,N_5805);
or U5899 (N_5899,N_5758,N_5731);
or U5900 (N_5900,N_5831,N_5840);
nor U5901 (N_5901,N_5750,N_5797);
or U5902 (N_5902,N_5771,N_5722);
and U5903 (N_5903,N_5828,N_5790);
and U5904 (N_5904,N_5732,N_5793);
or U5905 (N_5905,N_5780,N_5811);
nor U5906 (N_5906,N_5741,N_5745);
nand U5907 (N_5907,N_5733,N_5841);
nor U5908 (N_5908,N_5772,N_5844);
and U5909 (N_5909,N_5761,N_5762);
and U5910 (N_5910,N_5809,N_5746);
xnor U5911 (N_5911,N_5834,N_5767);
xor U5912 (N_5912,N_5708,N_5833);
nor U5913 (N_5913,N_5837,N_5753);
xnor U5914 (N_5914,N_5720,N_5777);
nor U5915 (N_5915,N_5830,N_5836);
and U5916 (N_5916,N_5726,N_5848);
or U5917 (N_5917,N_5715,N_5824);
xor U5918 (N_5918,N_5799,N_5801);
nand U5919 (N_5919,N_5803,N_5847);
and U5920 (N_5920,N_5810,N_5786);
and U5921 (N_5921,N_5788,N_5759);
nor U5922 (N_5922,N_5719,N_5738);
nand U5923 (N_5923,N_5701,N_5778);
nor U5924 (N_5924,N_5765,N_5849);
nand U5925 (N_5925,N_5737,N_5719);
and U5926 (N_5926,N_5722,N_5754);
nor U5927 (N_5927,N_5738,N_5715);
nand U5928 (N_5928,N_5701,N_5747);
nand U5929 (N_5929,N_5790,N_5738);
or U5930 (N_5930,N_5798,N_5781);
xnor U5931 (N_5931,N_5805,N_5800);
xnor U5932 (N_5932,N_5833,N_5837);
nor U5933 (N_5933,N_5772,N_5833);
nor U5934 (N_5934,N_5743,N_5712);
and U5935 (N_5935,N_5771,N_5795);
and U5936 (N_5936,N_5813,N_5823);
xor U5937 (N_5937,N_5815,N_5754);
nor U5938 (N_5938,N_5809,N_5776);
or U5939 (N_5939,N_5809,N_5706);
nor U5940 (N_5940,N_5797,N_5810);
nor U5941 (N_5941,N_5701,N_5813);
xor U5942 (N_5942,N_5764,N_5702);
and U5943 (N_5943,N_5742,N_5799);
or U5944 (N_5944,N_5753,N_5734);
nor U5945 (N_5945,N_5705,N_5828);
and U5946 (N_5946,N_5840,N_5700);
or U5947 (N_5947,N_5821,N_5737);
nor U5948 (N_5948,N_5776,N_5773);
nand U5949 (N_5949,N_5844,N_5846);
xor U5950 (N_5950,N_5825,N_5738);
or U5951 (N_5951,N_5780,N_5782);
nor U5952 (N_5952,N_5801,N_5803);
and U5953 (N_5953,N_5790,N_5768);
or U5954 (N_5954,N_5741,N_5816);
nand U5955 (N_5955,N_5750,N_5723);
xnor U5956 (N_5956,N_5742,N_5840);
or U5957 (N_5957,N_5788,N_5771);
and U5958 (N_5958,N_5752,N_5779);
or U5959 (N_5959,N_5707,N_5785);
nand U5960 (N_5960,N_5830,N_5724);
nand U5961 (N_5961,N_5728,N_5733);
xor U5962 (N_5962,N_5739,N_5802);
nand U5963 (N_5963,N_5773,N_5779);
nand U5964 (N_5964,N_5725,N_5729);
nand U5965 (N_5965,N_5840,N_5797);
and U5966 (N_5966,N_5715,N_5807);
xor U5967 (N_5967,N_5782,N_5794);
and U5968 (N_5968,N_5831,N_5793);
or U5969 (N_5969,N_5775,N_5732);
and U5970 (N_5970,N_5800,N_5742);
and U5971 (N_5971,N_5718,N_5737);
and U5972 (N_5972,N_5824,N_5808);
and U5973 (N_5973,N_5719,N_5783);
nand U5974 (N_5974,N_5816,N_5805);
xor U5975 (N_5975,N_5730,N_5813);
nor U5976 (N_5976,N_5719,N_5833);
nand U5977 (N_5977,N_5785,N_5703);
nand U5978 (N_5978,N_5732,N_5713);
xnor U5979 (N_5979,N_5734,N_5726);
nor U5980 (N_5980,N_5833,N_5845);
nand U5981 (N_5981,N_5761,N_5780);
nor U5982 (N_5982,N_5714,N_5791);
nor U5983 (N_5983,N_5836,N_5800);
nor U5984 (N_5984,N_5744,N_5760);
nor U5985 (N_5985,N_5759,N_5820);
nand U5986 (N_5986,N_5729,N_5832);
nor U5987 (N_5987,N_5833,N_5712);
xor U5988 (N_5988,N_5815,N_5826);
or U5989 (N_5989,N_5805,N_5724);
and U5990 (N_5990,N_5728,N_5702);
nor U5991 (N_5991,N_5763,N_5839);
xnor U5992 (N_5992,N_5763,N_5830);
nor U5993 (N_5993,N_5753,N_5719);
or U5994 (N_5994,N_5726,N_5807);
nor U5995 (N_5995,N_5818,N_5806);
and U5996 (N_5996,N_5848,N_5710);
or U5997 (N_5997,N_5711,N_5794);
or U5998 (N_5998,N_5713,N_5764);
xor U5999 (N_5999,N_5799,N_5787);
nand U6000 (N_6000,N_5924,N_5957);
or U6001 (N_6001,N_5907,N_5855);
and U6002 (N_6002,N_5937,N_5895);
nand U6003 (N_6003,N_5999,N_5901);
and U6004 (N_6004,N_5860,N_5972);
or U6005 (N_6005,N_5906,N_5927);
nor U6006 (N_6006,N_5915,N_5951);
nand U6007 (N_6007,N_5880,N_5973);
xor U6008 (N_6008,N_5894,N_5938);
or U6009 (N_6009,N_5875,N_5869);
xnor U6010 (N_6010,N_5891,N_5934);
xnor U6011 (N_6011,N_5959,N_5867);
nor U6012 (N_6012,N_5931,N_5940);
nand U6013 (N_6013,N_5879,N_5917);
nand U6014 (N_6014,N_5984,N_5893);
and U6015 (N_6015,N_5864,N_5922);
or U6016 (N_6016,N_5939,N_5936);
and U6017 (N_6017,N_5863,N_5868);
or U6018 (N_6018,N_5956,N_5994);
xnor U6019 (N_6019,N_5920,N_5947);
nor U6020 (N_6020,N_5892,N_5919);
or U6021 (N_6021,N_5884,N_5882);
or U6022 (N_6022,N_5905,N_5913);
nor U6023 (N_6023,N_5996,N_5923);
nor U6024 (N_6024,N_5997,N_5995);
xnor U6025 (N_6025,N_5900,N_5970);
nor U6026 (N_6026,N_5989,N_5904);
or U6027 (N_6027,N_5878,N_5902);
and U6028 (N_6028,N_5949,N_5852);
xor U6029 (N_6029,N_5945,N_5916);
and U6030 (N_6030,N_5876,N_5914);
or U6031 (N_6031,N_5877,N_5952);
nor U6032 (N_6032,N_5953,N_5909);
xor U6033 (N_6033,N_5911,N_5992);
nor U6034 (N_6034,N_5975,N_5966);
nand U6035 (N_6035,N_5883,N_5941);
or U6036 (N_6036,N_5859,N_5955);
xor U6037 (N_6037,N_5964,N_5978);
xor U6038 (N_6038,N_5933,N_5946);
nand U6039 (N_6039,N_5993,N_5908);
and U6040 (N_6040,N_5881,N_5858);
or U6041 (N_6041,N_5888,N_5963);
or U6042 (N_6042,N_5854,N_5899);
xnor U6043 (N_6043,N_5974,N_5958);
nor U6044 (N_6044,N_5930,N_5874);
xor U6045 (N_6045,N_5950,N_5967);
and U6046 (N_6046,N_5857,N_5932);
xor U6047 (N_6047,N_5921,N_5896);
or U6048 (N_6048,N_5987,N_5856);
nor U6049 (N_6049,N_5965,N_5969);
xor U6050 (N_6050,N_5998,N_5925);
and U6051 (N_6051,N_5929,N_5981);
or U6052 (N_6052,N_5977,N_5935);
nand U6053 (N_6053,N_5886,N_5903);
nand U6054 (N_6054,N_5890,N_5850);
and U6055 (N_6055,N_5983,N_5926);
xor U6056 (N_6056,N_5871,N_5870);
nand U6057 (N_6057,N_5943,N_5898);
and U6058 (N_6058,N_5897,N_5866);
or U6059 (N_6059,N_5991,N_5872);
or U6060 (N_6060,N_5986,N_5961);
and U6061 (N_6061,N_5990,N_5985);
nand U6062 (N_6062,N_5885,N_5980);
nor U6063 (N_6063,N_5865,N_5912);
or U6064 (N_6064,N_5928,N_5948);
xnor U6065 (N_6065,N_5982,N_5942);
xor U6066 (N_6066,N_5979,N_5988);
xor U6067 (N_6067,N_5971,N_5887);
nand U6068 (N_6068,N_5968,N_5862);
nand U6069 (N_6069,N_5861,N_5962);
and U6070 (N_6070,N_5944,N_5910);
or U6071 (N_6071,N_5873,N_5918);
nand U6072 (N_6072,N_5954,N_5853);
nand U6073 (N_6073,N_5976,N_5851);
nand U6074 (N_6074,N_5889,N_5960);
nand U6075 (N_6075,N_5963,N_5880);
xor U6076 (N_6076,N_5930,N_5898);
nand U6077 (N_6077,N_5973,N_5981);
or U6078 (N_6078,N_5975,N_5937);
nor U6079 (N_6079,N_5856,N_5995);
nor U6080 (N_6080,N_5917,N_5937);
or U6081 (N_6081,N_5927,N_5907);
nor U6082 (N_6082,N_5850,N_5952);
xnor U6083 (N_6083,N_5943,N_5931);
xnor U6084 (N_6084,N_5947,N_5892);
xor U6085 (N_6085,N_5865,N_5857);
and U6086 (N_6086,N_5956,N_5985);
or U6087 (N_6087,N_5944,N_5894);
or U6088 (N_6088,N_5993,N_5963);
nand U6089 (N_6089,N_5964,N_5856);
nor U6090 (N_6090,N_5855,N_5888);
nor U6091 (N_6091,N_5924,N_5988);
and U6092 (N_6092,N_5966,N_5965);
xnor U6093 (N_6093,N_5917,N_5871);
and U6094 (N_6094,N_5883,N_5899);
nand U6095 (N_6095,N_5897,N_5896);
xnor U6096 (N_6096,N_5880,N_5951);
and U6097 (N_6097,N_5985,N_5871);
nor U6098 (N_6098,N_5975,N_5869);
or U6099 (N_6099,N_5981,N_5859);
nor U6100 (N_6100,N_5900,N_5864);
and U6101 (N_6101,N_5900,N_5902);
nand U6102 (N_6102,N_5906,N_5852);
or U6103 (N_6103,N_5869,N_5913);
nor U6104 (N_6104,N_5871,N_5891);
xor U6105 (N_6105,N_5917,N_5901);
nand U6106 (N_6106,N_5870,N_5977);
nor U6107 (N_6107,N_5903,N_5874);
or U6108 (N_6108,N_5852,N_5971);
nor U6109 (N_6109,N_5941,N_5964);
and U6110 (N_6110,N_5860,N_5951);
xor U6111 (N_6111,N_5954,N_5870);
or U6112 (N_6112,N_5993,N_5878);
or U6113 (N_6113,N_5862,N_5877);
and U6114 (N_6114,N_5991,N_5978);
nor U6115 (N_6115,N_5976,N_5884);
and U6116 (N_6116,N_5861,N_5928);
and U6117 (N_6117,N_5875,N_5939);
or U6118 (N_6118,N_5917,N_5946);
xor U6119 (N_6119,N_5875,N_5894);
nand U6120 (N_6120,N_5987,N_5960);
nor U6121 (N_6121,N_5904,N_5952);
and U6122 (N_6122,N_5950,N_5957);
or U6123 (N_6123,N_5994,N_5903);
nand U6124 (N_6124,N_5898,N_5950);
xor U6125 (N_6125,N_5850,N_5864);
and U6126 (N_6126,N_5896,N_5957);
xor U6127 (N_6127,N_5891,N_5931);
and U6128 (N_6128,N_5935,N_5865);
nand U6129 (N_6129,N_5876,N_5933);
xor U6130 (N_6130,N_5970,N_5953);
or U6131 (N_6131,N_5947,N_5954);
xnor U6132 (N_6132,N_5950,N_5965);
and U6133 (N_6133,N_5995,N_5927);
nand U6134 (N_6134,N_5949,N_5940);
nand U6135 (N_6135,N_5877,N_5867);
and U6136 (N_6136,N_5986,N_5889);
and U6137 (N_6137,N_5860,N_5961);
xnor U6138 (N_6138,N_5881,N_5983);
or U6139 (N_6139,N_5884,N_5854);
and U6140 (N_6140,N_5995,N_5931);
nand U6141 (N_6141,N_5852,N_5935);
nor U6142 (N_6142,N_5976,N_5882);
nand U6143 (N_6143,N_5936,N_5937);
nand U6144 (N_6144,N_5972,N_5859);
or U6145 (N_6145,N_5960,N_5914);
nor U6146 (N_6146,N_5916,N_5946);
nand U6147 (N_6147,N_5971,N_5939);
xnor U6148 (N_6148,N_5882,N_5944);
or U6149 (N_6149,N_5994,N_5895);
nand U6150 (N_6150,N_6049,N_6080);
nor U6151 (N_6151,N_6042,N_6017);
nor U6152 (N_6152,N_6109,N_6000);
and U6153 (N_6153,N_6142,N_6099);
xnor U6154 (N_6154,N_6029,N_6096);
xnor U6155 (N_6155,N_6100,N_6079);
or U6156 (N_6156,N_6120,N_6038);
nor U6157 (N_6157,N_6069,N_6115);
or U6158 (N_6158,N_6065,N_6083);
and U6159 (N_6159,N_6018,N_6057);
and U6160 (N_6160,N_6051,N_6074);
nand U6161 (N_6161,N_6062,N_6147);
nor U6162 (N_6162,N_6002,N_6022);
nand U6163 (N_6163,N_6048,N_6033);
and U6164 (N_6164,N_6039,N_6047);
or U6165 (N_6165,N_6144,N_6112);
and U6166 (N_6166,N_6108,N_6110);
xor U6167 (N_6167,N_6136,N_6082);
nor U6168 (N_6168,N_6034,N_6046);
nand U6169 (N_6169,N_6116,N_6055);
and U6170 (N_6170,N_6035,N_6043);
nand U6171 (N_6171,N_6012,N_6061);
nor U6172 (N_6172,N_6078,N_6119);
nand U6173 (N_6173,N_6124,N_6103);
or U6174 (N_6174,N_6032,N_6113);
nor U6175 (N_6175,N_6041,N_6107);
xnor U6176 (N_6176,N_6006,N_6084);
or U6177 (N_6177,N_6127,N_6092);
xor U6178 (N_6178,N_6016,N_6148);
and U6179 (N_6179,N_6102,N_6132);
or U6180 (N_6180,N_6126,N_6104);
xor U6181 (N_6181,N_6134,N_6141);
xor U6182 (N_6182,N_6011,N_6009);
or U6183 (N_6183,N_6072,N_6137);
and U6184 (N_6184,N_6088,N_6063);
xor U6185 (N_6185,N_6001,N_6005);
and U6186 (N_6186,N_6117,N_6138);
nand U6187 (N_6187,N_6027,N_6026);
xnor U6188 (N_6188,N_6024,N_6007);
or U6189 (N_6189,N_6060,N_6093);
xnor U6190 (N_6190,N_6066,N_6135);
nand U6191 (N_6191,N_6025,N_6053);
or U6192 (N_6192,N_6014,N_6028);
nor U6193 (N_6193,N_6067,N_6094);
nand U6194 (N_6194,N_6105,N_6097);
xnor U6195 (N_6195,N_6045,N_6122);
or U6196 (N_6196,N_6070,N_6020);
xnor U6197 (N_6197,N_6073,N_6149);
and U6198 (N_6198,N_6008,N_6081);
and U6199 (N_6199,N_6146,N_6023);
nor U6200 (N_6200,N_6118,N_6010);
or U6201 (N_6201,N_6095,N_6111);
nand U6202 (N_6202,N_6101,N_6013);
xnor U6203 (N_6203,N_6003,N_6071);
nor U6204 (N_6204,N_6086,N_6125);
nor U6205 (N_6205,N_6031,N_6121);
or U6206 (N_6206,N_6052,N_6004);
or U6207 (N_6207,N_6085,N_6059);
and U6208 (N_6208,N_6077,N_6015);
and U6209 (N_6209,N_6139,N_6131);
nand U6210 (N_6210,N_6106,N_6145);
nand U6211 (N_6211,N_6130,N_6036);
nor U6212 (N_6212,N_6089,N_6133);
nand U6213 (N_6213,N_6064,N_6075);
and U6214 (N_6214,N_6098,N_6050);
nand U6215 (N_6215,N_6091,N_6021);
nor U6216 (N_6216,N_6128,N_6123);
nor U6217 (N_6217,N_6040,N_6030);
xnor U6218 (N_6218,N_6054,N_6087);
xor U6219 (N_6219,N_6129,N_6140);
xor U6220 (N_6220,N_6076,N_6056);
nand U6221 (N_6221,N_6044,N_6090);
and U6222 (N_6222,N_6143,N_6068);
and U6223 (N_6223,N_6058,N_6114);
xor U6224 (N_6224,N_6019,N_6037);
or U6225 (N_6225,N_6145,N_6061);
nor U6226 (N_6226,N_6103,N_6112);
xor U6227 (N_6227,N_6045,N_6093);
nand U6228 (N_6228,N_6145,N_6139);
xor U6229 (N_6229,N_6025,N_6096);
and U6230 (N_6230,N_6074,N_6121);
or U6231 (N_6231,N_6072,N_6092);
or U6232 (N_6232,N_6131,N_6109);
and U6233 (N_6233,N_6045,N_6073);
xnor U6234 (N_6234,N_6039,N_6140);
and U6235 (N_6235,N_6063,N_6099);
nand U6236 (N_6236,N_6087,N_6056);
nand U6237 (N_6237,N_6067,N_6108);
xor U6238 (N_6238,N_6003,N_6041);
xor U6239 (N_6239,N_6146,N_6074);
nor U6240 (N_6240,N_6105,N_6050);
nor U6241 (N_6241,N_6074,N_6088);
nor U6242 (N_6242,N_6147,N_6059);
or U6243 (N_6243,N_6073,N_6129);
nor U6244 (N_6244,N_6026,N_6051);
or U6245 (N_6245,N_6120,N_6019);
nor U6246 (N_6246,N_6062,N_6040);
nor U6247 (N_6247,N_6036,N_6017);
nor U6248 (N_6248,N_6028,N_6043);
nand U6249 (N_6249,N_6083,N_6123);
and U6250 (N_6250,N_6065,N_6022);
xnor U6251 (N_6251,N_6032,N_6054);
nand U6252 (N_6252,N_6035,N_6054);
or U6253 (N_6253,N_6044,N_6127);
and U6254 (N_6254,N_6084,N_6075);
and U6255 (N_6255,N_6068,N_6111);
nand U6256 (N_6256,N_6082,N_6115);
and U6257 (N_6257,N_6124,N_6041);
or U6258 (N_6258,N_6069,N_6005);
nand U6259 (N_6259,N_6050,N_6124);
nor U6260 (N_6260,N_6058,N_6097);
nand U6261 (N_6261,N_6042,N_6104);
or U6262 (N_6262,N_6067,N_6148);
or U6263 (N_6263,N_6090,N_6050);
xor U6264 (N_6264,N_6086,N_6126);
or U6265 (N_6265,N_6072,N_6067);
nand U6266 (N_6266,N_6121,N_6013);
or U6267 (N_6267,N_6064,N_6092);
or U6268 (N_6268,N_6146,N_6087);
nand U6269 (N_6269,N_6011,N_6125);
and U6270 (N_6270,N_6082,N_6078);
nor U6271 (N_6271,N_6047,N_6102);
xnor U6272 (N_6272,N_6059,N_6122);
nor U6273 (N_6273,N_6072,N_6075);
or U6274 (N_6274,N_6103,N_6053);
or U6275 (N_6275,N_6043,N_6023);
or U6276 (N_6276,N_6148,N_6018);
or U6277 (N_6277,N_6002,N_6057);
and U6278 (N_6278,N_6041,N_6135);
nand U6279 (N_6279,N_6095,N_6092);
and U6280 (N_6280,N_6149,N_6065);
and U6281 (N_6281,N_6127,N_6077);
and U6282 (N_6282,N_6018,N_6106);
or U6283 (N_6283,N_6080,N_6051);
or U6284 (N_6284,N_6106,N_6000);
or U6285 (N_6285,N_6084,N_6055);
or U6286 (N_6286,N_6104,N_6034);
or U6287 (N_6287,N_6091,N_6132);
xor U6288 (N_6288,N_6121,N_6133);
or U6289 (N_6289,N_6063,N_6004);
xor U6290 (N_6290,N_6104,N_6142);
and U6291 (N_6291,N_6033,N_6057);
and U6292 (N_6292,N_6008,N_6076);
and U6293 (N_6293,N_6129,N_6061);
nor U6294 (N_6294,N_6120,N_6004);
and U6295 (N_6295,N_6076,N_6140);
or U6296 (N_6296,N_6067,N_6062);
or U6297 (N_6297,N_6027,N_6069);
nor U6298 (N_6298,N_6023,N_6124);
or U6299 (N_6299,N_6143,N_6135);
xnor U6300 (N_6300,N_6241,N_6255);
nor U6301 (N_6301,N_6250,N_6265);
nand U6302 (N_6302,N_6261,N_6285);
nor U6303 (N_6303,N_6284,N_6162);
and U6304 (N_6304,N_6259,N_6268);
nor U6305 (N_6305,N_6166,N_6158);
nand U6306 (N_6306,N_6172,N_6231);
xnor U6307 (N_6307,N_6191,N_6297);
xor U6308 (N_6308,N_6173,N_6267);
nand U6309 (N_6309,N_6164,N_6181);
or U6310 (N_6310,N_6154,N_6197);
and U6311 (N_6311,N_6274,N_6245);
or U6312 (N_6312,N_6249,N_6209);
nand U6313 (N_6313,N_6187,N_6206);
xor U6314 (N_6314,N_6228,N_6283);
or U6315 (N_6315,N_6253,N_6290);
nand U6316 (N_6316,N_6163,N_6183);
nor U6317 (N_6317,N_6160,N_6161);
nand U6318 (N_6318,N_6215,N_6214);
nand U6319 (N_6319,N_6272,N_6177);
and U6320 (N_6320,N_6294,N_6157);
or U6321 (N_6321,N_6202,N_6243);
nor U6322 (N_6322,N_6169,N_6170);
and U6323 (N_6323,N_6180,N_6251);
nand U6324 (N_6324,N_6263,N_6193);
nor U6325 (N_6325,N_6208,N_6168);
nor U6326 (N_6326,N_6198,N_6273);
nand U6327 (N_6327,N_6195,N_6229);
or U6328 (N_6328,N_6182,N_6280);
xor U6329 (N_6329,N_6210,N_6174);
nand U6330 (N_6330,N_6194,N_6221);
and U6331 (N_6331,N_6151,N_6244);
and U6332 (N_6332,N_6156,N_6213);
and U6333 (N_6333,N_6188,N_6207);
xor U6334 (N_6334,N_6165,N_6176);
and U6335 (N_6335,N_6204,N_6262);
or U6336 (N_6336,N_6222,N_6242);
nand U6337 (N_6337,N_6211,N_6270);
and U6338 (N_6338,N_6153,N_6282);
or U6339 (N_6339,N_6257,N_6240);
xor U6340 (N_6340,N_6246,N_6276);
nor U6341 (N_6341,N_6237,N_6277);
or U6342 (N_6342,N_6186,N_6150);
xor U6343 (N_6343,N_6235,N_6266);
or U6344 (N_6344,N_6260,N_6289);
nor U6345 (N_6345,N_6203,N_6178);
nor U6346 (N_6346,N_6252,N_6279);
nor U6347 (N_6347,N_6239,N_6291);
nand U6348 (N_6348,N_6220,N_6296);
nor U6349 (N_6349,N_6216,N_6212);
nor U6350 (N_6350,N_6256,N_6155);
xor U6351 (N_6351,N_6269,N_6200);
nor U6352 (N_6352,N_6264,N_6217);
and U6353 (N_6353,N_6190,N_6184);
nand U6354 (N_6354,N_6278,N_6254);
xnor U6355 (N_6355,N_6224,N_6258);
nand U6356 (N_6356,N_6225,N_6288);
and U6357 (N_6357,N_6189,N_6185);
and U6358 (N_6358,N_6230,N_6292);
and U6359 (N_6359,N_6226,N_6293);
nor U6360 (N_6360,N_6299,N_6192);
or U6361 (N_6361,N_6227,N_6232);
nand U6362 (N_6362,N_6218,N_6175);
xor U6363 (N_6363,N_6275,N_6234);
or U6364 (N_6364,N_6205,N_6199);
or U6365 (N_6365,N_6298,N_6201);
nor U6366 (N_6366,N_6295,N_6247);
nand U6367 (N_6367,N_6219,N_6248);
nand U6368 (N_6368,N_6171,N_6152);
nor U6369 (N_6369,N_6233,N_6286);
xor U6370 (N_6370,N_6179,N_6167);
nand U6371 (N_6371,N_6236,N_6196);
nor U6372 (N_6372,N_6238,N_6287);
nor U6373 (N_6373,N_6159,N_6281);
nand U6374 (N_6374,N_6271,N_6223);
nand U6375 (N_6375,N_6253,N_6241);
nand U6376 (N_6376,N_6230,N_6250);
nand U6377 (N_6377,N_6186,N_6225);
or U6378 (N_6378,N_6271,N_6199);
or U6379 (N_6379,N_6153,N_6212);
and U6380 (N_6380,N_6263,N_6188);
or U6381 (N_6381,N_6230,N_6285);
or U6382 (N_6382,N_6203,N_6285);
and U6383 (N_6383,N_6255,N_6181);
or U6384 (N_6384,N_6185,N_6249);
xor U6385 (N_6385,N_6276,N_6286);
or U6386 (N_6386,N_6261,N_6244);
nand U6387 (N_6387,N_6219,N_6210);
or U6388 (N_6388,N_6227,N_6158);
nor U6389 (N_6389,N_6207,N_6293);
nand U6390 (N_6390,N_6253,N_6185);
nand U6391 (N_6391,N_6196,N_6180);
nand U6392 (N_6392,N_6169,N_6298);
or U6393 (N_6393,N_6246,N_6251);
xnor U6394 (N_6394,N_6288,N_6296);
or U6395 (N_6395,N_6255,N_6197);
nor U6396 (N_6396,N_6164,N_6295);
or U6397 (N_6397,N_6298,N_6279);
xnor U6398 (N_6398,N_6183,N_6230);
xnor U6399 (N_6399,N_6157,N_6259);
or U6400 (N_6400,N_6260,N_6278);
xor U6401 (N_6401,N_6269,N_6185);
or U6402 (N_6402,N_6154,N_6298);
nor U6403 (N_6403,N_6184,N_6280);
nand U6404 (N_6404,N_6243,N_6166);
xnor U6405 (N_6405,N_6208,N_6276);
xor U6406 (N_6406,N_6165,N_6236);
nor U6407 (N_6407,N_6178,N_6233);
nor U6408 (N_6408,N_6227,N_6195);
xnor U6409 (N_6409,N_6196,N_6200);
nor U6410 (N_6410,N_6272,N_6235);
and U6411 (N_6411,N_6294,N_6188);
xnor U6412 (N_6412,N_6198,N_6252);
nand U6413 (N_6413,N_6184,N_6292);
nand U6414 (N_6414,N_6234,N_6239);
or U6415 (N_6415,N_6240,N_6282);
nand U6416 (N_6416,N_6242,N_6245);
nand U6417 (N_6417,N_6252,N_6271);
or U6418 (N_6418,N_6269,N_6205);
and U6419 (N_6419,N_6294,N_6263);
or U6420 (N_6420,N_6252,N_6267);
xnor U6421 (N_6421,N_6231,N_6283);
nor U6422 (N_6422,N_6296,N_6265);
xor U6423 (N_6423,N_6206,N_6231);
nand U6424 (N_6424,N_6201,N_6244);
nand U6425 (N_6425,N_6199,N_6226);
nor U6426 (N_6426,N_6298,N_6293);
nor U6427 (N_6427,N_6251,N_6255);
xor U6428 (N_6428,N_6222,N_6180);
nor U6429 (N_6429,N_6269,N_6165);
or U6430 (N_6430,N_6203,N_6247);
nor U6431 (N_6431,N_6212,N_6249);
nor U6432 (N_6432,N_6243,N_6224);
nand U6433 (N_6433,N_6290,N_6279);
nand U6434 (N_6434,N_6169,N_6264);
nor U6435 (N_6435,N_6237,N_6255);
or U6436 (N_6436,N_6167,N_6243);
nor U6437 (N_6437,N_6165,N_6285);
nor U6438 (N_6438,N_6229,N_6181);
or U6439 (N_6439,N_6218,N_6158);
and U6440 (N_6440,N_6201,N_6219);
xnor U6441 (N_6441,N_6188,N_6196);
and U6442 (N_6442,N_6221,N_6299);
nand U6443 (N_6443,N_6273,N_6219);
xnor U6444 (N_6444,N_6205,N_6292);
and U6445 (N_6445,N_6236,N_6163);
nand U6446 (N_6446,N_6172,N_6184);
nand U6447 (N_6447,N_6242,N_6293);
xor U6448 (N_6448,N_6192,N_6200);
nand U6449 (N_6449,N_6239,N_6271);
nand U6450 (N_6450,N_6383,N_6360);
and U6451 (N_6451,N_6422,N_6307);
nor U6452 (N_6452,N_6417,N_6394);
xor U6453 (N_6453,N_6319,N_6431);
xor U6454 (N_6454,N_6391,N_6312);
and U6455 (N_6455,N_6320,N_6359);
nor U6456 (N_6456,N_6435,N_6424);
nor U6457 (N_6457,N_6348,N_6304);
xnor U6458 (N_6458,N_6448,N_6306);
nand U6459 (N_6459,N_6334,N_6409);
or U6460 (N_6460,N_6336,N_6429);
nor U6461 (N_6461,N_6378,N_6329);
and U6462 (N_6462,N_6353,N_6367);
nand U6463 (N_6463,N_6311,N_6305);
nor U6464 (N_6464,N_6389,N_6405);
and U6465 (N_6465,N_6369,N_6321);
nor U6466 (N_6466,N_6423,N_6442);
nor U6467 (N_6467,N_6351,N_6364);
nor U6468 (N_6468,N_6421,N_6428);
xor U6469 (N_6469,N_6316,N_6434);
nor U6470 (N_6470,N_6408,N_6385);
nor U6471 (N_6471,N_6363,N_6355);
xor U6472 (N_6472,N_6386,N_6418);
xnor U6473 (N_6473,N_6390,N_6404);
nand U6474 (N_6474,N_6395,N_6380);
or U6475 (N_6475,N_6345,N_6433);
xor U6476 (N_6476,N_6436,N_6420);
xor U6477 (N_6477,N_6342,N_6384);
and U6478 (N_6478,N_6344,N_6358);
or U6479 (N_6479,N_6410,N_6432);
or U6480 (N_6480,N_6411,N_6349);
nand U6481 (N_6481,N_6443,N_6439);
nand U6482 (N_6482,N_6371,N_6375);
and U6483 (N_6483,N_6326,N_6396);
or U6484 (N_6484,N_6301,N_6343);
nor U6485 (N_6485,N_6315,N_6350);
or U6486 (N_6486,N_6317,N_6392);
and U6487 (N_6487,N_6346,N_6407);
and U6488 (N_6488,N_6400,N_6365);
xnor U6489 (N_6489,N_6366,N_6302);
nor U6490 (N_6490,N_6309,N_6425);
nand U6491 (N_6491,N_6310,N_6339);
and U6492 (N_6492,N_6340,N_6393);
and U6493 (N_6493,N_6446,N_6379);
nand U6494 (N_6494,N_6347,N_6413);
xor U6495 (N_6495,N_6427,N_6447);
nand U6496 (N_6496,N_6332,N_6303);
and U6497 (N_6497,N_6300,N_6357);
nand U6498 (N_6498,N_6376,N_6445);
or U6499 (N_6499,N_6324,N_6362);
and U6500 (N_6500,N_6361,N_6388);
or U6501 (N_6501,N_6314,N_6406);
xor U6502 (N_6502,N_6325,N_6426);
nor U6503 (N_6503,N_6412,N_6318);
xnor U6504 (N_6504,N_6437,N_6322);
nor U6505 (N_6505,N_6387,N_6330);
or U6506 (N_6506,N_6341,N_6430);
nor U6507 (N_6507,N_6449,N_6397);
xor U6508 (N_6508,N_6327,N_6352);
nor U6509 (N_6509,N_6377,N_6354);
xor U6510 (N_6510,N_6337,N_6356);
xor U6511 (N_6511,N_6328,N_6331);
and U6512 (N_6512,N_6403,N_6335);
xnor U6513 (N_6513,N_6416,N_6382);
xor U6514 (N_6514,N_6368,N_6333);
nand U6515 (N_6515,N_6374,N_6414);
or U6516 (N_6516,N_6402,N_6440);
and U6517 (N_6517,N_6441,N_6372);
or U6518 (N_6518,N_6308,N_6401);
xnor U6519 (N_6519,N_6323,N_6419);
nand U6520 (N_6520,N_6399,N_6438);
or U6521 (N_6521,N_6370,N_6398);
nand U6522 (N_6522,N_6313,N_6444);
or U6523 (N_6523,N_6381,N_6373);
xor U6524 (N_6524,N_6415,N_6338);
nand U6525 (N_6525,N_6400,N_6334);
and U6526 (N_6526,N_6397,N_6426);
and U6527 (N_6527,N_6345,N_6366);
and U6528 (N_6528,N_6446,N_6397);
nor U6529 (N_6529,N_6329,N_6426);
nor U6530 (N_6530,N_6302,N_6363);
nand U6531 (N_6531,N_6314,N_6421);
or U6532 (N_6532,N_6308,N_6424);
nand U6533 (N_6533,N_6365,N_6380);
and U6534 (N_6534,N_6378,N_6319);
or U6535 (N_6535,N_6304,N_6423);
xnor U6536 (N_6536,N_6383,N_6310);
and U6537 (N_6537,N_6358,N_6402);
xnor U6538 (N_6538,N_6395,N_6354);
and U6539 (N_6539,N_6425,N_6337);
nand U6540 (N_6540,N_6321,N_6309);
and U6541 (N_6541,N_6395,N_6355);
xor U6542 (N_6542,N_6312,N_6430);
or U6543 (N_6543,N_6379,N_6342);
and U6544 (N_6544,N_6335,N_6398);
nor U6545 (N_6545,N_6445,N_6395);
nand U6546 (N_6546,N_6307,N_6439);
xnor U6547 (N_6547,N_6437,N_6353);
nand U6548 (N_6548,N_6406,N_6319);
and U6549 (N_6549,N_6354,N_6410);
and U6550 (N_6550,N_6339,N_6334);
nand U6551 (N_6551,N_6363,N_6428);
nor U6552 (N_6552,N_6340,N_6417);
and U6553 (N_6553,N_6332,N_6345);
or U6554 (N_6554,N_6335,N_6302);
nor U6555 (N_6555,N_6385,N_6376);
and U6556 (N_6556,N_6357,N_6392);
nor U6557 (N_6557,N_6332,N_6419);
or U6558 (N_6558,N_6383,N_6351);
xnor U6559 (N_6559,N_6343,N_6387);
or U6560 (N_6560,N_6302,N_6442);
and U6561 (N_6561,N_6424,N_6395);
and U6562 (N_6562,N_6402,N_6308);
nand U6563 (N_6563,N_6347,N_6325);
nand U6564 (N_6564,N_6361,N_6400);
or U6565 (N_6565,N_6306,N_6344);
and U6566 (N_6566,N_6437,N_6339);
nand U6567 (N_6567,N_6394,N_6418);
or U6568 (N_6568,N_6439,N_6353);
and U6569 (N_6569,N_6439,N_6312);
nand U6570 (N_6570,N_6448,N_6314);
nand U6571 (N_6571,N_6319,N_6332);
xor U6572 (N_6572,N_6379,N_6419);
or U6573 (N_6573,N_6383,N_6342);
nor U6574 (N_6574,N_6354,N_6371);
xnor U6575 (N_6575,N_6401,N_6351);
nand U6576 (N_6576,N_6333,N_6419);
or U6577 (N_6577,N_6363,N_6309);
and U6578 (N_6578,N_6423,N_6438);
and U6579 (N_6579,N_6426,N_6395);
nand U6580 (N_6580,N_6349,N_6414);
and U6581 (N_6581,N_6384,N_6331);
xor U6582 (N_6582,N_6304,N_6388);
nand U6583 (N_6583,N_6448,N_6307);
and U6584 (N_6584,N_6407,N_6447);
xnor U6585 (N_6585,N_6406,N_6340);
nor U6586 (N_6586,N_6356,N_6411);
xor U6587 (N_6587,N_6439,N_6432);
xnor U6588 (N_6588,N_6406,N_6441);
nor U6589 (N_6589,N_6399,N_6439);
or U6590 (N_6590,N_6398,N_6408);
or U6591 (N_6591,N_6401,N_6314);
and U6592 (N_6592,N_6410,N_6318);
nand U6593 (N_6593,N_6400,N_6362);
xnor U6594 (N_6594,N_6304,N_6378);
nand U6595 (N_6595,N_6383,N_6305);
and U6596 (N_6596,N_6346,N_6312);
xnor U6597 (N_6597,N_6397,N_6406);
and U6598 (N_6598,N_6436,N_6327);
nand U6599 (N_6599,N_6441,N_6303);
xor U6600 (N_6600,N_6498,N_6537);
xor U6601 (N_6601,N_6493,N_6545);
or U6602 (N_6602,N_6465,N_6595);
nor U6603 (N_6603,N_6523,N_6520);
and U6604 (N_6604,N_6481,N_6473);
nand U6605 (N_6605,N_6486,N_6491);
and U6606 (N_6606,N_6578,N_6571);
and U6607 (N_6607,N_6457,N_6513);
nor U6608 (N_6608,N_6459,N_6532);
nand U6609 (N_6609,N_6560,N_6474);
nor U6610 (N_6610,N_6499,N_6508);
xnor U6611 (N_6611,N_6553,N_6480);
nand U6612 (N_6612,N_6562,N_6590);
nor U6613 (N_6613,N_6494,N_6582);
xnor U6614 (N_6614,N_6460,N_6502);
xnor U6615 (N_6615,N_6490,N_6495);
xor U6616 (N_6616,N_6470,N_6552);
nor U6617 (N_6617,N_6546,N_6462);
or U6618 (N_6618,N_6554,N_6584);
nand U6619 (N_6619,N_6558,N_6489);
or U6620 (N_6620,N_6514,N_6484);
nor U6621 (N_6621,N_6591,N_6540);
and U6622 (N_6622,N_6526,N_6570);
nor U6623 (N_6623,N_6556,N_6456);
nor U6624 (N_6624,N_6507,N_6544);
nand U6625 (N_6625,N_6469,N_6557);
and U6626 (N_6626,N_6451,N_6505);
nand U6627 (N_6627,N_6482,N_6521);
xor U6628 (N_6628,N_6463,N_6561);
and U6629 (N_6629,N_6565,N_6536);
nand U6630 (N_6630,N_6577,N_6568);
xnor U6631 (N_6631,N_6538,N_6551);
xor U6632 (N_6632,N_6478,N_6547);
xor U6633 (N_6633,N_6483,N_6496);
nand U6634 (N_6634,N_6468,N_6450);
or U6635 (N_6635,N_6454,N_6501);
and U6636 (N_6636,N_6572,N_6485);
xor U6637 (N_6637,N_6517,N_6510);
nand U6638 (N_6638,N_6472,N_6587);
nand U6639 (N_6639,N_6586,N_6476);
xnor U6640 (N_6640,N_6597,N_6524);
nand U6641 (N_6641,N_6539,N_6580);
and U6642 (N_6642,N_6464,N_6458);
or U6643 (N_6643,N_6549,N_6567);
nand U6644 (N_6644,N_6550,N_6529);
and U6645 (N_6645,N_6500,N_6576);
or U6646 (N_6646,N_6585,N_6555);
nand U6647 (N_6647,N_6592,N_6596);
and U6648 (N_6648,N_6455,N_6598);
xor U6649 (N_6649,N_6594,N_6509);
and U6650 (N_6650,N_6581,N_6515);
xor U6651 (N_6651,N_6522,N_6527);
nor U6652 (N_6652,N_6575,N_6471);
or U6653 (N_6653,N_6467,N_6488);
nand U6654 (N_6654,N_6530,N_6511);
and U6655 (N_6655,N_6531,N_6559);
nand U6656 (N_6656,N_6589,N_6543);
nor U6657 (N_6657,N_6588,N_6512);
nand U6658 (N_6658,N_6519,N_6492);
and U6659 (N_6659,N_6548,N_6487);
xnor U6660 (N_6660,N_6516,N_6533);
or U6661 (N_6661,N_6504,N_6475);
nor U6662 (N_6662,N_6466,N_6461);
and U6663 (N_6663,N_6579,N_6573);
or U6664 (N_6664,N_6583,N_6569);
or U6665 (N_6665,N_6452,N_6479);
xnor U6666 (N_6666,N_6506,N_6497);
and U6667 (N_6667,N_6542,N_6593);
nor U6668 (N_6668,N_6574,N_6541);
xor U6669 (N_6669,N_6534,N_6453);
or U6670 (N_6670,N_6518,N_6599);
xnor U6671 (N_6671,N_6503,N_6477);
or U6672 (N_6672,N_6566,N_6563);
and U6673 (N_6673,N_6564,N_6528);
and U6674 (N_6674,N_6535,N_6525);
and U6675 (N_6675,N_6594,N_6493);
nor U6676 (N_6676,N_6518,N_6595);
or U6677 (N_6677,N_6522,N_6474);
or U6678 (N_6678,N_6581,N_6462);
and U6679 (N_6679,N_6581,N_6460);
and U6680 (N_6680,N_6573,N_6598);
nand U6681 (N_6681,N_6548,N_6480);
nand U6682 (N_6682,N_6579,N_6536);
nand U6683 (N_6683,N_6496,N_6479);
nand U6684 (N_6684,N_6500,N_6526);
nor U6685 (N_6685,N_6532,N_6506);
or U6686 (N_6686,N_6543,N_6455);
nand U6687 (N_6687,N_6521,N_6451);
and U6688 (N_6688,N_6531,N_6562);
and U6689 (N_6689,N_6557,N_6543);
or U6690 (N_6690,N_6505,N_6572);
nand U6691 (N_6691,N_6531,N_6569);
nand U6692 (N_6692,N_6490,N_6502);
nand U6693 (N_6693,N_6533,N_6500);
nand U6694 (N_6694,N_6525,N_6565);
xor U6695 (N_6695,N_6492,N_6473);
nand U6696 (N_6696,N_6556,N_6538);
nand U6697 (N_6697,N_6547,N_6578);
nand U6698 (N_6698,N_6556,N_6589);
or U6699 (N_6699,N_6455,N_6527);
nand U6700 (N_6700,N_6585,N_6575);
nand U6701 (N_6701,N_6553,N_6564);
nor U6702 (N_6702,N_6523,N_6478);
nand U6703 (N_6703,N_6466,N_6535);
and U6704 (N_6704,N_6473,N_6457);
nor U6705 (N_6705,N_6591,N_6515);
or U6706 (N_6706,N_6491,N_6459);
xor U6707 (N_6707,N_6554,N_6522);
xor U6708 (N_6708,N_6556,N_6581);
xor U6709 (N_6709,N_6551,N_6567);
or U6710 (N_6710,N_6546,N_6545);
nor U6711 (N_6711,N_6463,N_6530);
or U6712 (N_6712,N_6519,N_6522);
nand U6713 (N_6713,N_6519,N_6529);
nand U6714 (N_6714,N_6550,N_6495);
nand U6715 (N_6715,N_6570,N_6596);
xnor U6716 (N_6716,N_6596,N_6516);
or U6717 (N_6717,N_6490,N_6589);
nor U6718 (N_6718,N_6452,N_6496);
nor U6719 (N_6719,N_6467,N_6470);
xor U6720 (N_6720,N_6535,N_6472);
or U6721 (N_6721,N_6527,N_6519);
nand U6722 (N_6722,N_6490,N_6571);
xor U6723 (N_6723,N_6480,N_6506);
or U6724 (N_6724,N_6474,N_6574);
and U6725 (N_6725,N_6568,N_6570);
nand U6726 (N_6726,N_6530,N_6519);
or U6727 (N_6727,N_6461,N_6589);
xor U6728 (N_6728,N_6546,N_6564);
or U6729 (N_6729,N_6467,N_6594);
or U6730 (N_6730,N_6503,N_6557);
nand U6731 (N_6731,N_6538,N_6576);
nand U6732 (N_6732,N_6567,N_6526);
and U6733 (N_6733,N_6506,N_6512);
nor U6734 (N_6734,N_6492,N_6531);
nand U6735 (N_6735,N_6489,N_6505);
nand U6736 (N_6736,N_6494,N_6568);
nand U6737 (N_6737,N_6513,N_6537);
nand U6738 (N_6738,N_6585,N_6525);
xor U6739 (N_6739,N_6493,N_6578);
nand U6740 (N_6740,N_6590,N_6555);
or U6741 (N_6741,N_6562,N_6492);
nor U6742 (N_6742,N_6592,N_6452);
xor U6743 (N_6743,N_6469,N_6456);
nor U6744 (N_6744,N_6535,N_6597);
xor U6745 (N_6745,N_6483,N_6566);
nand U6746 (N_6746,N_6539,N_6599);
nor U6747 (N_6747,N_6536,N_6585);
or U6748 (N_6748,N_6543,N_6596);
nand U6749 (N_6749,N_6522,N_6588);
and U6750 (N_6750,N_6645,N_6652);
and U6751 (N_6751,N_6654,N_6719);
or U6752 (N_6752,N_6702,N_6668);
nand U6753 (N_6753,N_6633,N_6647);
or U6754 (N_6754,N_6665,N_6722);
nor U6755 (N_6755,N_6679,N_6733);
nand U6756 (N_6756,N_6746,N_6691);
nand U6757 (N_6757,N_6607,N_6666);
xor U6758 (N_6758,N_6659,N_6677);
nor U6759 (N_6759,N_6723,N_6644);
and U6760 (N_6760,N_6735,N_6676);
xor U6761 (N_6761,N_6646,N_6673);
and U6762 (N_6762,N_6749,N_6720);
xor U6763 (N_6763,N_6726,N_6609);
or U6764 (N_6764,N_6636,N_6663);
and U6765 (N_6765,N_6614,N_6731);
nand U6766 (N_6766,N_6747,N_6724);
and U6767 (N_6767,N_6641,N_6718);
or U6768 (N_6768,N_6717,N_6648);
and U6769 (N_6769,N_6623,N_6627);
or U6770 (N_6770,N_6699,N_6701);
nand U6771 (N_6771,N_6670,N_6738);
nand U6772 (N_6772,N_6605,N_6704);
nand U6773 (N_6773,N_6671,N_6692);
and U6774 (N_6774,N_6730,N_6740);
nand U6775 (N_6775,N_6669,N_6656);
xor U6776 (N_6776,N_6721,N_6618);
or U6777 (N_6777,N_6682,N_6629);
or U6778 (N_6778,N_6684,N_6628);
or U6779 (N_6779,N_6615,N_6608);
and U6780 (N_6780,N_6634,N_6693);
nor U6781 (N_6781,N_6700,N_6606);
nand U6782 (N_6782,N_6620,N_6748);
nor U6783 (N_6783,N_6643,N_6617);
nand U6784 (N_6784,N_6743,N_6706);
and U6785 (N_6785,N_6680,N_6619);
or U6786 (N_6786,N_6660,N_6600);
and U6787 (N_6787,N_6672,N_6661);
xor U6788 (N_6788,N_6732,N_6639);
or U6789 (N_6789,N_6739,N_6637);
xnor U6790 (N_6790,N_6709,N_6621);
or U6791 (N_6791,N_6744,N_6694);
xnor U6792 (N_6792,N_6696,N_6626);
xnor U6793 (N_6793,N_6632,N_6667);
nor U6794 (N_6794,N_6745,N_6662);
nand U6795 (N_6795,N_6674,N_6604);
nand U6796 (N_6796,N_6707,N_6642);
xor U6797 (N_6797,N_6697,N_6729);
xnor U6798 (N_6798,N_6678,N_6630);
nor U6799 (N_6799,N_6716,N_6631);
or U6800 (N_6800,N_6708,N_6741);
and U6801 (N_6801,N_6601,N_6742);
or U6802 (N_6802,N_6736,N_6635);
and U6803 (N_6803,N_6651,N_6727);
or U6804 (N_6804,N_6650,N_6613);
nand U6805 (N_6805,N_6603,N_6689);
xor U6806 (N_6806,N_6687,N_6664);
and U6807 (N_6807,N_6711,N_6658);
nor U6808 (N_6808,N_6681,N_6622);
and U6809 (N_6809,N_6640,N_6690);
or U6810 (N_6810,N_6655,N_6695);
and U6811 (N_6811,N_6649,N_6685);
xor U6812 (N_6812,N_6657,N_6715);
nor U6813 (N_6813,N_6612,N_6705);
and U6814 (N_6814,N_6734,N_6616);
nor U6815 (N_6815,N_6714,N_6602);
nor U6816 (N_6816,N_6698,N_6688);
xor U6817 (N_6817,N_6611,N_6725);
or U6818 (N_6818,N_6703,N_6710);
or U6819 (N_6819,N_6624,N_6737);
xor U6820 (N_6820,N_6713,N_6675);
nand U6821 (N_6821,N_6638,N_6653);
nand U6822 (N_6822,N_6728,N_6683);
nand U6823 (N_6823,N_6625,N_6712);
nor U6824 (N_6824,N_6686,N_6610);
nor U6825 (N_6825,N_6628,N_6601);
xor U6826 (N_6826,N_6652,N_6712);
or U6827 (N_6827,N_6749,N_6683);
and U6828 (N_6828,N_6628,N_6698);
nand U6829 (N_6829,N_6635,N_6685);
or U6830 (N_6830,N_6620,N_6631);
and U6831 (N_6831,N_6635,N_6642);
or U6832 (N_6832,N_6646,N_6726);
and U6833 (N_6833,N_6708,N_6601);
or U6834 (N_6834,N_6605,N_6663);
or U6835 (N_6835,N_6732,N_6701);
xnor U6836 (N_6836,N_6691,N_6627);
xnor U6837 (N_6837,N_6604,N_6685);
and U6838 (N_6838,N_6688,N_6641);
or U6839 (N_6839,N_6662,N_6706);
nand U6840 (N_6840,N_6662,N_6613);
and U6841 (N_6841,N_6689,N_6612);
and U6842 (N_6842,N_6722,N_6738);
and U6843 (N_6843,N_6632,N_6657);
xnor U6844 (N_6844,N_6641,N_6648);
nand U6845 (N_6845,N_6736,N_6670);
xnor U6846 (N_6846,N_6720,N_6686);
nand U6847 (N_6847,N_6624,N_6662);
nor U6848 (N_6848,N_6676,N_6710);
nor U6849 (N_6849,N_6658,N_6624);
nand U6850 (N_6850,N_6706,N_6693);
xnor U6851 (N_6851,N_6670,N_6647);
or U6852 (N_6852,N_6651,N_6633);
xor U6853 (N_6853,N_6727,N_6746);
xnor U6854 (N_6854,N_6695,N_6642);
or U6855 (N_6855,N_6665,N_6676);
or U6856 (N_6856,N_6671,N_6614);
nand U6857 (N_6857,N_6747,N_6688);
nor U6858 (N_6858,N_6738,N_6701);
xnor U6859 (N_6859,N_6612,N_6639);
xnor U6860 (N_6860,N_6652,N_6665);
xnor U6861 (N_6861,N_6652,N_6655);
or U6862 (N_6862,N_6632,N_6721);
or U6863 (N_6863,N_6733,N_6665);
and U6864 (N_6864,N_6639,N_6660);
or U6865 (N_6865,N_6625,N_6743);
and U6866 (N_6866,N_6709,N_6671);
nor U6867 (N_6867,N_6638,N_6690);
nand U6868 (N_6868,N_6676,N_6611);
or U6869 (N_6869,N_6623,N_6749);
nor U6870 (N_6870,N_6741,N_6717);
nand U6871 (N_6871,N_6624,N_6692);
nand U6872 (N_6872,N_6687,N_6680);
and U6873 (N_6873,N_6711,N_6634);
or U6874 (N_6874,N_6747,N_6722);
xnor U6875 (N_6875,N_6706,N_6641);
or U6876 (N_6876,N_6613,N_6667);
nand U6877 (N_6877,N_6679,N_6744);
or U6878 (N_6878,N_6637,N_6631);
or U6879 (N_6879,N_6676,N_6718);
and U6880 (N_6880,N_6734,N_6694);
nor U6881 (N_6881,N_6698,N_6669);
xnor U6882 (N_6882,N_6626,N_6638);
nand U6883 (N_6883,N_6644,N_6666);
nor U6884 (N_6884,N_6657,N_6698);
nand U6885 (N_6885,N_6738,N_6636);
and U6886 (N_6886,N_6609,N_6712);
and U6887 (N_6887,N_6645,N_6721);
xor U6888 (N_6888,N_6624,N_6711);
or U6889 (N_6889,N_6653,N_6713);
xnor U6890 (N_6890,N_6728,N_6727);
xnor U6891 (N_6891,N_6726,N_6663);
nand U6892 (N_6892,N_6674,N_6717);
or U6893 (N_6893,N_6661,N_6639);
and U6894 (N_6894,N_6736,N_6626);
nor U6895 (N_6895,N_6708,N_6693);
xnor U6896 (N_6896,N_6711,N_6606);
and U6897 (N_6897,N_6695,N_6618);
or U6898 (N_6898,N_6633,N_6714);
nand U6899 (N_6899,N_6700,N_6630);
xnor U6900 (N_6900,N_6770,N_6799);
or U6901 (N_6901,N_6865,N_6824);
or U6902 (N_6902,N_6812,N_6878);
xor U6903 (N_6903,N_6875,N_6897);
or U6904 (N_6904,N_6795,N_6800);
or U6905 (N_6905,N_6874,N_6821);
or U6906 (N_6906,N_6898,N_6818);
or U6907 (N_6907,N_6850,N_6860);
nor U6908 (N_6908,N_6755,N_6830);
nand U6909 (N_6909,N_6788,N_6872);
and U6910 (N_6910,N_6817,N_6787);
xnor U6911 (N_6911,N_6884,N_6814);
or U6912 (N_6912,N_6801,N_6791);
or U6913 (N_6913,N_6892,N_6804);
or U6914 (N_6914,N_6774,N_6880);
and U6915 (N_6915,N_6782,N_6815);
and U6916 (N_6916,N_6851,N_6762);
and U6917 (N_6917,N_6843,N_6848);
and U6918 (N_6918,N_6772,N_6854);
xor U6919 (N_6919,N_6802,N_6834);
nor U6920 (N_6920,N_6823,N_6783);
or U6921 (N_6921,N_6803,N_6837);
nor U6922 (N_6922,N_6887,N_6869);
nor U6923 (N_6923,N_6857,N_6871);
and U6924 (N_6924,N_6882,N_6894);
and U6925 (N_6925,N_6816,N_6856);
or U6926 (N_6926,N_6893,N_6763);
nand U6927 (N_6927,N_6833,N_6750);
nand U6928 (N_6928,N_6790,N_6813);
and U6929 (N_6929,N_6861,N_6859);
or U6930 (N_6930,N_6792,N_6853);
or U6931 (N_6931,N_6771,N_6768);
xor U6932 (N_6932,N_6798,N_6873);
nand U6933 (N_6933,N_6844,N_6852);
and U6934 (N_6934,N_6888,N_6810);
nand U6935 (N_6935,N_6806,N_6849);
xnor U6936 (N_6936,N_6879,N_6855);
and U6937 (N_6937,N_6819,N_6753);
and U6938 (N_6938,N_6838,N_6896);
nand U6939 (N_6939,N_6769,N_6870);
nor U6940 (N_6940,N_6796,N_6883);
nor U6941 (N_6941,N_6751,N_6826);
nand U6942 (N_6942,N_6839,N_6758);
nor U6943 (N_6943,N_6847,N_6846);
xor U6944 (N_6944,N_6864,N_6807);
xnor U6945 (N_6945,N_6862,N_6775);
nor U6946 (N_6946,N_6876,N_6842);
xor U6947 (N_6947,N_6794,N_6828);
or U6948 (N_6948,N_6841,N_6778);
nand U6949 (N_6949,N_6895,N_6756);
nor U6950 (N_6950,N_6899,N_6845);
and U6951 (N_6951,N_6877,N_6827);
nand U6952 (N_6952,N_6780,N_6829);
xor U6953 (N_6953,N_6831,N_6766);
nand U6954 (N_6954,N_6776,N_6797);
xor U6955 (N_6955,N_6760,N_6757);
xor U6956 (N_6956,N_6789,N_6805);
xnor U6957 (N_6957,N_6890,N_6811);
nor U6958 (N_6958,N_6773,N_6808);
or U6959 (N_6959,N_6765,N_6858);
xor U6960 (N_6960,N_6863,N_6784);
nand U6961 (N_6961,N_6786,N_6822);
and U6962 (N_6962,N_6891,N_6761);
nor U6963 (N_6963,N_6881,N_6825);
xnor U6964 (N_6964,N_6809,N_6767);
nor U6965 (N_6965,N_6868,N_6867);
nand U6966 (N_6966,N_6886,N_6820);
nand U6967 (N_6967,N_6754,N_6889);
and U6968 (N_6968,N_6866,N_6840);
nand U6969 (N_6969,N_6777,N_6785);
xor U6970 (N_6970,N_6836,N_6764);
and U6971 (N_6971,N_6781,N_6779);
or U6972 (N_6972,N_6832,N_6759);
or U6973 (N_6973,N_6752,N_6885);
or U6974 (N_6974,N_6835,N_6793);
xnor U6975 (N_6975,N_6791,N_6770);
and U6976 (N_6976,N_6838,N_6890);
and U6977 (N_6977,N_6863,N_6890);
nand U6978 (N_6978,N_6786,N_6761);
or U6979 (N_6979,N_6812,N_6784);
xnor U6980 (N_6980,N_6843,N_6760);
and U6981 (N_6981,N_6789,N_6769);
and U6982 (N_6982,N_6830,N_6785);
nor U6983 (N_6983,N_6791,N_6852);
xor U6984 (N_6984,N_6756,N_6881);
xor U6985 (N_6985,N_6772,N_6806);
nor U6986 (N_6986,N_6872,N_6789);
nand U6987 (N_6987,N_6871,N_6778);
nand U6988 (N_6988,N_6850,N_6757);
and U6989 (N_6989,N_6897,N_6775);
nor U6990 (N_6990,N_6838,N_6808);
nand U6991 (N_6991,N_6875,N_6867);
and U6992 (N_6992,N_6798,N_6779);
nor U6993 (N_6993,N_6766,N_6834);
xnor U6994 (N_6994,N_6849,N_6851);
and U6995 (N_6995,N_6765,N_6775);
or U6996 (N_6996,N_6785,N_6764);
or U6997 (N_6997,N_6779,N_6806);
nor U6998 (N_6998,N_6863,N_6895);
xor U6999 (N_6999,N_6798,N_6801);
and U7000 (N_7000,N_6826,N_6874);
xor U7001 (N_7001,N_6800,N_6867);
nor U7002 (N_7002,N_6875,N_6812);
xor U7003 (N_7003,N_6841,N_6885);
and U7004 (N_7004,N_6764,N_6838);
nor U7005 (N_7005,N_6779,N_6897);
and U7006 (N_7006,N_6840,N_6753);
or U7007 (N_7007,N_6778,N_6849);
nor U7008 (N_7008,N_6868,N_6802);
or U7009 (N_7009,N_6872,N_6806);
and U7010 (N_7010,N_6761,N_6861);
nand U7011 (N_7011,N_6803,N_6854);
nor U7012 (N_7012,N_6846,N_6815);
nand U7013 (N_7013,N_6818,N_6872);
nor U7014 (N_7014,N_6829,N_6785);
and U7015 (N_7015,N_6866,N_6793);
or U7016 (N_7016,N_6792,N_6790);
nor U7017 (N_7017,N_6825,N_6857);
nand U7018 (N_7018,N_6822,N_6890);
and U7019 (N_7019,N_6802,N_6791);
nand U7020 (N_7020,N_6817,N_6819);
xnor U7021 (N_7021,N_6832,N_6880);
xor U7022 (N_7022,N_6877,N_6790);
and U7023 (N_7023,N_6882,N_6761);
and U7024 (N_7024,N_6891,N_6812);
or U7025 (N_7025,N_6868,N_6810);
nor U7026 (N_7026,N_6758,N_6823);
xnor U7027 (N_7027,N_6820,N_6862);
or U7028 (N_7028,N_6843,N_6757);
or U7029 (N_7029,N_6790,N_6801);
xor U7030 (N_7030,N_6850,N_6887);
nor U7031 (N_7031,N_6808,N_6854);
or U7032 (N_7032,N_6791,N_6827);
or U7033 (N_7033,N_6833,N_6817);
xor U7034 (N_7034,N_6799,N_6801);
nand U7035 (N_7035,N_6815,N_6819);
nor U7036 (N_7036,N_6783,N_6884);
nand U7037 (N_7037,N_6897,N_6818);
nor U7038 (N_7038,N_6805,N_6862);
nor U7039 (N_7039,N_6880,N_6861);
nor U7040 (N_7040,N_6832,N_6865);
nor U7041 (N_7041,N_6856,N_6887);
nand U7042 (N_7042,N_6895,N_6774);
and U7043 (N_7043,N_6806,N_6793);
nand U7044 (N_7044,N_6754,N_6857);
nor U7045 (N_7045,N_6874,N_6813);
xor U7046 (N_7046,N_6806,N_6802);
or U7047 (N_7047,N_6826,N_6804);
nor U7048 (N_7048,N_6827,N_6859);
xor U7049 (N_7049,N_6751,N_6894);
nand U7050 (N_7050,N_6916,N_6944);
and U7051 (N_7051,N_6975,N_6953);
nand U7052 (N_7052,N_7010,N_6988);
nand U7053 (N_7053,N_7023,N_6937);
xor U7054 (N_7054,N_6989,N_7013);
nand U7055 (N_7055,N_7040,N_7000);
and U7056 (N_7056,N_6904,N_7020);
nand U7057 (N_7057,N_6934,N_6909);
nand U7058 (N_7058,N_6900,N_7034);
nor U7059 (N_7059,N_7044,N_6917);
and U7060 (N_7060,N_7015,N_7012);
nor U7061 (N_7061,N_6921,N_6938);
xnor U7062 (N_7062,N_7024,N_7049);
or U7063 (N_7063,N_7028,N_6979);
or U7064 (N_7064,N_6923,N_6967);
and U7065 (N_7065,N_7048,N_6996);
xor U7066 (N_7066,N_6902,N_6912);
nor U7067 (N_7067,N_6903,N_6964);
nand U7068 (N_7068,N_6971,N_6943);
nor U7069 (N_7069,N_6922,N_7029);
and U7070 (N_7070,N_6957,N_6925);
xnor U7071 (N_7071,N_7041,N_6970);
nor U7072 (N_7072,N_7032,N_6926);
nand U7073 (N_7073,N_6949,N_6920);
nand U7074 (N_7074,N_7045,N_6911);
or U7075 (N_7075,N_7008,N_6982);
nand U7076 (N_7076,N_7019,N_6929);
or U7077 (N_7077,N_6907,N_6969);
nor U7078 (N_7078,N_6993,N_6948);
or U7079 (N_7079,N_6986,N_6994);
xor U7080 (N_7080,N_7030,N_7021);
nand U7081 (N_7081,N_7004,N_6983);
or U7082 (N_7082,N_7037,N_7039);
and U7083 (N_7083,N_7042,N_6991);
or U7084 (N_7084,N_6914,N_6915);
nor U7085 (N_7085,N_7014,N_6950);
xor U7086 (N_7086,N_6960,N_7009);
xor U7087 (N_7087,N_6959,N_6908);
nand U7088 (N_7088,N_6995,N_6997);
xor U7089 (N_7089,N_6998,N_6918);
nor U7090 (N_7090,N_7002,N_6978);
xnor U7091 (N_7091,N_6924,N_7005);
and U7092 (N_7092,N_6933,N_6919);
and U7093 (N_7093,N_6992,N_6977);
or U7094 (N_7094,N_6941,N_7017);
nand U7095 (N_7095,N_7036,N_6942);
nand U7096 (N_7096,N_6961,N_7001);
and U7097 (N_7097,N_6954,N_7016);
nor U7098 (N_7098,N_6952,N_6945);
nand U7099 (N_7099,N_6968,N_6935);
or U7100 (N_7100,N_6974,N_7003);
nand U7101 (N_7101,N_6966,N_7043);
and U7102 (N_7102,N_6965,N_6913);
nor U7103 (N_7103,N_7035,N_6930);
xnor U7104 (N_7104,N_7007,N_7033);
and U7105 (N_7105,N_6946,N_6910);
nand U7106 (N_7106,N_6987,N_6955);
nand U7107 (N_7107,N_7026,N_6976);
or U7108 (N_7108,N_6928,N_6972);
xnor U7109 (N_7109,N_6956,N_6981);
xor U7110 (N_7110,N_7025,N_6936);
or U7111 (N_7111,N_7031,N_6906);
xor U7112 (N_7112,N_6932,N_6990);
nor U7113 (N_7113,N_6962,N_6984);
or U7114 (N_7114,N_7018,N_6939);
or U7115 (N_7115,N_6958,N_6951);
nor U7116 (N_7116,N_6905,N_6999);
or U7117 (N_7117,N_6963,N_6927);
nand U7118 (N_7118,N_6901,N_6973);
or U7119 (N_7119,N_7022,N_7027);
or U7120 (N_7120,N_6947,N_7047);
nor U7121 (N_7121,N_6931,N_7046);
or U7122 (N_7122,N_6985,N_6940);
nor U7123 (N_7123,N_7006,N_7038);
and U7124 (N_7124,N_7011,N_6980);
and U7125 (N_7125,N_6985,N_6944);
and U7126 (N_7126,N_7011,N_6907);
nor U7127 (N_7127,N_6902,N_6940);
and U7128 (N_7128,N_6956,N_6922);
or U7129 (N_7129,N_6982,N_6935);
xor U7130 (N_7130,N_6904,N_6912);
and U7131 (N_7131,N_6925,N_6975);
xnor U7132 (N_7132,N_7031,N_6904);
nor U7133 (N_7133,N_7024,N_6937);
nor U7134 (N_7134,N_6989,N_6984);
xnor U7135 (N_7135,N_7045,N_6998);
xnor U7136 (N_7136,N_6993,N_7019);
xor U7137 (N_7137,N_7022,N_7041);
or U7138 (N_7138,N_7030,N_6950);
nor U7139 (N_7139,N_6908,N_6944);
xor U7140 (N_7140,N_6973,N_7001);
or U7141 (N_7141,N_6990,N_6934);
nor U7142 (N_7142,N_6977,N_6928);
or U7143 (N_7143,N_7011,N_6927);
and U7144 (N_7144,N_7034,N_7049);
nor U7145 (N_7145,N_6936,N_6979);
and U7146 (N_7146,N_7013,N_7009);
or U7147 (N_7147,N_6940,N_6936);
or U7148 (N_7148,N_7042,N_6998);
nand U7149 (N_7149,N_7022,N_6930);
or U7150 (N_7150,N_6922,N_6977);
xnor U7151 (N_7151,N_7038,N_6977);
nor U7152 (N_7152,N_7007,N_7030);
xnor U7153 (N_7153,N_7033,N_6916);
nor U7154 (N_7154,N_6945,N_7008);
nand U7155 (N_7155,N_6912,N_6943);
xor U7156 (N_7156,N_7018,N_6903);
or U7157 (N_7157,N_7047,N_6914);
or U7158 (N_7158,N_6971,N_6916);
nand U7159 (N_7159,N_6915,N_6904);
xnor U7160 (N_7160,N_6959,N_6989);
and U7161 (N_7161,N_6907,N_7044);
or U7162 (N_7162,N_7015,N_6943);
xor U7163 (N_7163,N_6949,N_7029);
or U7164 (N_7164,N_6926,N_6997);
nand U7165 (N_7165,N_6997,N_6908);
and U7166 (N_7166,N_6971,N_7008);
nand U7167 (N_7167,N_6942,N_6922);
and U7168 (N_7168,N_7014,N_7048);
or U7169 (N_7169,N_7008,N_6980);
xnor U7170 (N_7170,N_6917,N_6901);
xor U7171 (N_7171,N_7008,N_7011);
nor U7172 (N_7172,N_6960,N_6925);
nand U7173 (N_7173,N_6919,N_6917);
nor U7174 (N_7174,N_7047,N_6964);
or U7175 (N_7175,N_7046,N_7022);
or U7176 (N_7176,N_6910,N_6967);
and U7177 (N_7177,N_7044,N_7010);
nand U7178 (N_7178,N_6982,N_6904);
and U7179 (N_7179,N_7003,N_6982);
or U7180 (N_7180,N_7040,N_7004);
nand U7181 (N_7181,N_7030,N_6994);
nor U7182 (N_7182,N_7011,N_6995);
or U7183 (N_7183,N_7014,N_7016);
or U7184 (N_7184,N_6976,N_6954);
or U7185 (N_7185,N_7035,N_6983);
nor U7186 (N_7186,N_7049,N_6955);
xnor U7187 (N_7187,N_7024,N_6907);
xnor U7188 (N_7188,N_7022,N_7035);
nand U7189 (N_7189,N_6925,N_6927);
and U7190 (N_7190,N_7049,N_7030);
nor U7191 (N_7191,N_7006,N_6965);
nand U7192 (N_7192,N_7034,N_6920);
nor U7193 (N_7193,N_6971,N_6980);
and U7194 (N_7194,N_7005,N_7030);
xor U7195 (N_7195,N_7035,N_6914);
xor U7196 (N_7196,N_7043,N_6997);
or U7197 (N_7197,N_6966,N_6928);
nand U7198 (N_7198,N_6900,N_6950);
and U7199 (N_7199,N_6967,N_6975);
xor U7200 (N_7200,N_7161,N_7159);
nor U7201 (N_7201,N_7128,N_7174);
or U7202 (N_7202,N_7155,N_7120);
and U7203 (N_7203,N_7181,N_7132);
xnor U7204 (N_7204,N_7093,N_7077);
and U7205 (N_7205,N_7065,N_7136);
nand U7206 (N_7206,N_7169,N_7199);
nand U7207 (N_7207,N_7082,N_7130);
nor U7208 (N_7208,N_7182,N_7061);
nor U7209 (N_7209,N_7156,N_7103);
nor U7210 (N_7210,N_7186,N_7118);
nand U7211 (N_7211,N_7139,N_7151);
or U7212 (N_7212,N_7108,N_7123);
and U7213 (N_7213,N_7055,N_7083);
or U7214 (N_7214,N_7141,N_7196);
and U7215 (N_7215,N_7197,N_7179);
xnor U7216 (N_7216,N_7059,N_7122);
xnor U7217 (N_7217,N_7150,N_7127);
and U7218 (N_7218,N_7165,N_7153);
and U7219 (N_7219,N_7160,N_7111);
xor U7220 (N_7220,N_7146,N_7109);
nor U7221 (N_7221,N_7114,N_7094);
xnor U7222 (N_7222,N_7126,N_7062);
nand U7223 (N_7223,N_7090,N_7064);
nand U7224 (N_7224,N_7068,N_7152);
or U7225 (N_7225,N_7102,N_7084);
nor U7226 (N_7226,N_7138,N_7164);
or U7227 (N_7227,N_7080,N_7135);
nand U7228 (N_7228,N_7148,N_7180);
or U7229 (N_7229,N_7050,N_7106);
nand U7230 (N_7230,N_7175,N_7189);
xor U7231 (N_7231,N_7178,N_7195);
nand U7232 (N_7232,N_7125,N_7137);
and U7233 (N_7233,N_7110,N_7054);
nand U7234 (N_7234,N_7129,N_7154);
xor U7235 (N_7235,N_7113,N_7107);
and U7236 (N_7236,N_7184,N_7134);
nand U7237 (N_7237,N_7071,N_7086);
nor U7238 (N_7238,N_7190,N_7115);
nor U7239 (N_7239,N_7158,N_7099);
xnor U7240 (N_7240,N_7163,N_7142);
nand U7241 (N_7241,N_7192,N_7119);
and U7242 (N_7242,N_7143,N_7170);
nand U7243 (N_7243,N_7052,N_7187);
or U7244 (N_7244,N_7193,N_7176);
xor U7245 (N_7245,N_7124,N_7076);
xor U7246 (N_7246,N_7096,N_7101);
nand U7247 (N_7247,N_7105,N_7104);
nor U7248 (N_7248,N_7177,N_7191);
and U7249 (N_7249,N_7145,N_7168);
nand U7250 (N_7250,N_7053,N_7162);
nand U7251 (N_7251,N_7116,N_7087);
and U7252 (N_7252,N_7100,N_7079);
nand U7253 (N_7253,N_7072,N_7172);
and U7254 (N_7254,N_7185,N_7149);
nand U7255 (N_7255,N_7063,N_7091);
and U7256 (N_7256,N_7121,N_7056);
nor U7257 (N_7257,N_7140,N_7097);
xnor U7258 (N_7258,N_7173,N_7058);
nor U7259 (N_7259,N_7133,N_7131);
nand U7260 (N_7260,N_7081,N_7095);
nor U7261 (N_7261,N_7066,N_7166);
and U7262 (N_7262,N_7073,N_7171);
nand U7263 (N_7263,N_7089,N_7075);
nand U7264 (N_7264,N_7188,N_7098);
or U7265 (N_7265,N_7070,N_7051);
xor U7266 (N_7266,N_7067,N_7060);
nor U7267 (N_7267,N_7112,N_7088);
xor U7268 (N_7268,N_7144,N_7117);
nor U7269 (N_7269,N_7078,N_7074);
and U7270 (N_7270,N_7069,N_7183);
nand U7271 (N_7271,N_7194,N_7167);
xor U7272 (N_7272,N_7147,N_7057);
xnor U7273 (N_7273,N_7085,N_7092);
or U7274 (N_7274,N_7157,N_7198);
and U7275 (N_7275,N_7068,N_7159);
nor U7276 (N_7276,N_7079,N_7111);
and U7277 (N_7277,N_7103,N_7089);
nand U7278 (N_7278,N_7149,N_7102);
nor U7279 (N_7279,N_7087,N_7129);
nor U7280 (N_7280,N_7095,N_7120);
nand U7281 (N_7281,N_7198,N_7135);
xor U7282 (N_7282,N_7105,N_7144);
or U7283 (N_7283,N_7070,N_7084);
and U7284 (N_7284,N_7133,N_7179);
and U7285 (N_7285,N_7125,N_7186);
nand U7286 (N_7286,N_7170,N_7182);
nor U7287 (N_7287,N_7133,N_7092);
nand U7288 (N_7288,N_7199,N_7195);
nor U7289 (N_7289,N_7127,N_7166);
nor U7290 (N_7290,N_7131,N_7163);
nor U7291 (N_7291,N_7181,N_7071);
and U7292 (N_7292,N_7055,N_7191);
or U7293 (N_7293,N_7102,N_7118);
nand U7294 (N_7294,N_7100,N_7109);
or U7295 (N_7295,N_7138,N_7184);
nor U7296 (N_7296,N_7113,N_7188);
xor U7297 (N_7297,N_7093,N_7097);
nor U7298 (N_7298,N_7050,N_7117);
nor U7299 (N_7299,N_7091,N_7098);
nand U7300 (N_7300,N_7143,N_7131);
or U7301 (N_7301,N_7075,N_7095);
nor U7302 (N_7302,N_7063,N_7139);
or U7303 (N_7303,N_7198,N_7111);
xnor U7304 (N_7304,N_7198,N_7103);
nor U7305 (N_7305,N_7120,N_7187);
xnor U7306 (N_7306,N_7056,N_7125);
xor U7307 (N_7307,N_7103,N_7179);
xor U7308 (N_7308,N_7079,N_7119);
nand U7309 (N_7309,N_7056,N_7127);
nand U7310 (N_7310,N_7105,N_7163);
nor U7311 (N_7311,N_7051,N_7196);
xor U7312 (N_7312,N_7060,N_7103);
nor U7313 (N_7313,N_7173,N_7100);
nor U7314 (N_7314,N_7166,N_7087);
nor U7315 (N_7315,N_7051,N_7152);
or U7316 (N_7316,N_7161,N_7079);
nor U7317 (N_7317,N_7066,N_7174);
nor U7318 (N_7318,N_7124,N_7119);
xnor U7319 (N_7319,N_7170,N_7184);
nor U7320 (N_7320,N_7126,N_7085);
nor U7321 (N_7321,N_7184,N_7085);
xnor U7322 (N_7322,N_7093,N_7095);
or U7323 (N_7323,N_7089,N_7183);
xor U7324 (N_7324,N_7176,N_7076);
or U7325 (N_7325,N_7096,N_7193);
nor U7326 (N_7326,N_7198,N_7146);
and U7327 (N_7327,N_7173,N_7128);
and U7328 (N_7328,N_7091,N_7067);
nor U7329 (N_7329,N_7187,N_7158);
nor U7330 (N_7330,N_7121,N_7196);
or U7331 (N_7331,N_7142,N_7109);
nand U7332 (N_7332,N_7085,N_7105);
nand U7333 (N_7333,N_7119,N_7136);
or U7334 (N_7334,N_7088,N_7145);
nand U7335 (N_7335,N_7137,N_7181);
or U7336 (N_7336,N_7103,N_7144);
and U7337 (N_7337,N_7063,N_7148);
and U7338 (N_7338,N_7180,N_7091);
nor U7339 (N_7339,N_7050,N_7079);
xnor U7340 (N_7340,N_7196,N_7120);
or U7341 (N_7341,N_7162,N_7199);
nand U7342 (N_7342,N_7115,N_7176);
nand U7343 (N_7343,N_7108,N_7084);
nand U7344 (N_7344,N_7106,N_7081);
and U7345 (N_7345,N_7089,N_7158);
or U7346 (N_7346,N_7086,N_7089);
and U7347 (N_7347,N_7087,N_7187);
or U7348 (N_7348,N_7153,N_7152);
and U7349 (N_7349,N_7091,N_7155);
nor U7350 (N_7350,N_7286,N_7271);
xnor U7351 (N_7351,N_7246,N_7276);
and U7352 (N_7352,N_7258,N_7346);
nand U7353 (N_7353,N_7214,N_7227);
nand U7354 (N_7354,N_7277,N_7248);
and U7355 (N_7355,N_7342,N_7218);
xnor U7356 (N_7356,N_7280,N_7201);
xor U7357 (N_7357,N_7267,N_7344);
nor U7358 (N_7358,N_7299,N_7306);
nand U7359 (N_7359,N_7341,N_7327);
or U7360 (N_7360,N_7325,N_7295);
nor U7361 (N_7361,N_7297,N_7230);
nor U7362 (N_7362,N_7207,N_7251);
or U7363 (N_7363,N_7308,N_7323);
xor U7364 (N_7364,N_7238,N_7321);
and U7365 (N_7365,N_7289,N_7270);
and U7366 (N_7366,N_7339,N_7303);
nor U7367 (N_7367,N_7264,N_7311);
nand U7368 (N_7368,N_7283,N_7334);
or U7369 (N_7369,N_7343,N_7333);
xnor U7370 (N_7370,N_7210,N_7300);
xor U7371 (N_7371,N_7256,N_7222);
or U7372 (N_7372,N_7241,N_7310);
nor U7373 (N_7373,N_7205,N_7242);
xnor U7374 (N_7374,N_7260,N_7335);
nand U7375 (N_7375,N_7348,N_7292);
xnor U7376 (N_7376,N_7340,N_7221);
nand U7377 (N_7377,N_7253,N_7225);
xor U7378 (N_7378,N_7208,N_7275);
nor U7379 (N_7379,N_7349,N_7212);
or U7380 (N_7380,N_7245,N_7228);
xnor U7381 (N_7381,N_7204,N_7269);
nor U7382 (N_7382,N_7324,N_7320);
or U7383 (N_7383,N_7200,N_7237);
xor U7384 (N_7384,N_7274,N_7226);
xor U7385 (N_7385,N_7291,N_7317);
nor U7386 (N_7386,N_7290,N_7298);
xor U7387 (N_7387,N_7247,N_7250);
nor U7388 (N_7388,N_7252,N_7312);
and U7389 (N_7389,N_7233,N_7314);
nor U7390 (N_7390,N_7345,N_7203);
nand U7391 (N_7391,N_7316,N_7272);
nand U7392 (N_7392,N_7304,N_7281);
xnor U7393 (N_7393,N_7288,N_7209);
xnor U7394 (N_7394,N_7268,N_7337);
nand U7395 (N_7395,N_7217,N_7229);
nor U7396 (N_7396,N_7254,N_7347);
or U7397 (N_7397,N_7234,N_7223);
nor U7398 (N_7398,N_7315,N_7261);
or U7399 (N_7399,N_7224,N_7328);
nor U7400 (N_7400,N_7338,N_7326);
nand U7401 (N_7401,N_7236,N_7206);
nor U7402 (N_7402,N_7243,N_7319);
xnor U7403 (N_7403,N_7257,N_7282);
or U7404 (N_7404,N_7331,N_7284);
nor U7405 (N_7405,N_7285,N_7235);
or U7406 (N_7406,N_7330,N_7231);
and U7407 (N_7407,N_7313,N_7262);
or U7408 (N_7408,N_7202,N_7336);
nor U7409 (N_7409,N_7302,N_7279);
nand U7410 (N_7410,N_7332,N_7215);
xor U7411 (N_7411,N_7219,N_7301);
nand U7412 (N_7412,N_7296,N_7259);
nand U7413 (N_7413,N_7322,N_7220);
nand U7414 (N_7414,N_7249,N_7213);
nor U7415 (N_7415,N_7244,N_7273);
and U7416 (N_7416,N_7266,N_7278);
and U7417 (N_7417,N_7211,N_7232);
nand U7418 (N_7418,N_7263,N_7307);
or U7419 (N_7419,N_7216,N_7305);
xnor U7420 (N_7420,N_7293,N_7294);
or U7421 (N_7421,N_7240,N_7265);
or U7422 (N_7422,N_7318,N_7309);
nand U7423 (N_7423,N_7255,N_7287);
and U7424 (N_7424,N_7239,N_7329);
xor U7425 (N_7425,N_7290,N_7291);
nand U7426 (N_7426,N_7343,N_7250);
or U7427 (N_7427,N_7267,N_7258);
or U7428 (N_7428,N_7304,N_7258);
nor U7429 (N_7429,N_7281,N_7233);
and U7430 (N_7430,N_7274,N_7239);
xor U7431 (N_7431,N_7340,N_7349);
nor U7432 (N_7432,N_7274,N_7242);
xor U7433 (N_7433,N_7304,N_7320);
nand U7434 (N_7434,N_7306,N_7228);
nand U7435 (N_7435,N_7344,N_7329);
nand U7436 (N_7436,N_7223,N_7318);
nor U7437 (N_7437,N_7319,N_7223);
xnor U7438 (N_7438,N_7247,N_7212);
xor U7439 (N_7439,N_7308,N_7222);
nand U7440 (N_7440,N_7266,N_7348);
or U7441 (N_7441,N_7245,N_7215);
nand U7442 (N_7442,N_7299,N_7302);
nor U7443 (N_7443,N_7336,N_7290);
and U7444 (N_7444,N_7250,N_7338);
nand U7445 (N_7445,N_7219,N_7237);
nor U7446 (N_7446,N_7262,N_7326);
nor U7447 (N_7447,N_7215,N_7283);
and U7448 (N_7448,N_7326,N_7309);
or U7449 (N_7449,N_7216,N_7279);
xor U7450 (N_7450,N_7234,N_7248);
and U7451 (N_7451,N_7331,N_7247);
nor U7452 (N_7452,N_7233,N_7299);
nand U7453 (N_7453,N_7325,N_7336);
xor U7454 (N_7454,N_7257,N_7342);
xor U7455 (N_7455,N_7264,N_7243);
or U7456 (N_7456,N_7288,N_7200);
xor U7457 (N_7457,N_7231,N_7203);
nor U7458 (N_7458,N_7275,N_7337);
or U7459 (N_7459,N_7243,N_7312);
or U7460 (N_7460,N_7336,N_7217);
nor U7461 (N_7461,N_7280,N_7274);
nand U7462 (N_7462,N_7287,N_7206);
and U7463 (N_7463,N_7342,N_7247);
nor U7464 (N_7464,N_7347,N_7301);
nand U7465 (N_7465,N_7227,N_7315);
and U7466 (N_7466,N_7334,N_7276);
nor U7467 (N_7467,N_7241,N_7275);
xor U7468 (N_7468,N_7240,N_7254);
or U7469 (N_7469,N_7223,N_7242);
and U7470 (N_7470,N_7200,N_7208);
and U7471 (N_7471,N_7275,N_7256);
nand U7472 (N_7472,N_7287,N_7316);
and U7473 (N_7473,N_7310,N_7289);
nor U7474 (N_7474,N_7339,N_7225);
nand U7475 (N_7475,N_7286,N_7326);
nand U7476 (N_7476,N_7299,N_7203);
and U7477 (N_7477,N_7265,N_7327);
xor U7478 (N_7478,N_7212,N_7225);
nand U7479 (N_7479,N_7243,N_7263);
nor U7480 (N_7480,N_7299,N_7242);
or U7481 (N_7481,N_7276,N_7207);
or U7482 (N_7482,N_7253,N_7238);
nand U7483 (N_7483,N_7345,N_7318);
xnor U7484 (N_7484,N_7291,N_7225);
nand U7485 (N_7485,N_7254,N_7332);
nor U7486 (N_7486,N_7288,N_7218);
or U7487 (N_7487,N_7307,N_7203);
or U7488 (N_7488,N_7298,N_7222);
nand U7489 (N_7489,N_7232,N_7234);
and U7490 (N_7490,N_7289,N_7278);
and U7491 (N_7491,N_7314,N_7337);
nand U7492 (N_7492,N_7321,N_7273);
or U7493 (N_7493,N_7230,N_7329);
nor U7494 (N_7494,N_7205,N_7222);
or U7495 (N_7495,N_7232,N_7312);
and U7496 (N_7496,N_7218,N_7314);
and U7497 (N_7497,N_7289,N_7311);
xor U7498 (N_7498,N_7294,N_7321);
nor U7499 (N_7499,N_7244,N_7306);
and U7500 (N_7500,N_7417,N_7406);
xor U7501 (N_7501,N_7407,N_7498);
nor U7502 (N_7502,N_7422,N_7399);
and U7503 (N_7503,N_7429,N_7355);
xor U7504 (N_7504,N_7435,N_7387);
nor U7505 (N_7505,N_7472,N_7494);
nand U7506 (N_7506,N_7461,N_7386);
and U7507 (N_7507,N_7431,N_7479);
nor U7508 (N_7508,N_7467,N_7362);
nor U7509 (N_7509,N_7454,N_7482);
nor U7510 (N_7510,N_7361,N_7395);
and U7511 (N_7511,N_7449,N_7425);
or U7512 (N_7512,N_7483,N_7463);
nand U7513 (N_7513,N_7353,N_7490);
and U7514 (N_7514,N_7396,N_7432);
and U7515 (N_7515,N_7476,N_7426);
xnor U7516 (N_7516,N_7363,N_7377);
or U7517 (N_7517,N_7404,N_7354);
nand U7518 (N_7518,N_7402,N_7487);
nand U7519 (N_7519,N_7452,N_7365);
nand U7520 (N_7520,N_7364,N_7375);
or U7521 (N_7521,N_7484,N_7455);
xor U7522 (N_7522,N_7409,N_7456);
nand U7523 (N_7523,N_7421,N_7424);
nor U7524 (N_7524,N_7414,N_7356);
or U7525 (N_7525,N_7410,N_7478);
nor U7526 (N_7526,N_7489,N_7371);
and U7527 (N_7527,N_7372,N_7496);
nor U7528 (N_7528,N_7408,N_7445);
xnor U7529 (N_7529,N_7428,N_7420);
and U7530 (N_7530,N_7480,N_7469);
xnor U7531 (N_7531,N_7499,N_7464);
and U7532 (N_7532,N_7351,N_7473);
nand U7533 (N_7533,N_7470,N_7439);
nor U7534 (N_7534,N_7369,N_7357);
nand U7535 (N_7535,N_7442,N_7401);
nand U7536 (N_7536,N_7416,N_7376);
nor U7537 (N_7537,N_7380,N_7388);
xor U7538 (N_7538,N_7397,N_7415);
and U7539 (N_7539,N_7444,N_7443);
or U7540 (N_7540,N_7413,N_7418);
or U7541 (N_7541,N_7419,N_7385);
and U7542 (N_7542,N_7405,N_7358);
xnor U7543 (N_7543,N_7468,N_7441);
or U7544 (N_7544,N_7379,N_7368);
xor U7545 (N_7545,N_7446,N_7488);
nand U7546 (N_7546,N_7367,N_7438);
nor U7547 (N_7547,N_7350,N_7403);
or U7548 (N_7548,N_7391,N_7453);
and U7549 (N_7549,N_7434,N_7366);
nor U7550 (N_7550,N_7450,N_7466);
nand U7551 (N_7551,N_7411,N_7474);
or U7552 (N_7552,N_7477,N_7392);
xnor U7553 (N_7553,N_7393,N_7491);
and U7554 (N_7554,N_7437,N_7352);
or U7555 (N_7555,N_7384,N_7400);
nor U7556 (N_7556,N_7370,N_7373);
nand U7557 (N_7557,N_7430,N_7390);
nand U7558 (N_7558,N_7459,N_7495);
or U7559 (N_7559,N_7433,N_7378);
and U7560 (N_7560,N_7436,N_7475);
or U7561 (N_7561,N_7382,N_7460);
or U7562 (N_7562,N_7493,N_7360);
xnor U7563 (N_7563,N_7485,N_7394);
nand U7564 (N_7564,N_7383,N_7359);
and U7565 (N_7565,N_7492,N_7462);
xor U7566 (N_7566,N_7447,N_7481);
and U7567 (N_7567,N_7440,N_7412);
nor U7568 (N_7568,N_7471,N_7457);
or U7569 (N_7569,N_7423,N_7458);
nor U7570 (N_7570,N_7451,N_7486);
xor U7571 (N_7571,N_7398,N_7427);
nor U7572 (N_7572,N_7389,N_7381);
nor U7573 (N_7573,N_7465,N_7448);
or U7574 (N_7574,N_7497,N_7374);
xor U7575 (N_7575,N_7442,N_7386);
nand U7576 (N_7576,N_7386,N_7397);
and U7577 (N_7577,N_7388,N_7456);
xor U7578 (N_7578,N_7362,N_7455);
nor U7579 (N_7579,N_7485,N_7388);
and U7580 (N_7580,N_7363,N_7488);
nand U7581 (N_7581,N_7356,N_7380);
nand U7582 (N_7582,N_7410,N_7420);
and U7583 (N_7583,N_7482,N_7426);
xor U7584 (N_7584,N_7356,N_7411);
nand U7585 (N_7585,N_7355,N_7465);
nor U7586 (N_7586,N_7376,N_7425);
nor U7587 (N_7587,N_7476,N_7496);
and U7588 (N_7588,N_7408,N_7478);
nor U7589 (N_7589,N_7418,N_7463);
or U7590 (N_7590,N_7411,N_7371);
and U7591 (N_7591,N_7490,N_7434);
xnor U7592 (N_7592,N_7356,N_7497);
and U7593 (N_7593,N_7353,N_7360);
xor U7594 (N_7594,N_7476,N_7403);
nor U7595 (N_7595,N_7363,N_7491);
or U7596 (N_7596,N_7425,N_7459);
nor U7597 (N_7597,N_7417,N_7495);
nor U7598 (N_7598,N_7473,N_7363);
and U7599 (N_7599,N_7381,N_7416);
nor U7600 (N_7600,N_7418,N_7431);
nor U7601 (N_7601,N_7435,N_7431);
or U7602 (N_7602,N_7428,N_7413);
and U7603 (N_7603,N_7484,N_7417);
or U7604 (N_7604,N_7487,N_7437);
xnor U7605 (N_7605,N_7367,N_7475);
xor U7606 (N_7606,N_7481,N_7370);
nand U7607 (N_7607,N_7378,N_7354);
nand U7608 (N_7608,N_7446,N_7487);
nor U7609 (N_7609,N_7461,N_7397);
nand U7610 (N_7610,N_7470,N_7475);
xor U7611 (N_7611,N_7401,N_7465);
nand U7612 (N_7612,N_7439,N_7360);
or U7613 (N_7613,N_7492,N_7440);
or U7614 (N_7614,N_7411,N_7465);
xnor U7615 (N_7615,N_7416,N_7434);
xor U7616 (N_7616,N_7476,N_7368);
nor U7617 (N_7617,N_7447,N_7436);
and U7618 (N_7618,N_7464,N_7372);
nand U7619 (N_7619,N_7388,N_7453);
and U7620 (N_7620,N_7491,N_7406);
nand U7621 (N_7621,N_7428,N_7385);
and U7622 (N_7622,N_7387,N_7399);
or U7623 (N_7623,N_7416,N_7488);
and U7624 (N_7624,N_7369,N_7439);
xor U7625 (N_7625,N_7473,N_7474);
nor U7626 (N_7626,N_7474,N_7467);
nand U7627 (N_7627,N_7498,N_7404);
nand U7628 (N_7628,N_7447,N_7458);
xor U7629 (N_7629,N_7480,N_7380);
xor U7630 (N_7630,N_7364,N_7382);
and U7631 (N_7631,N_7402,N_7362);
xnor U7632 (N_7632,N_7443,N_7453);
and U7633 (N_7633,N_7474,N_7463);
nor U7634 (N_7634,N_7373,N_7364);
xor U7635 (N_7635,N_7470,N_7479);
xor U7636 (N_7636,N_7455,N_7411);
and U7637 (N_7637,N_7403,N_7398);
and U7638 (N_7638,N_7394,N_7437);
nor U7639 (N_7639,N_7493,N_7463);
nor U7640 (N_7640,N_7469,N_7468);
nand U7641 (N_7641,N_7485,N_7439);
nand U7642 (N_7642,N_7474,N_7468);
and U7643 (N_7643,N_7497,N_7465);
nor U7644 (N_7644,N_7463,N_7371);
and U7645 (N_7645,N_7358,N_7417);
xor U7646 (N_7646,N_7356,N_7405);
xor U7647 (N_7647,N_7362,N_7469);
nor U7648 (N_7648,N_7353,N_7414);
xnor U7649 (N_7649,N_7446,N_7376);
xnor U7650 (N_7650,N_7570,N_7550);
nor U7651 (N_7651,N_7625,N_7605);
and U7652 (N_7652,N_7639,N_7514);
and U7653 (N_7653,N_7631,N_7532);
nand U7654 (N_7654,N_7596,N_7610);
nand U7655 (N_7655,N_7540,N_7559);
xnor U7656 (N_7656,N_7568,N_7529);
nand U7657 (N_7657,N_7548,N_7607);
nand U7658 (N_7658,N_7551,N_7600);
nand U7659 (N_7659,N_7508,N_7587);
nand U7660 (N_7660,N_7504,N_7592);
or U7661 (N_7661,N_7593,N_7516);
nand U7662 (N_7662,N_7512,N_7555);
xnor U7663 (N_7663,N_7640,N_7583);
nand U7664 (N_7664,N_7599,N_7606);
and U7665 (N_7665,N_7575,N_7580);
nor U7666 (N_7666,N_7531,N_7547);
nor U7667 (N_7667,N_7623,N_7609);
xor U7668 (N_7668,N_7616,N_7546);
nor U7669 (N_7669,N_7538,N_7553);
nand U7670 (N_7670,N_7620,N_7515);
or U7671 (N_7671,N_7632,N_7564);
xor U7672 (N_7672,N_7535,N_7643);
nor U7673 (N_7673,N_7542,N_7622);
xnor U7674 (N_7674,N_7595,N_7597);
xor U7675 (N_7675,N_7524,N_7619);
or U7676 (N_7676,N_7577,N_7584);
and U7677 (N_7677,N_7520,N_7558);
nand U7678 (N_7678,N_7633,N_7604);
or U7679 (N_7679,N_7526,N_7528);
and U7680 (N_7680,N_7608,N_7505);
nand U7681 (N_7681,N_7556,N_7521);
nand U7682 (N_7682,N_7522,N_7573);
nor U7683 (N_7683,N_7603,N_7557);
nor U7684 (N_7684,N_7509,N_7590);
and U7685 (N_7685,N_7624,N_7510);
nand U7686 (N_7686,N_7598,N_7541);
or U7687 (N_7687,N_7560,N_7567);
nand U7688 (N_7688,N_7585,N_7636);
or U7689 (N_7689,N_7615,N_7626);
or U7690 (N_7690,N_7602,N_7578);
or U7691 (N_7691,N_7549,N_7612);
xor U7692 (N_7692,N_7519,N_7617);
nor U7693 (N_7693,N_7637,N_7507);
nand U7694 (N_7694,N_7635,N_7565);
or U7695 (N_7695,N_7601,N_7646);
nand U7696 (N_7696,N_7534,N_7642);
or U7697 (N_7697,N_7647,N_7500);
nand U7698 (N_7698,N_7611,N_7571);
nand U7699 (N_7699,N_7630,N_7591);
xnor U7700 (N_7700,N_7561,N_7627);
nor U7701 (N_7701,N_7649,N_7543);
xor U7702 (N_7702,N_7566,N_7586);
xor U7703 (N_7703,N_7648,N_7644);
nor U7704 (N_7704,N_7563,N_7523);
xor U7705 (N_7705,N_7594,N_7506);
or U7706 (N_7706,N_7618,N_7518);
and U7707 (N_7707,N_7621,N_7562);
or U7708 (N_7708,N_7634,N_7539);
and U7709 (N_7709,N_7579,N_7525);
and U7710 (N_7710,N_7545,N_7581);
or U7711 (N_7711,N_7582,N_7614);
xnor U7712 (N_7712,N_7574,N_7513);
and U7713 (N_7713,N_7501,N_7572);
or U7714 (N_7714,N_7588,N_7536);
or U7715 (N_7715,N_7544,N_7537);
xnor U7716 (N_7716,N_7554,N_7629);
nand U7717 (N_7717,N_7641,N_7511);
nand U7718 (N_7718,N_7589,N_7552);
xnor U7719 (N_7719,N_7527,N_7569);
or U7720 (N_7720,N_7638,N_7503);
or U7721 (N_7721,N_7613,N_7530);
xnor U7722 (N_7722,N_7533,N_7517);
xor U7723 (N_7723,N_7628,N_7645);
nand U7724 (N_7724,N_7576,N_7502);
nand U7725 (N_7725,N_7522,N_7562);
nor U7726 (N_7726,N_7568,N_7634);
and U7727 (N_7727,N_7553,N_7565);
nor U7728 (N_7728,N_7521,N_7516);
nand U7729 (N_7729,N_7521,N_7605);
xor U7730 (N_7730,N_7507,N_7577);
nor U7731 (N_7731,N_7530,N_7500);
or U7732 (N_7732,N_7602,N_7582);
or U7733 (N_7733,N_7588,N_7510);
nor U7734 (N_7734,N_7633,N_7562);
nand U7735 (N_7735,N_7628,N_7527);
nor U7736 (N_7736,N_7531,N_7561);
or U7737 (N_7737,N_7636,N_7591);
and U7738 (N_7738,N_7525,N_7531);
xnor U7739 (N_7739,N_7513,N_7581);
nor U7740 (N_7740,N_7520,N_7635);
nor U7741 (N_7741,N_7644,N_7565);
nor U7742 (N_7742,N_7542,N_7525);
nor U7743 (N_7743,N_7623,N_7549);
or U7744 (N_7744,N_7648,N_7580);
nand U7745 (N_7745,N_7544,N_7616);
or U7746 (N_7746,N_7520,N_7511);
and U7747 (N_7747,N_7634,N_7550);
or U7748 (N_7748,N_7556,N_7554);
or U7749 (N_7749,N_7506,N_7554);
and U7750 (N_7750,N_7537,N_7518);
xnor U7751 (N_7751,N_7556,N_7587);
or U7752 (N_7752,N_7553,N_7552);
or U7753 (N_7753,N_7568,N_7628);
and U7754 (N_7754,N_7649,N_7563);
or U7755 (N_7755,N_7631,N_7595);
or U7756 (N_7756,N_7576,N_7613);
xor U7757 (N_7757,N_7645,N_7518);
or U7758 (N_7758,N_7609,N_7599);
nor U7759 (N_7759,N_7526,N_7633);
or U7760 (N_7760,N_7601,N_7599);
xnor U7761 (N_7761,N_7536,N_7623);
xor U7762 (N_7762,N_7634,N_7649);
or U7763 (N_7763,N_7553,N_7545);
nand U7764 (N_7764,N_7519,N_7500);
nand U7765 (N_7765,N_7507,N_7581);
nand U7766 (N_7766,N_7515,N_7600);
or U7767 (N_7767,N_7556,N_7581);
nor U7768 (N_7768,N_7535,N_7533);
and U7769 (N_7769,N_7527,N_7593);
xor U7770 (N_7770,N_7612,N_7596);
xnor U7771 (N_7771,N_7632,N_7548);
nor U7772 (N_7772,N_7558,N_7568);
and U7773 (N_7773,N_7561,N_7519);
or U7774 (N_7774,N_7518,N_7511);
nand U7775 (N_7775,N_7631,N_7551);
nand U7776 (N_7776,N_7513,N_7642);
or U7777 (N_7777,N_7570,N_7618);
or U7778 (N_7778,N_7587,N_7557);
xnor U7779 (N_7779,N_7643,N_7634);
xor U7780 (N_7780,N_7508,N_7532);
or U7781 (N_7781,N_7501,N_7503);
nor U7782 (N_7782,N_7521,N_7597);
xor U7783 (N_7783,N_7626,N_7633);
nor U7784 (N_7784,N_7552,N_7532);
or U7785 (N_7785,N_7633,N_7579);
nand U7786 (N_7786,N_7605,N_7555);
xor U7787 (N_7787,N_7522,N_7549);
nor U7788 (N_7788,N_7500,N_7637);
or U7789 (N_7789,N_7608,N_7576);
nand U7790 (N_7790,N_7647,N_7511);
or U7791 (N_7791,N_7578,N_7571);
nor U7792 (N_7792,N_7565,N_7554);
or U7793 (N_7793,N_7536,N_7533);
or U7794 (N_7794,N_7615,N_7627);
nand U7795 (N_7795,N_7500,N_7548);
or U7796 (N_7796,N_7638,N_7550);
xor U7797 (N_7797,N_7525,N_7611);
xor U7798 (N_7798,N_7524,N_7539);
or U7799 (N_7799,N_7595,N_7574);
and U7800 (N_7800,N_7746,N_7701);
nor U7801 (N_7801,N_7722,N_7744);
or U7802 (N_7802,N_7788,N_7717);
nor U7803 (N_7803,N_7755,N_7707);
nor U7804 (N_7804,N_7778,N_7677);
and U7805 (N_7805,N_7691,N_7670);
and U7806 (N_7806,N_7723,N_7681);
nand U7807 (N_7807,N_7745,N_7771);
nor U7808 (N_7808,N_7772,N_7798);
nor U7809 (N_7809,N_7713,N_7672);
or U7810 (N_7810,N_7774,N_7768);
xnor U7811 (N_7811,N_7704,N_7665);
nor U7812 (N_7812,N_7775,N_7739);
and U7813 (N_7813,N_7715,N_7763);
or U7814 (N_7814,N_7758,N_7721);
and U7815 (N_7815,N_7796,N_7697);
xnor U7816 (N_7816,N_7655,N_7692);
nand U7817 (N_7817,N_7680,N_7678);
or U7818 (N_7818,N_7792,N_7776);
xnor U7819 (N_7819,N_7671,N_7673);
or U7820 (N_7820,N_7657,N_7695);
nand U7821 (N_7821,N_7685,N_7693);
nand U7822 (N_7822,N_7702,N_7762);
and U7823 (N_7823,N_7716,N_7750);
nor U7824 (N_7824,N_7764,N_7773);
nand U7825 (N_7825,N_7741,N_7689);
nand U7826 (N_7826,N_7783,N_7787);
nor U7827 (N_7827,N_7720,N_7679);
nand U7828 (N_7828,N_7719,N_7690);
or U7829 (N_7829,N_7683,N_7705);
and U7830 (N_7830,N_7786,N_7686);
nor U7831 (N_7831,N_7793,N_7766);
nand U7832 (N_7832,N_7688,N_7740);
nand U7833 (N_7833,N_7724,N_7726);
xnor U7834 (N_7834,N_7727,N_7682);
xnor U7835 (N_7835,N_7652,N_7794);
nor U7836 (N_7836,N_7770,N_7728);
xnor U7837 (N_7837,N_7676,N_7661);
nand U7838 (N_7838,N_7738,N_7760);
nand U7839 (N_7839,N_7732,N_7654);
and U7840 (N_7840,N_7718,N_7754);
and U7841 (N_7841,N_7669,N_7674);
xnor U7842 (N_7842,N_7765,N_7757);
and U7843 (N_7843,N_7658,N_7699);
or U7844 (N_7844,N_7785,N_7790);
and U7845 (N_7845,N_7666,N_7653);
and U7846 (N_7846,N_7698,N_7782);
xnor U7847 (N_7847,N_7662,N_7651);
nor U7848 (N_7848,N_7753,N_7694);
nand U7849 (N_7849,N_7725,N_7664);
nor U7850 (N_7850,N_7761,N_7731);
nor U7851 (N_7851,N_7742,N_7799);
nor U7852 (N_7852,N_7696,N_7729);
nor U7853 (N_7853,N_7756,N_7668);
or U7854 (N_7854,N_7769,N_7712);
nor U7855 (N_7855,N_7733,N_7747);
or U7856 (N_7856,N_7650,N_7791);
nand U7857 (N_7857,N_7734,N_7737);
xor U7858 (N_7858,N_7667,N_7789);
xnor U7859 (N_7859,N_7706,N_7743);
or U7860 (N_7860,N_7730,N_7781);
nor U7861 (N_7861,N_7759,N_7777);
nor U7862 (N_7862,N_7660,N_7709);
or U7863 (N_7863,N_7687,N_7784);
nor U7864 (N_7864,N_7779,N_7748);
nand U7865 (N_7865,N_7736,N_7710);
nand U7866 (N_7866,N_7700,N_7711);
nand U7867 (N_7867,N_7684,N_7703);
and U7868 (N_7868,N_7735,N_7714);
and U7869 (N_7869,N_7780,N_7675);
xnor U7870 (N_7870,N_7656,N_7795);
nand U7871 (N_7871,N_7752,N_7708);
xnor U7872 (N_7872,N_7797,N_7663);
nand U7873 (N_7873,N_7767,N_7749);
and U7874 (N_7874,N_7751,N_7659);
or U7875 (N_7875,N_7752,N_7741);
and U7876 (N_7876,N_7772,N_7707);
xnor U7877 (N_7877,N_7752,N_7704);
xnor U7878 (N_7878,N_7745,N_7749);
nand U7879 (N_7879,N_7710,N_7732);
nor U7880 (N_7880,N_7691,N_7751);
nand U7881 (N_7881,N_7657,N_7743);
or U7882 (N_7882,N_7745,N_7797);
xnor U7883 (N_7883,N_7693,N_7752);
or U7884 (N_7884,N_7742,N_7771);
xnor U7885 (N_7885,N_7797,N_7743);
xnor U7886 (N_7886,N_7678,N_7747);
and U7887 (N_7887,N_7782,N_7748);
nand U7888 (N_7888,N_7686,N_7667);
nand U7889 (N_7889,N_7676,N_7780);
nor U7890 (N_7890,N_7767,N_7780);
and U7891 (N_7891,N_7790,N_7724);
nand U7892 (N_7892,N_7761,N_7795);
and U7893 (N_7893,N_7761,N_7703);
nand U7894 (N_7894,N_7699,N_7765);
or U7895 (N_7895,N_7749,N_7776);
xnor U7896 (N_7896,N_7656,N_7704);
nor U7897 (N_7897,N_7725,N_7684);
nor U7898 (N_7898,N_7754,N_7755);
or U7899 (N_7899,N_7796,N_7650);
xnor U7900 (N_7900,N_7670,N_7771);
nand U7901 (N_7901,N_7653,N_7728);
nor U7902 (N_7902,N_7654,N_7713);
nor U7903 (N_7903,N_7797,N_7662);
and U7904 (N_7904,N_7760,N_7697);
nand U7905 (N_7905,N_7670,N_7672);
or U7906 (N_7906,N_7761,N_7756);
nand U7907 (N_7907,N_7673,N_7791);
xnor U7908 (N_7908,N_7732,N_7768);
and U7909 (N_7909,N_7760,N_7732);
nor U7910 (N_7910,N_7781,N_7764);
or U7911 (N_7911,N_7780,N_7666);
xor U7912 (N_7912,N_7725,N_7740);
and U7913 (N_7913,N_7694,N_7774);
and U7914 (N_7914,N_7772,N_7656);
and U7915 (N_7915,N_7668,N_7660);
nand U7916 (N_7916,N_7783,N_7760);
nand U7917 (N_7917,N_7792,N_7794);
nand U7918 (N_7918,N_7782,N_7795);
nand U7919 (N_7919,N_7733,N_7727);
nor U7920 (N_7920,N_7763,N_7762);
nand U7921 (N_7921,N_7668,N_7732);
or U7922 (N_7922,N_7677,N_7714);
xor U7923 (N_7923,N_7737,N_7730);
and U7924 (N_7924,N_7659,N_7722);
nor U7925 (N_7925,N_7709,N_7754);
xnor U7926 (N_7926,N_7653,N_7658);
nand U7927 (N_7927,N_7774,N_7716);
or U7928 (N_7928,N_7771,N_7675);
nor U7929 (N_7929,N_7687,N_7788);
nor U7930 (N_7930,N_7729,N_7721);
or U7931 (N_7931,N_7677,N_7689);
xor U7932 (N_7932,N_7730,N_7679);
xnor U7933 (N_7933,N_7775,N_7733);
nand U7934 (N_7934,N_7664,N_7737);
or U7935 (N_7935,N_7695,N_7714);
and U7936 (N_7936,N_7795,N_7742);
or U7937 (N_7937,N_7711,N_7760);
nand U7938 (N_7938,N_7724,N_7710);
or U7939 (N_7939,N_7736,N_7789);
nor U7940 (N_7940,N_7775,N_7753);
nor U7941 (N_7941,N_7787,N_7700);
and U7942 (N_7942,N_7689,N_7673);
or U7943 (N_7943,N_7727,N_7655);
nand U7944 (N_7944,N_7692,N_7660);
nand U7945 (N_7945,N_7776,N_7762);
nor U7946 (N_7946,N_7720,N_7762);
nor U7947 (N_7947,N_7773,N_7669);
and U7948 (N_7948,N_7665,N_7745);
nand U7949 (N_7949,N_7688,N_7704);
and U7950 (N_7950,N_7864,N_7835);
xnor U7951 (N_7951,N_7851,N_7923);
and U7952 (N_7952,N_7805,N_7813);
and U7953 (N_7953,N_7924,N_7872);
nor U7954 (N_7954,N_7804,N_7831);
or U7955 (N_7955,N_7814,N_7811);
xnor U7956 (N_7956,N_7948,N_7899);
nand U7957 (N_7957,N_7904,N_7861);
nand U7958 (N_7958,N_7856,N_7908);
xor U7959 (N_7959,N_7865,N_7800);
and U7960 (N_7960,N_7870,N_7847);
or U7961 (N_7961,N_7824,N_7852);
nor U7962 (N_7962,N_7817,N_7802);
nand U7963 (N_7963,N_7928,N_7808);
nor U7964 (N_7964,N_7873,N_7897);
or U7965 (N_7965,N_7930,N_7866);
and U7966 (N_7966,N_7819,N_7837);
xnor U7967 (N_7967,N_7853,N_7921);
nor U7968 (N_7968,N_7911,N_7826);
nor U7969 (N_7969,N_7903,N_7929);
and U7970 (N_7970,N_7936,N_7893);
and U7971 (N_7971,N_7886,N_7823);
nor U7972 (N_7972,N_7844,N_7877);
and U7973 (N_7973,N_7935,N_7898);
and U7974 (N_7974,N_7878,N_7910);
xor U7975 (N_7975,N_7916,N_7850);
xor U7976 (N_7976,N_7901,N_7879);
or U7977 (N_7977,N_7927,N_7832);
or U7978 (N_7978,N_7876,N_7891);
or U7979 (N_7979,N_7825,N_7942);
or U7980 (N_7980,N_7863,N_7818);
and U7981 (N_7981,N_7810,N_7933);
nand U7982 (N_7982,N_7827,N_7900);
and U7983 (N_7983,N_7834,N_7809);
or U7984 (N_7984,N_7885,N_7887);
nand U7985 (N_7985,N_7949,N_7862);
and U7986 (N_7986,N_7914,N_7868);
or U7987 (N_7987,N_7833,N_7855);
or U7988 (N_7988,N_7922,N_7880);
and U7989 (N_7989,N_7940,N_7890);
xor U7990 (N_7990,N_7895,N_7892);
nor U7991 (N_7991,N_7943,N_7828);
nor U7992 (N_7992,N_7830,N_7821);
or U7993 (N_7993,N_7857,N_7946);
xnor U7994 (N_7994,N_7913,N_7918);
nor U7995 (N_7995,N_7849,N_7845);
nor U7996 (N_7996,N_7816,N_7836);
and U7997 (N_7997,N_7858,N_7874);
or U7998 (N_7998,N_7812,N_7937);
xor U7999 (N_7999,N_7854,N_7839);
xnor U8000 (N_8000,N_7931,N_7939);
or U8001 (N_8001,N_7884,N_7902);
or U8002 (N_8002,N_7905,N_7894);
nand U8003 (N_8003,N_7925,N_7944);
or U8004 (N_8004,N_7883,N_7871);
or U8005 (N_8005,N_7919,N_7915);
nand U8006 (N_8006,N_7843,N_7842);
nor U8007 (N_8007,N_7841,N_7807);
nand U8008 (N_8008,N_7838,N_7881);
xnor U8009 (N_8009,N_7947,N_7888);
nand U8010 (N_8010,N_7909,N_7906);
and U8011 (N_8011,N_7840,N_7803);
or U8012 (N_8012,N_7907,N_7860);
xnor U8013 (N_8013,N_7859,N_7869);
nor U8014 (N_8014,N_7801,N_7875);
nand U8015 (N_8015,N_7815,N_7882);
nand U8016 (N_8016,N_7829,N_7867);
nand U8017 (N_8017,N_7941,N_7932);
xnor U8018 (N_8018,N_7889,N_7912);
nor U8019 (N_8019,N_7822,N_7934);
and U8020 (N_8020,N_7820,N_7896);
xnor U8021 (N_8021,N_7917,N_7920);
nor U8022 (N_8022,N_7846,N_7938);
and U8023 (N_8023,N_7945,N_7926);
and U8024 (N_8024,N_7848,N_7806);
xnor U8025 (N_8025,N_7909,N_7917);
nor U8026 (N_8026,N_7921,N_7891);
and U8027 (N_8027,N_7907,N_7923);
and U8028 (N_8028,N_7853,N_7920);
nor U8029 (N_8029,N_7823,N_7912);
or U8030 (N_8030,N_7824,N_7853);
or U8031 (N_8031,N_7943,N_7944);
nor U8032 (N_8032,N_7831,N_7898);
and U8033 (N_8033,N_7935,N_7919);
and U8034 (N_8034,N_7932,N_7825);
xor U8035 (N_8035,N_7906,N_7901);
or U8036 (N_8036,N_7809,N_7862);
nor U8037 (N_8037,N_7829,N_7907);
or U8038 (N_8038,N_7873,N_7836);
nor U8039 (N_8039,N_7852,N_7949);
nand U8040 (N_8040,N_7902,N_7812);
nor U8041 (N_8041,N_7805,N_7939);
or U8042 (N_8042,N_7846,N_7931);
and U8043 (N_8043,N_7806,N_7947);
or U8044 (N_8044,N_7921,N_7917);
xnor U8045 (N_8045,N_7802,N_7864);
nor U8046 (N_8046,N_7940,N_7874);
nor U8047 (N_8047,N_7820,N_7889);
and U8048 (N_8048,N_7920,N_7848);
or U8049 (N_8049,N_7904,N_7931);
nor U8050 (N_8050,N_7816,N_7851);
xor U8051 (N_8051,N_7810,N_7909);
nand U8052 (N_8052,N_7830,N_7831);
or U8053 (N_8053,N_7874,N_7942);
xor U8054 (N_8054,N_7860,N_7849);
xor U8055 (N_8055,N_7925,N_7892);
and U8056 (N_8056,N_7849,N_7909);
and U8057 (N_8057,N_7824,N_7820);
and U8058 (N_8058,N_7913,N_7933);
nand U8059 (N_8059,N_7864,N_7838);
nand U8060 (N_8060,N_7921,N_7836);
or U8061 (N_8061,N_7914,N_7876);
or U8062 (N_8062,N_7892,N_7944);
nor U8063 (N_8063,N_7850,N_7917);
xnor U8064 (N_8064,N_7847,N_7851);
xor U8065 (N_8065,N_7946,N_7917);
or U8066 (N_8066,N_7931,N_7858);
and U8067 (N_8067,N_7908,N_7811);
xor U8068 (N_8068,N_7805,N_7860);
nand U8069 (N_8069,N_7884,N_7924);
nand U8070 (N_8070,N_7885,N_7860);
or U8071 (N_8071,N_7876,N_7803);
xor U8072 (N_8072,N_7809,N_7941);
xnor U8073 (N_8073,N_7828,N_7927);
or U8074 (N_8074,N_7873,N_7813);
xor U8075 (N_8075,N_7889,N_7856);
xor U8076 (N_8076,N_7822,N_7871);
nand U8077 (N_8077,N_7901,N_7876);
or U8078 (N_8078,N_7878,N_7935);
nand U8079 (N_8079,N_7808,N_7899);
nand U8080 (N_8080,N_7828,N_7852);
or U8081 (N_8081,N_7839,N_7925);
nor U8082 (N_8082,N_7933,N_7868);
nand U8083 (N_8083,N_7904,N_7927);
xor U8084 (N_8084,N_7945,N_7918);
nor U8085 (N_8085,N_7821,N_7925);
and U8086 (N_8086,N_7929,N_7866);
or U8087 (N_8087,N_7822,N_7878);
nand U8088 (N_8088,N_7875,N_7838);
nor U8089 (N_8089,N_7911,N_7864);
xor U8090 (N_8090,N_7923,N_7919);
nand U8091 (N_8091,N_7846,N_7850);
or U8092 (N_8092,N_7811,N_7858);
nor U8093 (N_8093,N_7850,N_7861);
and U8094 (N_8094,N_7848,N_7802);
nand U8095 (N_8095,N_7844,N_7825);
xnor U8096 (N_8096,N_7932,N_7919);
xor U8097 (N_8097,N_7860,N_7821);
and U8098 (N_8098,N_7846,N_7827);
xnor U8099 (N_8099,N_7848,N_7844);
and U8100 (N_8100,N_7993,N_8032);
xor U8101 (N_8101,N_8018,N_7984);
xnor U8102 (N_8102,N_8041,N_8034);
nand U8103 (N_8103,N_7980,N_7958);
nand U8104 (N_8104,N_8043,N_8022);
nor U8105 (N_8105,N_8038,N_8097);
and U8106 (N_8106,N_7982,N_7994);
nand U8107 (N_8107,N_7974,N_8062);
xor U8108 (N_8108,N_8016,N_8010);
xor U8109 (N_8109,N_7951,N_7996);
and U8110 (N_8110,N_7975,N_8075);
nor U8111 (N_8111,N_8071,N_8098);
and U8112 (N_8112,N_7972,N_8030);
nand U8113 (N_8113,N_8024,N_8007);
and U8114 (N_8114,N_8060,N_7997);
nand U8115 (N_8115,N_8039,N_8077);
or U8116 (N_8116,N_8087,N_8074);
nor U8117 (N_8117,N_7961,N_8037);
xor U8118 (N_8118,N_7978,N_7977);
or U8119 (N_8119,N_7965,N_7963);
and U8120 (N_8120,N_8061,N_8057);
or U8121 (N_8121,N_8080,N_8036);
and U8122 (N_8122,N_7950,N_8025);
xor U8123 (N_8123,N_8083,N_7987);
or U8124 (N_8124,N_8005,N_7986);
or U8125 (N_8125,N_8052,N_7955);
xnor U8126 (N_8126,N_8058,N_8063);
nor U8127 (N_8127,N_8019,N_8065);
or U8128 (N_8128,N_7998,N_7989);
xor U8129 (N_8129,N_8045,N_8092);
xnor U8130 (N_8130,N_8090,N_8093);
and U8131 (N_8131,N_8050,N_8042);
nand U8132 (N_8132,N_8064,N_8070);
nand U8133 (N_8133,N_8051,N_7954);
nor U8134 (N_8134,N_7964,N_8084);
or U8135 (N_8135,N_8066,N_8095);
nand U8136 (N_8136,N_8078,N_7956);
nand U8137 (N_8137,N_8068,N_7973);
or U8138 (N_8138,N_7985,N_8086);
nor U8139 (N_8139,N_8040,N_8029);
nand U8140 (N_8140,N_8072,N_7976);
xnor U8141 (N_8141,N_8012,N_8082);
nand U8142 (N_8142,N_8085,N_7995);
or U8143 (N_8143,N_8028,N_8009);
xnor U8144 (N_8144,N_7979,N_8044);
and U8145 (N_8145,N_8079,N_7990);
nand U8146 (N_8146,N_7960,N_8023);
nand U8147 (N_8147,N_8031,N_8003);
nor U8148 (N_8148,N_8026,N_7999);
and U8149 (N_8149,N_7967,N_8091);
or U8150 (N_8150,N_7969,N_7971);
nand U8151 (N_8151,N_7981,N_7962);
xor U8152 (N_8152,N_8056,N_8033);
or U8153 (N_8153,N_8055,N_7991);
nor U8154 (N_8154,N_8013,N_8000);
xnor U8155 (N_8155,N_7988,N_8094);
or U8156 (N_8156,N_8006,N_7957);
nor U8157 (N_8157,N_8027,N_7968);
and U8158 (N_8158,N_8073,N_8067);
nand U8159 (N_8159,N_8008,N_8054);
or U8160 (N_8160,N_8047,N_8004);
and U8161 (N_8161,N_8001,N_7953);
xnor U8162 (N_8162,N_8099,N_8014);
or U8163 (N_8163,N_8053,N_8096);
or U8164 (N_8164,N_8017,N_8021);
and U8165 (N_8165,N_7992,N_8059);
nand U8166 (N_8166,N_8046,N_8020);
or U8167 (N_8167,N_7966,N_8011);
nand U8168 (N_8168,N_8069,N_8049);
or U8169 (N_8169,N_8089,N_7970);
nand U8170 (N_8170,N_8076,N_8081);
nor U8171 (N_8171,N_8002,N_8015);
or U8172 (N_8172,N_7959,N_7952);
nand U8173 (N_8173,N_8035,N_7983);
xnor U8174 (N_8174,N_8088,N_8048);
xnor U8175 (N_8175,N_8009,N_7979);
or U8176 (N_8176,N_8006,N_8008);
nand U8177 (N_8177,N_7973,N_7991);
and U8178 (N_8178,N_8066,N_8087);
and U8179 (N_8179,N_8043,N_8048);
nor U8180 (N_8180,N_8048,N_8003);
xnor U8181 (N_8181,N_8000,N_8094);
nand U8182 (N_8182,N_8076,N_7977);
nor U8183 (N_8183,N_8075,N_8044);
and U8184 (N_8184,N_8017,N_8038);
nor U8185 (N_8185,N_7979,N_8013);
nand U8186 (N_8186,N_8032,N_8043);
xor U8187 (N_8187,N_8073,N_8044);
xor U8188 (N_8188,N_7978,N_8061);
xor U8189 (N_8189,N_8017,N_8016);
and U8190 (N_8190,N_7956,N_8085);
or U8191 (N_8191,N_8024,N_8081);
xnor U8192 (N_8192,N_7990,N_8050);
xor U8193 (N_8193,N_7979,N_7953);
xor U8194 (N_8194,N_7952,N_8068);
and U8195 (N_8195,N_7967,N_8047);
or U8196 (N_8196,N_7990,N_8053);
and U8197 (N_8197,N_8072,N_8004);
and U8198 (N_8198,N_8039,N_8031);
and U8199 (N_8199,N_7969,N_8064);
xnor U8200 (N_8200,N_7989,N_8051);
and U8201 (N_8201,N_8089,N_7968);
or U8202 (N_8202,N_7956,N_8028);
and U8203 (N_8203,N_8067,N_7992);
xnor U8204 (N_8204,N_8081,N_8036);
xor U8205 (N_8205,N_8052,N_7984);
and U8206 (N_8206,N_8076,N_7952);
nor U8207 (N_8207,N_8011,N_8020);
nor U8208 (N_8208,N_8029,N_7970);
nor U8209 (N_8209,N_7984,N_8023);
xor U8210 (N_8210,N_7950,N_8003);
nor U8211 (N_8211,N_7961,N_8094);
and U8212 (N_8212,N_8048,N_8000);
nand U8213 (N_8213,N_7971,N_8057);
or U8214 (N_8214,N_7968,N_7957);
nor U8215 (N_8215,N_8020,N_7990);
nor U8216 (N_8216,N_7989,N_7952);
and U8217 (N_8217,N_7990,N_7972);
nand U8218 (N_8218,N_7998,N_8084);
nor U8219 (N_8219,N_8065,N_8058);
nand U8220 (N_8220,N_8006,N_8042);
and U8221 (N_8221,N_8015,N_8077);
nand U8222 (N_8222,N_7968,N_8086);
and U8223 (N_8223,N_8081,N_7973);
and U8224 (N_8224,N_8018,N_8020);
and U8225 (N_8225,N_8006,N_7987);
and U8226 (N_8226,N_8049,N_8009);
xnor U8227 (N_8227,N_8045,N_8006);
and U8228 (N_8228,N_8001,N_8083);
and U8229 (N_8229,N_7961,N_8089);
and U8230 (N_8230,N_8047,N_8040);
nor U8231 (N_8231,N_8066,N_8049);
nor U8232 (N_8232,N_7963,N_8031);
xnor U8233 (N_8233,N_8026,N_8071);
and U8234 (N_8234,N_8096,N_8001);
and U8235 (N_8235,N_7976,N_7973);
and U8236 (N_8236,N_7988,N_7971);
and U8237 (N_8237,N_8072,N_8060);
nor U8238 (N_8238,N_8071,N_7989);
and U8239 (N_8239,N_8011,N_8027);
and U8240 (N_8240,N_7968,N_8009);
or U8241 (N_8241,N_7983,N_8013);
nand U8242 (N_8242,N_8037,N_7977);
nor U8243 (N_8243,N_8081,N_8042);
nand U8244 (N_8244,N_7987,N_8001);
nor U8245 (N_8245,N_8092,N_8034);
nand U8246 (N_8246,N_7983,N_8093);
or U8247 (N_8247,N_8095,N_8079);
nand U8248 (N_8248,N_8059,N_8010);
and U8249 (N_8249,N_8024,N_8095);
nor U8250 (N_8250,N_8177,N_8165);
nor U8251 (N_8251,N_8154,N_8157);
xnor U8252 (N_8252,N_8144,N_8147);
nor U8253 (N_8253,N_8232,N_8136);
nor U8254 (N_8254,N_8238,N_8166);
nor U8255 (N_8255,N_8218,N_8241);
xor U8256 (N_8256,N_8248,N_8172);
nor U8257 (N_8257,N_8102,N_8100);
and U8258 (N_8258,N_8203,N_8223);
or U8259 (N_8259,N_8162,N_8148);
and U8260 (N_8260,N_8143,N_8122);
or U8261 (N_8261,N_8108,N_8197);
nand U8262 (N_8262,N_8133,N_8187);
or U8263 (N_8263,N_8135,N_8155);
and U8264 (N_8264,N_8201,N_8196);
xnor U8265 (N_8265,N_8236,N_8225);
and U8266 (N_8266,N_8184,N_8234);
nand U8267 (N_8267,N_8119,N_8137);
or U8268 (N_8268,N_8182,N_8204);
nor U8269 (N_8269,N_8142,N_8240);
nand U8270 (N_8270,N_8169,N_8126);
nand U8271 (N_8271,N_8115,N_8207);
and U8272 (N_8272,N_8216,N_8185);
or U8273 (N_8273,N_8239,N_8183);
nand U8274 (N_8274,N_8180,N_8167);
nand U8275 (N_8275,N_8249,N_8128);
nand U8276 (N_8276,N_8212,N_8176);
or U8277 (N_8277,N_8174,N_8200);
and U8278 (N_8278,N_8246,N_8149);
xnor U8279 (N_8279,N_8211,N_8171);
or U8280 (N_8280,N_8129,N_8151);
nand U8281 (N_8281,N_8202,N_8130);
nand U8282 (N_8282,N_8138,N_8146);
nand U8283 (N_8283,N_8134,N_8243);
nor U8284 (N_8284,N_8199,N_8164);
or U8285 (N_8285,N_8161,N_8231);
or U8286 (N_8286,N_8219,N_8117);
and U8287 (N_8287,N_8118,N_8139);
or U8288 (N_8288,N_8103,N_8215);
nand U8289 (N_8289,N_8229,N_8141);
xor U8290 (N_8290,N_8210,N_8107);
xnor U8291 (N_8291,N_8173,N_8163);
nand U8292 (N_8292,N_8230,N_8221);
and U8293 (N_8293,N_8244,N_8153);
or U8294 (N_8294,N_8245,N_8110);
nand U8295 (N_8295,N_8193,N_8208);
nand U8296 (N_8296,N_8140,N_8111);
and U8297 (N_8297,N_8220,N_8179);
nand U8298 (N_8298,N_8213,N_8168);
nor U8299 (N_8299,N_8237,N_8222);
nor U8300 (N_8300,N_8131,N_8233);
or U8301 (N_8301,N_8227,N_8132);
nor U8302 (N_8302,N_8109,N_8247);
xnor U8303 (N_8303,N_8116,N_8175);
nand U8304 (N_8304,N_8217,N_8181);
nor U8305 (N_8305,N_8206,N_8191);
or U8306 (N_8306,N_8159,N_8198);
xor U8307 (N_8307,N_8205,N_8226);
or U8308 (N_8308,N_8105,N_8152);
nand U8309 (N_8309,N_8209,N_8113);
or U8310 (N_8310,N_8195,N_8192);
xnor U8311 (N_8311,N_8178,N_8124);
nand U8312 (N_8312,N_8101,N_8214);
nand U8313 (N_8313,N_8106,N_8158);
nand U8314 (N_8314,N_8125,N_8114);
xor U8315 (N_8315,N_8190,N_8224);
and U8316 (N_8316,N_8228,N_8160);
and U8317 (N_8317,N_8112,N_8120);
or U8318 (N_8318,N_8235,N_8121);
or U8319 (N_8319,N_8189,N_8145);
and U8320 (N_8320,N_8170,N_8194);
nand U8321 (N_8321,N_8242,N_8127);
xor U8322 (N_8322,N_8156,N_8104);
nor U8323 (N_8323,N_8150,N_8186);
xor U8324 (N_8324,N_8123,N_8188);
or U8325 (N_8325,N_8129,N_8216);
nand U8326 (N_8326,N_8150,N_8112);
or U8327 (N_8327,N_8221,N_8134);
nand U8328 (N_8328,N_8145,N_8123);
and U8329 (N_8329,N_8204,N_8145);
nor U8330 (N_8330,N_8151,N_8137);
or U8331 (N_8331,N_8209,N_8157);
or U8332 (N_8332,N_8146,N_8240);
nor U8333 (N_8333,N_8163,N_8241);
xnor U8334 (N_8334,N_8218,N_8150);
or U8335 (N_8335,N_8102,N_8132);
nand U8336 (N_8336,N_8162,N_8131);
and U8337 (N_8337,N_8228,N_8227);
xor U8338 (N_8338,N_8144,N_8227);
xnor U8339 (N_8339,N_8167,N_8208);
and U8340 (N_8340,N_8138,N_8175);
or U8341 (N_8341,N_8209,N_8129);
or U8342 (N_8342,N_8245,N_8209);
and U8343 (N_8343,N_8239,N_8131);
nand U8344 (N_8344,N_8232,N_8157);
nor U8345 (N_8345,N_8232,N_8100);
nor U8346 (N_8346,N_8111,N_8150);
xor U8347 (N_8347,N_8179,N_8176);
xnor U8348 (N_8348,N_8185,N_8157);
or U8349 (N_8349,N_8129,N_8145);
nand U8350 (N_8350,N_8206,N_8221);
or U8351 (N_8351,N_8137,N_8162);
xnor U8352 (N_8352,N_8188,N_8162);
xor U8353 (N_8353,N_8124,N_8136);
nand U8354 (N_8354,N_8152,N_8205);
or U8355 (N_8355,N_8232,N_8187);
nor U8356 (N_8356,N_8177,N_8230);
nor U8357 (N_8357,N_8244,N_8102);
or U8358 (N_8358,N_8234,N_8249);
nand U8359 (N_8359,N_8117,N_8171);
nand U8360 (N_8360,N_8163,N_8142);
nand U8361 (N_8361,N_8107,N_8189);
nand U8362 (N_8362,N_8230,N_8211);
or U8363 (N_8363,N_8218,N_8120);
nand U8364 (N_8364,N_8191,N_8233);
or U8365 (N_8365,N_8121,N_8172);
nand U8366 (N_8366,N_8115,N_8222);
xor U8367 (N_8367,N_8178,N_8246);
xor U8368 (N_8368,N_8156,N_8112);
xnor U8369 (N_8369,N_8199,N_8136);
nand U8370 (N_8370,N_8175,N_8180);
nand U8371 (N_8371,N_8226,N_8212);
nand U8372 (N_8372,N_8119,N_8146);
xor U8373 (N_8373,N_8170,N_8184);
and U8374 (N_8374,N_8152,N_8177);
xnor U8375 (N_8375,N_8211,N_8204);
nor U8376 (N_8376,N_8143,N_8210);
or U8377 (N_8377,N_8179,N_8180);
nor U8378 (N_8378,N_8175,N_8117);
and U8379 (N_8379,N_8177,N_8166);
or U8380 (N_8380,N_8217,N_8188);
xnor U8381 (N_8381,N_8247,N_8102);
nor U8382 (N_8382,N_8130,N_8207);
xor U8383 (N_8383,N_8119,N_8112);
and U8384 (N_8384,N_8177,N_8187);
nor U8385 (N_8385,N_8204,N_8189);
nor U8386 (N_8386,N_8125,N_8127);
nand U8387 (N_8387,N_8235,N_8168);
or U8388 (N_8388,N_8202,N_8200);
xnor U8389 (N_8389,N_8163,N_8170);
or U8390 (N_8390,N_8169,N_8242);
and U8391 (N_8391,N_8110,N_8120);
nor U8392 (N_8392,N_8236,N_8230);
nand U8393 (N_8393,N_8244,N_8107);
nand U8394 (N_8394,N_8135,N_8217);
nand U8395 (N_8395,N_8104,N_8138);
xnor U8396 (N_8396,N_8151,N_8236);
xnor U8397 (N_8397,N_8191,N_8176);
nand U8398 (N_8398,N_8219,N_8132);
and U8399 (N_8399,N_8154,N_8106);
and U8400 (N_8400,N_8390,N_8285);
xor U8401 (N_8401,N_8326,N_8258);
nor U8402 (N_8402,N_8317,N_8274);
or U8403 (N_8403,N_8280,N_8360);
nand U8404 (N_8404,N_8295,N_8385);
or U8405 (N_8405,N_8270,N_8395);
or U8406 (N_8406,N_8296,N_8349);
nor U8407 (N_8407,N_8352,N_8333);
nand U8408 (N_8408,N_8346,N_8377);
nand U8409 (N_8409,N_8345,N_8311);
xor U8410 (N_8410,N_8332,N_8253);
or U8411 (N_8411,N_8392,N_8373);
and U8412 (N_8412,N_8279,N_8272);
xnor U8413 (N_8413,N_8366,N_8355);
xnor U8414 (N_8414,N_8267,N_8251);
and U8415 (N_8415,N_8320,N_8268);
or U8416 (N_8416,N_8287,N_8310);
xor U8417 (N_8417,N_8353,N_8271);
nor U8418 (N_8418,N_8291,N_8262);
and U8419 (N_8419,N_8259,N_8257);
or U8420 (N_8420,N_8380,N_8281);
nand U8421 (N_8421,N_8396,N_8264);
nor U8422 (N_8422,N_8312,N_8398);
or U8423 (N_8423,N_8273,N_8315);
or U8424 (N_8424,N_8293,N_8382);
and U8425 (N_8425,N_8278,N_8364);
nand U8426 (N_8426,N_8391,N_8260);
or U8427 (N_8427,N_8277,N_8358);
nor U8428 (N_8428,N_8322,N_8276);
nand U8429 (N_8429,N_8284,N_8359);
or U8430 (N_8430,N_8265,N_8368);
or U8431 (N_8431,N_8339,N_8314);
nand U8432 (N_8432,N_8361,N_8250);
or U8433 (N_8433,N_8350,N_8301);
nor U8434 (N_8434,N_8338,N_8288);
or U8435 (N_8435,N_8351,N_8397);
or U8436 (N_8436,N_8297,N_8254);
xor U8437 (N_8437,N_8393,N_8354);
nand U8438 (N_8438,N_8399,N_8263);
or U8439 (N_8439,N_8266,N_8302);
xor U8440 (N_8440,N_8356,N_8367);
xor U8441 (N_8441,N_8292,N_8341);
or U8442 (N_8442,N_8289,N_8389);
and U8443 (N_8443,N_8337,N_8376);
nor U8444 (N_8444,N_8298,N_8307);
and U8445 (N_8445,N_8379,N_8316);
xor U8446 (N_8446,N_8256,N_8275);
and U8447 (N_8447,N_8381,N_8363);
xnor U8448 (N_8448,N_8304,N_8255);
xor U8449 (N_8449,N_8303,N_8374);
nor U8450 (N_8450,N_8283,N_8369);
nand U8451 (N_8451,N_8387,N_8261);
nand U8452 (N_8452,N_8318,N_8313);
or U8453 (N_8453,N_8334,N_8331);
nand U8454 (N_8454,N_8372,N_8323);
nor U8455 (N_8455,N_8347,N_8299);
nand U8456 (N_8456,N_8342,N_8357);
and U8457 (N_8457,N_8335,N_8394);
xor U8458 (N_8458,N_8383,N_8252);
and U8459 (N_8459,N_8321,N_8329);
xnor U8460 (N_8460,N_8336,N_8378);
nand U8461 (N_8461,N_8371,N_8282);
or U8462 (N_8462,N_8343,N_8344);
xor U8463 (N_8463,N_8388,N_8340);
xnor U8464 (N_8464,N_8300,N_8384);
nand U8465 (N_8465,N_8290,N_8362);
or U8466 (N_8466,N_8286,N_8375);
xnor U8467 (N_8467,N_8309,N_8328);
nor U8468 (N_8468,N_8294,N_8269);
nand U8469 (N_8469,N_8324,N_8305);
nor U8470 (N_8470,N_8330,N_8306);
or U8471 (N_8471,N_8319,N_8370);
xnor U8472 (N_8472,N_8386,N_8348);
and U8473 (N_8473,N_8325,N_8308);
or U8474 (N_8474,N_8365,N_8327);
and U8475 (N_8475,N_8366,N_8356);
or U8476 (N_8476,N_8388,N_8390);
nor U8477 (N_8477,N_8288,N_8284);
and U8478 (N_8478,N_8251,N_8341);
or U8479 (N_8479,N_8332,N_8340);
nor U8480 (N_8480,N_8304,N_8326);
or U8481 (N_8481,N_8379,N_8293);
and U8482 (N_8482,N_8340,N_8348);
and U8483 (N_8483,N_8324,N_8330);
nand U8484 (N_8484,N_8319,N_8312);
nor U8485 (N_8485,N_8289,N_8287);
xor U8486 (N_8486,N_8281,N_8280);
and U8487 (N_8487,N_8336,N_8304);
nand U8488 (N_8488,N_8367,N_8297);
and U8489 (N_8489,N_8327,N_8263);
nor U8490 (N_8490,N_8383,N_8366);
or U8491 (N_8491,N_8371,N_8314);
xor U8492 (N_8492,N_8300,N_8263);
nand U8493 (N_8493,N_8399,N_8306);
xnor U8494 (N_8494,N_8278,N_8288);
nand U8495 (N_8495,N_8253,N_8381);
nor U8496 (N_8496,N_8382,N_8326);
xnor U8497 (N_8497,N_8376,N_8275);
and U8498 (N_8498,N_8333,N_8255);
and U8499 (N_8499,N_8287,N_8321);
xnor U8500 (N_8500,N_8338,N_8293);
and U8501 (N_8501,N_8398,N_8346);
xnor U8502 (N_8502,N_8379,N_8342);
or U8503 (N_8503,N_8385,N_8307);
xor U8504 (N_8504,N_8283,N_8270);
and U8505 (N_8505,N_8346,N_8372);
or U8506 (N_8506,N_8349,N_8320);
and U8507 (N_8507,N_8361,N_8350);
and U8508 (N_8508,N_8287,N_8260);
or U8509 (N_8509,N_8272,N_8293);
xnor U8510 (N_8510,N_8355,N_8299);
and U8511 (N_8511,N_8396,N_8363);
xor U8512 (N_8512,N_8374,N_8265);
or U8513 (N_8513,N_8291,N_8362);
nand U8514 (N_8514,N_8352,N_8390);
and U8515 (N_8515,N_8292,N_8294);
nor U8516 (N_8516,N_8316,N_8305);
or U8517 (N_8517,N_8377,N_8276);
nand U8518 (N_8518,N_8355,N_8277);
or U8519 (N_8519,N_8352,N_8256);
nor U8520 (N_8520,N_8280,N_8304);
and U8521 (N_8521,N_8261,N_8388);
or U8522 (N_8522,N_8311,N_8266);
xnor U8523 (N_8523,N_8292,N_8310);
xnor U8524 (N_8524,N_8279,N_8384);
or U8525 (N_8525,N_8265,N_8341);
or U8526 (N_8526,N_8345,N_8267);
or U8527 (N_8527,N_8373,N_8352);
xnor U8528 (N_8528,N_8263,N_8344);
nand U8529 (N_8529,N_8370,N_8373);
nand U8530 (N_8530,N_8357,N_8360);
xor U8531 (N_8531,N_8268,N_8289);
and U8532 (N_8532,N_8322,N_8304);
or U8533 (N_8533,N_8292,N_8385);
nand U8534 (N_8534,N_8379,N_8363);
nand U8535 (N_8535,N_8266,N_8340);
or U8536 (N_8536,N_8330,N_8368);
and U8537 (N_8537,N_8377,N_8399);
or U8538 (N_8538,N_8273,N_8338);
and U8539 (N_8539,N_8380,N_8294);
or U8540 (N_8540,N_8324,N_8346);
nor U8541 (N_8541,N_8286,N_8264);
nand U8542 (N_8542,N_8265,N_8337);
nor U8543 (N_8543,N_8381,N_8390);
nand U8544 (N_8544,N_8387,N_8301);
and U8545 (N_8545,N_8383,N_8254);
nand U8546 (N_8546,N_8272,N_8253);
or U8547 (N_8547,N_8385,N_8254);
or U8548 (N_8548,N_8341,N_8373);
nand U8549 (N_8549,N_8392,N_8308);
or U8550 (N_8550,N_8414,N_8462);
nor U8551 (N_8551,N_8536,N_8465);
and U8552 (N_8552,N_8458,N_8519);
nand U8553 (N_8553,N_8432,N_8491);
xor U8554 (N_8554,N_8540,N_8548);
and U8555 (N_8555,N_8404,N_8401);
and U8556 (N_8556,N_8406,N_8507);
xor U8557 (N_8557,N_8433,N_8533);
nand U8558 (N_8558,N_8488,N_8480);
or U8559 (N_8559,N_8419,N_8439);
or U8560 (N_8560,N_8485,N_8466);
and U8561 (N_8561,N_8441,N_8454);
and U8562 (N_8562,N_8509,N_8434);
xnor U8563 (N_8563,N_8522,N_8421);
nand U8564 (N_8564,N_8436,N_8407);
xnor U8565 (N_8565,N_8526,N_8424);
xnor U8566 (N_8566,N_8475,N_8410);
nand U8567 (N_8567,N_8409,N_8531);
xnor U8568 (N_8568,N_8517,N_8473);
xor U8569 (N_8569,N_8506,N_8513);
xor U8570 (N_8570,N_8493,N_8455);
or U8571 (N_8571,N_8515,N_8511);
and U8572 (N_8572,N_8464,N_8476);
nor U8573 (N_8573,N_8463,N_8541);
or U8574 (N_8574,N_8435,N_8415);
nor U8575 (N_8575,N_8474,N_8411);
xor U8576 (N_8576,N_8484,N_8448);
nand U8577 (N_8577,N_8451,N_8481);
nor U8578 (N_8578,N_8518,N_8446);
and U8579 (N_8579,N_8537,N_8489);
or U8580 (N_8580,N_8437,N_8461);
xor U8581 (N_8581,N_8445,N_8505);
xnor U8582 (N_8582,N_8490,N_8542);
or U8583 (N_8583,N_8494,N_8539);
nor U8584 (N_8584,N_8479,N_8472);
xor U8585 (N_8585,N_8524,N_8449);
or U8586 (N_8586,N_8525,N_8413);
or U8587 (N_8587,N_8516,N_8402);
nor U8588 (N_8588,N_8440,N_8460);
or U8589 (N_8589,N_8504,N_8529);
or U8590 (N_8590,N_8423,N_8544);
xnor U8591 (N_8591,N_8412,N_8532);
or U8592 (N_8592,N_8501,N_8444);
nand U8593 (N_8593,N_8500,N_8503);
and U8594 (N_8594,N_8416,N_8502);
nor U8595 (N_8595,N_8523,N_8450);
nor U8596 (N_8596,N_8534,N_8510);
xor U8597 (N_8597,N_8405,N_8477);
and U8598 (N_8598,N_8438,N_8549);
and U8599 (N_8599,N_8520,N_8425);
nor U8600 (N_8600,N_8420,N_8497);
nor U8601 (N_8601,N_8547,N_8478);
or U8602 (N_8602,N_8470,N_8442);
and U8603 (N_8603,N_8512,N_8443);
and U8604 (N_8604,N_8498,N_8456);
and U8605 (N_8605,N_8459,N_8508);
nand U8606 (N_8606,N_8543,N_8528);
nand U8607 (N_8607,N_8545,N_8417);
nor U8608 (N_8608,N_8452,N_8487);
or U8609 (N_8609,N_8431,N_8527);
nand U8610 (N_8610,N_8403,N_8483);
nor U8611 (N_8611,N_8486,N_8427);
nand U8612 (N_8612,N_8535,N_8499);
nand U8613 (N_8613,N_8495,N_8453);
nand U8614 (N_8614,N_8492,N_8418);
nand U8615 (N_8615,N_8400,N_8430);
nand U8616 (N_8616,N_8538,N_8521);
and U8617 (N_8617,N_8426,N_8429);
and U8618 (N_8618,N_8496,N_8530);
xor U8619 (N_8619,N_8546,N_8469);
nand U8620 (N_8620,N_8471,N_8428);
or U8621 (N_8621,N_8447,N_8408);
xor U8622 (N_8622,N_8514,N_8468);
and U8623 (N_8623,N_8457,N_8422);
xnor U8624 (N_8624,N_8482,N_8467);
and U8625 (N_8625,N_8548,N_8533);
nor U8626 (N_8626,N_8415,N_8487);
xor U8627 (N_8627,N_8443,N_8403);
or U8628 (N_8628,N_8462,N_8540);
nand U8629 (N_8629,N_8507,N_8414);
nor U8630 (N_8630,N_8481,N_8400);
nor U8631 (N_8631,N_8469,N_8501);
nand U8632 (N_8632,N_8512,N_8439);
nand U8633 (N_8633,N_8431,N_8484);
nand U8634 (N_8634,N_8510,N_8506);
xnor U8635 (N_8635,N_8524,N_8438);
xnor U8636 (N_8636,N_8519,N_8422);
or U8637 (N_8637,N_8430,N_8442);
nand U8638 (N_8638,N_8471,N_8506);
xor U8639 (N_8639,N_8409,N_8427);
or U8640 (N_8640,N_8421,N_8455);
nand U8641 (N_8641,N_8401,N_8549);
xor U8642 (N_8642,N_8480,N_8512);
nand U8643 (N_8643,N_8444,N_8502);
or U8644 (N_8644,N_8440,N_8523);
nand U8645 (N_8645,N_8435,N_8533);
nand U8646 (N_8646,N_8407,N_8405);
or U8647 (N_8647,N_8462,N_8468);
nor U8648 (N_8648,N_8419,N_8479);
xor U8649 (N_8649,N_8402,N_8425);
nor U8650 (N_8650,N_8547,N_8454);
nand U8651 (N_8651,N_8458,N_8434);
nor U8652 (N_8652,N_8510,N_8443);
and U8653 (N_8653,N_8410,N_8428);
and U8654 (N_8654,N_8528,N_8409);
and U8655 (N_8655,N_8443,N_8549);
or U8656 (N_8656,N_8440,N_8448);
xor U8657 (N_8657,N_8515,N_8545);
nor U8658 (N_8658,N_8458,N_8401);
nand U8659 (N_8659,N_8401,N_8423);
or U8660 (N_8660,N_8465,N_8493);
or U8661 (N_8661,N_8430,N_8493);
nand U8662 (N_8662,N_8524,N_8526);
or U8663 (N_8663,N_8533,N_8515);
nor U8664 (N_8664,N_8454,N_8467);
and U8665 (N_8665,N_8483,N_8525);
or U8666 (N_8666,N_8433,N_8445);
nand U8667 (N_8667,N_8458,N_8491);
or U8668 (N_8668,N_8410,N_8510);
nand U8669 (N_8669,N_8463,N_8515);
xnor U8670 (N_8670,N_8493,N_8511);
nor U8671 (N_8671,N_8494,N_8530);
or U8672 (N_8672,N_8474,N_8402);
and U8673 (N_8673,N_8414,N_8486);
xor U8674 (N_8674,N_8514,N_8459);
or U8675 (N_8675,N_8536,N_8467);
or U8676 (N_8676,N_8430,N_8525);
nor U8677 (N_8677,N_8513,N_8452);
nand U8678 (N_8678,N_8483,N_8401);
or U8679 (N_8679,N_8491,N_8533);
nor U8680 (N_8680,N_8479,N_8436);
nand U8681 (N_8681,N_8417,N_8443);
or U8682 (N_8682,N_8480,N_8427);
and U8683 (N_8683,N_8506,N_8507);
nand U8684 (N_8684,N_8402,N_8489);
nand U8685 (N_8685,N_8509,N_8520);
and U8686 (N_8686,N_8436,N_8432);
nor U8687 (N_8687,N_8529,N_8427);
xor U8688 (N_8688,N_8514,N_8519);
nand U8689 (N_8689,N_8510,N_8430);
xnor U8690 (N_8690,N_8493,N_8494);
and U8691 (N_8691,N_8547,N_8465);
xnor U8692 (N_8692,N_8534,N_8463);
and U8693 (N_8693,N_8518,N_8491);
and U8694 (N_8694,N_8462,N_8506);
or U8695 (N_8695,N_8471,N_8472);
nand U8696 (N_8696,N_8470,N_8404);
or U8697 (N_8697,N_8545,N_8465);
nor U8698 (N_8698,N_8502,N_8420);
nor U8699 (N_8699,N_8496,N_8510);
or U8700 (N_8700,N_8645,N_8661);
or U8701 (N_8701,N_8616,N_8672);
or U8702 (N_8702,N_8583,N_8551);
xor U8703 (N_8703,N_8642,N_8613);
xnor U8704 (N_8704,N_8691,N_8608);
or U8705 (N_8705,N_8654,N_8678);
and U8706 (N_8706,N_8669,N_8657);
xor U8707 (N_8707,N_8597,N_8658);
and U8708 (N_8708,N_8580,N_8681);
and U8709 (N_8709,N_8664,N_8600);
xnor U8710 (N_8710,N_8632,N_8559);
nand U8711 (N_8711,N_8556,N_8698);
or U8712 (N_8712,N_8574,N_8618);
xor U8713 (N_8713,N_8635,N_8594);
nand U8714 (N_8714,N_8550,N_8655);
or U8715 (N_8715,N_8629,N_8590);
nand U8716 (N_8716,N_8586,N_8566);
xnor U8717 (N_8717,N_8578,N_8606);
nand U8718 (N_8718,N_8628,N_8640);
or U8719 (N_8719,N_8568,N_8679);
xor U8720 (N_8720,N_8572,N_8588);
nor U8721 (N_8721,N_8693,N_8584);
nand U8722 (N_8722,N_8697,N_8569);
or U8723 (N_8723,N_8633,N_8620);
xor U8724 (N_8724,N_8627,N_8682);
or U8725 (N_8725,N_8675,N_8601);
xor U8726 (N_8726,N_8611,N_8663);
nor U8727 (N_8727,N_8687,N_8621);
or U8728 (N_8728,N_8587,N_8619);
nand U8729 (N_8729,N_8579,N_8636);
nor U8730 (N_8730,N_8596,N_8667);
nor U8731 (N_8731,N_8685,N_8607);
or U8732 (N_8732,N_8638,N_8650);
and U8733 (N_8733,N_8576,N_8646);
nor U8734 (N_8734,N_8552,N_8603);
xor U8735 (N_8735,N_8564,N_8592);
and U8736 (N_8736,N_8557,N_8692);
xor U8737 (N_8737,N_8575,N_8615);
xor U8738 (N_8738,N_8688,N_8625);
nand U8739 (N_8739,N_8585,N_8674);
nand U8740 (N_8740,N_8609,N_8602);
nor U8741 (N_8741,N_8589,N_8660);
and U8742 (N_8742,N_8604,N_8652);
and U8743 (N_8743,N_8623,N_8555);
nand U8744 (N_8744,N_8651,N_8573);
or U8745 (N_8745,N_8659,N_8570);
nand U8746 (N_8746,N_8553,N_8641);
nor U8747 (N_8747,N_8591,N_8631);
nand U8748 (N_8748,N_8662,N_8673);
or U8749 (N_8749,N_8690,N_8665);
xor U8750 (N_8750,N_8643,N_8581);
nand U8751 (N_8751,N_8622,N_8595);
and U8752 (N_8752,N_8626,N_8637);
nor U8753 (N_8753,N_8605,N_8617);
xnor U8754 (N_8754,N_8695,N_8577);
nand U8755 (N_8755,N_8639,N_8554);
and U8756 (N_8756,N_8582,N_8567);
nor U8757 (N_8757,N_8647,N_8653);
and U8758 (N_8758,N_8684,N_8699);
xnor U8759 (N_8759,N_8677,N_8696);
and U8760 (N_8760,N_8649,N_8610);
and U8761 (N_8761,N_8683,N_8560);
nand U8762 (N_8762,N_8561,N_8656);
nor U8763 (N_8763,N_8644,N_8671);
and U8764 (N_8764,N_8612,N_8571);
xnor U8765 (N_8765,N_8676,N_8562);
and U8766 (N_8766,N_8666,N_8686);
xnor U8767 (N_8767,N_8563,N_8565);
xnor U8768 (N_8768,N_8593,N_8648);
xnor U8769 (N_8769,N_8599,N_8634);
nand U8770 (N_8770,N_8694,N_8630);
nor U8771 (N_8771,N_8670,N_8689);
nand U8772 (N_8772,N_8598,N_8668);
nor U8773 (N_8773,N_8558,N_8680);
nand U8774 (N_8774,N_8624,N_8614);
nand U8775 (N_8775,N_8673,N_8615);
and U8776 (N_8776,N_8641,N_8688);
xor U8777 (N_8777,N_8558,N_8646);
xor U8778 (N_8778,N_8613,N_8639);
nor U8779 (N_8779,N_8663,N_8652);
and U8780 (N_8780,N_8589,N_8614);
and U8781 (N_8781,N_8566,N_8579);
xnor U8782 (N_8782,N_8613,N_8634);
nor U8783 (N_8783,N_8551,N_8696);
nand U8784 (N_8784,N_8569,N_8554);
or U8785 (N_8785,N_8555,N_8696);
nor U8786 (N_8786,N_8643,N_8633);
nor U8787 (N_8787,N_8677,N_8620);
and U8788 (N_8788,N_8607,N_8650);
nor U8789 (N_8789,N_8618,N_8678);
nand U8790 (N_8790,N_8571,N_8619);
nand U8791 (N_8791,N_8601,N_8551);
nand U8792 (N_8792,N_8608,N_8649);
and U8793 (N_8793,N_8582,N_8562);
xnor U8794 (N_8794,N_8557,N_8561);
or U8795 (N_8795,N_8671,N_8683);
nand U8796 (N_8796,N_8606,N_8664);
or U8797 (N_8797,N_8553,N_8652);
nor U8798 (N_8798,N_8692,N_8551);
nor U8799 (N_8799,N_8661,N_8578);
or U8800 (N_8800,N_8689,N_8584);
nand U8801 (N_8801,N_8663,N_8697);
nand U8802 (N_8802,N_8571,N_8563);
nor U8803 (N_8803,N_8684,N_8558);
nor U8804 (N_8804,N_8682,N_8683);
or U8805 (N_8805,N_8607,N_8612);
nor U8806 (N_8806,N_8694,N_8693);
and U8807 (N_8807,N_8615,N_8693);
xor U8808 (N_8808,N_8593,N_8672);
and U8809 (N_8809,N_8636,N_8620);
nor U8810 (N_8810,N_8641,N_8626);
nor U8811 (N_8811,N_8626,N_8673);
or U8812 (N_8812,N_8633,N_8668);
and U8813 (N_8813,N_8660,N_8632);
or U8814 (N_8814,N_8643,N_8639);
or U8815 (N_8815,N_8683,N_8614);
nand U8816 (N_8816,N_8656,N_8609);
nand U8817 (N_8817,N_8656,N_8576);
nand U8818 (N_8818,N_8676,N_8679);
and U8819 (N_8819,N_8626,N_8577);
nor U8820 (N_8820,N_8601,N_8679);
or U8821 (N_8821,N_8692,N_8600);
xor U8822 (N_8822,N_8554,N_8662);
xnor U8823 (N_8823,N_8598,N_8627);
xnor U8824 (N_8824,N_8694,N_8574);
xor U8825 (N_8825,N_8643,N_8692);
xnor U8826 (N_8826,N_8604,N_8553);
or U8827 (N_8827,N_8639,N_8657);
and U8828 (N_8828,N_8694,N_8686);
and U8829 (N_8829,N_8563,N_8682);
xnor U8830 (N_8830,N_8693,N_8575);
or U8831 (N_8831,N_8699,N_8692);
or U8832 (N_8832,N_8678,N_8580);
or U8833 (N_8833,N_8684,N_8675);
nor U8834 (N_8834,N_8646,N_8605);
nor U8835 (N_8835,N_8656,N_8600);
xor U8836 (N_8836,N_8591,N_8564);
and U8837 (N_8837,N_8661,N_8558);
or U8838 (N_8838,N_8589,N_8550);
xor U8839 (N_8839,N_8576,N_8677);
nor U8840 (N_8840,N_8647,N_8685);
and U8841 (N_8841,N_8684,N_8579);
nor U8842 (N_8842,N_8675,N_8618);
nor U8843 (N_8843,N_8608,N_8555);
or U8844 (N_8844,N_8597,N_8662);
nor U8845 (N_8845,N_8630,N_8672);
and U8846 (N_8846,N_8606,N_8588);
nand U8847 (N_8847,N_8616,N_8580);
nand U8848 (N_8848,N_8676,N_8554);
nand U8849 (N_8849,N_8679,N_8680);
and U8850 (N_8850,N_8748,N_8792);
or U8851 (N_8851,N_8712,N_8831);
xor U8852 (N_8852,N_8846,N_8807);
or U8853 (N_8853,N_8710,N_8827);
nor U8854 (N_8854,N_8845,N_8772);
and U8855 (N_8855,N_8821,N_8787);
xnor U8856 (N_8856,N_8747,N_8711);
nand U8857 (N_8857,N_8806,N_8797);
or U8858 (N_8858,N_8840,N_8804);
nand U8859 (N_8859,N_8795,N_8733);
nor U8860 (N_8860,N_8829,N_8836);
nand U8861 (N_8861,N_8734,N_8841);
and U8862 (N_8862,N_8774,N_8702);
nor U8863 (N_8863,N_8781,N_8720);
nand U8864 (N_8864,N_8833,N_8713);
nor U8865 (N_8865,N_8732,N_8849);
xnor U8866 (N_8866,N_8761,N_8729);
nor U8867 (N_8867,N_8718,N_8763);
or U8868 (N_8868,N_8701,N_8791);
or U8869 (N_8869,N_8750,N_8819);
and U8870 (N_8870,N_8728,N_8751);
or U8871 (N_8871,N_8758,N_8842);
nor U8872 (N_8872,N_8796,N_8768);
nand U8873 (N_8873,N_8838,N_8706);
xor U8874 (N_8874,N_8779,N_8808);
nand U8875 (N_8875,N_8805,N_8783);
xnor U8876 (N_8876,N_8752,N_8730);
nor U8877 (N_8877,N_8812,N_8746);
nor U8878 (N_8878,N_8739,N_8832);
or U8879 (N_8879,N_8816,N_8790);
and U8880 (N_8880,N_8755,N_8828);
xnor U8881 (N_8881,N_8707,N_8731);
or U8882 (N_8882,N_8737,N_8715);
nand U8883 (N_8883,N_8834,N_8825);
and U8884 (N_8884,N_8843,N_8709);
and U8885 (N_8885,N_8817,N_8724);
nand U8886 (N_8886,N_8723,N_8784);
or U8887 (N_8887,N_8800,N_8844);
or U8888 (N_8888,N_8818,N_8754);
nand U8889 (N_8889,N_8837,N_8738);
nor U8890 (N_8890,N_8810,N_8740);
xor U8891 (N_8891,N_8786,N_8704);
nand U8892 (N_8892,N_8764,N_8802);
and U8893 (N_8893,N_8700,N_8780);
and U8894 (N_8894,N_8741,N_8789);
or U8895 (N_8895,N_8756,N_8744);
nand U8896 (N_8896,N_8839,N_8820);
or U8897 (N_8897,N_8703,N_8815);
and U8898 (N_8898,N_8771,N_8778);
or U8899 (N_8899,N_8826,N_8813);
xor U8900 (N_8900,N_8777,N_8801);
or U8901 (N_8901,N_8794,N_8766);
nand U8902 (N_8902,N_8770,N_8762);
nor U8903 (N_8903,N_8705,N_8822);
nor U8904 (N_8904,N_8708,N_8799);
nand U8905 (N_8905,N_8830,N_8725);
xnor U8906 (N_8906,N_8823,N_8760);
or U8907 (N_8907,N_8798,N_8735);
nor U8908 (N_8908,N_8736,N_8785);
nor U8909 (N_8909,N_8726,N_8714);
xnor U8910 (N_8910,N_8775,N_8773);
xor U8911 (N_8911,N_8835,N_8793);
and U8912 (N_8912,N_8753,N_8722);
and U8913 (N_8913,N_8716,N_8814);
nand U8914 (N_8914,N_8824,N_8765);
or U8915 (N_8915,N_8767,N_8742);
and U8916 (N_8916,N_8719,N_8759);
nor U8917 (N_8917,N_8743,N_8803);
and U8918 (N_8918,N_8749,N_8721);
or U8919 (N_8919,N_8782,N_8717);
nand U8920 (N_8920,N_8776,N_8809);
and U8921 (N_8921,N_8811,N_8788);
xnor U8922 (N_8922,N_8848,N_8745);
nor U8923 (N_8923,N_8757,N_8727);
or U8924 (N_8924,N_8769,N_8847);
or U8925 (N_8925,N_8848,N_8715);
or U8926 (N_8926,N_8828,N_8712);
nand U8927 (N_8927,N_8712,N_8827);
nor U8928 (N_8928,N_8778,N_8849);
xor U8929 (N_8929,N_8708,N_8719);
and U8930 (N_8930,N_8765,N_8766);
and U8931 (N_8931,N_8848,N_8765);
xnor U8932 (N_8932,N_8723,N_8773);
xnor U8933 (N_8933,N_8789,N_8731);
and U8934 (N_8934,N_8791,N_8811);
nor U8935 (N_8935,N_8713,N_8759);
nor U8936 (N_8936,N_8828,N_8763);
nor U8937 (N_8937,N_8838,N_8779);
xnor U8938 (N_8938,N_8820,N_8710);
and U8939 (N_8939,N_8737,N_8845);
or U8940 (N_8940,N_8752,N_8756);
nand U8941 (N_8941,N_8720,N_8785);
or U8942 (N_8942,N_8817,N_8835);
nor U8943 (N_8943,N_8772,N_8808);
or U8944 (N_8944,N_8746,N_8744);
xnor U8945 (N_8945,N_8819,N_8777);
nand U8946 (N_8946,N_8811,N_8734);
or U8947 (N_8947,N_8831,N_8731);
nor U8948 (N_8948,N_8725,N_8806);
and U8949 (N_8949,N_8842,N_8834);
nand U8950 (N_8950,N_8762,N_8806);
nand U8951 (N_8951,N_8738,N_8706);
nor U8952 (N_8952,N_8742,N_8795);
xnor U8953 (N_8953,N_8824,N_8775);
nor U8954 (N_8954,N_8815,N_8784);
nor U8955 (N_8955,N_8733,N_8707);
nand U8956 (N_8956,N_8814,N_8837);
xnor U8957 (N_8957,N_8780,N_8755);
nor U8958 (N_8958,N_8765,N_8733);
xnor U8959 (N_8959,N_8798,N_8750);
nand U8960 (N_8960,N_8763,N_8706);
and U8961 (N_8961,N_8804,N_8841);
nor U8962 (N_8962,N_8826,N_8806);
nor U8963 (N_8963,N_8742,N_8807);
nor U8964 (N_8964,N_8749,N_8718);
nand U8965 (N_8965,N_8745,N_8711);
or U8966 (N_8966,N_8750,N_8767);
xor U8967 (N_8967,N_8729,N_8751);
nor U8968 (N_8968,N_8749,N_8793);
nor U8969 (N_8969,N_8733,N_8770);
nor U8970 (N_8970,N_8733,N_8753);
nand U8971 (N_8971,N_8792,N_8843);
xor U8972 (N_8972,N_8745,N_8755);
or U8973 (N_8973,N_8700,N_8827);
xor U8974 (N_8974,N_8822,N_8826);
xnor U8975 (N_8975,N_8791,N_8802);
nand U8976 (N_8976,N_8848,N_8767);
nor U8977 (N_8977,N_8846,N_8703);
or U8978 (N_8978,N_8724,N_8745);
and U8979 (N_8979,N_8839,N_8771);
or U8980 (N_8980,N_8771,N_8814);
and U8981 (N_8981,N_8739,N_8732);
or U8982 (N_8982,N_8829,N_8751);
and U8983 (N_8983,N_8798,N_8763);
xor U8984 (N_8984,N_8815,N_8824);
nand U8985 (N_8985,N_8848,N_8795);
and U8986 (N_8986,N_8703,N_8766);
xor U8987 (N_8987,N_8816,N_8765);
xnor U8988 (N_8988,N_8810,N_8728);
and U8989 (N_8989,N_8756,N_8732);
nor U8990 (N_8990,N_8838,N_8778);
nand U8991 (N_8991,N_8822,N_8815);
nor U8992 (N_8992,N_8725,N_8714);
nand U8993 (N_8993,N_8849,N_8760);
xnor U8994 (N_8994,N_8764,N_8776);
nor U8995 (N_8995,N_8833,N_8759);
xor U8996 (N_8996,N_8801,N_8838);
xnor U8997 (N_8997,N_8761,N_8819);
nor U8998 (N_8998,N_8743,N_8732);
xor U8999 (N_8999,N_8746,N_8745);
and U9000 (N_9000,N_8961,N_8933);
nand U9001 (N_9001,N_8926,N_8900);
or U9002 (N_9002,N_8936,N_8884);
or U9003 (N_9003,N_8937,N_8990);
or U9004 (N_9004,N_8890,N_8927);
and U9005 (N_9005,N_8942,N_8941);
or U9006 (N_9006,N_8921,N_8995);
or U9007 (N_9007,N_8932,N_8973);
nor U9008 (N_9008,N_8859,N_8969);
nand U9009 (N_9009,N_8910,N_8914);
and U9010 (N_9010,N_8875,N_8863);
xnor U9011 (N_9011,N_8905,N_8950);
nand U9012 (N_9012,N_8966,N_8982);
and U9013 (N_9013,N_8899,N_8864);
and U9014 (N_9014,N_8882,N_8984);
nand U9015 (N_9015,N_8851,N_8949);
nand U9016 (N_9016,N_8868,N_8869);
nand U9017 (N_9017,N_8971,N_8871);
nor U9018 (N_9018,N_8935,N_8887);
nand U9019 (N_9019,N_8893,N_8854);
nor U9020 (N_9020,N_8979,N_8852);
and U9021 (N_9021,N_8931,N_8872);
nand U9022 (N_9022,N_8881,N_8976);
nand U9023 (N_9023,N_8867,N_8934);
nand U9024 (N_9024,N_8994,N_8960);
nor U9025 (N_9025,N_8962,N_8860);
nor U9026 (N_9026,N_8904,N_8930);
nand U9027 (N_9027,N_8873,N_8878);
nand U9028 (N_9028,N_8891,N_8876);
nand U9029 (N_9029,N_8958,N_8968);
or U9030 (N_9030,N_8929,N_8922);
nor U9031 (N_9031,N_8879,N_8855);
xor U9032 (N_9032,N_8894,N_8877);
nor U9033 (N_9033,N_8943,N_8870);
and U9034 (N_9034,N_8858,N_8957);
or U9035 (N_9035,N_8948,N_8896);
xnor U9036 (N_9036,N_8883,N_8997);
nand U9037 (N_9037,N_8917,N_8902);
nor U9038 (N_9038,N_8951,N_8866);
or U9039 (N_9039,N_8985,N_8928);
nand U9040 (N_9040,N_8944,N_8956);
and U9041 (N_9041,N_8987,N_8964);
nor U9042 (N_9042,N_8919,N_8912);
xor U9043 (N_9043,N_8939,N_8998);
nor U9044 (N_9044,N_8888,N_8978);
or U9045 (N_9045,N_8913,N_8974);
nor U9046 (N_9046,N_8983,N_8980);
or U9047 (N_9047,N_8856,N_8850);
nand U9048 (N_9048,N_8924,N_8963);
and U9049 (N_9049,N_8925,N_8909);
nand U9050 (N_9050,N_8898,N_8901);
nand U9051 (N_9051,N_8947,N_8938);
or U9052 (N_9052,N_8853,N_8996);
nor U9053 (N_9053,N_8916,N_8986);
or U9054 (N_9054,N_8885,N_8874);
xor U9055 (N_9055,N_8999,N_8865);
nand U9056 (N_9056,N_8923,N_8907);
nor U9057 (N_9057,N_8940,N_8895);
nand U9058 (N_9058,N_8857,N_8908);
and U9059 (N_9059,N_8988,N_8897);
and U9060 (N_9060,N_8945,N_8903);
nand U9061 (N_9061,N_8861,N_8946);
nor U9062 (N_9062,N_8970,N_8981);
xor U9063 (N_9063,N_8862,N_8892);
nand U9064 (N_9064,N_8918,N_8915);
and U9065 (N_9065,N_8952,N_8886);
xor U9066 (N_9066,N_8975,N_8959);
xnor U9067 (N_9067,N_8906,N_8977);
or U9068 (N_9068,N_8993,N_8953);
or U9069 (N_9069,N_8920,N_8989);
nor U9070 (N_9070,N_8965,N_8972);
xor U9071 (N_9071,N_8992,N_8955);
and U9072 (N_9072,N_8889,N_8911);
xor U9073 (N_9073,N_8991,N_8967);
or U9074 (N_9074,N_8880,N_8954);
xor U9075 (N_9075,N_8942,N_8877);
xnor U9076 (N_9076,N_8855,N_8884);
or U9077 (N_9077,N_8860,N_8959);
nor U9078 (N_9078,N_8888,N_8859);
and U9079 (N_9079,N_8940,N_8874);
nand U9080 (N_9080,N_8970,N_8989);
xor U9081 (N_9081,N_8920,N_8961);
nor U9082 (N_9082,N_8894,N_8932);
nor U9083 (N_9083,N_8865,N_8985);
and U9084 (N_9084,N_8880,N_8929);
or U9085 (N_9085,N_8871,N_8976);
and U9086 (N_9086,N_8966,N_8922);
or U9087 (N_9087,N_8968,N_8941);
and U9088 (N_9088,N_8900,N_8967);
xnor U9089 (N_9089,N_8983,N_8994);
or U9090 (N_9090,N_8978,N_8954);
xnor U9091 (N_9091,N_8862,N_8993);
nor U9092 (N_9092,N_8879,N_8884);
xor U9093 (N_9093,N_8969,N_8868);
nor U9094 (N_9094,N_8970,N_8878);
nor U9095 (N_9095,N_8976,N_8910);
xnor U9096 (N_9096,N_8916,N_8884);
xnor U9097 (N_9097,N_8900,N_8987);
or U9098 (N_9098,N_8941,N_8862);
nand U9099 (N_9099,N_8872,N_8987);
nand U9100 (N_9100,N_8992,N_8961);
xor U9101 (N_9101,N_8986,N_8908);
or U9102 (N_9102,N_8937,N_8905);
and U9103 (N_9103,N_8986,N_8865);
xnor U9104 (N_9104,N_8976,N_8878);
xor U9105 (N_9105,N_8952,N_8989);
and U9106 (N_9106,N_8859,N_8912);
and U9107 (N_9107,N_8913,N_8985);
nor U9108 (N_9108,N_8934,N_8860);
or U9109 (N_9109,N_8945,N_8957);
xnor U9110 (N_9110,N_8941,N_8893);
or U9111 (N_9111,N_8932,N_8875);
xor U9112 (N_9112,N_8972,N_8885);
nor U9113 (N_9113,N_8977,N_8937);
and U9114 (N_9114,N_8904,N_8914);
xnor U9115 (N_9115,N_8956,N_8941);
nor U9116 (N_9116,N_8992,N_8985);
xnor U9117 (N_9117,N_8879,N_8874);
or U9118 (N_9118,N_8886,N_8993);
nand U9119 (N_9119,N_8958,N_8892);
and U9120 (N_9120,N_8859,N_8899);
nand U9121 (N_9121,N_8997,N_8900);
nor U9122 (N_9122,N_8877,N_8863);
nor U9123 (N_9123,N_8885,N_8990);
or U9124 (N_9124,N_8983,N_8981);
nor U9125 (N_9125,N_8967,N_8901);
and U9126 (N_9126,N_8933,N_8964);
nor U9127 (N_9127,N_8999,N_8980);
nor U9128 (N_9128,N_8911,N_8880);
nand U9129 (N_9129,N_8972,N_8974);
or U9130 (N_9130,N_8993,N_8991);
xor U9131 (N_9131,N_8880,N_8983);
or U9132 (N_9132,N_8852,N_8916);
nor U9133 (N_9133,N_8866,N_8881);
nand U9134 (N_9134,N_8875,N_8887);
or U9135 (N_9135,N_8882,N_8896);
and U9136 (N_9136,N_8898,N_8946);
nand U9137 (N_9137,N_8916,N_8892);
and U9138 (N_9138,N_8956,N_8884);
nor U9139 (N_9139,N_8932,N_8955);
nor U9140 (N_9140,N_8943,N_8878);
nor U9141 (N_9141,N_8963,N_8919);
and U9142 (N_9142,N_8857,N_8873);
nor U9143 (N_9143,N_8862,N_8856);
or U9144 (N_9144,N_8961,N_8926);
nand U9145 (N_9145,N_8876,N_8908);
xor U9146 (N_9146,N_8975,N_8860);
or U9147 (N_9147,N_8877,N_8885);
and U9148 (N_9148,N_8920,N_8982);
or U9149 (N_9149,N_8873,N_8941);
nand U9150 (N_9150,N_9023,N_9087);
and U9151 (N_9151,N_9003,N_9054);
nor U9152 (N_9152,N_9081,N_9124);
xnor U9153 (N_9153,N_9016,N_9102);
xnor U9154 (N_9154,N_9083,N_9004);
or U9155 (N_9155,N_9138,N_9093);
nand U9156 (N_9156,N_9085,N_9105);
or U9157 (N_9157,N_9026,N_9106);
and U9158 (N_9158,N_9049,N_9052);
xnor U9159 (N_9159,N_9019,N_9103);
or U9160 (N_9160,N_9134,N_9065);
or U9161 (N_9161,N_9009,N_9128);
nor U9162 (N_9162,N_9060,N_9114);
or U9163 (N_9163,N_9110,N_9121);
or U9164 (N_9164,N_9127,N_9118);
and U9165 (N_9165,N_9047,N_9012);
or U9166 (N_9166,N_9001,N_9045);
nand U9167 (N_9167,N_9139,N_9013);
nor U9168 (N_9168,N_9039,N_9082);
or U9169 (N_9169,N_9064,N_9090);
or U9170 (N_9170,N_9107,N_9108);
and U9171 (N_9171,N_9066,N_9020);
xnor U9172 (N_9172,N_9041,N_9100);
nand U9173 (N_9173,N_9069,N_9046);
or U9174 (N_9174,N_9006,N_9131);
nor U9175 (N_9175,N_9002,N_9077);
and U9176 (N_9176,N_9099,N_9068);
nor U9177 (N_9177,N_9115,N_9089);
and U9178 (N_9178,N_9050,N_9112);
and U9179 (N_9179,N_9126,N_9148);
nor U9180 (N_9180,N_9141,N_9101);
and U9181 (N_9181,N_9059,N_9030);
nor U9182 (N_9182,N_9043,N_9145);
nor U9183 (N_9183,N_9007,N_9074);
nand U9184 (N_9184,N_9117,N_9036);
and U9185 (N_9185,N_9008,N_9031);
nand U9186 (N_9186,N_9011,N_9079);
and U9187 (N_9187,N_9129,N_9146);
or U9188 (N_9188,N_9073,N_9057);
or U9189 (N_9189,N_9092,N_9072);
or U9190 (N_9190,N_9097,N_9123);
or U9191 (N_9191,N_9080,N_9048);
or U9192 (N_9192,N_9125,N_9042);
nand U9193 (N_9193,N_9096,N_9051);
nand U9194 (N_9194,N_9076,N_9062);
xnor U9195 (N_9195,N_9022,N_9005);
xor U9196 (N_9196,N_9130,N_9063);
xor U9197 (N_9197,N_9071,N_9109);
nand U9198 (N_9198,N_9142,N_9143);
or U9199 (N_9199,N_9119,N_9037);
xnor U9200 (N_9200,N_9104,N_9040);
xnor U9201 (N_9201,N_9133,N_9014);
nand U9202 (N_9202,N_9018,N_9044);
nand U9203 (N_9203,N_9135,N_9034);
or U9204 (N_9204,N_9095,N_9113);
or U9205 (N_9205,N_9078,N_9025);
or U9206 (N_9206,N_9010,N_9056);
or U9207 (N_9207,N_9024,N_9144);
or U9208 (N_9208,N_9091,N_9111);
xnor U9209 (N_9209,N_9029,N_9035);
nor U9210 (N_9210,N_9021,N_9028);
and U9211 (N_9211,N_9075,N_9116);
nor U9212 (N_9212,N_9067,N_9147);
and U9213 (N_9213,N_9061,N_9086);
nand U9214 (N_9214,N_9033,N_9058);
or U9215 (N_9215,N_9088,N_9084);
xor U9216 (N_9216,N_9017,N_9120);
xnor U9217 (N_9217,N_9149,N_9070);
nor U9218 (N_9218,N_9132,N_9137);
and U9219 (N_9219,N_9094,N_9027);
and U9220 (N_9220,N_9136,N_9032);
nor U9221 (N_9221,N_9053,N_9140);
and U9222 (N_9222,N_9055,N_9038);
or U9223 (N_9223,N_9000,N_9122);
nor U9224 (N_9224,N_9098,N_9015);
nor U9225 (N_9225,N_9090,N_9005);
xnor U9226 (N_9226,N_9129,N_9147);
or U9227 (N_9227,N_9087,N_9112);
nor U9228 (N_9228,N_9069,N_9029);
nand U9229 (N_9229,N_9075,N_9125);
xnor U9230 (N_9230,N_9074,N_9101);
nor U9231 (N_9231,N_9100,N_9078);
xor U9232 (N_9232,N_9042,N_9045);
xor U9233 (N_9233,N_9060,N_9025);
and U9234 (N_9234,N_9068,N_9147);
xnor U9235 (N_9235,N_9104,N_9108);
nand U9236 (N_9236,N_9060,N_9142);
nand U9237 (N_9237,N_9006,N_9073);
or U9238 (N_9238,N_9048,N_9122);
nor U9239 (N_9239,N_9112,N_9109);
nand U9240 (N_9240,N_9042,N_9005);
and U9241 (N_9241,N_9069,N_9075);
nor U9242 (N_9242,N_9072,N_9139);
or U9243 (N_9243,N_9053,N_9030);
nor U9244 (N_9244,N_9031,N_9104);
nor U9245 (N_9245,N_9104,N_9145);
nand U9246 (N_9246,N_9113,N_9010);
and U9247 (N_9247,N_9110,N_9062);
and U9248 (N_9248,N_9071,N_9007);
xor U9249 (N_9249,N_9067,N_9137);
or U9250 (N_9250,N_9108,N_9134);
nor U9251 (N_9251,N_9148,N_9082);
nand U9252 (N_9252,N_9016,N_9123);
xnor U9253 (N_9253,N_9043,N_9014);
or U9254 (N_9254,N_9115,N_9012);
nor U9255 (N_9255,N_9034,N_9095);
or U9256 (N_9256,N_9091,N_9013);
xor U9257 (N_9257,N_9033,N_9056);
nor U9258 (N_9258,N_9004,N_9088);
nor U9259 (N_9259,N_9146,N_9131);
nand U9260 (N_9260,N_9114,N_9067);
or U9261 (N_9261,N_9133,N_9017);
and U9262 (N_9262,N_9115,N_9103);
xnor U9263 (N_9263,N_9122,N_9087);
nand U9264 (N_9264,N_9088,N_9081);
and U9265 (N_9265,N_9069,N_9130);
xnor U9266 (N_9266,N_9028,N_9133);
nand U9267 (N_9267,N_9139,N_9056);
nand U9268 (N_9268,N_9061,N_9101);
or U9269 (N_9269,N_9033,N_9091);
nand U9270 (N_9270,N_9027,N_9074);
nand U9271 (N_9271,N_9094,N_9007);
nand U9272 (N_9272,N_9078,N_9040);
xor U9273 (N_9273,N_9110,N_9020);
nand U9274 (N_9274,N_9131,N_9132);
xor U9275 (N_9275,N_9079,N_9101);
or U9276 (N_9276,N_9108,N_9040);
nor U9277 (N_9277,N_9044,N_9116);
nor U9278 (N_9278,N_9019,N_9077);
nand U9279 (N_9279,N_9089,N_9016);
nand U9280 (N_9280,N_9117,N_9061);
or U9281 (N_9281,N_9055,N_9134);
and U9282 (N_9282,N_9043,N_9102);
nor U9283 (N_9283,N_9069,N_9146);
xor U9284 (N_9284,N_9143,N_9116);
nor U9285 (N_9285,N_9077,N_9124);
nand U9286 (N_9286,N_9042,N_9095);
xor U9287 (N_9287,N_9046,N_9106);
nor U9288 (N_9288,N_9062,N_9113);
and U9289 (N_9289,N_9139,N_9006);
or U9290 (N_9290,N_9025,N_9000);
xor U9291 (N_9291,N_9088,N_9040);
or U9292 (N_9292,N_9108,N_9015);
nand U9293 (N_9293,N_9008,N_9102);
xnor U9294 (N_9294,N_9025,N_9013);
or U9295 (N_9295,N_9020,N_9133);
nor U9296 (N_9296,N_9019,N_9129);
xor U9297 (N_9297,N_9121,N_9049);
and U9298 (N_9298,N_9010,N_9070);
and U9299 (N_9299,N_9083,N_9131);
xor U9300 (N_9300,N_9151,N_9209);
xor U9301 (N_9301,N_9285,N_9264);
or U9302 (N_9302,N_9188,N_9215);
nand U9303 (N_9303,N_9197,N_9171);
nand U9304 (N_9304,N_9210,N_9168);
xor U9305 (N_9305,N_9225,N_9177);
xor U9306 (N_9306,N_9218,N_9241);
xnor U9307 (N_9307,N_9274,N_9253);
xor U9308 (N_9308,N_9292,N_9262);
or U9309 (N_9309,N_9206,N_9170);
xnor U9310 (N_9310,N_9265,N_9259);
and U9311 (N_9311,N_9266,N_9261);
xnor U9312 (N_9312,N_9243,N_9165);
nor U9313 (N_9313,N_9228,N_9257);
and U9314 (N_9314,N_9169,N_9247);
and U9315 (N_9315,N_9273,N_9217);
xnor U9316 (N_9316,N_9186,N_9175);
and U9317 (N_9317,N_9258,N_9270);
nor U9318 (N_9318,N_9182,N_9154);
nor U9319 (N_9319,N_9211,N_9296);
nand U9320 (N_9320,N_9254,N_9208);
or U9321 (N_9321,N_9160,N_9157);
and U9322 (N_9322,N_9181,N_9167);
nand U9323 (N_9323,N_9189,N_9267);
and U9324 (N_9324,N_9194,N_9248);
nand U9325 (N_9325,N_9179,N_9230);
nand U9326 (N_9326,N_9176,N_9180);
nor U9327 (N_9327,N_9293,N_9224);
nor U9328 (N_9328,N_9203,N_9185);
and U9329 (N_9329,N_9164,N_9271);
and U9330 (N_9330,N_9299,N_9159);
or U9331 (N_9331,N_9289,N_9213);
nand U9332 (N_9332,N_9227,N_9174);
nand U9333 (N_9333,N_9260,N_9178);
or U9334 (N_9334,N_9190,N_9288);
nand U9335 (N_9335,N_9237,N_9163);
and U9336 (N_9336,N_9193,N_9232);
xor U9337 (N_9337,N_9278,N_9161);
nor U9338 (N_9338,N_9269,N_9226);
xor U9339 (N_9339,N_9279,N_9295);
nor U9340 (N_9340,N_9242,N_9240);
and U9341 (N_9341,N_9184,N_9195);
nand U9342 (N_9342,N_9239,N_9287);
or U9343 (N_9343,N_9276,N_9198);
nor U9344 (N_9344,N_9272,N_9155);
nand U9345 (N_9345,N_9246,N_9238);
and U9346 (N_9346,N_9234,N_9249);
nor U9347 (N_9347,N_9191,N_9219);
nand U9348 (N_9348,N_9212,N_9256);
xnor U9349 (N_9349,N_9173,N_9290);
xnor U9350 (N_9350,N_9220,N_9156);
xnor U9351 (N_9351,N_9207,N_9281);
xnor U9352 (N_9352,N_9268,N_9152);
nand U9353 (N_9353,N_9221,N_9283);
or U9354 (N_9354,N_9294,N_9150);
nor U9355 (N_9355,N_9199,N_9205);
or U9356 (N_9356,N_9251,N_9231);
xor U9357 (N_9357,N_9216,N_9236);
xnor U9358 (N_9358,N_9204,N_9153);
and U9359 (N_9359,N_9183,N_9192);
nand U9360 (N_9360,N_9223,N_9297);
nand U9361 (N_9361,N_9166,N_9187);
or U9362 (N_9362,N_9222,N_9214);
nand U9363 (N_9363,N_9250,N_9172);
xnor U9364 (N_9364,N_9275,N_9233);
nand U9365 (N_9365,N_9201,N_9291);
nand U9366 (N_9366,N_9280,N_9158);
xnor U9367 (N_9367,N_9229,N_9244);
or U9368 (N_9368,N_9298,N_9282);
or U9369 (N_9369,N_9255,N_9286);
nand U9370 (N_9370,N_9245,N_9284);
or U9371 (N_9371,N_9162,N_9202);
xnor U9372 (N_9372,N_9277,N_9200);
xnor U9373 (N_9373,N_9252,N_9263);
or U9374 (N_9374,N_9196,N_9235);
or U9375 (N_9375,N_9239,N_9220);
nand U9376 (N_9376,N_9208,N_9209);
and U9377 (N_9377,N_9223,N_9150);
nand U9378 (N_9378,N_9197,N_9220);
nor U9379 (N_9379,N_9252,N_9270);
xnor U9380 (N_9380,N_9197,N_9238);
nand U9381 (N_9381,N_9234,N_9261);
nand U9382 (N_9382,N_9203,N_9218);
xnor U9383 (N_9383,N_9283,N_9222);
xor U9384 (N_9384,N_9274,N_9226);
xor U9385 (N_9385,N_9281,N_9201);
xor U9386 (N_9386,N_9282,N_9265);
xor U9387 (N_9387,N_9231,N_9252);
nor U9388 (N_9388,N_9200,N_9164);
nor U9389 (N_9389,N_9265,N_9285);
nand U9390 (N_9390,N_9211,N_9156);
nor U9391 (N_9391,N_9248,N_9295);
nor U9392 (N_9392,N_9247,N_9171);
and U9393 (N_9393,N_9170,N_9298);
xnor U9394 (N_9394,N_9224,N_9176);
xnor U9395 (N_9395,N_9205,N_9221);
or U9396 (N_9396,N_9221,N_9235);
and U9397 (N_9397,N_9254,N_9270);
nand U9398 (N_9398,N_9210,N_9266);
xnor U9399 (N_9399,N_9265,N_9220);
nand U9400 (N_9400,N_9200,N_9219);
and U9401 (N_9401,N_9281,N_9172);
xnor U9402 (N_9402,N_9210,N_9187);
nand U9403 (N_9403,N_9240,N_9219);
xnor U9404 (N_9404,N_9296,N_9249);
or U9405 (N_9405,N_9235,N_9243);
nor U9406 (N_9406,N_9264,N_9244);
or U9407 (N_9407,N_9285,N_9177);
or U9408 (N_9408,N_9194,N_9170);
or U9409 (N_9409,N_9276,N_9294);
and U9410 (N_9410,N_9279,N_9231);
xnor U9411 (N_9411,N_9291,N_9250);
and U9412 (N_9412,N_9227,N_9287);
nand U9413 (N_9413,N_9179,N_9236);
or U9414 (N_9414,N_9163,N_9243);
and U9415 (N_9415,N_9270,N_9155);
or U9416 (N_9416,N_9177,N_9153);
xor U9417 (N_9417,N_9283,N_9213);
xnor U9418 (N_9418,N_9182,N_9191);
or U9419 (N_9419,N_9269,N_9184);
or U9420 (N_9420,N_9240,N_9174);
and U9421 (N_9421,N_9169,N_9228);
xnor U9422 (N_9422,N_9226,N_9262);
xnor U9423 (N_9423,N_9207,N_9167);
nand U9424 (N_9424,N_9287,N_9168);
nand U9425 (N_9425,N_9288,N_9269);
and U9426 (N_9426,N_9179,N_9188);
and U9427 (N_9427,N_9268,N_9297);
and U9428 (N_9428,N_9279,N_9200);
xnor U9429 (N_9429,N_9212,N_9174);
nor U9430 (N_9430,N_9165,N_9192);
nor U9431 (N_9431,N_9252,N_9186);
xor U9432 (N_9432,N_9160,N_9183);
nor U9433 (N_9433,N_9265,N_9163);
and U9434 (N_9434,N_9284,N_9156);
or U9435 (N_9435,N_9155,N_9170);
xor U9436 (N_9436,N_9233,N_9298);
or U9437 (N_9437,N_9152,N_9265);
or U9438 (N_9438,N_9296,N_9234);
nand U9439 (N_9439,N_9249,N_9223);
nand U9440 (N_9440,N_9205,N_9235);
or U9441 (N_9441,N_9203,N_9238);
nand U9442 (N_9442,N_9233,N_9271);
and U9443 (N_9443,N_9286,N_9163);
or U9444 (N_9444,N_9210,N_9220);
nand U9445 (N_9445,N_9162,N_9195);
nor U9446 (N_9446,N_9176,N_9190);
nor U9447 (N_9447,N_9215,N_9255);
or U9448 (N_9448,N_9291,N_9192);
and U9449 (N_9449,N_9252,N_9241);
nand U9450 (N_9450,N_9412,N_9375);
nor U9451 (N_9451,N_9388,N_9409);
nand U9452 (N_9452,N_9323,N_9318);
nand U9453 (N_9453,N_9377,N_9354);
nand U9454 (N_9454,N_9414,N_9327);
or U9455 (N_9455,N_9366,N_9398);
nand U9456 (N_9456,N_9405,N_9333);
nand U9457 (N_9457,N_9345,N_9433);
or U9458 (N_9458,N_9313,N_9352);
nand U9459 (N_9459,N_9426,N_9332);
xnor U9460 (N_9460,N_9419,N_9404);
nor U9461 (N_9461,N_9307,N_9413);
xnor U9462 (N_9462,N_9309,N_9379);
and U9463 (N_9463,N_9342,N_9306);
nand U9464 (N_9464,N_9384,N_9365);
or U9465 (N_9465,N_9401,N_9382);
nor U9466 (N_9466,N_9374,N_9443);
xor U9467 (N_9467,N_9320,N_9344);
xor U9468 (N_9468,N_9300,N_9407);
or U9469 (N_9469,N_9326,N_9429);
nor U9470 (N_9470,N_9370,N_9302);
nand U9471 (N_9471,N_9380,N_9403);
or U9472 (N_9472,N_9303,N_9317);
xnor U9473 (N_9473,N_9340,N_9315);
or U9474 (N_9474,N_9434,N_9329);
nand U9475 (N_9475,N_9325,N_9408);
nand U9476 (N_9476,N_9301,N_9449);
nand U9477 (N_9477,N_9362,N_9397);
nor U9478 (N_9478,N_9436,N_9319);
and U9479 (N_9479,N_9438,N_9421);
nor U9480 (N_9480,N_9439,N_9328);
and U9481 (N_9481,N_9394,N_9410);
or U9482 (N_9482,N_9311,N_9361);
or U9483 (N_9483,N_9314,N_9444);
xnor U9484 (N_9484,N_9392,N_9396);
nand U9485 (N_9485,N_9348,N_9432);
nand U9486 (N_9486,N_9395,N_9339);
nand U9487 (N_9487,N_9381,N_9331);
nand U9488 (N_9488,N_9351,N_9341);
nor U9489 (N_9489,N_9446,N_9416);
nand U9490 (N_9490,N_9378,N_9371);
nor U9491 (N_9491,N_9393,N_9420);
and U9492 (N_9492,N_9383,N_9427);
xnor U9493 (N_9493,N_9338,N_9357);
xor U9494 (N_9494,N_9431,N_9355);
and U9495 (N_9495,N_9389,N_9418);
nand U9496 (N_9496,N_9402,N_9312);
nor U9497 (N_9497,N_9399,N_9445);
xnor U9498 (N_9498,N_9360,N_9447);
or U9499 (N_9499,N_9437,N_9425);
or U9500 (N_9500,N_9350,N_9334);
and U9501 (N_9501,N_9387,N_9390);
nor U9502 (N_9502,N_9347,N_9305);
xnor U9503 (N_9503,N_9415,N_9411);
or U9504 (N_9504,N_9424,N_9310);
and U9505 (N_9505,N_9346,N_9321);
or U9506 (N_9506,N_9336,N_9356);
nand U9507 (N_9507,N_9337,N_9442);
and U9508 (N_9508,N_9417,N_9423);
xor U9509 (N_9509,N_9308,N_9422);
nor U9510 (N_9510,N_9330,N_9304);
xnor U9511 (N_9511,N_9428,N_9359);
xor U9512 (N_9512,N_9343,N_9448);
or U9513 (N_9513,N_9353,N_9335);
xor U9514 (N_9514,N_9440,N_9367);
nand U9515 (N_9515,N_9400,N_9430);
and U9516 (N_9516,N_9358,N_9406);
nor U9517 (N_9517,N_9324,N_9376);
or U9518 (N_9518,N_9372,N_9435);
xnor U9519 (N_9519,N_9385,N_9369);
nor U9520 (N_9520,N_9349,N_9368);
and U9521 (N_9521,N_9364,N_9373);
or U9522 (N_9522,N_9386,N_9441);
nand U9523 (N_9523,N_9391,N_9322);
or U9524 (N_9524,N_9316,N_9363);
xor U9525 (N_9525,N_9337,N_9398);
or U9526 (N_9526,N_9391,N_9416);
nand U9527 (N_9527,N_9360,N_9419);
nor U9528 (N_9528,N_9430,N_9380);
xnor U9529 (N_9529,N_9350,N_9435);
nand U9530 (N_9530,N_9431,N_9352);
or U9531 (N_9531,N_9322,N_9419);
nor U9532 (N_9532,N_9395,N_9389);
and U9533 (N_9533,N_9403,N_9419);
and U9534 (N_9534,N_9325,N_9347);
nor U9535 (N_9535,N_9409,N_9428);
or U9536 (N_9536,N_9336,N_9445);
xnor U9537 (N_9537,N_9386,N_9390);
xor U9538 (N_9538,N_9328,N_9336);
nor U9539 (N_9539,N_9327,N_9373);
xor U9540 (N_9540,N_9416,N_9443);
and U9541 (N_9541,N_9393,N_9436);
nand U9542 (N_9542,N_9426,N_9444);
nand U9543 (N_9543,N_9358,N_9300);
and U9544 (N_9544,N_9444,N_9414);
or U9545 (N_9545,N_9372,N_9446);
nand U9546 (N_9546,N_9314,N_9437);
nor U9547 (N_9547,N_9328,N_9304);
nand U9548 (N_9548,N_9442,N_9310);
xor U9549 (N_9549,N_9313,N_9367);
or U9550 (N_9550,N_9405,N_9444);
or U9551 (N_9551,N_9361,N_9331);
nor U9552 (N_9552,N_9316,N_9366);
and U9553 (N_9553,N_9319,N_9334);
and U9554 (N_9554,N_9373,N_9368);
xor U9555 (N_9555,N_9443,N_9404);
and U9556 (N_9556,N_9328,N_9401);
nand U9557 (N_9557,N_9429,N_9434);
nor U9558 (N_9558,N_9434,N_9307);
nand U9559 (N_9559,N_9448,N_9381);
nor U9560 (N_9560,N_9307,N_9444);
and U9561 (N_9561,N_9364,N_9428);
xnor U9562 (N_9562,N_9391,N_9431);
nand U9563 (N_9563,N_9443,N_9338);
nand U9564 (N_9564,N_9310,N_9374);
nand U9565 (N_9565,N_9324,N_9430);
xnor U9566 (N_9566,N_9313,N_9429);
or U9567 (N_9567,N_9381,N_9340);
nor U9568 (N_9568,N_9350,N_9440);
nor U9569 (N_9569,N_9390,N_9435);
nor U9570 (N_9570,N_9333,N_9383);
nand U9571 (N_9571,N_9441,N_9424);
xnor U9572 (N_9572,N_9376,N_9446);
nand U9573 (N_9573,N_9407,N_9307);
nand U9574 (N_9574,N_9360,N_9394);
and U9575 (N_9575,N_9390,N_9406);
nand U9576 (N_9576,N_9405,N_9345);
xnor U9577 (N_9577,N_9319,N_9322);
nor U9578 (N_9578,N_9350,N_9381);
nor U9579 (N_9579,N_9337,N_9412);
and U9580 (N_9580,N_9446,N_9413);
and U9581 (N_9581,N_9353,N_9318);
xor U9582 (N_9582,N_9404,N_9366);
nor U9583 (N_9583,N_9418,N_9365);
and U9584 (N_9584,N_9448,N_9310);
or U9585 (N_9585,N_9390,N_9307);
nand U9586 (N_9586,N_9340,N_9375);
nor U9587 (N_9587,N_9406,N_9341);
and U9588 (N_9588,N_9362,N_9380);
or U9589 (N_9589,N_9395,N_9332);
and U9590 (N_9590,N_9306,N_9414);
xor U9591 (N_9591,N_9441,N_9423);
or U9592 (N_9592,N_9300,N_9432);
or U9593 (N_9593,N_9430,N_9444);
nand U9594 (N_9594,N_9432,N_9325);
nand U9595 (N_9595,N_9409,N_9372);
or U9596 (N_9596,N_9314,N_9339);
nand U9597 (N_9597,N_9440,N_9382);
xor U9598 (N_9598,N_9429,N_9446);
or U9599 (N_9599,N_9416,N_9417);
and U9600 (N_9600,N_9536,N_9527);
nand U9601 (N_9601,N_9455,N_9531);
or U9602 (N_9602,N_9483,N_9490);
or U9603 (N_9603,N_9534,N_9506);
and U9604 (N_9604,N_9471,N_9575);
nand U9605 (N_9605,N_9554,N_9552);
or U9606 (N_9606,N_9541,N_9478);
xor U9607 (N_9607,N_9460,N_9526);
or U9608 (N_9608,N_9461,N_9599);
nand U9609 (N_9609,N_9547,N_9588);
xor U9610 (N_9610,N_9535,N_9597);
xnor U9611 (N_9611,N_9537,N_9519);
nand U9612 (N_9612,N_9458,N_9543);
nor U9613 (N_9613,N_9574,N_9453);
nand U9614 (N_9614,N_9589,N_9581);
or U9615 (N_9615,N_9558,N_9544);
or U9616 (N_9616,N_9463,N_9493);
and U9617 (N_9617,N_9533,N_9516);
and U9618 (N_9618,N_9592,N_9521);
xor U9619 (N_9619,N_9591,N_9482);
or U9620 (N_9620,N_9560,N_9467);
nor U9621 (N_9621,N_9494,N_9487);
or U9622 (N_9622,N_9465,N_9515);
and U9623 (N_9623,N_9542,N_9457);
or U9624 (N_9624,N_9479,N_9571);
and U9625 (N_9625,N_9499,N_9504);
and U9626 (N_9626,N_9485,N_9492);
xor U9627 (N_9627,N_9529,N_9476);
or U9628 (N_9628,N_9503,N_9570);
xnor U9629 (N_9629,N_9459,N_9469);
xnor U9630 (N_9630,N_9472,N_9462);
or U9631 (N_9631,N_9518,N_9572);
nor U9632 (N_9632,N_9496,N_9566);
nand U9633 (N_9633,N_9454,N_9450);
xnor U9634 (N_9634,N_9520,N_9556);
nand U9635 (N_9635,N_9584,N_9579);
nor U9636 (N_9636,N_9551,N_9456);
or U9637 (N_9637,N_9538,N_9550);
or U9638 (N_9638,N_9517,N_9546);
nor U9639 (N_9639,N_9470,N_9580);
nand U9640 (N_9640,N_9475,N_9569);
nor U9641 (N_9641,N_9577,N_9545);
nand U9642 (N_9642,N_9498,N_9583);
xor U9643 (N_9643,N_9539,N_9525);
xor U9644 (N_9644,N_9593,N_9488);
and U9645 (N_9645,N_9598,N_9452);
xor U9646 (N_9646,N_9557,N_9530);
or U9647 (N_9647,N_9500,N_9573);
and U9648 (N_9648,N_9524,N_9555);
nor U9649 (N_9649,N_9590,N_9510);
xor U9650 (N_9650,N_9468,N_9489);
and U9651 (N_9651,N_9451,N_9559);
or U9652 (N_9652,N_9564,N_9594);
or U9653 (N_9653,N_9481,N_9511);
or U9654 (N_9654,N_9553,N_9497);
or U9655 (N_9655,N_9568,N_9548);
nand U9656 (N_9656,N_9502,N_9484);
xnor U9657 (N_9657,N_9561,N_9508);
and U9658 (N_9658,N_9464,N_9473);
nand U9659 (N_9659,N_9505,N_9507);
xor U9660 (N_9660,N_9586,N_9513);
nand U9661 (N_9661,N_9514,N_9480);
xor U9662 (N_9662,N_9501,N_9596);
xnor U9663 (N_9663,N_9567,N_9477);
and U9664 (N_9664,N_9491,N_9582);
and U9665 (N_9665,N_9549,N_9540);
xor U9666 (N_9666,N_9466,N_9585);
nand U9667 (N_9667,N_9562,N_9565);
xnor U9668 (N_9668,N_9576,N_9587);
xor U9669 (N_9669,N_9522,N_9495);
or U9670 (N_9670,N_9578,N_9512);
and U9671 (N_9671,N_9595,N_9509);
or U9672 (N_9672,N_9474,N_9563);
nor U9673 (N_9673,N_9528,N_9486);
xnor U9674 (N_9674,N_9523,N_9532);
or U9675 (N_9675,N_9472,N_9523);
xnor U9676 (N_9676,N_9518,N_9507);
xor U9677 (N_9677,N_9555,N_9566);
nand U9678 (N_9678,N_9588,N_9540);
and U9679 (N_9679,N_9536,N_9598);
and U9680 (N_9680,N_9509,N_9513);
or U9681 (N_9681,N_9513,N_9491);
and U9682 (N_9682,N_9562,N_9499);
or U9683 (N_9683,N_9577,N_9569);
or U9684 (N_9684,N_9570,N_9495);
and U9685 (N_9685,N_9559,N_9506);
or U9686 (N_9686,N_9548,N_9571);
xor U9687 (N_9687,N_9492,N_9518);
and U9688 (N_9688,N_9529,N_9561);
xor U9689 (N_9689,N_9587,N_9528);
or U9690 (N_9690,N_9556,N_9554);
nor U9691 (N_9691,N_9510,N_9513);
nor U9692 (N_9692,N_9569,N_9597);
nor U9693 (N_9693,N_9598,N_9563);
or U9694 (N_9694,N_9530,N_9484);
and U9695 (N_9695,N_9538,N_9533);
nor U9696 (N_9696,N_9584,N_9598);
or U9697 (N_9697,N_9534,N_9592);
nand U9698 (N_9698,N_9578,N_9565);
xor U9699 (N_9699,N_9578,N_9496);
nand U9700 (N_9700,N_9595,N_9463);
and U9701 (N_9701,N_9598,N_9560);
or U9702 (N_9702,N_9470,N_9525);
or U9703 (N_9703,N_9470,N_9513);
nor U9704 (N_9704,N_9499,N_9477);
nor U9705 (N_9705,N_9452,N_9555);
nand U9706 (N_9706,N_9494,N_9569);
and U9707 (N_9707,N_9552,N_9456);
or U9708 (N_9708,N_9501,N_9555);
nand U9709 (N_9709,N_9597,N_9566);
or U9710 (N_9710,N_9494,N_9527);
nand U9711 (N_9711,N_9553,N_9588);
or U9712 (N_9712,N_9573,N_9499);
nand U9713 (N_9713,N_9514,N_9456);
and U9714 (N_9714,N_9504,N_9573);
nand U9715 (N_9715,N_9594,N_9501);
nand U9716 (N_9716,N_9511,N_9494);
nand U9717 (N_9717,N_9466,N_9519);
xnor U9718 (N_9718,N_9563,N_9490);
nor U9719 (N_9719,N_9585,N_9574);
or U9720 (N_9720,N_9522,N_9471);
and U9721 (N_9721,N_9453,N_9500);
nor U9722 (N_9722,N_9562,N_9463);
or U9723 (N_9723,N_9568,N_9598);
or U9724 (N_9724,N_9450,N_9554);
or U9725 (N_9725,N_9579,N_9551);
nand U9726 (N_9726,N_9479,N_9460);
xor U9727 (N_9727,N_9489,N_9555);
and U9728 (N_9728,N_9583,N_9460);
nand U9729 (N_9729,N_9529,N_9482);
or U9730 (N_9730,N_9572,N_9593);
nor U9731 (N_9731,N_9537,N_9478);
xnor U9732 (N_9732,N_9551,N_9516);
or U9733 (N_9733,N_9575,N_9590);
nor U9734 (N_9734,N_9562,N_9505);
xor U9735 (N_9735,N_9533,N_9477);
and U9736 (N_9736,N_9595,N_9510);
nand U9737 (N_9737,N_9477,N_9586);
or U9738 (N_9738,N_9529,N_9517);
nand U9739 (N_9739,N_9555,N_9513);
xnor U9740 (N_9740,N_9557,N_9544);
xor U9741 (N_9741,N_9509,N_9555);
xnor U9742 (N_9742,N_9549,N_9528);
or U9743 (N_9743,N_9581,N_9498);
or U9744 (N_9744,N_9475,N_9548);
or U9745 (N_9745,N_9513,N_9536);
nor U9746 (N_9746,N_9520,N_9566);
or U9747 (N_9747,N_9566,N_9503);
nor U9748 (N_9748,N_9538,N_9485);
and U9749 (N_9749,N_9579,N_9482);
nor U9750 (N_9750,N_9720,N_9681);
nand U9751 (N_9751,N_9728,N_9707);
nor U9752 (N_9752,N_9613,N_9708);
or U9753 (N_9753,N_9605,N_9660);
nor U9754 (N_9754,N_9648,N_9730);
and U9755 (N_9755,N_9734,N_9665);
xor U9756 (N_9756,N_9718,N_9619);
nand U9757 (N_9757,N_9692,N_9656);
nand U9758 (N_9758,N_9749,N_9686);
xor U9759 (N_9759,N_9612,N_9735);
nor U9760 (N_9760,N_9661,N_9606);
nor U9761 (N_9761,N_9693,N_9727);
or U9762 (N_9762,N_9699,N_9677);
nand U9763 (N_9763,N_9655,N_9726);
and U9764 (N_9764,N_9622,N_9625);
or U9765 (N_9765,N_9675,N_9670);
nand U9766 (N_9766,N_9706,N_9696);
xnor U9767 (N_9767,N_9682,N_9617);
and U9768 (N_9768,N_9714,N_9673);
and U9769 (N_9769,N_9614,N_9643);
nand U9770 (N_9770,N_9610,N_9657);
nor U9771 (N_9771,N_9701,N_9628);
nand U9772 (N_9772,N_9641,N_9633);
xor U9773 (N_9773,N_9748,N_9674);
or U9774 (N_9774,N_9672,N_9719);
nand U9775 (N_9775,N_9635,N_9663);
and U9776 (N_9776,N_9704,N_9658);
and U9777 (N_9777,N_9639,N_9710);
xor U9778 (N_9778,N_9615,N_9724);
nor U9779 (N_9779,N_9638,N_9601);
and U9780 (N_9780,N_9746,N_9632);
nor U9781 (N_9781,N_9689,N_9671);
xor U9782 (N_9782,N_9680,N_9649);
nor U9783 (N_9783,N_9713,N_9659);
and U9784 (N_9784,N_9740,N_9733);
nor U9785 (N_9785,N_9627,N_9640);
nand U9786 (N_9786,N_9664,N_9703);
and U9787 (N_9787,N_9684,N_9620);
xnor U9788 (N_9788,N_9616,N_9624);
xor U9789 (N_9789,N_9630,N_9744);
and U9790 (N_9790,N_9712,N_9723);
and U9791 (N_9791,N_9603,N_9626);
or U9792 (N_9792,N_9745,N_9647);
xor U9793 (N_9793,N_9687,N_9690);
nor U9794 (N_9794,N_9618,N_9669);
and U9795 (N_9795,N_9721,N_9636);
xor U9796 (N_9796,N_9607,N_9600);
or U9797 (N_9797,N_9651,N_9741);
and U9798 (N_9798,N_9683,N_9743);
xor U9799 (N_9799,N_9739,N_9729);
and U9800 (N_9800,N_9668,N_9700);
nand U9801 (N_9801,N_9725,N_9742);
and U9802 (N_9802,N_9650,N_9715);
nor U9803 (N_9803,N_9705,N_9653);
nand U9804 (N_9804,N_9698,N_9694);
nor U9805 (N_9805,N_9631,N_9688);
xor U9806 (N_9806,N_9695,N_9678);
or U9807 (N_9807,N_9685,N_9602);
nor U9808 (N_9808,N_9709,N_9711);
xor U9809 (N_9809,N_9676,N_9666);
nor U9810 (N_9810,N_9608,N_9634);
nand U9811 (N_9811,N_9621,N_9637);
or U9812 (N_9812,N_9731,N_9629);
xnor U9813 (N_9813,N_9738,N_9604);
nand U9814 (N_9814,N_9702,N_9623);
nand U9815 (N_9815,N_9732,N_9736);
and U9816 (N_9816,N_9667,N_9691);
xnor U9817 (N_9817,N_9697,N_9645);
nand U9818 (N_9818,N_9654,N_9652);
nand U9819 (N_9819,N_9722,N_9747);
nor U9820 (N_9820,N_9737,N_9644);
nor U9821 (N_9821,N_9717,N_9662);
nor U9822 (N_9822,N_9646,N_9679);
xnor U9823 (N_9823,N_9642,N_9609);
nand U9824 (N_9824,N_9716,N_9611);
nor U9825 (N_9825,N_9726,N_9693);
and U9826 (N_9826,N_9738,N_9620);
nand U9827 (N_9827,N_9695,N_9626);
and U9828 (N_9828,N_9693,N_9658);
nor U9829 (N_9829,N_9606,N_9649);
nor U9830 (N_9830,N_9628,N_9679);
or U9831 (N_9831,N_9652,N_9648);
nand U9832 (N_9832,N_9690,N_9672);
nor U9833 (N_9833,N_9738,N_9626);
nand U9834 (N_9834,N_9698,N_9628);
nand U9835 (N_9835,N_9670,N_9715);
nor U9836 (N_9836,N_9670,N_9678);
xnor U9837 (N_9837,N_9746,N_9651);
nand U9838 (N_9838,N_9724,N_9707);
nor U9839 (N_9839,N_9619,N_9722);
and U9840 (N_9840,N_9732,N_9725);
or U9841 (N_9841,N_9669,N_9619);
nand U9842 (N_9842,N_9634,N_9668);
xor U9843 (N_9843,N_9747,N_9734);
or U9844 (N_9844,N_9679,N_9674);
nor U9845 (N_9845,N_9707,N_9695);
nor U9846 (N_9846,N_9652,N_9678);
nor U9847 (N_9847,N_9694,N_9677);
nor U9848 (N_9848,N_9705,N_9695);
nand U9849 (N_9849,N_9719,N_9675);
or U9850 (N_9850,N_9747,N_9656);
or U9851 (N_9851,N_9733,N_9693);
nand U9852 (N_9852,N_9731,N_9688);
or U9853 (N_9853,N_9620,N_9721);
nor U9854 (N_9854,N_9736,N_9636);
xnor U9855 (N_9855,N_9674,N_9737);
nand U9856 (N_9856,N_9648,N_9670);
nor U9857 (N_9857,N_9657,N_9660);
and U9858 (N_9858,N_9658,N_9743);
and U9859 (N_9859,N_9684,N_9714);
and U9860 (N_9860,N_9744,N_9746);
xor U9861 (N_9861,N_9668,N_9685);
nand U9862 (N_9862,N_9625,N_9633);
and U9863 (N_9863,N_9662,N_9659);
xor U9864 (N_9864,N_9665,N_9694);
nand U9865 (N_9865,N_9604,N_9713);
xnor U9866 (N_9866,N_9629,N_9696);
or U9867 (N_9867,N_9613,N_9743);
or U9868 (N_9868,N_9661,N_9633);
nand U9869 (N_9869,N_9702,N_9709);
nor U9870 (N_9870,N_9674,N_9684);
and U9871 (N_9871,N_9689,N_9625);
and U9872 (N_9872,N_9651,N_9633);
xor U9873 (N_9873,N_9640,N_9636);
nor U9874 (N_9874,N_9640,N_9631);
or U9875 (N_9875,N_9737,N_9647);
nand U9876 (N_9876,N_9690,N_9707);
nand U9877 (N_9877,N_9686,N_9728);
or U9878 (N_9878,N_9664,N_9746);
nand U9879 (N_9879,N_9668,N_9747);
and U9880 (N_9880,N_9641,N_9704);
xnor U9881 (N_9881,N_9603,N_9619);
or U9882 (N_9882,N_9604,N_9627);
or U9883 (N_9883,N_9631,N_9742);
xor U9884 (N_9884,N_9692,N_9714);
xor U9885 (N_9885,N_9741,N_9680);
xnor U9886 (N_9886,N_9656,N_9685);
or U9887 (N_9887,N_9629,N_9649);
nand U9888 (N_9888,N_9652,N_9740);
nand U9889 (N_9889,N_9650,N_9688);
xor U9890 (N_9890,N_9645,N_9661);
nand U9891 (N_9891,N_9704,N_9703);
nor U9892 (N_9892,N_9649,N_9662);
xnor U9893 (N_9893,N_9619,N_9663);
xnor U9894 (N_9894,N_9639,N_9641);
nand U9895 (N_9895,N_9649,N_9706);
nor U9896 (N_9896,N_9638,N_9669);
and U9897 (N_9897,N_9624,N_9734);
xor U9898 (N_9898,N_9697,N_9704);
and U9899 (N_9899,N_9639,N_9646);
nor U9900 (N_9900,N_9867,N_9836);
and U9901 (N_9901,N_9835,N_9818);
and U9902 (N_9902,N_9875,N_9784);
or U9903 (N_9903,N_9831,N_9761);
xor U9904 (N_9904,N_9787,N_9883);
or U9905 (N_9905,N_9877,N_9764);
and U9906 (N_9906,N_9821,N_9785);
nor U9907 (N_9907,N_9811,N_9803);
xor U9908 (N_9908,N_9894,N_9862);
and U9909 (N_9909,N_9852,N_9873);
xnor U9910 (N_9910,N_9880,N_9762);
or U9911 (N_9911,N_9804,N_9773);
or U9912 (N_9912,N_9829,N_9828);
nor U9913 (N_9913,N_9795,N_9778);
xor U9914 (N_9914,N_9752,N_9895);
or U9915 (N_9915,N_9899,N_9827);
nor U9916 (N_9916,N_9791,N_9807);
and U9917 (N_9917,N_9792,N_9767);
or U9918 (N_9918,N_9892,N_9871);
xor U9919 (N_9919,N_9859,N_9757);
xor U9920 (N_9920,N_9798,N_9843);
or U9921 (N_9921,N_9812,N_9758);
xnor U9922 (N_9922,N_9885,N_9805);
xnor U9923 (N_9923,N_9822,N_9870);
nor U9924 (N_9924,N_9813,N_9786);
and U9925 (N_9925,N_9806,N_9856);
xor U9926 (N_9926,N_9847,N_9754);
xnor U9927 (N_9927,N_9800,N_9833);
and U9928 (N_9928,N_9797,N_9780);
nand U9929 (N_9929,N_9830,N_9872);
nor U9930 (N_9930,N_9881,N_9775);
and U9931 (N_9931,N_9889,N_9810);
nand U9932 (N_9932,N_9781,N_9816);
and U9933 (N_9933,N_9887,N_9845);
and U9934 (N_9934,N_9890,N_9770);
nor U9935 (N_9935,N_9853,N_9876);
nor U9936 (N_9936,N_9794,N_9865);
or U9937 (N_9937,N_9753,N_9782);
nor U9938 (N_9938,N_9789,N_9861);
and U9939 (N_9939,N_9815,N_9817);
nor U9940 (N_9940,N_9793,N_9855);
or U9941 (N_9941,N_9878,N_9790);
and U9942 (N_9942,N_9799,N_9891);
nor U9943 (N_9943,N_9886,N_9774);
or U9944 (N_9944,N_9846,N_9874);
xnor U9945 (N_9945,N_9824,N_9888);
nand U9946 (N_9946,N_9849,N_9776);
and U9947 (N_9947,N_9819,N_9879);
and U9948 (N_9948,N_9808,N_9834);
and U9949 (N_9949,N_9823,N_9809);
or U9950 (N_9950,N_9788,N_9898);
nor U9951 (N_9951,N_9850,N_9796);
and U9952 (N_9952,N_9783,N_9802);
nand U9953 (N_9953,N_9882,N_9893);
xor U9954 (N_9954,N_9863,N_9751);
and U9955 (N_9955,N_9864,N_9820);
xnor U9956 (N_9956,N_9842,N_9896);
or U9957 (N_9957,N_9765,N_9848);
nand U9958 (N_9958,N_9884,N_9750);
xnor U9959 (N_9959,N_9838,N_9755);
xor U9960 (N_9960,N_9858,N_9779);
and U9961 (N_9961,N_9860,N_9854);
and U9962 (N_9962,N_9825,N_9897);
and U9963 (N_9963,N_9851,N_9772);
nand U9964 (N_9964,N_9826,N_9801);
nor U9965 (N_9965,N_9769,N_9832);
xor U9966 (N_9966,N_9777,N_9844);
or U9967 (N_9967,N_9841,N_9759);
xor U9968 (N_9968,N_9768,N_9766);
xnor U9969 (N_9969,N_9839,N_9840);
xnor U9970 (N_9970,N_9756,N_9763);
nor U9971 (N_9971,N_9814,N_9857);
nand U9972 (N_9972,N_9869,N_9866);
xor U9973 (N_9973,N_9868,N_9837);
and U9974 (N_9974,N_9771,N_9760);
xor U9975 (N_9975,N_9869,N_9783);
xnor U9976 (N_9976,N_9832,N_9793);
and U9977 (N_9977,N_9831,N_9873);
nand U9978 (N_9978,N_9839,N_9780);
or U9979 (N_9979,N_9785,N_9868);
nor U9980 (N_9980,N_9767,N_9770);
or U9981 (N_9981,N_9806,N_9764);
nor U9982 (N_9982,N_9875,N_9816);
nand U9983 (N_9983,N_9772,N_9782);
nor U9984 (N_9984,N_9805,N_9897);
nor U9985 (N_9985,N_9827,N_9829);
xnor U9986 (N_9986,N_9796,N_9802);
nor U9987 (N_9987,N_9859,N_9813);
or U9988 (N_9988,N_9788,N_9759);
nor U9989 (N_9989,N_9841,N_9878);
nor U9990 (N_9990,N_9801,N_9807);
xnor U9991 (N_9991,N_9850,N_9768);
nand U9992 (N_9992,N_9766,N_9811);
and U9993 (N_9993,N_9826,N_9775);
and U9994 (N_9994,N_9788,N_9833);
or U9995 (N_9995,N_9797,N_9890);
and U9996 (N_9996,N_9808,N_9813);
nor U9997 (N_9997,N_9809,N_9894);
or U9998 (N_9998,N_9892,N_9894);
or U9999 (N_9999,N_9760,N_9830);
nand U10000 (N_10000,N_9785,N_9763);
or U10001 (N_10001,N_9769,N_9771);
xnor U10002 (N_10002,N_9780,N_9752);
xor U10003 (N_10003,N_9888,N_9817);
xnor U10004 (N_10004,N_9799,N_9811);
or U10005 (N_10005,N_9888,N_9862);
or U10006 (N_10006,N_9820,N_9808);
xnor U10007 (N_10007,N_9803,N_9864);
xor U10008 (N_10008,N_9787,N_9876);
xnor U10009 (N_10009,N_9878,N_9754);
nand U10010 (N_10010,N_9894,N_9882);
xnor U10011 (N_10011,N_9870,N_9848);
nand U10012 (N_10012,N_9878,N_9787);
nor U10013 (N_10013,N_9896,N_9814);
and U10014 (N_10014,N_9772,N_9806);
and U10015 (N_10015,N_9790,N_9853);
and U10016 (N_10016,N_9847,N_9823);
and U10017 (N_10017,N_9878,N_9753);
nand U10018 (N_10018,N_9770,N_9863);
xnor U10019 (N_10019,N_9814,N_9893);
xor U10020 (N_10020,N_9792,N_9808);
and U10021 (N_10021,N_9870,N_9781);
or U10022 (N_10022,N_9878,N_9891);
and U10023 (N_10023,N_9752,N_9851);
nor U10024 (N_10024,N_9891,N_9866);
and U10025 (N_10025,N_9870,N_9772);
or U10026 (N_10026,N_9857,N_9852);
or U10027 (N_10027,N_9808,N_9880);
nand U10028 (N_10028,N_9864,N_9875);
nor U10029 (N_10029,N_9775,N_9815);
and U10030 (N_10030,N_9849,N_9831);
or U10031 (N_10031,N_9798,N_9831);
xor U10032 (N_10032,N_9828,N_9797);
and U10033 (N_10033,N_9835,N_9780);
and U10034 (N_10034,N_9851,N_9806);
and U10035 (N_10035,N_9833,N_9846);
and U10036 (N_10036,N_9813,N_9846);
or U10037 (N_10037,N_9864,N_9846);
nand U10038 (N_10038,N_9894,N_9863);
nand U10039 (N_10039,N_9840,N_9869);
nand U10040 (N_10040,N_9889,N_9819);
or U10041 (N_10041,N_9815,N_9802);
xor U10042 (N_10042,N_9776,N_9828);
or U10043 (N_10043,N_9777,N_9895);
and U10044 (N_10044,N_9802,N_9812);
or U10045 (N_10045,N_9780,N_9754);
and U10046 (N_10046,N_9878,N_9779);
nand U10047 (N_10047,N_9768,N_9819);
or U10048 (N_10048,N_9758,N_9882);
xnor U10049 (N_10049,N_9871,N_9821);
and U10050 (N_10050,N_9929,N_9909);
and U10051 (N_10051,N_10005,N_9962);
nor U10052 (N_10052,N_10040,N_9906);
nand U10053 (N_10053,N_10039,N_9928);
nor U10054 (N_10054,N_9977,N_9975);
and U10055 (N_10055,N_10025,N_9986);
nand U10056 (N_10056,N_10003,N_9946);
and U10057 (N_10057,N_10015,N_9913);
xor U10058 (N_10058,N_9949,N_9902);
xnor U10059 (N_10059,N_10010,N_9985);
nor U10060 (N_10060,N_9961,N_9979);
nor U10061 (N_10061,N_10021,N_9937);
xnor U10062 (N_10062,N_9934,N_9999);
nand U10063 (N_10063,N_9982,N_9998);
xor U10064 (N_10064,N_9940,N_10024);
nor U10065 (N_10065,N_9989,N_9951);
nor U10066 (N_10066,N_10032,N_10022);
nand U10067 (N_10067,N_9959,N_9996);
nor U10068 (N_10068,N_10047,N_9991);
nor U10069 (N_10069,N_9938,N_9969);
nand U10070 (N_10070,N_9917,N_10016);
nor U10071 (N_10071,N_9974,N_10001);
xnor U10072 (N_10072,N_9958,N_9919);
nor U10073 (N_10073,N_9922,N_9967);
or U10074 (N_10074,N_9904,N_9973);
xnor U10075 (N_10075,N_9954,N_9953);
nand U10076 (N_10076,N_10004,N_10020);
nor U10077 (N_10077,N_10043,N_10041);
nor U10078 (N_10078,N_9988,N_9965);
nand U10079 (N_10079,N_10026,N_9941);
or U10080 (N_10080,N_9950,N_10018);
nor U10081 (N_10081,N_10008,N_10012);
and U10082 (N_10082,N_10035,N_9923);
or U10083 (N_10083,N_9915,N_9921);
nand U10084 (N_10084,N_10029,N_10042);
xnor U10085 (N_10085,N_9920,N_10034);
xor U10086 (N_10086,N_9925,N_9908);
nor U10087 (N_10087,N_9983,N_9935);
nor U10088 (N_10088,N_9980,N_10033);
nand U10089 (N_10089,N_9943,N_10046);
nand U10090 (N_10090,N_9942,N_9994);
nor U10091 (N_10091,N_10017,N_9956);
and U10092 (N_10092,N_10044,N_9903);
and U10093 (N_10093,N_9933,N_10014);
xor U10094 (N_10094,N_10013,N_9981);
or U10095 (N_10095,N_9901,N_10011);
nand U10096 (N_10096,N_9939,N_10049);
xnor U10097 (N_10097,N_9932,N_10031);
and U10098 (N_10098,N_9972,N_9960);
nor U10099 (N_10099,N_9992,N_10030);
xnor U10100 (N_10100,N_9924,N_9952);
nor U10101 (N_10101,N_9945,N_9905);
and U10102 (N_10102,N_10019,N_9993);
nand U10103 (N_10103,N_9936,N_9916);
nor U10104 (N_10104,N_9931,N_10048);
nand U10105 (N_10105,N_9964,N_9971);
nor U10106 (N_10106,N_9970,N_9976);
nand U10107 (N_10107,N_9914,N_10009);
nor U10108 (N_10108,N_9947,N_9987);
or U10109 (N_10109,N_9900,N_9918);
nand U10110 (N_10110,N_9997,N_9990);
or U10111 (N_10111,N_10028,N_9910);
or U10112 (N_10112,N_10002,N_9984);
or U10113 (N_10113,N_9963,N_9944);
and U10114 (N_10114,N_10037,N_10007);
xnor U10115 (N_10115,N_10006,N_10027);
nand U10116 (N_10116,N_9930,N_9968);
or U10117 (N_10117,N_9912,N_10045);
xor U10118 (N_10118,N_10038,N_10036);
and U10119 (N_10119,N_9957,N_9995);
nor U10120 (N_10120,N_9966,N_10000);
and U10121 (N_10121,N_9907,N_9978);
nor U10122 (N_10122,N_9926,N_10023);
xnor U10123 (N_10123,N_9948,N_9927);
xor U10124 (N_10124,N_9911,N_9955);
xor U10125 (N_10125,N_9974,N_9977);
nand U10126 (N_10126,N_10036,N_9934);
nand U10127 (N_10127,N_9954,N_10010);
nand U10128 (N_10128,N_9950,N_9926);
nand U10129 (N_10129,N_10049,N_10029);
or U10130 (N_10130,N_10023,N_9967);
or U10131 (N_10131,N_10049,N_10008);
xor U10132 (N_10132,N_10044,N_9974);
and U10133 (N_10133,N_9905,N_9900);
xor U10134 (N_10134,N_10002,N_9905);
xnor U10135 (N_10135,N_10021,N_9942);
and U10136 (N_10136,N_10010,N_10038);
or U10137 (N_10137,N_9999,N_9964);
nor U10138 (N_10138,N_9961,N_9909);
or U10139 (N_10139,N_9968,N_10005);
or U10140 (N_10140,N_9901,N_9910);
nand U10141 (N_10141,N_9950,N_9904);
or U10142 (N_10142,N_9920,N_9934);
xor U10143 (N_10143,N_10025,N_10028);
nor U10144 (N_10144,N_10004,N_9955);
nor U10145 (N_10145,N_9923,N_10033);
nand U10146 (N_10146,N_9914,N_9900);
and U10147 (N_10147,N_10047,N_9902);
or U10148 (N_10148,N_9926,N_9982);
nand U10149 (N_10149,N_10012,N_10040);
or U10150 (N_10150,N_9950,N_9938);
or U10151 (N_10151,N_9930,N_9912);
and U10152 (N_10152,N_10042,N_10000);
nor U10153 (N_10153,N_9938,N_9904);
nand U10154 (N_10154,N_10026,N_9995);
or U10155 (N_10155,N_9977,N_9910);
nor U10156 (N_10156,N_9956,N_10026);
nand U10157 (N_10157,N_9961,N_9935);
xor U10158 (N_10158,N_9962,N_9933);
nand U10159 (N_10159,N_9918,N_9928);
or U10160 (N_10160,N_9919,N_9915);
nand U10161 (N_10161,N_10032,N_9973);
nor U10162 (N_10162,N_10030,N_10018);
nand U10163 (N_10163,N_10035,N_9947);
nand U10164 (N_10164,N_10000,N_9967);
xnor U10165 (N_10165,N_9907,N_10011);
or U10166 (N_10166,N_9966,N_9903);
nor U10167 (N_10167,N_10010,N_9929);
and U10168 (N_10168,N_9915,N_9950);
or U10169 (N_10169,N_9970,N_9925);
and U10170 (N_10170,N_10042,N_9933);
nand U10171 (N_10171,N_10027,N_9929);
or U10172 (N_10172,N_9998,N_9943);
and U10173 (N_10173,N_10039,N_9971);
xnor U10174 (N_10174,N_10012,N_10037);
or U10175 (N_10175,N_9976,N_10026);
xor U10176 (N_10176,N_9920,N_10037);
nor U10177 (N_10177,N_9995,N_9984);
nor U10178 (N_10178,N_9977,N_9946);
or U10179 (N_10179,N_10006,N_10028);
xor U10180 (N_10180,N_10024,N_10006);
and U10181 (N_10181,N_9929,N_9907);
or U10182 (N_10182,N_10040,N_9974);
or U10183 (N_10183,N_9991,N_9934);
nand U10184 (N_10184,N_9905,N_9970);
or U10185 (N_10185,N_9989,N_9911);
nor U10186 (N_10186,N_9960,N_9918);
and U10187 (N_10187,N_10047,N_9931);
or U10188 (N_10188,N_9927,N_9975);
or U10189 (N_10189,N_9920,N_9941);
and U10190 (N_10190,N_9994,N_9903);
or U10191 (N_10191,N_9963,N_9912);
and U10192 (N_10192,N_9926,N_9987);
or U10193 (N_10193,N_9956,N_9941);
xor U10194 (N_10194,N_10015,N_9943);
nand U10195 (N_10195,N_9929,N_9971);
nand U10196 (N_10196,N_10037,N_9982);
nor U10197 (N_10197,N_9901,N_9937);
nor U10198 (N_10198,N_9960,N_9944);
xnor U10199 (N_10199,N_10040,N_9926);
and U10200 (N_10200,N_10154,N_10172);
xnor U10201 (N_10201,N_10087,N_10059);
xnor U10202 (N_10202,N_10062,N_10177);
or U10203 (N_10203,N_10152,N_10099);
and U10204 (N_10204,N_10178,N_10193);
and U10205 (N_10205,N_10066,N_10072);
or U10206 (N_10206,N_10084,N_10142);
and U10207 (N_10207,N_10167,N_10131);
nand U10208 (N_10208,N_10116,N_10093);
and U10209 (N_10209,N_10160,N_10094);
and U10210 (N_10210,N_10100,N_10188);
and U10211 (N_10211,N_10095,N_10122);
xor U10212 (N_10212,N_10067,N_10135);
nor U10213 (N_10213,N_10077,N_10191);
and U10214 (N_10214,N_10189,N_10120);
or U10215 (N_10215,N_10165,N_10136);
and U10216 (N_10216,N_10151,N_10103);
nor U10217 (N_10217,N_10169,N_10159);
xor U10218 (N_10218,N_10065,N_10185);
nor U10219 (N_10219,N_10076,N_10056);
xor U10220 (N_10220,N_10164,N_10088);
xnor U10221 (N_10221,N_10158,N_10146);
or U10222 (N_10222,N_10055,N_10109);
xor U10223 (N_10223,N_10186,N_10199);
or U10224 (N_10224,N_10166,N_10081);
or U10225 (N_10225,N_10075,N_10192);
xor U10226 (N_10226,N_10061,N_10114);
nor U10227 (N_10227,N_10145,N_10183);
or U10228 (N_10228,N_10098,N_10053);
or U10229 (N_10229,N_10130,N_10123);
and U10230 (N_10230,N_10163,N_10126);
or U10231 (N_10231,N_10108,N_10182);
nand U10232 (N_10232,N_10073,N_10079);
nand U10233 (N_10233,N_10090,N_10082);
xor U10234 (N_10234,N_10176,N_10070);
or U10235 (N_10235,N_10052,N_10110);
xor U10236 (N_10236,N_10128,N_10155);
xnor U10237 (N_10237,N_10132,N_10113);
and U10238 (N_10238,N_10057,N_10068);
and U10239 (N_10239,N_10144,N_10156);
and U10240 (N_10240,N_10063,N_10137);
nand U10241 (N_10241,N_10089,N_10117);
xor U10242 (N_10242,N_10175,N_10104);
nor U10243 (N_10243,N_10180,N_10187);
or U10244 (N_10244,N_10161,N_10138);
or U10245 (N_10245,N_10085,N_10106);
xor U10246 (N_10246,N_10080,N_10190);
xnor U10247 (N_10247,N_10092,N_10194);
and U10248 (N_10248,N_10170,N_10091);
or U10249 (N_10249,N_10071,N_10139);
or U10250 (N_10250,N_10197,N_10125);
xor U10251 (N_10251,N_10101,N_10069);
xor U10252 (N_10252,N_10162,N_10195);
or U10253 (N_10253,N_10112,N_10150);
nor U10254 (N_10254,N_10105,N_10153);
nor U10255 (N_10255,N_10141,N_10058);
xor U10256 (N_10256,N_10086,N_10078);
xnor U10257 (N_10257,N_10051,N_10184);
and U10258 (N_10258,N_10064,N_10097);
nand U10259 (N_10259,N_10198,N_10168);
nor U10260 (N_10260,N_10181,N_10134);
and U10261 (N_10261,N_10157,N_10118);
xor U10262 (N_10262,N_10129,N_10115);
xor U10263 (N_10263,N_10127,N_10119);
nand U10264 (N_10264,N_10147,N_10196);
nand U10265 (N_10265,N_10140,N_10050);
nand U10266 (N_10266,N_10179,N_10149);
and U10267 (N_10267,N_10124,N_10174);
xor U10268 (N_10268,N_10102,N_10121);
or U10269 (N_10269,N_10143,N_10054);
xor U10270 (N_10270,N_10148,N_10171);
and U10271 (N_10271,N_10173,N_10133);
nand U10272 (N_10272,N_10111,N_10107);
nor U10273 (N_10273,N_10074,N_10060);
xnor U10274 (N_10274,N_10083,N_10096);
or U10275 (N_10275,N_10140,N_10104);
or U10276 (N_10276,N_10199,N_10135);
or U10277 (N_10277,N_10060,N_10055);
nand U10278 (N_10278,N_10091,N_10183);
or U10279 (N_10279,N_10103,N_10114);
and U10280 (N_10280,N_10125,N_10073);
and U10281 (N_10281,N_10162,N_10129);
nand U10282 (N_10282,N_10089,N_10057);
and U10283 (N_10283,N_10197,N_10103);
or U10284 (N_10284,N_10080,N_10125);
nand U10285 (N_10285,N_10061,N_10147);
nor U10286 (N_10286,N_10093,N_10076);
and U10287 (N_10287,N_10104,N_10090);
and U10288 (N_10288,N_10163,N_10188);
nand U10289 (N_10289,N_10094,N_10087);
nor U10290 (N_10290,N_10059,N_10074);
nand U10291 (N_10291,N_10085,N_10188);
and U10292 (N_10292,N_10072,N_10096);
nor U10293 (N_10293,N_10181,N_10120);
nor U10294 (N_10294,N_10161,N_10196);
xor U10295 (N_10295,N_10077,N_10114);
and U10296 (N_10296,N_10198,N_10130);
xor U10297 (N_10297,N_10163,N_10111);
nor U10298 (N_10298,N_10183,N_10178);
nand U10299 (N_10299,N_10062,N_10078);
nand U10300 (N_10300,N_10172,N_10051);
nand U10301 (N_10301,N_10157,N_10129);
or U10302 (N_10302,N_10199,N_10189);
and U10303 (N_10303,N_10144,N_10163);
nand U10304 (N_10304,N_10056,N_10084);
nor U10305 (N_10305,N_10077,N_10134);
xor U10306 (N_10306,N_10184,N_10062);
xnor U10307 (N_10307,N_10095,N_10175);
xnor U10308 (N_10308,N_10156,N_10160);
nand U10309 (N_10309,N_10165,N_10118);
or U10310 (N_10310,N_10161,N_10128);
nor U10311 (N_10311,N_10153,N_10081);
nor U10312 (N_10312,N_10149,N_10101);
or U10313 (N_10313,N_10100,N_10165);
or U10314 (N_10314,N_10120,N_10145);
or U10315 (N_10315,N_10152,N_10081);
xnor U10316 (N_10316,N_10168,N_10084);
nand U10317 (N_10317,N_10110,N_10100);
nand U10318 (N_10318,N_10081,N_10053);
or U10319 (N_10319,N_10181,N_10115);
and U10320 (N_10320,N_10068,N_10181);
nor U10321 (N_10321,N_10157,N_10187);
nand U10322 (N_10322,N_10171,N_10189);
or U10323 (N_10323,N_10192,N_10157);
nor U10324 (N_10324,N_10139,N_10122);
nand U10325 (N_10325,N_10137,N_10160);
xor U10326 (N_10326,N_10126,N_10093);
nor U10327 (N_10327,N_10104,N_10153);
xor U10328 (N_10328,N_10088,N_10171);
and U10329 (N_10329,N_10191,N_10090);
or U10330 (N_10330,N_10129,N_10070);
or U10331 (N_10331,N_10091,N_10134);
nor U10332 (N_10332,N_10159,N_10067);
or U10333 (N_10333,N_10148,N_10098);
nor U10334 (N_10334,N_10122,N_10089);
xnor U10335 (N_10335,N_10113,N_10052);
nand U10336 (N_10336,N_10193,N_10121);
nand U10337 (N_10337,N_10158,N_10098);
and U10338 (N_10338,N_10096,N_10076);
nand U10339 (N_10339,N_10109,N_10076);
and U10340 (N_10340,N_10056,N_10081);
xor U10341 (N_10341,N_10103,N_10094);
xor U10342 (N_10342,N_10121,N_10052);
nor U10343 (N_10343,N_10065,N_10129);
or U10344 (N_10344,N_10084,N_10153);
xnor U10345 (N_10345,N_10090,N_10098);
nor U10346 (N_10346,N_10062,N_10089);
and U10347 (N_10347,N_10170,N_10126);
xor U10348 (N_10348,N_10092,N_10143);
nand U10349 (N_10349,N_10148,N_10118);
nor U10350 (N_10350,N_10263,N_10318);
or U10351 (N_10351,N_10203,N_10234);
or U10352 (N_10352,N_10249,N_10317);
or U10353 (N_10353,N_10331,N_10233);
or U10354 (N_10354,N_10316,N_10258);
and U10355 (N_10355,N_10228,N_10298);
and U10356 (N_10356,N_10325,N_10240);
and U10357 (N_10357,N_10227,N_10342);
nor U10358 (N_10358,N_10256,N_10200);
xor U10359 (N_10359,N_10276,N_10322);
nand U10360 (N_10360,N_10344,N_10265);
xnor U10361 (N_10361,N_10210,N_10204);
nand U10362 (N_10362,N_10205,N_10246);
or U10363 (N_10363,N_10224,N_10267);
xnor U10364 (N_10364,N_10297,N_10217);
or U10365 (N_10365,N_10313,N_10226);
and U10366 (N_10366,N_10283,N_10348);
nand U10367 (N_10367,N_10274,N_10266);
xor U10368 (N_10368,N_10334,N_10216);
or U10369 (N_10369,N_10248,N_10264);
nand U10370 (N_10370,N_10251,N_10326);
xnor U10371 (N_10371,N_10245,N_10333);
xor U10372 (N_10372,N_10229,N_10314);
nand U10373 (N_10373,N_10338,N_10304);
nor U10374 (N_10374,N_10312,N_10328);
nand U10375 (N_10375,N_10315,N_10296);
and U10376 (N_10376,N_10242,N_10201);
and U10377 (N_10377,N_10280,N_10332);
nor U10378 (N_10378,N_10213,N_10250);
nand U10379 (N_10379,N_10273,N_10335);
and U10380 (N_10380,N_10215,N_10239);
nor U10381 (N_10381,N_10287,N_10269);
and U10382 (N_10382,N_10236,N_10295);
and U10383 (N_10383,N_10285,N_10202);
and U10384 (N_10384,N_10341,N_10214);
nand U10385 (N_10385,N_10320,N_10294);
or U10386 (N_10386,N_10271,N_10241);
nand U10387 (N_10387,N_10225,N_10219);
nor U10388 (N_10388,N_10207,N_10279);
or U10389 (N_10389,N_10293,N_10339);
nor U10390 (N_10390,N_10221,N_10222);
nand U10391 (N_10391,N_10288,N_10218);
nand U10392 (N_10392,N_10347,N_10232);
and U10393 (N_10393,N_10327,N_10300);
xnor U10394 (N_10394,N_10211,N_10291);
and U10395 (N_10395,N_10286,N_10329);
xor U10396 (N_10396,N_10336,N_10257);
nand U10397 (N_10397,N_10301,N_10244);
and U10398 (N_10398,N_10206,N_10261);
and U10399 (N_10399,N_10337,N_10282);
and U10400 (N_10400,N_10305,N_10275);
nand U10401 (N_10401,N_10323,N_10309);
nor U10402 (N_10402,N_10284,N_10237);
nor U10403 (N_10403,N_10290,N_10330);
nor U10404 (N_10404,N_10262,N_10278);
or U10405 (N_10405,N_10308,N_10306);
or U10406 (N_10406,N_10303,N_10349);
and U10407 (N_10407,N_10259,N_10307);
xnor U10408 (N_10408,N_10260,N_10340);
xor U10409 (N_10409,N_10343,N_10252);
nand U10410 (N_10410,N_10254,N_10220);
or U10411 (N_10411,N_10243,N_10310);
nand U10412 (N_10412,N_10345,N_10289);
nor U10413 (N_10413,N_10321,N_10253);
and U10414 (N_10414,N_10346,N_10277);
xnor U10415 (N_10415,N_10268,N_10231);
and U10416 (N_10416,N_10209,N_10302);
nor U10417 (N_10417,N_10311,N_10270);
or U10418 (N_10418,N_10247,N_10238);
or U10419 (N_10419,N_10235,N_10208);
nor U10420 (N_10420,N_10255,N_10292);
or U10421 (N_10421,N_10272,N_10281);
nor U10422 (N_10422,N_10324,N_10223);
or U10423 (N_10423,N_10299,N_10212);
or U10424 (N_10424,N_10230,N_10319);
nor U10425 (N_10425,N_10282,N_10313);
or U10426 (N_10426,N_10208,N_10233);
xnor U10427 (N_10427,N_10274,N_10321);
nand U10428 (N_10428,N_10318,N_10301);
or U10429 (N_10429,N_10218,N_10296);
nor U10430 (N_10430,N_10233,N_10340);
and U10431 (N_10431,N_10243,N_10290);
or U10432 (N_10432,N_10278,N_10219);
and U10433 (N_10433,N_10255,N_10294);
and U10434 (N_10434,N_10345,N_10330);
xor U10435 (N_10435,N_10332,N_10325);
and U10436 (N_10436,N_10255,N_10200);
xnor U10437 (N_10437,N_10284,N_10348);
nor U10438 (N_10438,N_10245,N_10272);
and U10439 (N_10439,N_10262,N_10312);
nor U10440 (N_10440,N_10304,N_10229);
nor U10441 (N_10441,N_10227,N_10229);
nor U10442 (N_10442,N_10209,N_10327);
and U10443 (N_10443,N_10215,N_10236);
and U10444 (N_10444,N_10317,N_10274);
xor U10445 (N_10445,N_10233,N_10271);
xnor U10446 (N_10446,N_10219,N_10321);
nor U10447 (N_10447,N_10298,N_10237);
and U10448 (N_10448,N_10321,N_10250);
and U10449 (N_10449,N_10229,N_10221);
nor U10450 (N_10450,N_10205,N_10347);
nor U10451 (N_10451,N_10246,N_10322);
xnor U10452 (N_10452,N_10244,N_10212);
xor U10453 (N_10453,N_10224,N_10296);
and U10454 (N_10454,N_10229,N_10214);
or U10455 (N_10455,N_10223,N_10308);
and U10456 (N_10456,N_10247,N_10315);
nand U10457 (N_10457,N_10280,N_10294);
nand U10458 (N_10458,N_10270,N_10203);
nor U10459 (N_10459,N_10262,N_10344);
xnor U10460 (N_10460,N_10340,N_10222);
and U10461 (N_10461,N_10292,N_10337);
nand U10462 (N_10462,N_10214,N_10239);
nand U10463 (N_10463,N_10313,N_10210);
xnor U10464 (N_10464,N_10332,N_10341);
nor U10465 (N_10465,N_10330,N_10225);
nand U10466 (N_10466,N_10320,N_10240);
xnor U10467 (N_10467,N_10203,N_10222);
nand U10468 (N_10468,N_10318,N_10222);
xnor U10469 (N_10469,N_10324,N_10319);
xnor U10470 (N_10470,N_10245,N_10213);
and U10471 (N_10471,N_10269,N_10273);
xnor U10472 (N_10472,N_10348,N_10312);
nand U10473 (N_10473,N_10317,N_10296);
or U10474 (N_10474,N_10312,N_10258);
nor U10475 (N_10475,N_10347,N_10258);
and U10476 (N_10476,N_10324,N_10216);
and U10477 (N_10477,N_10336,N_10263);
nand U10478 (N_10478,N_10214,N_10212);
xnor U10479 (N_10479,N_10327,N_10339);
nor U10480 (N_10480,N_10326,N_10296);
and U10481 (N_10481,N_10299,N_10236);
nor U10482 (N_10482,N_10329,N_10209);
nor U10483 (N_10483,N_10325,N_10300);
nand U10484 (N_10484,N_10284,N_10279);
and U10485 (N_10485,N_10286,N_10230);
nor U10486 (N_10486,N_10213,N_10305);
nand U10487 (N_10487,N_10249,N_10251);
nor U10488 (N_10488,N_10241,N_10279);
xor U10489 (N_10489,N_10227,N_10344);
nand U10490 (N_10490,N_10279,N_10324);
and U10491 (N_10491,N_10247,N_10221);
and U10492 (N_10492,N_10264,N_10327);
nor U10493 (N_10493,N_10283,N_10257);
nand U10494 (N_10494,N_10294,N_10293);
and U10495 (N_10495,N_10223,N_10249);
nand U10496 (N_10496,N_10279,N_10283);
and U10497 (N_10497,N_10227,N_10207);
nor U10498 (N_10498,N_10263,N_10274);
and U10499 (N_10499,N_10332,N_10216);
and U10500 (N_10500,N_10425,N_10499);
and U10501 (N_10501,N_10431,N_10381);
xnor U10502 (N_10502,N_10351,N_10495);
nand U10503 (N_10503,N_10372,N_10396);
or U10504 (N_10504,N_10398,N_10446);
nand U10505 (N_10505,N_10494,N_10453);
xnor U10506 (N_10506,N_10395,N_10358);
nand U10507 (N_10507,N_10374,N_10422);
xor U10508 (N_10508,N_10365,N_10362);
xnor U10509 (N_10509,N_10355,N_10463);
xnor U10510 (N_10510,N_10437,N_10384);
xor U10511 (N_10511,N_10410,N_10389);
nand U10512 (N_10512,N_10475,N_10392);
xnor U10513 (N_10513,N_10370,N_10443);
and U10514 (N_10514,N_10361,N_10429);
nor U10515 (N_10515,N_10373,N_10383);
or U10516 (N_10516,N_10407,N_10455);
nand U10517 (N_10517,N_10460,N_10428);
nand U10518 (N_10518,N_10382,N_10408);
and U10519 (N_10519,N_10484,N_10445);
or U10520 (N_10520,N_10457,N_10473);
and U10521 (N_10521,N_10421,N_10447);
nand U10522 (N_10522,N_10405,N_10385);
xnor U10523 (N_10523,N_10424,N_10356);
nor U10524 (N_10524,N_10458,N_10353);
xor U10525 (N_10525,N_10386,N_10417);
xor U10526 (N_10526,N_10468,N_10465);
nor U10527 (N_10527,N_10413,N_10488);
and U10528 (N_10528,N_10450,N_10489);
nor U10529 (N_10529,N_10497,N_10472);
or U10530 (N_10530,N_10487,N_10426);
and U10531 (N_10531,N_10491,N_10403);
or U10532 (N_10532,N_10394,N_10482);
nor U10533 (N_10533,N_10368,N_10485);
nor U10534 (N_10534,N_10415,N_10496);
xnor U10535 (N_10535,N_10363,N_10404);
nand U10536 (N_10536,N_10430,N_10483);
and U10537 (N_10537,N_10439,N_10493);
xnor U10538 (N_10538,N_10451,N_10391);
nor U10539 (N_10539,N_10448,N_10399);
or U10540 (N_10540,N_10388,N_10436);
nor U10541 (N_10541,N_10401,N_10478);
nand U10542 (N_10542,N_10357,N_10377);
and U10543 (N_10543,N_10481,N_10402);
nor U10544 (N_10544,N_10406,N_10474);
nand U10545 (N_10545,N_10486,N_10380);
or U10546 (N_10546,N_10416,N_10452);
nor U10547 (N_10547,N_10441,N_10498);
or U10548 (N_10548,N_10379,N_10459);
nand U10549 (N_10549,N_10418,N_10419);
nand U10550 (N_10550,N_10354,N_10467);
nand U10551 (N_10551,N_10440,N_10471);
nor U10552 (N_10552,N_10420,N_10393);
nor U10553 (N_10553,N_10490,N_10378);
and U10554 (N_10554,N_10369,N_10466);
nor U10555 (N_10555,N_10360,N_10449);
nor U10556 (N_10556,N_10438,N_10412);
xnor U10557 (N_10557,N_10414,N_10397);
or U10558 (N_10558,N_10442,N_10434);
and U10559 (N_10559,N_10350,N_10435);
or U10560 (N_10560,N_10409,N_10444);
xnor U10561 (N_10561,N_10432,N_10411);
nor U10562 (N_10562,N_10462,N_10364);
nor U10563 (N_10563,N_10479,N_10376);
nor U10564 (N_10564,N_10366,N_10375);
nor U10565 (N_10565,N_10464,N_10387);
or U10566 (N_10566,N_10480,N_10371);
and U10567 (N_10567,N_10427,N_10492);
nand U10568 (N_10568,N_10454,N_10367);
or U10569 (N_10569,N_10476,N_10359);
nor U10570 (N_10570,N_10352,N_10390);
xor U10571 (N_10571,N_10477,N_10400);
xnor U10572 (N_10572,N_10456,N_10469);
xor U10573 (N_10573,N_10461,N_10470);
or U10574 (N_10574,N_10433,N_10423);
nor U10575 (N_10575,N_10365,N_10442);
and U10576 (N_10576,N_10409,N_10485);
or U10577 (N_10577,N_10444,N_10480);
nor U10578 (N_10578,N_10360,N_10375);
and U10579 (N_10579,N_10451,N_10381);
and U10580 (N_10580,N_10380,N_10419);
and U10581 (N_10581,N_10412,N_10354);
nand U10582 (N_10582,N_10496,N_10373);
nor U10583 (N_10583,N_10382,N_10475);
xor U10584 (N_10584,N_10435,N_10498);
nand U10585 (N_10585,N_10496,N_10443);
or U10586 (N_10586,N_10395,N_10354);
xnor U10587 (N_10587,N_10359,N_10404);
nand U10588 (N_10588,N_10470,N_10494);
and U10589 (N_10589,N_10397,N_10379);
nand U10590 (N_10590,N_10385,N_10442);
and U10591 (N_10591,N_10365,N_10436);
and U10592 (N_10592,N_10431,N_10388);
nor U10593 (N_10593,N_10499,N_10355);
nor U10594 (N_10594,N_10492,N_10436);
or U10595 (N_10595,N_10378,N_10417);
nor U10596 (N_10596,N_10470,N_10388);
xnor U10597 (N_10597,N_10398,N_10384);
or U10598 (N_10598,N_10468,N_10393);
xor U10599 (N_10599,N_10451,N_10492);
nor U10600 (N_10600,N_10431,N_10402);
xnor U10601 (N_10601,N_10397,N_10410);
nand U10602 (N_10602,N_10465,N_10477);
xnor U10603 (N_10603,N_10377,N_10407);
nor U10604 (N_10604,N_10403,N_10486);
xor U10605 (N_10605,N_10362,N_10419);
xnor U10606 (N_10606,N_10486,N_10396);
nand U10607 (N_10607,N_10398,N_10406);
nand U10608 (N_10608,N_10425,N_10377);
and U10609 (N_10609,N_10455,N_10491);
or U10610 (N_10610,N_10472,N_10485);
nand U10611 (N_10611,N_10370,N_10487);
and U10612 (N_10612,N_10450,N_10490);
xnor U10613 (N_10613,N_10453,N_10499);
or U10614 (N_10614,N_10489,N_10460);
and U10615 (N_10615,N_10421,N_10406);
and U10616 (N_10616,N_10485,N_10498);
nand U10617 (N_10617,N_10417,N_10363);
xnor U10618 (N_10618,N_10465,N_10429);
xor U10619 (N_10619,N_10468,N_10417);
nor U10620 (N_10620,N_10487,N_10480);
nand U10621 (N_10621,N_10398,N_10393);
or U10622 (N_10622,N_10431,N_10499);
and U10623 (N_10623,N_10432,N_10496);
nand U10624 (N_10624,N_10380,N_10499);
or U10625 (N_10625,N_10481,N_10431);
xor U10626 (N_10626,N_10425,N_10423);
nand U10627 (N_10627,N_10387,N_10363);
xnor U10628 (N_10628,N_10409,N_10427);
and U10629 (N_10629,N_10462,N_10358);
nand U10630 (N_10630,N_10384,N_10365);
nand U10631 (N_10631,N_10488,N_10396);
nor U10632 (N_10632,N_10476,N_10369);
nand U10633 (N_10633,N_10463,N_10365);
or U10634 (N_10634,N_10413,N_10444);
and U10635 (N_10635,N_10493,N_10364);
xnor U10636 (N_10636,N_10497,N_10483);
xor U10637 (N_10637,N_10456,N_10373);
nor U10638 (N_10638,N_10351,N_10426);
and U10639 (N_10639,N_10351,N_10485);
xnor U10640 (N_10640,N_10451,N_10423);
nand U10641 (N_10641,N_10410,N_10398);
or U10642 (N_10642,N_10443,N_10499);
nand U10643 (N_10643,N_10370,N_10458);
and U10644 (N_10644,N_10424,N_10362);
or U10645 (N_10645,N_10480,N_10409);
nand U10646 (N_10646,N_10451,N_10416);
xor U10647 (N_10647,N_10405,N_10456);
nand U10648 (N_10648,N_10467,N_10481);
and U10649 (N_10649,N_10418,N_10464);
and U10650 (N_10650,N_10592,N_10625);
xor U10651 (N_10651,N_10584,N_10538);
and U10652 (N_10652,N_10640,N_10645);
and U10653 (N_10653,N_10517,N_10596);
xor U10654 (N_10654,N_10589,N_10563);
nand U10655 (N_10655,N_10603,N_10544);
xor U10656 (N_10656,N_10530,N_10593);
nand U10657 (N_10657,N_10630,N_10522);
and U10658 (N_10658,N_10548,N_10638);
and U10659 (N_10659,N_10604,N_10559);
nor U10660 (N_10660,N_10643,N_10610);
or U10661 (N_10661,N_10537,N_10510);
nor U10662 (N_10662,N_10597,N_10631);
nand U10663 (N_10663,N_10626,N_10527);
nand U10664 (N_10664,N_10639,N_10535);
nand U10665 (N_10665,N_10627,N_10533);
and U10666 (N_10666,N_10561,N_10591);
or U10667 (N_10667,N_10579,N_10542);
xnor U10668 (N_10668,N_10632,N_10614);
nor U10669 (N_10669,N_10621,N_10573);
nor U10670 (N_10670,N_10512,N_10556);
nand U10671 (N_10671,N_10607,N_10601);
xnor U10672 (N_10672,N_10511,N_10580);
and U10673 (N_10673,N_10606,N_10577);
and U10674 (N_10674,N_10618,N_10641);
and U10675 (N_10675,N_10555,N_10622);
xor U10676 (N_10676,N_10531,N_10629);
or U10677 (N_10677,N_10569,N_10609);
or U10678 (N_10678,N_10628,N_10600);
nor U10679 (N_10679,N_10649,N_10545);
nor U10680 (N_10680,N_10586,N_10567);
and U10681 (N_10681,N_10566,N_10541);
nor U10682 (N_10682,N_10565,N_10612);
nand U10683 (N_10683,N_10501,N_10594);
xor U10684 (N_10684,N_10602,N_10608);
xor U10685 (N_10685,N_10648,N_10528);
nand U10686 (N_10686,N_10587,N_10515);
nor U10687 (N_10687,N_10585,N_10553);
xnor U10688 (N_10688,N_10646,N_10503);
nand U10689 (N_10689,N_10543,N_10578);
or U10690 (N_10690,N_10647,N_10642);
nand U10691 (N_10691,N_10634,N_10611);
and U10692 (N_10692,N_10613,N_10571);
xor U10693 (N_10693,N_10526,N_10507);
or U10694 (N_10694,N_10505,N_10637);
and U10695 (N_10695,N_10644,N_10633);
nand U10696 (N_10696,N_10552,N_10557);
nor U10697 (N_10697,N_10506,N_10536);
nor U10698 (N_10698,N_10595,N_10525);
and U10699 (N_10699,N_10581,N_10636);
and U10700 (N_10700,N_10624,N_10620);
nor U10701 (N_10701,N_10598,N_10588);
nand U10702 (N_10702,N_10514,N_10560);
xnor U10703 (N_10703,N_10532,N_10616);
and U10704 (N_10704,N_10583,N_10549);
xnor U10705 (N_10705,N_10617,N_10570);
or U10706 (N_10706,N_10500,N_10572);
and U10707 (N_10707,N_10562,N_10623);
nand U10708 (N_10708,N_10529,N_10564);
nand U10709 (N_10709,N_10574,N_10550);
or U10710 (N_10710,N_10590,N_10582);
nand U10711 (N_10711,N_10523,N_10502);
xor U10712 (N_10712,N_10509,N_10504);
or U10713 (N_10713,N_10534,N_10576);
and U10714 (N_10714,N_10508,N_10635);
and U10715 (N_10715,N_10524,N_10539);
nor U10716 (N_10716,N_10568,N_10619);
and U10717 (N_10717,N_10516,N_10558);
nor U10718 (N_10718,N_10605,N_10513);
or U10719 (N_10719,N_10521,N_10575);
xor U10720 (N_10720,N_10520,N_10546);
and U10721 (N_10721,N_10554,N_10551);
or U10722 (N_10722,N_10599,N_10519);
nand U10723 (N_10723,N_10518,N_10615);
nand U10724 (N_10724,N_10540,N_10547);
and U10725 (N_10725,N_10624,N_10607);
and U10726 (N_10726,N_10581,N_10614);
nor U10727 (N_10727,N_10577,N_10514);
nor U10728 (N_10728,N_10524,N_10505);
xnor U10729 (N_10729,N_10519,N_10627);
nor U10730 (N_10730,N_10611,N_10539);
or U10731 (N_10731,N_10500,N_10611);
nand U10732 (N_10732,N_10512,N_10572);
xnor U10733 (N_10733,N_10607,N_10537);
nand U10734 (N_10734,N_10615,N_10609);
xor U10735 (N_10735,N_10525,N_10540);
nand U10736 (N_10736,N_10594,N_10608);
and U10737 (N_10737,N_10534,N_10556);
xor U10738 (N_10738,N_10621,N_10602);
nand U10739 (N_10739,N_10515,N_10579);
or U10740 (N_10740,N_10559,N_10574);
xnor U10741 (N_10741,N_10594,N_10514);
nor U10742 (N_10742,N_10588,N_10640);
nand U10743 (N_10743,N_10546,N_10625);
nor U10744 (N_10744,N_10568,N_10572);
xnor U10745 (N_10745,N_10556,N_10510);
xnor U10746 (N_10746,N_10518,N_10621);
xor U10747 (N_10747,N_10624,N_10533);
and U10748 (N_10748,N_10648,N_10631);
nand U10749 (N_10749,N_10627,N_10534);
nor U10750 (N_10750,N_10647,N_10574);
xor U10751 (N_10751,N_10523,N_10526);
xor U10752 (N_10752,N_10551,N_10529);
xnor U10753 (N_10753,N_10631,N_10530);
nand U10754 (N_10754,N_10508,N_10619);
nor U10755 (N_10755,N_10647,N_10558);
xor U10756 (N_10756,N_10647,N_10551);
or U10757 (N_10757,N_10595,N_10611);
nand U10758 (N_10758,N_10508,N_10626);
or U10759 (N_10759,N_10503,N_10556);
and U10760 (N_10760,N_10579,N_10607);
nor U10761 (N_10761,N_10605,N_10600);
nand U10762 (N_10762,N_10589,N_10521);
xor U10763 (N_10763,N_10549,N_10615);
xor U10764 (N_10764,N_10582,N_10533);
and U10765 (N_10765,N_10533,N_10583);
xor U10766 (N_10766,N_10628,N_10644);
and U10767 (N_10767,N_10616,N_10639);
and U10768 (N_10768,N_10560,N_10509);
and U10769 (N_10769,N_10639,N_10603);
nor U10770 (N_10770,N_10503,N_10527);
xor U10771 (N_10771,N_10647,N_10562);
xnor U10772 (N_10772,N_10522,N_10617);
xnor U10773 (N_10773,N_10619,N_10647);
or U10774 (N_10774,N_10629,N_10535);
nand U10775 (N_10775,N_10538,N_10557);
or U10776 (N_10776,N_10548,N_10574);
and U10777 (N_10777,N_10503,N_10619);
and U10778 (N_10778,N_10587,N_10517);
nor U10779 (N_10779,N_10525,N_10620);
and U10780 (N_10780,N_10522,N_10593);
nand U10781 (N_10781,N_10644,N_10526);
nor U10782 (N_10782,N_10553,N_10640);
nor U10783 (N_10783,N_10533,N_10517);
xor U10784 (N_10784,N_10509,N_10578);
or U10785 (N_10785,N_10589,N_10608);
or U10786 (N_10786,N_10567,N_10648);
nor U10787 (N_10787,N_10545,N_10622);
nand U10788 (N_10788,N_10585,N_10555);
nand U10789 (N_10789,N_10647,N_10578);
or U10790 (N_10790,N_10619,N_10598);
nor U10791 (N_10791,N_10507,N_10586);
nor U10792 (N_10792,N_10625,N_10605);
xor U10793 (N_10793,N_10515,N_10539);
and U10794 (N_10794,N_10549,N_10628);
nor U10795 (N_10795,N_10542,N_10636);
and U10796 (N_10796,N_10525,N_10563);
and U10797 (N_10797,N_10523,N_10501);
nand U10798 (N_10798,N_10517,N_10566);
nand U10799 (N_10799,N_10534,N_10631);
xor U10800 (N_10800,N_10749,N_10744);
and U10801 (N_10801,N_10710,N_10686);
and U10802 (N_10802,N_10776,N_10780);
nand U10803 (N_10803,N_10764,N_10735);
or U10804 (N_10804,N_10740,N_10722);
xnor U10805 (N_10805,N_10669,N_10737);
nand U10806 (N_10806,N_10704,N_10726);
and U10807 (N_10807,N_10766,N_10748);
or U10808 (N_10808,N_10676,N_10659);
nor U10809 (N_10809,N_10699,N_10653);
xnor U10810 (N_10810,N_10702,N_10689);
xor U10811 (N_10811,N_10670,N_10677);
or U10812 (N_10812,N_10660,N_10703);
nor U10813 (N_10813,N_10730,N_10658);
or U10814 (N_10814,N_10654,N_10758);
xnor U10815 (N_10815,N_10762,N_10687);
xor U10816 (N_10816,N_10727,N_10792);
or U10817 (N_10817,N_10716,N_10681);
and U10818 (N_10818,N_10650,N_10794);
and U10819 (N_10819,N_10753,N_10709);
nor U10820 (N_10820,N_10717,N_10784);
or U10821 (N_10821,N_10787,N_10663);
or U10822 (N_10822,N_10705,N_10680);
or U10823 (N_10823,N_10750,N_10739);
and U10824 (N_10824,N_10742,N_10672);
nor U10825 (N_10825,N_10746,N_10697);
and U10826 (N_10826,N_10791,N_10712);
or U10827 (N_10827,N_10668,N_10797);
nand U10828 (N_10828,N_10725,N_10711);
xor U10829 (N_10829,N_10798,N_10781);
xor U10830 (N_10830,N_10761,N_10718);
xnor U10831 (N_10831,N_10657,N_10788);
or U10832 (N_10832,N_10708,N_10664);
xor U10833 (N_10833,N_10661,N_10665);
and U10834 (N_10834,N_10651,N_10785);
nor U10835 (N_10835,N_10679,N_10724);
nor U10836 (N_10836,N_10698,N_10656);
or U10837 (N_10837,N_10775,N_10789);
and U10838 (N_10838,N_10738,N_10691);
or U10839 (N_10839,N_10729,N_10745);
nor U10840 (N_10840,N_10771,N_10770);
xnor U10841 (N_10841,N_10652,N_10695);
xor U10842 (N_10842,N_10678,N_10715);
and U10843 (N_10843,N_10682,N_10693);
or U10844 (N_10844,N_10719,N_10720);
or U10845 (N_10845,N_10694,N_10673);
xor U10846 (N_10846,N_10701,N_10741);
nor U10847 (N_10847,N_10688,N_10774);
nand U10848 (N_10848,N_10747,N_10684);
nand U10849 (N_10849,N_10706,N_10662);
xor U10850 (N_10850,N_10757,N_10713);
xnor U10851 (N_10851,N_10675,N_10765);
xor U10852 (N_10852,N_10707,N_10768);
and U10853 (N_10853,N_10767,N_10671);
and U10854 (N_10854,N_10728,N_10756);
and U10855 (N_10855,N_10733,N_10683);
or U10856 (N_10856,N_10755,N_10779);
and U10857 (N_10857,N_10793,N_10696);
or U10858 (N_10858,N_10732,N_10759);
nor U10859 (N_10859,N_10799,N_10783);
xor U10860 (N_10860,N_10790,N_10700);
and U10861 (N_10861,N_10786,N_10685);
nand U10862 (N_10862,N_10692,N_10769);
nor U10863 (N_10863,N_10721,N_10736);
nand U10864 (N_10864,N_10734,N_10723);
nor U10865 (N_10865,N_10731,N_10773);
and U10866 (N_10866,N_10667,N_10690);
nor U10867 (N_10867,N_10666,N_10795);
nand U10868 (N_10868,N_10777,N_10714);
xnor U10869 (N_10869,N_10778,N_10743);
nor U10870 (N_10870,N_10772,N_10782);
and U10871 (N_10871,N_10796,N_10754);
nor U10872 (N_10872,N_10674,N_10655);
nand U10873 (N_10873,N_10763,N_10752);
nand U10874 (N_10874,N_10751,N_10760);
or U10875 (N_10875,N_10729,N_10671);
nand U10876 (N_10876,N_10787,N_10773);
nand U10877 (N_10877,N_10710,N_10764);
nor U10878 (N_10878,N_10732,N_10768);
and U10879 (N_10879,N_10727,N_10712);
xor U10880 (N_10880,N_10679,N_10728);
xnor U10881 (N_10881,N_10744,N_10799);
or U10882 (N_10882,N_10664,N_10754);
xor U10883 (N_10883,N_10708,N_10669);
or U10884 (N_10884,N_10715,N_10685);
or U10885 (N_10885,N_10701,N_10652);
or U10886 (N_10886,N_10689,N_10753);
nor U10887 (N_10887,N_10772,N_10746);
or U10888 (N_10888,N_10794,N_10788);
or U10889 (N_10889,N_10695,N_10712);
xnor U10890 (N_10890,N_10653,N_10677);
and U10891 (N_10891,N_10695,N_10670);
nand U10892 (N_10892,N_10698,N_10670);
and U10893 (N_10893,N_10694,N_10733);
and U10894 (N_10894,N_10667,N_10657);
nand U10895 (N_10895,N_10773,N_10668);
and U10896 (N_10896,N_10679,N_10730);
nor U10897 (N_10897,N_10660,N_10783);
nor U10898 (N_10898,N_10679,N_10738);
nand U10899 (N_10899,N_10724,N_10722);
nor U10900 (N_10900,N_10780,N_10689);
nand U10901 (N_10901,N_10697,N_10739);
xor U10902 (N_10902,N_10663,N_10661);
nand U10903 (N_10903,N_10735,N_10661);
and U10904 (N_10904,N_10774,N_10668);
xor U10905 (N_10905,N_10740,N_10708);
nor U10906 (N_10906,N_10710,N_10673);
and U10907 (N_10907,N_10766,N_10721);
nor U10908 (N_10908,N_10699,N_10709);
and U10909 (N_10909,N_10764,N_10783);
nor U10910 (N_10910,N_10764,N_10723);
nor U10911 (N_10911,N_10794,N_10672);
nand U10912 (N_10912,N_10727,N_10759);
xor U10913 (N_10913,N_10791,N_10721);
nor U10914 (N_10914,N_10687,N_10742);
xnor U10915 (N_10915,N_10735,N_10797);
nand U10916 (N_10916,N_10677,N_10717);
and U10917 (N_10917,N_10684,N_10660);
nor U10918 (N_10918,N_10652,N_10678);
xnor U10919 (N_10919,N_10753,N_10707);
or U10920 (N_10920,N_10769,N_10783);
nand U10921 (N_10921,N_10704,N_10715);
and U10922 (N_10922,N_10714,N_10732);
xnor U10923 (N_10923,N_10756,N_10778);
nand U10924 (N_10924,N_10705,N_10722);
nand U10925 (N_10925,N_10798,N_10731);
nand U10926 (N_10926,N_10773,N_10714);
xnor U10927 (N_10927,N_10682,N_10666);
nand U10928 (N_10928,N_10685,N_10728);
nor U10929 (N_10929,N_10660,N_10677);
and U10930 (N_10930,N_10698,N_10734);
xnor U10931 (N_10931,N_10737,N_10730);
nand U10932 (N_10932,N_10660,N_10773);
or U10933 (N_10933,N_10770,N_10707);
nor U10934 (N_10934,N_10663,N_10678);
nand U10935 (N_10935,N_10785,N_10740);
nor U10936 (N_10936,N_10661,N_10746);
nand U10937 (N_10937,N_10705,N_10755);
and U10938 (N_10938,N_10743,N_10699);
or U10939 (N_10939,N_10742,N_10785);
and U10940 (N_10940,N_10652,N_10698);
or U10941 (N_10941,N_10659,N_10720);
nor U10942 (N_10942,N_10732,N_10795);
or U10943 (N_10943,N_10703,N_10689);
or U10944 (N_10944,N_10662,N_10770);
nand U10945 (N_10945,N_10660,N_10687);
or U10946 (N_10946,N_10753,N_10767);
xnor U10947 (N_10947,N_10741,N_10717);
nor U10948 (N_10948,N_10687,N_10696);
and U10949 (N_10949,N_10679,N_10680);
or U10950 (N_10950,N_10875,N_10939);
nand U10951 (N_10951,N_10867,N_10815);
xor U10952 (N_10952,N_10917,N_10934);
or U10953 (N_10953,N_10822,N_10912);
or U10954 (N_10954,N_10842,N_10836);
and U10955 (N_10955,N_10935,N_10904);
nand U10956 (N_10956,N_10940,N_10868);
nand U10957 (N_10957,N_10856,N_10819);
nand U10958 (N_10958,N_10808,N_10847);
nor U10959 (N_10959,N_10879,N_10941);
nor U10960 (N_10960,N_10897,N_10845);
nand U10961 (N_10961,N_10895,N_10802);
nor U10962 (N_10962,N_10841,N_10909);
or U10963 (N_10963,N_10869,N_10924);
xnor U10964 (N_10964,N_10929,N_10814);
and U10965 (N_10965,N_10886,N_10900);
xnor U10966 (N_10966,N_10820,N_10849);
or U10967 (N_10967,N_10949,N_10858);
nand U10968 (N_10968,N_10899,N_10887);
nand U10969 (N_10969,N_10848,N_10844);
nor U10970 (N_10970,N_10816,N_10916);
nor U10971 (N_10971,N_10838,N_10933);
nor U10972 (N_10972,N_10896,N_10920);
xor U10973 (N_10973,N_10829,N_10801);
and U10974 (N_10974,N_10811,N_10946);
nor U10975 (N_10975,N_10850,N_10833);
nand U10976 (N_10976,N_10905,N_10864);
and U10977 (N_10977,N_10882,N_10865);
or U10978 (N_10978,N_10945,N_10861);
nand U10979 (N_10979,N_10813,N_10884);
or U10980 (N_10980,N_10830,N_10928);
xnor U10981 (N_10981,N_10892,N_10910);
xnor U10982 (N_10982,N_10866,N_10821);
xor U10983 (N_10983,N_10834,N_10806);
xor U10984 (N_10984,N_10921,N_10872);
nand U10985 (N_10985,N_10938,N_10891);
and U10986 (N_10986,N_10889,N_10944);
or U10987 (N_10987,N_10800,N_10854);
nand U10988 (N_10988,N_10885,N_10930);
and U10989 (N_10989,N_10888,N_10831);
nor U10990 (N_10990,N_10852,N_10873);
nand U10991 (N_10991,N_10828,N_10862);
xor U10992 (N_10992,N_10870,N_10918);
nand U10993 (N_10993,N_10907,N_10926);
nand U10994 (N_10994,N_10809,N_10803);
xor U10995 (N_10995,N_10804,N_10810);
xnor U10996 (N_10996,N_10936,N_10898);
or U10997 (N_10997,N_10843,N_10937);
nand U10998 (N_10998,N_10859,N_10855);
or U10999 (N_10999,N_10948,N_10818);
nor U11000 (N_11000,N_10943,N_10927);
nand U11001 (N_11001,N_10835,N_10901);
nor U11002 (N_11002,N_10837,N_10863);
xor U11003 (N_11003,N_10902,N_10876);
nand U11004 (N_11004,N_10942,N_10817);
nor U11005 (N_11005,N_10846,N_10825);
nand U11006 (N_11006,N_10906,N_10871);
nand U11007 (N_11007,N_10913,N_10840);
and U11008 (N_11008,N_10832,N_10894);
and U11009 (N_11009,N_10923,N_10915);
nor U11010 (N_11010,N_10883,N_10911);
nand U11011 (N_11011,N_10947,N_10880);
or U11012 (N_11012,N_10826,N_10860);
nor U11013 (N_11013,N_10925,N_10890);
nor U11014 (N_11014,N_10903,N_10807);
nor U11015 (N_11015,N_10878,N_10908);
nand U11016 (N_11016,N_10853,N_10874);
or U11017 (N_11017,N_10805,N_10823);
nor U11018 (N_11018,N_10931,N_10839);
and U11019 (N_11019,N_10812,N_10824);
xor U11020 (N_11020,N_10893,N_10919);
or U11021 (N_11021,N_10914,N_10932);
nor U11022 (N_11022,N_10922,N_10877);
xor U11023 (N_11023,N_10881,N_10827);
nor U11024 (N_11024,N_10851,N_10857);
nand U11025 (N_11025,N_10847,N_10812);
xor U11026 (N_11026,N_10815,N_10809);
xnor U11027 (N_11027,N_10904,N_10903);
or U11028 (N_11028,N_10940,N_10886);
xnor U11029 (N_11029,N_10942,N_10833);
or U11030 (N_11030,N_10925,N_10876);
or U11031 (N_11031,N_10892,N_10800);
or U11032 (N_11032,N_10912,N_10824);
and U11033 (N_11033,N_10843,N_10821);
and U11034 (N_11034,N_10913,N_10875);
and U11035 (N_11035,N_10872,N_10825);
nand U11036 (N_11036,N_10854,N_10904);
nand U11037 (N_11037,N_10863,N_10804);
xnor U11038 (N_11038,N_10833,N_10871);
nor U11039 (N_11039,N_10816,N_10807);
and U11040 (N_11040,N_10852,N_10887);
and U11041 (N_11041,N_10898,N_10945);
and U11042 (N_11042,N_10902,N_10920);
xnor U11043 (N_11043,N_10945,N_10941);
xor U11044 (N_11044,N_10902,N_10842);
and U11045 (N_11045,N_10914,N_10895);
and U11046 (N_11046,N_10855,N_10913);
and U11047 (N_11047,N_10921,N_10938);
and U11048 (N_11048,N_10933,N_10852);
xnor U11049 (N_11049,N_10895,N_10933);
nand U11050 (N_11050,N_10889,N_10894);
nor U11051 (N_11051,N_10908,N_10839);
nor U11052 (N_11052,N_10923,N_10828);
nor U11053 (N_11053,N_10888,N_10800);
xnor U11054 (N_11054,N_10863,N_10833);
and U11055 (N_11055,N_10885,N_10822);
or U11056 (N_11056,N_10850,N_10852);
nor U11057 (N_11057,N_10912,N_10907);
nand U11058 (N_11058,N_10804,N_10940);
xnor U11059 (N_11059,N_10881,N_10893);
or U11060 (N_11060,N_10817,N_10856);
xor U11061 (N_11061,N_10879,N_10872);
xnor U11062 (N_11062,N_10928,N_10816);
or U11063 (N_11063,N_10892,N_10914);
and U11064 (N_11064,N_10868,N_10893);
and U11065 (N_11065,N_10898,N_10907);
nand U11066 (N_11066,N_10831,N_10833);
xor U11067 (N_11067,N_10926,N_10869);
nor U11068 (N_11068,N_10911,N_10908);
nand U11069 (N_11069,N_10897,N_10840);
and U11070 (N_11070,N_10820,N_10819);
or U11071 (N_11071,N_10925,N_10898);
nand U11072 (N_11072,N_10811,N_10805);
and U11073 (N_11073,N_10877,N_10934);
or U11074 (N_11074,N_10836,N_10841);
and U11075 (N_11075,N_10843,N_10906);
or U11076 (N_11076,N_10869,N_10806);
xor U11077 (N_11077,N_10949,N_10915);
nand U11078 (N_11078,N_10845,N_10909);
or U11079 (N_11079,N_10803,N_10921);
nand U11080 (N_11080,N_10862,N_10821);
or U11081 (N_11081,N_10931,N_10867);
nor U11082 (N_11082,N_10913,N_10899);
nor U11083 (N_11083,N_10918,N_10828);
nand U11084 (N_11084,N_10846,N_10938);
or U11085 (N_11085,N_10924,N_10897);
nand U11086 (N_11086,N_10838,N_10814);
or U11087 (N_11087,N_10932,N_10893);
or U11088 (N_11088,N_10948,N_10854);
xnor U11089 (N_11089,N_10886,N_10836);
nand U11090 (N_11090,N_10832,N_10807);
or U11091 (N_11091,N_10802,N_10827);
and U11092 (N_11092,N_10883,N_10919);
xnor U11093 (N_11093,N_10867,N_10823);
nor U11094 (N_11094,N_10891,N_10871);
or U11095 (N_11095,N_10869,N_10889);
nor U11096 (N_11096,N_10902,N_10937);
nand U11097 (N_11097,N_10886,N_10924);
nor U11098 (N_11098,N_10897,N_10884);
or U11099 (N_11099,N_10915,N_10907);
or U11100 (N_11100,N_10971,N_11020);
or U11101 (N_11101,N_11027,N_10976);
or U11102 (N_11102,N_11039,N_11053);
nand U11103 (N_11103,N_11097,N_10952);
and U11104 (N_11104,N_11089,N_11038);
or U11105 (N_11105,N_11047,N_10968);
and U11106 (N_11106,N_11067,N_11010);
or U11107 (N_11107,N_11045,N_11029);
nor U11108 (N_11108,N_10999,N_10963);
or U11109 (N_11109,N_11095,N_11012);
or U11110 (N_11110,N_10987,N_10973);
nor U11111 (N_11111,N_10961,N_11003);
nor U11112 (N_11112,N_11011,N_11034);
nand U11113 (N_11113,N_11057,N_11079);
or U11114 (N_11114,N_11071,N_11063);
nor U11115 (N_11115,N_10960,N_11052);
or U11116 (N_11116,N_11051,N_11030);
xnor U11117 (N_11117,N_10950,N_11078);
or U11118 (N_11118,N_11002,N_10974);
or U11119 (N_11119,N_11035,N_11069);
and U11120 (N_11120,N_11036,N_10955);
nand U11121 (N_11121,N_11028,N_10975);
nand U11122 (N_11122,N_11000,N_11022);
nand U11123 (N_11123,N_11065,N_11004);
or U11124 (N_11124,N_11080,N_11046);
or U11125 (N_11125,N_11043,N_10993);
and U11126 (N_11126,N_11096,N_10954);
and U11127 (N_11127,N_10967,N_11061);
nand U11128 (N_11128,N_11006,N_11016);
or U11129 (N_11129,N_11007,N_10977);
nand U11130 (N_11130,N_11032,N_11083);
nor U11131 (N_11131,N_11001,N_11018);
or U11132 (N_11132,N_11099,N_11040);
and U11133 (N_11133,N_11056,N_10959);
nand U11134 (N_11134,N_11091,N_11074);
and U11135 (N_11135,N_11021,N_10991);
nor U11136 (N_11136,N_10982,N_11055);
nor U11137 (N_11137,N_10957,N_10965);
and U11138 (N_11138,N_11009,N_11086);
and U11139 (N_11139,N_10994,N_11090);
nor U11140 (N_11140,N_11075,N_10962);
or U11141 (N_11141,N_11084,N_11026);
and U11142 (N_11142,N_10970,N_11054);
xnor U11143 (N_11143,N_10985,N_11094);
nor U11144 (N_11144,N_11014,N_11025);
nand U11145 (N_11145,N_11093,N_10964);
or U11146 (N_11146,N_11072,N_10956);
nand U11147 (N_11147,N_10986,N_11042);
nor U11148 (N_11148,N_11019,N_10978);
nand U11149 (N_11149,N_10996,N_11066);
nand U11150 (N_11150,N_11059,N_11037);
or U11151 (N_11151,N_11044,N_11058);
xor U11152 (N_11152,N_11024,N_11050);
and U11153 (N_11153,N_10980,N_10997);
and U11154 (N_11154,N_10990,N_10951);
and U11155 (N_11155,N_11031,N_11088);
or U11156 (N_11156,N_11008,N_11064);
or U11157 (N_11157,N_10989,N_10972);
nor U11158 (N_11158,N_11062,N_10992);
and U11159 (N_11159,N_10983,N_11098);
and U11160 (N_11160,N_10979,N_11023);
nand U11161 (N_11161,N_11005,N_11081);
and U11162 (N_11162,N_10988,N_10995);
nand U11163 (N_11163,N_11017,N_10998);
and U11164 (N_11164,N_11041,N_11092);
nand U11165 (N_11165,N_10981,N_11070);
or U11166 (N_11166,N_11033,N_11013);
nand U11167 (N_11167,N_10966,N_11049);
xnor U11168 (N_11168,N_11068,N_10969);
and U11169 (N_11169,N_11082,N_10984);
and U11170 (N_11170,N_11087,N_11015);
or U11171 (N_11171,N_11085,N_11076);
and U11172 (N_11172,N_11048,N_11077);
or U11173 (N_11173,N_11060,N_10958);
or U11174 (N_11174,N_11073,N_10953);
and U11175 (N_11175,N_11023,N_11041);
nor U11176 (N_11176,N_10988,N_11004);
or U11177 (N_11177,N_11015,N_11029);
or U11178 (N_11178,N_10998,N_11003);
xor U11179 (N_11179,N_10966,N_10952);
nor U11180 (N_11180,N_11097,N_11000);
nand U11181 (N_11181,N_10969,N_10987);
xnor U11182 (N_11182,N_10994,N_10952);
xnor U11183 (N_11183,N_10982,N_11062);
xor U11184 (N_11184,N_11043,N_11054);
nand U11185 (N_11185,N_10991,N_11097);
and U11186 (N_11186,N_11023,N_10980);
xnor U11187 (N_11187,N_11055,N_11020);
and U11188 (N_11188,N_11076,N_11011);
xor U11189 (N_11189,N_10997,N_11018);
xor U11190 (N_11190,N_11084,N_11069);
or U11191 (N_11191,N_11039,N_10977);
nand U11192 (N_11192,N_11070,N_11086);
nand U11193 (N_11193,N_11098,N_11096);
or U11194 (N_11194,N_11014,N_10951);
nand U11195 (N_11195,N_11005,N_10988);
and U11196 (N_11196,N_11001,N_10988);
xor U11197 (N_11197,N_11004,N_10985);
nand U11198 (N_11198,N_11079,N_11097);
or U11199 (N_11199,N_10992,N_11056);
or U11200 (N_11200,N_11026,N_10961);
nand U11201 (N_11201,N_10967,N_10995);
xor U11202 (N_11202,N_10964,N_11009);
and U11203 (N_11203,N_11078,N_11051);
xor U11204 (N_11204,N_11021,N_11090);
xor U11205 (N_11205,N_11012,N_11093);
and U11206 (N_11206,N_10958,N_10959);
nor U11207 (N_11207,N_11050,N_11082);
xnor U11208 (N_11208,N_11020,N_10955);
xor U11209 (N_11209,N_10987,N_11096);
and U11210 (N_11210,N_10992,N_11065);
or U11211 (N_11211,N_11001,N_11024);
xnor U11212 (N_11212,N_11044,N_11051);
nor U11213 (N_11213,N_11025,N_11042);
or U11214 (N_11214,N_11004,N_11075);
xor U11215 (N_11215,N_10960,N_11087);
nor U11216 (N_11216,N_11042,N_11021);
nand U11217 (N_11217,N_11086,N_11097);
xor U11218 (N_11218,N_11041,N_11054);
xor U11219 (N_11219,N_10990,N_11088);
and U11220 (N_11220,N_10954,N_10953);
nand U11221 (N_11221,N_11037,N_10950);
nor U11222 (N_11222,N_10987,N_11034);
or U11223 (N_11223,N_11092,N_11007);
and U11224 (N_11224,N_11060,N_11049);
nand U11225 (N_11225,N_11031,N_11050);
nand U11226 (N_11226,N_11054,N_10994);
and U11227 (N_11227,N_11038,N_11003);
nand U11228 (N_11228,N_10986,N_10978);
nor U11229 (N_11229,N_11083,N_10955);
or U11230 (N_11230,N_10972,N_11076);
or U11231 (N_11231,N_10995,N_11011);
and U11232 (N_11232,N_11022,N_11018);
nand U11233 (N_11233,N_11022,N_11090);
and U11234 (N_11234,N_10957,N_11002);
and U11235 (N_11235,N_11072,N_11006);
and U11236 (N_11236,N_11006,N_11030);
or U11237 (N_11237,N_10971,N_11028);
or U11238 (N_11238,N_11058,N_10987);
nor U11239 (N_11239,N_11014,N_11083);
and U11240 (N_11240,N_11084,N_11070);
nand U11241 (N_11241,N_11000,N_11014);
and U11242 (N_11242,N_10972,N_11037);
and U11243 (N_11243,N_10995,N_11087);
nor U11244 (N_11244,N_11036,N_11022);
and U11245 (N_11245,N_11029,N_10956);
nand U11246 (N_11246,N_11006,N_10966);
nor U11247 (N_11247,N_11072,N_11061);
nand U11248 (N_11248,N_11002,N_11055);
nor U11249 (N_11249,N_11070,N_11069);
or U11250 (N_11250,N_11165,N_11100);
nor U11251 (N_11251,N_11155,N_11151);
or U11252 (N_11252,N_11223,N_11131);
or U11253 (N_11253,N_11113,N_11207);
and U11254 (N_11254,N_11139,N_11211);
nor U11255 (N_11255,N_11200,N_11157);
nor U11256 (N_11256,N_11212,N_11105);
nor U11257 (N_11257,N_11232,N_11145);
and U11258 (N_11258,N_11176,N_11146);
xnor U11259 (N_11259,N_11134,N_11201);
nor U11260 (N_11260,N_11241,N_11199);
xnor U11261 (N_11261,N_11189,N_11156);
xnor U11262 (N_11262,N_11152,N_11205);
nor U11263 (N_11263,N_11138,N_11194);
nor U11264 (N_11264,N_11107,N_11214);
xnor U11265 (N_11265,N_11112,N_11160);
nand U11266 (N_11266,N_11153,N_11149);
and U11267 (N_11267,N_11221,N_11147);
nand U11268 (N_11268,N_11158,N_11116);
and U11269 (N_11269,N_11186,N_11137);
and U11270 (N_11270,N_11150,N_11249);
and U11271 (N_11271,N_11124,N_11173);
and U11272 (N_11272,N_11119,N_11120);
or U11273 (N_11273,N_11135,N_11210);
xor U11274 (N_11274,N_11202,N_11225);
and U11275 (N_11275,N_11180,N_11140);
and U11276 (N_11276,N_11148,N_11191);
xor U11277 (N_11277,N_11236,N_11233);
nor U11278 (N_11278,N_11170,N_11108);
xor U11279 (N_11279,N_11182,N_11215);
or U11280 (N_11280,N_11248,N_11118);
nor U11281 (N_11281,N_11141,N_11183);
nor U11282 (N_11282,N_11220,N_11187);
nor U11283 (N_11283,N_11122,N_11192);
nand U11284 (N_11284,N_11123,N_11101);
nand U11285 (N_11285,N_11216,N_11130);
or U11286 (N_11286,N_11197,N_11244);
nor U11287 (N_11287,N_11127,N_11240);
or U11288 (N_11288,N_11188,N_11247);
xor U11289 (N_11289,N_11229,N_11179);
and U11290 (N_11290,N_11204,N_11164);
xnor U11291 (N_11291,N_11174,N_11227);
nand U11292 (N_11292,N_11136,N_11195);
and U11293 (N_11293,N_11239,N_11129);
nor U11294 (N_11294,N_11208,N_11242);
nand U11295 (N_11295,N_11166,N_11217);
nand U11296 (N_11296,N_11198,N_11171);
or U11297 (N_11297,N_11163,N_11162);
or U11298 (N_11298,N_11161,N_11209);
xnor U11299 (N_11299,N_11237,N_11159);
xnor U11300 (N_11300,N_11111,N_11103);
nor U11301 (N_11301,N_11117,N_11109);
nor U11302 (N_11302,N_11193,N_11102);
xnor U11303 (N_11303,N_11178,N_11224);
xnor U11304 (N_11304,N_11169,N_11184);
or U11305 (N_11305,N_11190,N_11177);
xnor U11306 (N_11306,N_11106,N_11246);
xor U11307 (N_11307,N_11115,N_11167);
nand U11308 (N_11308,N_11230,N_11226);
xnor U11309 (N_11309,N_11185,N_11172);
nand U11310 (N_11310,N_11114,N_11231);
or U11311 (N_11311,N_11196,N_11175);
nor U11312 (N_11312,N_11125,N_11168);
nand U11313 (N_11313,N_11142,N_11132);
and U11314 (N_11314,N_11238,N_11110);
xnor U11315 (N_11315,N_11203,N_11245);
or U11316 (N_11316,N_11235,N_11213);
or U11317 (N_11317,N_11121,N_11234);
and U11318 (N_11318,N_11104,N_11243);
xor U11319 (N_11319,N_11218,N_11228);
and U11320 (N_11320,N_11206,N_11154);
nand U11321 (N_11321,N_11143,N_11128);
or U11322 (N_11322,N_11126,N_11219);
nor U11323 (N_11323,N_11181,N_11144);
nor U11324 (N_11324,N_11222,N_11133);
or U11325 (N_11325,N_11230,N_11105);
or U11326 (N_11326,N_11139,N_11220);
nor U11327 (N_11327,N_11186,N_11230);
and U11328 (N_11328,N_11203,N_11205);
or U11329 (N_11329,N_11161,N_11110);
nand U11330 (N_11330,N_11168,N_11117);
xnor U11331 (N_11331,N_11105,N_11243);
or U11332 (N_11332,N_11192,N_11112);
xnor U11333 (N_11333,N_11191,N_11165);
or U11334 (N_11334,N_11202,N_11207);
nand U11335 (N_11335,N_11103,N_11142);
and U11336 (N_11336,N_11155,N_11205);
nor U11337 (N_11337,N_11194,N_11245);
nand U11338 (N_11338,N_11168,N_11199);
nand U11339 (N_11339,N_11225,N_11110);
and U11340 (N_11340,N_11139,N_11173);
or U11341 (N_11341,N_11128,N_11208);
or U11342 (N_11342,N_11115,N_11151);
nand U11343 (N_11343,N_11182,N_11116);
nor U11344 (N_11344,N_11245,N_11112);
nand U11345 (N_11345,N_11227,N_11110);
nand U11346 (N_11346,N_11229,N_11205);
xor U11347 (N_11347,N_11239,N_11225);
nand U11348 (N_11348,N_11249,N_11156);
or U11349 (N_11349,N_11128,N_11227);
or U11350 (N_11350,N_11184,N_11120);
nor U11351 (N_11351,N_11249,N_11154);
nor U11352 (N_11352,N_11109,N_11227);
or U11353 (N_11353,N_11131,N_11143);
or U11354 (N_11354,N_11105,N_11109);
nor U11355 (N_11355,N_11239,N_11237);
xnor U11356 (N_11356,N_11194,N_11226);
xnor U11357 (N_11357,N_11144,N_11193);
xnor U11358 (N_11358,N_11219,N_11109);
nor U11359 (N_11359,N_11178,N_11142);
or U11360 (N_11360,N_11230,N_11106);
nand U11361 (N_11361,N_11224,N_11159);
nor U11362 (N_11362,N_11160,N_11243);
and U11363 (N_11363,N_11188,N_11105);
and U11364 (N_11364,N_11119,N_11162);
nor U11365 (N_11365,N_11116,N_11179);
nor U11366 (N_11366,N_11129,N_11183);
nor U11367 (N_11367,N_11167,N_11193);
and U11368 (N_11368,N_11211,N_11177);
xor U11369 (N_11369,N_11150,N_11136);
or U11370 (N_11370,N_11136,N_11123);
and U11371 (N_11371,N_11156,N_11117);
nand U11372 (N_11372,N_11209,N_11249);
nand U11373 (N_11373,N_11186,N_11238);
nor U11374 (N_11374,N_11188,N_11148);
nor U11375 (N_11375,N_11124,N_11203);
nand U11376 (N_11376,N_11126,N_11130);
or U11377 (N_11377,N_11144,N_11189);
nand U11378 (N_11378,N_11196,N_11217);
and U11379 (N_11379,N_11142,N_11147);
nor U11380 (N_11380,N_11186,N_11237);
nand U11381 (N_11381,N_11147,N_11167);
nor U11382 (N_11382,N_11125,N_11162);
nand U11383 (N_11383,N_11223,N_11129);
or U11384 (N_11384,N_11112,N_11105);
xnor U11385 (N_11385,N_11119,N_11227);
and U11386 (N_11386,N_11219,N_11124);
and U11387 (N_11387,N_11173,N_11143);
nand U11388 (N_11388,N_11131,N_11182);
or U11389 (N_11389,N_11118,N_11128);
xnor U11390 (N_11390,N_11212,N_11156);
nand U11391 (N_11391,N_11173,N_11107);
or U11392 (N_11392,N_11185,N_11100);
xnor U11393 (N_11393,N_11184,N_11156);
xor U11394 (N_11394,N_11142,N_11149);
and U11395 (N_11395,N_11192,N_11235);
or U11396 (N_11396,N_11128,N_11129);
nor U11397 (N_11397,N_11156,N_11169);
nand U11398 (N_11398,N_11153,N_11137);
and U11399 (N_11399,N_11185,N_11247);
nand U11400 (N_11400,N_11326,N_11271);
or U11401 (N_11401,N_11316,N_11353);
xor U11402 (N_11402,N_11373,N_11253);
nand U11403 (N_11403,N_11375,N_11277);
nand U11404 (N_11404,N_11259,N_11365);
xor U11405 (N_11405,N_11343,N_11389);
xor U11406 (N_11406,N_11301,N_11341);
or U11407 (N_11407,N_11305,N_11297);
or U11408 (N_11408,N_11381,N_11325);
xnor U11409 (N_11409,N_11289,N_11399);
xnor U11410 (N_11410,N_11314,N_11269);
xor U11411 (N_11411,N_11318,N_11355);
and U11412 (N_11412,N_11321,N_11279);
or U11413 (N_11413,N_11327,N_11354);
or U11414 (N_11414,N_11283,N_11296);
nor U11415 (N_11415,N_11308,N_11350);
and U11416 (N_11416,N_11292,N_11342);
nor U11417 (N_11417,N_11303,N_11336);
nand U11418 (N_11418,N_11281,N_11357);
and U11419 (N_11419,N_11364,N_11309);
nor U11420 (N_11420,N_11284,N_11311);
nand U11421 (N_11421,N_11310,N_11356);
and U11422 (N_11422,N_11258,N_11291);
nor U11423 (N_11423,N_11319,N_11278);
xnor U11424 (N_11424,N_11387,N_11392);
or U11425 (N_11425,N_11359,N_11377);
xor U11426 (N_11426,N_11393,N_11367);
and U11427 (N_11427,N_11374,N_11264);
nand U11428 (N_11428,N_11280,N_11252);
nand U11429 (N_11429,N_11371,N_11391);
or U11430 (N_11430,N_11340,N_11385);
or U11431 (N_11431,N_11332,N_11388);
nand U11432 (N_11432,N_11282,N_11302);
nand U11433 (N_11433,N_11329,N_11363);
and U11434 (N_11434,N_11338,N_11304);
nand U11435 (N_11435,N_11260,N_11299);
xnor U11436 (N_11436,N_11382,N_11267);
and U11437 (N_11437,N_11268,N_11306);
nor U11438 (N_11438,N_11369,N_11315);
xor U11439 (N_11439,N_11257,N_11368);
or U11440 (N_11440,N_11294,N_11361);
or U11441 (N_11441,N_11328,N_11300);
nand U11442 (N_11442,N_11345,N_11394);
xor U11443 (N_11443,N_11396,N_11372);
xor U11444 (N_11444,N_11376,N_11288);
and U11445 (N_11445,N_11322,N_11285);
nor U11446 (N_11446,N_11378,N_11358);
xnor U11447 (N_11447,N_11380,N_11383);
and U11448 (N_11448,N_11255,N_11276);
xor U11449 (N_11449,N_11251,N_11379);
xnor U11450 (N_11450,N_11333,N_11397);
nand U11451 (N_11451,N_11348,N_11395);
xor U11452 (N_11452,N_11256,N_11324);
and U11453 (N_11453,N_11320,N_11262);
and U11454 (N_11454,N_11335,N_11265);
and U11455 (N_11455,N_11366,N_11312);
nor U11456 (N_11456,N_11286,N_11293);
nand U11457 (N_11457,N_11274,N_11384);
xnor U11458 (N_11458,N_11370,N_11347);
xnor U11459 (N_11459,N_11272,N_11287);
xnor U11460 (N_11460,N_11337,N_11254);
nor U11461 (N_11461,N_11261,N_11351);
or U11462 (N_11462,N_11330,N_11250);
xor U11463 (N_11463,N_11360,N_11263);
xor U11464 (N_11464,N_11386,N_11390);
and U11465 (N_11465,N_11298,N_11339);
nor U11466 (N_11466,N_11313,N_11317);
or U11467 (N_11467,N_11275,N_11307);
or U11468 (N_11468,N_11352,N_11331);
nor U11469 (N_11469,N_11270,N_11362);
xor U11470 (N_11470,N_11349,N_11344);
nand U11471 (N_11471,N_11334,N_11273);
xor U11472 (N_11472,N_11290,N_11295);
nand U11473 (N_11473,N_11323,N_11346);
or U11474 (N_11474,N_11398,N_11266);
xor U11475 (N_11475,N_11316,N_11292);
nand U11476 (N_11476,N_11317,N_11378);
xor U11477 (N_11477,N_11273,N_11329);
xor U11478 (N_11478,N_11374,N_11306);
or U11479 (N_11479,N_11396,N_11255);
nor U11480 (N_11480,N_11360,N_11274);
and U11481 (N_11481,N_11362,N_11374);
nor U11482 (N_11482,N_11272,N_11359);
xnor U11483 (N_11483,N_11394,N_11264);
or U11484 (N_11484,N_11382,N_11362);
and U11485 (N_11485,N_11252,N_11384);
xor U11486 (N_11486,N_11285,N_11308);
nand U11487 (N_11487,N_11353,N_11282);
and U11488 (N_11488,N_11334,N_11258);
nand U11489 (N_11489,N_11330,N_11254);
xnor U11490 (N_11490,N_11270,N_11300);
and U11491 (N_11491,N_11301,N_11286);
nand U11492 (N_11492,N_11355,N_11295);
nand U11493 (N_11493,N_11290,N_11277);
nor U11494 (N_11494,N_11332,N_11285);
or U11495 (N_11495,N_11385,N_11341);
xor U11496 (N_11496,N_11375,N_11309);
xnor U11497 (N_11497,N_11262,N_11275);
nor U11498 (N_11498,N_11382,N_11358);
nor U11499 (N_11499,N_11370,N_11337);
xnor U11500 (N_11500,N_11324,N_11363);
nor U11501 (N_11501,N_11331,N_11372);
nor U11502 (N_11502,N_11257,N_11326);
xor U11503 (N_11503,N_11343,N_11325);
nand U11504 (N_11504,N_11397,N_11309);
or U11505 (N_11505,N_11318,N_11364);
or U11506 (N_11506,N_11280,N_11372);
or U11507 (N_11507,N_11272,N_11345);
nor U11508 (N_11508,N_11320,N_11303);
and U11509 (N_11509,N_11342,N_11251);
nor U11510 (N_11510,N_11371,N_11281);
and U11511 (N_11511,N_11339,N_11335);
nor U11512 (N_11512,N_11304,N_11339);
nor U11513 (N_11513,N_11398,N_11293);
nor U11514 (N_11514,N_11385,N_11395);
xor U11515 (N_11515,N_11309,N_11314);
and U11516 (N_11516,N_11268,N_11255);
and U11517 (N_11517,N_11339,N_11317);
xnor U11518 (N_11518,N_11254,N_11290);
or U11519 (N_11519,N_11393,N_11386);
or U11520 (N_11520,N_11332,N_11264);
nor U11521 (N_11521,N_11310,N_11288);
nor U11522 (N_11522,N_11384,N_11310);
nand U11523 (N_11523,N_11325,N_11371);
or U11524 (N_11524,N_11399,N_11312);
or U11525 (N_11525,N_11330,N_11378);
or U11526 (N_11526,N_11371,N_11268);
and U11527 (N_11527,N_11273,N_11351);
nand U11528 (N_11528,N_11365,N_11345);
nand U11529 (N_11529,N_11319,N_11375);
xnor U11530 (N_11530,N_11267,N_11354);
or U11531 (N_11531,N_11349,N_11347);
nor U11532 (N_11532,N_11315,N_11318);
xor U11533 (N_11533,N_11383,N_11371);
and U11534 (N_11534,N_11377,N_11252);
nand U11535 (N_11535,N_11279,N_11253);
or U11536 (N_11536,N_11364,N_11382);
or U11537 (N_11537,N_11360,N_11299);
nor U11538 (N_11538,N_11262,N_11279);
nand U11539 (N_11539,N_11377,N_11313);
and U11540 (N_11540,N_11337,N_11264);
or U11541 (N_11541,N_11350,N_11256);
nand U11542 (N_11542,N_11371,N_11287);
nor U11543 (N_11543,N_11252,N_11258);
and U11544 (N_11544,N_11397,N_11292);
and U11545 (N_11545,N_11265,N_11352);
nand U11546 (N_11546,N_11300,N_11271);
xor U11547 (N_11547,N_11257,N_11299);
or U11548 (N_11548,N_11355,N_11277);
nand U11549 (N_11549,N_11364,N_11320);
or U11550 (N_11550,N_11463,N_11543);
nor U11551 (N_11551,N_11447,N_11528);
xnor U11552 (N_11552,N_11436,N_11459);
nand U11553 (N_11553,N_11465,N_11413);
and U11554 (N_11554,N_11522,N_11549);
nor U11555 (N_11555,N_11441,N_11501);
nor U11556 (N_11556,N_11416,N_11453);
and U11557 (N_11557,N_11456,N_11542);
and U11558 (N_11558,N_11534,N_11492);
nand U11559 (N_11559,N_11427,N_11530);
nand U11560 (N_11560,N_11423,N_11420);
or U11561 (N_11561,N_11434,N_11428);
or U11562 (N_11562,N_11460,N_11502);
and U11563 (N_11563,N_11514,N_11446);
xor U11564 (N_11564,N_11499,N_11497);
or U11565 (N_11565,N_11476,N_11535);
or U11566 (N_11566,N_11520,N_11517);
or U11567 (N_11567,N_11518,N_11412);
xnor U11568 (N_11568,N_11479,N_11449);
nor U11569 (N_11569,N_11506,N_11452);
xor U11570 (N_11570,N_11400,N_11486);
or U11571 (N_11571,N_11414,N_11471);
and U11572 (N_11572,N_11533,N_11536);
nor U11573 (N_11573,N_11515,N_11541);
nor U11574 (N_11574,N_11487,N_11401);
nor U11575 (N_11575,N_11407,N_11405);
nand U11576 (N_11576,N_11538,N_11418);
or U11577 (N_11577,N_11509,N_11417);
and U11578 (N_11578,N_11488,N_11429);
and U11579 (N_11579,N_11500,N_11433);
nor U11580 (N_11580,N_11482,N_11450);
or U11581 (N_11581,N_11448,N_11512);
xnor U11582 (N_11582,N_11409,N_11466);
and U11583 (N_11583,N_11451,N_11524);
xnor U11584 (N_11584,N_11510,N_11516);
or U11585 (N_11585,N_11489,N_11521);
nor U11586 (N_11586,N_11472,N_11508);
nand U11587 (N_11587,N_11504,N_11493);
and U11588 (N_11588,N_11546,N_11519);
nand U11589 (N_11589,N_11545,N_11505);
nor U11590 (N_11590,N_11495,N_11547);
or U11591 (N_11591,N_11415,N_11437);
xor U11592 (N_11592,N_11511,N_11445);
nand U11593 (N_11593,N_11419,N_11531);
nor U11594 (N_11594,N_11426,N_11503);
nor U11595 (N_11595,N_11411,N_11540);
xor U11596 (N_11596,N_11457,N_11484);
xor U11597 (N_11597,N_11548,N_11478);
or U11598 (N_11598,N_11527,N_11431);
nand U11599 (N_11599,N_11422,N_11403);
or U11600 (N_11600,N_11438,N_11485);
or U11601 (N_11601,N_11539,N_11458);
or U11602 (N_11602,N_11523,N_11408);
or U11603 (N_11603,N_11532,N_11462);
nand U11604 (N_11604,N_11498,N_11402);
nand U11605 (N_11605,N_11469,N_11490);
or U11606 (N_11606,N_11442,N_11425);
xor U11607 (N_11607,N_11410,N_11421);
nand U11608 (N_11608,N_11481,N_11475);
nor U11609 (N_11609,N_11439,N_11496);
or U11610 (N_11610,N_11529,N_11443);
nand U11611 (N_11611,N_11526,N_11473);
and U11612 (N_11612,N_11544,N_11513);
xnor U11613 (N_11613,N_11537,N_11435);
or U11614 (N_11614,N_11424,N_11430);
and U11615 (N_11615,N_11483,N_11474);
or U11616 (N_11616,N_11432,N_11468);
nor U11617 (N_11617,N_11477,N_11444);
and U11618 (N_11618,N_11461,N_11406);
and U11619 (N_11619,N_11454,N_11470);
xor U11620 (N_11620,N_11525,N_11404);
xnor U11621 (N_11621,N_11494,N_11455);
or U11622 (N_11622,N_11467,N_11464);
xnor U11623 (N_11623,N_11507,N_11440);
or U11624 (N_11624,N_11480,N_11491);
nand U11625 (N_11625,N_11523,N_11401);
and U11626 (N_11626,N_11532,N_11540);
or U11627 (N_11627,N_11403,N_11488);
and U11628 (N_11628,N_11540,N_11510);
xnor U11629 (N_11629,N_11540,N_11529);
xnor U11630 (N_11630,N_11408,N_11450);
nand U11631 (N_11631,N_11547,N_11549);
and U11632 (N_11632,N_11469,N_11459);
nor U11633 (N_11633,N_11416,N_11437);
or U11634 (N_11634,N_11469,N_11463);
or U11635 (N_11635,N_11506,N_11412);
xor U11636 (N_11636,N_11427,N_11406);
and U11637 (N_11637,N_11488,N_11406);
and U11638 (N_11638,N_11409,N_11539);
xnor U11639 (N_11639,N_11511,N_11432);
or U11640 (N_11640,N_11484,N_11449);
and U11641 (N_11641,N_11517,N_11475);
or U11642 (N_11642,N_11515,N_11453);
and U11643 (N_11643,N_11530,N_11409);
nand U11644 (N_11644,N_11430,N_11537);
or U11645 (N_11645,N_11421,N_11480);
nand U11646 (N_11646,N_11474,N_11545);
nor U11647 (N_11647,N_11444,N_11438);
and U11648 (N_11648,N_11436,N_11455);
nand U11649 (N_11649,N_11480,N_11439);
xor U11650 (N_11650,N_11535,N_11478);
nand U11651 (N_11651,N_11422,N_11416);
or U11652 (N_11652,N_11420,N_11464);
or U11653 (N_11653,N_11503,N_11545);
nor U11654 (N_11654,N_11538,N_11421);
xnor U11655 (N_11655,N_11486,N_11431);
or U11656 (N_11656,N_11507,N_11413);
and U11657 (N_11657,N_11547,N_11548);
and U11658 (N_11658,N_11478,N_11526);
xnor U11659 (N_11659,N_11437,N_11500);
nor U11660 (N_11660,N_11452,N_11534);
and U11661 (N_11661,N_11400,N_11519);
xor U11662 (N_11662,N_11548,N_11515);
nand U11663 (N_11663,N_11511,N_11435);
nand U11664 (N_11664,N_11495,N_11540);
and U11665 (N_11665,N_11401,N_11529);
nand U11666 (N_11666,N_11457,N_11531);
xor U11667 (N_11667,N_11402,N_11485);
xnor U11668 (N_11668,N_11499,N_11434);
nand U11669 (N_11669,N_11469,N_11440);
nor U11670 (N_11670,N_11519,N_11527);
or U11671 (N_11671,N_11447,N_11536);
nor U11672 (N_11672,N_11516,N_11502);
nor U11673 (N_11673,N_11466,N_11487);
and U11674 (N_11674,N_11540,N_11515);
xor U11675 (N_11675,N_11433,N_11443);
and U11676 (N_11676,N_11535,N_11505);
xnor U11677 (N_11677,N_11496,N_11532);
nand U11678 (N_11678,N_11433,N_11446);
nand U11679 (N_11679,N_11478,N_11536);
xnor U11680 (N_11680,N_11454,N_11478);
and U11681 (N_11681,N_11548,N_11549);
xnor U11682 (N_11682,N_11424,N_11439);
and U11683 (N_11683,N_11472,N_11529);
xor U11684 (N_11684,N_11447,N_11494);
nand U11685 (N_11685,N_11533,N_11400);
nand U11686 (N_11686,N_11500,N_11401);
or U11687 (N_11687,N_11418,N_11411);
nand U11688 (N_11688,N_11538,N_11426);
nor U11689 (N_11689,N_11436,N_11406);
nand U11690 (N_11690,N_11412,N_11409);
xor U11691 (N_11691,N_11433,N_11414);
xnor U11692 (N_11692,N_11534,N_11521);
xor U11693 (N_11693,N_11482,N_11479);
and U11694 (N_11694,N_11481,N_11549);
or U11695 (N_11695,N_11416,N_11414);
nand U11696 (N_11696,N_11441,N_11455);
nand U11697 (N_11697,N_11548,N_11493);
xnor U11698 (N_11698,N_11427,N_11468);
nand U11699 (N_11699,N_11480,N_11535);
xnor U11700 (N_11700,N_11675,N_11626);
or U11701 (N_11701,N_11649,N_11584);
xnor U11702 (N_11702,N_11680,N_11555);
xnor U11703 (N_11703,N_11678,N_11639);
nand U11704 (N_11704,N_11607,N_11598);
and U11705 (N_11705,N_11662,N_11660);
xnor U11706 (N_11706,N_11677,N_11617);
nor U11707 (N_11707,N_11581,N_11663);
nand U11708 (N_11708,N_11577,N_11631);
nand U11709 (N_11709,N_11633,N_11627);
nand U11710 (N_11710,N_11676,N_11600);
nand U11711 (N_11711,N_11624,N_11654);
and U11712 (N_11712,N_11593,N_11690);
and U11713 (N_11713,N_11602,N_11621);
and U11714 (N_11714,N_11687,N_11636);
xnor U11715 (N_11715,N_11592,N_11559);
or U11716 (N_11716,N_11553,N_11669);
nand U11717 (N_11717,N_11688,N_11657);
nor U11718 (N_11718,N_11638,N_11562);
and U11719 (N_11719,N_11557,N_11574);
and U11720 (N_11720,N_11670,N_11618);
nand U11721 (N_11721,N_11583,N_11647);
nor U11722 (N_11722,N_11629,N_11685);
and U11723 (N_11723,N_11613,N_11697);
or U11724 (N_11724,N_11573,N_11561);
xnor U11725 (N_11725,N_11619,N_11576);
or U11726 (N_11726,N_11643,N_11665);
and U11727 (N_11727,N_11595,N_11637);
or U11728 (N_11728,N_11611,N_11601);
xnor U11729 (N_11729,N_11625,N_11578);
nor U11730 (N_11730,N_11692,N_11644);
or U11731 (N_11731,N_11575,N_11572);
or U11732 (N_11732,N_11566,N_11653);
nand U11733 (N_11733,N_11668,N_11696);
xor U11734 (N_11734,N_11609,N_11604);
nor U11735 (N_11735,N_11641,N_11579);
or U11736 (N_11736,N_11642,N_11655);
nand U11737 (N_11737,N_11664,N_11659);
xor U11738 (N_11738,N_11610,N_11686);
or U11739 (N_11739,N_11605,N_11681);
or U11740 (N_11740,N_11674,N_11556);
nor U11741 (N_11741,N_11567,N_11623);
nand U11742 (N_11742,N_11563,N_11699);
nand U11743 (N_11743,N_11606,N_11558);
nor U11744 (N_11744,N_11596,N_11672);
xnor U11745 (N_11745,N_11679,N_11634);
nand U11746 (N_11746,N_11661,N_11698);
nand U11747 (N_11747,N_11691,N_11586);
and U11748 (N_11748,N_11622,N_11694);
xor U11749 (N_11749,N_11569,N_11554);
xor U11750 (N_11750,N_11570,N_11552);
and U11751 (N_11751,N_11614,N_11652);
or U11752 (N_11752,N_11599,N_11673);
nand U11753 (N_11753,N_11615,N_11571);
and U11754 (N_11754,N_11565,N_11648);
xor U11755 (N_11755,N_11628,N_11588);
xnor U11756 (N_11756,N_11568,N_11589);
nand U11757 (N_11757,N_11630,N_11587);
and U11758 (N_11758,N_11551,N_11656);
and U11759 (N_11759,N_11645,N_11671);
nand U11760 (N_11760,N_11646,N_11612);
nor U11761 (N_11761,N_11684,N_11640);
xor U11762 (N_11762,N_11590,N_11608);
nand U11763 (N_11763,N_11580,N_11667);
xnor U11764 (N_11764,N_11620,N_11582);
and U11765 (N_11765,N_11650,N_11666);
or U11766 (N_11766,N_11635,N_11560);
nor U11767 (N_11767,N_11594,N_11658);
nor U11768 (N_11768,N_11651,N_11603);
xor U11769 (N_11769,N_11564,N_11616);
and U11770 (N_11770,N_11597,N_11693);
xor U11771 (N_11771,N_11591,N_11695);
nand U11772 (N_11772,N_11550,N_11682);
and U11773 (N_11773,N_11632,N_11585);
xnor U11774 (N_11774,N_11683,N_11689);
nand U11775 (N_11775,N_11696,N_11663);
and U11776 (N_11776,N_11643,N_11590);
nor U11777 (N_11777,N_11685,N_11683);
and U11778 (N_11778,N_11658,N_11684);
xnor U11779 (N_11779,N_11657,N_11645);
or U11780 (N_11780,N_11615,N_11576);
nor U11781 (N_11781,N_11654,N_11687);
nand U11782 (N_11782,N_11595,N_11649);
nor U11783 (N_11783,N_11629,N_11696);
and U11784 (N_11784,N_11610,N_11697);
nand U11785 (N_11785,N_11674,N_11569);
nor U11786 (N_11786,N_11696,N_11598);
or U11787 (N_11787,N_11588,N_11680);
and U11788 (N_11788,N_11592,N_11670);
xnor U11789 (N_11789,N_11628,N_11584);
nor U11790 (N_11790,N_11562,N_11678);
xor U11791 (N_11791,N_11594,N_11678);
xnor U11792 (N_11792,N_11633,N_11676);
and U11793 (N_11793,N_11657,N_11565);
nand U11794 (N_11794,N_11626,N_11597);
nor U11795 (N_11795,N_11644,N_11624);
nand U11796 (N_11796,N_11602,N_11676);
or U11797 (N_11797,N_11647,N_11676);
and U11798 (N_11798,N_11570,N_11576);
nor U11799 (N_11799,N_11691,N_11639);
xnor U11800 (N_11800,N_11635,N_11601);
and U11801 (N_11801,N_11551,N_11563);
or U11802 (N_11802,N_11554,N_11692);
and U11803 (N_11803,N_11565,N_11558);
and U11804 (N_11804,N_11632,N_11649);
xnor U11805 (N_11805,N_11687,N_11658);
xnor U11806 (N_11806,N_11625,N_11676);
xor U11807 (N_11807,N_11637,N_11663);
nand U11808 (N_11808,N_11591,N_11698);
nand U11809 (N_11809,N_11670,N_11558);
nand U11810 (N_11810,N_11571,N_11651);
nor U11811 (N_11811,N_11686,N_11564);
nor U11812 (N_11812,N_11550,N_11571);
nor U11813 (N_11813,N_11661,N_11629);
nand U11814 (N_11814,N_11583,N_11690);
nand U11815 (N_11815,N_11627,N_11647);
xor U11816 (N_11816,N_11624,N_11657);
xor U11817 (N_11817,N_11614,N_11551);
or U11818 (N_11818,N_11572,N_11678);
and U11819 (N_11819,N_11630,N_11632);
and U11820 (N_11820,N_11587,N_11624);
nand U11821 (N_11821,N_11684,N_11634);
and U11822 (N_11822,N_11565,N_11556);
nor U11823 (N_11823,N_11649,N_11573);
nor U11824 (N_11824,N_11612,N_11650);
xor U11825 (N_11825,N_11638,N_11633);
xor U11826 (N_11826,N_11561,N_11682);
or U11827 (N_11827,N_11559,N_11634);
or U11828 (N_11828,N_11664,N_11551);
xor U11829 (N_11829,N_11696,N_11586);
xnor U11830 (N_11830,N_11609,N_11573);
xor U11831 (N_11831,N_11687,N_11612);
nand U11832 (N_11832,N_11607,N_11656);
nand U11833 (N_11833,N_11646,N_11692);
xnor U11834 (N_11834,N_11638,N_11636);
and U11835 (N_11835,N_11576,N_11583);
or U11836 (N_11836,N_11615,N_11622);
nor U11837 (N_11837,N_11629,N_11591);
xnor U11838 (N_11838,N_11674,N_11551);
and U11839 (N_11839,N_11689,N_11622);
and U11840 (N_11840,N_11577,N_11632);
nor U11841 (N_11841,N_11566,N_11659);
or U11842 (N_11842,N_11636,N_11671);
nor U11843 (N_11843,N_11620,N_11642);
xor U11844 (N_11844,N_11674,N_11616);
nand U11845 (N_11845,N_11588,N_11603);
xnor U11846 (N_11846,N_11611,N_11660);
nor U11847 (N_11847,N_11670,N_11555);
xor U11848 (N_11848,N_11685,N_11567);
and U11849 (N_11849,N_11587,N_11572);
and U11850 (N_11850,N_11783,N_11740);
nand U11851 (N_11851,N_11793,N_11736);
and U11852 (N_11852,N_11755,N_11718);
nand U11853 (N_11853,N_11727,N_11819);
and U11854 (N_11854,N_11763,N_11708);
and U11855 (N_11855,N_11838,N_11807);
nor U11856 (N_11856,N_11753,N_11757);
and U11857 (N_11857,N_11713,N_11787);
and U11858 (N_11858,N_11833,N_11800);
xor U11859 (N_11859,N_11804,N_11811);
and U11860 (N_11860,N_11728,N_11743);
or U11861 (N_11861,N_11821,N_11704);
or U11862 (N_11862,N_11845,N_11817);
or U11863 (N_11863,N_11789,N_11762);
xor U11864 (N_11864,N_11812,N_11836);
nor U11865 (N_11865,N_11810,N_11813);
or U11866 (N_11866,N_11780,N_11831);
nand U11867 (N_11867,N_11742,N_11828);
xor U11868 (N_11868,N_11802,N_11825);
or U11869 (N_11869,N_11735,N_11798);
nor U11870 (N_11870,N_11722,N_11786);
nand U11871 (N_11871,N_11805,N_11771);
nand U11872 (N_11872,N_11705,N_11794);
nor U11873 (N_11873,N_11814,N_11826);
or U11874 (N_11874,N_11760,N_11806);
nand U11875 (N_11875,N_11772,N_11830);
nand U11876 (N_11876,N_11710,N_11840);
xor U11877 (N_11877,N_11792,N_11748);
nor U11878 (N_11878,N_11839,N_11779);
or U11879 (N_11879,N_11775,N_11732);
and U11880 (N_11880,N_11721,N_11774);
xor U11881 (N_11881,N_11818,N_11754);
and U11882 (N_11882,N_11797,N_11803);
xor U11883 (N_11883,N_11758,N_11752);
and U11884 (N_11884,N_11791,N_11824);
or U11885 (N_11885,N_11843,N_11730);
nor U11886 (N_11886,N_11846,N_11745);
or U11887 (N_11887,N_11799,N_11749);
or U11888 (N_11888,N_11820,N_11773);
nand U11889 (N_11889,N_11808,N_11747);
xor U11890 (N_11890,N_11734,N_11785);
nand U11891 (N_11891,N_11709,N_11823);
nor U11892 (N_11892,N_11790,N_11844);
and U11893 (N_11893,N_11795,N_11827);
xnor U11894 (N_11894,N_11767,N_11781);
nor U11895 (N_11895,N_11848,N_11724);
or U11896 (N_11896,N_11782,N_11822);
xnor U11897 (N_11897,N_11719,N_11741);
and U11898 (N_11898,N_11834,N_11744);
nor U11899 (N_11899,N_11725,N_11849);
or U11900 (N_11900,N_11738,N_11723);
nand U11901 (N_11901,N_11701,N_11715);
xnor U11902 (N_11902,N_11711,N_11770);
nor U11903 (N_11903,N_11768,N_11842);
and U11904 (N_11904,N_11769,N_11717);
nor U11905 (N_11905,N_11750,N_11816);
and U11906 (N_11906,N_11714,N_11796);
nand U11907 (N_11907,N_11777,N_11702);
nor U11908 (N_11908,N_11801,N_11739);
xor U11909 (N_11909,N_11815,N_11703);
or U11910 (N_11910,N_11764,N_11756);
or U11911 (N_11911,N_11832,N_11778);
xnor U11912 (N_11912,N_11784,N_11731);
xor U11913 (N_11913,N_11712,N_11729);
xor U11914 (N_11914,N_11837,N_11766);
xnor U11915 (N_11915,N_11776,N_11765);
and U11916 (N_11916,N_11847,N_11759);
or U11917 (N_11917,N_11726,N_11716);
and U11918 (N_11918,N_11700,N_11746);
xor U11919 (N_11919,N_11706,N_11707);
or U11920 (N_11920,N_11835,N_11761);
nor U11921 (N_11921,N_11829,N_11733);
nor U11922 (N_11922,N_11809,N_11788);
nor U11923 (N_11923,N_11737,N_11751);
and U11924 (N_11924,N_11841,N_11720);
nor U11925 (N_11925,N_11740,N_11830);
nand U11926 (N_11926,N_11840,N_11799);
xnor U11927 (N_11927,N_11735,N_11792);
or U11928 (N_11928,N_11821,N_11760);
and U11929 (N_11929,N_11791,N_11810);
xnor U11930 (N_11930,N_11725,N_11830);
or U11931 (N_11931,N_11778,N_11716);
or U11932 (N_11932,N_11829,N_11802);
nor U11933 (N_11933,N_11795,N_11714);
and U11934 (N_11934,N_11839,N_11721);
nor U11935 (N_11935,N_11733,N_11849);
xnor U11936 (N_11936,N_11761,N_11773);
xnor U11937 (N_11937,N_11804,N_11715);
xnor U11938 (N_11938,N_11792,N_11758);
nand U11939 (N_11939,N_11774,N_11819);
or U11940 (N_11940,N_11833,N_11728);
nand U11941 (N_11941,N_11810,N_11838);
nand U11942 (N_11942,N_11800,N_11771);
nand U11943 (N_11943,N_11703,N_11752);
or U11944 (N_11944,N_11712,N_11811);
and U11945 (N_11945,N_11764,N_11835);
and U11946 (N_11946,N_11720,N_11790);
and U11947 (N_11947,N_11727,N_11824);
nand U11948 (N_11948,N_11764,N_11791);
and U11949 (N_11949,N_11783,N_11799);
xnor U11950 (N_11950,N_11792,N_11788);
nor U11951 (N_11951,N_11809,N_11798);
nand U11952 (N_11952,N_11787,N_11719);
and U11953 (N_11953,N_11749,N_11794);
or U11954 (N_11954,N_11726,N_11770);
xnor U11955 (N_11955,N_11800,N_11701);
and U11956 (N_11956,N_11841,N_11721);
or U11957 (N_11957,N_11822,N_11753);
nor U11958 (N_11958,N_11733,N_11724);
xnor U11959 (N_11959,N_11846,N_11821);
xor U11960 (N_11960,N_11753,N_11800);
nor U11961 (N_11961,N_11838,N_11738);
nor U11962 (N_11962,N_11701,N_11739);
xor U11963 (N_11963,N_11813,N_11828);
or U11964 (N_11964,N_11774,N_11812);
or U11965 (N_11965,N_11734,N_11732);
xor U11966 (N_11966,N_11739,N_11711);
and U11967 (N_11967,N_11711,N_11805);
nand U11968 (N_11968,N_11827,N_11822);
or U11969 (N_11969,N_11814,N_11743);
nor U11970 (N_11970,N_11755,N_11733);
or U11971 (N_11971,N_11765,N_11799);
nand U11972 (N_11972,N_11759,N_11755);
or U11973 (N_11973,N_11734,N_11779);
or U11974 (N_11974,N_11776,N_11794);
nand U11975 (N_11975,N_11751,N_11707);
xnor U11976 (N_11976,N_11761,N_11775);
and U11977 (N_11977,N_11806,N_11773);
or U11978 (N_11978,N_11735,N_11826);
nand U11979 (N_11979,N_11789,N_11721);
xor U11980 (N_11980,N_11754,N_11712);
and U11981 (N_11981,N_11807,N_11713);
or U11982 (N_11982,N_11837,N_11844);
nand U11983 (N_11983,N_11767,N_11814);
or U11984 (N_11984,N_11777,N_11787);
nor U11985 (N_11985,N_11743,N_11830);
or U11986 (N_11986,N_11823,N_11797);
nor U11987 (N_11987,N_11796,N_11845);
nand U11988 (N_11988,N_11746,N_11844);
or U11989 (N_11989,N_11705,N_11830);
and U11990 (N_11990,N_11741,N_11776);
nor U11991 (N_11991,N_11704,N_11838);
xor U11992 (N_11992,N_11721,N_11833);
nor U11993 (N_11993,N_11717,N_11765);
nand U11994 (N_11994,N_11742,N_11780);
xnor U11995 (N_11995,N_11743,N_11794);
and U11996 (N_11996,N_11718,N_11776);
nor U11997 (N_11997,N_11742,N_11787);
nor U11998 (N_11998,N_11705,N_11729);
or U11999 (N_11999,N_11837,N_11748);
or U12000 (N_12000,N_11863,N_11943);
nor U12001 (N_12001,N_11897,N_11945);
xor U12002 (N_12002,N_11974,N_11856);
nand U12003 (N_12003,N_11902,N_11916);
and U12004 (N_12004,N_11870,N_11875);
nand U12005 (N_12005,N_11930,N_11978);
nand U12006 (N_12006,N_11862,N_11927);
nor U12007 (N_12007,N_11877,N_11932);
and U12008 (N_12008,N_11938,N_11882);
xnor U12009 (N_12009,N_11979,N_11933);
or U12010 (N_12010,N_11941,N_11861);
xnor U12011 (N_12011,N_11908,N_11967);
nor U12012 (N_12012,N_11984,N_11859);
and U12013 (N_12013,N_11850,N_11998);
and U12014 (N_12014,N_11851,N_11940);
xor U12015 (N_12015,N_11963,N_11993);
and U12016 (N_12016,N_11890,N_11985);
nor U12017 (N_12017,N_11924,N_11950);
or U12018 (N_12018,N_11868,N_11899);
xor U12019 (N_12019,N_11855,N_11910);
or U12020 (N_12020,N_11860,N_11905);
nand U12021 (N_12021,N_11946,N_11925);
nor U12022 (N_12022,N_11891,N_11997);
and U12023 (N_12023,N_11878,N_11903);
or U12024 (N_12024,N_11951,N_11895);
nor U12025 (N_12025,N_11919,N_11907);
and U12026 (N_12026,N_11922,N_11889);
and U12027 (N_12027,N_11957,N_11992);
and U12028 (N_12028,N_11964,N_11944);
nand U12029 (N_12029,N_11883,N_11947);
xnor U12030 (N_12030,N_11935,N_11937);
and U12031 (N_12031,N_11880,N_11975);
xor U12032 (N_12032,N_11952,N_11898);
nor U12033 (N_12033,N_11896,N_11983);
xnor U12034 (N_12034,N_11921,N_11972);
xnor U12035 (N_12035,N_11973,N_11965);
nor U12036 (N_12036,N_11876,N_11961);
and U12037 (N_12037,N_11887,N_11929);
xor U12038 (N_12038,N_11981,N_11864);
nor U12039 (N_12039,N_11962,N_11857);
or U12040 (N_12040,N_11867,N_11865);
or U12041 (N_12041,N_11912,N_11956);
xor U12042 (N_12042,N_11915,N_11980);
nand U12043 (N_12043,N_11988,N_11904);
nor U12044 (N_12044,N_11999,N_11881);
nor U12045 (N_12045,N_11958,N_11953);
nand U12046 (N_12046,N_11900,N_11936);
and U12047 (N_12047,N_11968,N_11971);
nor U12048 (N_12048,N_11989,N_11885);
nor U12049 (N_12049,N_11913,N_11942);
and U12050 (N_12050,N_11954,N_11852);
nor U12051 (N_12051,N_11892,N_11966);
and U12052 (N_12052,N_11911,N_11872);
nand U12053 (N_12053,N_11982,N_11931);
or U12054 (N_12054,N_11869,N_11884);
and U12055 (N_12055,N_11894,N_11879);
xor U12056 (N_12056,N_11990,N_11996);
nand U12057 (N_12057,N_11901,N_11969);
nor U12058 (N_12058,N_11888,N_11960);
and U12059 (N_12059,N_11955,N_11918);
or U12060 (N_12060,N_11854,N_11926);
or U12061 (N_12061,N_11948,N_11920);
or U12062 (N_12062,N_11906,N_11987);
nor U12063 (N_12063,N_11871,N_11928);
or U12064 (N_12064,N_11853,N_11917);
nand U12065 (N_12065,N_11893,N_11909);
xor U12066 (N_12066,N_11995,N_11977);
or U12067 (N_12067,N_11934,N_11873);
and U12068 (N_12068,N_11959,N_11886);
nand U12069 (N_12069,N_11923,N_11914);
or U12070 (N_12070,N_11976,N_11970);
or U12071 (N_12071,N_11994,N_11986);
and U12072 (N_12072,N_11939,N_11991);
xor U12073 (N_12073,N_11874,N_11949);
nand U12074 (N_12074,N_11866,N_11858);
nand U12075 (N_12075,N_11862,N_11994);
nor U12076 (N_12076,N_11946,N_11904);
xor U12077 (N_12077,N_11959,N_11869);
and U12078 (N_12078,N_11859,N_11971);
nor U12079 (N_12079,N_11965,N_11866);
nor U12080 (N_12080,N_11916,N_11904);
xnor U12081 (N_12081,N_11923,N_11892);
and U12082 (N_12082,N_11964,N_11903);
and U12083 (N_12083,N_11981,N_11986);
or U12084 (N_12084,N_11964,N_11993);
nand U12085 (N_12085,N_11864,N_11892);
nand U12086 (N_12086,N_11920,N_11983);
or U12087 (N_12087,N_11876,N_11935);
or U12088 (N_12088,N_11976,N_11916);
or U12089 (N_12089,N_11900,N_11962);
or U12090 (N_12090,N_11953,N_11929);
nor U12091 (N_12091,N_11905,N_11945);
and U12092 (N_12092,N_11859,N_11882);
and U12093 (N_12093,N_11929,N_11987);
or U12094 (N_12094,N_11930,N_11961);
nand U12095 (N_12095,N_11883,N_11914);
nand U12096 (N_12096,N_11885,N_11937);
nor U12097 (N_12097,N_11978,N_11944);
xnor U12098 (N_12098,N_11888,N_11947);
nand U12099 (N_12099,N_11938,N_11936);
or U12100 (N_12100,N_11914,N_11905);
or U12101 (N_12101,N_11865,N_11905);
or U12102 (N_12102,N_11906,N_11852);
and U12103 (N_12103,N_11883,N_11993);
and U12104 (N_12104,N_11984,N_11855);
xnor U12105 (N_12105,N_11936,N_11976);
and U12106 (N_12106,N_11856,N_11984);
xnor U12107 (N_12107,N_11996,N_11872);
nor U12108 (N_12108,N_11940,N_11911);
nor U12109 (N_12109,N_11915,N_11865);
nor U12110 (N_12110,N_11957,N_11892);
and U12111 (N_12111,N_11979,N_11989);
and U12112 (N_12112,N_11997,N_11863);
or U12113 (N_12113,N_11934,N_11975);
nand U12114 (N_12114,N_11933,N_11988);
and U12115 (N_12115,N_11887,N_11944);
and U12116 (N_12116,N_11886,N_11938);
nor U12117 (N_12117,N_11856,N_11852);
xor U12118 (N_12118,N_11867,N_11949);
nand U12119 (N_12119,N_11949,N_11972);
and U12120 (N_12120,N_11903,N_11869);
nor U12121 (N_12121,N_11910,N_11922);
and U12122 (N_12122,N_11912,N_11921);
or U12123 (N_12123,N_11851,N_11890);
xnor U12124 (N_12124,N_11925,N_11920);
nor U12125 (N_12125,N_11933,N_11986);
nand U12126 (N_12126,N_11894,N_11937);
or U12127 (N_12127,N_11860,N_11984);
xnor U12128 (N_12128,N_11977,N_11932);
or U12129 (N_12129,N_11873,N_11865);
nor U12130 (N_12130,N_11910,N_11885);
and U12131 (N_12131,N_11868,N_11983);
or U12132 (N_12132,N_11910,N_11958);
nand U12133 (N_12133,N_11970,N_11887);
or U12134 (N_12134,N_11976,N_11886);
xnor U12135 (N_12135,N_11978,N_11851);
xnor U12136 (N_12136,N_11877,N_11938);
and U12137 (N_12137,N_11871,N_11988);
or U12138 (N_12138,N_11917,N_11971);
nand U12139 (N_12139,N_11936,N_11884);
nor U12140 (N_12140,N_11974,N_11865);
nand U12141 (N_12141,N_11966,N_11908);
xnor U12142 (N_12142,N_11908,N_11863);
and U12143 (N_12143,N_11979,N_11929);
nor U12144 (N_12144,N_11852,N_11908);
nor U12145 (N_12145,N_11946,N_11927);
nand U12146 (N_12146,N_11959,N_11926);
xor U12147 (N_12147,N_11976,N_11910);
nor U12148 (N_12148,N_11901,N_11995);
xor U12149 (N_12149,N_11935,N_11901);
nand U12150 (N_12150,N_12043,N_12007);
xnor U12151 (N_12151,N_12035,N_12044);
or U12152 (N_12152,N_12080,N_12112);
and U12153 (N_12153,N_12034,N_12074);
or U12154 (N_12154,N_12060,N_12086);
nor U12155 (N_12155,N_12076,N_12103);
xor U12156 (N_12156,N_12017,N_12135);
xnor U12157 (N_12157,N_12097,N_12016);
nand U12158 (N_12158,N_12115,N_12118);
nand U12159 (N_12159,N_12029,N_12079);
and U12160 (N_12160,N_12039,N_12126);
nand U12161 (N_12161,N_12058,N_12005);
xnor U12162 (N_12162,N_12063,N_12041);
nor U12163 (N_12163,N_12095,N_12089);
or U12164 (N_12164,N_12025,N_12067);
nand U12165 (N_12165,N_12010,N_12072);
nor U12166 (N_12166,N_12140,N_12062);
or U12167 (N_12167,N_12141,N_12116);
and U12168 (N_12168,N_12053,N_12093);
nand U12169 (N_12169,N_12091,N_12096);
nand U12170 (N_12170,N_12134,N_12106);
nand U12171 (N_12171,N_12014,N_12136);
or U12172 (N_12172,N_12033,N_12050);
xnor U12173 (N_12173,N_12143,N_12018);
nand U12174 (N_12174,N_12087,N_12139);
xor U12175 (N_12175,N_12069,N_12123);
nor U12176 (N_12176,N_12068,N_12142);
and U12177 (N_12177,N_12037,N_12065);
xor U12178 (N_12178,N_12040,N_12026);
xnor U12179 (N_12179,N_12008,N_12031);
and U12180 (N_12180,N_12090,N_12022);
nor U12181 (N_12181,N_12082,N_12149);
xnor U12182 (N_12182,N_12094,N_12104);
and U12183 (N_12183,N_12003,N_12110);
xor U12184 (N_12184,N_12015,N_12111);
nor U12185 (N_12185,N_12049,N_12070);
nand U12186 (N_12186,N_12059,N_12131);
or U12187 (N_12187,N_12020,N_12001);
nand U12188 (N_12188,N_12052,N_12145);
nand U12189 (N_12189,N_12119,N_12028);
and U12190 (N_12190,N_12024,N_12004);
xor U12191 (N_12191,N_12114,N_12121);
nand U12192 (N_12192,N_12066,N_12137);
xnor U12193 (N_12193,N_12099,N_12085);
and U12194 (N_12194,N_12147,N_12113);
nand U12195 (N_12195,N_12000,N_12073);
nor U12196 (N_12196,N_12100,N_12105);
or U12197 (N_12197,N_12042,N_12027);
and U12198 (N_12198,N_12101,N_12146);
nand U12199 (N_12199,N_12045,N_12083);
or U12200 (N_12200,N_12002,N_12038);
nor U12201 (N_12201,N_12081,N_12102);
and U12202 (N_12202,N_12012,N_12036);
nand U12203 (N_12203,N_12117,N_12075);
and U12204 (N_12204,N_12127,N_12011);
and U12205 (N_12205,N_12108,N_12109);
nor U12206 (N_12206,N_12148,N_12046);
nor U12207 (N_12207,N_12084,N_12032);
nand U12208 (N_12208,N_12061,N_12051);
nor U12209 (N_12209,N_12009,N_12056);
xnor U12210 (N_12210,N_12130,N_12092);
or U12211 (N_12211,N_12088,N_12124);
nand U12212 (N_12212,N_12013,N_12078);
xnor U12213 (N_12213,N_12071,N_12138);
and U12214 (N_12214,N_12098,N_12144);
nor U12215 (N_12215,N_12129,N_12133);
nor U12216 (N_12216,N_12077,N_12023);
and U12217 (N_12217,N_12047,N_12054);
nand U12218 (N_12218,N_12019,N_12122);
or U12219 (N_12219,N_12048,N_12030);
and U12220 (N_12220,N_12055,N_12107);
or U12221 (N_12221,N_12125,N_12057);
or U12222 (N_12222,N_12128,N_12006);
nand U12223 (N_12223,N_12132,N_12021);
nand U12224 (N_12224,N_12064,N_12120);
xnor U12225 (N_12225,N_12144,N_12064);
nor U12226 (N_12226,N_12111,N_12000);
xnor U12227 (N_12227,N_12066,N_12023);
nand U12228 (N_12228,N_12029,N_12110);
or U12229 (N_12229,N_12087,N_12147);
and U12230 (N_12230,N_12062,N_12063);
xor U12231 (N_12231,N_12019,N_12042);
nand U12232 (N_12232,N_12100,N_12145);
nand U12233 (N_12233,N_12021,N_12097);
nand U12234 (N_12234,N_12115,N_12129);
nand U12235 (N_12235,N_12062,N_12020);
and U12236 (N_12236,N_12043,N_12041);
xor U12237 (N_12237,N_12035,N_12068);
nand U12238 (N_12238,N_12012,N_12066);
xor U12239 (N_12239,N_12089,N_12015);
and U12240 (N_12240,N_12087,N_12004);
or U12241 (N_12241,N_12041,N_12016);
nand U12242 (N_12242,N_12044,N_12104);
nor U12243 (N_12243,N_12060,N_12034);
and U12244 (N_12244,N_12119,N_12105);
nor U12245 (N_12245,N_12137,N_12050);
or U12246 (N_12246,N_12015,N_12047);
nand U12247 (N_12247,N_12103,N_12016);
nor U12248 (N_12248,N_12023,N_12102);
nor U12249 (N_12249,N_12134,N_12096);
or U12250 (N_12250,N_12072,N_12009);
nand U12251 (N_12251,N_12110,N_12147);
nor U12252 (N_12252,N_12023,N_12116);
xor U12253 (N_12253,N_12096,N_12113);
and U12254 (N_12254,N_12117,N_12092);
or U12255 (N_12255,N_12071,N_12146);
nor U12256 (N_12256,N_12120,N_12079);
and U12257 (N_12257,N_12049,N_12041);
or U12258 (N_12258,N_12018,N_12047);
nand U12259 (N_12259,N_12007,N_12033);
and U12260 (N_12260,N_12003,N_12011);
nor U12261 (N_12261,N_12003,N_12052);
or U12262 (N_12262,N_12128,N_12111);
and U12263 (N_12263,N_12129,N_12096);
nor U12264 (N_12264,N_12094,N_12006);
and U12265 (N_12265,N_12115,N_12108);
or U12266 (N_12266,N_12137,N_12128);
nand U12267 (N_12267,N_12111,N_12102);
xor U12268 (N_12268,N_12033,N_12085);
or U12269 (N_12269,N_12004,N_12076);
nand U12270 (N_12270,N_12056,N_12015);
or U12271 (N_12271,N_12064,N_12076);
xor U12272 (N_12272,N_12033,N_12077);
nor U12273 (N_12273,N_12122,N_12069);
nand U12274 (N_12274,N_12019,N_12045);
xor U12275 (N_12275,N_12141,N_12124);
or U12276 (N_12276,N_12050,N_12078);
nor U12277 (N_12277,N_12077,N_12047);
xor U12278 (N_12278,N_12055,N_12038);
xor U12279 (N_12279,N_12037,N_12118);
or U12280 (N_12280,N_12044,N_12026);
and U12281 (N_12281,N_12124,N_12043);
or U12282 (N_12282,N_12133,N_12143);
nor U12283 (N_12283,N_12127,N_12122);
nor U12284 (N_12284,N_12145,N_12116);
nand U12285 (N_12285,N_12007,N_12054);
and U12286 (N_12286,N_12072,N_12074);
nand U12287 (N_12287,N_12095,N_12146);
nand U12288 (N_12288,N_12008,N_12026);
or U12289 (N_12289,N_12050,N_12060);
nand U12290 (N_12290,N_12027,N_12064);
nor U12291 (N_12291,N_12075,N_12001);
nor U12292 (N_12292,N_12127,N_12078);
nand U12293 (N_12293,N_12023,N_12030);
and U12294 (N_12294,N_12108,N_12003);
nor U12295 (N_12295,N_12030,N_12138);
nor U12296 (N_12296,N_12142,N_12111);
nand U12297 (N_12297,N_12031,N_12083);
xnor U12298 (N_12298,N_12147,N_12131);
and U12299 (N_12299,N_12043,N_12115);
nand U12300 (N_12300,N_12235,N_12245);
nor U12301 (N_12301,N_12231,N_12298);
or U12302 (N_12302,N_12153,N_12188);
and U12303 (N_12303,N_12175,N_12198);
xnor U12304 (N_12304,N_12196,N_12226);
xnor U12305 (N_12305,N_12274,N_12209);
or U12306 (N_12306,N_12189,N_12272);
xnor U12307 (N_12307,N_12238,N_12240);
and U12308 (N_12308,N_12178,N_12160);
and U12309 (N_12309,N_12225,N_12150);
or U12310 (N_12310,N_12215,N_12244);
nor U12311 (N_12311,N_12254,N_12218);
nand U12312 (N_12312,N_12193,N_12260);
nor U12313 (N_12313,N_12159,N_12294);
xor U12314 (N_12314,N_12182,N_12234);
xnor U12315 (N_12315,N_12230,N_12284);
nand U12316 (N_12316,N_12291,N_12280);
and U12317 (N_12317,N_12247,N_12184);
and U12318 (N_12318,N_12216,N_12293);
xor U12319 (N_12319,N_12210,N_12236);
xnor U12320 (N_12320,N_12166,N_12192);
nand U12321 (N_12321,N_12268,N_12269);
and U12322 (N_12322,N_12157,N_12264);
xnor U12323 (N_12323,N_12287,N_12176);
xor U12324 (N_12324,N_12194,N_12233);
nand U12325 (N_12325,N_12241,N_12282);
or U12326 (N_12326,N_12250,N_12161);
or U12327 (N_12327,N_12278,N_12168);
and U12328 (N_12328,N_12248,N_12259);
or U12329 (N_12329,N_12249,N_12286);
or U12330 (N_12330,N_12190,N_12199);
and U12331 (N_12331,N_12202,N_12219);
nor U12332 (N_12332,N_12223,N_12285);
xnor U12333 (N_12333,N_12296,N_12201);
or U12334 (N_12334,N_12173,N_12265);
xor U12335 (N_12335,N_12256,N_12297);
nor U12336 (N_12336,N_12222,N_12261);
nand U12337 (N_12337,N_12191,N_12180);
nor U12338 (N_12338,N_12271,N_12299);
nor U12339 (N_12339,N_12203,N_12243);
and U12340 (N_12340,N_12151,N_12162);
nand U12341 (N_12341,N_12276,N_12174);
xnor U12342 (N_12342,N_12266,N_12187);
xor U12343 (N_12343,N_12185,N_12267);
nor U12344 (N_12344,N_12273,N_12205);
and U12345 (N_12345,N_12224,N_12262);
xor U12346 (N_12346,N_12169,N_12212);
or U12347 (N_12347,N_12181,N_12195);
nand U12348 (N_12348,N_12227,N_12255);
nor U12349 (N_12349,N_12186,N_12295);
nor U12350 (N_12350,N_12179,N_12211);
or U12351 (N_12351,N_12213,N_12155);
or U12352 (N_12352,N_12251,N_12163);
xor U12353 (N_12353,N_12239,N_12228);
and U12354 (N_12354,N_12171,N_12242);
xor U12355 (N_12355,N_12279,N_12208);
or U12356 (N_12356,N_12229,N_12172);
xor U12357 (N_12357,N_12288,N_12167);
nor U12358 (N_12358,N_12152,N_12170);
nor U12359 (N_12359,N_12237,N_12207);
nor U12360 (N_12360,N_12290,N_12164);
nor U12361 (N_12361,N_12220,N_12204);
nor U12362 (N_12362,N_12270,N_12200);
and U12363 (N_12363,N_12206,N_12158);
xnor U12364 (N_12364,N_12283,N_12281);
nand U12365 (N_12365,N_12292,N_12253);
nand U12366 (N_12366,N_12197,N_12183);
xnor U12367 (N_12367,N_12214,N_12232);
and U12368 (N_12368,N_12258,N_12217);
and U12369 (N_12369,N_12221,N_12246);
nand U12370 (N_12370,N_12263,N_12177);
nand U12371 (N_12371,N_12156,N_12257);
and U12372 (N_12372,N_12252,N_12277);
xnor U12373 (N_12373,N_12165,N_12289);
xnor U12374 (N_12374,N_12154,N_12275);
and U12375 (N_12375,N_12228,N_12182);
nand U12376 (N_12376,N_12173,N_12275);
or U12377 (N_12377,N_12281,N_12182);
nand U12378 (N_12378,N_12210,N_12280);
nand U12379 (N_12379,N_12179,N_12270);
or U12380 (N_12380,N_12240,N_12152);
xnor U12381 (N_12381,N_12271,N_12188);
xor U12382 (N_12382,N_12220,N_12286);
nand U12383 (N_12383,N_12252,N_12267);
or U12384 (N_12384,N_12163,N_12257);
or U12385 (N_12385,N_12189,N_12198);
or U12386 (N_12386,N_12205,N_12270);
and U12387 (N_12387,N_12156,N_12220);
nand U12388 (N_12388,N_12233,N_12242);
xnor U12389 (N_12389,N_12254,N_12157);
and U12390 (N_12390,N_12205,N_12199);
nor U12391 (N_12391,N_12269,N_12204);
xor U12392 (N_12392,N_12242,N_12267);
and U12393 (N_12393,N_12173,N_12289);
nand U12394 (N_12394,N_12221,N_12282);
or U12395 (N_12395,N_12163,N_12247);
and U12396 (N_12396,N_12208,N_12291);
and U12397 (N_12397,N_12186,N_12176);
and U12398 (N_12398,N_12272,N_12255);
nand U12399 (N_12399,N_12262,N_12230);
nand U12400 (N_12400,N_12212,N_12156);
nor U12401 (N_12401,N_12270,N_12154);
nor U12402 (N_12402,N_12278,N_12250);
nand U12403 (N_12403,N_12158,N_12182);
xnor U12404 (N_12404,N_12280,N_12188);
or U12405 (N_12405,N_12158,N_12280);
xor U12406 (N_12406,N_12201,N_12274);
and U12407 (N_12407,N_12279,N_12250);
nor U12408 (N_12408,N_12296,N_12262);
or U12409 (N_12409,N_12223,N_12220);
or U12410 (N_12410,N_12221,N_12228);
nor U12411 (N_12411,N_12183,N_12160);
nand U12412 (N_12412,N_12276,N_12258);
and U12413 (N_12413,N_12181,N_12200);
nand U12414 (N_12414,N_12177,N_12236);
or U12415 (N_12415,N_12170,N_12281);
xnor U12416 (N_12416,N_12204,N_12196);
and U12417 (N_12417,N_12201,N_12276);
or U12418 (N_12418,N_12205,N_12229);
xor U12419 (N_12419,N_12152,N_12282);
or U12420 (N_12420,N_12292,N_12236);
xnor U12421 (N_12421,N_12227,N_12203);
and U12422 (N_12422,N_12291,N_12244);
nor U12423 (N_12423,N_12231,N_12195);
and U12424 (N_12424,N_12153,N_12263);
and U12425 (N_12425,N_12175,N_12158);
nor U12426 (N_12426,N_12170,N_12268);
and U12427 (N_12427,N_12212,N_12267);
xnor U12428 (N_12428,N_12191,N_12266);
or U12429 (N_12429,N_12205,N_12178);
xnor U12430 (N_12430,N_12161,N_12286);
nor U12431 (N_12431,N_12176,N_12254);
or U12432 (N_12432,N_12161,N_12154);
or U12433 (N_12433,N_12157,N_12261);
and U12434 (N_12434,N_12275,N_12270);
nor U12435 (N_12435,N_12210,N_12260);
and U12436 (N_12436,N_12174,N_12199);
or U12437 (N_12437,N_12197,N_12278);
or U12438 (N_12438,N_12272,N_12214);
xnor U12439 (N_12439,N_12226,N_12289);
nand U12440 (N_12440,N_12210,N_12187);
and U12441 (N_12441,N_12152,N_12286);
or U12442 (N_12442,N_12159,N_12185);
xnor U12443 (N_12443,N_12246,N_12178);
or U12444 (N_12444,N_12253,N_12268);
nand U12445 (N_12445,N_12187,N_12180);
and U12446 (N_12446,N_12203,N_12220);
and U12447 (N_12447,N_12203,N_12154);
nand U12448 (N_12448,N_12263,N_12199);
nor U12449 (N_12449,N_12181,N_12222);
xnor U12450 (N_12450,N_12372,N_12316);
nor U12451 (N_12451,N_12318,N_12362);
nand U12452 (N_12452,N_12449,N_12445);
xnor U12453 (N_12453,N_12350,N_12309);
or U12454 (N_12454,N_12305,N_12345);
and U12455 (N_12455,N_12442,N_12327);
and U12456 (N_12456,N_12341,N_12402);
and U12457 (N_12457,N_12412,N_12404);
xor U12458 (N_12458,N_12375,N_12423);
or U12459 (N_12459,N_12340,N_12302);
xnor U12460 (N_12460,N_12430,N_12414);
nor U12461 (N_12461,N_12419,N_12417);
and U12462 (N_12462,N_12320,N_12334);
xor U12463 (N_12463,N_12398,N_12317);
or U12464 (N_12464,N_12343,N_12371);
nor U12465 (N_12465,N_12310,N_12360);
and U12466 (N_12466,N_12313,N_12365);
nand U12467 (N_12467,N_12324,N_12429);
xnor U12468 (N_12468,N_12407,N_12377);
and U12469 (N_12469,N_12331,N_12357);
nor U12470 (N_12470,N_12363,N_12380);
or U12471 (N_12471,N_12431,N_12439);
or U12472 (N_12472,N_12415,N_12426);
or U12473 (N_12473,N_12373,N_12386);
nand U12474 (N_12474,N_12403,N_12444);
nor U12475 (N_12475,N_12322,N_12387);
nand U12476 (N_12476,N_12356,N_12338);
xor U12477 (N_12477,N_12358,N_12370);
and U12478 (N_12478,N_12353,N_12332);
nand U12479 (N_12479,N_12443,N_12409);
or U12480 (N_12480,N_12384,N_12308);
nand U12481 (N_12481,N_12441,N_12383);
nor U12482 (N_12482,N_12311,N_12300);
nor U12483 (N_12483,N_12382,N_12389);
and U12484 (N_12484,N_12411,N_12348);
or U12485 (N_12485,N_12319,N_12399);
nand U12486 (N_12486,N_12351,N_12440);
nor U12487 (N_12487,N_12446,N_12397);
nor U12488 (N_12488,N_12368,N_12413);
or U12489 (N_12489,N_12347,N_12421);
and U12490 (N_12490,N_12364,N_12378);
nor U12491 (N_12491,N_12395,N_12391);
xnor U12492 (N_12492,N_12333,N_12447);
or U12493 (N_12493,N_12436,N_12361);
and U12494 (N_12494,N_12418,N_12428);
and U12495 (N_12495,N_12304,N_12315);
and U12496 (N_12496,N_12307,N_12335);
or U12497 (N_12497,N_12337,N_12306);
nand U12498 (N_12498,N_12406,N_12381);
and U12499 (N_12499,N_12420,N_12374);
xnor U12500 (N_12500,N_12435,N_12354);
or U12501 (N_12501,N_12432,N_12339);
nor U12502 (N_12502,N_12388,N_12367);
and U12503 (N_12503,N_12416,N_12408);
nand U12504 (N_12504,N_12410,N_12314);
or U12505 (N_12505,N_12385,N_12400);
xnor U12506 (N_12506,N_12344,N_12326);
xor U12507 (N_12507,N_12325,N_12425);
and U12508 (N_12508,N_12392,N_12369);
nand U12509 (N_12509,N_12437,N_12303);
nand U12510 (N_12510,N_12438,N_12396);
nor U12511 (N_12511,N_12366,N_12330);
xnor U12512 (N_12512,N_12376,N_12329);
and U12513 (N_12513,N_12355,N_12312);
and U12514 (N_12514,N_12352,N_12328);
and U12515 (N_12515,N_12390,N_12301);
and U12516 (N_12516,N_12433,N_12427);
or U12517 (N_12517,N_12346,N_12405);
and U12518 (N_12518,N_12349,N_12321);
and U12519 (N_12519,N_12323,N_12424);
or U12520 (N_12520,N_12336,N_12379);
and U12521 (N_12521,N_12401,N_12448);
nor U12522 (N_12522,N_12394,N_12393);
xor U12523 (N_12523,N_12422,N_12359);
xor U12524 (N_12524,N_12342,N_12434);
xnor U12525 (N_12525,N_12411,N_12438);
or U12526 (N_12526,N_12405,N_12314);
or U12527 (N_12527,N_12440,N_12372);
nand U12528 (N_12528,N_12419,N_12333);
nand U12529 (N_12529,N_12400,N_12379);
xnor U12530 (N_12530,N_12330,N_12308);
nor U12531 (N_12531,N_12360,N_12313);
xnor U12532 (N_12532,N_12391,N_12304);
nor U12533 (N_12533,N_12392,N_12413);
and U12534 (N_12534,N_12317,N_12336);
or U12535 (N_12535,N_12357,N_12339);
nand U12536 (N_12536,N_12405,N_12333);
nor U12537 (N_12537,N_12427,N_12435);
and U12538 (N_12538,N_12376,N_12351);
and U12539 (N_12539,N_12355,N_12415);
and U12540 (N_12540,N_12341,N_12336);
xor U12541 (N_12541,N_12404,N_12428);
xor U12542 (N_12542,N_12317,N_12444);
and U12543 (N_12543,N_12352,N_12432);
nand U12544 (N_12544,N_12306,N_12402);
and U12545 (N_12545,N_12405,N_12356);
or U12546 (N_12546,N_12425,N_12318);
and U12547 (N_12547,N_12418,N_12311);
nand U12548 (N_12548,N_12396,N_12371);
or U12549 (N_12549,N_12347,N_12378);
or U12550 (N_12550,N_12350,N_12433);
or U12551 (N_12551,N_12375,N_12368);
or U12552 (N_12552,N_12357,N_12428);
and U12553 (N_12553,N_12435,N_12325);
or U12554 (N_12554,N_12446,N_12316);
xor U12555 (N_12555,N_12327,N_12415);
nor U12556 (N_12556,N_12344,N_12447);
nor U12557 (N_12557,N_12339,N_12364);
nor U12558 (N_12558,N_12432,N_12408);
nor U12559 (N_12559,N_12320,N_12326);
and U12560 (N_12560,N_12418,N_12434);
xor U12561 (N_12561,N_12366,N_12407);
xor U12562 (N_12562,N_12331,N_12392);
nand U12563 (N_12563,N_12402,N_12323);
xor U12564 (N_12564,N_12426,N_12432);
nand U12565 (N_12565,N_12384,N_12316);
and U12566 (N_12566,N_12351,N_12410);
nor U12567 (N_12567,N_12393,N_12408);
xor U12568 (N_12568,N_12326,N_12423);
xor U12569 (N_12569,N_12417,N_12347);
xor U12570 (N_12570,N_12381,N_12389);
xnor U12571 (N_12571,N_12424,N_12358);
and U12572 (N_12572,N_12324,N_12340);
or U12573 (N_12573,N_12353,N_12419);
nand U12574 (N_12574,N_12368,N_12328);
xnor U12575 (N_12575,N_12325,N_12379);
xnor U12576 (N_12576,N_12319,N_12305);
nand U12577 (N_12577,N_12313,N_12301);
nand U12578 (N_12578,N_12396,N_12398);
nor U12579 (N_12579,N_12437,N_12352);
or U12580 (N_12580,N_12424,N_12446);
and U12581 (N_12581,N_12340,N_12320);
or U12582 (N_12582,N_12343,N_12366);
or U12583 (N_12583,N_12309,N_12420);
and U12584 (N_12584,N_12430,N_12352);
nor U12585 (N_12585,N_12363,N_12301);
nor U12586 (N_12586,N_12390,N_12345);
and U12587 (N_12587,N_12305,N_12382);
and U12588 (N_12588,N_12378,N_12374);
xor U12589 (N_12589,N_12417,N_12311);
and U12590 (N_12590,N_12358,N_12342);
xor U12591 (N_12591,N_12309,N_12417);
and U12592 (N_12592,N_12336,N_12373);
and U12593 (N_12593,N_12418,N_12372);
nor U12594 (N_12594,N_12320,N_12408);
and U12595 (N_12595,N_12414,N_12357);
and U12596 (N_12596,N_12311,N_12349);
nor U12597 (N_12597,N_12391,N_12445);
nor U12598 (N_12598,N_12353,N_12391);
xnor U12599 (N_12599,N_12320,N_12435);
or U12600 (N_12600,N_12589,N_12527);
and U12601 (N_12601,N_12514,N_12522);
nand U12602 (N_12602,N_12466,N_12565);
and U12603 (N_12603,N_12562,N_12557);
xnor U12604 (N_12604,N_12517,N_12505);
xnor U12605 (N_12605,N_12460,N_12454);
or U12606 (N_12606,N_12474,N_12516);
nor U12607 (N_12607,N_12596,N_12475);
or U12608 (N_12608,N_12591,N_12546);
xnor U12609 (N_12609,N_12551,N_12552);
xor U12610 (N_12610,N_12497,N_12478);
and U12611 (N_12611,N_12467,N_12571);
nand U12612 (N_12612,N_12508,N_12566);
nor U12613 (N_12613,N_12510,N_12587);
xor U12614 (N_12614,N_12494,N_12493);
or U12615 (N_12615,N_12461,N_12553);
nor U12616 (N_12616,N_12483,N_12468);
nand U12617 (N_12617,N_12583,N_12463);
or U12618 (N_12618,N_12568,N_12585);
nand U12619 (N_12619,N_12532,N_12530);
nor U12620 (N_12620,N_12543,N_12567);
nand U12621 (N_12621,N_12534,N_12520);
nor U12622 (N_12622,N_12599,N_12536);
or U12623 (N_12623,N_12485,N_12561);
xnor U12624 (N_12624,N_12537,N_12488);
and U12625 (N_12625,N_12594,N_12515);
and U12626 (N_12626,N_12503,N_12570);
nor U12627 (N_12627,N_12542,N_12577);
and U12628 (N_12628,N_12453,N_12593);
and U12629 (N_12629,N_12555,N_12554);
or U12630 (N_12630,N_12579,N_12486);
and U12631 (N_12631,N_12506,N_12465);
xor U12632 (N_12632,N_12592,N_12482);
or U12633 (N_12633,N_12524,N_12495);
nor U12634 (N_12634,N_12531,N_12451);
or U12635 (N_12635,N_12575,N_12450);
xor U12636 (N_12636,N_12504,N_12533);
and U12637 (N_12637,N_12535,N_12525);
nand U12638 (N_12638,N_12513,N_12588);
nand U12639 (N_12639,N_12544,N_12564);
and U12640 (N_12640,N_12509,N_12526);
nand U12641 (N_12641,N_12455,N_12597);
or U12642 (N_12642,N_12462,N_12572);
nor U12643 (N_12643,N_12539,N_12563);
nand U12644 (N_12644,N_12472,N_12481);
or U12645 (N_12645,N_12523,N_12489);
and U12646 (N_12646,N_12550,N_12473);
and U12647 (N_12647,N_12558,N_12560);
or U12648 (N_12648,N_12501,N_12502);
xor U12649 (N_12649,N_12521,N_12540);
xor U12650 (N_12650,N_12581,N_12470);
or U12651 (N_12651,N_12499,N_12496);
and U12652 (N_12652,N_12541,N_12547);
xnor U12653 (N_12653,N_12459,N_12584);
nand U12654 (N_12654,N_12573,N_12511);
nand U12655 (N_12655,N_12578,N_12464);
nor U12656 (N_12656,N_12491,N_12469);
and U12657 (N_12657,N_12498,N_12500);
or U12658 (N_12658,N_12452,N_12492);
xnor U12659 (N_12659,N_12548,N_12484);
and U12660 (N_12660,N_12598,N_12471);
or U12661 (N_12661,N_12549,N_12576);
or U12662 (N_12662,N_12582,N_12580);
and U12663 (N_12663,N_12512,N_12569);
xor U12664 (N_12664,N_12574,N_12595);
and U12665 (N_12665,N_12545,N_12559);
or U12666 (N_12666,N_12556,N_12518);
or U12667 (N_12667,N_12457,N_12476);
and U12668 (N_12668,N_12458,N_12487);
or U12669 (N_12669,N_12586,N_12480);
nor U12670 (N_12670,N_12529,N_12477);
and U12671 (N_12671,N_12456,N_12507);
and U12672 (N_12672,N_12519,N_12490);
xor U12673 (N_12673,N_12528,N_12590);
nand U12674 (N_12674,N_12479,N_12538);
nand U12675 (N_12675,N_12506,N_12479);
or U12676 (N_12676,N_12575,N_12458);
nor U12677 (N_12677,N_12489,N_12490);
or U12678 (N_12678,N_12581,N_12544);
and U12679 (N_12679,N_12495,N_12576);
nor U12680 (N_12680,N_12497,N_12581);
nor U12681 (N_12681,N_12514,N_12573);
and U12682 (N_12682,N_12535,N_12511);
nand U12683 (N_12683,N_12529,N_12517);
and U12684 (N_12684,N_12540,N_12474);
nor U12685 (N_12685,N_12463,N_12595);
nor U12686 (N_12686,N_12528,N_12512);
nand U12687 (N_12687,N_12521,N_12587);
xnor U12688 (N_12688,N_12467,N_12456);
and U12689 (N_12689,N_12538,N_12488);
and U12690 (N_12690,N_12522,N_12474);
xnor U12691 (N_12691,N_12541,N_12520);
or U12692 (N_12692,N_12562,N_12597);
or U12693 (N_12693,N_12577,N_12485);
or U12694 (N_12694,N_12522,N_12511);
and U12695 (N_12695,N_12589,N_12523);
nand U12696 (N_12696,N_12507,N_12457);
xnor U12697 (N_12697,N_12494,N_12548);
and U12698 (N_12698,N_12563,N_12505);
nand U12699 (N_12699,N_12594,N_12521);
nand U12700 (N_12700,N_12453,N_12526);
and U12701 (N_12701,N_12561,N_12556);
and U12702 (N_12702,N_12561,N_12536);
and U12703 (N_12703,N_12523,N_12587);
nor U12704 (N_12704,N_12576,N_12577);
xnor U12705 (N_12705,N_12563,N_12466);
nor U12706 (N_12706,N_12504,N_12524);
nor U12707 (N_12707,N_12485,N_12575);
and U12708 (N_12708,N_12515,N_12505);
xnor U12709 (N_12709,N_12508,N_12480);
nand U12710 (N_12710,N_12457,N_12462);
and U12711 (N_12711,N_12453,N_12498);
and U12712 (N_12712,N_12586,N_12577);
and U12713 (N_12713,N_12581,N_12542);
xnor U12714 (N_12714,N_12579,N_12531);
xnor U12715 (N_12715,N_12596,N_12597);
xor U12716 (N_12716,N_12475,N_12560);
nand U12717 (N_12717,N_12487,N_12583);
xnor U12718 (N_12718,N_12572,N_12532);
nand U12719 (N_12719,N_12511,N_12576);
nor U12720 (N_12720,N_12471,N_12545);
or U12721 (N_12721,N_12516,N_12586);
and U12722 (N_12722,N_12577,N_12481);
nor U12723 (N_12723,N_12506,N_12519);
or U12724 (N_12724,N_12545,N_12546);
xnor U12725 (N_12725,N_12580,N_12551);
nor U12726 (N_12726,N_12543,N_12537);
xnor U12727 (N_12727,N_12563,N_12574);
and U12728 (N_12728,N_12536,N_12592);
xnor U12729 (N_12729,N_12542,N_12469);
nor U12730 (N_12730,N_12534,N_12501);
or U12731 (N_12731,N_12537,N_12475);
nor U12732 (N_12732,N_12590,N_12513);
xor U12733 (N_12733,N_12545,N_12593);
nand U12734 (N_12734,N_12477,N_12499);
and U12735 (N_12735,N_12476,N_12592);
nor U12736 (N_12736,N_12477,N_12510);
and U12737 (N_12737,N_12495,N_12519);
or U12738 (N_12738,N_12585,N_12491);
and U12739 (N_12739,N_12580,N_12460);
or U12740 (N_12740,N_12516,N_12580);
and U12741 (N_12741,N_12451,N_12573);
nor U12742 (N_12742,N_12580,N_12486);
nand U12743 (N_12743,N_12515,N_12517);
xor U12744 (N_12744,N_12460,N_12540);
or U12745 (N_12745,N_12464,N_12459);
nand U12746 (N_12746,N_12494,N_12455);
nor U12747 (N_12747,N_12529,N_12462);
xor U12748 (N_12748,N_12590,N_12576);
and U12749 (N_12749,N_12490,N_12505);
nand U12750 (N_12750,N_12678,N_12690);
xnor U12751 (N_12751,N_12718,N_12691);
nand U12752 (N_12752,N_12693,N_12670);
and U12753 (N_12753,N_12710,N_12709);
and U12754 (N_12754,N_12640,N_12673);
nor U12755 (N_12755,N_12720,N_12695);
or U12756 (N_12756,N_12630,N_12745);
nand U12757 (N_12757,N_12610,N_12740);
nor U12758 (N_12758,N_12659,N_12611);
xnor U12759 (N_12759,N_12737,N_12624);
xor U12760 (N_12760,N_12604,N_12620);
xor U12761 (N_12761,N_12618,N_12636);
xnor U12762 (N_12762,N_12644,N_12734);
nor U12763 (N_12763,N_12664,N_12739);
xnor U12764 (N_12764,N_12680,N_12742);
nor U12765 (N_12765,N_12615,N_12622);
xnor U12766 (N_12766,N_12667,N_12717);
and U12767 (N_12767,N_12602,N_12735);
nor U12768 (N_12768,N_12650,N_12703);
xnor U12769 (N_12769,N_12660,N_12689);
xnor U12770 (N_12770,N_12614,N_12635);
and U12771 (N_12771,N_12712,N_12617);
xor U12772 (N_12772,N_12738,N_12608);
xor U12773 (N_12773,N_12747,N_12649);
nand U12774 (N_12774,N_12697,N_12731);
and U12775 (N_12775,N_12707,N_12621);
xnor U12776 (N_12776,N_12662,N_12651);
nor U12777 (N_12777,N_12656,N_12623);
xor U12778 (N_12778,N_12696,N_12672);
nand U12779 (N_12779,N_12619,N_12666);
nand U12780 (N_12780,N_12679,N_12665);
nand U12781 (N_12781,N_12634,N_12741);
or U12782 (N_12782,N_12729,N_12653);
xor U12783 (N_12783,N_12727,N_12724);
nor U12784 (N_12784,N_12600,N_12674);
or U12785 (N_12785,N_12688,N_12645);
xor U12786 (N_12786,N_12705,N_12669);
nor U12787 (N_12787,N_12642,N_12725);
xor U12788 (N_12788,N_12748,N_12694);
and U12789 (N_12789,N_12652,N_12704);
xnor U12790 (N_12790,N_12629,N_12713);
and U12791 (N_12791,N_12722,N_12733);
xnor U12792 (N_12792,N_12657,N_12671);
xor U12793 (N_12793,N_12719,N_12677);
nor U12794 (N_12794,N_12609,N_12648);
or U12795 (N_12795,N_12607,N_12744);
or U12796 (N_12796,N_12627,N_12639);
nand U12797 (N_12797,N_12631,N_12723);
nand U12798 (N_12798,N_12628,N_12726);
nor U12799 (N_12799,N_12702,N_12654);
xnor U12800 (N_12800,N_12684,N_12601);
nand U12801 (N_12801,N_12701,N_12728);
nor U12802 (N_12802,N_12683,N_12626);
nor U12803 (N_12803,N_12686,N_12663);
nand U12804 (N_12804,N_12711,N_12655);
xor U12805 (N_12805,N_12681,N_12612);
nand U12806 (N_12806,N_12708,N_12668);
or U12807 (N_12807,N_12687,N_12746);
nand U12808 (N_12808,N_12638,N_12641);
or U12809 (N_12809,N_12732,N_12700);
nand U12810 (N_12810,N_12676,N_12706);
and U12811 (N_12811,N_12637,N_12632);
xor U12812 (N_12812,N_12714,N_12715);
or U12813 (N_12813,N_12743,N_12625);
nor U12814 (N_12814,N_12699,N_12616);
or U12815 (N_12815,N_12613,N_12698);
and U12816 (N_12816,N_12633,N_12605);
nor U12817 (N_12817,N_12692,N_12721);
nand U12818 (N_12818,N_12647,N_12646);
nand U12819 (N_12819,N_12661,N_12749);
or U12820 (N_12820,N_12685,N_12643);
nand U12821 (N_12821,N_12736,N_12658);
xnor U12822 (N_12822,N_12730,N_12682);
and U12823 (N_12823,N_12675,N_12716);
nor U12824 (N_12824,N_12606,N_12603);
or U12825 (N_12825,N_12640,N_12739);
nor U12826 (N_12826,N_12670,N_12610);
and U12827 (N_12827,N_12729,N_12636);
xnor U12828 (N_12828,N_12612,N_12615);
and U12829 (N_12829,N_12666,N_12670);
nand U12830 (N_12830,N_12733,N_12623);
xor U12831 (N_12831,N_12668,N_12682);
nand U12832 (N_12832,N_12730,N_12679);
xnor U12833 (N_12833,N_12671,N_12674);
nand U12834 (N_12834,N_12628,N_12617);
and U12835 (N_12835,N_12703,N_12715);
and U12836 (N_12836,N_12657,N_12620);
or U12837 (N_12837,N_12683,N_12659);
and U12838 (N_12838,N_12692,N_12724);
xor U12839 (N_12839,N_12603,N_12683);
or U12840 (N_12840,N_12652,N_12738);
or U12841 (N_12841,N_12625,N_12682);
or U12842 (N_12842,N_12672,N_12625);
xnor U12843 (N_12843,N_12651,N_12724);
nand U12844 (N_12844,N_12718,N_12674);
xor U12845 (N_12845,N_12684,N_12678);
and U12846 (N_12846,N_12732,N_12647);
nor U12847 (N_12847,N_12613,N_12693);
and U12848 (N_12848,N_12646,N_12607);
and U12849 (N_12849,N_12731,N_12671);
or U12850 (N_12850,N_12685,N_12610);
and U12851 (N_12851,N_12602,N_12634);
or U12852 (N_12852,N_12675,N_12618);
nand U12853 (N_12853,N_12616,N_12719);
or U12854 (N_12854,N_12704,N_12705);
or U12855 (N_12855,N_12714,N_12605);
nor U12856 (N_12856,N_12689,N_12637);
nand U12857 (N_12857,N_12664,N_12642);
nor U12858 (N_12858,N_12600,N_12648);
and U12859 (N_12859,N_12749,N_12678);
nand U12860 (N_12860,N_12613,N_12683);
xnor U12861 (N_12861,N_12659,N_12703);
nand U12862 (N_12862,N_12600,N_12728);
and U12863 (N_12863,N_12613,N_12656);
and U12864 (N_12864,N_12723,N_12612);
xor U12865 (N_12865,N_12601,N_12715);
nand U12866 (N_12866,N_12747,N_12643);
xnor U12867 (N_12867,N_12730,N_12659);
and U12868 (N_12868,N_12687,N_12740);
nor U12869 (N_12869,N_12734,N_12720);
and U12870 (N_12870,N_12629,N_12668);
nand U12871 (N_12871,N_12685,N_12706);
or U12872 (N_12872,N_12714,N_12717);
and U12873 (N_12873,N_12693,N_12708);
and U12874 (N_12874,N_12607,N_12700);
nor U12875 (N_12875,N_12732,N_12685);
nor U12876 (N_12876,N_12710,N_12655);
nand U12877 (N_12877,N_12720,N_12652);
and U12878 (N_12878,N_12726,N_12643);
xor U12879 (N_12879,N_12604,N_12741);
xor U12880 (N_12880,N_12683,N_12694);
xor U12881 (N_12881,N_12609,N_12646);
or U12882 (N_12882,N_12656,N_12736);
and U12883 (N_12883,N_12615,N_12718);
or U12884 (N_12884,N_12728,N_12699);
nand U12885 (N_12885,N_12688,N_12661);
nor U12886 (N_12886,N_12631,N_12709);
and U12887 (N_12887,N_12619,N_12728);
nor U12888 (N_12888,N_12682,N_12692);
nor U12889 (N_12889,N_12701,N_12661);
nor U12890 (N_12890,N_12610,N_12615);
nand U12891 (N_12891,N_12675,N_12714);
and U12892 (N_12892,N_12657,N_12670);
and U12893 (N_12893,N_12601,N_12636);
xor U12894 (N_12894,N_12698,N_12747);
nor U12895 (N_12895,N_12714,N_12744);
xnor U12896 (N_12896,N_12700,N_12635);
nand U12897 (N_12897,N_12646,N_12626);
nor U12898 (N_12898,N_12705,N_12604);
and U12899 (N_12899,N_12736,N_12632);
or U12900 (N_12900,N_12853,N_12833);
or U12901 (N_12901,N_12784,N_12818);
nor U12902 (N_12902,N_12863,N_12874);
xor U12903 (N_12903,N_12854,N_12866);
and U12904 (N_12904,N_12865,N_12823);
or U12905 (N_12905,N_12819,N_12831);
or U12906 (N_12906,N_12851,N_12829);
nor U12907 (N_12907,N_12862,N_12797);
and U12908 (N_12908,N_12894,N_12801);
xnor U12909 (N_12909,N_12806,N_12888);
and U12910 (N_12910,N_12834,N_12792);
nand U12911 (N_12911,N_12824,N_12849);
nand U12912 (N_12912,N_12892,N_12870);
xor U12913 (N_12913,N_12864,N_12813);
nor U12914 (N_12914,N_12790,N_12771);
nor U12915 (N_12915,N_12846,N_12879);
nand U12916 (N_12916,N_12825,N_12798);
nor U12917 (N_12917,N_12876,N_12763);
or U12918 (N_12918,N_12860,N_12852);
and U12919 (N_12919,N_12855,N_12817);
nor U12920 (N_12920,N_12802,N_12884);
nand U12921 (N_12921,N_12767,N_12885);
xor U12922 (N_12922,N_12761,N_12857);
xor U12923 (N_12923,N_12832,N_12880);
and U12924 (N_12924,N_12783,N_12780);
nand U12925 (N_12925,N_12753,N_12858);
nor U12926 (N_12926,N_12848,N_12899);
nor U12927 (N_12927,N_12886,N_12873);
xor U12928 (N_12928,N_12845,N_12786);
nand U12929 (N_12929,N_12856,N_12755);
and U12930 (N_12930,N_12777,N_12882);
xnor U12931 (N_12931,N_12807,N_12838);
and U12932 (N_12932,N_12835,N_12809);
nand U12933 (N_12933,N_12859,N_12781);
xor U12934 (N_12934,N_12800,N_12768);
nor U12935 (N_12935,N_12841,N_12757);
and U12936 (N_12936,N_12822,N_12787);
and U12937 (N_12937,N_12872,N_12896);
xnor U12938 (N_12938,N_12789,N_12890);
nand U12939 (N_12939,N_12760,N_12821);
xnor U12940 (N_12940,N_12772,N_12750);
nand U12941 (N_12941,N_12816,N_12847);
xnor U12942 (N_12942,N_12808,N_12837);
nor U12943 (N_12943,N_12765,N_12889);
nand U12944 (N_12944,N_12871,N_12881);
or U12945 (N_12945,N_12811,N_12814);
xnor U12946 (N_12946,N_12812,N_12895);
xnor U12947 (N_12947,N_12898,N_12785);
and U12948 (N_12948,N_12788,N_12751);
and U12949 (N_12949,N_12754,N_12867);
nor U12950 (N_12950,N_12773,N_12869);
and U12951 (N_12951,N_12810,N_12778);
nor U12952 (N_12952,N_12794,N_12766);
nand U12953 (N_12953,N_12759,N_12782);
and U12954 (N_12954,N_12878,N_12887);
nor U12955 (N_12955,N_12793,N_12799);
and U12956 (N_12956,N_12827,N_12805);
or U12957 (N_12957,N_12776,N_12828);
or U12958 (N_12958,N_12752,N_12843);
and U12959 (N_12959,N_12769,N_12836);
and U12960 (N_12960,N_12796,N_12774);
nor U12961 (N_12961,N_12891,N_12844);
nor U12962 (N_12962,N_12839,N_12791);
or U12963 (N_12963,N_12762,N_12775);
nand U12964 (N_12964,N_12842,N_12883);
and U12965 (N_12965,N_12779,N_12897);
and U12966 (N_12966,N_12820,N_12877);
nor U12967 (N_12967,N_12868,N_12850);
or U12968 (N_12968,N_12875,N_12815);
and U12969 (N_12969,N_12804,N_12826);
or U12970 (N_12970,N_12830,N_12758);
xor U12971 (N_12971,N_12840,N_12795);
nand U12972 (N_12972,N_12770,N_12861);
and U12973 (N_12973,N_12893,N_12764);
xnor U12974 (N_12974,N_12756,N_12803);
xnor U12975 (N_12975,N_12804,N_12774);
nand U12976 (N_12976,N_12802,N_12768);
or U12977 (N_12977,N_12822,N_12823);
and U12978 (N_12978,N_12840,N_12753);
nand U12979 (N_12979,N_12835,N_12851);
nor U12980 (N_12980,N_12828,N_12822);
or U12981 (N_12981,N_12790,N_12897);
and U12982 (N_12982,N_12803,N_12814);
xnor U12983 (N_12983,N_12758,N_12815);
nand U12984 (N_12984,N_12896,N_12801);
xnor U12985 (N_12985,N_12862,N_12865);
nand U12986 (N_12986,N_12815,N_12885);
nand U12987 (N_12987,N_12852,N_12759);
or U12988 (N_12988,N_12830,N_12818);
nand U12989 (N_12989,N_12866,N_12896);
or U12990 (N_12990,N_12810,N_12879);
and U12991 (N_12991,N_12783,N_12837);
nor U12992 (N_12992,N_12854,N_12877);
nand U12993 (N_12993,N_12780,N_12889);
nand U12994 (N_12994,N_12862,N_12822);
or U12995 (N_12995,N_12793,N_12859);
xor U12996 (N_12996,N_12762,N_12798);
xor U12997 (N_12997,N_12750,N_12755);
xnor U12998 (N_12998,N_12855,N_12802);
nor U12999 (N_12999,N_12878,N_12870);
nor U13000 (N_13000,N_12888,N_12776);
or U13001 (N_13001,N_12774,N_12871);
xor U13002 (N_13002,N_12888,N_12798);
xor U13003 (N_13003,N_12868,N_12755);
xor U13004 (N_13004,N_12870,N_12811);
nand U13005 (N_13005,N_12848,N_12843);
nor U13006 (N_13006,N_12895,N_12779);
nand U13007 (N_13007,N_12767,N_12783);
and U13008 (N_13008,N_12831,N_12784);
and U13009 (N_13009,N_12782,N_12797);
nor U13010 (N_13010,N_12803,N_12839);
xor U13011 (N_13011,N_12847,N_12866);
nand U13012 (N_13012,N_12872,N_12885);
xor U13013 (N_13013,N_12801,N_12833);
and U13014 (N_13014,N_12789,N_12754);
xnor U13015 (N_13015,N_12835,N_12844);
nor U13016 (N_13016,N_12850,N_12792);
or U13017 (N_13017,N_12786,N_12767);
nand U13018 (N_13018,N_12812,N_12752);
xnor U13019 (N_13019,N_12774,N_12770);
or U13020 (N_13020,N_12751,N_12823);
or U13021 (N_13021,N_12836,N_12825);
xnor U13022 (N_13022,N_12801,N_12829);
nand U13023 (N_13023,N_12848,N_12866);
and U13024 (N_13024,N_12826,N_12876);
and U13025 (N_13025,N_12895,N_12873);
nor U13026 (N_13026,N_12796,N_12823);
xnor U13027 (N_13027,N_12895,N_12754);
xnor U13028 (N_13028,N_12869,N_12838);
xnor U13029 (N_13029,N_12832,N_12814);
nor U13030 (N_13030,N_12831,N_12753);
and U13031 (N_13031,N_12801,N_12826);
or U13032 (N_13032,N_12894,N_12866);
and U13033 (N_13033,N_12856,N_12775);
nand U13034 (N_13034,N_12890,N_12827);
and U13035 (N_13035,N_12783,N_12877);
or U13036 (N_13036,N_12832,N_12774);
nor U13037 (N_13037,N_12766,N_12878);
or U13038 (N_13038,N_12873,N_12807);
or U13039 (N_13039,N_12808,N_12750);
xnor U13040 (N_13040,N_12881,N_12897);
nor U13041 (N_13041,N_12840,N_12765);
xnor U13042 (N_13042,N_12823,N_12811);
xor U13043 (N_13043,N_12868,N_12874);
xnor U13044 (N_13044,N_12852,N_12835);
or U13045 (N_13045,N_12875,N_12840);
nor U13046 (N_13046,N_12798,N_12768);
and U13047 (N_13047,N_12863,N_12821);
nor U13048 (N_13048,N_12774,N_12785);
xnor U13049 (N_13049,N_12777,N_12843);
and U13050 (N_13050,N_12992,N_12946);
xnor U13051 (N_13051,N_12928,N_13010);
nand U13052 (N_13052,N_12990,N_13038);
or U13053 (N_13053,N_12931,N_12934);
or U13054 (N_13054,N_13032,N_12966);
and U13055 (N_13055,N_13021,N_12981);
nor U13056 (N_13056,N_13033,N_12912);
xnor U13057 (N_13057,N_12913,N_12922);
nand U13058 (N_13058,N_12910,N_13036);
and U13059 (N_13059,N_13001,N_13027);
and U13060 (N_13060,N_13013,N_12907);
or U13061 (N_13061,N_12900,N_12983);
and U13062 (N_13062,N_13043,N_12943);
xor U13063 (N_13063,N_13049,N_12933);
nand U13064 (N_13064,N_13037,N_12961);
or U13065 (N_13065,N_12955,N_13015);
and U13066 (N_13066,N_12915,N_12987);
and U13067 (N_13067,N_13026,N_12942);
xor U13068 (N_13068,N_12918,N_12996);
or U13069 (N_13069,N_12984,N_12967);
nand U13070 (N_13070,N_13009,N_12973);
or U13071 (N_13071,N_12976,N_12953);
xor U13072 (N_13072,N_12998,N_12901);
nand U13073 (N_13073,N_13041,N_12989);
xor U13074 (N_13074,N_12963,N_13014);
xor U13075 (N_13075,N_12950,N_12991);
xor U13076 (N_13076,N_13002,N_12916);
nor U13077 (N_13077,N_12937,N_12979);
nor U13078 (N_13078,N_12908,N_13031);
nor U13079 (N_13079,N_12959,N_12972);
nor U13080 (N_13080,N_12919,N_12954);
nor U13081 (N_13081,N_12904,N_12936);
nand U13082 (N_13082,N_12964,N_12965);
xnor U13083 (N_13083,N_12995,N_12938);
nand U13084 (N_13084,N_13019,N_12960);
and U13085 (N_13085,N_13034,N_12999);
or U13086 (N_13086,N_12914,N_13007);
nor U13087 (N_13087,N_12929,N_12988);
and U13088 (N_13088,N_13040,N_12923);
or U13089 (N_13089,N_13048,N_13017);
nand U13090 (N_13090,N_13004,N_12993);
and U13091 (N_13091,N_12985,N_13016);
or U13092 (N_13092,N_12969,N_12994);
nand U13093 (N_13093,N_13012,N_12940);
or U13094 (N_13094,N_12903,N_12939);
nand U13095 (N_13095,N_12952,N_13035);
or U13096 (N_13096,N_13025,N_13039);
and U13097 (N_13097,N_12971,N_12978);
and U13098 (N_13098,N_13005,N_12956);
nand U13099 (N_13099,N_13020,N_12911);
nor U13100 (N_13100,N_12980,N_12974);
nor U13101 (N_13101,N_12920,N_12932);
or U13102 (N_13102,N_13000,N_12944);
and U13103 (N_13103,N_12962,N_12947);
nand U13104 (N_13104,N_12975,N_13023);
and U13105 (N_13105,N_13018,N_12970);
xnor U13106 (N_13106,N_13030,N_13006);
nor U13107 (N_13107,N_12986,N_13008);
xnor U13108 (N_13108,N_12906,N_12925);
nand U13109 (N_13109,N_13045,N_13003);
nand U13110 (N_13110,N_13046,N_12902);
xor U13111 (N_13111,N_12905,N_13047);
nand U13112 (N_13112,N_12935,N_12917);
and U13113 (N_13113,N_12951,N_12957);
nand U13114 (N_13114,N_13044,N_12926);
nand U13115 (N_13115,N_12930,N_13028);
xor U13116 (N_13116,N_12949,N_12997);
nor U13117 (N_13117,N_12909,N_12941);
and U13118 (N_13118,N_12927,N_12968);
or U13119 (N_13119,N_13042,N_13022);
nor U13120 (N_13120,N_12921,N_12948);
nand U13121 (N_13121,N_12977,N_13024);
or U13122 (N_13122,N_12982,N_12945);
nor U13123 (N_13123,N_13029,N_13011);
nand U13124 (N_13124,N_12958,N_12924);
or U13125 (N_13125,N_12922,N_12943);
xor U13126 (N_13126,N_13032,N_12926);
nand U13127 (N_13127,N_12961,N_12931);
nand U13128 (N_13128,N_13023,N_12933);
or U13129 (N_13129,N_12916,N_12924);
nand U13130 (N_13130,N_13032,N_12997);
or U13131 (N_13131,N_12998,N_12991);
xor U13132 (N_13132,N_12929,N_13029);
nor U13133 (N_13133,N_13024,N_12986);
xor U13134 (N_13134,N_12921,N_13008);
or U13135 (N_13135,N_13000,N_12942);
nand U13136 (N_13136,N_13044,N_12965);
nor U13137 (N_13137,N_13004,N_12976);
or U13138 (N_13138,N_12935,N_13043);
and U13139 (N_13139,N_13036,N_12996);
nor U13140 (N_13140,N_12974,N_13046);
xnor U13141 (N_13141,N_12924,N_12903);
nand U13142 (N_13142,N_12971,N_12909);
xor U13143 (N_13143,N_12958,N_12925);
and U13144 (N_13144,N_13041,N_12974);
xnor U13145 (N_13145,N_12995,N_12973);
or U13146 (N_13146,N_13048,N_12903);
and U13147 (N_13147,N_13045,N_13011);
nor U13148 (N_13148,N_13041,N_12972);
nor U13149 (N_13149,N_13007,N_12950);
nor U13150 (N_13150,N_12954,N_13035);
nor U13151 (N_13151,N_12965,N_12963);
nor U13152 (N_13152,N_12962,N_13015);
or U13153 (N_13153,N_13038,N_12985);
nand U13154 (N_13154,N_12949,N_12989);
and U13155 (N_13155,N_12987,N_12925);
nand U13156 (N_13156,N_12934,N_12992);
or U13157 (N_13157,N_13041,N_12957);
and U13158 (N_13158,N_12934,N_13038);
or U13159 (N_13159,N_12962,N_12942);
and U13160 (N_13160,N_12907,N_12977);
or U13161 (N_13161,N_12911,N_13002);
or U13162 (N_13162,N_12998,N_13045);
or U13163 (N_13163,N_12987,N_13013);
and U13164 (N_13164,N_12956,N_12949);
and U13165 (N_13165,N_12935,N_12976);
nand U13166 (N_13166,N_12996,N_12939);
nor U13167 (N_13167,N_13026,N_12981);
xnor U13168 (N_13168,N_13048,N_12907);
nand U13169 (N_13169,N_12955,N_13030);
nor U13170 (N_13170,N_13012,N_12926);
and U13171 (N_13171,N_12997,N_12958);
xnor U13172 (N_13172,N_12943,N_12991);
or U13173 (N_13173,N_13035,N_12908);
nand U13174 (N_13174,N_13016,N_12994);
and U13175 (N_13175,N_13040,N_12969);
nor U13176 (N_13176,N_12954,N_13046);
nor U13177 (N_13177,N_12916,N_12979);
nor U13178 (N_13178,N_12981,N_13000);
and U13179 (N_13179,N_12934,N_12947);
xor U13180 (N_13180,N_12996,N_13011);
nor U13181 (N_13181,N_12979,N_13041);
and U13182 (N_13182,N_13012,N_12963);
xor U13183 (N_13183,N_13033,N_12992);
nor U13184 (N_13184,N_12993,N_12953);
or U13185 (N_13185,N_12923,N_12905);
xnor U13186 (N_13186,N_12932,N_12961);
and U13187 (N_13187,N_13041,N_13044);
or U13188 (N_13188,N_12971,N_12934);
nor U13189 (N_13189,N_12962,N_13012);
and U13190 (N_13190,N_13004,N_13036);
xor U13191 (N_13191,N_12915,N_12985);
nor U13192 (N_13192,N_13037,N_13030);
and U13193 (N_13193,N_12948,N_12938);
nor U13194 (N_13194,N_13006,N_13011);
nor U13195 (N_13195,N_13034,N_12966);
nand U13196 (N_13196,N_13041,N_13047);
nand U13197 (N_13197,N_13015,N_12971);
nand U13198 (N_13198,N_12966,N_12997);
xnor U13199 (N_13199,N_12966,N_12921);
and U13200 (N_13200,N_13190,N_13107);
and U13201 (N_13201,N_13070,N_13073);
xnor U13202 (N_13202,N_13184,N_13100);
nand U13203 (N_13203,N_13164,N_13122);
and U13204 (N_13204,N_13153,N_13099);
nand U13205 (N_13205,N_13054,N_13067);
nand U13206 (N_13206,N_13063,N_13147);
and U13207 (N_13207,N_13088,N_13165);
xnor U13208 (N_13208,N_13155,N_13050);
xnor U13209 (N_13209,N_13149,N_13182);
nor U13210 (N_13210,N_13186,N_13196);
xnor U13211 (N_13211,N_13144,N_13118);
and U13212 (N_13212,N_13093,N_13151);
xor U13213 (N_13213,N_13148,N_13058);
and U13214 (N_13214,N_13171,N_13136);
or U13215 (N_13215,N_13095,N_13142);
nor U13216 (N_13216,N_13178,N_13121);
xor U13217 (N_13217,N_13119,N_13176);
and U13218 (N_13218,N_13077,N_13198);
xnor U13219 (N_13219,N_13168,N_13113);
and U13220 (N_13220,N_13120,N_13154);
nor U13221 (N_13221,N_13084,N_13111);
nor U13222 (N_13222,N_13081,N_13064);
nand U13223 (N_13223,N_13065,N_13087);
and U13224 (N_13224,N_13195,N_13108);
nor U13225 (N_13225,N_13090,N_13072);
nor U13226 (N_13226,N_13132,N_13083);
and U13227 (N_13227,N_13157,N_13059);
or U13228 (N_13228,N_13085,N_13160);
nor U13229 (N_13229,N_13173,N_13152);
nor U13230 (N_13230,N_13078,N_13109);
xor U13231 (N_13231,N_13066,N_13055);
and U13232 (N_13232,N_13141,N_13075);
nand U13233 (N_13233,N_13193,N_13053);
xnor U13234 (N_13234,N_13146,N_13102);
nor U13235 (N_13235,N_13076,N_13130);
nor U13236 (N_13236,N_13123,N_13129);
nor U13237 (N_13237,N_13098,N_13140);
and U13238 (N_13238,N_13180,N_13194);
nand U13239 (N_13239,N_13057,N_13061);
or U13240 (N_13240,N_13069,N_13110);
xnor U13241 (N_13241,N_13089,N_13117);
nand U13242 (N_13242,N_13051,N_13188);
nand U13243 (N_13243,N_13137,N_13172);
nand U13244 (N_13244,N_13127,N_13133);
nand U13245 (N_13245,N_13125,N_13162);
nand U13246 (N_13246,N_13163,N_13096);
and U13247 (N_13247,N_13092,N_13101);
nand U13248 (N_13248,N_13128,N_13179);
xnor U13249 (N_13249,N_13114,N_13103);
or U13250 (N_13250,N_13169,N_13056);
or U13251 (N_13251,N_13192,N_13097);
nor U13252 (N_13252,N_13071,N_13052);
or U13253 (N_13253,N_13183,N_13124);
and U13254 (N_13254,N_13197,N_13150);
or U13255 (N_13255,N_13126,N_13167);
nand U13256 (N_13256,N_13185,N_13094);
nand U13257 (N_13257,N_13115,N_13131);
and U13258 (N_13258,N_13199,N_13086);
nand U13259 (N_13259,N_13106,N_13105);
or U13260 (N_13260,N_13074,N_13091);
nor U13261 (N_13261,N_13060,N_13082);
nor U13262 (N_13262,N_13143,N_13191);
nand U13263 (N_13263,N_13080,N_13181);
nand U13264 (N_13264,N_13145,N_13161);
nand U13265 (N_13265,N_13177,N_13068);
or U13266 (N_13266,N_13138,N_13135);
nand U13267 (N_13267,N_13166,N_13159);
nor U13268 (N_13268,N_13134,N_13189);
xor U13269 (N_13269,N_13175,N_13187);
xor U13270 (N_13270,N_13062,N_13104);
and U13271 (N_13271,N_13156,N_13116);
and U13272 (N_13272,N_13158,N_13174);
nor U13273 (N_13273,N_13112,N_13139);
or U13274 (N_13274,N_13170,N_13079);
or U13275 (N_13275,N_13161,N_13059);
xor U13276 (N_13276,N_13141,N_13156);
xor U13277 (N_13277,N_13075,N_13175);
nor U13278 (N_13278,N_13083,N_13087);
nor U13279 (N_13279,N_13067,N_13068);
xnor U13280 (N_13280,N_13052,N_13102);
nor U13281 (N_13281,N_13150,N_13194);
or U13282 (N_13282,N_13114,N_13150);
or U13283 (N_13283,N_13139,N_13117);
or U13284 (N_13284,N_13192,N_13105);
and U13285 (N_13285,N_13171,N_13094);
nor U13286 (N_13286,N_13133,N_13160);
and U13287 (N_13287,N_13133,N_13177);
xnor U13288 (N_13288,N_13054,N_13175);
nand U13289 (N_13289,N_13137,N_13133);
xnor U13290 (N_13290,N_13142,N_13109);
nand U13291 (N_13291,N_13098,N_13084);
nor U13292 (N_13292,N_13069,N_13190);
nor U13293 (N_13293,N_13164,N_13131);
nor U13294 (N_13294,N_13071,N_13182);
nor U13295 (N_13295,N_13052,N_13091);
nand U13296 (N_13296,N_13128,N_13083);
and U13297 (N_13297,N_13113,N_13126);
or U13298 (N_13298,N_13114,N_13139);
xor U13299 (N_13299,N_13136,N_13064);
or U13300 (N_13300,N_13077,N_13084);
nor U13301 (N_13301,N_13116,N_13142);
xor U13302 (N_13302,N_13058,N_13144);
and U13303 (N_13303,N_13093,N_13190);
or U13304 (N_13304,N_13184,N_13117);
xnor U13305 (N_13305,N_13052,N_13069);
nand U13306 (N_13306,N_13185,N_13097);
and U13307 (N_13307,N_13140,N_13058);
or U13308 (N_13308,N_13142,N_13075);
or U13309 (N_13309,N_13198,N_13104);
and U13310 (N_13310,N_13080,N_13170);
nand U13311 (N_13311,N_13109,N_13098);
and U13312 (N_13312,N_13074,N_13071);
or U13313 (N_13313,N_13063,N_13162);
nor U13314 (N_13314,N_13172,N_13093);
nand U13315 (N_13315,N_13086,N_13193);
nor U13316 (N_13316,N_13112,N_13075);
xor U13317 (N_13317,N_13066,N_13089);
xnor U13318 (N_13318,N_13135,N_13120);
nand U13319 (N_13319,N_13112,N_13104);
nor U13320 (N_13320,N_13195,N_13142);
nor U13321 (N_13321,N_13121,N_13080);
nor U13322 (N_13322,N_13074,N_13127);
nor U13323 (N_13323,N_13147,N_13104);
nor U13324 (N_13324,N_13173,N_13177);
nand U13325 (N_13325,N_13176,N_13093);
nor U13326 (N_13326,N_13182,N_13168);
nand U13327 (N_13327,N_13176,N_13060);
and U13328 (N_13328,N_13172,N_13057);
and U13329 (N_13329,N_13072,N_13149);
nor U13330 (N_13330,N_13145,N_13184);
xor U13331 (N_13331,N_13157,N_13055);
nand U13332 (N_13332,N_13099,N_13081);
and U13333 (N_13333,N_13116,N_13115);
xor U13334 (N_13334,N_13074,N_13075);
xnor U13335 (N_13335,N_13056,N_13071);
and U13336 (N_13336,N_13127,N_13097);
xor U13337 (N_13337,N_13112,N_13064);
nand U13338 (N_13338,N_13114,N_13132);
or U13339 (N_13339,N_13174,N_13177);
nor U13340 (N_13340,N_13091,N_13084);
or U13341 (N_13341,N_13148,N_13149);
nand U13342 (N_13342,N_13074,N_13141);
and U13343 (N_13343,N_13123,N_13161);
and U13344 (N_13344,N_13172,N_13173);
or U13345 (N_13345,N_13131,N_13139);
nand U13346 (N_13346,N_13072,N_13176);
nor U13347 (N_13347,N_13059,N_13096);
and U13348 (N_13348,N_13143,N_13180);
xnor U13349 (N_13349,N_13130,N_13181);
and U13350 (N_13350,N_13250,N_13276);
and U13351 (N_13351,N_13237,N_13227);
and U13352 (N_13352,N_13293,N_13267);
or U13353 (N_13353,N_13261,N_13311);
xor U13354 (N_13354,N_13304,N_13228);
xnor U13355 (N_13355,N_13294,N_13266);
and U13356 (N_13356,N_13326,N_13215);
and U13357 (N_13357,N_13256,N_13305);
and U13358 (N_13358,N_13283,N_13341);
or U13359 (N_13359,N_13285,N_13342);
or U13360 (N_13360,N_13345,N_13322);
or U13361 (N_13361,N_13269,N_13264);
and U13362 (N_13362,N_13275,N_13253);
nor U13363 (N_13363,N_13235,N_13254);
xnor U13364 (N_13364,N_13248,N_13218);
nand U13365 (N_13365,N_13244,N_13329);
xnor U13366 (N_13366,N_13299,N_13200);
xor U13367 (N_13367,N_13330,N_13204);
xor U13368 (N_13368,N_13317,N_13316);
or U13369 (N_13369,N_13309,N_13335);
nor U13370 (N_13370,N_13222,N_13270);
nor U13371 (N_13371,N_13224,N_13277);
xnor U13372 (N_13372,N_13312,N_13231);
xor U13373 (N_13373,N_13320,N_13259);
nor U13374 (N_13374,N_13336,N_13296);
nor U13375 (N_13375,N_13246,N_13298);
nor U13376 (N_13376,N_13306,N_13297);
nand U13377 (N_13377,N_13233,N_13287);
or U13378 (N_13378,N_13242,N_13308);
and U13379 (N_13379,N_13301,N_13258);
xnor U13380 (N_13380,N_13313,N_13347);
and U13381 (N_13381,N_13230,N_13315);
xnor U13382 (N_13382,N_13289,N_13257);
or U13383 (N_13383,N_13300,N_13262);
nand U13384 (N_13384,N_13273,N_13274);
and U13385 (N_13385,N_13290,N_13349);
or U13386 (N_13386,N_13201,N_13241);
nor U13387 (N_13387,N_13327,N_13221);
and U13388 (N_13388,N_13260,N_13234);
xnor U13389 (N_13389,N_13314,N_13214);
or U13390 (N_13390,N_13229,N_13265);
nor U13391 (N_13391,N_13205,N_13226);
and U13392 (N_13392,N_13339,N_13292);
nand U13393 (N_13393,N_13249,N_13279);
nand U13394 (N_13394,N_13245,N_13225);
xnor U13395 (N_13395,N_13321,N_13303);
nor U13396 (N_13396,N_13232,N_13272);
xor U13397 (N_13397,N_13211,N_13247);
or U13398 (N_13398,N_13282,N_13307);
nand U13399 (N_13399,N_13216,N_13203);
xnor U13400 (N_13400,N_13286,N_13344);
xor U13401 (N_13401,N_13243,N_13202);
xnor U13402 (N_13402,N_13323,N_13251);
and U13403 (N_13403,N_13209,N_13310);
or U13404 (N_13404,N_13288,N_13263);
or U13405 (N_13405,N_13328,N_13337);
xor U13406 (N_13406,N_13239,N_13324);
or U13407 (N_13407,N_13332,N_13252);
and U13408 (N_13408,N_13340,N_13331);
xor U13409 (N_13409,N_13302,N_13238);
nand U13410 (N_13410,N_13271,N_13295);
nand U13411 (N_13411,N_13291,N_13236);
xnor U13412 (N_13412,N_13334,N_13207);
or U13413 (N_13413,N_13325,N_13343);
nand U13414 (N_13414,N_13318,N_13284);
nor U13415 (N_13415,N_13220,N_13219);
or U13416 (N_13416,N_13212,N_13213);
or U13417 (N_13417,N_13338,N_13268);
and U13418 (N_13418,N_13348,N_13333);
nand U13419 (N_13419,N_13210,N_13240);
and U13420 (N_13420,N_13319,N_13280);
and U13421 (N_13421,N_13206,N_13255);
nand U13422 (N_13422,N_13208,N_13278);
or U13423 (N_13423,N_13223,N_13217);
and U13424 (N_13424,N_13346,N_13281);
and U13425 (N_13425,N_13348,N_13321);
and U13426 (N_13426,N_13332,N_13330);
and U13427 (N_13427,N_13313,N_13290);
nor U13428 (N_13428,N_13238,N_13245);
xor U13429 (N_13429,N_13299,N_13310);
and U13430 (N_13430,N_13347,N_13222);
xor U13431 (N_13431,N_13244,N_13219);
nand U13432 (N_13432,N_13239,N_13258);
and U13433 (N_13433,N_13330,N_13250);
nand U13434 (N_13434,N_13275,N_13231);
nor U13435 (N_13435,N_13280,N_13344);
nand U13436 (N_13436,N_13244,N_13281);
nor U13437 (N_13437,N_13255,N_13334);
and U13438 (N_13438,N_13276,N_13283);
xor U13439 (N_13439,N_13231,N_13294);
nor U13440 (N_13440,N_13233,N_13300);
or U13441 (N_13441,N_13263,N_13313);
nor U13442 (N_13442,N_13333,N_13323);
nor U13443 (N_13443,N_13306,N_13320);
xnor U13444 (N_13444,N_13349,N_13272);
and U13445 (N_13445,N_13280,N_13322);
xnor U13446 (N_13446,N_13289,N_13248);
and U13447 (N_13447,N_13228,N_13274);
or U13448 (N_13448,N_13314,N_13280);
or U13449 (N_13449,N_13245,N_13264);
and U13450 (N_13450,N_13327,N_13273);
nand U13451 (N_13451,N_13265,N_13347);
nor U13452 (N_13452,N_13334,N_13289);
nor U13453 (N_13453,N_13212,N_13320);
nand U13454 (N_13454,N_13343,N_13275);
nor U13455 (N_13455,N_13265,N_13246);
xnor U13456 (N_13456,N_13317,N_13328);
nand U13457 (N_13457,N_13249,N_13319);
nor U13458 (N_13458,N_13281,N_13217);
nand U13459 (N_13459,N_13255,N_13216);
or U13460 (N_13460,N_13202,N_13209);
nand U13461 (N_13461,N_13208,N_13201);
and U13462 (N_13462,N_13292,N_13336);
xnor U13463 (N_13463,N_13273,N_13321);
xor U13464 (N_13464,N_13293,N_13249);
nand U13465 (N_13465,N_13305,N_13343);
nand U13466 (N_13466,N_13286,N_13247);
nor U13467 (N_13467,N_13339,N_13333);
nand U13468 (N_13468,N_13308,N_13329);
and U13469 (N_13469,N_13236,N_13311);
nor U13470 (N_13470,N_13290,N_13317);
nor U13471 (N_13471,N_13238,N_13288);
or U13472 (N_13472,N_13288,N_13330);
or U13473 (N_13473,N_13305,N_13346);
nor U13474 (N_13474,N_13343,N_13330);
or U13475 (N_13475,N_13296,N_13280);
or U13476 (N_13476,N_13205,N_13329);
nand U13477 (N_13477,N_13211,N_13217);
xor U13478 (N_13478,N_13260,N_13325);
nor U13479 (N_13479,N_13202,N_13337);
nand U13480 (N_13480,N_13271,N_13286);
nand U13481 (N_13481,N_13338,N_13217);
or U13482 (N_13482,N_13291,N_13296);
nor U13483 (N_13483,N_13336,N_13210);
or U13484 (N_13484,N_13297,N_13233);
xor U13485 (N_13485,N_13215,N_13232);
or U13486 (N_13486,N_13283,N_13325);
nor U13487 (N_13487,N_13207,N_13231);
nand U13488 (N_13488,N_13312,N_13277);
nand U13489 (N_13489,N_13236,N_13300);
nor U13490 (N_13490,N_13342,N_13283);
and U13491 (N_13491,N_13214,N_13327);
nand U13492 (N_13492,N_13347,N_13238);
nand U13493 (N_13493,N_13292,N_13205);
or U13494 (N_13494,N_13323,N_13258);
xor U13495 (N_13495,N_13270,N_13291);
nor U13496 (N_13496,N_13305,N_13254);
nor U13497 (N_13497,N_13290,N_13325);
and U13498 (N_13498,N_13326,N_13292);
and U13499 (N_13499,N_13302,N_13280);
xor U13500 (N_13500,N_13474,N_13489);
and U13501 (N_13501,N_13463,N_13486);
and U13502 (N_13502,N_13453,N_13396);
or U13503 (N_13503,N_13446,N_13499);
and U13504 (N_13504,N_13424,N_13440);
nand U13505 (N_13505,N_13389,N_13401);
nand U13506 (N_13506,N_13471,N_13428);
nor U13507 (N_13507,N_13398,N_13400);
xnor U13508 (N_13508,N_13384,N_13448);
nor U13509 (N_13509,N_13394,N_13383);
and U13510 (N_13510,N_13481,N_13435);
or U13511 (N_13511,N_13455,N_13442);
xor U13512 (N_13512,N_13414,N_13483);
xor U13513 (N_13513,N_13487,N_13492);
nor U13514 (N_13514,N_13472,N_13377);
nor U13515 (N_13515,N_13498,N_13422);
and U13516 (N_13516,N_13452,N_13352);
nor U13517 (N_13517,N_13355,N_13477);
xor U13518 (N_13518,N_13399,N_13460);
and U13519 (N_13519,N_13393,N_13454);
nor U13520 (N_13520,N_13359,N_13470);
or U13521 (N_13521,N_13404,N_13370);
nor U13522 (N_13522,N_13386,N_13391);
nor U13523 (N_13523,N_13411,N_13485);
and U13524 (N_13524,N_13387,N_13430);
and U13525 (N_13525,N_13439,N_13368);
and U13526 (N_13526,N_13436,N_13479);
or U13527 (N_13527,N_13390,N_13350);
or U13528 (N_13528,N_13488,N_13365);
nand U13529 (N_13529,N_13409,N_13388);
and U13530 (N_13530,N_13433,N_13491);
or U13531 (N_13531,N_13497,N_13447);
xor U13532 (N_13532,N_13410,N_13438);
nand U13533 (N_13533,N_13403,N_13351);
or U13534 (N_13534,N_13372,N_13465);
nor U13535 (N_13535,N_13445,N_13364);
nor U13536 (N_13536,N_13379,N_13484);
nor U13537 (N_13537,N_13417,N_13407);
and U13538 (N_13538,N_13367,N_13434);
and U13539 (N_13539,N_13413,N_13462);
or U13540 (N_13540,N_13444,N_13361);
or U13541 (N_13541,N_13354,N_13419);
nor U13542 (N_13542,N_13397,N_13469);
nand U13543 (N_13543,N_13468,N_13353);
and U13544 (N_13544,N_13357,N_13380);
or U13545 (N_13545,N_13475,N_13362);
nand U13546 (N_13546,N_13405,N_13427);
nor U13547 (N_13547,N_13363,N_13443);
nor U13548 (N_13548,N_13418,N_13432);
and U13549 (N_13549,N_13423,N_13382);
nand U13550 (N_13550,N_13378,N_13385);
xnor U13551 (N_13551,N_13360,N_13369);
and U13552 (N_13552,N_13406,N_13358);
nand U13553 (N_13553,N_13429,N_13461);
or U13554 (N_13554,N_13457,N_13458);
or U13555 (N_13555,N_13421,N_13431);
nand U13556 (N_13556,N_13408,N_13426);
xnor U13557 (N_13557,N_13466,N_13482);
nand U13558 (N_13558,N_13459,N_13496);
or U13559 (N_13559,N_13425,N_13495);
nand U13560 (N_13560,N_13456,N_13494);
nor U13561 (N_13561,N_13366,N_13467);
and U13562 (N_13562,N_13450,N_13395);
and U13563 (N_13563,N_13356,N_13449);
xnor U13564 (N_13564,N_13437,N_13371);
nand U13565 (N_13565,N_13493,N_13476);
or U13566 (N_13566,N_13392,N_13464);
xor U13567 (N_13567,N_13374,N_13420);
nor U13568 (N_13568,N_13375,N_13412);
nand U13569 (N_13569,N_13381,N_13478);
nor U13570 (N_13570,N_13373,N_13490);
or U13571 (N_13571,N_13473,N_13376);
nand U13572 (N_13572,N_13415,N_13480);
nor U13573 (N_13573,N_13441,N_13416);
xnor U13574 (N_13574,N_13402,N_13451);
nor U13575 (N_13575,N_13478,N_13438);
xor U13576 (N_13576,N_13385,N_13372);
xor U13577 (N_13577,N_13390,N_13465);
nand U13578 (N_13578,N_13489,N_13350);
or U13579 (N_13579,N_13387,N_13476);
and U13580 (N_13580,N_13416,N_13390);
xnor U13581 (N_13581,N_13424,N_13388);
xor U13582 (N_13582,N_13462,N_13466);
nand U13583 (N_13583,N_13493,N_13431);
and U13584 (N_13584,N_13429,N_13365);
xnor U13585 (N_13585,N_13391,N_13448);
xnor U13586 (N_13586,N_13461,N_13372);
nor U13587 (N_13587,N_13375,N_13351);
nor U13588 (N_13588,N_13404,N_13449);
and U13589 (N_13589,N_13498,N_13461);
and U13590 (N_13590,N_13413,N_13355);
xnor U13591 (N_13591,N_13499,N_13368);
nand U13592 (N_13592,N_13490,N_13472);
nor U13593 (N_13593,N_13387,N_13477);
or U13594 (N_13594,N_13425,N_13366);
and U13595 (N_13595,N_13434,N_13483);
nand U13596 (N_13596,N_13361,N_13454);
nand U13597 (N_13597,N_13495,N_13435);
nor U13598 (N_13598,N_13364,N_13401);
nor U13599 (N_13599,N_13420,N_13463);
and U13600 (N_13600,N_13405,N_13358);
xor U13601 (N_13601,N_13377,N_13367);
or U13602 (N_13602,N_13385,N_13459);
nand U13603 (N_13603,N_13441,N_13356);
and U13604 (N_13604,N_13431,N_13435);
nor U13605 (N_13605,N_13453,N_13417);
nor U13606 (N_13606,N_13473,N_13350);
or U13607 (N_13607,N_13426,N_13377);
xnor U13608 (N_13608,N_13486,N_13395);
and U13609 (N_13609,N_13498,N_13399);
xor U13610 (N_13610,N_13419,N_13424);
xor U13611 (N_13611,N_13411,N_13495);
xnor U13612 (N_13612,N_13390,N_13381);
xor U13613 (N_13613,N_13384,N_13438);
nor U13614 (N_13614,N_13479,N_13463);
or U13615 (N_13615,N_13382,N_13498);
or U13616 (N_13616,N_13397,N_13375);
xor U13617 (N_13617,N_13390,N_13387);
and U13618 (N_13618,N_13476,N_13414);
xnor U13619 (N_13619,N_13387,N_13499);
xor U13620 (N_13620,N_13488,N_13466);
xor U13621 (N_13621,N_13403,N_13399);
nor U13622 (N_13622,N_13427,N_13491);
or U13623 (N_13623,N_13378,N_13492);
and U13624 (N_13624,N_13457,N_13424);
or U13625 (N_13625,N_13441,N_13398);
nand U13626 (N_13626,N_13496,N_13389);
nand U13627 (N_13627,N_13476,N_13468);
xnor U13628 (N_13628,N_13420,N_13361);
xnor U13629 (N_13629,N_13466,N_13472);
or U13630 (N_13630,N_13499,N_13420);
or U13631 (N_13631,N_13496,N_13406);
or U13632 (N_13632,N_13467,N_13466);
or U13633 (N_13633,N_13410,N_13489);
or U13634 (N_13634,N_13460,N_13456);
nor U13635 (N_13635,N_13497,N_13357);
nand U13636 (N_13636,N_13454,N_13473);
or U13637 (N_13637,N_13362,N_13361);
nor U13638 (N_13638,N_13449,N_13355);
nand U13639 (N_13639,N_13365,N_13399);
or U13640 (N_13640,N_13371,N_13469);
or U13641 (N_13641,N_13385,N_13397);
nor U13642 (N_13642,N_13352,N_13469);
or U13643 (N_13643,N_13384,N_13445);
and U13644 (N_13644,N_13372,N_13423);
and U13645 (N_13645,N_13359,N_13448);
nor U13646 (N_13646,N_13361,N_13441);
nor U13647 (N_13647,N_13459,N_13488);
and U13648 (N_13648,N_13443,N_13468);
or U13649 (N_13649,N_13467,N_13418);
nand U13650 (N_13650,N_13543,N_13639);
xnor U13651 (N_13651,N_13600,N_13615);
and U13652 (N_13652,N_13560,N_13568);
xnor U13653 (N_13653,N_13572,N_13637);
xor U13654 (N_13654,N_13588,N_13532);
and U13655 (N_13655,N_13565,N_13536);
nor U13656 (N_13656,N_13598,N_13576);
xor U13657 (N_13657,N_13601,N_13500);
nand U13658 (N_13658,N_13544,N_13566);
or U13659 (N_13659,N_13570,N_13592);
xor U13660 (N_13660,N_13623,N_13522);
nand U13661 (N_13661,N_13524,N_13552);
nor U13662 (N_13662,N_13642,N_13518);
nand U13663 (N_13663,N_13649,N_13527);
and U13664 (N_13664,N_13507,N_13562);
xnor U13665 (N_13665,N_13545,N_13614);
or U13666 (N_13666,N_13624,N_13627);
and U13667 (N_13667,N_13505,N_13547);
nor U13668 (N_13668,N_13534,N_13510);
or U13669 (N_13669,N_13550,N_13611);
and U13670 (N_13670,N_13533,N_13542);
or U13671 (N_13671,N_13525,N_13602);
nand U13672 (N_13672,N_13628,N_13573);
nor U13673 (N_13673,N_13634,N_13563);
nor U13674 (N_13674,N_13594,N_13553);
or U13675 (N_13675,N_13521,N_13513);
and U13676 (N_13676,N_13638,N_13535);
or U13677 (N_13677,N_13636,N_13559);
nor U13678 (N_13678,N_13583,N_13617);
and U13679 (N_13679,N_13515,N_13610);
and U13680 (N_13680,N_13564,N_13538);
and U13681 (N_13681,N_13540,N_13577);
and U13682 (N_13682,N_13620,N_13582);
nor U13683 (N_13683,N_13569,N_13643);
xor U13684 (N_13684,N_13506,N_13630);
nand U13685 (N_13685,N_13590,N_13539);
xnor U13686 (N_13686,N_13575,N_13580);
or U13687 (N_13687,N_13635,N_13604);
xnor U13688 (N_13688,N_13593,N_13551);
nor U13689 (N_13689,N_13523,N_13502);
or U13690 (N_13690,N_13585,N_13626);
nand U13691 (N_13691,N_13574,N_13501);
or U13692 (N_13692,N_13579,N_13520);
and U13693 (N_13693,N_13504,N_13607);
xor U13694 (N_13694,N_13609,N_13648);
xnor U13695 (N_13695,N_13586,N_13519);
nand U13696 (N_13696,N_13512,N_13616);
xnor U13697 (N_13697,N_13608,N_13644);
xor U13698 (N_13698,N_13541,N_13612);
and U13699 (N_13699,N_13549,N_13629);
xnor U13700 (N_13700,N_13625,N_13528);
or U13701 (N_13701,N_13595,N_13603);
and U13702 (N_13702,N_13647,N_13618);
or U13703 (N_13703,N_13621,N_13578);
and U13704 (N_13704,N_13599,N_13619);
xnor U13705 (N_13705,N_13555,N_13640);
or U13706 (N_13706,N_13587,N_13509);
nor U13707 (N_13707,N_13645,N_13546);
or U13708 (N_13708,N_13613,N_13508);
and U13709 (N_13709,N_13503,N_13537);
and U13710 (N_13710,N_13605,N_13633);
xnor U13711 (N_13711,N_13606,N_13557);
and U13712 (N_13712,N_13591,N_13526);
or U13713 (N_13713,N_13589,N_13558);
xor U13714 (N_13714,N_13517,N_13596);
or U13715 (N_13715,N_13631,N_13581);
xnor U13716 (N_13716,N_13531,N_13548);
and U13717 (N_13717,N_13511,N_13567);
and U13718 (N_13718,N_13571,N_13646);
nand U13719 (N_13719,N_13554,N_13622);
nor U13720 (N_13720,N_13530,N_13641);
or U13721 (N_13721,N_13561,N_13584);
and U13722 (N_13722,N_13632,N_13529);
and U13723 (N_13723,N_13556,N_13516);
and U13724 (N_13724,N_13514,N_13597);
and U13725 (N_13725,N_13520,N_13601);
and U13726 (N_13726,N_13586,N_13564);
xnor U13727 (N_13727,N_13609,N_13618);
or U13728 (N_13728,N_13515,N_13525);
nor U13729 (N_13729,N_13589,N_13510);
and U13730 (N_13730,N_13619,N_13552);
or U13731 (N_13731,N_13600,N_13559);
or U13732 (N_13732,N_13553,N_13555);
nand U13733 (N_13733,N_13522,N_13524);
xnor U13734 (N_13734,N_13613,N_13512);
nand U13735 (N_13735,N_13527,N_13610);
xor U13736 (N_13736,N_13576,N_13585);
or U13737 (N_13737,N_13596,N_13576);
and U13738 (N_13738,N_13598,N_13575);
xor U13739 (N_13739,N_13567,N_13639);
xor U13740 (N_13740,N_13594,N_13524);
or U13741 (N_13741,N_13515,N_13585);
nand U13742 (N_13742,N_13568,N_13623);
nor U13743 (N_13743,N_13507,N_13613);
and U13744 (N_13744,N_13628,N_13568);
or U13745 (N_13745,N_13628,N_13562);
xnor U13746 (N_13746,N_13500,N_13630);
and U13747 (N_13747,N_13646,N_13510);
nor U13748 (N_13748,N_13532,N_13634);
nor U13749 (N_13749,N_13628,N_13586);
xor U13750 (N_13750,N_13598,N_13604);
or U13751 (N_13751,N_13638,N_13607);
nor U13752 (N_13752,N_13556,N_13555);
xnor U13753 (N_13753,N_13639,N_13584);
nor U13754 (N_13754,N_13604,N_13501);
xor U13755 (N_13755,N_13594,N_13598);
and U13756 (N_13756,N_13594,N_13648);
or U13757 (N_13757,N_13574,N_13587);
nor U13758 (N_13758,N_13594,N_13557);
nor U13759 (N_13759,N_13513,N_13543);
xnor U13760 (N_13760,N_13516,N_13512);
nor U13761 (N_13761,N_13568,N_13624);
nand U13762 (N_13762,N_13540,N_13526);
nand U13763 (N_13763,N_13593,N_13544);
and U13764 (N_13764,N_13647,N_13626);
nor U13765 (N_13765,N_13580,N_13585);
and U13766 (N_13766,N_13617,N_13530);
xnor U13767 (N_13767,N_13574,N_13593);
xnor U13768 (N_13768,N_13556,N_13538);
nand U13769 (N_13769,N_13546,N_13519);
xnor U13770 (N_13770,N_13503,N_13613);
or U13771 (N_13771,N_13539,N_13626);
or U13772 (N_13772,N_13612,N_13533);
nor U13773 (N_13773,N_13525,N_13597);
nand U13774 (N_13774,N_13506,N_13593);
or U13775 (N_13775,N_13608,N_13537);
and U13776 (N_13776,N_13553,N_13595);
and U13777 (N_13777,N_13599,N_13516);
and U13778 (N_13778,N_13614,N_13638);
nor U13779 (N_13779,N_13613,N_13615);
nor U13780 (N_13780,N_13586,N_13566);
xor U13781 (N_13781,N_13574,N_13645);
xnor U13782 (N_13782,N_13573,N_13544);
and U13783 (N_13783,N_13521,N_13564);
or U13784 (N_13784,N_13545,N_13628);
nand U13785 (N_13785,N_13531,N_13634);
nand U13786 (N_13786,N_13566,N_13523);
nand U13787 (N_13787,N_13635,N_13526);
nor U13788 (N_13788,N_13624,N_13647);
or U13789 (N_13789,N_13572,N_13516);
nand U13790 (N_13790,N_13505,N_13589);
nand U13791 (N_13791,N_13577,N_13625);
nand U13792 (N_13792,N_13613,N_13609);
nor U13793 (N_13793,N_13573,N_13627);
or U13794 (N_13794,N_13548,N_13565);
xnor U13795 (N_13795,N_13567,N_13598);
or U13796 (N_13796,N_13619,N_13605);
and U13797 (N_13797,N_13536,N_13586);
xor U13798 (N_13798,N_13541,N_13628);
or U13799 (N_13799,N_13597,N_13626);
or U13800 (N_13800,N_13788,N_13703);
nand U13801 (N_13801,N_13682,N_13680);
or U13802 (N_13802,N_13796,N_13692);
and U13803 (N_13803,N_13717,N_13787);
nand U13804 (N_13804,N_13792,N_13661);
and U13805 (N_13805,N_13668,N_13666);
nor U13806 (N_13806,N_13707,N_13701);
nand U13807 (N_13807,N_13681,N_13718);
xor U13808 (N_13808,N_13657,N_13663);
nand U13809 (N_13809,N_13757,N_13704);
or U13810 (N_13810,N_13655,N_13695);
and U13811 (N_13811,N_13727,N_13764);
nor U13812 (N_13812,N_13784,N_13769);
or U13813 (N_13813,N_13786,N_13720);
or U13814 (N_13814,N_13674,N_13746);
nor U13815 (N_13815,N_13728,N_13650);
nand U13816 (N_13816,N_13712,N_13675);
and U13817 (N_13817,N_13689,N_13726);
nand U13818 (N_13818,N_13706,N_13740);
nor U13819 (N_13819,N_13658,N_13716);
nor U13820 (N_13820,N_13662,N_13710);
nor U13821 (N_13821,N_13795,N_13673);
nor U13822 (N_13822,N_13709,N_13799);
or U13823 (N_13823,N_13651,N_13794);
nand U13824 (N_13824,N_13761,N_13722);
or U13825 (N_13825,N_13763,N_13750);
or U13826 (N_13826,N_13711,N_13687);
and U13827 (N_13827,N_13659,N_13783);
or U13828 (N_13828,N_13653,N_13767);
xor U13829 (N_13829,N_13774,N_13694);
nand U13830 (N_13830,N_13729,N_13797);
and U13831 (N_13831,N_13789,N_13782);
or U13832 (N_13832,N_13672,N_13715);
nand U13833 (N_13833,N_13790,N_13777);
nand U13834 (N_13834,N_13739,N_13765);
nor U13835 (N_13835,N_13677,N_13768);
xnor U13836 (N_13836,N_13678,N_13691);
or U13837 (N_13837,N_13664,N_13676);
nor U13838 (N_13838,N_13702,N_13736);
and U13839 (N_13839,N_13766,N_13700);
xor U13840 (N_13840,N_13669,N_13679);
and U13841 (N_13841,N_13779,N_13798);
or U13842 (N_13842,N_13686,N_13770);
nor U13843 (N_13843,N_13697,N_13743);
nand U13844 (N_13844,N_13654,N_13721);
nand U13845 (N_13845,N_13771,N_13744);
and U13846 (N_13846,N_13785,N_13665);
xnor U13847 (N_13847,N_13749,N_13699);
nand U13848 (N_13848,N_13735,N_13754);
or U13849 (N_13849,N_13780,N_13742);
or U13850 (N_13850,N_13723,N_13688);
nor U13851 (N_13851,N_13747,N_13733);
xor U13852 (N_13852,N_13745,N_13652);
nor U13853 (N_13853,N_13683,N_13772);
nor U13854 (N_13854,N_13760,N_13753);
nand U13855 (N_13855,N_13684,N_13756);
and U13856 (N_13856,N_13708,N_13690);
and U13857 (N_13857,N_13781,N_13714);
nand U13858 (N_13858,N_13791,N_13696);
or U13859 (N_13859,N_13778,N_13775);
nor U13860 (N_13860,N_13734,N_13755);
or U13861 (N_13861,N_13713,N_13793);
nand U13862 (N_13862,N_13725,N_13773);
and U13863 (N_13863,N_13732,N_13748);
and U13864 (N_13864,N_13737,N_13667);
nand U13865 (N_13865,N_13741,N_13730);
or U13866 (N_13866,N_13685,N_13671);
nor U13867 (N_13867,N_13758,N_13724);
xnor U13868 (N_13868,N_13762,N_13759);
xor U13869 (N_13869,N_13776,N_13705);
and U13870 (N_13870,N_13693,N_13738);
nand U13871 (N_13871,N_13719,N_13751);
nand U13872 (N_13872,N_13752,N_13656);
or U13873 (N_13873,N_13698,N_13731);
nand U13874 (N_13874,N_13670,N_13660);
and U13875 (N_13875,N_13766,N_13724);
nand U13876 (N_13876,N_13665,N_13686);
or U13877 (N_13877,N_13795,N_13699);
and U13878 (N_13878,N_13666,N_13764);
nand U13879 (N_13879,N_13701,N_13658);
xor U13880 (N_13880,N_13777,N_13679);
or U13881 (N_13881,N_13682,N_13718);
and U13882 (N_13882,N_13753,N_13798);
nor U13883 (N_13883,N_13733,N_13727);
or U13884 (N_13884,N_13666,N_13704);
and U13885 (N_13885,N_13715,N_13724);
nand U13886 (N_13886,N_13687,N_13771);
and U13887 (N_13887,N_13730,N_13771);
or U13888 (N_13888,N_13758,N_13686);
nor U13889 (N_13889,N_13702,N_13717);
nand U13890 (N_13890,N_13779,N_13684);
xor U13891 (N_13891,N_13762,N_13670);
nor U13892 (N_13892,N_13665,N_13783);
nand U13893 (N_13893,N_13771,N_13656);
xnor U13894 (N_13894,N_13688,N_13736);
nand U13895 (N_13895,N_13742,N_13729);
nor U13896 (N_13896,N_13673,N_13719);
and U13897 (N_13897,N_13720,N_13727);
and U13898 (N_13898,N_13755,N_13783);
or U13899 (N_13899,N_13785,N_13769);
or U13900 (N_13900,N_13786,N_13797);
xor U13901 (N_13901,N_13735,N_13658);
xor U13902 (N_13902,N_13786,N_13676);
nand U13903 (N_13903,N_13665,N_13767);
or U13904 (N_13904,N_13745,N_13689);
nor U13905 (N_13905,N_13778,N_13743);
or U13906 (N_13906,N_13737,N_13666);
nor U13907 (N_13907,N_13796,N_13655);
nand U13908 (N_13908,N_13714,N_13738);
or U13909 (N_13909,N_13668,N_13681);
and U13910 (N_13910,N_13650,N_13737);
nand U13911 (N_13911,N_13683,N_13764);
or U13912 (N_13912,N_13670,N_13700);
or U13913 (N_13913,N_13688,N_13691);
xnor U13914 (N_13914,N_13677,N_13690);
nor U13915 (N_13915,N_13655,N_13776);
xor U13916 (N_13916,N_13674,N_13720);
nor U13917 (N_13917,N_13716,N_13798);
or U13918 (N_13918,N_13735,N_13652);
nand U13919 (N_13919,N_13660,N_13773);
xor U13920 (N_13920,N_13675,N_13780);
or U13921 (N_13921,N_13672,N_13652);
nand U13922 (N_13922,N_13774,N_13739);
nor U13923 (N_13923,N_13671,N_13651);
xor U13924 (N_13924,N_13793,N_13700);
nand U13925 (N_13925,N_13738,N_13773);
nand U13926 (N_13926,N_13681,N_13776);
nand U13927 (N_13927,N_13716,N_13714);
or U13928 (N_13928,N_13790,N_13733);
or U13929 (N_13929,N_13728,N_13794);
nor U13930 (N_13930,N_13751,N_13701);
nand U13931 (N_13931,N_13775,N_13782);
or U13932 (N_13932,N_13757,N_13726);
nor U13933 (N_13933,N_13653,N_13689);
or U13934 (N_13934,N_13766,N_13789);
nand U13935 (N_13935,N_13773,N_13731);
or U13936 (N_13936,N_13669,N_13776);
nor U13937 (N_13937,N_13659,N_13788);
nor U13938 (N_13938,N_13781,N_13712);
or U13939 (N_13939,N_13760,N_13684);
or U13940 (N_13940,N_13782,N_13797);
and U13941 (N_13941,N_13673,N_13761);
nand U13942 (N_13942,N_13653,N_13682);
or U13943 (N_13943,N_13729,N_13749);
and U13944 (N_13944,N_13759,N_13692);
and U13945 (N_13945,N_13682,N_13747);
nor U13946 (N_13946,N_13700,N_13704);
nor U13947 (N_13947,N_13702,N_13733);
xnor U13948 (N_13948,N_13717,N_13744);
nand U13949 (N_13949,N_13673,N_13715);
and U13950 (N_13950,N_13946,N_13820);
and U13951 (N_13951,N_13937,N_13849);
xnor U13952 (N_13952,N_13932,N_13845);
or U13953 (N_13953,N_13862,N_13826);
and U13954 (N_13954,N_13818,N_13843);
nand U13955 (N_13955,N_13856,N_13899);
xor U13956 (N_13956,N_13815,N_13854);
xnor U13957 (N_13957,N_13851,N_13915);
xnor U13958 (N_13958,N_13924,N_13900);
and U13959 (N_13959,N_13803,N_13922);
nor U13960 (N_13960,N_13887,N_13941);
and U13961 (N_13961,N_13920,N_13813);
nand U13962 (N_13962,N_13875,N_13864);
nor U13963 (N_13963,N_13945,N_13866);
xnor U13964 (N_13964,N_13858,N_13931);
or U13965 (N_13965,N_13800,N_13833);
nand U13966 (N_13966,N_13828,N_13810);
xnor U13967 (N_13967,N_13933,N_13916);
and U13968 (N_13968,N_13879,N_13872);
and U13969 (N_13969,N_13834,N_13919);
nand U13970 (N_13970,N_13906,N_13892);
or U13971 (N_13971,N_13901,N_13831);
and U13972 (N_13972,N_13801,N_13809);
and U13973 (N_13973,N_13830,N_13948);
or U13974 (N_13974,N_13921,N_13848);
or U13975 (N_13975,N_13897,N_13808);
or U13976 (N_13976,N_13832,N_13914);
or U13977 (N_13977,N_13827,N_13934);
xor U13978 (N_13978,N_13918,N_13877);
or U13979 (N_13979,N_13816,N_13838);
xor U13980 (N_13980,N_13861,N_13891);
or U13981 (N_13981,N_13909,N_13927);
and U13982 (N_13982,N_13942,N_13944);
or U13983 (N_13983,N_13853,N_13847);
and U13984 (N_13984,N_13926,N_13884);
xor U13985 (N_13985,N_13893,N_13902);
nand U13986 (N_13986,N_13860,N_13894);
or U13987 (N_13987,N_13855,N_13844);
nand U13988 (N_13988,N_13881,N_13850);
or U13989 (N_13989,N_13841,N_13913);
nand U13990 (N_13990,N_13928,N_13903);
and U13991 (N_13991,N_13859,N_13911);
or U13992 (N_13992,N_13867,N_13824);
nand U13993 (N_13993,N_13836,N_13837);
nor U13994 (N_13994,N_13938,N_13923);
nand U13995 (N_13995,N_13839,N_13822);
xor U13996 (N_13996,N_13806,N_13929);
xnor U13997 (N_13997,N_13873,N_13870);
nand U13998 (N_13998,N_13882,N_13817);
and U13999 (N_13999,N_13910,N_13852);
or U14000 (N_14000,N_13805,N_13888);
and U14001 (N_14001,N_13896,N_13874);
nand U14002 (N_14002,N_13819,N_13949);
xnor U14003 (N_14003,N_13804,N_13895);
or U14004 (N_14004,N_13883,N_13846);
and U14005 (N_14005,N_13823,N_13912);
nor U14006 (N_14006,N_13925,N_13886);
nor U14007 (N_14007,N_13936,N_13898);
or U14008 (N_14008,N_13940,N_13930);
and U14009 (N_14009,N_13876,N_13802);
nand U14010 (N_14010,N_13871,N_13869);
and U14011 (N_14011,N_13907,N_13829);
xnor U14012 (N_14012,N_13821,N_13890);
nand U14013 (N_14013,N_13917,N_13904);
and U14014 (N_14014,N_13825,N_13889);
nor U14015 (N_14015,N_13814,N_13835);
xnor U14016 (N_14016,N_13868,N_13811);
nor U14017 (N_14017,N_13863,N_13840);
or U14018 (N_14018,N_13865,N_13939);
or U14019 (N_14019,N_13812,N_13842);
or U14020 (N_14020,N_13857,N_13880);
nor U14021 (N_14021,N_13935,N_13905);
nor U14022 (N_14022,N_13943,N_13908);
or U14023 (N_14023,N_13885,N_13878);
nand U14024 (N_14024,N_13807,N_13947);
or U14025 (N_14025,N_13845,N_13897);
or U14026 (N_14026,N_13911,N_13845);
nand U14027 (N_14027,N_13924,N_13922);
nand U14028 (N_14028,N_13814,N_13908);
and U14029 (N_14029,N_13899,N_13864);
or U14030 (N_14030,N_13902,N_13872);
or U14031 (N_14031,N_13831,N_13812);
and U14032 (N_14032,N_13920,N_13800);
xor U14033 (N_14033,N_13858,N_13920);
or U14034 (N_14034,N_13828,N_13843);
xor U14035 (N_14035,N_13863,N_13814);
xor U14036 (N_14036,N_13844,N_13829);
xnor U14037 (N_14037,N_13809,N_13810);
nor U14038 (N_14038,N_13800,N_13939);
xnor U14039 (N_14039,N_13903,N_13830);
nand U14040 (N_14040,N_13898,N_13814);
xor U14041 (N_14041,N_13940,N_13816);
xnor U14042 (N_14042,N_13859,N_13873);
or U14043 (N_14043,N_13855,N_13851);
nand U14044 (N_14044,N_13870,N_13934);
nand U14045 (N_14045,N_13911,N_13828);
xnor U14046 (N_14046,N_13935,N_13923);
xnor U14047 (N_14047,N_13824,N_13833);
xor U14048 (N_14048,N_13884,N_13931);
or U14049 (N_14049,N_13864,N_13858);
xnor U14050 (N_14050,N_13828,N_13857);
xor U14051 (N_14051,N_13884,N_13923);
or U14052 (N_14052,N_13868,N_13923);
nand U14053 (N_14053,N_13889,N_13810);
xnor U14054 (N_14054,N_13944,N_13856);
nand U14055 (N_14055,N_13863,N_13912);
or U14056 (N_14056,N_13831,N_13846);
and U14057 (N_14057,N_13939,N_13935);
and U14058 (N_14058,N_13859,N_13825);
xnor U14059 (N_14059,N_13852,N_13829);
nor U14060 (N_14060,N_13939,N_13846);
xor U14061 (N_14061,N_13811,N_13815);
xnor U14062 (N_14062,N_13946,N_13886);
or U14063 (N_14063,N_13883,N_13910);
xnor U14064 (N_14064,N_13861,N_13914);
or U14065 (N_14065,N_13848,N_13816);
xor U14066 (N_14066,N_13830,N_13816);
or U14067 (N_14067,N_13804,N_13852);
nor U14068 (N_14068,N_13915,N_13881);
xor U14069 (N_14069,N_13889,N_13861);
xnor U14070 (N_14070,N_13830,N_13866);
xor U14071 (N_14071,N_13839,N_13825);
nand U14072 (N_14072,N_13809,N_13949);
or U14073 (N_14073,N_13908,N_13931);
and U14074 (N_14074,N_13860,N_13881);
xnor U14075 (N_14075,N_13893,N_13835);
nor U14076 (N_14076,N_13838,N_13804);
or U14077 (N_14077,N_13830,N_13845);
nand U14078 (N_14078,N_13855,N_13814);
nand U14079 (N_14079,N_13853,N_13895);
xnor U14080 (N_14080,N_13913,N_13805);
xor U14081 (N_14081,N_13916,N_13825);
nor U14082 (N_14082,N_13879,N_13920);
nand U14083 (N_14083,N_13830,N_13921);
nor U14084 (N_14084,N_13902,N_13905);
or U14085 (N_14085,N_13892,N_13939);
and U14086 (N_14086,N_13939,N_13856);
nand U14087 (N_14087,N_13940,N_13898);
and U14088 (N_14088,N_13870,N_13887);
or U14089 (N_14089,N_13866,N_13871);
nor U14090 (N_14090,N_13921,N_13929);
nand U14091 (N_14091,N_13945,N_13885);
and U14092 (N_14092,N_13928,N_13939);
and U14093 (N_14093,N_13855,N_13837);
nor U14094 (N_14094,N_13949,N_13896);
nand U14095 (N_14095,N_13903,N_13932);
nand U14096 (N_14096,N_13930,N_13915);
and U14097 (N_14097,N_13813,N_13850);
xor U14098 (N_14098,N_13884,N_13824);
and U14099 (N_14099,N_13853,N_13834);
xor U14100 (N_14100,N_14009,N_14024);
and U14101 (N_14101,N_14033,N_14010);
or U14102 (N_14102,N_13954,N_14028);
or U14103 (N_14103,N_14054,N_14053);
nand U14104 (N_14104,N_13970,N_14038);
nor U14105 (N_14105,N_14031,N_14015);
nor U14106 (N_14106,N_14044,N_13986);
and U14107 (N_14107,N_14037,N_14011);
nand U14108 (N_14108,N_14098,N_14089);
xnor U14109 (N_14109,N_14016,N_14055);
nand U14110 (N_14110,N_13990,N_14021);
xor U14111 (N_14111,N_13997,N_13963);
and U14112 (N_14112,N_14027,N_14062);
and U14113 (N_14113,N_14099,N_14070);
nand U14114 (N_14114,N_13965,N_13982);
or U14115 (N_14115,N_14094,N_14036);
or U14116 (N_14116,N_14046,N_14018);
xor U14117 (N_14117,N_14000,N_14014);
nand U14118 (N_14118,N_14085,N_14040);
nand U14119 (N_14119,N_14029,N_14050);
and U14120 (N_14120,N_14084,N_14096);
nand U14121 (N_14121,N_14082,N_14019);
or U14122 (N_14122,N_14090,N_14012);
xnor U14123 (N_14123,N_14013,N_13955);
nand U14124 (N_14124,N_14097,N_14049);
xor U14125 (N_14125,N_13979,N_14043);
xor U14126 (N_14126,N_14026,N_13996);
nand U14127 (N_14127,N_13995,N_14091);
nor U14128 (N_14128,N_14066,N_13981);
or U14129 (N_14129,N_13968,N_14079);
xor U14130 (N_14130,N_13972,N_14006);
nor U14131 (N_14131,N_13993,N_13989);
nand U14132 (N_14132,N_14039,N_14081);
xor U14133 (N_14133,N_13966,N_13998);
xor U14134 (N_14134,N_13967,N_13983);
nand U14135 (N_14135,N_14078,N_14063);
xor U14136 (N_14136,N_13962,N_14076);
and U14137 (N_14137,N_13959,N_13987);
xor U14138 (N_14138,N_14008,N_13953);
nor U14139 (N_14139,N_14072,N_14086);
xnor U14140 (N_14140,N_14005,N_13994);
xnor U14141 (N_14141,N_14032,N_14052);
or U14142 (N_14142,N_14022,N_13985);
xnor U14143 (N_14143,N_13992,N_14025);
nand U14144 (N_14144,N_14034,N_13971);
nand U14145 (N_14145,N_14064,N_14083);
nand U14146 (N_14146,N_13976,N_14020);
and U14147 (N_14147,N_13980,N_14060);
xnor U14148 (N_14148,N_13973,N_14001);
or U14149 (N_14149,N_14058,N_14023);
or U14150 (N_14150,N_14047,N_14007);
or U14151 (N_14151,N_14051,N_14059);
nand U14152 (N_14152,N_14095,N_13991);
xor U14153 (N_14153,N_14077,N_13977);
nand U14154 (N_14154,N_14068,N_13964);
nand U14155 (N_14155,N_13974,N_13984);
nor U14156 (N_14156,N_14087,N_13999);
nand U14157 (N_14157,N_14002,N_14074);
nand U14158 (N_14158,N_13957,N_13969);
or U14159 (N_14159,N_14030,N_14065);
nor U14160 (N_14160,N_14041,N_14004);
nand U14161 (N_14161,N_14045,N_14069);
xor U14162 (N_14162,N_14093,N_14056);
nor U14163 (N_14163,N_14067,N_13988);
nor U14164 (N_14164,N_14088,N_13952);
or U14165 (N_14165,N_13960,N_14071);
xnor U14166 (N_14166,N_14035,N_13961);
or U14167 (N_14167,N_14057,N_14092);
nor U14168 (N_14168,N_14017,N_13958);
nor U14169 (N_14169,N_14080,N_13951);
and U14170 (N_14170,N_14003,N_14048);
xor U14171 (N_14171,N_13950,N_13956);
and U14172 (N_14172,N_13978,N_14061);
xor U14173 (N_14173,N_13975,N_14042);
nand U14174 (N_14174,N_14075,N_14073);
nand U14175 (N_14175,N_14025,N_14098);
xnor U14176 (N_14176,N_13959,N_13989);
nand U14177 (N_14177,N_14076,N_14060);
and U14178 (N_14178,N_13966,N_14058);
and U14179 (N_14179,N_14072,N_13991);
xor U14180 (N_14180,N_13993,N_14040);
and U14181 (N_14181,N_14048,N_14092);
or U14182 (N_14182,N_14024,N_13998);
nand U14183 (N_14183,N_14058,N_13961);
nand U14184 (N_14184,N_13959,N_14033);
and U14185 (N_14185,N_14099,N_14075);
nor U14186 (N_14186,N_13980,N_14056);
nor U14187 (N_14187,N_14001,N_13966);
nand U14188 (N_14188,N_14022,N_14048);
or U14189 (N_14189,N_13996,N_13976);
nand U14190 (N_14190,N_14016,N_13971);
nor U14191 (N_14191,N_14098,N_14047);
nor U14192 (N_14192,N_14093,N_13960);
nor U14193 (N_14193,N_13972,N_14056);
or U14194 (N_14194,N_13978,N_14031);
nand U14195 (N_14195,N_13997,N_14022);
and U14196 (N_14196,N_13966,N_14048);
nor U14197 (N_14197,N_13991,N_14040);
or U14198 (N_14198,N_14031,N_14054);
xor U14199 (N_14199,N_14037,N_13958);
nand U14200 (N_14200,N_14095,N_14035);
and U14201 (N_14201,N_13999,N_14039);
nor U14202 (N_14202,N_14057,N_14059);
xnor U14203 (N_14203,N_13954,N_13994);
and U14204 (N_14204,N_14008,N_14009);
and U14205 (N_14205,N_14095,N_13989);
nor U14206 (N_14206,N_14096,N_13999);
or U14207 (N_14207,N_13987,N_14095);
or U14208 (N_14208,N_14018,N_13955);
xnor U14209 (N_14209,N_14080,N_13966);
nand U14210 (N_14210,N_13962,N_14053);
and U14211 (N_14211,N_14071,N_13956);
and U14212 (N_14212,N_13967,N_13978);
and U14213 (N_14213,N_13990,N_13965);
or U14214 (N_14214,N_14031,N_14065);
and U14215 (N_14215,N_14029,N_14082);
nor U14216 (N_14216,N_14040,N_14049);
nand U14217 (N_14217,N_13966,N_13950);
nor U14218 (N_14218,N_14026,N_14017);
xnor U14219 (N_14219,N_14043,N_13973);
nand U14220 (N_14220,N_14015,N_14007);
xor U14221 (N_14221,N_14077,N_14012);
nand U14222 (N_14222,N_14081,N_14029);
and U14223 (N_14223,N_14090,N_14077);
or U14224 (N_14224,N_14027,N_14055);
nor U14225 (N_14225,N_14013,N_14092);
xor U14226 (N_14226,N_14003,N_14043);
and U14227 (N_14227,N_14096,N_13976);
and U14228 (N_14228,N_13986,N_14053);
xnor U14229 (N_14229,N_13995,N_14062);
nor U14230 (N_14230,N_14089,N_14094);
nand U14231 (N_14231,N_13952,N_13994);
xnor U14232 (N_14232,N_13963,N_14036);
and U14233 (N_14233,N_14039,N_14098);
or U14234 (N_14234,N_13956,N_13957);
nor U14235 (N_14235,N_14051,N_14096);
or U14236 (N_14236,N_13965,N_14059);
nand U14237 (N_14237,N_13951,N_14077);
or U14238 (N_14238,N_14049,N_14034);
and U14239 (N_14239,N_14044,N_13990);
nor U14240 (N_14240,N_13960,N_13991);
xnor U14241 (N_14241,N_14049,N_14082);
or U14242 (N_14242,N_14042,N_14061);
or U14243 (N_14243,N_14043,N_13959);
or U14244 (N_14244,N_14024,N_14060);
and U14245 (N_14245,N_13974,N_14080);
and U14246 (N_14246,N_14087,N_13975);
or U14247 (N_14247,N_14017,N_14086);
nand U14248 (N_14248,N_13962,N_13987);
or U14249 (N_14249,N_14032,N_14095);
or U14250 (N_14250,N_14245,N_14238);
and U14251 (N_14251,N_14186,N_14220);
or U14252 (N_14252,N_14115,N_14169);
nor U14253 (N_14253,N_14164,N_14226);
or U14254 (N_14254,N_14204,N_14193);
or U14255 (N_14255,N_14249,N_14235);
nand U14256 (N_14256,N_14113,N_14131);
nand U14257 (N_14257,N_14111,N_14213);
and U14258 (N_14258,N_14130,N_14221);
nand U14259 (N_14259,N_14228,N_14158);
and U14260 (N_14260,N_14241,N_14152);
xor U14261 (N_14261,N_14244,N_14151);
xnor U14262 (N_14262,N_14168,N_14108);
or U14263 (N_14263,N_14248,N_14137);
and U14264 (N_14264,N_14148,N_14163);
nand U14265 (N_14265,N_14142,N_14135);
nand U14266 (N_14266,N_14196,N_14246);
xnor U14267 (N_14267,N_14106,N_14211);
and U14268 (N_14268,N_14160,N_14149);
and U14269 (N_14269,N_14140,N_14145);
and U14270 (N_14270,N_14105,N_14179);
xor U14271 (N_14271,N_14155,N_14147);
and U14272 (N_14272,N_14236,N_14205);
or U14273 (N_14273,N_14206,N_14170);
nand U14274 (N_14274,N_14119,N_14100);
xnor U14275 (N_14275,N_14132,N_14219);
or U14276 (N_14276,N_14188,N_14172);
nand U14277 (N_14277,N_14102,N_14185);
nand U14278 (N_14278,N_14209,N_14203);
and U14279 (N_14279,N_14109,N_14187);
xnor U14280 (N_14280,N_14165,N_14167);
nand U14281 (N_14281,N_14150,N_14194);
or U14282 (N_14282,N_14227,N_14190);
or U14283 (N_14283,N_14240,N_14138);
nor U14284 (N_14284,N_14153,N_14200);
or U14285 (N_14285,N_14133,N_14175);
xor U14286 (N_14286,N_14184,N_14117);
xnor U14287 (N_14287,N_14129,N_14210);
and U14288 (N_14288,N_14122,N_14217);
and U14289 (N_14289,N_14141,N_14197);
xor U14290 (N_14290,N_14139,N_14191);
nand U14291 (N_14291,N_14237,N_14178);
and U14292 (N_14292,N_14114,N_14201);
xnor U14293 (N_14293,N_14216,N_14181);
nor U14294 (N_14294,N_14177,N_14192);
xor U14295 (N_14295,N_14128,N_14173);
and U14296 (N_14296,N_14247,N_14162);
or U14297 (N_14297,N_14159,N_14208);
nand U14298 (N_14298,N_14127,N_14234);
nand U14299 (N_14299,N_14223,N_14230);
or U14300 (N_14300,N_14154,N_14157);
xor U14301 (N_14301,N_14224,N_14104);
xor U14302 (N_14302,N_14218,N_14120);
xor U14303 (N_14303,N_14225,N_14123);
xor U14304 (N_14304,N_14182,N_14195);
or U14305 (N_14305,N_14124,N_14166);
or U14306 (N_14306,N_14161,N_14125);
or U14307 (N_14307,N_14174,N_14118);
and U14308 (N_14308,N_14136,N_14180);
xnor U14309 (N_14309,N_14229,N_14222);
nor U14310 (N_14310,N_14107,N_14176);
or U14311 (N_14311,N_14189,N_14215);
and U14312 (N_14312,N_14110,N_14243);
nor U14313 (N_14313,N_14144,N_14232);
xor U14314 (N_14314,N_14198,N_14156);
or U14315 (N_14315,N_14214,N_14126);
xnor U14316 (N_14316,N_14207,N_14212);
xor U14317 (N_14317,N_14231,N_14112);
or U14318 (N_14318,N_14171,N_14101);
xnor U14319 (N_14319,N_14202,N_14242);
and U14320 (N_14320,N_14183,N_14143);
or U14321 (N_14321,N_14116,N_14233);
xnor U14322 (N_14322,N_14199,N_14239);
nor U14323 (N_14323,N_14121,N_14146);
and U14324 (N_14324,N_14103,N_14134);
and U14325 (N_14325,N_14105,N_14164);
nor U14326 (N_14326,N_14176,N_14127);
or U14327 (N_14327,N_14194,N_14134);
or U14328 (N_14328,N_14201,N_14120);
xor U14329 (N_14329,N_14239,N_14163);
nor U14330 (N_14330,N_14160,N_14170);
and U14331 (N_14331,N_14105,N_14200);
nand U14332 (N_14332,N_14135,N_14140);
nand U14333 (N_14333,N_14212,N_14127);
and U14334 (N_14334,N_14244,N_14197);
nand U14335 (N_14335,N_14132,N_14175);
and U14336 (N_14336,N_14236,N_14208);
nor U14337 (N_14337,N_14249,N_14215);
or U14338 (N_14338,N_14152,N_14105);
and U14339 (N_14339,N_14133,N_14193);
xnor U14340 (N_14340,N_14211,N_14138);
nand U14341 (N_14341,N_14125,N_14128);
or U14342 (N_14342,N_14175,N_14118);
nor U14343 (N_14343,N_14109,N_14108);
xor U14344 (N_14344,N_14110,N_14177);
and U14345 (N_14345,N_14229,N_14125);
nand U14346 (N_14346,N_14241,N_14238);
xor U14347 (N_14347,N_14114,N_14130);
xnor U14348 (N_14348,N_14158,N_14138);
and U14349 (N_14349,N_14194,N_14239);
or U14350 (N_14350,N_14231,N_14179);
nand U14351 (N_14351,N_14183,N_14155);
nand U14352 (N_14352,N_14124,N_14223);
or U14353 (N_14353,N_14233,N_14190);
or U14354 (N_14354,N_14213,N_14135);
xnor U14355 (N_14355,N_14245,N_14162);
xor U14356 (N_14356,N_14169,N_14127);
and U14357 (N_14357,N_14221,N_14139);
nor U14358 (N_14358,N_14183,N_14236);
nand U14359 (N_14359,N_14211,N_14154);
nor U14360 (N_14360,N_14230,N_14191);
or U14361 (N_14361,N_14213,N_14160);
xnor U14362 (N_14362,N_14182,N_14178);
nor U14363 (N_14363,N_14161,N_14133);
and U14364 (N_14364,N_14229,N_14195);
xor U14365 (N_14365,N_14125,N_14179);
or U14366 (N_14366,N_14132,N_14138);
nand U14367 (N_14367,N_14238,N_14147);
nor U14368 (N_14368,N_14176,N_14179);
xor U14369 (N_14369,N_14201,N_14110);
and U14370 (N_14370,N_14124,N_14208);
nor U14371 (N_14371,N_14135,N_14155);
or U14372 (N_14372,N_14232,N_14184);
or U14373 (N_14373,N_14228,N_14176);
nor U14374 (N_14374,N_14107,N_14120);
nand U14375 (N_14375,N_14212,N_14239);
and U14376 (N_14376,N_14203,N_14137);
nor U14377 (N_14377,N_14171,N_14211);
nand U14378 (N_14378,N_14165,N_14236);
and U14379 (N_14379,N_14134,N_14110);
or U14380 (N_14380,N_14228,N_14153);
nor U14381 (N_14381,N_14205,N_14179);
xor U14382 (N_14382,N_14242,N_14106);
xnor U14383 (N_14383,N_14114,N_14211);
nand U14384 (N_14384,N_14140,N_14124);
xor U14385 (N_14385,N_14184,N_14134);
nand U14386 (N_14386,N_14100,N_14207);
and U14387 (N_14387,N_14194,N_14117);
xnor U14388 (N_14388,N_14246,N_14101);
and U14389 (N_14389,N_14150,N_14206);
nand U14390 (N_14390,N_14210,N_14209);
xnor U14391 (N_14391,N_14176,N_14177);
xor U14392 (N_14392,N_14209,N_14220);
or U14393 (N_14393,N_14246,N_14231);
xor U14394 (N_14394,N_14191,N_14228);
and U14395 (N_14395,N_14124,N_14100);
xor U14396 (N_14396,N_14146,N_14174);
nand U14397 (N_14397,N_14183,N_14139);
nand U14398 (N_14398,N_14122,N_14170);
nand U14399 (N_14399,N_14187,N_14196);
nand U14400 (N_14400,N_14367,N_14355);
nor U14401 (N_14401,N_14298,N_14309);
nand U14402 (N_14402,N_14264,N_14361);
nand U14403 (N_14403,N_14273,N_14344);
nor U14404 (N_14404,N_14349,N_14313);
nand U14405 (N_14405,N_14323,N_14319);
and U14406 (N_14406,N_14254,N_14320);
xnor U14407 (N_14407,N_14272,N_14389);
nor U14408 (N_14408,N_14281,N_14270);
xnor U14409 (N_14409,N_14336,N_14398);
xnor U14410 (N_14410,N_14373,N_14311);
nand U14411 (N_14411,N_14283,N_14292);
nand U14412 (N_14412,N_14370,N_14382);
nand U14413 (N_14413,N_14315,N_14326);
nor U14414 (N_14414,N_14258,N_14275);
xor U14415 (N_14415,N_14364,N_14280);
nor U14416 (N_14416,N_14377,N_14286);
nor U14417 (N_14417,N_14356,N_14288);
nor U14418 (N_14418,N_14337,N_14322);
xor U14419 (N_14419,N_14329,N_14372);
or U14420 (N_14420,N_14385,N_14274);
and U14421 (N_14421,N_14331,N_14278);
and U14422 (N_14422,N_14251,N_14363);
or U14423 (N_14423,N_14332,N_14334);
nor U14424 (N_14424,N_14257,N_14348);
nor U14425 (N_14425,N_14330,N_14396);
or U14426 (N_14426,N_14339,N_14289);
or U14427 (N_14427,N_14267,N_14342);
or U14428 (N_14428,N_14276,N_14386);
xor U14429 (N_14429,N_14345,N_14265);
and U14430 (N_14430,N_14271,N_14358);
nor U14431 (N_14431,N_14378,N_14287);
nand U14432 (N_14432,N_14296,N_14293);
nor U14433 (N_14433,N_14362,N_14302);
nor U14434 (N_14434,N_14335,N_14261);
xnor U14435 (N_14435,N_14327,N_14317);
and U14436 (N_14436,N_14250,N_14253);
nor U14437 (N_14437,N_14266,N_14365);
nand U14438 (N_14438,N_14294,N_14290);
xor U14439 (N_14439,N_14325,N_14353);
nand U14440 (N_14440,N_14310,N_14384);
xor U14441 (N_14441,N_14369,N_14381);
nor U14442 (N_14442,N_14341,N_14395);
nand U14443 (N_14443,N_14383,N_14374);
nor U14444 (N_14444,N_14295,N_14368);
or U14445 (N_14445,N_14291,N_14262);
nor U14446 (N_14446,N_14379,N_14387);
nor U14447 (N_14447,N_14376,N_14360);
nor U14448 (N_14448,N_14340,N_14259);
nand U14449 (N_14449,N_14333,N_14391);
xor U14450 (N_14450,N_14350,N_14297);
and U14451 (N_14451,N_14397,N_14307);
or U14452 (N_14452,N_14359,N_14343);
and U14453 (N_14453,N_14279,N_14366);
nor U14454 (N_14454,N_14256,N_14346);
nor U14455 (N_14455,N_14388,N_14312);
nand U14456 (N_14456,N_14371,N_14347);
or U14457 (N_14457,N_14393,N_14380);
or U14458 (N_14458,N_14268,N_14354);
nand U14459 (N_14459,N_14263,N_14352);
xor U14460 (N_14460,N_14390,N_14306);
nor U14461 (N_14461,N_14316,N_14277);
xor U14462 (N_14462,N_14285,N_14318);
nand U14463 (N_14463,N_14300,N_14314);
or U14464 (N_14464,N_14351,N_14338);
nor U14465 (N_14465,N_14255,N_14301);
nand U14466 (N_14466,N_14284,N_14357);
or U14467 (N_14467,N_14303,N_14304);
xnor U14468 (N_14468,N_14305,N_14321);
nand U14469 (N_14469,N_14260,N_14308);
or U14470 (N_14470,N_14399,N_14394);
nand U14471 (N_14471,N_14299,N_14328);
and U14472 (N_14472,N_14392,N_14252);
and U14473 (N_14473,N_14324,N_14269);
xor U14474 (N_14474,N_14375,N_14282);
xor U14475 (N_14475,N_14317,N_14362);
xnor U14476 (N_14476,N_14360,N_14280);
and U14477 (N_14477,N_14346,N_14292);
xnor U14478 (N_14478,N_14381,N_14356);
and U14479 (N_14479,N_14271,N_14326);
xnor U14480 (N_14480,N_14269,N_14252);
nand U14481 (N_14481,N_14348,N_14371);
xnor U14482 (N_14482,N_14263,N_14270);
xnor U14483 (N_14483,N_14364,N_14373);
nor U14484 (N_14484,N_14270,N_14254);
or U14485 (N_14485,N_14257,N_14366);
nand U14486 (N_14486,N_14262,N_14253);
nor U14487 (N_14487,N_14357,N_14305);
or U14488 (N_14488,N_14290,N_14381);
xnor U14489 (N_14489,N_14345,N_14299);
nand U14490 (N_14490,N_14349,N_14354);
nand U14491 (N_14491,N_14365,N_14339);
and U14492 (N_14492,N_14284,N_14278);
xor U14493 (N_14493,N_14262,N_14318);
or U14494 (N_14494,N_14260,N_14364);
and U14495 (N_14495,N_14275,N_14372);
nor U14496 (N_14496,N_14321,N_14363);
and U14497 (N_14497,N_14325,N_14277);
or U14498 (N_14498,N_14276,N_14271);
or U14499 (N_14499,N_14351,N_14315);
and U14500 (N_14500,N_14378,N_14390);
xor U14501 (N_14501,N_14328,N_14396);
nor U14502 (N_14502,N_14337,N_14365);
and U14503 (N_14503,N_14360,N_14322);
nor U14504 (N_14504,N_14305,N_14257);
xor U14505 (N_14505,N_14309,N_14361);
xnor U14506 (N_14506,N_14316,N_14341);
and U14507 (N_14507,N_14260,N_14283);
xnor U14508 (N_14508,N_14354,N_14337);
or U14509 (N_14509,N_14367,N_14325);
xnor U14510 (N_14510,N_14369,N_14265);
or U14511 (N_14511,N_14304,N_14367);
nand U14512 (N_14512,N_14262,N_14365);
nor U14513 (N_14513,N_14345,N_14310);
xnor U14514 (N_14514,N_14261,N_14284);
nand U14515 (N_14515,N_14386,N_14395);
or U14516 (N_14516,N_14395,N_14311);
and U14517 (N_14517,N_14315,N_14343);
nor U14518 (N_14518,N_14352,N_14312);
or U14519 (N_14519,N_14395,N_14252);
and U14520 (N_14520,N_14396,N_14302);
or U14521 (N_14521,N_14381,N_14392);
nand U14522 (N_14522,N_14276,N_14367);
and U14523 (N_14523,N_14339,N_14265);
nand U14524 (N_14524,N_14277,N_14321);
xor U14525 (N_14525,N_14323,N_14327);
nand U14526 (N_14526,N_14338,N_14350);
or U14527 (N_14527,N_14356,N_14375);
nor U14528 (N_14528,N_14302,N_14342);
nand U14529 (N_14529,N_14373,N_14320);
nor U14530 (N_14530,N_14306,N_14264);
and U14531 (N_14531,N_14349,N_14389);
xor U14532 (N_14532,N_14338,N_14256);
nor U14533 (N_14533,N_14336,N_14389);
xnor U14534 (N_14534,N_14288,N_14258);
or U14535 (N_14535,N_14279,N_14397);
or U14536 (N_14536,N_14355,N_14381);
nand U14537 (N_14537,N_14379,N_14344);
nand U14538 (N_14538,N_14268,N_14270);
nor U14539 (N_14539,N_14354,N_14280);
nor U14540 (N_14540,N_14305,N_14302);
and U14541 (N_14541,N_14280,N_14373);
and U14542 (N_14542,N_14270,N_14269);
nor U14543 (N_14543,N_14330,N_14372);
nor U14544 (N_14544,N_14266,N_14372);
or U14545 (N_14545,N_14355,N_14351);
and U14546 (N_14546,N_14393,N_14277);
nor U14547 (N_14547,N_14302,N_14325);
xnor U14548 (N_14548,N_14310,N_14333);
and U14549 (N_14549,N_14277,N_14326);
xor U14550 (N_14550,N_14414,N_14459);
xnor U14551 (N_14551,N_14443,N_14436);
or U14552 (N_14552,N_14489,N_14471);
xor U14553 (N_14553,N_14449,N_14522);
or U14554 (N_14554,N_14539,N_14476);
xnor U14555 (N_14555,N_14432,N_14485);
xnor U14556 (N_14556,N_14492,N_14447);
xor U14557 (N_14557,N_14525,N_14517);
or U14558 (N_14558,N_14509,N_14502);
and U14559 (N_14559,N_14543,N_14411);
nor U14560 (N_14560,N_14452,N_14475);
nor U14561 (N_14561,N_14435,N_14453);
nand U14562 (N_14562,N_14526,N_14501);
nor U14563 (N_14563,N_14505,N_14477);
or U14564 (N_14564,N_14513,N_14470);
and U14565 (N_14565,N_14491,N_14472);
nand U14566 (N_14566,N_14402,N_14404);
and U14567 (N_14567,N_14512,N_14407);
nand U14568 (N_14568,N_14507,N_14544);
and U14569 (N_14569,N_14523,N_14425);
nand U14570 (N_14570,N_14483,N_14403);
xor U14571 (N_14571,N_14429,N_14454);
xnor U14572 (N_14572,N_14417,N_14531);
nand U14573 (N_14573,N_14487,N_14548);
nand U14574 (N_14574,N_14540,N_14442);
or U14575 (N_14575,N_14529,N_14545);
xor U14576 (N_14576,N_14437,N_14457);
nor U14577 (N_14577,N_14479,N_14467);
and U14578 (N_14578,N_14445,N_14520);
xor U14579 (N_14579,N_14474,N_14500);
nor U14580 (N_14580,N_14463,N_14532);
xor U14581 (N_14581,N_14462,N_14418);
nor U14582 (N_14582,N_14516,N_14537);
nand U14583 (N_14583,N_14515,N_14521);
and U14584 (N_14584,N_14469,N_14541);
or U14585 (N_14585,N_14519,N_14488);
or U14586 (N_14586,N_14496,N_14480);
nor U14587 (N_14587,N_14460,N_14466);
and U14588 (N_14588,N_14450,N_14546);
xnor U14589 (N_14589,N_14508,N_14433);
nand U14590 (N_14590,N_14497,N_14494);
nand U14591 (N_14591,N_14503,N_14518);
nand U14592 (N_14592,N_14536,N_14444);
or U14593 (N_14593,N_14538,N_14455);
nand U14594 (N_14594,N_14419,N_14416);
or U14595 (N_14595,N_14439,N_14511);
nor U14596 (N_14596,N_14448,N_14498);
or U14597 (N_14597,N_14401,N_14451);
and U14598 (N_14598,N_14547,N_14506);
nand U14599 (N_14599,N_14431,N_14528);
nand U14600 (N_14600,N_14421,N_14461);
or U14601 (N_14601,N_14456,N_14504);
nand U14602 (N_14602,N_14533,N_14468);
nor U14603 (N_14603,N_14410,N_14400);
xnor U14604 (N_14604,N_14482,N_14486);
or U14605 (N_14605,N_14413,N_14420);
xnor U14606 (N_14606,N_14542,N_14423);
and U14607 (N_14607,N_14434,N_14490);
xor U14608 (N_14608,N_14481,N_14415);
or U14609 (N_14609,N_14530,N_14412);
or U14610 (N_14610,N_14495,N_14422);
nand U14611 (N_14611,N_14424,N_14427);
nand U14612 (N_14612,N_14438,N_14493);
and U14613 (N_14613,N_14535,N_14430);
xor U14614 (N_14614,N_14473,N_14405);
or U14615 (N_14615,N_14408,N_14441);
and U14616 (N_14616,N_14409,N_14426);
or U14617 (N_14617,N_14524,N_14510);
nor U14618 (N_14618,N_14484,N_14478);
and U14619 (N_14619,N_14527,N_14406);
xor U14620 (N_14620,N_14499,N_14446);
or U14621 (N_14621,N_14458,N_14549);
or U14622 (N_14622,N_14514,N_14534);
and U14623 (N_14623,N_14465,N_14440);
nor U14624 (N_14624,N_14428,N_14464);
nor U14625 (N_14625,N_14501,N_14469);
xnor U14626 (N_14626,N_14476,N_14526);
or U14627 (N_14627,N_14500,N_14443);
or U14628 (N_14628,N_14431,N_14508);
or U14629 (N_14629,N_14448,N_14438);
nand U14630 (N_14630,N_14457,N_14511);
or U14631 (N_14631,N_14479,N_14486);
nand U14632 (N_14632,N_14423,N_14443);
or U14633 (N_14633,N_14490,N_14405);
nor U14634 (N_14634,N_14415,N_14435);
xor U14635 (N_14635,N_14532,N_14540);
nand U14636 (N_14636,N_14402,N_14462);
or U14637 (N_14637,N_14471,N_14530);
nor U14638 (N_14638,N_14491,N_14539);
and U14639 (N_14639,N_14425,N_14405);
and U14640 (N_14640,N_14521,N_14407);
xor U14641 (N_14641,N_14518,N_14455);
and U14642 (N_14642,N_14405,N_14427);
nand U14643 (N_14643,N_14548,N_14537);
or U14644 (N_14644,N_14403,N_14519);
xnor U14645 (N_14645,N_14538,N_14542);
nand U14646 (N_14646,N_14434,N_14405);
or U14647 (N_14647,N_14513,N_14437);
nand U14648 (N_14648,N_14507,N_14450);
nand U14649 (N_14649,N_14483,N_14533);
or U14650 (N_14650,N_14472,N_14521);
xor U14651 (N_14651,N_14540,N_14446);
and U14652 (N_14652,N_14466,N_14410);
nand U14653 (N_14653,N_14440,N_14470);
nor U14654 (N_14654,N_14532,N_14497);
and U14655 (N_14655,N_14443,N_14502);
or U14656 (N_14656,N_14468,N_14426);
and U14657 (N_14657,N_14519,N_14466);
nand U14658 (N_14658,N_14439,N_14536);
nor U14659 (N_14659,N_14521,N_14506);
or U14660 (N_14660,N_14425,N_14516);
xor U14661 (N_14661,N_14435,N_14494);
nand U14662 (N_14662,N_14506,N_14486);
xor U14663 (N_14663,N_14518,N_14487);
nor U14664 (N_14664,N_14436,N_14468);
and U14665 (N_14665,N_14452,N_14474);
xor U14666 (N_14666,N_14492,N_14480);
and U14667 (N_14667,N_14463,N_14437);
xnor U14668 (N_14668,N_14431,N_14430);
xor U14669 (N_14669,N_14430,N_14417);
nor U14670 (N_14670,N_14436,N_14464);
and U14671 (N_14671,N_14538,N_14522);
xnor U14672 (N_14672,N_14430,N_14465);
and U14673 (N_14673,N_14449,N_14466);
nand U14674 (N_14674,N_14403,N_14477);
nand U14675 (N_14675,N_14406,N_14549);
nand U14676 (N_14676,N_14528,N_14416);
xnor U14677 (N_14677,N_14538,N_14480);
or U14678 (N_14678,N_14546,N_14504);
or U14679 (N_14679,N_14481,N_14513);
or U14680 (N_14680,N_14447,N_14486);
xnor U14681 (N_14681,N_14457,N_14549);
nor U14682 (N_14682,N_14433,N_14464);
xor U14683 (N_14683,N_14404,N_14473);
or U14684 (N_14684,N_14420,N_14407);
and U14685 (N_14685,N_14429,N_14500);
nand U14686 (N_14686,N_14535,N_14528);
xor U14687 (N_14687,N_14508,N_14520);
and U14688 (N_14688,N_14539,N_14501);
nand U14689 (N_14689,N_14492,N_14478);
nand U14690 (N_14690,N_14417,N_14440);
or U14691 (N_14691,N_14442,N_14479);
nand U14692 (N_14692,N_14514,N_14465);
xnor U14693 (N_14693,N_14444,N_14422);
and U14694 (N_14694,N_14481,N_14456);
and U14695 (N_14695,N_14440,N_14405);
and U14696 (N_14696,N_14466,N_14451);
or U14697 (N_14697,N_14513,N_14512);
xor U14698 (N_14698,N_14519,N_14460);
nor U14699 (N_14699,N_14496,N_14440);
xor U14700 (N_14700,N_14680,N_14681);
xor U14701 (N_14701,N_14655,N_14582);
or U14702 (N_14702,N_14672,N_14640);
and U14703 (N_14703,N_14561,N_14650);
or U14704 (N_14704,N_14669,N_14563);
xor U14705 (N_14705,N_14578,N_14590);
nand U14706 (N_14706,N_14641,N_14594);
nor U14707 (N_14707,N_14628,N_14558);
nor U14708 (N_14708,N_14573,N_14636);
or U14709 (N_14709,N_14626,N_14580);
xor U14710 (N_14710,N_14649,N_14668);
or U14711 (N_14711,N_14585,N_14694);
or U14712 (N_14712,N_14620,N_14679);
xnor U14713 (N_14713,N_14607,N_14553);
nand U14714 (N_14714,N_14646,N_14695);
xnor U14715 (N_14715,N_14622,N_14629);
nand U14716 (N_14716,N_14645,N_14555);
or U14717 (N_14717,N_14644,N_14604);
xnor U14718 (N_14718,N_14608,N_14583);
nand U14719 (N_14719,N_14657,N_14688);
xnor U14720 (N_14720,N_14613,N_14687);
xor U14721 (N_14721,N_14564,N_14550);
or U14722 (N_14722,N_14568,N_14665);
or U14723 (N_14723,N_14581,N_14676);
or U14724 (N_14724,N_14632,N_14598);
nand U14725 (N_14725,N_14601,N_14683);
and U14726 (N_14726,N_14652,N_14663);
or U14727 (N_14727,N_14686,N_14662);
nor U14728 (N_14728,N_14648,N_14571);
xnor U14729 (N_14729,N_14691,N_14677);
nand U14730 (N_14730,N_14682,N_14659);
nand U14731 (N_14731,N_14557,N_14675);
nand U14732 (N_14732,N_14625,N_14637);
xnor U14733 (N_14733,N_14584,N_14559);
nor U14734 (N_14734,N_14654,N_14599);
xnor U14735 (N_14735,N_14595,N_14616);
and U14736 (N_14736,N_14653,N_14624);
or U14737 (N_14737,N_14664,N_14627);
or U14738 (N_14738,N_14619,N_14603);
nor U14739 (N_14739,N_14658,N_14651);
nor U14740 (N_14740,N_14689,N_14666);
xnor U14741 (N_14741,N_14639,N_14670);
nor U14742 (N_14742,N_14609,N_14575);
nor U14743 (N_14743,N_14596,N_14693);
and U14744 (N_14744,N_14656,N_14566);
nor U14745 (N_14745,N_14588,N_14605);
or U14746 (N_14746,N_14630,N_14692);
xor U14747 (N_14747,N_14660,N_14698);
or U14748 (N_14748,N_14699,N_14661);
nor U14749 (N_14749,N_14623,N_14638);
xnor U14750 (N_14750,N_14606,N_14671);
and U14751 (N_14751,N_14612,N_14574);
xnor U14752 (N_14752,N_14678,N_14615);
nand U14753 (N_14753,N_14587,N_14697);
nand U14754 (N_14754,N_14556,N_14610);
nand U14755 (N_14755,N_14690,N_14602);
nor U14756 (N_14756,N_14562,N_14635);
or U14757 (N_14757,N_14643,N_14572);
nor U14758 (N_14758,N_14617,N_14667);
nand U14759 (N_14759,N_14600,N_14577);
or U14760 (N_14760,N_14633,N_14591);
or U14761 (N_14761,N_14569,N_14631);
nand U14762 (N_14762,N_14684,N_14592);
nand U14763 (N_14763,N_14642,N_14696);
xnor U14764 (N_14764,N_14597,N_14593);
nand U14765 (N_14765,N_14570,N_14674);
nand U14766 (N_14766,N_14576,N_14685);
and U14767 (N_14767,N_14634,N_14586);
nand U14768 (N_14768,N_14621,N_14552);
and U14769 (N_14769,N_14579,N_14589);
and U14770 (N_14770,N_14614,N_14618);
xnor U14771 (N_14771,N_14647,N_14551);
or U14772 (N_14772,N_14673,N_14554);
xnor U14773 (N_14773,N_14567,N_14560);
and U14774 (N_14774,N_14565,N_14611);
and U14775 (N_14775,N_14569,N_14626);
or U14776 (N_14776,N_14687,N_14694);
nand U14777 (N_14777,N_14588,N_14557);
nand U14778 (N_14778,N_14655,N_14680);
xor U14779 (N_14779,N_14569,N_14661);
and U14780 (N_14780,N_14615,N_14590);
and U14781 (N_14781,N_14562,N_14614);
xnor U14782 (N_14782,N_14668,N_14570);
or U14783 (N_14783,N_14568,N_14598);
or U14784 (N_14784,N_14679,N_14644);
nand U14785 (N_14785,N_14593,N_14585);
or U14786 (N_14786,N_14608,N_14686);
nand U14787 (N_14787,N_14641,N_14671);
and U14788 (N_14788,N_14560,N_14605);
xnor U14789 (N_14789,N_14589,N_14663);
and U14790 (N_14790,N_14580,N_14617);
nor U14791 (N_14791,N_14595,N_14665);
and U14792 (N_14792,N_14661,N_14557);
or U14793 (N_14793,N_14696,N_14618);
or U14794 (N_14794,N_14683,N_14675);
or U14795 (N_14795,N_14568,N_14683);
xor U14796 (N_14796,N_14685,N_14607);
nor U14797 (N_14797,N_14631,N_14593);
xor U14798 (N_14798,N_14600,N_14685);
and U14799 (N_14799,N_14576,N_14552);
nand U14800 (N_14800,N_14640,N_14600);
and U14801 (N_14801,N_14582,N_14697);
xnor U14802 (N_14802,N_14565,N_14557);
and U14803 (N_14803,N_14587,N_14615);
and U14804 (N_14804,N_14604,N_14659);
and U14805 (N_14805,N_14603,N_14653);
nor U14806 (N_14806,N_14610,N_14607);
and U14807 (N_14807,N_14662,N_14691);
or U14808 (N_14808,N_14602,N_14629);
xnor U14809 (N_14809,N_14646,N_14626);
or U14810 (N_14810,N_14688,N_14690);
xor U14811 (N_14811,N_14650,N_14564);
or U14812 (N_14812,N_14566,N_14682);
or U14813 (N_14813,N_14637,N_14587);
nor U14814 (N_14814,N_14576,N_14657);
xor U14815 (N_14815,N_14595,N_14578);
xnor U14816 (N_14816,N_14583,N_14639);
nand U14817 (N_14817,N_14685,N_14589);
xnor U14818 (N_14818,N_14558,N_14647);
nor U14819 (N_14819,N_14629,N_14578);
or U14820 (N_14820,N_14691,N_14641);
nand U14821 (N_14821,N_14662,N_14591);
and U14822 (N_14822,N_14592,N_14639);
nand U14823 (N_14823,N_14688,N_14664);
nor U14824 (N_14824,N_14618,N_14684);
xor U14825 (N_14825,N_14686,N_14677);
nor U14826 (N_14826,N_14639,N_14644);
xnor U14827 (N_14827,N_14627,N_14679);
nor U14828 (N_14828,N_14591,N_14686);
or U14829 (N_14829,N_14662,N_14699);
nor U14830 (N_14830,N_14662,N_14567);
or U14831 (N_14831,N_14697,N_14687);
nor U14832 (N_14832,N_14604,N_14631);
nand U14833 (N_14833,N_14666,N_14639);
or U14834 (N_14834,N_14670,N_14559);
nand U14835 (N_14835,N_14556,N_14573);
xor U14836 (N_14836,N_14586,N_14624);
nand U14837 (N_14837,N_14568,N_14624);
xor U14838 (N_14838,N_14642,N_14560);
xnor U14839 (N_14839,N_14627,N_14590);
xor U14840 (N_14840,N_14673,N_14686);
nand U14841 (N_14841,N_14688,N_14672);
xnor U14842 (N_14842,N_14638,N_14695);
nor U14843 (N_14843,N_14578,N_14616);
and U14844 (N_14844,N_14688,N_14578);
and U14845 (N_14845,N_14590,N_14555);
xor U14846 (N_14846,N_14598,N_14668);
and U14847 (N_14847,N_14687,N_14625);
or U14848 (N_14848,N_14556,N_14560);
nand U14849 (N_14849,N_14554,N_14666);
xor U14850 (N_14850,N_14728,N_14701);
nor U14851 (N_14851,N_14785,N_14812);
and U14852 (N_14852,N_14800,N_14708);
nor U14853 (N_14853,N_14740,N_14741);
and U14854 (N_14854,N_14844,N_14791);
or U14855 (N_14855,N_14720,N_14709);
or U14856 (N_14856,N_14705,N_14807);
xor U14857 (N_14857,N_14768,N_14732);
and U14858 (N_14858,N_14826,N_14840);
and U14859 (N_14859,N_14811,N_14827);
and U14860 (N_14860,N_14841,N_14744);
nand U14861 (N_14861,N_14765,N_14838);
xor U14862 (N_14862,N_14763,N_14724);
and U14863 (N_14863,N_14719,N_14778);
or U14864 (N_14864,N_14794,N_14803);
and U14865 (N_14865,N_14750,N_14786);
and U14866 (N_14866,N_14714,N_14836);
nand U14867 (N_14867,N_14833,N_14815);
xor U14868 (N_14868,N_14804,N_14810);
or U14869 (N_14869,N_14760,N_14771);
nor U14870 (N_14870,N_14761,N_14755);
or U14871 (N_14871,N_14735,N_14801);
nor U14872 (N_14872,N_14706,N_14753);
and U14873 (N_14873,N_14776,N_14824);
or U14874 (N_14874,N_14817,N_14828);
or U14875 (N_14875,N_14843,N_14832);
nand U14876 (N_14876,N_14834,N_14730);
or U14877 (N_14877,N_14781,N_14792);
nand U14878 (N_14878,N_14777,N_14769);
nand U14879 (N_14879,N_14802,N_14700);
nor U14880 (N_14880,N_14752,N_14845);
and U14881 (N_14881,N_14770,N_14788);
nor U14882 (N_14882,N_14733,N_14842);
xor U14883 (N_14883,N_14715,N_14754);
or U14884 (N_14884,N_14703,N_14775);
and U14885 (N_14885,N_14835,N_14716);
nor U14886 (N_14886,N_14783,N_14746);
and U14887 (N_14887,N_14767,N_14848);
or U14888 (N_14888,N_14742,N_14723);
xor U14889 (N_14889,N_14774,N_14847);
nand U14890 (N_14890,N_14779,N_14766);
nor U14891 (N_14891,N_14789,N_14734);
nand U14892 (N_14892,N_14816,N_14738);
nand U14893 (N_14893,N_14757,N_14839);
nand U14894 (N_14894,N_14822,N_14756);
or U14895 (N_14895,N_14837,N_14731);
xnor U14896 (N_14896,N_14806,N_14846);
nor U14897 (N_14897,N_14711,N_14747);
xnor U14898 (N_14898,N_14796,N_14809);
xnor U14899 (N_14899,N_14821,N_14710);
or U14900 (N_14900,N_14790,N_14805);
nor U14901 (N_14901,N_14721,N_14818);
nor U14902 (N_14902,N_14729,N_14759);
or U14903 (N_14903,N_14758,N_14825);
xor U14904 (N_14904,N_14702,N_14749);
or U14905 (N_14905,N_14762,N_14726);
xor U14906 (N_14906,N_14739,N_14808);
xnor U14907 (N_14907,N_14798,N_14795);
and U14908 (N_14908,N_14722,N_14707);
xor U14909 (N_14909,N_14773,N_14819);
and U14910 (N_14910,N_14784,N_14748);
xnor U14911 (N_14911,N_14814,N_14787);
xor U14912 (N_14912,N_14737,N_14799);
or U14913 (N_14913,N_14718,N_14849);
or U14914 (N_14914,N_14725,N_14751);
or U14915 (N_14915,N_14813,N_14793);
or U14916 (N_14916,N_14727,N_14830);
and U14917 (N_14917,N_14717,N_14823);
or U14918 (N_14918,N_14820,N_14829);
nand U14919 (N_14919,N_14736,N_14782);
and U14920 (N_14920,N_14797,N_14743);
and U14921 (N_14921,N_14764,N_14713);
or U14922 (N_14922,N_14745,N_14780);
or U14923 (N_14923,N_14712,N_14772);
and U14924 (N_14924,N_14831,N_14704);
and U14925 (N_14925,N_14835,N_14843);
xnor U14926 (N_14926,N_14731,N_14734);
and U14927 (N_14927,N_14747,N_14732);
nand U14928 (N_14928,N_14735,N_14814);
or U14929 (N_14929,N_14732,N_14773);
or U14930 (N_14930,N_14819,N_14824);
or U14931 (N_14931,N_14798,N_14808);
nor U14932 (N_14932,N_14729,N_14745);
xnor U14933 (N_14933,N_14838,N_14704);
or U14934 (N_14934,N_14749,N_14802);
nor U14935 (N_14935,N_14715,N_14709);
xor U14936 (N_14936,N_14789,N_14834);
xor U14937 (N_14937,N_14832,N_14702);
and U14938 (N_14938,N_14841,N_14806);
and U14939 (N_14939,N_14706,N_14739);
or U14940 (N_14940,N_14833,N_14759);
nand U14941 (N_14941,N_14787,N_14723);
nor U14942 (N_14942,N_14735,N_14730);
or U14943 (N_14943,N_14741,N_14825);
and U14944 (N_14944,N_14754,N_14788);
nand U14945 (N_14945,N_14750,N_14806);
and U14946 (N_14946,N_14789,N_14784);
or U14947 (N_14947,N_14814,N_14756);
and U14948 (N_14948,N_14833,N_14775);
nor U14949 (N_14949,N_14736,N_14731);
or U14950 (N_14950,N_14743,N_14739);
nand U14951 (N_14951,N_14712,N_14724);
or U14952 (N_14952,N_14766,N_14773);
nand U14953 (N_14953,N_14838,N_14735);
or U14954 (N_14954,N_14779,N_14792);
nor U14955 (N_14955,N_14708,N_14733);
xor U14956 (N_14956,N_14817,N_14811);
nand U14957 (N_14957,N_14823,N_14832);
xnor U14958 (N_14958,N_14833,N_14755);
nor U14959 (N_14959,N_14700,N_14728);
nor U14960 (N_14960,N_14730,N_14746);
or U14961 (N_14961,N_14782,N_14759);
nor U14962 (N_14962,N_14817,N_14755);
nor U14963 (N_14963,N_14799,N_14782);
or U14964 (N_14964,N_14717,N_14810);
xnor U14965 (N_14965,N_14840,N_14707);
or U14966 (N_14966,N_14780,N_14770);
xnor U14967 (N_14967,N_14821,N_14826);
and U14968 (N_14968,N_14836,N_14769);
or U14969 (N_14969,N_14750,N_14797);
and U14970 (N_14970,N_14754,N_14702);
or U14971 (N_14971,N_14783,N_14777);
and U14972 (N_14972,N_14709,N_14744);
and U14973 (N_14973,N_14821,N_14832);
or U14974 (N_14974,N_14722,N_14761);
and U14975 (N_14975,N_14747,N_14824);
or U14976 (N_14976,N_14789,N_14709);
nand U14977 (N_14977,N_14790,N_14772);
and U14978 (N_14978,N_14707,N_14708);
nand U14979 (N_14979,N_14813,N_14786);
xor U14980 (N_14980,N_14715,N_14776);
and U14981 (N_14981,N_14831,N_14775);
and U14982 (N_14982,N_14844,N_14776);
nand U14983 (N_14983,N_14729,N_14711);
nand U14984 (N_14984,N_14740,N_14771);
nor U14985 (N_14985,N_14827,N_14831);
and U14986 (N_14986,N_14797,N_14727);
nand U14987 (N_14987,N_14750,N_14805);
xor U14988 (N_14988,N_14716,N_14808);
xor U14989 (N_14989,N_14777,N_14715);
or U14990 (N_14990,N_14788,N_14780);
xor U14991 (N_14991,N_14701,N_14748);
nand U14992 (N_14992,N_14756,N_14743);
nand U14993 (N_14993,N_14749,N_14711);
nand U14994 (N_14994,N_14773,N_14717);
or U14995 (N_14995,N_14713,N_14746);
xor U14996 (N_14996,N_14766,N_14754);
xnor U14997 (N_14997,N_14769,N_14738);
nor U14998 (N_14998,N_14708,N_14837);
and U14999 (N_14999,N_14725,N_14825);
nand UO_0 (O_0,N_14981,N_14956);
nor UO_1 (O_1,N_14906,N_14953);
xnor UO_2 (O_2,N_14904,N_14993);
xor UO_3 (O_3,N_14995,N_14855);
nand UO_4 (O_4,N_14909,N_14891);
and UO_5 (O_5,N_14896,N_14872);
nor UO_6 (O_6,N_14974,N_14985);
nand UO_7 (O_7,N_14980,N_14943);
or UO_8 (O_8,N_14913,N_14964);
nor UO_9 (O_9,N_14863,N_14895);
nand UO_10 (O_10,N_14900,N_14886);
nand UO_11 (O_11,N_14928,N_14888);
and UO_12 (O_12,N_14983,N_14989);
xnor UO_13 (O_13,N_14910,N_14991);
nor UO_14 (O_14,N_14887,N_14941);
nor UO_15 (O_15,N_14946,N_14967);
nand UO_16 (O_16,N_14873,N_14984);
nor UO_17 (O_17,N_14876,N_14977);
nor UO_18 (O_18,N_14965,N_14894);
xnor UO_19 (O_19,N_14911,N_14898);
nor UO_20 (O_20,N_14878,N_14933);
or UO_21 (O_21,N_14871,N_14973);
nand UO_22 (O_22,N_14999,N_14936);
nand UO_23 (O_23,N_14851,N_14955);
xnor UO_24 (O_24,N_14959,N_14882);
xor UO_25 (O_25,N_14963,N_14958);
nor UO_26 (O_26,N_14992,N_14901);
xor UO_27 (O_27,N_14951,N_14986);
nand UO_28 (O_28,N_14970,N_14982);
nor UO_29 (O_29,N_14978,N_14923);
and UO_30 (O_30,N_14877,N_14918);
nor UO_31 (O_31,N_14939,N_14949);
nand UO_32 (O_32,N_14926,N_14908);
and UO_33 (O_33,N_14868,N_14927);
xnor UO_34 (O_34,N_14937,N_14944);
nand UO_35 (O_35,N_14915,N_14945);
or UO_36 (O_36,N_14997,N_14902);
and UO_37 (O_37,N_14938,N_14935);
nor UO_38 (O_38,N_14920,N_14867);
nor UO_39 (O_39,N_14859,N_14899);
nand UO_40 (O_40,N_14931,N_14971);
or UO_41 (O_41,N_14914,N_14856);
or UO_42 (O_42,N_14921,N_14972);
nand UO_43 (O_43,N_14853,N_14930);
xnor UO_44 (O_44,N_14874,N_14885);
and UO_45 (O_45,N_14919,N_14892);
nand UO_46 (O_46,N_14932,N_14866);
or UO_47 (O_47,N_14881,N_14942);
or UO_48 (O_48,N_14934,N_14854);
xor UO_49 (O_49,N_14957,N_14869);
nand UO_50 (O_50,N_14952,N_14948);
xor UO_51 (O_51,N_14998,N_14917);
xnor UO_52 (O_52,N_14947,N_14875);
nand UO_53 (O_53,N_14925,N_14962);
and UO_54 (O_54,N_14966,N_14969);
nor UO_55 (O_55,N_14870,N_14990);
or UO_56 (O_56,N_14988,N_14864);
nor UO_57 (O_57,N_14865,N_14897);
xor UO_58 (O_58,N_14905,N_14976);
or UO_59 (O_59,N_14883,N_14994);
and UO_60 (O_60,N_14950,N_14862);
nand UO_61 (O_61,N_14979,N_14857);
xnor UO_62 (O_62,N_14929,N_14861);
xor UO_63 (O_63,N_14960,N_14987);
xnor UO_64 (O_64,N_14954,N_14907);
nand UO_65 (O_65,N_14912,N_14968);
nor UO_66 (O_66,N_14924,N_14975);
and UO_67 (O_67,N_14890,N_14922);
nand UO_68 (O_68,N_14860,N_14852);
nor UO_69 (O_69,N_14903,N_14889);
xnor UO_70 (O_70,N_14996,N_14880);
nor UO_71 (O_71,N_14893,N_14858);
nor UO_72 (O_72,N_14879,N_14940);
or UO_73 (O_73,N_14884,N_14916);
nor UO_74 (O_74,N_14961,N_14850);
and UO_75 (O_75,N_14930,N_14939);
xnor UO_76 (O_76,N_14971,N_14880);
nor UO_77 (O_77,N_14949,N_14953);
nor UO_78 (O_78,N_14949,N_14901);
xnor UO_79 (O_79,N_14942,N_14925);
nor UO_80 (O_80,N_14944,N_14931);
and UO_81 (O_81,N_14905,N_14980);
and UO_82 (O_82,N_14999,N_14983);
nor UO_83 (O_83,N_14902,N_14942);
nand UO_84 (O_84,N_14887,N_14936);
xor UO_85 (O_85,N_14868,N_14907);
or UO_86 (O_86,N_14924,N_14892);
xor UO_87 (O_87,N_14938,N_14901);
xor UO_88 (O_88,N_14943,N_14872);
nor UO_89 (O_89,N_14853,N_14896);
nand UO_90 (O_90,N_14929,N_14891);
and UO_91 (O_91,N_14863,N_14951);
nor UO_92 (O_92,N_14994,N_14967);
nand UO_93 (O_93,N_14930,N_14965);
or UO_94 (O_94,N_14999,N_14870);
nor UO_95 (O_95,N_14894,N_14970);
or UO_96 (O_96,N_14953,N_14918);
or UO_97 (O_97,N_14915,N_14971);
xnor UO_98 (O_98,N_14980,N_14960);
or UO_99 (O_99,N_14966,N_14920);
nor UO_100 (O_100,N_14920,N_14919);
or UO_101 (O_101,N_14873,N_14897);
nor UO_102 (O_102,N_14887,N_14913);
and UO_103 (O_103,N_14973,N_14979);
nor UO_104 (O_104,N_14880,N_14976);
xnor UO_105 (O_105,N_14874,N_14913);
and UO_106 (O_106,N_14925,N_14886);
nor UO_107 (O_107,N_14959,N_14977);
and UO_108 (O_108,N_14912,N_14870);
and UO_109 (O_109,N_14939,N_14923);
or UO_110 (O_110,N_14905,N_14934);
or UO_111 (O_111,N_14939,N_14943);
nand UO_112 (O_112,N_14918,N_14862);
nand UO_113 (O_113,N_14865,N_14884);
xor UO_114 (O_114,N_14881,N_14986);
nor UO_115 (O_115,N_14854,N_14974);
nand UO_116 (O_116,N_14969,N_14945);
nor UO_117 (O_117,N_14946,N_14930);
or UO_118 (O_118,N_14964,N_14867);
and UO_119 (O_119,N_14943,N_14990);
and UO_120 (O_120,N_14890,N_14929);
nor UO_121 (O_121,N_14853,N_14872);
and UO_122 (O_122,N_14927,N_14993);
nand UO_123 (O_123,N_14891,N_14855);
xnor UO_124 (O_124,N_14975,N_14946);
or UO_125 (O_125,N_14998,N_14953);
or UO_126 (O_126,N_14865,N_14879);
xor UO_127 (O_127,N_14986,N_14880);
or UO_128 (O_128,N_14885,N_14971);
nand UO_129 (O_129,N_14978,N_14862);
and UO_130 (O_130,N_14897,N_14867);
and UO_131 (O_131,N_14856,N_14931);
and UO_132 (O_132,N_14894,N_14891);
and UO_133 (O_133,N_14920,N_14971);
xor UO_134 (O_134,N_14910,N_14942);
nand UO_135 (O_135,N_14892,N_14968);
or UO_136 (O_136,N_14961,N_14872);
and UO_137 (O_137,N_14940,N_14948);
nor UO_138 (O_138,N_14904,N_14937);
and UO_139 (O_139,N_14850,N_14867);
nand UO_140 (O_140,N_14892,N_14870);
nor UO_141 (O_141,N_14991,N_14925);
or UO_142 (O_142,N_14942,N_14993);
xnor UO_143 (O_143,N_14951,N_14869);
xor UO_144 (O_144,N_14917,N_14978);
nor UO_145 (O_145,N_14963,N_14860);
and UO_146 (O_146,N_14887,N_14883);
or UO_147 (O_147,N_14908,N_14938);
xor UO_148 (O_148,N_14998,N_14938);
nand UO_149 (O_149,N_14894,N_14916);
or UO_150 (O_150,N_14945,N_14861);
or UO_151 (O_151,N_14966,N_14949);
nand UO_152 (O_152,N_14935,N_14976);
and UO_153 (O_153,N_14892,N_14923);
or UO_154 (O_154,N_14915,N_14909);
xnor UO_155 (O_155,N_14893,N_14983);
and UO_156 (O_156,N_14892,N_14859);
nand UO_157 (O_157,N_14996,N_14976);
and UO_158 (O_158,N_14934,N_14864);
or UO_159 (O_159,N_14948,N_14919);
nand UO_160 (O_160,N_14871,N_14923);
xnor UO_161 (O_161,N_14979,N_14964);
nand UO_162 (O_162,N_14933,N_14870);
xnor UO_163 (O_163,N_14988,N_14986);
nor UO_164 (O_164,N_14964,N_14880);
nand UO_165 (O_165,N_14951,N_14874);
xor UO_166 (O_166,N_14855,N_14955);
nor UO_167 (O_167,N_14934,N_14965);
xnor UO_168 (O_168,N_14952,N_14957);
nor UO_169 (O_169,N_14942,N_14933);
and UO_170 (O_170,N_14964,N_14948);
or UO_171 (O_171,N_14959,N_14893);
and UO_172 (O_172,N_14858,N_14875);
xnor UO_173 (O_173,N_14881,N_14935);
nor UO_174 (O_174,N_14895,N_14905);
or UO_175 (O_175,N_14951,N_14871);
xor UO_176 (O_176,N_14866,N_14968);
xnor UO_177 (O_177,N_14910,N_14890);
or UO_178 (O_178,N_14978,N_14891);
or UO_179 (O_179,N_14926,N_14891);
and UO_180 (O_180,N_14999,N_14858);
xor UO_181 (O_181,N_14984,N_14982);
nand UO_182 (O_182,N_14946,N_14994);
and UO_183 (O_183,N_14950,N_14937);
nor UO_184 (O_184,N_14970,N_14866);
xor UO_185 (O_185,N_14914,N_14905);
and UO_186 (O_186,N_14997,N_14915);
or UO_187 (O_187,N_14856,N_14881);
or UO_188 (O_188,N_14905,N_14998);
xnor UO_189 (O_189,N_14905,N_14944);
or UO_190 (O_190,N_14861,N_14908);
nand UO_191 (O_191,N_14943,N_14944);
or UO_192 (O_192,N_14980,N_14999);
xnor UO_193 (O_193,N_14898,N_14979);
nand UO_194 (O_194,N_14888,N_14944);
nor UO_195 (O_195,N_14940,N_14964);
xnor UO_196 (O_196,N_14913,N_14893);
nand UO_197 (O_197,N_14888,N_14934);
xnor UO_198 (O_198,N_14924,N_14997);
or UO_199 (O_199,N_14962,N_14967);
and UO_200 (O_200,N_14921,N_14854);
nor UO_201 (O_201,N_14905,N_14873);
or UO_202 (O_202,N_14869,N_14859);
or UO_203 (O_203,N_14855,N_14864);
xor UO_204 (O_204,N_14892,N_14914);
and UO_205 (O_205,N_14912,N_14899);
or UO_206 (O_206,N_14923,N_14925);
xnor UO_207 (O_207,N_14952,N_14873);
or UO_208 (O_208,N_14975,N_14936);
xor UO_209 (O_209,N_14953,N_14880);
xor UO_210 (O_210,N_14945,N_14982);
or UO_211 (O_211,N_14952,N_14977);
xnor UO_212 (O_212,N_14879,N_14956);
or UO_213 (O_213,N_14874,N_14995);
and UO_214 (O_214,N_14991,N_14850);
nand UO_215 (O_215,N_14938,N_14867);
xnor UO_216 (O_216,N_14972,N_14962);
xor UO_217 (O_217,N_14934,N_14946);
nand UO_218 (O_218,N_14925,N_14943);
and UO_219 (O_219,N_14984,N_14970);
xnor UO_220 (O_220,N_14944,N_14913);
or UO_221 (O_221,N_14992,N_14925);
nor UO_222 (O_222,N_14946,N_14947);
or UO_223 (O_223,N_14889,N_14854);
xor UO_224 (O_224,N_14919,N_14995);
xor UO_225 (O_225,N_14908,N_14901);
xor UO_226 (O_226,N_14918,N_14996);
xnor UO_227 (O_227,N_14881,N_14965);
or UO_228 (O_228,N_14862,N_14881);
and UO_229 (O_229,N_14947,N_14914);
or UO_230 (O_230,N_14999,N_14923);
xor UO_231 (O_231,N_14925,N_14931);
or UO_232 (O_232,N_14981,N_14928);
or UO_233 (O_233,N_14969,N_14974);
and UO_234 (O_234,N_14866,N_14938);
or UO_235 (O_235,N_14970,N_14858);
or UO_236 (O_236,N_14986,N_14897);
xor UO_237 (O_237,N_14880,N_14892);
and UO_238 (O_238,N_14879,N_14962);
or UO_239 (O_239,N_14943,N_14884);
and UO_240 (O_240,N_14908,N_14882);
xnor UO_241 (O_241,N_14881,N_14912);
xnor UO_242 (O_242,N_14972,N_14887);
nor UO_243 (O_243,N_14897,N_14898);
nand UO_244 (O_244,N_14903,N_14928);
nand UO_245 (O_245,N_14938,N_14937);
and UO_246 (O_246,N_14932,N_14980);
nand UO_247 (O_247,N_14951,N_14953);
nand UO_248 (O_248,N_14861,N_14997);
xnor UO_249 (O_249,N_14891,N_14948);
and UO_250 (O_250,N_14965,N_14916);
and UO_251 (O_251,N_14948,N_14975);
xor UO_252 (O_252,N_14855,N_14944);
nand UO_253 (O_253,N_14860,N_14911);
or UO_254 (O_254,N_14850,N_14871);
and UO_255 (O_255,N_14882,N_14881);
xnor UO_256 (O_256,N_14987,N_14978);
nor UO_257 (O_257,N_14903,N_14975);
nor UO_258 (O_258,N_14905,N_14978);
and UO_259 (O_259,N_14955,N_14966);
xnor UO_260 (O_260,N_14930,N_14947);
or UO_261 (O_261,N_14854,N_14868);
or UO_262 (O_262,N_14930,N_14978);
xnor UO_263 (O_263,N_14976,N_14888);
nor UO_264 (O_264,N_14909,N_14959);
nand UO_265 (O_265,N_14991,N_14964);
nand UO_266 (O_266,N_14915,N_14949);
or UO_267 (O_267,N_14908,N_14985);
xnor UO_268 (O_268,N_14950,N_14984);
xnor UO_269 (O_269,N_14990,N_14973);
and UO_270 (O_270,N_14933,N_14911);
xor UO_271 (O_271,N_14888,N_14963);
xnor UO_272 (O_272,N_14905,N_14927);
xnor UO_273 (O_273,N_14879,N_14985);
xor UO_274 (O_274,N_14866,N_14967);
or UO_275 (O_275,N_14870,N_14998);
nand UO_276 (O_276,N_14881,N_14873);
xor UO_277 (O_277,N_14852,N_14881);
nand UO_278 (O_278,N_14920,N_14855);
and UO_279 (O_279,N_14940,N_14884);
nand UO_280 (O_280,N_14881,N_14911);
nand UO_281 (O_281,N_14896,N_14883);
and UO_282 (O_282,N_14877,N_14939);
or UO_283 (O_283,N_14863,N_14866);
and UO_284 (O_284,N_14955,N_14869);
nor UO_285 (O_285,N_14922,N_14913);
nor UO_286 (O_286,N_14940,N_14927);
xor UO_287 (O_287,N_14896,N_14869);
nand UO_288 (O_288,N_14931,N_14929);
xor UO_289 (O_289,N_14886,N_14860);
or UO_290 (O_290,N_14965,N_14952);
or UO_291 (O_291,N_14991,N_14935);
or UO_292 (O_292,N_14990,N_14897);
xor UO_293 (O_293,N_14897,N_14936);
xor UO_294 (O_294,N_14903,N_14979);
nor UO_295 (O_295,N_14999,N_14907);
xor UO_296 (O_296,N_14891,N_14872);
and UO_297 (O_297,N_14991,N_14941);
and UO_298 (O_298,N_14900,N_14891);
xnor UO_299 (O_299,N_14908,N_14951);
and UO_300 (O_300,N_14991,N_14921);
and UO_301 (O_301,N_14906,N_14995);
nand UO_302 (O_302,N_14915,N_14883);
xor UO_303 (O_303,N_14878,N_14996);
and UO_304 (O_304,N_14965,N_14863);
xnor UO_305 (O_305,N_14881,N_14998);
nand UO_306 (O_306,N_14964,N_14956);
nand UO_307 (O_307,N_14868,N_14981);
or UO_308 (O_308,N_14907,N_14956);
nand UO_309 (O_309,N_14867,N_14979);
and UO_310 (O_310,N_14952,N_14931);
nand UO_311 (O_311,N_14929,N_14928);
and UO_312 (O_312,N_14902,N_14896);
or UO_313 (O_313,N_14883,N_14969);
nand UO_314 (O_314,N_14870,N_14994);
nand UO_315 (O_315,N_14946,N_14884);
nand UO_316 (O_316,N_14983,N_14981);
or UO_317 (O_317,N_14976,N_14850);
xor UO_318 (O_318,N_14983,N_14954);
or UO_319 (O_319,N_14876,N_14966);
nand UO_320 (O_320,N_14989,N_14875);
and UO_321 (O_321,N_14922,N_14888);
nand UO_322 (O_322,N_14850,N_14893);
or UO_323 (O_323,N_14857,N_14865);
or UO_324 (O_324,N_14976,N_14925);
or UO_325 (O_325,N_14869,N_14853);
and UO_326 (O_326,N_14962,N_14853);
xor UO_327 (O_327,N_14956,N_14916);
nor UO_328 (O_328,N_14913,N_14951);
nor UO_329 (O_329,N_14933,N_14853);
or UO_330 (O_330,N_14950,N_14944);
or UO_331 (O_331,N_14912,N_14867);
nand UO_332 (O_332,N_14986,N_14878);
xor UO_333 (O_333,N_14930,N_14903);
and UO_334 (O_334,N_14900,N_14866);
or UO_335 (O_335,N_14927,N_14982);
nor UO_336 (O_336,N_14876,N_14983);
and UO_337 (O_337,N_14861,N_14937);
or UO_338 (O_338,N_14985,N_14929);
xor UO_339 (O_339,N_14918,N_14903);
xnor UO_340 (O_340,N_14861,N_14886);
or UO_341 (O_341,N_14854,N_14850);
nand UO_342 (O_342,N_14851,N_14882);
and UO_343 (O_343,N_14883,N_14859);
and UO_344 (O_344,N_14911,N_14861);
nor UO_345 (O_345,N_14940,N_14905);
nand UO_346 (O_346,N_14854,N_14853);
and UO_347 (O_347,N_14973,N_14860);
nand UO_348 (O_348,N_14966,N_14918);
nand UO_349 (O_349,N_14932,N_14991);
and UO_350 (O_350,N_14962,N_14856);
or UO_351 (O_351,N_14976,N_14928);
nand UO_352 (O_352,N_14868,N_14890);
nor UO_353 (O_353,N_14910,N_14896);
and UO_354 (O_354,N_14949,N_14881);
or UO_355 (O_355,N_14950,N_14939);
nor UO_356 (O_356,N_14957,N_14962);
or UO_357 (O_357,N_14891,N_14994);
xor UO_358 (O_358,N_14905,N_14942);
or UO_359 (O_359,N_14865,N_14921);
nand UO_360 (O_360,N_14995,N_14854);
xor UO_361 (O_361,N_14912,N_14935);
nand UO_362 (O_362,N_14896,N_14867);
nor UO_363 (O_363,N_14874,N_14965);
nand UO_364 (O_364,N_14893,N_14949);
xor UO_365 (O_365,N_14959,N_14944);
xnor UO_366 (O_366,N_14939,N_14996);
nand UO_367 (O_367,N_14933,N_14998);
xor UO_368 (O_368,N_14917,N_14879);
nor UO_369 (O_369,N_14851,N_14934);
xor UO_370 (O_370,N_14935,N_14939);
xor UO_371 (O_371,N_14897,N_14900);
xnor UO_372 (O_372,N_14914,N_14929);
xnor UO_373 (O_373,N_14907,N_14920);
xor UO_374 (O_374,N_14993,N_14950);
xnor UO_375 (O_375,N_14878,N_14924);
and UO_376 (O_376,N_14952,N_14930);
nor UO_377 (O_377,N_14870,N_14995);
xnor UO_378 (O_378,N_14999,N_14996);
xor UO_379 (O_379,N_14882,N_14978);
nand UO_380 (O_380,N_14856,N_14972);
xor UO_381 (O_381,N_14855,N_14940);
xor UO_382 (O_382,N_14962,N_14951);
nor UO_383 (O_383,N_14988,N_14914);
xnor UO_384 (O_384,N_14892,N_14918);
xor UO_385 (O_385,N_14857,N_14905);
nor UO_386 (O_386,N_14884,N_14911);
nand UO_387 (O_387,N_14886,N_14973);
or UO_388 (O_388,N_14859,N_14851);
xor UO_389 (O_389,N_14892,N_14860);
or UO_390 (O_390,N_14971,N_14863);
xor UO_391 (O_391,N_14970,N_14886);
nor UO_392 (O_392,N_14936,N_14978);
and UO_393 (O_393,N_14975,N_14853);
or UO_394 (O_394,N_14931,N_14887);
and UO_395 (O_395,N_14982,N_14971);
nor UO_396 (O_396,N_14923,N_14994);
xnor UO_397 (O_397,N_14926,N_14943);
and UO_398 (O_398,N_14912,N_14958);
nand UO_399 (O_399,N_14868,N_14979);
or UO_400 (O_400,N_14916,N_14872);
and UO_401 (O_401,N_14941,N_14910);
nand UO_402 (O_402,N_14983,N_14913);
nor UO_403 (O_403,N_14874,N_14941);
xor UO_404 (O_404,N_14852,N_14886);
and UO_405 (O_405,N_14988,N_14862);
nand UO_406 (O_406,N_14856,N_14951);
xor UO_407 (O_407,N_14921,N_14968);
xnor UO_408 (O_408,N_14892,N_14887);
or UO_409 (O_409,N_14985,N_14887);
nor UO_410 (O_410,N_14855,N_14907);
xnor UO_411 (O_411,N_14880,N_14859);
and UO_412 (O_412,N_14863,N_14993);
or UO_413 (O_413,N_14862,N_14951);
nand UO_414 (O_414,N_14914,N_14878);
and UO_415 (O_415,N_14902,N_14970);
xnor UO_416 (O_416,N_14910,N_14857);
nor UO_417 (O_417,N_14851,N_14855);
nor UO_418 (O_418,N_14968,N_14944);
xnor UO_419 (O_419,N_14950,N_14852);
nor UO_420 (O_420,N_14853,N_14858);
and UO_421 (O_421,N_14907,N_14857);
xor UO_422 (O_422,N_14986,N_14987);
and UO_423 (O_423,N_14934,N_14900);
nand UO_424 (O_424,N_14977,N_14945);
nand UO_425 (O_425,N_14968,N_14956);
or UO_426 (O_426,N_14870,N_14900);
nor UO_427 (O_427,N_14877,N_14953);
or UO_428 (O_428,N_14921,N_14943);
and UO_429 (O_429,N_14918,N_14938);
xor UO_430 (O_430,N_14893,N_14904);
nor UO_431 (O_431,N_14866,N_14982);
xor UO_432 (O_432,N_14990,N_14966);
or UO_433 (O_433,N_14861,N_14895);
or UO_434 (O_434,N_14980,N_14914);
nand UO_435 (O_435,N_14931,N_14923);
and UO_436 (O_436,N_14977,N_14869);
nand UO_437 (O_437,N_14977,N_14918);
nor UO_438 (O_438,N_14949,N_14913);
nand UO_439 (O_439,N_14917,N_14983);
nor UO_440 (O_440,N_14936,N_14994);
and UO_441 (O_441,N_14897,N_14917);
nor UO_442 (O_442,N_14953,N_14868);
nand UO_443 (O_443,N_14966,N_14961);
xor UO_444 (O_444,N_14943,N_14935);
and UO_445 (O_445,N_14969,N_14891);
nor UO_446 (O_446,N_14948,N_14978);
nor UO_447 (O_447,N_14938,N_14974);
xnor UO_448 (O_448,N_14903,N_14885);
nor UO_449 (O_449,N_14904,N_14899);
nand UO_450 (O_450,N_14934,N_14876);
and UO_451 (O_451,N_14887,N_14899);
or UO_452 (O_452,N_14940,N_14986);
nand UO_453 (O_453,N_14911,N_14853);
or UO_454 (O_454,N_14904,N_14883);
xnor UO_455 (O_455,N_14916,N_14979);
xnor UO_456 (O_456,N_14897,N_14925);
xor UO_457 (O_457,N_14850,N_14998);
nor UO_458 (O_458,N_14922,N_14875);
and UO_459 (O_459,N_14920,N_14859);
xnor UO_460 (O_460,N_14981,N_14991);
nor UO_461 (O_461,N_14876,N_14879);
xnor UO_462 (O_462,N_14947,N_14971);
nand UO_463 (O_463,N_14964,N_14903);
and UO_464 (O_464,N_14898,N_14963);
xnor UO_465 (O_465,N_14933,N_14939);
and UO_466 (O_466,N_14880,N_14918);
or UO_467 (O_467,N_14931,N_14985);
xor UO_468 (O_468,N_14966,N_14989);
nand UO_469 (O_469,N_14867,N_14936);
or UO_470 (O_470,N_14918,N_14949);
nor UO_471 (O_471,N_14892,N_14927);
and UO_472 (O_472,N_14946,N_14865);
nand UO_473 (O_473,N_14877,N_14962);
or UO_474 (O_474,N_14896,N_14984);
or UO_475 (O_475,N_14964,N_14995);
nor UO_476 (O_476,N_14883,N_14942);
nor UO_477 (O_477,N_14957,N_14890);
nor UO_478 (O_478,N_14999,N_14944);
and UO_479 (O_479,N_14908,N_14990);
or UO_480 (O_480,N_14890,N_14901);
nand UO_481 (O_481,N_14948,N_14994);
and UO_482 (O_482,N_14936,N_14890);
and UO_483 (O_483,N_14852,N_14974);
nand UO_484 (O_484,N_14941,N_14919);
nand UO_485 (O_485,N_14952,N_14990);
nor UO_486 (O_486,N_14913,N_14939);
and UO_487 (O_487,N_14946,N_14892);
or UO_488 (O_488,N_14885,N_14924);
and UO_489 (O_489,N_14979,N_14974);
and UO_490 (O_490,N_14964,N_14932);
nor UO_491 (O_491,N_14905,N_14872);
xnor UO_492 (O_492,N_14975,N_14885);
or UO_493 (O_493,N_14881,N_14853);
xor UO_494 (O_494,N_14862,N_14860);
nand UO_495 (O_495,N_14894,N_14919);
and UO_496 (O_496,N_14903,N_14944);
and UO_497 (O_497,N_14935,N_14862);
nand UO_498 (O_498,N_14990,N_14957);
nor UO_499 (O_499,N_14925,N_14918);
nand UO_500 (O_500,N_14941,N_14917);
xor UO_501 (O_501,N_14964,N_14934);
nand UO_502 (O_502,N_14906,N_14904);
and UO_503 (O_503,N_14854,N_14942);
nor UO_504 (O_504,N_14970,N_14937);
or UO_505 (O_505,N_14955,N_14975);
nand UO_506 (O_506,N_14960,N_14958);
nor UO_507 (O_507,N_14982,N_14948);
nor UO_508 (O_508,N_14914,N_14864);
and UO_509 (O_509,N_14949,N_14974);
or UO_510 (O_510,N_14888,N_14997);
nor UO_511 (O_511,N_14930,N_14956);
and UO_512 (O_512,N_14939,N_14870);
or UO_513 (O_513,N_14865,N_14896);
or UO_514 (O_514,N_14865,N_14996);
xnor UO_515 (O_515,N_14933,N_14915);
and UO_516 (O_516,N_14931,N_14893);
nand UO_517 (O_517,N_14913,N_14989);
or UO_518 (O_518,N_14953,N_14939);
nor UO_519 (O_519,N_14877,N_14927);
and UO_520 (O_520,N_14977,N_14897);
and UO_521 (O_521,N_14898,N_14985);
xnor UO_522 (O_522,N_14954,N_14877);
nor UO_523 (O_523,N_14880,N_14867);
and UO_524 (O_524,N_14974,N_14986);
nor UO_525 (O_525,N_14963,N_14961);
or UO_526 (O_526,N_14850,N_14981);
xnor UO_527 (O_527,N_14916,N_14912);
nand UO_528 (O_528,N_14984,N_14859);
and UO_529 (O_529,N_14865,N_14872);
and UO_530 (O_530,N_14969,N_14940);
xnor UO_531 (O_531,N_14954,N_14895);
nand UO_532 (O_532,N_14977,N_14981);
nand UO_533 (O_533,N_14942,N_14893);
or UO_534 (O_534,N_14925,N_14853);
or UO_535 (O_535,N_14945,N_14904);
nor UO_536 (O_536,N_14939,N_14951);
and UO_537 (O_537,N_14964,N_14917);
nor UO_538 (O_538,N_14900,N_14896);
or UO_539 (O_539,N_14943,N_14918);
xor UO_540 (O_540,N_14876,N_14936);
or UO_541 (O_541,N_14977,N_14887);
or UO_542 (O_542,N_14934,N_14980);
or UO_543 (O_543,N_14944,N_14936);
and UO_544 (O_544,N_14915,N_14924);
xnor UO_545 (O_545,N_14966,N_14924);
nand UO_546 (O_546,N_14850,N_14988);
or UO_547 (O_547,N_14886,N_14978);
nor UO_548 (O_548,N_14980,N_14986);
nand UO_549 (O_549,N_14989,N_14948);
nand UO_550 (O_550,N_14983,N_14934);
nand UO_551 (O_551,N_14979,N_14854);
nor UO_552 (O_552,N_14931,N_14896);
xor UO_553 (O_553,N_14857,N_14994);
nor UO_554 (O_554,N_14977,N_14854);
nand UO_555 (O_555,N_14898,N_14909);
or UO_556 (O_556,N_14953,N_14969);
or UO_557 (O_557,N_14965,N_14933);
and UO_558 (O_558,N_14904,N_14947);
nand UO_559 (O_559,N_14964,N_14910);
nor UO_560 (O_560,N_14906,N_14980);
and UO_561 (O_561,N_14851,N_14856);
or UO_562 (O_562,N_14934,N_14925);
and UO_563 (O_563,N_14915,N_14864);
nand UO_564 (O_564,N_14906,N_14946);
or UO_565 (O_565,N_14900,N_14964);
nor UO_566 (O_566,N_14876,N_14923);
nand UO_567 (O_567,N_14990,N_14989);
or UO_568 (O_568,N_14864,N_14876);
nand UO_569 (O_569,N_14946,N_14921);
or UO_570 (O_570,N_14954,N_14977);
and UO_571 (O_571,N_14851,N_14901);
nand UO_572 (O_572,N_14944,N_14907);
nor UO_573 (O_573,N_14982,N_14884);
xnor UO_574 (O_574,N_14915,N_14887);
nor UO_575 (O_575,N_14967,N_14971);
and UO_576 (O_576,N_14920,N_14961);
nand UO_577 (O_577,N_14866,N_14875);
nand UO_578 (O_578,N_14905,N_14887);
nor UO_579 (O_579,N_14859,N_14956);
or UO_580 (O_580,N_14911,N_14970);
and UO_581 (O_581,N_14975,N_14867);
or UO_582 (O_582,N_14966,N_14890);
and UO_583 (O_583,N_14912,N_14986);
nand UO_584 (O_584,N_14901,N_14860);
nor UO_585 (O_585,N_14985,N_14987);
xor UO_586 (O_586,N_14882,N_14929);
xnor UO_587 (O_587,N_14892,N_14988);
nand UO_588 (O_588,N_14962,N_14871);
or UO_589 (O_589,N_14931,N_14872);
or UO_590 (O_590,N_14863,N_14902);
nor UO_591 (O_591,N_14906,N_14882);
xor UO_592 (O_592,N_14927,N_14878);
and UO_593 (O_593,N_14932,N_14996);
xor UO_594 (O_594,N_14926,N_14860);
and UO_595 (O_595,N_14907,N_14962);
xnor UO_596 (O_596,N_14985,N_14882);
nor UO_597 (O_597,N_14980,N_14865);
xor UO_598 (O_598,N_14964,N_14955);
nor UO_599 (O_599,N_14991,N_14904);
nand UO_600 (O_600,N_14959,N_14870);
xnor UO_601 (O_601,N_14938,N_14885);
nand UO_602 (O_602,N_14979,N_14913);
and UO_603 (O_603,N_14953,N_14862);
xnor UO_604 (O_604,N_14878,N_14889);
xnor UO_605 (O_605,N_14876,N_14892);
or UO_606 (O_606,N_14869,N_14959);
or UO_607 (O_607,N_14855,N_14931);
and UO_608 (O_608,N_14852,N_14961);
nor UO_609 (O_609,N_14942,N_14874);
and UO_610 (O_610,N_14884,N_14878);
xor UO_611 (O_611,N_14963,N_14869);
and UO_612 (O_612,N_14954,N_14924);
nor UO_613 (O_613,N_14871,N_14852);
and UO_614 (O_614,N_14923,N_14921);
and UO_615 (O_615,N_14935,N_14953);
nor UO_616 (O_616,N_14997,N_14876);
and UO_617 (O_617,N_14921,N_14851);
or UO_618 (O_618,N_14928,N_14853);
xnor UO_619 (O_619,N_14919,N_14896);
nand UO_620 (O_620,N_14856,N_14869);
or UO_621 (O_621,N_14904,N_14921);
and UO_622 (O_622,N_14902,N_14906);
nand UO_623 (O_623,N_14968,N_14941);
nor UO_624 (O_624,N_14987,N_14865);
nand UO_625 (O_625,N_14943,N_14955);
and UO_626 (O_626,N_14965,N_14938);
nor UO_627 (O_627,N_14946,N_14873);
nand UO_628 (O_628,N_14903,N_14994);
or UO_629 (O_629,N_14988,N_14904);
nor UO_630 (O_630,N_14998,N_14893);
nand UO_631 (O_631,N_14993,N_14924);
nand UO_632 (O_632,N_14860,N_14918);
or UO_633 (O_633,N_14914,N_14854);
or UO_634 (O_634,N_14958,N_14860);
xnor UO_635 (O_635,N_14941,N_14883);
nand UO_636 (O_636,N_14877,N_14982);
or UO_637 (O_637,N_14869,N_14904);
nand UO_638 (O_638,N_14951,N_14890);
and UO_639 (O_639,N_14964,N_14883);
and UO_640 (O_640,N_14987,N_14903);
or UO_641 (O_641,N_14895,N_14858);
nand UO_642 (O_642,N_14894,N_14937);
nand UO_643 (O_643,N_14925,N_14965);
xnor UO_644 (O_644,N_14930,N_14858);
nand UO_645 (O_645,N_14918,N_14850);
nand UO_646 (O_646,N_14964,N_14989);
nand UO_647 (O_647,N_14867,N_14909);
nand UO_648 (O_648,N_14859,N_14967);
nor UO_649 (O_649,N_14965,N_14905);
or UO_650 (O_650,N_14997,N_14857);
or UO_651 (O_651,N_14945,N_14981);
or UO_652 (O_652,N_14922,N_14932);
or UO_653 (O_653,N_14913,N_14864);
xnor UO_654 (O_654,N_14863,N_14959);
and UO_655 (O_655,N_14869,N_14958);
nand UO_656 (O_656,N_14966,N_14975);
or UO_657 (O_657,N_14941,N_14988);
nand UO_658 (O_658,N_14907,N_14890);
nand UO_659 (O_659,N_14919,N_14886);
xnor UO_660 (O_660,N_14951,N_14943);
nor UO_661 (O_661,N_14948,N_14869);
or UO_662 (O_662,N_14869,N_14871);
and UO_663 (O_663,N_14906,N_14955);
nor UO_664 (O_664,N_14941,N_14895);
and UO_665 (O_665,N_14853,N_14892);
or UO_666 (O_666,N_14959,N_14967);
or UO_667 (O_667,N_14998,N_14992);
nand UO_668 (O_668,N_14908,N_14899);
and UO_669 (O_669,N_14875,N_14973);
and UO_670 (O_670,N_14916,N_14907);
xor UO_671 (O_671,N_14965,N_14942);
nor UO_672 (O_672,N_14989,N_14953);
or UO_673 (O_673,N_14883,N_14977);
nor UO_674 (O_674,N_14994,N_14998);
xor UO_675 (O_675,N_14942,N_14894);
or UO_676 (O_676,N_14941,N_14906);
xor UO_677 (O_677,N_14890,N_14896);
or UO_678 (O_678,N_14913,N_14918);
xnor UO_679 (O_679,N_14951,N_14979);
nor UO_680 (O_680,N_14977,N_14940);
xor UO_681 (O_681,N_14935,N_14980);
or UO_682 (O_682,N_14871,N_14937);
nor UO_683 (O_683,N_14978,N_14944);
nand UO_684 (O_684,N_14979,N_14896);
nand UO_685 (O_685,N_14994,N_14897);
nor UO_686 (O_686,N_14979,N_14990);
nand UO_687 (O_687,N_14873,N_14864);
nand UO_688 (O_688,N_14960,N_14866);
or UO_689 (O_689,N_14980,N_14950);
and UO_690 (O_690,N_14861,N_14956);
xnor UO_691 (O_691,N_14906,N_14852);
and UO_692 (O_692,N_14985,N_14855);
nor UO_693 (O_693,N_14934,N_14986);
nand UO_694 (O_694,N_14930,N_14856);
or UO_695 (O_695,N_14964,N_14862);
nand UO_696 (O_696,N_14886,N_14894);
xnor UO_697 (O_697,N_14993,N_14979);
or UO_698 (O_698,N_14944,N_14857);
nor UO_699 (O_699,N_14903,N_14867);
nand UO_700 (O_700,N_14879,N_14974);
or UO_701 (O_701,N_14985,N_14948);
and UO_702 (O_702,N_14959,N_14924);
xor UO_703 (O_703,N_14951,N_14868);
xnor UO_704 (O_704,N_14959,N_14994);
nor UO_705 (O_705,N_14900,N_14942);
or UO_706 (O_706,N_14974,N_14981);
and UO_707 (O_707,N_14893,N_14908);
nor UO_708 (O_708,N_14917,N_14863);
nor UO_709 (O_709,N_14985,N_14873);
or UO_710 (O_710,N_14865,N_14894);
nand UO_711 (O_711,N_14867,N_14866);
or UO_712 (O_712,N_14969,N_14952);
nand UO_713 (O_713,N_14895,N_14862);
and UO_714 (O_714,N_14856,N_14996);
and UO_715 (O_715,N_14983,N_14973);
nand UO_716 (O_716,N_14986,N_14926);
nand UO_717 (O_717,N_14870,N_14871);
or UO_718 (O_718,N_14892,N_14897);
xor UO_719 (O_719,N_14945,N_14899);
xnor UO_720 (O_720,N_14909,N_14934);
xnor UO_721 (O_721,N_14994,N_14875);
nand UO_722 (O_722,N_14853,N_14886);
or UO_723 (O_723,N_14936,N_14862);
nor UO_724 (O_724,N_14915,N_14852);
and UO_725 (O_725,N_14994,N_14949);
nor UO_726 (O_726,N_14931,N_14895);
and UO_727 (O_727,N_14850,N_14884);
and UO_728 (O_728,N_14889,N_14897);
and UO_729 (O_729,N_14973,N_14939);
and UO_730 (O_730,N_14911,N_14997);
nor UO_731 (O_731,N_14872,N_14877);
xor UO_732 (O_732,N_14957,N_14868);
or UO_733 (O_733,N_14948,N_14918);
and UO_734 (O_734,N_14914,N_14851);
nor UO_735 (O_735,N_14858,N_14975);
and UO_736 (O_736,N_14995,N_14979);
and UO_737 (O_737,N_14936,N_14959);
and UO_738 (O_738,N_14956,N_14986);
xor UO_739 (O_739,N_14933,N_14904);
nor UO_740 (O_740,N_14886,N_14864);
or UO_741 (O_741,N_14971,N_14861);
nand UO_742 (O_742,N_14992,N_14979);
and UO_743 (O_743,N_14895,N_14909);
and UO_744 (O_744,N_14934,N_14917);
or UO_745 (O_745,N_14900,N_14912);
nor UO_746 (O_746,N_14902,N_14850);
and UO_747 (O_747,N_14893,N_14946);
or UO_748 (O_748,N_14889,N_14918);
and UO_749 (O_749,N_14966,N_14985);
nand UO_750 (O_750,N_14957,N_14949);
nor UO_751 (O_751,N_14951,N_14987);
or UO_752 (O_752,N_14984,N_14976);
xnor UO_753 (O_753,N_14928,N_14918);
or UO_754 (O_754,N_14981,N_14926);
and UO_755 (O_755,N_14962,N_14944);
nand UO_756 (O_756,N_14917,N_14850);
nand UO_757 (O_757,N_14870,N_14897);
nor UO_758 (O_758,N_14857,N_14924);
xnor UO_759 (O_759,N_14932,N_14963);
nand UO_760 (O_760,N_14877,N_14908);
xnor UO_761 (O_761,N_14907,N_14880);
xnor UO_762 (O_762,N_14862,N_14962);
nand UO_763 (O_763,N_14866,N_14879);
nand UO_764 (O_764,N_14989,N_14993);
xnor UO_765 (O_765,N_14937,N_14890);
and UO_766 (O_766,N_14852,N_14983);
nor UO_767 (O_767,N_14951,N_14870);
or UO_768 (O_768,N_14889,N_14992);
and UO_769 (O_769,N_14997,N_14989);
nor UO_770 (O_770,N_14920,N_14902);
nand UO_771 (O_771,N_14977,N_14932);
nor UO_772 (O_772,N_14991,N_14879);
and UO_773 (O_773,N_14917,N_14868);
nor UO_774 (O_774,N_14927,N_14901);
or UO_775 (O_775,N_14874,N_14877);
nand UO_776 (O_776,N_14901,N_14869);
nor UO_777 (O_777,N_14858,N_14935);
xnor UO_778 (O_778,N_14932,N_14882);
and UO_779 (O_779,N_14915,N_14942);
or UO_780 (O_780,N_14934,N_14995);
nor UO_781 (O_781,N_14983,N_14975);
and UO_782 (O_782,N_14875,N_14855);
nor UO_783 (O_783,N_14886,N_14862);
xnor UO_784 (O_784,N_14904,N_14925);
xnor UO_785 (O_785,N_14918,N_14920);
or UO_786 (O_786,N_14894,N_14907);
xor UO_787 (O_787,N_14989,N_14924);
or UO_788 (O_788,N_14925,N_14862);
and UO_789 (O_789,N_14919,N_14982);
nand UO_790 (O_790,N_14924,N_14850);
and UO_791 (O_791,N_14865,N_14984);
or UO_792 (O_792,N_14875,N_14992);
or UO_793 (O_793,N_14861,N_14963);
xor UO_794 (O_794,N_14958,N_14923);
nor UO_795 (O_795,N_14897,N_14930);
xor UO_796 (O_796,N_14863,N_14947);
xnor UO_797 (O_797,N_14922,N_14866);
and UO_798 (O_798,N_14870,N_14922);
or UO_799 (O_799,N_14969,N_14951);
nand UO_800 (O_800,N_14950,N_14965);
or UO_801 (O_801,N_14931,N_14972);
and UO_802 (O_802,N_14908,N_14876);
or UO_803 (O_803,N_14956,N_14911);
and UO_804 (O_804,N_14969,N_14943);
nor UO_805 (O_805,N_14855,N_14951);
nand UO_806 (O_806,N_14863,N_14864);
and UO_807 (O_807,N_14935,N_14947);
nor UO_808 (O_808,N_14980,N_14900);
nor UO_809 (O_809,N_14922,N_14967);
xor UO_810 (O_810,N_14861,N_14865);
nor UO_811 (O_811,N_14932,N_14979);
or UO_812 (O_812,N_14889,N_14935);
nor UO_813 (O_813,N_14977,N_14965);
or UO_814 (O_814,N_14988,N_14867);
nand UO_815 (O_815,N_14911,N_14891);
nor UO_816 (O_816,N_14987,N_14864);
and UO_817 (O_817,N_14966,N_14997);
or UO_818 (O_818,N_14990,N_14933);
or UO_819 (O_819,N_14969,N_14919);
nand UO_820 (O_820,N_14904,N_14928);
and UO_821 (O_821,N_14952,N_14885);
xor UO_822 (O_822,N_14982,N_14911);
xnor UO_823 (O_823,N_14892,N_14965);
nor UO_824 (O_824,N_14942,N_14903);
and UO_825 (O_825,N_14859,N_14973);
or UO_826 (O_826,N_14876,N_14907);
and UO_827 (O_827,N_14994,N_14990);
and UO_828 (O_828,N_14979,N_14853);
nor UO_829 (O_829,N_14870,N_14911);
nor UO_830 (O_830,N_14900,N_14907);
and UO_831 (O_831,N_14970,N_14878);
and UO_832 (O_832,N_14854,N_14915);
xor UO_833 (O_833,N_14951,N_14879);
nand UO_834 (O_834,N_14962,N_14894);
nor UO_835 (O_835,N_14985,N_14941);
xor UO_836 (O_836,N_14965,N_14861);
and UO_837 (O_837,N_14944,N_14946);
nand UO_838 (O_838,N_14870,N_14971);
xnor UO_839 (O_839,N_14941,N_14998);
and UO_840 (O_840,N_14919,N_14976);
or UO_841 (O_841,N_14940,N_14886);
xnor UO_842 (O_842,N_14920,N_14992);
nand UO_843 (O_843,N_14907,N_14909);
nor UO_844 (O_844,N_14864,N_14970);
nor UO_845 (O_845,N_14871,N_14991);
nor UO_846 (O_846,N_14930,N_14960);
and UO_847 (O_847,N_14969,N_14855);
and UO_848 (O_848,N_14873,N_14910);
xor UO_849 (O_849,N_14923,N_14959);
nand UO_850 (O_850,N_14927,N_14971);
and UO_851 (O_851,N_14863,N_14880);
or UO_852 (O_852,N_14927,N_14885);
and UO_853 (O_853,N_14892,N_14961);
nor UO_854 (O_854,N_14910,N_14893);
and UO_855 (O_855,N_14919,N_14991);
nor UO_856 (O_856,N_14875,N_14909);
nand UO_857 (O_857,N_14976,N_14973);
nand UO_858 (O_858,N_14862,N_14985);
or UO_859 (O_859,N_14982,N_14864);
xnor UO_860 (O_860,N_14937,N_14858);
or UO_861 (O_861,N_14954,N_14955);
nand UO_862 (O_862,N_14890,N_14912);
or UO_863 (O_863,N_14954,N_14971);
xor UO_864 (O_864,N_14927,N_14879);
xor UO_865 (O_865,N_14903,N_14920);
and UO_866 (O_866,N_14877,N_14879);
nand UO_867 (O_867,N_14998,N_14950);
xnor UO_868 (O_868,N_14961,N_14914);
nand UO_869 (O_869,N_14850,N_14985);
nor UO_870 (O_870,N_14942,N_14979);
nand UO_871 (O_871,N_14900,N_14944);
xnor UO_872 (O_872,N_14872,N_14988);
xor UO_873 (O_873,N_14854,N_14861);
xnor UO_874 (O_874,N_14910,N_14946);
and UO_875 (O_875,N_14936,N_14883);
nor UO_876 (O_876,N_14964,N_14894);
xnor UO_877 (O_877,N_14990,N_14942);
nor UO_878 (O_878,N_14893,N_14973);
or UO_879 (O_879,N_14964,N_14961);
xnor UO_880 (O_880,N_14956,N_14976);
and UO_881 (O_881,N_14854,N_14966);
nor UO_882 (O_882,N_14867,N_14917);
or UO_883 (O_883,N_14962,N_14956);
and UO_884 (O_884,N_14872,N_14990);
and UO_885 (O_885,N_14950,N_14943);
nor UO_886 (O_886,N_14992,N_14898);
and UO_887 (O_887,N_14882,N_14910);
xor UO_888 (O_888,N_14900,N_14913);
nand UO_889 (O_889,N_14908,N_14892);
and UO_890 (O_890,N_14958,N_14937);
xnor UO_891 (O_891,N_14916,N_14903);
or UO_892 (O_892,N_14939,N_14857);
and UO_893 (O_893,N_14902,N_14974);
xor UO_894 (O_894,N_14954,N_14970);
or UO_895 (O_895,N_14919,N_14899);
xor UO_896 (O_896,N_14927,N_14967);
nand UO_897 (O_897,N_14952,N_14893);
nor UO_898 (O_898,N_14853,N_14987);
nand UO_899 (O_899,N_14909,N_14938);
or UO_900 (O_900,N_14933,N_14951);
nor UO_901 (O_901,N_14928,N_14974);
or UO_902 (O_902,N_14952,N_14973);
xnor UO_903 (O_903,N_14854,N_14877);
or UO_904 (O_904,N_14992,N_14916);
xnor UO_905 (O_905,N_14934,N_14860);
nor UO_906 (O_906,N_14894,N_14994);
and UO_907 (O_907,N_14916,N_14977);
or UO_908 (O_908,N_14886,N_14958);
and UO_909 (O_909,N_14988,N_14919);
nand UO_910 (O_910,N_14896,N_14959);
nor UO_911 (O_911,N_14918,N_14990);
nand UO_912 (O_912,N_14988,N_14994);
nor UO_913 (O_913,N_14983,N_14903);
and UO_914 (O_914,N_14961,N_14905);
nand UO_915 (O_915,N_14934,N_14870);
xor UO_916 (O_916,N_14864,N_14973);
xnor UO_917 (O_917,N_14976,N_14934);
xnor UO_918 (O_918,N_14882,N_14914);
or UO_919 (O_919,N_14869,N_14944);
nand UO_920 (O_920,N_14950,N_14992);
nor UO_921 (O_921,N_14873,N_14940);
and UO_922 (O_922,N_14888,N_14866);
xnor UO_923 (O_923,N_14863,N_14920);
nor UO_924 (O_924,N_14990,N_14876);
nor UO_925 (O_925,N_14873,N_14866);
xor UO_926 (O_926,N_14894,N_14981);
nand UO_927 (O_927,N_14894,N_14854);
xnor UO_928 (O_928,N_14907,N_14991);
and UO_929 (O_929,N_14888,N_14973);
and UO_930 (O_930,N_14855,N_14949);
nor UO_931 (O_931,N_14883,N_14997);
nand UO_932 (O_932,N_14942,N_14986);
nor UO_933 (O_933,N_14992,N_14993);
nor UO_934 (O_934,N_14861,N_14943);
nor UO_935 (O_935,N_14902,N_14858);
and UO_936 (O_936,N_14907,N_14925);
nand UO_937 (O_937,N_14854,N_14945);
xor UO_938 (O_938,N_14998,N_14974);
nand UO_939 (O_939,N_14850,N_14986);
xor UO_940 (O_940,N_14993,N_14874);
xor UO_941 (O_941,N_14944,N_14927);
or UO_942 (O_942,N_14918,N_14868);
and UO_943 (O_943,N_14916,N_14923);
xnor UO_944 (O_944,N_14980,N_14909);
nand UO_945 (O_945,N_14896,N_14898);
xnor UO_946 (O_946,N_14964,N_14921);
or UO_947 (O_947,N_14940,N_14990);
xor UO_948 (O_948,N_14863,N_14896);
and UO_949 (O_949,N_14975,N_14944);
xor UO_950 (O_950,N_14862,N_14970);
or UO_951 (O_951,N_14867,N_14960);
nand UO_952 (O_952,N_14992,N_14850);
nor UO_953 (O_953,N_14952,N_14972);
or UO_954 (O_954,N_14974,N_14930);
or UO_955 (O_955,N_14902,N_14883);
xnor UO_956 (O_956,N_14897,N_14902);
nand UO_957 (O_957,N_14859,N_14931);
xnor UO_958 (O_958,N_14856,N_14917);
or UO_959 (O_959,N_14960,N_14850);
xnor UO_960 (O_960,N_14913,N_14919);
or UO_961 (O_961,N_14928,N_14906);
nand UO_962 (O_962,N_14880,N_14887);
nor UO_963 (O_963,N_14972,N_14854);
xor UO_964 (O_964,N_14959,N_14976);
and UO_965 (O_965,N_14888,N_14966);
nor UO_966 (O_966,N_14988,N_14957);
nor UO_967 (O_967,N_14929,N_14970);
and UO_968 (O_968,N_14965,N_14901);
nor UO_969 (O_969,N_14865,N_14855);
and UO_970 (O_970,N_14852,N_14882);
nor UO_971 (O_971,N_14854,N_14946);
and UO_972 (O_972,N_14912,N_14901);
nor UO_973 (O_973,N_14877,N_14890);
nor UO_974 (O_974,N_14874,N_14892);
nor UO_975 (O_975,N_14897,N_14866);
and UO_976 (O_976,N_14925,N_14957);
nor UO_977 (O_977,N_14953,N_14875);
nand UO_978 (O_978,N_14989,N_14862);
xnor UO_979 (O_979,N_14888,N_14912);
or UO_980 (O_980,N_14867,N_14928);
nand UO_981 (O_981,N_14896,N_14960);
or UO_982 (O_982,N_14857,N_14953);
or UO_983 (O_983,N_14910,N_14894);
xor UO_984 (O_984,N_14874,N_14907);
nand UO_985 (O_985,N_14937,N_14999);
or UO_986 (O_986,N_14967,N_14886);
or UO_987 (O_987,N_14965,N_14920);
xor UO_988 (O_988,N_14993,N_14856);
or UO_989 (O_989,N_14911,N_14987);
xnor UO_990 (O_990,N_14926,N_14974);
nand UO_991 (O_991,N_14853,N_14867);
or UO_992 (O_992,N_14936,N_14964);
nand UO_993 (O_993,N_14899,N_14979);
and UO_994 (O_994,N_14924,N_14958);
or UO_995 (O_995,N_14898,N_14854);
nor UO_996 (O_996,N_14984,N_14870);
nor UO_997 (O_997,N_14963,N_14943);
nand UO_998 (O_998,N_14892,N_14962);
nor UO_999 (O_999,N_14981,N_14924);
xor UO_1000 (O_1000,N_14946,N_14855);
xor UO_1001 (O_1001,N_14881,N_14851);
nor UO_1002 (O_1002,N_14863,N_14970);
and UO_1003 (O_1003,N_14950,N_14941);
and UO_1004 (O_1004,N_14863,N_14911);
or UO_1005 (O_1005,N_14935,N_14975);
and UO_1006 (O_1006,N_14950,N_14868);
nand UO_1007 (O_1007,N_14958,N_14893);
or UO_1008 (O_1008,N_14864,N_14939);
and UO_1009 (O_1009,N_14920,N_14990);
nand UO_1010 (O_1010,N_14980,N_14863);
nand UO_1011 (O_1011,N_14893,N_14986);
nand UO_1012 (O_1012,N_14997,N_14860);
and UO_1013 (O_1013,N_14974,N_14931);
nand UO_1014 (O_1014,N_14940,N_14949);
nand UO_1015 (O_1015,N_14933,N_14869);
nand UO_1016 (O_1016,N_14912,N_14962);
or UO_1017 (O_1017,N_14925,N_14902);
nor UO_1018 (O_1018,N_14991,N_14861);
nor UO_1019 (O_1019,N_14893,N_14960);
or UO_1020 (O_1020,N_14898,N_14878);
and UO_1021 (O_1021,N_14951,N_14994);
nand UO_1022 (O_1022,N_14857,N_14963);
xnor UO_1023 (O_1023,N_14880,N_14993);
nor UO_1024 (O_1024,N_14963,N_14895);
or UO_1025 (O_1025,N_14969,N_14972);
and UO_1026 (O_1026,N_14919,N_14858);
or UO_1027 (O_1027,N_14961,N_14922);
and UO_1028 (O_1028,N_14860,N_14888);
xnor UO_1029 (O_1029,N_14899,N_14941);
xor UO_1030 (O_1030,N_14969,N_14956);
xor UO_1031 (O_1031,N_14989,N_14916);
xor UO_1032 (O_1032,N_14999,N_14992);
nor UO_1033 (O_1033,N_14934,N_14958);
or UO_1034 (O_1034,N_14955,N_14977);
nor UO_1035 (O_1035,N_14957,N_14860);
xnor UO_1036 (O_1036,N_14973,N_14889);
nor UO_1037 (O_1037,N_14983,N_14877);
or UO_1038 (O_1038,N_14878,N_14868);
nand UO_1039 (O_1039,N_14969,N_14858);
and UO_1040 (O_1040,N_14943,N_14853);
or UO_1041 (O_1041,N_14853,N_14850);
nor UO_1042 (O_1042,N_14934,N_14868);
nand UO_1043 (O_1043,N_14916,N_14946);
or UO_1044 (O_1044,N_14908,N_14852);
nand UO_1045 (O_1045,N_14939,N_14955);
xor UO_1046 (O_1046,N_14945,N_14987);
nor UO_1047 (O_1047,N_14853,N_14976);
or UO_1048 (O_1048,N_14980,N_14936);
xor UO_1049 (O_1049,N_14994,N_14968);
xnor UO_1050 (O_1050,N_14971,N_14996);
or UO_1051 (O_1051,N_14893,N_14856);
or UO_1052 (O_1052,N_14903,N_14890);
xor UO_1053 (O_1053,N_14905,N_14963);
xor UO_1054 (O_1054,N_14962,N_14919);
and UO_1055 (O_1055,N_14972,N_14928);
nor UO_1056 (O_1056,N_14869,N_14915);
or UO_1057 (O_1057,N_14867,N_14987);
nor UO_1058 (O_1058,N_14975,N_14992);
nand UO_1059 (O_1059,N_14920,N_14985);
xor UO_1060 (O_1060,N_14902,N_14861);
nand UO_1061 (O_1061,N_14946,N_14920);
nor UO_1062 (O_1062,N_14939,N_14875);
xnor UO_1063 (O_1063,N_14932,N_14893);
and UO_1064 (O_1064,N_14912,N_14942);
or UO_1065 (O_1065,N_14882,N_14980);
and UO_1066 (O_1066,N_14977,N_14877);
xor UO_1067 (O_1067,N_14944,N_14904);
xnor UO_1068 (O_1068,N_14854,N_14984);
and UO_1069 (O_1069,N_14939,N_14874);
nor UO_1070 (O_1070,N_14893,N_14899);
xnor UO_1071 (O_1071,N_14904,N_14919);
and UO_1072 (O_1072,N_14870,N_14886);
nor UO_1073 (O_1073,N_14945,N_14954);
or UO_1074 (O_1074,N_14948,N_14884);
and UO_1075 (O_1075,N_14960,N_14879);
and UO_1076 (O_1076,N_14990,N_14938);
xnor UO_1077 (O_1077,N_14967,N_14865);
nand UO_1078 (O_1078,N_14910,N_14897);
and UO_1079 (O_1079,N_14893,N_14940);
xnor UO_1080 (O_1080,N_14894,N_14995);
or UO_1081 (O_1081,N_14953,N_14866);
and UO_1082 (O_1082,N_14928,N_14979);
xnor UO_1083 (O_1083,N_14987,N_14949);
nor UO_1084 (O_1084,N_14986,N_14886);
or UO_1085 (O_1085,N_14863,N_14939);
or UO_1086 (O_1086,N_14998,N_14946);
and UO_1087 (O_1087,N_14942,N_14923);
nand UO_1088 (O_1088,N_14987,N_14943);
and UO_1089 (O_1089,N_14870,N_14891);
and UO_1090 (O_1090,N_14995,N_14986);
xnor UO_1091 (O_1091,N_14912,N_14910);
or UO_1092 (O_1092,N_14983,N_14996);
nand UO_1093 (O_1093,N_14940,N_14997);
or UO_1094 (O_1094,N_14912,N_14946);
or UO_1095 (O_1095,N_14889,N_14936);
or UO_1096 (O_1096,N_14892,N_14907);
xnor UO_1097 (O_1097,N_14889,N_14969);
and UO_1098 (O_1098,N_14898,N_14945);
xnor UO_1099 (O_1099,N_14926,N_14870);
xnor UO_1100 (O_1100,N_14965,N_14960);
xor UO_1101 (O_1101,N_14858,N_14903);
or UO_1102 (O_1102,N_14873,N_14876);
or UO_1103 (O_1103,N_14974,N_14978);
nand UO_1104 (O_1104,N_14950,N_14888);
and UO_1105 (O_1105,N_14857,N_14882);
xor UO_1106 (O_1106,N_14904,N_14888);
nor UO_1107 (O_1107,N_14863,N_14926);
and UO_1108 (O_1108,N_14876,N_14956);
nor UO_1109 (O_1109,N_14905,N_14953);
or UO_1110 (O_1110,N_14911,N_14925);
and UO_1111 (O_1111,N_14930,N_14873);
nor UO_1112 (O_1112,N_14862,N_14923);
and UO_1113 (O_1113,N_14919,N_14972);
nand UO_1114 (O_1114,N_14892,N_14893);
or UO_1115 (O_1115,N_14978,N_14956);
and UO_1116 (O_1116,N_14986,N_14903);
xor UO_1117 (O_1117,N_14992,N_14980);
or UO_1118 (O_1118,N_14968,N_14943);
nor UO_1119 (O_1119,N_14992,N_14995);
or UO_1120 (O_1120,N_14912,N_14919);
or UO_1121 (O_1121,N_14869,N_14893);
or UO_1122 (O_1122,N_14873,N_14922);
xnor UO_1123 (O_1123,N_14924,N_14979);
or UO_1124 (O_1124,N_14865,N_14979);
xor UO_1125 (O_1125,N_14931,N_14988);
nand UO_1126 (O_1126,N_14912,N_14872);
and UO_1127 (O_1127,N_14900,N_14859);
or UO_1128 (O_1128,N_14875,N_14990);
nand UO_1129 (O_1129,N_14960,N_14954);
and UO_1130 (O_1130,N_14962,N_14921);
and UO_1131 (O_1131,N_14970,N_14999);
xnor UO_1132 (O_1132,N_14994,N_14954);
xnor UO_1133 (O_1133,N_14949,N_14931);
nor UO_1134 (O_1134,N_14931,N_14858);
or UO_1135 (O_1135,N_14857,N_14863);
and UO_1136 (O_1136,N_14898,N_14868);
or UO_1137 (O_1137,N_14868,N_14923);
nand UO_1138 (O_1138,N_14854,N_14983);
and UO_1139 (O_1139,N_14970,N_14949);
nand UO_1140 (O_1140,N_14951,N_14978);
and UO_1141 (O_1141,N_14980,N_14869);
and UO_1142 (O_1142,N_14878,N_14873);
nand UO_1143 (O_1143,N_14961,N_14975);
nand UO_1144 (O_1144,N_14969,N_14878);
xor UO_1145 (O_1145,N_14868,N_14870);
or UO_1146 (O_1146,N_14947,N_14948);
xnor UO_1147 (O_1147,N_14854,N_14912);
xnor UO_1148 (O_1148,N_14909,N_14882);
and UO_1149 (O_1149,N_14895,N_14989);
nand UO_1150 (O_1150,N_14982,N_14859);
nor UO_1151 (O_1151,N_14892,N_14952);
or UO_1152 (O_1152,N_14851,N_14890);
nand UO_1153 (O_1153,N_14917,N_14957);
or UO_1154 (O_1154,N_14940,N_14982);
nor UO_1155 (O_1155,N_14929,N_14995);
nand UO_1156 (O_1156,N_14961,N_14913);
xnor UO_1157 (O_1157,N_14938,N_14970);
nor UO_1158 (O_1158,N_14855,N_14869);
and UO_1159 (O_1159,N_14874,N_14950);
and UO_1160 (O_1160,N_14922,N_14898);
xnor UO_1161 (O_1161,N_14959,N_14852);
xnor UO_1162 (O_1162,N_14891,N_14982);
or UO_1163 (O_1163,N_14940,N_14861);
nor UO_1164 (O_1164,N_14923,N_14998);
and UO_1165 (O_1165,N_14914,N_14863);
nor UO_1166 (O_1166,N_14898,N_14946);
nor UO_1167 (O_1167,N_14919,N_14968);
nor UO_1168 (O_1168,N_14914,N_14938);
xor UO_1169 (O_1169,N_14976,N_14957);
nor UO_1170 (O_1170,N_14897,N_14884);
xor UO_1171 (O_1171,N_14981,N_14975);
xnor UO_1172 (O_1172,N_14887,N_14900);
xor UO_1173 (O_1173,N_14963,N_14891);
or UO_1174 (O_1174,N_14910,N_14970);
xor UO_1175 (O_1175,N_14854,N_14962);
and UO_1176 (O_1176,N_14981,N_14900);
or UO_1177 (O_1177,N_14989,N_14952);
or UO_1178 (O_1178,N_14988,N_14925);
xor UO_1179 (O_1179,N_14983,N_14950);
or UO_1180 (O_1180,N_14936,N_14891);
nor UO_1181 (O_1181,N_14990,N_14893);
and UO_1182 (O_1182,N_14899,N_14872);
xor UO_1183 (O_1183,N_14873,N_14953);
nand UO_1184 (O_1184,N_14869,N_14967);
nor UO_1185 (O_1185,N_14894,N_14978);
and UO_1186 (O_1186,N_14925,N_14854);
and UO_1187 (O_1187,N_14987,N_14981);
nand UO_1188 (O_1188,N_14986,N_14858);
nor UO_1189 (O_1189,N_14973,N_14913);
nor UO_1190 (O_1190,N_14979,N_14869);
or UO_1191 (O_1191,N_14879,N_14873);
nor UO_1192 (O_1192,N_14945,N_14911);
nor UO_1193 (O_1193,N_14974,N_14948);
xor UO_1194 (O_1194,N_14883,N_14950);
and UO_1195 (O_1195,N_14868,N_14911);
xor UO_1196 (O_1196,N_14954,N_14940);
nand UO_1197 (O_1197,N_14933,N_14999);
nand UO_1198 (O_1198,N_14906,N_14993);
and UO_1199 (O_1199,N_14999,N_14856);
nand UO_1200 (O_1200,N_14973,N_14947);
nand UO_1201 (O_1201,N_14876,N_14965);
and UO_1202 (O_1202,N_14926,N_14856);
nand UO_1203 (O_1203,N_14965,N_14856);
or UO_1204 (O_1204,N_14984,N_14868);
nor UO_1205 (O_1205,N_14876,N_14905);
nand UO_1206 (O_1206,N_14862,N_14937);
or UO_1207 (O_1207,N_14987,N_14927);
nor UO_1208 (O_1208,N_14939,N_14876);
xor UO_1209 (O_1209,N_14939,N_14886);
nand UO_1210 (O_1210,N_14942,N_14850);
nor UO_1211 (O_1211,N_14929,N_14866);
or UO_1212 (O_1212,N_14996,N_14863);
nand UO_1213 (O_1213,N_14946,N_14927);
xnor UO_1214 (O_1214,N_14966,N_14904);
nand UO_1215 (O_1215,N_14959,N_14911);
xor UO_1216 (O_1216,N_14960,N_14932);
nor UO_1217 (O_1217,N_14993,N_14933);
and UO_1218 (O_1218,N_14926,N_14872);
nand UO_1219 (O_1219,N_14951,N_14998);
or UO_1220 (O_1220,N_14898,N_14981);
xor UO_1221 (O_1221,N_14978,N_14897);
and UO_1222 (O_1222,N_14909,N_14946);
nand UO_1223 (O_1223,N_14878,N_14937);
xor UO_1224 (O_1224,N_14900,N_14852);
or UO_1225 (O_1225,N_14919,N_14878);
or UO_1226 (O_1226,N_14936,N_14942);
xor UO_1227 (O_1227,N_14960,N_14910);
and UO_1228 (O_1228,N_14886,N_14898);
nand UO_1229 (O_1229,N_14900,N_14974);
or UO_1230 (O_1230,N_14931,N_14880);
nand UO_1231 (O_1231,N_14861,N_14990);
or UO_1232 (O_1232,N_14883,N_14851);
nand UO_1233 (O_1233,N_14908,N_14895);
nand UO_1234 (O_1234,N_14935,N_14925);
nand UO_1235 (O_1235,N_14947,N_14893);
and UO_1236 (O_1236,N_14956,N_14924);
nor UO_1237 (O_1237,N_14923,N_14864);
nand UO_1238 (O_1238,N_14941,N_14958);
nand UO_1239 (O_1239,N_14986,N_14922);
or UO_1240 (O_1240,N_14883,N_14852);
nor UO_1241 (O_1241,N_14923,N_14981);
or UO_1242 (O_1242,N_14851,N_14941);
nand UO_1243 (O_1243,N_14969,N_14938);
xor UO_1244 (O_1244,N_14893,N_14917);
or UO_1245 (O_1245,N_14998,N_14861);
or UO_1246 (O_1246,N_14985,N_14932);
and UO_1247 (O_1247,N_14964,N_14922);
or UO_1248 (O_1248,N_14952,N_14961);
nand UO_1249 (O_1249,N_14944,N_14916);
nor UO_1250 (O_1250,N_14866,N_14891);
xor UO_1251 (O_1251,N_14998,N_14986);
xnor UO_1252 (O_1252,N_14870,N_14873);
xnor UO_1253 (O_1253,N_14876,N_14877);
and UO_1254 (O_1254,N_14906,N_14874);
nand UO_1255 (O_1255,N_14897,N_14887);
xnor UO_1256 (O_1256,N_14935,N_14860);
nand UO_1257 (O_1257,N_14861,N_14852);
and UO_1258 (O_1258,N_14989,N_14991);
nor UO_1259 (O_1259,N_14911,N_14889);
or UO_1260 (O_1260,N_14883,N_14992);
xnor UO_1261 (O_1261,N_14900,N_14901);
nand UO_1262 (O_1262,N_14986,N_14992);
nand UO_1263 (O_1263,N_14940,N_14946);
or UO_1264 (O_1264,N_14936,N_14857);
xor UO_1265 (O_1265,N_14958,N_14865);
or UO_1266 (O_1266,N_14931,N_14868);
or UO_1267 (O_1267,N_14963,N_14907);
or UO_1268 (O_1268,N_14996,N_14901);
nand UO_1269 (O_1269,N_14937,N_14926);
and UO_1270 (O_1270,N_14975,N_14943);
and UO_1271 (O_1271,N_14917,N_14921);
and UO_1272 (O_1272,N_14932,N_14876);
nor UO_1273 (O_1273,N_14987,N_14888);
or UO_1274 (O_1274,N_14889,N_14882);
nand UO_1275 (O_1275,N_14950,N_14961);
and UO_1276 (O_1276,N_14913,N_14987);
xor UO_1277 (O_1277,N_14999,N_14875);
nand UO_1278 (O_1278,N_14928,N_14870);
nand UO_1279 (O_1279,N_14975,N_14916);
nor UO_1280 (O_1280,N_14897,N_14888);
nor UO_1281 (O_1281,N_14962,N_14985);
nor UO_1282 (O_1282,N_14937,N_14959);
nor UO_1283 (O_1283,N_14978,N_14979);
xnor UO_1284 (O_1284,N_14877,N_14907);
xnor UO_1285 (O_1285,N_14907,N_14884);
xor UO_1286 (O_1286,N_14969,N_14994);
or UO_1287 (O_1287,N_14907,N_14930);
nand UO_1288 (O_1288,N_14930,N_14973);
nor UO_1289 (O_1289,N_14887,N_14980);
or UO_1290 (O_1290,N_14941,N_14916);
xor UO_1291 (O_1291,N_14983,N_14987);
or UO_1292 (O_1292,N_14891,N_14893);
xor UO_1293 (O_1293,N_14985,N_14897);
and UO_1294 (O_1294,N_14948,N_14871);
or UO_1295 (O_1295,N_14955,N_14950);
or UO_1296 (O_1296,N_14931,N_14981);
and UO_1297 (O_1297,N_14852,N_14885);
nand UO_1298 (O_1298,N_14918,N_14921);
or UO_1299 (O_1299,N_14966,N_14979);
and UO_1300 (O_1300,N_14886,N_14917);
or UO_1301 (O_1301,N_14944,N_14971);
and UO_1302 (O_1302,N_14956,N_14880);
or UO_1303 (O_1303,N_14854,N_14968);
and UO_1304 (O_1304,N_14916,N_14861);
nand UO_1305 (O_1305,N_14976,N_14851);
nor UO_1306 (O_1306,N_14863,N_14874);
nor UO_1307 (O_1307,N_14924,N_14983);
nor UO_1308 (O_1308,N_14993,N_14897);
nor UO_1309 (O_1309,N_14897,N_14879);
and UO_1310 (O_1310,N_14912,N_14992);
nor UO_1311 (O_1311,N_14969,N_14867);
and UO_1312 (O_1312,N_14914,N_14970);
nand UO_1313 (O_1313,N_14877,N_14895);
xnor UO_1314 (O_1314,N_14855,N_14885);
xor UO_1315 (O_1315,N_14908,N_14896);
and UO_1316 (O_1316,N_14898,N_14865);
and UO_1317 (O_1317,N_14893,N_14954);
xor UO_1318 (O_1318,N_14913,N_14852);
xor UO_1319 (O_1319,N_14953,N_14987);
and UO_1320 (O_1320,N_14879,N_14964);
xnor UO_1321 (O_1321,N_14923,N_14873);
or UO_1322 (O_1322,N_14974,N_14927);
or UO_1323 (O_1323,N_14958,N_14998);
or UO_1324 (O_1324,N_14918,N_14861);
and UO_1325 (O_1325,N_14931,N_14878);
xnor UO_1326 (O_1326,N_14926,N_14973);
or UO_1327 (O_1327,N_14905,N_14958);
and UO_1328 (O_1328,N_14886,N_14873);
and UO_1329 (O_1329,N_14957,N_14948);
nand UO_1330 (O_1330,N_14948,N_14889);
and UO_1331 (O_1331,N_14927,N_14960);
and UO_1332 (O_1332,N_14947,N_14995);
and UO_1333 (O_1333,N_14997,N_14970);
nand UO_1334 (O_1334,N_14910,N_14962);
nand UO_1335 (O_1335,N_14929,N_14864);
nor UO_1336 (O_1336,N_14983,N_14861);
xor UO_1337 (O_1337,N_14972,N_14877);
and UO_1338 (O_1338,N_14895,N_14937);
and UO_1339 (O_1339,N_14879,N_14882);
and UO_1340 (O_1340,N_14938,N_14869);
nand UO_1341 (O_1341,N_14872,N_14983);
and UO_1342 (O_1342,N_14854,N_14883);
xnor UO_1343 (O_1343,N_14973,N_14866);
xor UO_1344 (O_1344,N_14869,N_14866);
nand UO_1345 (O_1345,N_14855,N_14968);
xnor UO_1346 (O_1346,N_14905,N_14855);
or UO_1347 (O_1347,N_14886,N_14968);
nand UO_1348 (O_1348,N_14880,N_14909);
nor UO_1349 (O_1349,N_14951,N_14885);
and UO_1350 (O_1350,N_14884,N_14949);
nand UO_1351 (O_1351,N_14936,N_14946);
nand UO_1352 (O_1352,N_14938,N_14945);
and UO_1353 (O_1353,N_14972,N_14935);
nor UO_1354 (O_1354,N_14931,N_14959);
nor UO_1355 (O_1355,N_14903,N_14850);
xor UO_1356 (O_1356,N_14894,N_14946);
xor UO_1357 (O_1357,N_14866,N_14942);
or UO_1358 (O_1358,N_14940,N_14937);
nand UO_1359 (O_1359,N_14969,N_14963);
nor UO_1360 (O_1360,N_14925,N_14998);
xor UO_1361 (O_1361,N_14852,N_14855);
xor UO_1362 (O_1362,N_14882,N_14878);
xnor UO_1363 (O_1363,N_14896,N_14882);
xnor UO_1364 (O_1364,N_14996,N_14885);
nor UO_1365 (O_1365,N_14938,N_14968);
or UO_1366 (O_1366,N_14985,N_14965);
nor UO_1367 (O_1367,N_14874,N_14899);
nor UO_1368 (O_1368,N_14984,N_14903);
and UO_1369 (O_1369,N_14889,N_14938);
xor UO_1370 (O_1370,N_14861,N_14867);
xnor UO_1371 (O_1371,N_14854,N_14987);
xnor UO_1372 (O_1372,N_14884,N_14971);
xor UO_1373 (O_1373,N_14997,N_14863);
nand UO_1374 (O_1374,N_14984,N_14951);
and UO_1375 (O_1375,N_14991,N_14946);
and UO_1376 (O_1376,N_14928,N_14958);
xnor UO_1377 (O_1377,N_14993,N_14936);
and UO_1378 (O_1378,N_14990,N_14923);
nand UO_1379 (O_1379,N_14931,N_14894);
or UO_1380 (O_1380,N_14950,N_14895);
or UO_1381 (O_1381,N_14997,N_14944);
and UO_1382 (O_1382,N_14960,N_14953);
or UO_1383 (O_1383,N_14963,N_14998);
nor UO_1384 (O_1384,N_14897,N_14905);
xor UO_1385 (O_1385,N_14982,N_14862);
nor UO_1386 (O_1386,N_14941,N_14936);
nor UO_1387 (O_1387,N_14883,N_14927);
nand UO_1388 (O_1388,N_14936,N_14907);
and UO_1389 (O_1389,N_14949,N_14930);
nand UO_1390 (O_1390,N_14931,N_14910);
nand UO_1391 (O_1391,N_14982,N_14990);
nor UO_1392 (O_1392,N_14856,N_14960);
xnor UO_1393 (O_1393,N_14860,N_14909);
or UO_1394 (O_1394,N_14851,N_14863);
xor UO_1395 (O_1395,N_14986,N_14948);
or UO_1396 (O_1396,N_14878,N_14861);
nor UO_1397 (O_1397,N_14975,N_14953);
nand UO_1398 (O_1398,N_14941,N_14879);
and UO_1399 (O_1399,N_14898,N_14888);
nor UO_1400 (O_1400,N_14963,N_14900);
nand UO_1401 (O_1401,N_14912,N_14883);
nor UO_1402 (O_1402,N_14990,N_14881);
and UO_1403 (O_1403,N_14952,N_14897);
xnor UO_1404 (O_1404,N_14964,N_14924);
or UO_1405 (O_1405,N_14863,N_14861);
and UO_1406 (O_1406,N_14976,N_14874);
or UO_1407 (O_1407,N_14966,N_14958);
or UO_1408 (O_1408,N_14888,N_14916);
and UO_1409 (O_1409,N_14902,N_14984);
nand UO_1410 (O_1410,N_14905,N_14860);
and UO_1411 (O_1411,N_14925,N_14903);
or UO_1412 (O_1412,N_14866,N_14954);
nand UO_1413 (O_1413,N_14863,N_14948);
xor UO_1414 (O_1414,N_14935,N_14911);
or UO_1415 (O_1415,N_14884,N_14947);
and UO_1416 (O_1416,N_14906,N_14876);
or UO_1417 (O_1417,N_14895,N_14871);
nor UO_1418 (O_1418,N_14907,N_14889);
or UO_1419 (O_1419,N_14868,N_14922);
or UO_1420 (O_1420,N_14998,N_14878);
and UO_1421 (O_1421,N_14958,N_14857);
nand UO_1422 (O_1422,N_14938,N_14890);
or UO_1423 (O_1423,N_14961,N_14957);
or UO_1424 (O_1424,N_14944,N_14871);
and UO_1425 (O_1425,N_14870,N_14993);
nand UO_1426 (O_1426,N_14998,N_14932);
xor UO_1427 (O_1427,N_14921,N_14974);
xor UO_1428 (O_1428,N_14885,N_14887);
and UO_1429 (O_1429,N_14875,N_14954);
nor UO_1430 (O_1430,N_14936,N_14933);
and UO_1431 (O_1431,N_14942,N_14876);
nand UO_1432 (O_1432,N_14929,N_14887);
nor UO_1433 (O_1433,N_14973,N_14891);
or UO_1434 (O_1434,N_14939,N_14947);
nor UO_1435 (O_1435,N_14888,N_14953);
nand UO_1436 (O_1436,N_14939,N_14956);
nor UO_1437 (O_1437,N_14916,N_14878);
nor UO_1438 (O_1438,N_14857,N_14906);
xor UO_1439 (O_1439,N_14933,N_14918);
nand UO_1440 (O_1440,N_14874,N_14922);
nor UO_1441 (O_1441,N_14860,N_14904);
xnor UO_1442 (O_1442,N_14994,N_14905);
nor UO_1443 (O_1443,N_14892,N_14855);
and UO_1444 (O_1444,N_14974,N_14905);
or UO_1445 (O_1445,N_14957,N_14850);
nand UO_1446 (O_1446,N_14879,N_14901);
and UO_1447 (O_1447,N_14915,N_14871);
nand UO_1448 (O_1448,N_14944,N_14867);
nand UO_1449 (O_1449,N_14861,N_14906);
and UO_1450 (O_1450,N_14865,N_14853);
nor UO_1451 (O_1451,N_14879,N_14906);
and UO_1452 (O_1452,N_14855,N_14863);
nor UO_1453 (O_1453,N_14956,N_14987);
xor UO_1454 (O_1454,N_14869,N_14914);
nor UO_1455 (O_1455,N_14941,N_14977);
and UO_1456 (O_1456,N_14884,N_14868);
nand UO_1457 (O_1457,N_14969,N_14978);
xnor UO_1458 (O_1458,N_14953,N_14976);
and UO_1459 (O_1459,N_14929,N_14966);
xor UO_1460 (O_1460,N_14888,N_14919);
nor UO_1461 (O_1461,N_14891,N_14966);
nor UO_1462 (O_1462,N_14912,N_14898);
nand UO_1463 (O_1463,N_14920,N_14854);
xnor UO_1464 (O_1464,N_14890,N_14872);
nor UO_1465 (O_1465,N_14973,N_14884);
or UO_1466 (O_1466,N_14960,N_14914);
nor UO_1467 (O_1467,N_14979,N_14954);
or UO_1468 (O_1468,N_14947,N_14888);
or UO_1469 (O_1469,N_14926,N_14941);
nor UO_1470 (O_1470,N_14903,N_14999);
or UO_1471 (O_1471,N_14903,N_14919);
or UO_1472 (O_1472,N_14872,N_14949);
or UO_1473 (O_1473,N_14975,N_14900);
or UO_1474 (O_1474,N_14910,N_14881);
nand UO_1475 (O_1475,N_14882,N_14916);
and UO_1476 (O_1476,N_14980,N_14940);
nor UO_1477 (O_1477,N_14933,N_14948);
nand UO_1478 (O_1478,N_14947,N_14970);
nor UO_1479 (O_1479,N_14961,N_14876);
nand UO_1480 (O_1480,N_14988,N_14860);
or UO_1481 (O_1481,N_14931,N_14977);
nand UO_1482 (O_1482,N_14877,N_14929);
nor UO_1483 (O_1483,N_14882,N_14989);
nor UO_1484 (O_1484,N_14976,N_14913);
xor UO_1485 (O_1485,N_14858,N_14876);
nand UO_1486 (O_1486,N_14951,N_14924);
nand UO_1487 (O_1487,N_14878,N_14917);
xnor UO_1488 (O_1488,N_14982,N_14958);
nand UO_1489 (O_1489,N_14928,N_14887);
and UO_1490 (O_1490,N_14868,N_14958);
xnor UO_1491 (O_1491,N_14925,N_14997);
and UO_1492 (O_1492,N_14876,N_14931);
xor UO_1493 (O_1493,N_14919,N_14867);
and UO_1494 (O_1494,N_14971,N_14965);
nor UO_1495 (O_1495,N_14975,N_14938);
and UO_1496 (O_1496,N_14926,N_14858);
or UO_1497 (O_1497,N_14988,N_14961);
nand UO_1498 (O_1498,N_14859,N_14857);
or UO_1499 (O_1499,N_14944,N_14878);
nor UO_1500 (O_1500,N_14898,N_14856);
or UO_1501 (O_1501,N_14876,N_14926);
nand UO_1502 (O_1502,N_14926,N_14989);
xnor UO_1503 (O_1503,N_14874,N_14986);
nor UO_1504 (O_1504,N_14871,N_14943);
xnor UO_1505 (O_1505,N_14934,N_14857);
nor UO_1506 (O_1506,N_14994,N_14995);
nand UO_1507 (O_1507,N_14920,N_14924);
nor UO_1508 (O_1508,N_14961,N_14903);
nand UO_1509 (O_1509,N_14865,N_14952);
or UO_1510 (O_1510,N_14911,N_14909);
nor UO_1511 (O_1511,N_14927,N_14881);
nand UO_1512 (O_1512,N_14998,N_14918);
and UO_1513 (O_1513,N_14880,N_14873);
nor UO_1514 (O_1514,N_14993,N_14952);
nor UO_1515 (O_1515,N_14989,N_14937);
xor UO_1516 (O_1516,N_14966,N_14991);
nand UO_1517 (O_1517,N_14934,N_14962);
or UO_1518 (O_1518,N_14959,N_14898);
or UO_1519 (O_1519,N_14942,N_14950);
nor UO_1520 (O_1520,N_14867,N_14868);
xor UO_1521 (O_1521,N_14973,N_14969);
xor UO_1522 (O_1522,N_14910,N_14979);
xnor UO_1523 (O_1523,N_14975,N_14866);
nor UO_1524 (O_1524,N_14994,N_14860);
or UO_1525 (O_1525,N_14900,N_14919);
xor UO_1526 (O_1526,N_14851,N_14987);
nor UO_1527 (O_1527,N_14944,N_14880);
nand UO_1528 (O_1528,N_14992,N_14966);
nand UO_1529 (O_1529,N_14991,N_14942);
xor UO_1530 (O_1530,N_14996,N_14935);
and UO_1531 (O_1531,N_14855,N_14994);
or UO_1532 (O_1532,N_14968,N_14987);
or UO_1533 (O_1533,N_14883,N_14968);
or UO_1534 (O_1534,N_14932,N_14913);
and UO_1535 (O_1535,N_14984,N_14932);
or UO_1536 (O_1536,N_14887,N_14906);
xor UO_1537 (O_1537,N_14951,N_14971);
nand UO_1538 (O_1538,N_14867,N_14953);
or UO_1539 (O_1539,N_14857,N_14896);
nand UO_1540 (O_1540,N_14937,N_14974);
xor UO_1541 (O_1541,N_14928,N_14938);
nor UO_1542 (O_1542,N_14920,N_14861);
nor UO_1543 (O_1543,N_14948,N_14900);
nand UO_1544 (O_1544,N_14979,N_14934);
and UO_1545 (O_1545,N_14945,N_14864);
xor UO_1546 (O_1546,N_14959,N_14960);
and UO_1547 (O_1547,N_14887,N_14948);
or UO_1548 (O_1548,N_14952,N_14960);
or UO_1549 (O_1549,N_14935,N_14961);
and UO_1550 (O_1550,N_14901,N_14853);
xor UO_1551 (O_1551,N_14853,N_14929);
or UO_1552 (O_1552,N_14912,N_14963);
xnor UO_1553 (O_1553,N_14867,N_14972);
xor UO_1554 (O_1554,N_14881,N_14995);
nor UO_1555 (O_1555,N_14949,N_14924);
and UO_1556 (O_1556,N_14879,N_14894);
nand UO_1557 (O_1557,N_14946,N_14963);
or UO_1558 (O_1558,N_14905,N_14926);
or UO_1559 (O_1559,N_14912,N_14921);
xnor UO_1560 (O_1560,N_14922,N_14894);
xor UO_1561 (O_1561,N_14950,N_14864);
and UO_1562 (O_1562,N_14877,N_14959);
and UO_1563 (O_1563,N_14989,N_14928);
nor UO_1564 (O_1564,N_14885,N_14850);
nand UO_1565 (O_1565,N_14896,N_14941);
xor UO_1566 (O_1566,N_14897,N_14882);
and UO_1567 (O_1567,N_14951,N_14941);
xnor UO_1568 (O_1568,N_14891,N_14975);
nor UO_1569 (O_1569,N_14956,N_14860);
and UO_1570 (O_1570,N_14992,N_14886);
xnor UO_1571 (O_1571,N_14900,N_14920);
nor UO_1572 (O_1572,N_14978,N_14896);
nor UO_1573 (O_1573,N_14861,N_14900);
xnor UO_1574 (O_1574,N_14914,N_14950);
xnor UO_1575 (O_1575,N_14939,N_14908);
or UO_1576 (O_1576,N_14932,N_14906);
and UO_1577 (O_1577,N_14937,N_14943);
nor UO_1578 (O_1578,N_14886,N_14984);
nor UO_1579 (O_1579,N_14969,N_14917);
nor UO_1580 (O_1580,N_14988,N_14901);
xor UO_1581 (O_1581,N_14858,N_14991);
and UO_1582 (O_1582,N_14886,N_14877);
or UO_1583 (O_1583,N_14861,N_14951);
and UO_1584 (O_1584,N_14885,N_14925);
or UO_1585 (O_1585,N_14888,N_14995);
and UO_1586 (O_1586,N_14876,N_14885);
nor UO_1587 (O_1587,N_14882,N_14912);
xnor UO_1588 (O_1588,N_14863,N_14906);
or UO_1589 (O_1589,N_14978,N_14934);
and UO_1590 (O_1590,N_14957,N_14955);
xnor UO_1591 (O_1591,N_14983,N_14990);
and UO_1592 (O_1592,N_14988,N_14913);
nand UO_1593 (O_1593,N_14870,N_14867);
and UO_1594 (O_1594,N_14937,N_14995);
xor UO_1595 (O_1595,N_14911,N_14941);
nor UO_1596 (O_1596,N_14870,N_14881);
and UO_1597 (O_1597,N_14948,N_14929);
or UO_1598 (O_1598,N_14905,N_14938);
nor UO_1599 (O_1599,N_14879,N_14990);
and UO_1600 (O_1600,N_14976,N_14869);
and UO_1601 (O_1601,N_14992,N_14911);
or UO_1602 (O_1602,N_14905,N_14960);
and UO_1603 (O_1603,N_14987,N_14882);
nand UO_1604 (O_1604,N_14855,N_14906);
and UO_1605 (O_1605,N_14939,N_14889);
xnor UO_1606 (O_1606,N_14981,N_14869);
nor UO_1607 (O_1607,N_14909,N_14876);
or UO_1608 (O_1608,N_14912,N_14999);
nand UO_1609 (O_1609,N_14888,N_14854);
xnor UO_1610 (O_1610,N_14870,N_14893);
nor UO_1611 (O_1611,N_14858,N_14971);
nand UO_1612 (O_1612,N_14913,N_14876);
nand UO_1613 (O_1613,N_14964,N_14937);
or UO_1614 (O_1614,N_14997,N_14979);
xnor UO_1615 (O_1615,N_14949,N_14922);
or UO_1616 (O_1616,N_14974,N_14885);
xor UO_1617 (O_1617,N_14855,N_14966);
nand UO_1618 (O_1618,N_14980,N_14875);
and UO_1619 (O_1619,N_14861,N_14933);
and UO_1620 (O_1620,N_14962,N_14914);
or UO_1621 (O_1621,N_14852,N_14909);
and UO_1622 (O_1622,N_14852,N_14952);
nand UO_1623 (O_1623,N_14924,N_14976);
nor UO_1624 (O_1624,N_14852,N_14999);
xnor UO_1625 (O_1625,N_14871,N_14888);
xnor UO_1626 (O_1626,N_14996,N_14936);
and UO_1627 (O_1627,N_14949,N_14988);
xnor UO_1628 (O_1628,N_14898,N_14884);
or UO_1629 (O_1629,N_14986,N_14967);
and UO_1630 (O_1630,N_14874,N_14852);
xnor UO_1631 (O_1631,N_14891,N_14877);
and UO_1632 (O_1632,N_14914,N_14995);
or UO_1633 (O_1633,N_14946,N_14875);
or UO_1634 (O_1634,N_14986,N_14961);
xnor UO_1635 (O_1635,N_14908,N_14925);
nand UO_1636 (O_1636,N_14885,N_14880);
nand UO_1637 (O_1637,N_14993,N_14946);
and UO_1638 (O_1638,N_14977,N_14986);
or UO_1639 (O_1639,N_14987,N_14910);
or UO_1640 (O_1640,N_14914,N_14915);
nand UO_1641 (O_1641,N_14930,N_14901);
or UO_1642 (O_1642,N_14974,N_14920);
nand UO_1643 (O_1643,N_14866,N_14972);
nand UO_1644 (O_1644,N_14968,N_14965);
nor UO_1645 (O_1645,N_14965,N_14858);
and UO_1646 (O_1646,N_14945,N_14964);
or UO_1647 (O_1647,N_14893,N_14982);
nor UO_1648 (O_1648,N_14948,N_14910);
xor UO_1649 (O_1649,N_14892,N_14980);
xor UO_1650 (O_1650,N_14958,N_14884);
or UO_1651 (O_1651,N_14918,N_14899);
nand UO_1652 (O_1652,N_14973,N_14927);
and UO_1653 (O_1653,N_14981,N_14918);
xnor UO_1654 (O_1654,N_14917,N_14982);
xnor UO_1655 (O_1655,N_14864,N_14959);
and UO_1656 (O_1656,N_14853,N_14855);
nor UO_1657 (O_1657,N_14967,N_14864);
and UO_1658 (O_1658,N_14959,N_14996);
nand UO_1659 (O_1659,N_14910,N_14888);
and UO_1660 (O_1660,N_14898,N_14929);
nand UO_1661 (O_1661,N_14945,N_14994);
or UO_1662 (O_1662,N_14922,N_14998);
or UO_1663 (O_1663,N_14908,N_14953);
nand UO_1664 (O_1664,N_14901,N_14919);
or UO_1665 (O_1665,N_14853,N_14877);
xor UO_1666 (O_1666,N_14963,N_14902);
and UO_1667 (O_1667,N_14936,N_14997);
nor UO_1668 (O_1668,N_14936,N_14962);
or UO_1669 (O_1669,N_14878,N_14940);
xor UO_1670 (O_1670,N_14875,N_14936);
nand UO_1671 (O_1671,N_14971,N_14851);
and UO_1672 (O_1672,N_14973,N_14850);
or UO_1673 (O_1673,N_14921,N_14998);
nand UO_1674 (O_1674,N_14983,N_14875);
or UO_1675 (O_1675,N_14862,N_14941);
or UO_1676 (O_1676,N_14932,N_14867);
xor UO_1677 (O_1677,N_14943,N_14976);
xor UO_1678 (O_1678,N_14876,N_14945);
xor UO_1679 (O_1679,N_14982,N_14943);
or UO_1680 (O_1680,N_14883,N_14931);
xnor UO_1681 (O_1681,N_14868,N_14972);
xor UO_1682 (O_1682,N_14931,N_14874);
and UO_1683 (O_1683,N_14974,N_14954);
or UO_1684 (O_1684,N_14886,N_14869);
or UO_1685 (O_1685,N_14923,N_14875);
nand UO_1686 (O_1686,N_14852,N_14934);
and UO_1687 (O_1687,N_14970,N_14961);
or UO_1688 (O_1688,N_14914,N_14909);
nor UO_1689 (O_1689,N_14937,N_14977);
and UO_1690 (O_1690,N_14904,N_14896);
nand UO_1691 (O_1691,N_14912,N_14933);
or UO_1692 (O_1692,N_14893,N_14920);
nor UO_1693 (O_1693,N_14971,N_14936);
nor UO_1694 (O_1694,N_14951,N_14991);
xor UO_1695 (O_1695,N_14981,N_14884);
nand UO_1696 (O_1696,N_14865,N_14905);
nor UO_1697 (O_1697,N_14927,N_14856);
and UO_1698 (O_1698,N_14879,N_14872);
xor UO_1699 (O_1699,N_14996,N_14952);
nand UO_1700 (O_1700,N_14884,N_14889);
or UO_1701 (O_1701,N_14908,N_14986);
nand UO_1702 (O_1702,N_14915,N_14894);
xor UO_1703 (O_1703,N_14891,N_14867);
xnor UO_1704 (O_1704,N_14999,N_14908);
nor UO_1705 (O_1705,N_14957,N_14989);
nor UO_1706 (O_1706,N_14935,N_14870);
or UO_1707 (O_1707,N_14963,N_14872);
or UO_1708 (O_1708,N_14888,N_14971);
xnor UO_1709 (O_1709,N_14936,N_14984);
nand UO_1710 (O_1710,N_14944,N_14859);
xor UO_1711 (O_1711,N_14957,N_14853);
xnor UO_1712 (O_1712,N_14859,N_14916);
nand UO_1713 (O_1713,N_14869,N_14878);
and UO_1714 (O_1714,N_14870,N_14890);
and UO_1715 (O_1715,N_14893,N_14971);
and UO_1716 (O_1716,N_14959,N_14983);
and UO_1717 (O_1717,N_14872,N_14967);
xnor UO_1718 (O_1718,N_14956,N_14945);
xnor UO_1719 (O_1719,N_14881,N_14855);
nand UO_1720 (O_1720,N_14911,N_14918);
or UO_1721 (O_1721,N_14867,N_14911);
nand UO_1722 (O_1722,N_14905,N_14888);
and UO_1723 (O_1723,N_14926,N_14871);
or UO_1724 (O_1724,N_14985,N_14911);
or UO_1725 (O_1725,N_14983,N_14871);
nand UO_1726 (O_1726,N_14942,N_14855);
xnor UO_1727 (O_1727,N_14969,N_14987);
nor UO_1728 (O_1728,N_14993,N_14935);
and UO_1729 (O_1729,N_14871,N_14964);
nor UO_1730 (O_1730,N_14859,N_14947);
nand UO_1731 (O_1731,N_14890,N_14956);
nand UO_1732 (O_1732,N_14906,N_14901);
or UO_1733 (O_1733,N_14886,N_14930);
nor UO_1734 (O_1734,N_14962,N_14922);
or UO_1735 (O_1735,N_14856,N_14910);
xnor UO_1736 (O_1736,N_14946,N_14853);
nor UO_1737 (O_1737,N_14930,N_14996);
or UO_1738 (O_1738,N_14931,N_14967);
nand UO_1739 (O_1739,N_14999,N_14887);
or UO_1740 (O_1740,N_14926,N_14900);
xor UO_1741 (O_1741,N_14896,N_14877);
or UO_1742 (O_1742,N_14865,N_14869);
nor UO_1743 (O_1743,N_14854,N_14937);
nor UO_1744 (O_1744,N_14941,N_14973);
nor UO_1745 (O_1745,N_14994,N_14939);
nor UO_1746 (O_1746,N_14900,N_14997);
nor UO_1747 (O_1747,N_14995,N_14985);
nand UO_1748 (O_1748,N_14852,N_14880);
xor UO_1749 (O_1749,N_14940,N_14887);
nor UO_1750 (O_1750,N_14999,N_14941);
nand UO_1751 (O_1751,N_14921,N_14915);
nor UO_1752 (O_1752,N_14956,N_14948);
or UO_1753 (O_1753,N_14882,N_14872);
nand UO_1754 (O_1754,N_14913,N_14861);
nand UO_1755 (O_1755,N_14995,N_14950);
nand UO_1756 (O_1756,N_14916,N_14873);
nor UO_1757 (O_1757,N_14946,N_14949);
nor UO_1758 (O_1758,N_14946,N_14883);
nand UO_1759 (O_1759,N_14866,N_14995);
nand UO_1760 (O_1760,N_14923,N_14972);
nand UO_1761 (O_1761,N_14870,N_14945);
xnor UO_1762 (O_1762,N_14961,N_14958);
xor UO_1763 (O_1763,N_14952,N_14945);
and UO_1764 (O_1764,N_14872,N_14911);
nand UO_1765 (O_1765,N_14918,N_14945);
nand UO_1766 (O_1766,N_14931,N_14905);
xor UO_1767 (O_1767,N_14912,N_14893);
or UO_1768 (O_1768,N_14936,N_14870);
nor UO_1769 (O_1769,N_14918,N_14970);
or UO_1770 (O_1770,N_14877,N_14863);
nand UO_1771 (O_1771,N_14948,N_14873);
or UO_1772 (O_1772,N_14989,N_14866);
nand UO_1773 (O_1773,N_14891,N_14987);
nor UO_1774 (O_1774,N_14914,N_14959);
nand UO_1775 (O_1775,N_14894,N_14969);
and UO_1776 (O_1776,N_14970,N_14927);
and UO_1777 (O_1777,N_14932,N_14877);
or UO_1778 (O_1778,N_14982,N_14853);
nor UO_1779 (O_1779,N_14875,N_14851);
nand UO_1780 (O_1780,N_14992,N_14878);
or UO_1781 (O_1781,N_14915,N_14862);
or UO_1782 (O_1782,N_14940,N_14947);
nor UO_1783 (O_1783,N_14868,N_14947);
and UO_1784 (O_1784,N_14945,N_14919);
and UO_1785 (O_1785,N_14882,N_14988);
nor UO_1786 (O_1786,N_14878,N_14939);
nand UO_1787 (O_1787,N_14902,N_14874);
xor UO_1788 (O_1788,N_14970,N_14991);
or UO_1789 (O_1789,N_14924,N_14894);
and UO_1790 (O_1790,N_14931,N_14922);
nor UO_1791 (O_1791,N_14899,N_14966);
or UO_1792 (O_1792,N_14875,N_14998);
or UO_1793 (O_1793,N_14889,N_14934);
nand UO_1794 (O_1794,N_14986,N_14952);
nor UO_1795 (O_1795,N_14995,N_14918);
or UO_1796 (O_1796,N_14935,N_14909);
and UO_1797 (O_1797,N_14875,N_14861);
nor UO_1798 (O_1798,N_14934,N_14987);
nor UO_1799 (O_1799,N_14954,N_14992);
xnor UO_1800 (O_1800,N_14923,N_14947);
xor UO_1801 (O_1801,N_14967,N_14911);
or UO_1802 (O_1802,N_14946,N_14911);
and UO_1803 (O_1803,N_14930,N_14869);
and UO_1804 (O_1804,N_14974,N_14960);
nand UO_1805 (O_1805,N_14953,N_14925);
xor UO_1806 (O_1806,N_14963,N_14906);
nand UO_1807 (O_1807,N_14863,N_14858);
and UO_1808 (O_1808,N_14889,N_14892);
and UO_1809 (O_1809,N_14882,N_14950);
xor UO_1810 (O_1810,N_14892,N_14920);
or UO_1811 (O_1811,N_14882,N_14993);
nand UO_1812 (O_1812,N_14998,N_14975);
and UO_1813 (O_1813,N_14950,N_14861);
and UO_1814 (O_1814,N_14940,N_14894);
or UO_1815 (O_1815,N_14898,N_14926);
and UO_1816 (O_1816,N_14869,N_14873);
or UO_1817 (O_1817,N_14955,N_14998);
or UO_1818 (O_1818,N_14969,N_14903);
xnor UO_1819 (O_1819,N_14997,N_14969);
xnor UO_1820 (O_1820,N_14968,N_14887);
nand UO_1821 (O_1821,N_14945,N_14973);
nand UO_1822 (O_1822,N_14856,N_14904);
nand UO_1823 (O_1823,N_14880,N_14966);
and UO_1824 (O_1824,N_14902,N_14865);
and UO_1825 (O_1825,N_14899,N_14929);
xnor UO_1826 (O_1826,N_14885,N_14892);
and UO_1827 (O_1827,N_14901,N_14932);
and UO_1828 (O_1828,N_14928,N_14978);
nand UO_1829 (O_1829,N_14957,N_14910);
nor UO_1830 (O_1830,N_14938,N_14932);
nor UO_1831 (O_1831,N_14858,N_14877);
or UO_1832 (O_1832,N_14995,N_14882);
nand UO_1833 (O_1833,N_14889,N_14941);
nand UO_1834 (O_1834,N_14896,N_14899);
xnor UO_1835 (O_1835,N_14904,N_14880);
xnor UO_1836 (O_1836,N_14915,N_14992);
xor UO_1837 (O_1837,N_14897,N_14896);
and UO_1838 (O_1838,N_14943,N_14877);
xnor UO_1839 (O_1839,N_14971,N_14948);
nand UO_1840 (O_1840,N_14891,N_14912);
and UO_1841 (O_1841,N_14985,N_14875);
and UO_1842 (O_1842,N_14981,N_14897);
or UO_1843 (O_1843,N_14882,N_14869);
or UO_1844 (O_1844,N_14940,N_14890);
nand UO_1845 (O_1845,N_14854,N_14981);
and UO_1846 (O_1846,N_14988,N_14929);
nand UO_1847 (O_1847,N_14871,N_14970);
nor UO_1848 (O_1848,N_14913,N_14855);
nor UO_1849 (O_1849,N_14927,N_14884);
or UO_1850 (O_1850,N_14977,N_14917);
xor UO_1851 (O_1851,N_14924,N_14967);
nor UO_1852 (O_1852,N_14885,N_14904);
and UO_1853 (O_1853,N_14850,N_14994);
or UO_1854 (O_1854,N_14962,N_14953);
xor UO_1855 (O_1855,N_14899,N_14971);
nor UO_1856 (O_1856,N_14953,N_14921);
nor UO_1857 (O_1857,N_14978,N_14999);
nand UO_1858 (O_1858,N_14880,N_14992);
nand UO_1859 (O_1859,N_14891,N_14955);
or UO_1860 (O_1860,N_14957,N_14993);
nor UO_1861 (O_1861,N_14895,N_14980);
and UO_1862 (O_1862,N_14855,N_14919);
nand UO_1863 (O_1863,N_14891,N_14974);
and UO_1864 (O_1864,N_14884,N_14895);
or UO_1865 (O_1865,N_14859,N_14894);
and UO_1866 (O_1866,N_14941,N_14949);
and UO_1867 (O_1867,N_14947,N_14996);
xor UO_1868 (O_1868,N_14922,N_14975);
xor UO_1869 (O_1869,N_14942,N_14927);
nor UO_1870 (O_1870,N_14868,N_14919);
xor UO_1871 (O_1871,N_14989,N_14935);
nand UO_1872 (O_1872,N_14931,N_14963);
nand UO_1873 (O_1873,N_14979,N_14893);
or UO_1874 (O_1874,N_14922,N_14899);
nor UO_1875 (O_1875,N_14895,N_14974);
and UO_1876 (O_1876,N_14853,N_14921);
or UO_1877 (O_1877,N_14914,N_14921);
xor UO_1878 (O_1878,N_14974,N_14933);
nor UO_1879 (O_1879,N_14908,N_14965);
or UO_1880 (O_1880,N_14861,N_14985);
nand UO_1881 (O_1881,N_14982,N_14965);
or UO_1882 (O_1882,N_14916,N_14881);
xor UO_1883 (O_1883,N_14953,N_14966);
xor UO_1884 (O_1884,N_14933,N_14895);
and UO_1885 (O_1885,N_14969,N_14859);
nand UO_1886 (O_1886,N_14974,N_14950);
or UO_1887 (O_1887,N_14944,N_14951);
and UO_1888 (O_1888,N_14928,N_14988);
nor UO_1889 (O_1889,N_14941,N_14956);
or UO_1890 (O_1890,N_14879,N_14973);
nor UO_1891 (O_1891,N_14855,N_14945);
nand UO_1892 (O_1892,N_14878,N_14925);
or UO_1893 (O_1893,N_14990,N_14894);
nor UO_1894 (O_1894,N_14893,N_14934);
xnor UO_1895 (O_1895,N_14895,N_14875);
or UO_1896 (O_1896,N_14865,N_14900);
xor UO_1897 (O_1897,N_14865,N_14878);
xor UO_1898 (O_1898,N_14858,N_14966);
and UO_1899 (O_1899,N_14967,N_14974);
nand UO_1900 (O_1900,N_14974,N_14911);
xor UO_1901 (O_1901,N_14907,N_14864);
nor UO_1902 (O_1902,N_14919,N_14908);
nor UO_1903 (O_1903,N_14893,N_14862);
or UO_1904 (O_1904,N_14973,N_14932);
nand UO_1905 (O_1905,N_14902,N_14926);
and UO_1906 (O_1906,N_14983,N_14905);
or UO_1907 (O_1907,N_14978,N_14864);
or UO_1908 (O_1908,N_14984,N_14914);
and UO_1909 (O_1909,N_14920,N_14962);
xnor UO_1910 (O_1910,N_14978,N_14924);
nor UO_1911 (O_1911,N_14948,N_14984);
and UO_1912 (O_1912,N_14982,N_14851);
nand UO_1913 (O_1913,N_14872,N_14940);
or UO_1914 (O_1914,N_14976,N_14899);
xor UO_1915 (O_1915,N_14922,N_14930);
xor UO_1916 (O_1916,N_14908,N_14948);
and UO_1917 (O_1917,N_14968,N_14976);
nand UO_1918 (O_1918,N_14939,N_14887);
and UO_1919 (O_1919,N_14997,N_14886);
or UO_1920 (O_1920,N_14885,N_14902);
xnor UO_1921 (O_1921,N_14873,N_14872);
or UO_1922 (O_1922,N_14946,N_14996);
nand UO_1923 (O_1923,N_14984,N_14938);
and UO_1924 (O_1924,N_14890,N_14915);
and UO_1925 (O_1925,N_14904,N_14927);
nor UO_1926 (O_1926,N_14873,N_14924);
nor UO_1927 (O_1927,N_14883,N_14898);
and UO_1928 (O_1928,N_14964,N_14999);
and UO_1929 (O_1929,N_14961,N_14965);
nand UO_1930 (O_1930,N_14867,N_14877);
nor UO_1931 (O_1931,N_14997,N_14999);
nand UO_1932 (O_1932,N_14967,N_14918);
nand UO_1933 (O_1933,N_14959,N_14871);
and UO_1934 (O_1934,N_14959,N_14928);
or UO_1935 (O_1935,N_14899,N_14930);
or UO_1936 (O_1936,N_14952,N_14991);
and UO_1937 (O_1937,N_14994,N_14920);
or UO_1938 (O_1938,N_14894,N_14872);
nor UO_1939 (O_1939,N_14941,N_14870);
xor UO_1940 (O_1940,N_14953,N_14898);
nor UO_1941 (O_1941,N_14961,N_14936);
or UO_1942 (O_1942,N_14922,N_14881);
nor UO_1943 (O_1943,N_14961,N_14881);
nand UO_1944 (O_1944,N_14861,N_14880);
or UO_1945 (O_1945,N_14929,N_14870);
nand UO_1946 (O_1946,N_14987,N_14961);
nand UO_1947 (O_1947,N_14930,N_14988);
or UO_1948 (O_1948,N_14888,N_14921);
nand UO_1949 (O_1949,N_14977,N_14861);
and UO_1950 (O_1950,N_14973,N_14904);
and UO_1951 (O_1951,N_14939,N_14904);
nor UO_1952 (O_1952,N_14894,N_14976);
nor UO_1953 (O_1953,N_14937,N_14911);
nand UO_1954 (O_1954,N_14876,N_14896);
or UO_1955 (O_1955,N_14885,N_14856);
and UO_1956 (O_1956,N_14952,N_14962);
nand UO_1957 (O_1957,N_14901,N_14917);
nand UO_1958 (O_1958,N_14963,N_14975);
xnor UO_1959 (O_1959,N_14955,N_14983);
nand UO_1960 (O_1960,N_14992,N_14961);
nor UO_1961 (O_1961,N_14872,N_14999);
and UO_1962 (O_1962,N_14945,N_14908);
nor UO_1963 (O_1963,N_14922,N_14897);
nor UO_1964 (O_1964,N_14977,N_14979);
and UO_1965 (O_1965,N_14913,N_14975);
nand UO_1966 (O_1966,N_14967,N_14905);
nor UO_1967 (O_1967,N_14969,N_14890);
and UO_1968 (O_1968,N_14942,N_14887);
and UO_1969 (O_1969,N_14901,N_14983);
and UO_1970 (O_1970,N_14866,N_14963);
or UO_1971 (O_1971,N_14915,N_14860);
xor UO_1972 (O_1972,N_14927,N_14979);
nor UO_1973 (O_1973,N_14914,N_14957);
nor UO_1974 (O_1974,N_14889,N_14914);
or UO_1975 (O_1975,N_14971,N_14916);
nor UO_1976 (O_1976,N_14947,N_14928);
or UO_1977 (O_1977,N_14967,N_14877);
nor UO_1978 (O_1978,N_14932,N_14943);
xor UO_1979 (O_1979,N_14912,N_14987);
or UO_1980 (O_1980,N_14985,N_14992);
nand UO_1981 (O_1981,N_14992,N_14884);
or UO_1982 (O_1982,N_14900,N_14924);
and UO_1983 (O_1983,N_14899,N_14870);
nor UO_1984 (O_1984,N_14856,N_14864);
xor UO_1985 (O_1985,N_14964,N_14943);
nor UO_1986 (O_1986,N_14986,N_14972);
nor UO_1987 (O_1987,N_14926,N_14880);
and UO_1988 (O_1988,N_14951,N_14897);
xnor UO_1989 (O_1989,N_14952,N_14913);
nor UO_1990 (O_1990,N_14936,N_14913);
or UO_1991 (O_1991,N_14863,N_14850);
nand UO_1992 (O_1992,N_14926,N_14964);
nor UO_1993 (O_1993,N_14873,N_14970);
or UO_1994 (O_1994,N_14919,N_14902);
xnor UO_1995 (O_1995,N_14950,N_14930);
and UO_1996 (O_1996,N_14913,N_14882);
and UO_1997 (O_1997,N_14882,N_14966);
nand UO_1998 (O_1998,N_14974,N_14989);
xnor UO_1999 (O_1999,N_14887,N_14878);
endmodule