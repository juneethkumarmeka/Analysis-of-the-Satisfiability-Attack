module basic_1000_10000_1500_10_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_637,In_168);
nor U1 (N_1,In_409,In_965);
and U2 (N_2,In_684,In_745);
nor U3 (N_3,In_662,In_672);
and U4 (N_4,In_382,In_929);
nor U5 (N_5,In_432,In_402);
nor U6 (N_6,In_883,In_738);
or U7 (N_7,In_481,In_102);
nand U8 (N_8,In_322,In_850);
or U9 (N_9,In_593,In_868);
nand U10 (N_10,In_75,In_874);
nand U11 (N_11,In_68,In_72);
xnor U12 (N_12,In_59,In_332);
nand U13 (N_13,In_587,In_649);
and U14 (N_14,In_426,In_911);
nand U15 (N_15,In_331,In_363);
nand U16 (N_16,In_241,In_293);
nor U17 (N_17,In_209,In_132);
nand U18 (N_18,In_873,In_586);
nor U19 (N_19,In_477,In_414);
or U20 (N_20,In_324,In_595);
or U21 (N_21,In_990,In_840);
nand U22 (N_22,In_884,In_392);
nand U23 (N_23,In_664,In_216);
nand U24 (N_24,In_553,In_858);
and U25 (N_25,In_939,In_895);
or U26 (N_26,In_403,In_145);
nor U27 (N_27,In_696,In_694);
or U28 (N_28,In_786,In_615);
xor U29 (N_29,In_267,In_397);
or U30 (N_30,In_571,In_959);
nor U31 (N_31,In_940,In_314);
and U32 (N_32,In_967,In_651);
nor U33 (N_33,In_345,In_105);
and U34 (N_34,In_909,In_668);
or U35 (N_35,In_380,In_872);
or U36 (N_36,In_278,In_531);
or U37 (N_37,In_801,In_765);
nor U38 (N_38,In_435,In_635);
nor U39 (N_39,In_588,In_565);
nor U40 (N_40,In_141,In_408);
or U41 (N_41,In_761,In_783);
and U42 (N_42,In_172,In_308);
nor U43 (N_43,In_286,In_865);
or U44 (N_44,In_458,In_636);
and U45 (N_45,In_415,In_468);
nand U46 (N_46,In_576,In_735);
nand U47 (N_47,In_767,In_643);
and U48 (N_48,In_585,In_584);
or U49 (N_49,In_390,In_50);
or U50 (N_50,In_508,In_838);
and U51 (N_51,In_856,In_301);
and U52 (N_52,In_846,In_825);
nor U53 (N_53,In_712,In_474);
nor U54 (N_54,In_368,In_726);
nand U55 (N_55,In_673,In_614);
and U56 (N_56,In_600,In_741);
nor U57 (N_57,In_710,In_151);
and U58 (N_58,In_570,In_291);
nor U59 (N_59,In_357,In_289);
or U60 (N_60,In_819,In_303);
nand U61 (N_61,In_921,In_176);
nand U62 (N_62,In_70,In_193);
or U63 (N_63,In_948,In_785);
nand U64 (N_64,In_457,In_861);
nand U65 (N_65,In_628,In_416);
and U66 (N_66,In_171,In_732);
and U67 (N_67,In_894,In_487);
nand U68 (N_68,In_158,In_453);
or U69 (N_69,In_561,In_827);
and U70 (N_70,In_916,In_857);
nor U71 (N_71,In_410,In_656);
nand U72 (N_72,In_714,In_211);
or U73 (N_73,In_495,In_233);
or U74 (N_74,In_613,In_923);
nor U75 (N_75,In_796,In_279);
and U76 (N_76,In_752,In_315);
and U77 (N_77,In_904,In_455);
or U78 (N_78,In_913,In_190);
or U79 (N_79,In_890,In_52);
and U80 (N_80,In_864,In_21);
or U81 (N_81,In_244,In_483);
nand U82 (N_82,In_725,In_994);
or U83 (N_83,In_797,In_496);
nor U84 (N_84,In_67,In_356);
xor U85 (N_85,In_688,In_533);
or U86 (N_86,In_146,In_599);
nor U87 (N_87,In_442,In_339);
nor U88 (N_88,In_683,In_882);
nand U89 (N_89,In_43,In_124);
nand U90 (N_90,In_138,In_762);
nor U91 (N_91,In_606,In_104);
nand U92 (N_92,In_790,In_309);
and U93 (N_93,In_343,In_37);
nand U94 (N_94,In_731,In_188);
or U95 (N_95,In_659,In_969);
or U96 (N_96,In_706,In_154);
nor U97 (N_97,In_80,In_754);
nor U98 (N_98,In_552,In_54);
or U99 (N_99,In_33,In_624);
nor U100 (N_100,In_323,In_389);
xor U101 (N_101,In_451,In_941);
nor U102 (N_102,In_95,In_272);
or U103 (N_103,In_167,In_310);
or U104 (N_104,In_963,In_985);
nor U105 (N_105,In_181,In_527);
and U106 (N_106,In_564,In_629);
and U107 (N_107,In_250,In_329);
and U108 (N_108,In_321,In_805);
nor U109 (N_109,In_157,In_325);
nand U110 (N_110,In_358,In_648);
and U111 (N_111,In_748,In_702);
nor U112 (N_112,In_887,In_34);
and U113 (N_113,In_930,In_798);
nor U114 (N_114,In_354,In_422);
or U115 (N_115,In_313,In_718);
and U116 (N_116,In_543,In_888);
and U117 (N_117,In_81,In_133);
nor U118 (N_118,In_812,In_544);
and U119 (N_119,In_842,In_341);
and U120 (N_120,In_802,In_811);
and U121 (N_121,In_891,In_851);
nand U122 (N_122,In_778,In_192);
and U123 (N_123,In_195,In_189);
nor U124 (N_124,In_505,In_632);
nor U125 (N_125,In_263,In_692);
or U126 (N_126,In_198,In_788);
nor U127 (N_127,In_924,In_537);
and U128 (N_128,In_434,In_660);
nand U129 (N_129,In_384,In_758);
xor U130 (N_130,In_524,In_256);
and U131 (N_131,In_283,In_973);
nand U132 (N_132,In_834,In_722);
and U133 (N_133,In_680,In_130);
nor U134 (N_134,In_196,In_947);
nand U135 (N_135,In_258,In_55);
nor U136 (N_136,In_208,In_346);
nor U137 (N_137,In_954,In_266);
nand U138 (N_138,In_619,In_123);
nor U139 (N_139,In_918,In_445);
nor U140 (N_140,In_523,In_885);
nand U141 (N_141,In_40,In_821);
or U142 (N_142,In_685,In_525);
and U143 (N_143,In_113,In_946);
nor U144 (N_144,In_436,In_106);
nand U145 (N_145,In_330,In_10);
nand U146 (N_146,In_367,In_74);
nand U147 (N_147,In_347,In_627);
or U148 (N_148,In_177,In_831);
or U149 (N_149,In_781,In_980);
or U150 (N_150,In_534,In_213);
nand U151 (N_151,In_603,In_53);
xnor U152 (N_152,In_934,In_184);
nor U153 (N_153,In_504,In_697);
and U154 (N_154,In_832,In_642);
nor U155 (N_155,In_623,In_406);
or U156 (N_156,In_791,In_806);
xnor U157 (N_157,In_862,In_567);
or U158 (N_158,In_489,In_787);
nor U159 (N_159,In_449,In_290);
or U160 (N_160,In_413,In_704);
nor U161 (N_161,In_983,In_542);
or U162 (N_162,In_476,In_665);
and U163 (N_163,In_679,In_641);
and U164 (N_164,In_503,In_404);
nor U165 (N_165,In_378,In_931);
nor U166 (N_166,In_23,In_405);
nand U167 (N_167,In_516,In_369);
nand U168 (N_168,In_695,In_342);
or U169 (N_169,In_15,In_937);
and U170 (N_170,In_161,In_917);
and U171 (N_171,In_14,In_264);
nand U172 (N_172,In_554,In_82);
or U173 (N_173,In_608,In_589);
nor U174 (N_174,In_548,In_943);
nand U175 (N_175,In_610,In_254);
or U176 (N_176,In_48,In_149);
nand U177 (N_177,In_803,In_807);
or U178 (N_178,In_804,In_621);
or U179 (N_179,In_232,In_425);
nand U180 (N_180,In_817,In_920);
nor U181 (N_181,In_120,In_225);
or U182 (N_182,In_529,In_860);
and U183 (N_183,In_156,In_285);
nor U184 (N_184,In_228,In_5);
nand U185 (N_185,In_427,In_925);
nand U186 (N_186,In_515,In_951);
nor U187 (N_187,In_655,In_550);
or U188 (N_188,In_900,In_764);
xor U189 (N_189,In_964,In_763);
nor U190 (N_190,In_9,In_818);
nand U191 (N_191,In_898,In_179);
nor U192 (N_192,In_957,In_446);
nand U193 (N_193,In_85,In_127);
or U194 (N_194,In_876,In_978);
or U195 (N_195,In_926,In_312);
nand U196 (N_196,In_150,In_297);
and U197 (N_197,In_746,In_908);
nand U198 (N_198,In_31,In_792);
or U199 (N_199,In_607,In_109);
and U200 (N_200,In_604,In_78);
nand U201 (N_201,In_517,In_273);
nand U202 (N_202,In_852,In_488);
nor U203 (N_203,In_676,In_903);
nand U204 (N_204,In_234,In_675);
nand U205 (N_205,In_139,In_337);
nor U206 (N_206,In_497,In_97);
nor U207 (N_207,In_287,In_777);
or U208 (N_208,In_693,In_372);
nor U209 (N_209,In_653,In_956);
nor U210 (N_210,In_248,In_633);
and U211 (N_211,In_243,In_597);
nand U212 (N_212,In_845,In_56);
nor U213 (N_213,In_219,In_465);
nor U214 (N_214,In_439,In_574);
or U215 (N_215,In_148,In_238);
or U216 (N_216,In_601,In_393);
nand U217 (N_217,In_265,In_30);
and U218 (N_218,In_217,In_936);
nor U219 (N_219,In_955,In_870);
and U220 (N_220,In_461,In_839);
and U221 (N_221,In_340,In_582);
and U222 (N_222,In_979,In_147);
and U223 (N_223,In_547,In_430);
nor U224 (N_224,In_905,In_799);
nand U225 (N_225,In_249,In_766);
or U226 (N_226,In_375,In_13);
or U227 (N_227,In_511,In_443);
nand U228 (N_228,In_828,In_528);
or U229 (N_229,In_51,In_720);
nand U230 (N_230,In_809,In_304);
or U231 (N_231,In_793,In_681);
nand U232 (N_232,In_867,In_899);
and U233 (N_233,In_494,In_591);
nor U234 (N_234,In_92,In_779);
or U235 (N_235,In_901,In_578);
nand U236 (N_236,In_407,In_237);
nor U237 (N_237,In_119,In_353);
nor U238 (N_238,In_159,In_60);
and U239 (N_239,In_999,In_448);
nand U240 (N_240,In_514,In_723);
or U241 (N_241,In_42,In_419);
xnor U242 (N_242,In_893,In_907);
or U243 (N_243,In_438,In_709);
nor U244 (N_244,In_640,In_412);
nor U245 (N_245,In_73,In_160);
and U246 (N_246,In_774,In_251);
or U247 (N_247,In_348,In_622);
or U248 (N_248,In_630,In_753);
nor U249 (N_249,In_486,In_535);
nand U250 (N_250,In_395,In_493);
nor U251 (N_251,In_919,In_462);
nand U252 (N_252,In_987,In_522);
or U253 (N_253,In_993,In_736);
nand U254 (N_254,In_536,In_57);
and U255 (N_255,In_970,In_563);
or U256 (N_256,In_485,In_560);
nand U257 (N_257,In_906,In_558);
and U258 (N_258,In_960,In_260);
nand U259 (N_259,In_747,In_236);
nand U260 (N_260,In_780,In_539);
nand U261 (N_261,In_327,In_829);
and U262 (N_262,In_207,In_271);
nand U263 (N_263,In_91,In_99);
or U264 (N_264,In_569,In_111);
and U265 (N_265,In_230,In_351);
or U266 (N_266,In_84,In_201);
and U267 (N_267,In_221,In_83);
nor U268 (N_268,In_775,In_117);
and U269 (N_269,In_750,In_863);
and U270 (N_270,In_444,In_252);
nor U271 (N_271,In_125,In_545);
or U272 (N_272,In_220,In_942);
nor U273 (N_273,In_713,In_938);
and U274 (N_274,In_482,In_253);
and U275 (N_275,In_773,In_751);
nand U276 (N_276,In_733,In_39);
and U277 (N_277,In_617,In_226);
and U278 (N_278,In_914,In_822);
or U279 (N_279,In_305,In_506);
and U280 (N_280,In_17,In_566);
and U281 (N_281,In_374,In_927);
nand U282 (N_282,In_240,In_813);
nor U283 (N_283,In_45,In_789);
nor U284 (N_284,In_118,In_944);
and U285 (N_285,In_996,In_326);
or U286 (N_286,In_114,In_381);
or U287 (N_287,In_28,In_815);
and U288 (N_288,In_966,In_365);
or U289 (N_289,In_246,In_187);
and U290 (N_290,In_371,In_32);
nand U291 (N_291,In_336,In_837);
nand U292 (N_292,In_460,In_616);
or U293 (N_293,In_450,In_950);
and U294 (N_294,In_879,In_47);
or U295 (N_295,In_134,In_344);
nor U296 (N_296,In_721,In_769);
nor U297 (N_297,In_214,In_816);
nor U298 (N_298,In_269,In_502);
and U299 (N_299,In_479,In_682);
nand U300 (N_300,In_810,In_428);
and U301 (N_301,In_878,In_88);
xor U302 (N_302,In_11,In_581);
xnor U303 (N_303,In_652,In_771);
or U304 (N_304,In_701,In_480);
nor U305 (N_305,In_398,In_311);
nor U306 (N_306,In_708,In_847);
and U307 (N_307,In_170,In_513);
nand U308 (N_308,In_270,In_631);
or U309 (N_309,In_352,In_647);
or U310 (N_310,In_532,In_173);
nor U311 (N_311,In_19,In_100);
nand U312 (N_312,In_259,In_307);
xnor U313 (N_313,In_359,In_526);
and U314 (N_314,In_540,In_759);
nand U315 (N_315,In_671,In_275);
nor U316 (N_316,In_152,In_98);
or U317 (N_317,In_743,In_49);
nor U318 (N_318,In_433,In_296);
or U319 (N_319,In_848,In_666);
xnor U320 (N_320,In_820,In_364);
nand U321 (N_321,In_379,In_478);
nand U322 (N_322,In_974,In_674);
and U323 (N_323,In_231,In_64);
nor U324 (N_324,In_853,In_730);
or U325 (N_325,In_361,In_247);
and U326 (N_326,In_541,In_44);
nand U327 (N_327,In_896,In_441);
nand U328 (N_328,In_245,In_222);
or U329 (N_329,In_981,In_855);
nand U330 (N_330,In_137,In_135);
and U331 (N_331,In_501,In_509);
nor U332 (N_332,In_334,In_657);
or U333 (N_333,In_194,In_770);
and U334 (N_334,In_218,In_995);
nor U335 (N_335,In_328,In_215);
or U336 (N_336,In_391,In_800);
and U337 (N_337,In_583,In_300);
and U338 (N_338,In_592,In_20);
xnor U339 (N_339,In_89,In_577);
nand U340 (N_340,In_459,In_206);
nand U341 (N_341,In_129,In_274);
nand U342 (N_342,In_962,In_205);
nand U343 (N_343,In_734,In_932);
or U344 (N_344,In_492,In_808);
and U345 (N_345,In_634,In_605);
xnor U346 (N_346,In_897,In_115);
and U347 (N_347,In_638,In_429);
and U348 (N_348,In_877,In_142);
and U349 (N_349,In_26,In_191);
or U350 (N_350,In_411,In_112);
and U351 (N_351,In_169,In_93);
nor U352 (N_352,In_650,In_699);
xor U353 (N_353,In_594,In_71);
and U354 (N_354,In_719,In_678);
nand U355 (N_355,In_318,In_262);
nor U356 (N_356,In_96,In_355);
or U357 (N_357,In_575,In_982);
nand U358 (N_358,In_711,In_202);
nor U359 (N_359,In_185,In_830);
and U360 (N_360,In_27,In_625);
and U361 (N_361,In_952,In_366);
and U362 (N_362,In_288,In_620);
nor U363 (N_363,In_349,In_386);
and U364 (N_364,In_242,In_223);
or U365 (N_365,In_654,In_166);
nor U366 (N_366,In_2,In_178);
and U367 (N_367,In_257,In_784);
nand U368 (N_368,In_997,In_500);
nand U369 (N_369,In_1,In_16);
nor U370 (N_370,In_700,In_742);
and U371 (N_371,In_175,In_38);
nor U372 (N_372,In_740,In_79);
and U373 (N_373,In_689,In_122);
and U374 (N_374,In_886,In_690);
nor U375 (N_375,In_128,In_121);
or U376 (N_376,In_484,In_350);
xnor U377 (N_377,In_469,In_399);
nor U378 (N_378,In_843,In_556);
and U379 (N_379,In_546,In_58);
nand U380 (N_380,In_25,In_464);
xor U381 (N_381,In_174,In_383);
or U382 (N_382,In_454,In_977);
or U383 (N_383,In_724,In_136);
or U384 (N_384,In_463,In_144);
and U385 (N_385,In_153,In_424);
and U386 (N_386,In_835,In_470);
and U387 (N_387,In_182,In_0);
and U388 (N_388,In_729,In_686);
or U389 (N_389,In_276,In_338);
nor U390 (N_390,In_46,In_551);
and U391 (N_391,In_875,In_555);
and U392 (N_392,In_4,In_298);
or U393 (N_393,In_715,In_186);
or U394 (N_394,In_580,In_110);
or U395 (N_395,In_7,In_507);
or U396 (N_396,In_609,In_744);
nor U397 (N_397,In_992,In_61);
nand U398 (N_398,In_317,In_975);
and U399 (N_399,In_373,In_935);
nand U400 (N_400,In_94,In_299);
nor U401 (N_401,In_210,In_306);
nand U402 (N_402,In_512,In_90);
xnor U403 (N_403,In_490,In_661);
and U404 (N_404,In_108,In_521);
nor U405 (N_405,In_612,In_116);
and U406 (N_406,In_41,In_663);
or U407 (N_407,In_958,In_644);
xnor U408 (N_408,In_949,In_639);
nand U409 (N_409,In_836,In_431);
nand U410 (N_410,In_519,In_698);
or U411 (N_411,In_183,In_645);
and U412 (N_412,In_658,In_670);
nor U413 (N_413,In_491,In_6);
or U414 (N_414,In_971,In_755);
nor U415 (N_415,In_646,In_823);
or U416 (N_416,In_335,In_87);
nor U417 (N_417,In_772,In_437);
and U418 (N_418,In_705,In_826);
or U419 (N_419,In_107,In_360);
nor U420 (N_420,In_669,In_155);
and U421 (N_421,In_370,In_164);
nor U422 (N_422,In_131,In_596);
nor U423 (N_423,In_86,In_849);
or U424 (N_424,In_871,In_892);
nand U425 (N_425,In_691,In_472);
nor U426 (N_426,In_385,In_261);
nand U427 (N_427,In_824,In_387);
and U428 (N_428,In_255,In_396);
or U429 (N_429,In_573,In_986);
nor U430 (N_430,In_199,In_530);
nand U431 (N_431,In_880,In_282);
nor U432 (N_432,In_626,In_869);
nand U433 (N_433,In_36,In_126);
or U434 (N_434,In_881,In_320);
xor U435 (N_435,In_602,In_953);
nor U436 (N_436,In_292,In_866);
nand U437 (N_437,In_498,In_376);
nor U438 (N_438,In_677,In_163);
nor U439 (N_439,In_557,In_590);
or U440 (N_440,In_418,In_559);
or U441 (N_441,In_200,In_8);
nor U442 (N_442,In_281,In_915);
nand U443 (N_443,In_972,In_760);
and U444 (N_444,In_162,In_401);
nor U445 (N_445,In_945,In_388);
or U446 (N_446,In_928,In_611);
and U447 (N_447,In_794,In_212);
xnor U448 (N_448,In_456,In_316);
nand U449 (N_449,In_229,In_922);
and U450 (N_450,In_737,In_717);
nor U451 (N_451,In_29,In_421);
xnor U452 (N_452,In_727,In_568);
and U453 (N_453,In_302,In_394);
nand U454 (N_454,In_66,In_579);
and U455 (N_455,In_197,In_988);
and U456 (N_456,In_203,In_510);
nor U457 (N_457,In_814,In_284);
and U458 (N_458,In_562,In_859);
and U459 (N_459,In_466,In_224);
nor U460 (N_460,In_968,In_77);
and U461 (N_461,In_989,In_377);
and U462 (N_462,In_35,In_984);
nand U463 (N_463,In_618,In_235);
nor U464 (N_464,In_933,In_707);
nand U465 (N_465,In_467,In_687);
and U466 (N_466,In_549,In_69);
and U467 (N_467,In_333,In_280);
or U468 (N_468,In_473,In_452);
nand U469 (N_469,In_143,In_3);
nor U470 (N_470,In_277,In_18);
nor U471 (N_471,In_776,In_998);
nor U472 (N_472,In_362,In_572);
or U473 (N_473,In_140,In_447);
nand U474 (N_474,In_227,In_103);
nor U475 (N_475,In_76,In_703);
and U476 (N_476,In_499,In_844);
or U477 (N_477,In_598,In_739);
nor U478 (N_478,In_749,In_420);
nor U479 (N_479,In_912,In_518);
nor U480 (N_480,In_991,In_757);
nor U481 (N_481,In_768,In_165);
nand U482 (N_482,In_319,In_902);
xnor U483 (N_483,In_440,In_268);
nand U484 (N_484,In_471,In_204);
nor U485 (N_485,In_538,In_63);
or U486 (N_486,In_756,In_101);
or U487 (N_487,In_62,In_295);
or U488 (N_488,In_423,In_841);
or U489 (N_489,In_716,In_782);
and U490 (N_490,In_180,In_961);
nor U491 (N_491,In_239,In_728);
nand U492 (N_492,In_795,In_976);
nand U493 (N_493,In_12,In_22);
nor U494 (N_494,In_475,In_400);
nor U495 (N_495,In_65,In_889);
nand U496 (N_496,In_854,In_24);
and U497 (N_497,In_520,In_667);
or U498 (N_498,In_910,In_294);
nand U499 (N_499,In_417,In_833);
or U500 (N_500,In_987,In_555);
nand U501 (N_501,In_926,In_218);
nor U502 (N_502,In_614,In_609);
or U503 (N_503,In_552,In_982);
nor U504 (N_504,In_350,In_365);
nand U505 (N_505,In_229,In_680);
nand U506 (N_506,In_472,In_193);
nor U507 (N_507,In_220,In_508);
or U508 (N_508,In_924,In_172);
and U509 (N_509,In_886,In_211);
nor U510 (N_510,In_179,In_251);
nand U511 (N_511,In_744,In_549);
and U512 (N_512,In_463,In_828);
nor U513 (N_513,In_730,In_444);
nor U514 (N_514,In_816,In_564);
nor U515 (N_515,In_165,In_513);
nor U516 (N_516,In_855,In_921);
nand U517 (N_517,In_2,In_966);
nor U518 (N_518,In_738,In_119);
and U519 (N_519,In_950,In_84);
nand U520 (N_520,In_866,In_741);
or U521 (N_521,In_208,In_204);
nand U522 (N_522,In_128,In_450);
and U523 (N_523,In_119,In_724);
and U524 (N_524,In_357,In_954);
nor U525 (N_525,In_65,In_955);
nand U526 (N_526,In_499,In_23);
nand U527 (N_527,In_642,In_646);
nand U528 (N_528,In_75,In_998);
nor U529 (N_529,In_944,In_279);
nor U530 (N_530,In_908,In_340);
or U531 (N_531,In_693,In_832);
nand U532 (N_532,In_830,In_975);
and U533 (N_533,In_57,In_252);
and U534 (N_534,In_265,In_650);
nor U535 (N_535,In_301,In_547);
and U536 (N_536,In_823,In_732);
or U537 (N_537,In_242,In_870);
nor U538 (N_538,In_247,In_256);
nand U539 (N_539,In_935,In_545);
or U540 (N_540,In_950,In_54);
nor U541 (N_541,In_163,In_331);
and U542 (N_542,In_599,In_31);
nand U543 (N_543,In_943,In_78);
nand U544 (N_544,In_243,In_648);
or U545 (N_545,In_746,In_410);
or U546 (N_546,In_322,In_369);
or U547 (N_547,In_432,In_594);
or U548 (N_548,In_668,In_16);
or U549 (N_549,In_344,In_576);
nand U550 (N_550,In_9,In_707);
nor U551 (N_551,In_793,In_555);
and U552 (N_552,In_396,In_870);
nor U553 (N_553,In_5,In_528);
and U554 (N_554,In_923,In_884);
and U555 (N_555,In_921,In_40);
nand U556 (N_556,In_988,In_257);
nor U557 (N_557,In_778,In_544);
and U558 (N_558,In_280,In_95);
nor U559 (N_559,In_417,In_595);
and U560 (N_560,In_781,In_570);
nor U561 (N_561,In_580,In_985);
nor U562 (N_562,In_925,In_461);
nor U563 (N_563,In_342,In_541);
or U564 (N_564,In_929,In_13);
or U565 (N_565,In_68,In_690);
nor U566 (N_566,In_370,In_472);
nand U567 (N_567,In_871,In_400);
and U568 (N_568,In_210,In_877);
xor U569 (N_569,In_925,In_308);
and U570 (N_570,In_197,In_169);
nor U571 (N_571,In_95,In_664);
nand U572 (N_572,In_698,In_847);
nand U573 (N_573,In_708,In_545);
nor U574 (N_574,In_261,In_920);
and U575 (N_575,In_506,In_26);
or U576 (N_576,In_298,In_338);
nand U577 (N_577,In_950,In_851);
nor U578 (N_578,In_384,In_117);
nand U579 (N_579,In_68,In_970);
nand U580 (N_580,In_193,In_323);
nor U581 (N_581,In_860,In_66);
or U582 (N_582,In_702,In_453);
or U583 (N_583,In_293,In_959);
and U584 (N_584,In_946,In_273);
or U585 (N_585,In_648,In_154);
nand U586 (N_586,In_40,In_477);
nor U587 (N_587,In_359,In_985);
and U588 (N_588,In_512,In_770);
or U589 (N_589,In_880,In_233);
nand U590 (N_590,In_725,In_90);
and U591 (N_591,In_603,In_472);
nand U592 (N_592,In_882,In_793);
or U593 (N_593,In_884,In_358);
nand U594 (N_594,In_86,In_347);
or U595 (N_595,In_435,In_747);
nor U596 (N_596,In_942,In_292);
or U597 (N_597,In_808,In_220);
or U598 (N_598,In_932,In_233);
nand U599 (N_599,In_955,In_702);
or U600 (N_600,In_564,In_482);
xor U601 (N_601,In_361,In_458);
xor U602 (N_602,In_367,In_935);
or U603 (N_603,In_345,In_17);
and U604 (N_604,In_33,In_266);
and U605 (N_605,In_615,In_151);
nor U606 (N_606,In_187,In_984);
or U607 (N_607,In_805,In_658);
and U608 (N_608,In_553,In_804);
or U609 (N_609,In_449,In_726);
nand U610 (N_610,In_215,In_397);
or U611 (N_611,In_185,In_611);
or U612 (N_612,In_859,In_58);
or U613 (N_613,In_198,In_155);
xor U614 (N_614,In_989,In_511);
nor U615 (N_615,In_485,In_904);
nand U616 (N_616,In_153,In_126);
or U617 (N_617,In_244,In_692);
or U618 (N_618,In_3,In_379);
xor U619 (N_619,In_793,In_786);
nor U620 (N_620,In_208,In_579);
or U621 (N_621,In_23,In_223);
nor U622 (N_622,In_382,In_16);
and U623 (N_623,In_402,In_189);
or U624 (N_624,In_439,In_698);
xnor U625 (N_625,In_369,In_367);
or U626 (N_626,In_730,In_937);
or U627 (N_627,In_71,In_222);
and U628 (N_628,In_417,In_557);
or U629 (N_629,In_790,In_470);
nor U630 (N_630,In_430,In_42);
and U631 (N_631,In_251,In_379);
xor U632 (N_632,In_649,In_851);
nand U633 (N_633,In_365,In_993);
and U634 (N_634,In_772,In_339);
and U635 (N_635,In_630,In_807);
or U636 (N_636,In_959,In_104);
nor U637 (N_637,In_754,In_943);
or U638 (N_638,In_477,In_593);
or U639 (N_639,In_355,In_272);
or U640 (N_640,In_193,In_110);
and U641 (N_641,In_462,In_302);
or U642 (N_642,In_572,In_821);
or U643 (N_643,In_349,In_522);
nand U644 (N_644,In_972,In_532);
nand U645 (N_645,In_272,In_433);
nand U646 (N_646,In_304,In_458);
and U647 (N_647,In_937,In_211);
or U648 (N_648,In_593,In_754);
nor U649 (N_649,In_91,In_900);
nand U650 (N_650,In_125,In_362);
and U651 (N_651,In_639,In_901);
nor U652 (N_652,In_150,In_918);
or U653 (N_653,In_882,In_407);
or U654 (N_654,In_338,In_47);
and U655 (N_655,In_924,In_134);
nor U656 (N_656,In_334,In_977);
and U657 (N_657,In_926,In_593);
nand U658 (N_658,In_44,In_84);
and U659 (N_659,In_408,In_566);
nor U660 (N_660,In_584,In_898);
and U661 (N_661,In_517,In_433);
nor U662 (N_662,In_553,In_690);
nor U663 (N_663,In_742,In_947);
or U664 (N_664,In_598,In_796);
or U665 (N_665,In_764,In_787);
nor U666 (N_666,In_250,In_593);
nand U667 (N_667,In_339,In_761);
and U668 (N_668,In_796,In_942);
nand U669 (N_669,In_126,In_773);
xor U670 (N_670,In_768,In_60);
nor U671 (N_671,In_211,In_981);
nor U672 (N_672,In_459,In_857);
and U673 (N_673,In_825,In_668);
or U674 (N_674,In_766,In_52);
or U675 (N_675,In_3,In_720);
nor U676 (N_676,In_904,In_240);
nor U677 (N_677,In_612,In_8);
and U678 (N_678,In_369,In_121);
and U679 (N_679,In_731,In_952);
nand U680 (N_680,In_446,In_94);
or U681 (N_681,In_248,In_366);
nor U682 (N_682,In_982,In_758);
nand U683 (N_683,In_285,In_891);
or U684 (N_684,In_384,In_500);
nor U685 (N_685,In_751,In_209);
or U686 (N_686,In_927,In_142);
or U687 (N_687,In_456,In_444);
nor U688 (N_688,In_457,In_310);
or U689 (N_689,In_420,In_611);
nor U690 (N_690,In_80,In_240);
nand U691 (N_691,In_577,In_835);
and U692 (N_692,In_972,In_625);
nand U693 (N_693,In_687,In_952);
and U694 (N_694,In_426,In_47);
nand U695 (N_695,In_968,In_636);
or U696 (N_696,In_585,In_109);
or U697 (N_697,In_63,In_194);
nand U698 (N_698,In_528,In_638);
nand U699 (N_699,In_500,In_494);
xnor U700 (N_700,In_289,In_422);
and U701 (N_701,In_43,In_837);
nor U702 (N_702,In_154,In_657);
nor U703 (N_703,In_811,In_961);
and U704 (N_704,In_338,In_57);
nand U705 (N_705,In_459,In_175);
nand U706 (N_706,In_816,In_457);
nand U707 (N_707,In_218,In_836);
and U708 (N_708,In_857,In_639);
nand U709 (N_709,In_167,In_553);
or U710 (N_710,In_669,In_538);
and U711 (N_711,In_775,In_917);
nor U712 (N_712,In_252,In_565);
or U713 (N_713,In_967,In_383);
or U714 (N_714,In_341,In_906);
nor U715 (N_715,In_833,In_802);
nand U716 (N_716,In_990,In_649);
nand U717 (N_717,In_973,In_450);
nor U718 (N_718,In_293,In_351);
nor U719 (N_719,In_706,In_35);
or U720 (N_720,In_506,In_798);
or U721 (N_721,In_918,In_446);
nand U722 (N_722,In_195,In_936);
and U723 (N_723,In_921,In_974);
nor U724 (N_724,In_369,In_613);
xnor U725 (N_725,In_546,In_227);
nand U726 (N_726,In_13,In_57);
nor U727 (N_727,In_692,In_839);
nand U728 (N_728,In_847,In_632);
and U729 (N_729,In_591,In_539);
nor U730 (N_730,In_456,In_721);
nand U731 (N_731,In_543,In_602);
or U732 (N_732,In_723,In_957);
nor U733 (N_733,In_22,In_296);
and U734 (N_734,In_130,In_576);
nand U735 (N_735,In_39,In_643);
nand U736 (N_736,In_350,In_642);
and U737 (N_737,In_341,In_857);
nand U738 (N_738,In_476,In_128);
nor U739 (N_739,In_316,In_549);
nor U740 (N_740,In_990,In_787);
nand U741 (N_741,In_514,In_985);
nand U742 (N_742,In_94,In_199);
and U743 (N_743,In_361,In_394);
nand U744 (N_744,In_535,In_39);
nor U745 (N_745,In_709,In_740);
xnor U746 (N_746,In_494,In_903);
nand U747 (N_747,In_471,In_243);
nor U748 (N_748,In_903,In_594);
nand U749 (N_749,In_606,In_771);
nand U750 (N_750,In_964,In_411);
nand U751 (N_751,In_438,In_273);
or U752 (N_752,In_96,In_292);
nand U753 (N_753,In_646,In_104);
nand U754 (N_754,In_376,In_258);
nand U755 (N_755,In_827,In_818);
nor U756 (N_756,In_140,In_341);
nand U757 (N_757,In_66,In_756);
and U758 (N_758,In_438,In_658);
nand U759 (N_759,In_496,In_612);
and U760 (N_760,In_250,In_373);
and U761 (N_761,In_827,In_730);
or U762 (N_762,In_630,In_232);
nand U763 (N_763,In_702,In_546);
or U764 (N_764,In_452,In_536);
and U765 (N_765,In_651,In_852);
nor U766 (N_766,In_717,In_943);
or U767 (N_767,In_399,In_935);
nor U768 (N_768,In_139,In_449);
nor U769 (N_769,In_312,In_592);
nand U770 (N_770,In_772,In_655);
nor U771 (N_771,In_20,In_342);
and U772 (N_772,In_385,In_280);
and U773 (N_773,In_487,In_618);
xnor U774 (N_774,In_135,In_667);
nand U775 (N_775,In_590,In_485);
or U776 (N_776,In_846,In_36);
nor U777 (N_777,In_89,In_948);
and U778 (N_778,In_413,In_599);
nor U779 (N_779,In_36,In_7);
or U780 (N_780,In_220,In_986);
nand U781 (N_781,In_665,In_418);
xnor U782 (N_782,In_451,In_10);
nor U783 (N_783,In_848,In_613);
nor U784 (N_784,In_502,In_513);
xor U785 (N_785,In_260,In_737);
nand U786 (N_786,In_178,In_968);
or U787 (N_787,In_677,In_432);
and U788 (N_788,In_820,In_422);
or U789 (N_789,In_852,In_798);
nor U790 (N_790,In_707,In_254);
or U791 (N_791,In_620,In_251);
nand U792 (N_792,In_847,In_715);
nand U793 (N_793,In_847,In_801);
or U794 (N_794,In_637,In_178);
and U795 (N_795,In_819,In_928);
nor U796 (N_796,In_989,In_983);
or U797 (N_797,In_755,In_259);
nand U798 (N_798,In_684,In_739);
nand U799 (N_799,In_624,In_742);
nand U800 (N_800,In_516,In_634);
or U801 (N_801,In_599,In_40);
nand U802 (N_802,In_207,In_764);
nor U803 (N_803,In_639,In_385);
and U804 (N_804,In_73,In_622);
xnor U805 (N_805,In_460,In_952);
xor U806 (N_806,In_838,In_770);
nor U807 (N_807,In_698,In_37);
nor U808 (N_808,In_79,In_330);
nor U809 (N_809,In_449,In_378);
nand U810 (N_810,In_214,In_925);
nand U811 (N_811,In_126,In_631);
or U812 (N_812,In_137,In_200);
nor U813 (N_813,In_164,In_327);
and U814 (N_814,In_439,In_826);
or U815 (N_815,In_517,In_718);
nor U816 (N_816,In_9,In_548);
nand U817 (N_817,In_384,In_786);
nand U818 (N_818,In_738,In_250);
nand U819 (N_819,In_120,In_334);
and U820 (N_820,In_941,In_320);
or U821 (N_821,In_924,In_481);
nor U822 (N_822,In_820,In_119);
xor U823 (N_823,In_565,In_562);
nand U824 (N_824,In_366,In_652);
or U825 (N_825,In_695,In_675);
nand U826 (N_826,In_463,In_655);
nand U827 (N_827,In_12,In_664);
nand U828 (N_828,In_113,In_611);
and U829 (N_829,In_13,In_453);
or U830 (N_830,In_609,In_224);
and U831 (N_831,In_785,In_568);
or U832 (N_832,In_940,In_150);
nor U833 (N_833,In_142,In_832);
nor U834 (N_834,In_218,In_749);
nand U835 (N_835,In_895,In_63);
nand U836 (N_836,In_679,In_791);
or U837 (N_837,In_780,In_49);
and U838 (N_838,In_467,In_373);
or U839 (N_839,In_518,In_707);
nand U840 (N_840,In_678,In_186);
nor U841 (N_841,In_654,In_855);
nor U842 (N_842,In_723,In_35);
nor U843 (N_843,In_478,In_437);
and U844 (N_844,In_235,In_142);
nor U845 (N_845,In_311,In_230);
and U846 (N_846,In_304,In_363);
nand U847 (N_847,In_786,In_276);
nor U848 (N_848,In_234,In_640);
and U849 (N_849,In_446,In_522);
or U850 (N_850,In_692,In_600);
and U851 (N_851,In_505,In_72);
and U852 (N_852,In_406,In_39);
nand U853 (N_853,In_321,In_982);
and U854 (N_854,In_823,In_678);
nor U855 (N_855,In_17,In_337);
xor U856 (N_856,In_322,In_280);
nand U857 (N_857,In_537,In_162);
nand U858 (N_858,In_941,In_332);
nor U859 (N_859,In_532,In_946);
and U860 (N_860,In_678,In_353);
and U861 (N_861,In_737,In_589);
nor U862 (N_862,In_282,In_985);
and U863 (N_863,In_400,In_138);
nand U864 (N_864,In_556,In_729);
and U865 (N_865,In_528,In_355);
nand U866 (N_866,In_702,In_859);
nand U867 (N_867,In_825,In_872);
nand U868 (N_868,In_211,In_970);
nand U869 (N_869,In_783,In_245);
and U870 (N_870,In_624,In_506);
and U871 (N_871,In_303,In_155);
nor U872 (N_872,In_36,In_180);
and U873 (N_873,In_66,In_44);
and U874 (N_874,In_569,In_332);
nor U875 (N_875,In_115,In_164);
and U876 (N_876,In_550,In_541);
nand U877 (N_877,In_266,In_733);
nand U878 (N_878,In_490,In_497);
and U879 (N_879,In_28,In_107);
or U880 (N_880,In_161,In_335);
nand U881 (N_881,In_610,In_746);
nand U882 (N_882,In_41,In_888);
or U883 (N_883,In_214,In_576);
or U884 (N_884,In_270,In_525);
nand U885 (N_885,In_274,In_942);
nand U886 (N_886,In_292,In_157);
nor U887 (N_887,In_752,In_823);
xnor U888 (N_888,In_408,In_234);
nand U889 (N_889,In_665,In_47);
or U890 (N_890,In_946,In_155);
or U891 (N_891,In_977,In_239);
and U892 (N_892,In_98,In_194);
nand U893 (N_893,In_421,In_772);
and U894 (N_894,In_926,In_290);
and U895 (N_895,In_454,In_205);
or U896 (N_896,In_358,In_165);
nand U897 (N_897,In_28,In_384);
and U898 (N_898,In_361,In_990);
nor U899 (N_899,In_600,In_423);
and U900 (N_900,In_591,In_618);
and U901 (N_901,In_660,In_880);
and U902 (N_902,In_743,In_882);
nand U903 (N_903,In_916,In_726);
or U904 (N_904,In_995,In_700);
xor U905 (N_905,In_226,In_795);
and U906 (N_906,In_321,In_941);
nor U907 (N_907,In_690,In_936);
or U908 (N_908,In_575,In_585);
nand U909 (N_909,In_323,In_938);
nand U910 (N_910,In_249,In_533);
nor U911 (N_911,In_791,In_339);
or U912 (N_912,In_893,In_434);
and U913 (N_913,In_474,In_587);
or U914 (N_914,In_863,In_259);
or U915 (N_915,In_99,In_402);
and U916 (N_916,In_759,In_14);
or U917 (N_917,In_602,In_812);
or U918 (N_918,In_301,In_742);
or U919 (N_919,In_785,In_612);
nand U920 (N_920,In_846,In_208);
and U921 (N_921,In_274,In_235);
or U922 (N_922,In_424,In_811);
nor U923 (N_923,In_676,In_665);
nand U924 (N_924,In_377,In_181);
nand U925 (N_925,In_189,In_464);
nand U926 (N_926,In_162,In_879);
and U927 (N_927,In_870,In_490);
nor U928 (N_928,In_395,In_624);
nand U929 (N_929,In_596,In_219);
nand U930 (N_930,In_856,In_811);
nand U931 (N_931,In_632,In_85);
and U932 (N_932,In_114,In_382);
nor U933 (N_933,In_710,In_260);
and U934 (N_934,In_603,In_588);
or U935 (N_935,In_463,In_347);
and U936 (N_936,In_975,In_269);
nand U937 (N_937,In_328,In_568);
and U938 (N_938,In_407,In_607);
nor U939 (N_939,In_13,In_490);
nand U940 (N_940,In_309,In_942);
nor U941 (N_941,In_196,In_956);
nor U942 (N_942,In_250,In_140);
and U943 (N_943,In_951,In_106);
nor U944 (N_944,In_722,In_881);
or U945 (N_945,In_302,In_819);
nor U946 (N_946,In_942,In_812);
or U947 (N_947,In_932,In_498);
or U948 (N_948,In_317,In_724);
or U949 (N_949,In_144,In_940);
and U950 (N_950,In_47,In_193);
and U951 (N_951,In_114,In_666);
nand U952 (N_952,In_602,In_418);
nor U953 (N_953,In_641,In_995);
and U954 (N_954,In_249,In_957);
nor U955 (N_955,In_340,In_959);
and U956 (N_956,In_597,In_639);
nand U957 (N_957,In_458,In_620);
and U958 (N_958,In_374,In_661);
nor U959 (N_959,In_648,In_443);
and U960 (N_960,In_711,In_720);
and U961 (N_961,In_852,In_207);
and U962 (N_962,In_750,In_92);
nor U963 (N_963,In_284,In_616);
nor U964 (N_964,In_25,In_10);
or U965 (N_965,In_467,In_405);
nor U966 (N_966,In_901,In_339);
or U967 (N_967,In_763,In_617);
xnor U968 (N_968,In_730,In_657);
nor U969 (N_969,In_697,In_766);
or U970 (N_970,In_426,In_206);
nand U971 (N_971,In_77,In_933);
and U972 (N_972,In_307,In_636);
and U973 (N_973,In_226,In_815);
nor U974 (N_974,In_882,In_256);
and U975 (N_975,In_450,In_631);
nor U976 (N_976,In_789,In_366);
and U977 (N_977,In_480,In_617);
nor U978 (N_978,In_639,In_892);
nand U979 (N_979,In_747,In_968);
nand U980 (N_980,In_730,In_432);
and U981 (N_981,In_983,In_844);
nor U982 (N_982,In_205,In_563);
or U983 (N_983,In_735,In_252);
nor U984 (N_984,In_369,In_716);
nor U985 (N_985,In_33,In_138);
nand U986 (N_986,In_180,In_196);
and U987 (N_987,In_338,In_645);
nand U988 (N_988,In_132,In_765);
nor U989 (N_989,In_371,In_293);
and U990 (N_990,In_733,In_6);
or U991 (N_991,In_474,In_289);
and U992 (N_992,In_715,In_245);
or U993 (N_993,In_123,In_672);
nand U994 (N_994,In_816,In_217);
and U995 (N_995,In_648,In_317);
nor U996 (N_996,In_984,In_706);
nor U997 (N_997,In_302,In_925);
and U998 (N_998,In_463,In_269);
and U999 (N_999,In_913,In_649);
and U1000 (N_1000,N_414,N_740);
nor U1001 (N_1001,N_201,N_364);
or U1002 (N_1002,N_62,N_61);
xnor U1003 (N_1003,N_816,N_175);
and U1004 (N_1004,N_46,N_709);
nand U1005 (N_1005,N_322,N_165);
and U1006 (N_1006,N_95,N_408);
and U1007 (N_1007,N_524,N_944);
and U1008 (N_1008,N_794,N_616);
xor U1009 (N_1009,N_673,N_749);
or U1010 (N_1010,N_739,N_42);
or U1011 (N_1011,N_539,N_589);
nand U1012 (N_1012,N_987,N_263);
or U1013 (N_1013,N_857,N_438);
or U1014 (N_1014,N_587,N_16);
and U1015 (N_1015,N_181,N_343);
nand U1016 (N_1016,N_972,N_394);
nor U1017 (N_1017,N_724,N_492);
xor U1018 (N_1018,N_427,N_534);
nand U1019 (N_1019,N_865,N_475);
and U1020 (N_1020,N_168,N_847);
or U1021 (N_1021,N_300,N_639);
and U1022 (N_1022,N_247,N_308);
nand U1023 (N_1023,N_715,N_549);
and U1024 (N_1024,N_785,N_914);
or U1025 (N_1025,N_951,N_852);
nand U1026 (N_1026,N_114,N_943);
nand U1027 (N_1027,N_69,N_289);
and U1028 (N_1028,N_927,N_957);
nand U1029 (N_1029,N_478,N_52);
and U1030 (N_1030,N_615,N_331);
and U1031 (N_1031,N_407,N_541);
nor U1032 (N_1032,N_409,N_545);
and U1033 (N_1033,N_837,N_568);
nor U1034 (N_1034,N_937,N_258);
nor U1035 (N_1035,N_31,N_783);
or U1036 (N_1036,N_89,N_295);
or U1037 (N_1037,N_814,N_88);
or U1038 (N_1038,N_251,N_646);
nand U1039 (N_1039,N_695,N_22);
and U1040 (N_1040,N_554,N_202);
xnor U1041 (N_1041,N_81,N_894);
nand U1042 (N_1042,N_84,N_306);
and U1043 (N_1043,N_150,N_471);
and U1044 (N_1044,N_864,N_517);
nand U1045 (N_1045,N_981,N_451);
nor U1046 (N_1046,N_352,N_361);
nand U1047 (N_1047,N_618,N_463);
or U1048 (N_1048,N_912,N_638);
nand U1049 (N_1049,N_321,N_756);
or U1050 (N_1050,N_930,N_571);
or U1051 (N_1051,N_397,N_782);
nand U1052 (N_1052,N_932,N_706);
nand U1053 (N_1053,N_130,N_330);
and U1054 (N_1054,N_708,N_260);
nand U1055 (N_1055,N_45,N_462);
xnor U1056 (N_1056,N_174,N_860);
or U1057 (N_1057,N_692,N_106);
nand U1058 (N_1058,N_85,N_629);
nor U1059 (N_1059,N_167,N_34);
nor U1060 (N_1060,N_422,N_928);
and U1061 (N_1061,N_867,N_40);
and U1062 (N_1062,N_74,N_226);
nand U1063 (N_1063,N_291,N_873);
nor U1064 (N_1064,N_365,N_193);
xor U1065 (N_1065,N_983,N_390);
or U1066 (N_1066,N_48,N_523);
nor U1067 (N_1067,N_311,N_498);
and U1068 (N_1068,N_854,N_214);
and U1069 (N_1069,N_86,N_841);
nand U1070 (N_1070,N_730,N_955);
nor U1071 (N_1071,N_127,N_425);
nand U1072 (N_1072,N_36,N_466);
or U1073 (N_1073,N_173,N_994);
or U1074 (N_1074,N_242,N_387);
or U1075 (N_1075,N_578,N_237);
and U1076 (N_1076,N_148,N_869);
xnor U1077 (N_1077,N_598,N_839);
or U1078 (N_1078,N_810,N_101);
nand U1079 (N_1079,N_126,N_519);
nor U1080 (N_1080,N_372,N_354);
and U1081 (N_1081,N_536,N_107);
nand U1082 (N_1082,N_603,N_817);
xor U1083 (N_1083,N_391,N_583);
nor U1084 (N_1084,N_801,N_23);
and U1085 (N_1085,N_163,N_887);
or U1086 (N_1086,N_788,N_65);
nor U1087 (N_1087,N_921,N_888);
or U1088 (N_1088,N_131,N_129);
and U1089 (N_1089,N_297,N_593);
and U1090 (N_1090,N_848,N_191);
and U1091 (N_1091,N_787,N_218);
nand U1092 (N_1092,N_49,N_188);
or U1093 (N_1093,N_828,N_641);
nor U1094 (N_1094,N_123,N_373);
nand U1095 (N_1095,N_736,N_866);
and U1096 (N_1096,N_171,N_940);
or U1097 (N_1097,N_90,N_870);
nor U1098 (N_1098,N_102,N_820);
nor U1099 (N_1099,N_184,N_845);
or U1100 (N_1100,N_136,N_179);
nand U1101 (N_1101,N_923,N_43);
or U1102 (N_1102,N_273,N_780);
or U1103 (N_1103,N_378,N_241);
nand U1104 (N_1104,N_895,N_604);
nor U1105 (N_1105,N_590,N_39);
nand U1106 (N_1106,N_973,N_721);
nor U1107 (N_1107,N_185,N_815);
nor U1108 (N_1108,N_161,N_8);
nor U1109 (N_1109,N_356,N_797);
and U1110 (N_1110,N_720,N_454);
nand U1111 (N_1111,N_959,N_26);
nand U1112 (N_1112,N_314,N_876);
xor U1113 (N_1113,N_430,N_982);
or U1114 (N_1114,N_936,N_978);
or U1115 (N_1115,N_694,N_747);
nor U1116 (N_1116,N_11,N_200);
nor U1117 (N_1117,N_490,N_770);
or U1118 (N_1118,N_384,N_3);
nor U1119 (N_1119,N_376,N_644);
and U1120 (N_1120,N_71,N_953);
nor U1121 (N_1121,N_893,N_264);
or U1122 (N_1122,N_117,N_647);
or U1123 (N_1123,N_856,N_779);
nor U1124 (N_1124,N_905,N_135);
nor U1125 (N_1125,N_298,N_19);
and U1126 (N_1126,N_212,N_180);
nor U1127 (N_1127,N_890,N_217);
or U1128 (N_1128,N_717,N_566);
or U1129 (N_1129,N_155,N_124);
nand U1130 (N_1130,N_51,N_675);
nor U1131 (N_1131,N_952,N_547);
xnor U1132 (N_1132,N_455,N_299);
and U1133 (N_1133,N_614,N_500);
xnor U1134 (N_1134,N_388,N_778);
or U1135 (N_1135,N_626,N_336);
nand U1136 (N_1136,N_702,N_871);
xor U1137 (N_1137,N_934,N_746);
nand U1138 (N_1138,N_279,N_555);
xor U1139 (N_1139,N_170,N_872);
nor U1140 (N_1140,N_685,N_77);
or U1141 (N_1141,N_553,N_514);
and U1142 (N_1142,N_623,N_444);
and U1143 (N_1143,N_111,N_911);
nor U1144 (N_1144,N_268,N_690);
nand U1145 (N_1145,N_346,N_964);
nand U1146 (N_1146,N_682,N_328);
nor U1147 (N_1147,N_296,N_883);
nor U1148 (N_1148,N_924,N_960);
nand U1149 (N_1149,N_47,N_24);
and U1150 (N_1150,N_503,N_389);
or U1151 (N_1151,N_581,N_758);
or U1152 (N_1152,N_431,N_183);
nor U1153 (N_1153,N_488,N_222);
or U1154 (N_1154,N_320,N_812);
xor U1155 (N_1155,N_467,N_293);
or U1156 (N_1156,N_881,N_683);
or U1157 (N_1157,N_235,N_274);
nand U1158 (N_1158,N_433,N_803);
nand U1159 (N_1159,N_836,N_252);
nor U1160 (N_1160,N_548,N_544);
nand U1161 (N_1161,N_935,N_406);
or U1162 (N_1162,N_283,N_120);
nand U1163 (N_1163,N_383,N_696);
and U1164 (N_1164,N_502,N_680);
nand U1165 (N_1165,N_115,N_521);
or U1166 (N_1166,N_842,N_961);
and U1167 (N_1167,N_699,N_14);
nor U1168 (N_1168,N_759,N_197);
nand U1169 (N_1169,N_974,N_97);
nor U1170 (N_1170,N_177,N_760);
nand U1171 (N_1171,N_585,N_979);
or U1172 (N_1172,N_13,N_775);
and U1173 (N_1173,N_574,N_642);
and U1174 (N_1174,N_906,N_162);
and U1175 (N_1175,N_899,N_832);
or U1176 (N_1176,N_653,N_248);
nand U1177 (N_1177,N_59,N_510);
and U1178 (N_1178,N_851,N_528);
xnor U1179 (N_1179,N_579,N_711);
nor U1180 (N_1180,N_662,N_942);
or U1181 (N_1181,N_231,N_302);
nor U1182 (N_1182,N_651,N_530);
nor U1183 (N_1183,N_681,N_316);
nor U1184 (N_1184,N_993,N_344);
nor U1185 (N_1185,N_32,N_450);
or U1186 (N_1186,N_325,N_508);
nor U1187 (N_1187,N_791,N_259);
or U1188 (N_1188,N_573,N_221);
and U1189 (N_1189,N_435,N_904);
nor U1190 (N_1190,N_68,N_358);
nand U1191 (N_1191,N_975,N_417);
or U1192 (N_1192,N_381,N_307);
nor U1193 (N_1193,N_194,N_215);
nor U1194 (N_1194,N_948,N_434);
nor U1195 (N_1195,N_80,N_831);
nand U1196 (N_1196,N_35,N_954);
or U1197 (N_1197,N_947,N_657);
nand U1198 (N_1198,N_652,N_668);
nand U1199 (N_1199,N_700,N_412);
nor U1200 (N_1200,N_154,N_400);
nand U1201 (N_1201,N_613,N_456);
or U1202 (N_1202,N_984,N_827);
nand U1203 (N_1203,N_12,N_158);
or U1204 (N_1204,N_357,N_501);
and U1205 (N_1205,N_596,N_900);
nor U1206 (N_1206,N_375,N_113);
and U1207 (N_1207,N_920,N_977);
nor U1208 (N_1208,N_989,N_660);
nand U1209 (N_1209,N_239,N_569);
nor U1210 (N_1210,N_728,N_472);
nand U1211 (N_1211,N_774,N_710);
nand U1212 (N_1212,N_679,N_654);
nand U1213 (N_1213,N_511,N_476);
or U1214 (N_1214,N_572,N_725);
nand U1215 (N_1215,N_103,N_976);
and U1216 (N_1216,N_908,N_335);
nand U1217 (N_1217,N_527,N_83);
nand U1218 (N_1218,N_439,N_257);
nor U1219 (N_1219,N_495,N_773);
nand U1220 (N_1220,N_766,N_285);
xor U1221 (N_1221,N_665,N_601);
xor U1222 (N_1222,N_228,N_206);
nor U1223 (N_1223,N_727,N_386);
nor U1224 (N_1224,N_768,N_634);
nand U1225 (N_1225,N_802,N_37);
nand U1226 (N_1226,N_838,N_342);
and U1227 (N_1227,N_515,N_448);
nand U1228 (N_1228,N_104,N_341);
nor U1229 (N_1229,N_825,N_351);
and U1230 (N_1230,N_956,N_853);
nand U1231 (N_1231,N_835,N_73);
or U1232 (N_1232,N_823,N_55);
and U1233 (N_1233,N_477,N_671);
or U1234 (N_1234,N_275,N_997);
nor U1235 (N_1235,N_687,N_703);
nor U1236 (N_1236,N_677,N_885);
or U1237 (N_1237,N_499,N_305);
and U1238 (N_1238,N_238,N_965);
nor U1239 (N_1239,N_323,N_350);
and U1240 (N_1240,N_784,N_143);
nand U1241 (N_1241,N_428,N_112);
and U1242 (N_1242,N_966,N_140);
nor U1243 (N_1243,N_292,N_243);
or U1244 (N_1244,N_230,N_337);
and U1245 (N_1245,N_631,N_855);
nand U1246 (N_1246,N_506,N_368);
nor U1247 (N_1247,N_664,N_769);
nor U1248 (N_1248,N_863,N_538);
nor U1249 (N_1249,N_693,N_470);
and U1250 (N_1250,N_624,N_63);
nor U1251 (N_1251,N_850,N_421);
and U1252 (N_1252,N_922,N_907);
nand U1253 (N_1253,N_182,N_271);
nand U1254 (N_1254,N_891,N_423);
or U1255 (N_1255,N_482,N_110);
nor U1256 (N_1256,N_892,N_712);
nand U1257 (N_1257,N_594,N_99);
or U1258 (N_1258,N_269,N_220);
or U1259 (N_1259,N_21,N_209);
or U1260 (N_1260,N_575,N_277);
nand U1261 (N_1261,N_882,N_286);
nor U1262 (N_1262,N_166,N_78);
and U1263 (N_1263,N_754,N_755);
and U1264 (N_1264,N_862,N_591);
nand U1265 (N_1265,N_561,N_118);
or U1266 (N_1266,N_707,N_125);
or U1267 (N_1267,N_632,N_44);
and U1268 (N_1268,N_460,N_877);
and U1269 (N_1269,N_599,N_216);
nand U1270 (N_1270,N_98,N_985);
xnor U1271 (N_1271,N_332,N_303);
nor U1272 (N_1272,N_100,N_809);
or U1273 (N_1273,N_93,N_689);
or U1274 (N_1274,N_326,N_232);
nand U1275 (N_1275,N_748,N_520);
and U1276 (N_1276,N_645,N_830);
and U1277 (N_1277,N_586,N_790);
or U1278 (N_1278,N_868,N_805);
nand U1279 (N_1279,N_189,N_595);
or U1280 (N_1280,N_840,N_109);
nand U1281 (N_1281,N_910,N_447);
nor U1282 (N_1282,N_996,N_532);
or U1283 (N_1283,N_338,N_886);
nand U1284 (N_1284,N_419,N_236);
and U1285 (N_1285,N_245,N_600);
nor U1286 (N_1286,N_190,N_410);
nand U1287 (N_1287,N_9,N_276);
nor U1288 (N_1288,N_543,N_516);
nor U1289 (N_1289,N_990,N_436);
and U1290 (N_1290,N_884,N_192);
xor U1291 (N_1291,N_440,N_558);
nor U1292 (N_1292,N_781,N_958);
nand U1293 (N_1293,N_795,N_811);
and U1294 (N_1294,N_496,N_2);
nand U1295 (N_1295,N_211,N_280);
and U1296 (N_1296,N_819,N_382);
nand U1297 (N_1297,N_762,N_79);
or U1298 (N_1298,N_329,N_902);
nor U1299 (N_1299,N_526,N_7);
or U1300 (N_1300,N_315,N_761);
and U1301 (N_1301,N_160,N_915);
nand U1302 (N_1302,N_418,N_963);
and U1303 (N_1303,N_327,N_385);
nand U1304 (N_1304,N_648,N_546);
or U1305 (N_1305,N_663,N_735);
xor U1306 (N_1306,N_808,N_666);
or U1307 (N_1307,N_146,N_29);
nor U1308 (N_1308,N_659,N_324);
nand U1309 (N_1309,N_901,N_186);
or U1310 (N_1310,N_255,N_254);
or U1311 (N_1311,N_941,N_878);
or U1312 (N_1312,N_898,N_301);
nor U1313 (N_1313,N_287,N_729);
nor U1314 (N_1314,N_333,N_550);
nand U1315 (N_1315,N_225,N_834);
and U1316 (N_1316,N_610,N_429);
and U1317 (N_1317,N_310,N_992);
or U1318 (N_1318,N_493,N_437);
nand U1319 (N_1319,N_5,N_741);
nand U1320 (N_1320,N_38,N_334);
nand U1321 (N_1321,N_187,N_757);
nand U1322 (N_1322,N_988,N_826);
and U1323 (N_1323,N_938,N_612);
nand U1324 (N_1324,N_25,N_443);
or U1325 (N_1325,N_317,N_91);
nand U1326 (N_1326,N_620,N_92);
nor U1327 (N_1327,N_844,N_818);
nand U1328 (N_1328,N_265,N_157);
or U1329 (N_1329,N_584,N_227);
or U1330 (N_1330,N_874,N_319);
and U1331 (N_1331,N_946,N_945);
or U1332 (N_1332,N_147,N_967);
and U1333 (N_1333,N_244,N_658);
nand U1334 (N_1334,N_76,N_733);
nand U1335 (N_1335,N_1,N_531);
nor U1336 (N_1336,N_272,N_786);
or U1337 (N_1337,N_504,N_716);
or U1338 (N_1338,N_743,N_58);
and U1339 (N_1339,N_141,N_701);
nor U1340 (N_1340,N_497,N_619);
xor U1341 (N_1341,N_796,N_288);
nand U1342 (N_1342,N_176,N_402);
nand U1343 (N_1343,N_420,N_15);
nand U1344 (N_1344,N_156,N_793);
and U1345 (N_1345,N_734,N_349);
or U1346 (N_1346,N_33,N_261);
nor U1347 (N_1347,N_995,N_557);
or U1348 (N_1348,N_968,N_153);
or U1349 (N_1349,N_643,N_152);
nand U1350 (N_1350,N_731,N_142);
or U1351 (N_1351,N_672,N_843);
and U1352 (N_1352,N_369,N_522);
nand U1353 (N_1353,N_50,N_404);
nand U1354 (N_1354,N_128,N_453);
nor U1355 (N_1355,N_10,N_403);
nor U1356 (N_1356,N_213,N_925);
nor U1357 (N_1357,N_688,N_897);
or U1358 (N_1358,N_70,N_379);
nor U1359 (N_1359,N_464,N_207);
or U1360 (N_1360,N_137,N_576);
nand U1361 (N_1361,N_159,N_792);
nor U1362 (N_1362,N_813,N_340);
and U1363 (N_1363,N_611,N_875);
nor U1364 (N_1364,N_649,N_723);
and U1365 (N_1365,N_469,N_540);
and U1366 (N_1366,N_377,N_208);
and U1367 (N_1367,N_763,N_726);
nor U1368 (N_1368,N_822,N_392);
nand U1369 (N_1369,N_367,N_752);
nand U1370 (N_1370,N_732,N_18);
nand U1371 (N_1371,N_933,N_608);
nor U1372 (N_1372,N_432,N_398);
nand U1373 (N_1373,N_75,N_588);
or U1374 (N_1374,N_602,N_628);
and U1375 (N_1375,N_452,N_804);
and U1376 (N_1376,N_627,N_290);
or U1377 (N_1377,N_481,N_57);
and U1378 (N_1378,N_345,N_931);
or U1379 (N_1379,N_318,N_304);
nand U1380 (N_1380,N_718,N_577);
and U1381 (N_1381,N_371,N_309);
nor U1382 (N_1382,N_196,N_861);
nand U1383 (N_1383,N_473,N_169);
nor U1384 (N_1384,N_737,N_705);
or U1385 (N_1385,N_284,N_41);
nand U1386 (N_1386,N_744,N_393);
nand U1387 (N_1387,N_374,N_580);
or U1388 (N_1388,N_234,N_138);
and U1389 (N_1389,N_348,N_203);
nand U1390 (N_1390,N_262,N_30);
nor U1391 (N_1391,N_607,N_551);
nor U1392 (N_1392,N_635,N_363);
or U1393 (N_1393,N_445,N_401);
or U1394 (N_1394,N_353,N_480);
and U1395 (N_1395,N_789,N_800);
and U1396 (N_1396,N_424,N_474);
nand U1397 (N_1397,N_950,N_461);
nor U1398 (N_1398,N_53,N_750);
nor U1399 (N_1399,N_533,N_224);
nor U1400 (N_1400,N_560,N_916);
nor U1401 (N_1401,N_281,N_606);
nor U1402 (N_1402,N_676,N_67);
nor U1403 (N_1403,N_625,N_108);
nand U1404 (N_1404,N_777,N_542);
nor U1405 (N_1405,N_859,N_909);
or U1406 (N_1406,N_637,N_806);
nand U1407 (N_1407,N_929,N_413);
or U1408 (N_1408,N_655,N_172);
and U1409 (N_1409,N_879,N_742);
nor U1410 (N_1410,N_798,N_426);
nand U1411 (N_1411,N_807,N_278);
or U1412 (N_1412,N_347,N_537);
nor U1413 (N_1413,N_479,N_396);
nor U1414 (N_1414,N_829,N_411);
and U1415 (N_1415,N_833,N_552);
nor U1416 (N_1416,N_745,N_27);
nor U1417 (N_1417,N_582,N_266);
or U1418 (N_1418,N_567,N_205);
xor U1419 (N_1419,N_94,N_210);
nor U1420 (N_1420,N_366,N_54);
nand U1421 (N_1421,N_441,N_339);
or U1422 (N_1422,N_233,N_512);
nand U1423 (N_1423,N_661,N_458);
nand U1424 (N_1424,N_999,N_229);
or U1425 (N_1425,N_556,N_223);
nand U1426 (N_1426,N_294,N_670);
or U1427 (N_1427,N_139,N_998);
nand U1428 (N_1428,N_116,N_713);
or U1429 (N_1429,N_267,N_597);
nand U1430 (N_1430,N_684,N_518);
nor U1431 (N_1431,N_903,N_969);
or U1432 (N_1432,N_697,N_719);
and U1433 (N_1433,N_87,N_355);
and U1434 (N_1434,N_96,N_246);
nand U1435 (N_1435,N_764,N_939);
or U1436 (N_1436,N_256,N_535);
or U1437 (N_1437,N_399,N_970);
or U1438 (N_1438,N_449,N_105);
xor U1439 (N_1439,N_962,N_219);
and U1440 (N_1440,N_119,N_282);
and U1441 (N_1441,N_270,N_56);
nand U1442 (N_1442,N_28,N_483);
nor U1443 (N_1443,N_765,N_751);
nor U1444 (N_1444,N_195,N_505);
nand U1445 (N_1445,N_134,N_66);
and U1446 (N_1446,N_370,N_980);
or U1447 (N_1447,N_380,N_564);
or U1448 (N_1448,N_359,N_132);
nand U1449 (N_1449,N_714,N_151);
nor U1450 (N_1450,N_489,N_565);
nor U1451 (N_1451,N_667,N_633);
xnor U1452 (N_1452,N_824,N_529);
and U1453 (N_1453,N_896,N_772);
and U1454 (N_1454,N_698,N_691);
nand U1455 (N_1455,N_674,N_617);
nor U1456 (N_1456,N_621,N_525);
nor U1457 (N_1457,N_64,N_570);
nand U1458 (N_1458,N_630,N_82);
nand U1459 (N_1459,N_313,N_17);
or U1460 (N_1460,N_416,N_917);
nand U1461 (N_1461,N_144,N_636);
nand U1462 (N_1462,N_767,N_249);
nor U1463 (N_1463,N_442,N_704);
nand U1464 (N_1464,N_821,N_4);
or U1465 (N_1465,N_889,N_60);
nand U1466 (N_1466,N_486,N_459);
or U1467 (N_1467,N_858,N_986);
nand U1468 (N_1468,N_253,N_485);
and U1469 (N_1469,N_562,N_971);
nor U1470 (N_1470,N_846,N_771);
or U1471 (N_1471,N_722,N_622);
nor U1472 (N_1472,N_6,N_656);
nor U1473 (N_1473,N_465,N_509);
nor U1474 (N_1474,N_880,N_849);
nand U1475 (N_1475,N_362,N_122);
xor U1476 (N_1476,N_563,N_360);
nor U1477 (N_1477,N_72,N_494);
nand U1478 (N_1478,N_121,N_415);
and U1479 (N_1479,N_559,N_487);
or U1480 (N_1480,N_145,N_605);
nor U1481 (N_1481,N_457,N_799);
nand U1482 (N_1482,N_468,N_949);
and U1483 (N_1483,N_513,N_491);
nand U1484 (N_1484,N_753,N_0);
or U1485 (N_1485,N_918,N_405);
or U1486 (N_1486,N_395,N_609);
nor U1487 (N_1487,N_669,N_484);
nor U1488 (N_1488,N_650,N_776);
and U1489 (N_1489,N_198,N_592);
or U1490 (N_1490,N_640,N_678);
nor U1491 (N_1491,N_164,N_913);
nand U1492 (N_1492,N_204,N_919);
and U1493 (N_1493,N_250,N_178);
nor U1494 (N_1494,N_133,N_991);
or U1495 (N_1495,N_199,N_20);
nand U1496 (N_1496,N_240,N_686);
and U1497 (N_1497,N_149,N_738);
nand U1498 (N_1498,N_507,N_926);
or U1499 (N_1499,N_446,N_312);
or U1500 (N_1500,N_247,N_598);
nor U1501 (N_1501,N_159,N_576);
and U1502 (N_1502,N_658,N_366);
nor U1503 (N_1503,N_819,N_513);
and U1504 (N_1504,N_438,N_947);
nor U1505 (N_1505,N_648,N_447);
and U1506 (N_1506,N_161,N_654);
or U1507 (N_1507,N_128,N_618);
or U1508 (N_1508,N_225,N_275);
xor U1509 (N_1509,N_115,N_877);
and U1510 (N_1510,N_724,N_336);
or U1511 (N_1511,N_852,N_517);
nand U1512 (N_1512,N_208,N_434);
xor U1513 (N_1513,N_642,N_18);
nor U1514 (N_1514,N_90,N_139);
and U1515 (N_1515,N_14,N_454);
nor U1516 (N_1516,N_852,N_960);
or U1517 (N_1517,N_606,N_891);
nor U1518 (N_1518,N_751,N_154);
or U1519 (N_1519,N_173,N_303);
or U1520 (N_1520,N_170,N_680);
nor U1521 (N_1521,N_294,N_208);
nor U1522 (N_1522,N_12,N_873);
and U1523 (N_1523,N_37,N_219);
or U1524 (N_1524,N_728,N_710);
and U1525 (N_1525,N_683,N_816);
and U1526 (N_1526,N_778,N_20);
and U1527 (N_1527,N_860,N_167);
and U1528 (N_1528,N_643,N_713);
or U1529 (N_1529,N_776,N_280);
xor U1530 (N_1530,N_992,N_289);
nand U1531 (N_1531,N_558,N_22);
nor U1532 (N_1532,N_131,N_426);
nand U1533 (N_1533,N_992,N_284);
nor U1534 (N_1534,N_210,N_928);
nor U1535 (N_1535,N_460,N_605);
nor U1536 (N_1536,N_604,N_256);
nand U1537 (N_1537,N_274,N_715);
or U1538 (N_1538,N_547,N_545);
nand U1539 (N_1539,N_991,N_329);
or U1540 (N_1540,N_854,N_200);
nor U1541 (N_1541,N_352,N_548);
nand U1542 (N_1542,N_115,N_742);
nor U1543 (N_1543,N_968,N_517);
nand U1544 (N_1544,N_267,N_458);
and U1545 (N_1545,N_213,N_724);
nor U1546 (N_1546,N_329,N_951);
nor U1547 (N_1547,N_582,N_242);
and U1548 (N_1548,N_58,N_391);
nand U1549 (N_1549,N_701,N_378);
or U1550 (N_1550,N_77,N_441);
or U1551 (N_1551,N_252,N_170);
and U1552 (N_1552,N_984,N_220);
or U1553 (N_1553,N_292,N_618);
and U1554 (N_1554,N_829,N_626);
nand U1555 (N_1555,N_588,N_128);
or U1556 (N_1556,N_71,N_501);
or U1557 (N_1557,N_212,N_808);
and U1558 (N_1558,N_62,N_581);
and U1559 (N_1559,N_360,N_712);
nand U1560 (N_1560,N_201,N_839);
nor U1561 (N_1561,N_178,N_934);
and U1562 (N_1562,N_741,N_994);
and U1563 (N_1563,N_673,N_410);
or U1564 (N_1564,N_998,N_173);
or U1565 (N_1565,N_897,N_591);
or U1566 (N_1566,N_624,N_678);
or U1567 (N_1567,N_741,N_898);
nand U1568 (N_1568,N_150,N_250);
xnor U1569 (N_1569,N_353,N_243);
or U1570 (N_1570,N_785,N_425);
and U1571 (N_1571,N_902,N_721);
nor U1572 (N_1572,N_88,N_854);
nand U1573 (N_1573,N_648,N_582);
nand U1574 (N_1574,N_494,N_32);
and U1575 (N_1575,N_809,N_414);
xor U1576 (N_1576,N_241,N_786);
nor U1577 (N_1577,N_141,N_774);
and U1578 (N_1578,N_893,N_422);
and U1579 (N_1579,N_602,N_781);
or U1580 (N_1580,N_245,N_948);
and U1581 (N_1581,N_534,N_151);
and U1582 (N_1582,N_325,N_925);
nor U1583 (N_1583,N_954,N_792);
and U1584 (N_1584,N_760,N_902);
or U1585 (N_1585,N_711,N_74);
and U1586 (N_1586,N_289,N_365);
and U1587 (N_1587,N_423,N_214);
nor U1588 (N_1588,N_166,N_896);
nand U1589 (N_1589,N_764,N_633);
nand U1590 (N_1590,N_558,N_415);
nor U1591 (N_1591,N_529,N_342);
nor U1592 (N_1592,N_372,N_429);
and U1593 (N_1593,N_842,N_791);
nor U1594 (N_1594,N_172,N_29);
or U1595 (N_1595,N_481,N_584);
nor U1596 (N_1596,N_205,N_836);
nor U1597 (N_1597,N_800,N_258);
or U1598 (N_1598,N_404,N_17);
nor U1599 (N_1599,N_233,N_796);
nand U1600 (N_1600,N_663,N_652);
and U1601 (N_1601,N_393,N_864);
nand U1602 (N_1602,N_233,N_927);
nor U1603 (N_1603,N_899,N_668);
nor U1604 (N_1604,N_712,N_151);
nor U1605 (N_1605,N_220,N_532);
and U1606 (N_1606,N_311,N_622);
nor U1607 (N_1607,N_320,N_167);
nand U1608 (N_1608,N_918,N_606);
nand U1609 (N_1609,N_55,N_234);
xor U1610 (N_1610,N_271,N_172);
nand U1611 (N_1611,N_773,N_804);
and U1612 (N_1612,N_343,N_312);
and U1613 (N_1613,N_650,N_186);
nand U1614 (N_1614,N_237,N_207);
nor U1615 (N_1615,N_735,N_873);
and U1616 (N_1616,N_190,N_908);
or U1617 (N_1617,N_972,N_385);
nor U1618 (N_1618,N_481,N_771);
or U1619 (N_1619,N_263,N_441);
and U1620 (N_1620,N_948,N_982);
or U1621 (N_1621,N_597,N_494);
and U1622 (N_1622,N_483,N_640);
or U1623 (N_1623,N_408,N_377);
nor U1624 (N_1624,N_659,N_662);
nand U1625 (N_1625,N_284,N_869);
nand U1626 (N_1626,N_287,N_192);
nand U1627 (N_1627,N_425,N_60);
or U1628 (N_1628,N_297,N_266);
or U1629 (N_1629,N_504,N_613);
nor U1630 (N_1630,N_363,N_815);
and U1631 (N_1631,N_672,N_263);
nand U1632 (N_1632,N_349,N_51);
nor U1633 (N_1633,N_689,N_468);
and U1634 (N_1634,N_989,N_595);
or U1635 (N_1635,N_389,N_74);
nand U1636 (N_1636,N_251,N_242);
nor U1637 (N_1637,N_653,N_553);
nor U1638 (N_1638,N_52,N_559);
and U1639 (N_1639,N_6,N_422);
or U1640 (N_1640,N_487,N_496);
nand U1641 (N_1641,N_279,N_688);
nor U1642 (N_1642,N_84,N_539);
nand U1643 (N_1643,N_229,N_957);
or U1644 (N_1644,N_497,N_633);
nor U1645 (N_1645,N_546,N_699);
nand U1646 (N_1646,N_461,N_368);
or U1647 (N_1647,N_66,N_174);
or U1648 (N_1648,N_772,N_546);
nand U1649 (N_1649,N_684,N_169);
nand U1650 (N_1650,N_88,N_219);
or U1651 (N_1651,N_557,N_651);
and U1652 (N_1652,N_135,N_284);
nor U1653 (N_1653,N_796,N_896);
or U1654 (N_1654,N_872,N_72);
and U1655 (N_1655,N_2,N_339);
or U1656 (N_1656,N_259,N_293);
or U1657 (N_1657,N_210,N_228);
nor U1658 (N_1658,N_590,N_682);
and U1659 (N_1659,N_529,N_692);
nor U1660 (N_1660,N_563,N_436);
nor U1661 (N_1661,N_497,N_357);
or U1662 (N_1662,N_193,N_824);
or U1663 (N_1663,N_453,N_908);
or U1664 (N_1664,N_118,N_469);
nor U1665 (N_1665,N_644,N_54);
nor U1666 (N_1666,N_250,N_402);
nand U1667 (N_1667,N_298,N_794);
and U1668 (N_1668,N_32,N_779);
nor U1669 (N_1669,N_157,N_233);
or U1670 (N_1670,N_647,N_363);
nand U1671 (N_1671,N_423,N_658);
or U1672 (N_1672,N_766,N_533);
nor U1673 (N_1673,N_375,N_689);
or U1674 (N_1674,N_664,N_72);
or U1675 (N_1675,N_560,N_448);
nor U1676 (N_1676,N_875,N_737);
and U1677 (N_1677,N_821,N_209);
or U1678 (N_1678,N_208,N_340);
nand U1679 (N_1679,N_85,N_62);
and U1680 (N_1680,N_436,N_694);
and U1681 (N_1681,N_789,N_73);
or U1682 (N_1682,N_875,N_801);
nand U1683 (N_1683,N_70,N_943);
or U1684 (N_1684,N_615,N_747);
and U1685 (N_1685,N_375,N_711);
nand U1686 (N_1686,N_333,N_858);
nand U1687 (N_1687,N_457,N_885);
nor U1688 (N_1688,N_458,N_962);
nand U1689 (N_1689,N_131,N_626);
and U1690 (N_1690,N_470,N_129);
nand U1691 (N_1691,N_546,N_885);
nor U1692 (N_1692,N_121,N_713);
xnor U1693 (N_1693,N_364,N_642);
or U1694 (N_1694,N_292,N_883);
and U1695 (N_1695,N_680,N_822);
nand U1696 (N_1696,N_615,N_325);
nor U1697 (N_1697,N_928,N_776);
and U1698 (N_1698,N_113,N_127);
nor U1699 (N_1699,N_406,N_452);
and U1700 (N_1700,N_739,N_742);
nand U1701 (N_1701,N_512,N_492);
nand U1702 (N_1702,N_310,N_420);
nand U1703 (N_1703,N_336,N_796);
or U1704 (N_1704,N_960,N_894);
and U1705 (N_1705,N_834,N_643);
nand U1706 (N_1706,N_1,N_686);
nor U1707 (N_1707,N_701,N_86);
and U1708 (N_1708,N_56,N_952);
nor U1709 (N_1709,N_286,N_728);
or U1710 (N_1710,N_785,N_736);
and U1711 (N_1711,N_92,N_50);
nand U1712 (N_1712,N_767,N_489);
and U1713 (N_1713,N_855,N_808);
or U1714 (N_1714,N_770,N_721);
or U1715 (N_1715,N_395,N_745);
or U1716 (N_1716,N_15,N_466);
and U1717 (N_1717,N_654,N_432);
nand U1718 (N_1718,N_425,N_353);
nand U1719 (N_1719,N_614,N_827);
nor U1720 (N_1720,N_628,N_618);
and U1721 (N_1721,N_226,N_862);
nor U1722 (N_1722,N_256,N_345);
or U1723 (N_1723,N_35,N_187);
and U1724 (N_1724,N_764,N_79);
nand U1725 (N_1725,N_490,N_237);
nand U1726 (N_1726,N_111,N_98);
or U1727 (N_1727,N_126,N_350);
or U1728 (N_1728,N_464,N_63);
or U1729 (N_1729,N_39,N_177);
and U1730 (N_1730,N_696,N_552);
nand U1731 (N_1731,N_165,N_771);
and U1732 (N_1732,N_123,N_246);
xor U1733 (N_1733,N_981,N_884);
or U1734 (N_1734,N_734,N_466);
nand U1735 (N_1735,N_65,N_360);
and U1736 (N_1736,N_917,N_504);
or U1737 (N_1737,N_536,N_505);
or U1738 (N_1738,N_815,N_941);
xnor U1739 (N_1739,N_833,N_791);
and U1740 (N_1740,N_375,N_908);
nand U1741 (N_1741,N_391,N_220);
and U1742 (N_1742,N_414,N_267);
and U1743 (N_1743,N_905,N_593);
and U1744 (N_1744,N_819,N_926);
and U1745 (N_1745,N_444,N_121);
or U1746 (N_1746,N_837,N_673);
nor U1747 (N_1747,N_171,N_366);
nand U1748 (N_1748,N_953,N_601);
and U1749 (N_1749,N_8,N_420);
nor U1750 (N_1750,N_502,N_18);
nand U1751 (N_1751,N_482,N_550);
nand U1752 (N_1752,N_437,N_204);
or U1753 (N_1753,N_930,N_69);
and U1754 (N_1754,N_297,N_569);
nor U1755 (N_1755,N_234,N_450);
nor U1756 (N_1756,N_912,N_457);
nand U1757 (N_1757,N_831,N_954);
or U1758 (N_1758,N_982,N_58);
and U1759 (N_1759,N_86,N_432);
nor U1760 (N_1760,N_642,N_705);
or U1761 (N_1761,N_165,N_856);
nor U1762 (N_1762,N_889,N_137);
and U1763 (N_1763,N_393,N_86);
or U1764 (N_1764,N_823,N_639);
or U1765 (N_1765,N_655,N_155);
and U1766 (N_1766,N_761,N_355);
nand U1767 (N_1767,N_961,N_128);
and U1768 (N_1768,N_639,N_873);
nor U1769 (N_1769,N_571,N_218);
or U1770 (N_1770,N_27,N_587);
and U1771 (N_1771,N_771,N_398);
and U1772 (N_1772,N_697,N_361);
and U1773 (N_1773,N_23,N_38);
nand U1774 (N_1774,N_562,N_619);
and U1775 (N_1775,N_524,N_715);
nand U1776 (N_1776,N_286,N_284);
nor U1777 (N_1777,N_615,N_224);
and U1778 (N_1778,N_25,N_38);
nor U1779 (N_1779,N_545,N_612);
nor U1780 (N_1780,N_208,N_142);
nor U1781 (N_1781,N_301,N_438);
or U1782 (N_1782,N_782,N_455);
or U1783 (N_1783,N_215,N_117);
nor U1784 (N_1784,N_263,N_24);
nand U1785 (N_1785,N_118,N_499);
nand U1786 (N_1786,N_165,N_979);
or U1787 (N_1787,N_807,N_803);
nand U1788 (N_1788,N_977,N_735);
or U1789 (N_1789,N_416,N_672);
or U1790 (N_1790,N_33,N_547);
nand U1791 (N_1791,N_241,N_994);
or U1792 (N_1792,N_712,N_980);
nor U1793 (N_1793,N_690,N_481);
or U1794 (N_1794,N_993,N_431);
nand U1795 (N_1795,N_585,N_563);
nand U1796 (N_1796,N_588,N_882);
nand U1797 (N_1797,N_115,N_72);
or U1798 (N_1798,N_962,N_863);
nor U1799 (N_1799,N_356,N_908);
and U1800 (N_1800,N_163,N_232);
nor U1801 (N_1801,N_248,N_601);
xnor U1802 (N_1802,N_391,N_135);
or U1803 (N_1803,N_286,N_912);
xor U1804 (N_1804,N_445,N_188);
nor U1805 (N_1805,N_420,N_121);
or U1806 (N_1806,N_791,N_727);
or U1807 (N_1807,N_91,N_102);
nor U1808 (N_1808,N_745,N_512);
nand U1809 (N_1809,N_257,N_708);
and U1810 (N_1810,N_202,N_281);
and U1811 (N_1811,N_827,N_892);
or U1812 (N_1812,N_353,N_177);
and U1813 (N_1813,N_738,N_315);
or U1814 (N_1814,N_118,N_477);
or U1815 (N_1815,N_9,N_888);
and U1816 (N_1816,N_305,N_662);
and U1817 (N_1817,N_919,N_754);
or U1818 (N_1818,N_325,N_969);
nor U1819 (N_1819,N_205,N_494);
or U1820 (N_1820,N_237,N_156);
or U1821 (N_1821,N_916,N_397);
or U1822 (N_1822,N_663,N_364);
nor U1823 (N_1823,N_750,N_919);
and U1824 (N_1824,N_807,N_840);
nand U1825 (N_1825,N_838,N_971);
or U1826 (N_1826,N_26,N_105);
and U1827 (N_1827,N_611,N_175);
and U1828 (N_1828,N_705,N_319);
or U1829 (N_1829,N_778,N_97);
and U1830 (N_1830,N_133,N_787);
and U1831 (N_1831,N_981,N_753);
or U1832 (N_1832,N_644,N_42);
or U1833 (N_1833,N_752,N_244);
nor U1834 (N_1834,N_675,N_238);
and U1835 (N_1835,N_611,N_131);
nand U1836 (N_1836,N_22,N_667);
nand U1837 (N_1837,N_764,N_997);
and U1838 (N_1838,N_435,N_909);
nor U1839 (N_1839,N_659,N_159);
and U1840 (N_1840,N_273,N_905);
nand U1841 (N_1841,N_46,N_417);
nand U1842 (N_1842,N_917,N_132);
or U1843 (N_1843,N_46,N_856);
nor U1844 (N_1844,N_731,N_252);
or U1845 (N_1845,N_123,N_182);
and U1846 (N_1846,N_485,N_385);
and U1847 (N_1847,N_275,N_210);
nand U1848 (N_1848,N_827,N_883);
nor U1849 (N_1849,N_122,N_325);
and U1850 (N_1850,N_300,N_955);
xnor U1851 (N_1851,N_113,N_78);
or U1852 (N_1852,N_705,N_197);
nor U1853 (N_1853,N_78,N_843);
and U1854 (N_1854,N_801,N_710);
and U1855 (N_1855,N_623,N_232);
nand U1856 (N_1856,N_807,N_962);
and U1857 (N_1857,N_352,N_972);
nand U1858 (N_1858,N_242,N_834);
and U1859 (N_1859,N_792,N_836);
or U1860 (N_1860,N_859,N_734);
nand U1861 (N_1861,N_236,N_813);
xor U1862 (N_1862,N_4,N_184);
or U1863 (N_1863,N_372,N_835);
nand U1864 (N_1864,N_105,N_116);
and U1865 (N_1865,N_279,N_432);
nor U1866 (N_1866,N_281,N_660);
nand U1867 (N_1867,N_515,N_366);
nand U1868 (N_1868,N_66,N_242);
and U1869 (N_1869,N_92,N_331);
xor U1870 (N_1870,N_366,N_962);
and U1871 (N_1871,N_496,N_578);
or U1872 (N_1872,N_788,N_529);
or U1873 (N_1873,N_624,N_450);
nor U1874 (N_1874,N_478,N_645);
nand U1875 (N_1875,N_252,N_521);
nand U1876 (N_1876,N_9,N_619);
nor U1877 (N_1877,N_466,N_327);
nor U1878 (N_1878,N_932,N_163);
and U1879 (N_1879,N_844,N_436);
nand U1880 (N_1880,N_155,N_472);
or U1881 (N_1881,N_190,N_788);
nor U1882 (N_1882,N_623,N_546);
nand U1883 (N_1883,N_989,N_30);
nor U1884 (N_1884,N_904,N_320);
or U1885 (N_1885,N_561,N_479);
nor U1886 (N_1886,N_918,N_344);
or U1887 (N_1887,N_560,N_143);
and U1888 (N_1888,N_243,N_427);
or U1889 (N_1889,N_339,N_646);
nor U1890 (N_1890,N_904,N_905);
nor U1891 (N_1891,N_1,N_974);
nor U1892 (N_1892,N_935,N_268);
xnor U1893 (N_1893,N_96,N_380);
nor U1894 (N_1894,N_745,N_344);
nand U1895 (N_1895,N_79,N_439);
nand U1896 (N_1896,N_299,N_647);
nor U1897 (N_1897,N_783,N_80);
nand U1898 (N_1898,N_979,N_773);
nand U1899 (N_1899,N_154,N_537);
or U1900 (N_1900,N_434,N_449);
or U1901 (N_1901,N_214,N_391);
nor U1902 (N_1902,N_944,N_933);
nor U1903 (N_1903,N_929,N_986);
nand U1904 (N_1904,N_163,N_869);
nand U1905 (N_1905,N_631,N_593);
nand U1906 (N_1906,N_358,N_328);
nand U1907 (N_1907,N_631,N_747);
nand U1908 (N_1908,N_547,N_482);
nor U1909 (N_1909,N_320,N_332);
and U1910 (N_1910,N_289,N_444);
and U1911 (N_1911,N_266,N_389);
and U1912 (N_1912,N_210,N_797);
or U1913 (N_1913,N_406,N_629);
or U1914 (N_1914,N_308,N_266);
or U1915 (N_1915,N_301,N_523);
or U1916 (N_1916,N_837,N_25);
nor U1917 (N_1917,N_3,N_907);
and U1918 (N_1918,N_531,N_726);
nand U1919 (N_1919,N_314,N_640);
nor U1920 (N_1920,N_569,N_551);
xnor U1921 (N_1921,N_862,N_960);
nand U1922 (N_1922,N_986,N_652);
nor U1923 (N_1923,N_202,N_994);
and U1924 (N_1924,N_646,N_117);
nor U1925 (N_1925,N_468,N_503);
nand U1926 (N_1926,N_396,N_997);
nor U1927 (N_1927,N_190,N_191);
nor U1928 (N_1928,N_317,N_387);
nand U1929 (N_1929,N_999,N_723);
nand U1930 (N_1930,N_56,N_921);
xor U1931 (N_1931,N_433,N_831);
or U1932 (N_1932,N_105,N_576);
nor U1933 (N_1933,N_106,N_951);
or U1934 (N_1934,N_238,N_569);
nand U1935 (N_1935,N_778,N_381);
nand U1936 (N_1936,N_388,N_491);
and U1937 (N_1937,N_280,N_770);
or U1938 (N_1938,N_675,N_102);
nor U1939 (N_1939,N_478,N_627);
and U1940 (N_1940,N_519,N_723);
nand U1941 (N_1941,N_102,N_359);
nand U1942 (N_1942,N_419,N_353);
or U1943 (N_1943,N_408,N_585);
xnor U1944 (N_1944,N_184,N_233);
or U1945 (N_1945,N_262,N_59);
nand U1946 (N_1946,N_410,N_814);
or U1947 (N_1947,N_25,N_850);
or U1948 (N_1948,N_625,N_206);
or U1949 (N_1949,N_346,N_199);
nand U1950 (N_1950,N_194,N_891);
nand U1951 (N_1951,N_594,N_322);
nor U1952 (N_1952,N_730,N_899);
nand U1953 (N_1953,N_493,N_341);
nor U1954 (N_1954,N_252,N_0);
or U1955 (N_1955,N_861,N_326);
nand U1956 (N_1956,N_120,N_358);
or U1957 (N_1957,N_444,N_614);
nor U1958 (N_1958,N_342,N_216);
or U1959 (N_1959,N_622,N_18);
and U1960 (N_1960,N_494,N_325);
xnor U1961 (N_1961,N_66,N_207);
or U1962 (N_1962,N_481,N_857);
or U1963 (N_1963,N_756,N_899);
nand U1964 (N_1964,N_836,N_102);
and U1965 (N_1965,N_959,N_662);
or U1966 (N_1966,N_479,N_790);
nor U1967 (N_1967,N_572,N_85);
and U1968 (N_1968,N_308,N_476);
nor U1969 (N_1969,N_852,N_13);
nor U1970 (N_1970,N_572,N_284);
nor U1971 (N_1971,N_986,N_227);
or U1972 (N_1972,N_436,N_505);
nand U1973 (N_1973,N_214,N_470);
nand U1974 (N_1974,N_951,N_497);
or U1975 (N_1975,N_274,N_894);
nor U1976 (N_1976,N_917,N_189);
and U1977 (N_1977,N_933,N_955);
nand U1978 (N_1978,N_176,N_836);
nor U1979 (N_1979,N_552,N_243);
or U1980 (N_1980,N_491,N_387);
nor U1981 (N_1981,N_666,N_723);
nand U1982 (N_1982,N_450,N_38);
or U1983 (N_1983,N_240,N_713);
or U1984 (N_1984,N_129,N_836);
or U1985 (N_1985,N_809,N_443);
or U1986 (N_1986,N_494,N_889);
nor U1987 (N_1987,N_400,N_590);
and U1988 (N_1988,N_161,N_874);
nand U1989 (N_1989,N_678,N_781);
or U1990 (N_1990,N_491,N_266);
nor U1991 (N_1991,N_357,N_565);
and U1992 (N_1992,N_500,N_783);
and U1993 (N_1993,N_574,N_146);
and U1994 (N_1994,N_477,N_217);
nand U1995 (N_1995,N_954,N_692);
nor U1996 (N_1996,N_47,N_814);
nor U1997 (N_1997,N_372,N_873);
or U1998 (N_1998,N_861,N_217);
nor U1999 (N_1999,N_836,N_304);
nand U2000 (N_2000,N_1363,N_1808);
nor U2001 (N_2001,N_1019,N_1612);
xor U2002 (N_2002,N_1995,N_1846);
or U2003 (N_2003,N_1993,N_1024);
or U2004 (N_2004,N_1869,N_1634);
or U2005 (N_2005,N_1134,N_1112);
or U2006 (N_2006,N_1294,N_1262);
nor U2007 (N_2007,N_1248,N_1959);
nor U2008 (N_2008,N_1898,N_1657);
or U2009 (N_2009,N_1289,N_1978);
nor U2010 (N_2010,N_1949,N_1989);
and U2011 (N_2011,N_1558,N_1584);
nor U2012 (N_2012,N_1072,N_1255);
nand U2013 (N_2013,N_1656,N_1958);
nand U2014 (N_2014,N_1256,N_1912);
nand U2015 (N_2015,N_1629,N_1088);
nor U2016 (N_2016,N_1849,N_1827);
xor U2017 (N_2017,N_1644,N_1353);
nor U2018 (N_2018,N_1118,N_1204);
and U2019 (N_2019,N_1382,N_1527);
and U2020 (N_2020,N_1415,N_1573);
nand U2021 (N_2021,N_1461,N_1055);
nor U2022 (N_2022,N_1409,N_1696);
nor U2023 (N_2023,N_1392,N_1329);
and U2024 (N_2024,N_1891,N_1040);
nand U2025 (N_2025,N_1609,N_1886);
and U2026 (N_2026,N_1467,N_1041);
nand U2027 (N_2027,N_1483,N_1351);
and U2028 (N_2028,N_1525,N_1709);
and U2029 (N_2029,N_1556,N_1954);
nor U2030 (N_2030,N_1571,N_1726);
nor U2031 (N_2031,N_1951,N_1970);
or U2032 (N_2032,N_1154,N_1037);
nor U2033 (N_2033,N_1356,N_1602);
nor U2034 (N_2034,N_1606,N_1457);
or U2035 (N_2035,N_1651,N_1401);
and U2036 (N_2036,N_1851,N_1840);
nor U2037 (N_2037,N_1038,N_1318);
and U2038 (N_2038,N_1099,N_1747);
and U2039 (N_2039,N_1812,N_1131);
and U2040 (N_2040,N_1281,N_1589);
nand U2041 (N_2041,N_1463,N_1716);
or U2042 (N_2042,N_1637,N_1981);
and U2043 (N_2043,N_1877,N_1526);
nand U2044 (N_2044,N_1247,N_1101);
and U2045 (N_2045,N_1772,N_1331);
or U2046 (N_2046,N_1321,N_1945);
or U2047 (N_2047,N_1355,N_1374);
nor U2048 (N_2048,N_1199,N_1446);
nor U2049 (N_2049,N_1727,N_1142);
and U2050 (N_2050,N_1883,N_1557);
nand U2051 (N_2051,N_1311,N_1767);
nor U2052 (N_2052,N_1383,N_1505);
and U2053 (N_2053,N_1487,N_1292);
nor U2054 (N_2054,N_1962,N_1855);
and U2055 (N_2055,N_1793,N_1626);
nand U2056 (N_2056,N_1802,N_1701);
nor U2057 (N_2057,N_1964,N_1439);
or U2058 (N_2058,N_1650,N_1595);
and U2059 (N_2059,N_1820,N_1391);
or U2060 (N_2060,N_1371,N_1147);
nor U2061 (N_2061,N_1049,N_1502);
xnor U2062 (N_2062,N_1313,N_1358);
and U2063 (N_2063,N_1148,N_1575);
nor U2064 (N_2064,N_1937,N_1717);
nand U2065 (N_2065,N_1053,N_1455);
and U2066 (N_2066,N_1619,N_1264);
nand U2067 (N_2067,N_1296,N_1744);
nand U2068 (N_2068,N_1544,N_1865);
nor U2069 (N_2069,N_1508,N_1452);
or U2070 (N_2070,N_1210,N_1996);
nor U2071 (N_2071,N_1690,N_1639);
or U2072 (N_2072,N_1135,N_1672);
and U2073 (N_2073,N_1509,N_1089);
or U2074 (N_2074,N_1122,N_1555);
nand U2075 (N_2075,N_1934,N_1233);
nor U2076 (N_2076,N_1938,N_1769);
nand U2077 (N_2077,N_1221,N_1532);
and U2078 (N_2078,N_1149,N_1316);
nor U2079 (N_2079,N_1218,N_1920);
and U2080 (N_2080,N_1939,N_1488);
or U2081 (N_2081,N_1910,N_1501);
or U2082 (N_2082,N_1539,N_1841);
nor U2083 (N_2083,N_1976,N_1381);
nand U2084 (N_2084,N_1577,N_1469);
nand U2085 (N_2085,N_1194,N_1493);
xnor U2086 (N_2086,N_1043,N_1163);
nand U2087 (N_2087,N_1359,N_1139);
nand U2088 (N_2088,N_1424,N_1327);
or U2089 (N_2089,N_1064,N_1832);
nor U2090 (N_2090,N_1087,N_1432);
or U2091 (N_2091,N_1091,N_1715);
nor U2092 (N_2092,N_1541,N_1155);
and U2093 (N_2093,N_1343,N_1130);
nand U2094 (N_2094,N_1216,N_1412);
or U2095 (N_2095,N_1279,N_1414);
or U2096 (N_2096,N_1816,N_1896);
nor U2097 (N_2097,N_1132,N_1404);
nor U2098 (N_2098,N_1591,N_1862);
nor U2099 (N_2099,N_1025,N_1385);
and U2100 (N_2100,N_1295,N_1029);
and U2101 (N_2101,N_1164,N_1031);
nand U2102 (N_2102,N_1004,N_1915);
nor U2103 (N_2103,N_1092,N_1000);
and U2104 (N_2104,N_1007,N_1572);
or U2105 (N_2105,N_1106,N_1514);
xnor U2106 (N_2106,N_1183,N_1309);
or U2107 (N_2107,N_1528,N_1018);
nand U2108 (N_2108,N_1687,N_1021);
or U2109 (N_2109,N_1330,N_1740);
nor U2110 (N_2110,N_1341,N_1593);
or U2111 (N_2111,N_1789,N_1080);
nor U2112 (N_2112,N_1983,N_1608);
nor U2113 (N_2113,N_1357,N_1227);
and U2114 (N_2114,N_1002,N_1839);
and U2115 (N_2115,N_1073,N_1235);
nand U2116 (N_2116,N_1834,N_1868);
nor U2117 (N_2117,N_1662,N_1418);
or U2118 (N_2118,N_1748,N_1536);
and U2119 (N_2119,N_1731,N_1523);
and U2120 (N_2120,N_1465,N_1624);
nor U2121 (N_2121,N_1191,N_1882);
nand U2122 (N_2122,N_1923,N_1686);
and U2123 (N_2123,N_1746,N_1105);
nor U2124 (N_2124,N_1429,N_1047);
or U2125 (N_2125,N_1873,N_1678);
nand U2126 (N_2126,N_1236,N_1177);
nand U2127 (N_2127,N_1638,N_1046);
or U2128 (N_2128,N_1661,N_1518);
and U2129 (N_2129,N_1943,N_1707);
and U2130 (N_2130,N_1157,N_1395);
nor U2131 (N_2131,N_1187,N_1704);
and U2132 (N_2132,N_1110,N_1322);
nand U2133 (N_2133,N_1421,N_1909);
nand U2134 (N_2134,N_1553,N_1646);
nor U2135 (N_2135,N_1984,N_1173);
nor U2136 (N_2136,N_1082,N_1090);
or U2137 (N_2137,N_1334,N_1766);
and U2138 (N_2138,N_1585,N_1876);
and U2139 (N_2139,N_1344,N_1141);
nor U2140 (N_2140,N_1145,N_1688);
and U2141 (N_2141,N_1914,N_1997);
or U2142 (N_2142,N_1534,N_1160);
or U2143 (N_2143,N_1115,N_1339);
nand U2144 (N_2144,N_1551,N_1070);
and U2145 (N_2145,N_1538,N_1211);
nor U2146 (N_2146,N_1590,N_1314);
or U2147 (N_2147,N_1396,N_1197);
and U2148 (N_2148,N_1420,N_1710);
or U2149 (N_2149,N_1621,N_1161);
nor U2150 (N_2150,N_1611,N_1172);
nand U2151 (N_2151,N_1065,N_1928);
or U2152 (N_2152,N_1213,N_1918);
and U2153 (N_2153,N_1966,N_1084);
or U2154 (N_2154,N_1299,N_1464);
nand U2155 (N_2155,N_1794,N_1857);
or U2156 (N_2156,N_1494,N_1228);
or U2157 (N_2157,N_1773,N_1323);
or U2158 (N_2158,N_1474,N_1618);
xor U2159 (N_2159,N_1016,N_1947);
and U2160 (N_2160,N_1471,N_1006);
or U2161 (N_2161,N_1009,N_1725);
nor U2162 (N_2162,N_1360,N_1413);
nor U2163 (N_2163,N_1893,N_1307);
xor U2164 (N_2164,N_1998,N_1133);
xnor U2165 (N_2165,N_1231,N_1114);
or U2166 (N_2166,N_1922,N_1303);
xnor U2167 (N_2167,N_1033,N_1535);
and U2168 (N_2168,N_1480,N_1190);
and U2169 (N_2169,N_1765,N_1908);
or U2170 (N_2170,N_1251,N_1434);
nand U2171 (N_2171,N_1079,N_1955);
and U2172 (N_2172,N_1890,N_1200);
nor U2173 (N_2173,N_1430,N_1614);
xor U2174 (N_2174,N_1405,N_1306);
nor U2175 (N_2175,N_1921,N_1506);
or U2176 (N_2176,N_1482,N_1859);
or U2177 (N_2177,N_1692,N_1833);
nor U2178 (N_2178,N_1278,N_1179);
or U2179 (N_2179,N_1174,N_1346);
and U2180 (N_2180,N_1677,N_1596);
nand U2181 (N_2181,N_1290,N_1098);
nor U2182 (N_2182,N_1705,N_1856);
or U2183 (N_2183,N_1689,N_1598);
nand U2184 (N_2184,N_1987,N_1270);
and U2185 (N_2185,N_1843,N_1051);
or U2186 (N_2186,N_1991,N_1074);
nor U2187 (N_2187,N_1354,N_1529);
and U2188 (N_2188,N_1503,N_1979);
and U2189 (N_2189,N_1932,N_1762);
nor U2190 (N_2190,N_1673,N_1953);
and U2191 (N_2191,N_1887,N_1874);
nand U2192 (N_2192,N_1718,N_1956);
and U2193 (N_2193,N_1260,N_1653);
or U2194 (N_2194,N_1108,N_1237);
and U2195 (N_2195,N_1837,N_1165);
nor U2196 (N_2196,N_1060,N_1378);
and U2197 (N_2197,N_1836,N_1974);
and U2198 (N_2198,N_1445,N_1902);
and U2199 (N_2199,N_1504,N_1093);
or U2200 (N_2200,N_1205,N_1076);
nor U2201 (N_2201,N_1096,N_1950);
nand U2202 (N_2202,N_1048,N_1340);
nand U2203 (N_2203,N_1436,N_1623);
or U2204 (N_2204,N_1522,N_1500);
and U2205 (N_2205,N_1805,N_1138);
nor U2206 (N_2206,N_1790,N_1507);
and U2207 (N_2207,N_1610,N_1783);
and U2208 (N_2208,N_1771,N_1062);
or U2209 (N_2209,N_1711,N_1150);
and U2210 (N_2210,N_1086,N_1485);
nor U2211 (N_2211,N_1659,N_1977);
nor U2212 (N_2212,N_1971,N_1906);
and U2213 (N_2213,N_1581,N_1751);
or U2214 (N_2214,N_1652,N_1636);
or U2215 (N_2215,N_1373,N_1389);
nor U2216 (N_2216,N_1015,N_1817);
or U2217 (N_2217,N_1261,N_1372);
nor U2218 (N_2218,N_1103,N_1540);
nor U2219 (N_2219,N_1907,N_1472);
or U2220 (N_2220,N_1450,N_1333);
nand U2221 (N_2221,N_1775,N_1369);
nor U2222 (N_2222,N_1246,N_1059);
or U2223 (N_2223,N_1056,N_1215);
or U2224 (N_2224,N_1599,N_1022);
nor U2225 (N_2225,N_1470,N_1967);
and U2226 (N_2226,N_1100,N_1752);
or U2227 (N_2227,N_1377,N_1753);
nand U2228 (N_2228,N_1668,N_1604);
and U2229 (N_2229,N_1824,N_1738);
and U2230 (N_2230,N_1061,N_1444);
nor U2231 (N_2231,N_1083,N_1592);
and U2232 (N_2232,N_1328,N_1517);
nand U2233 (N_2233,N_1003,N_1380);
xor U2234 (N_2234,N_1714,N_1230);
and U2235 (N_2235,N_1315,N_1800);
nor U2236 (N_2236,N_1326,N_1742);
nand U2237 (N_2237,N_1274,N_1858);
or U2238 (N_2238,N_1900,N_1588);
and U2239 (N_2239,N_1104,N_1167);
and U2240 (N_2240,N_1933,N_1854);
or U2241 (N_2241,N_1969,N_1466);
nor U2242 (N_2242,N_1630,N_1224);
nand U2243 (N_2243,N_1397,N_1437);
nand U2244 (N_2244,N_1683,N_1697);
nor U2245 (N_2245,N_1669,N_1613);
nor U2246 (N_2246,N_1667,N_1510);
nand U2247 (N_2247,N_1497,N_1885);
nor U2248 (N_2248,N_1407,N_1879);
nor U2249 (N_2249,N_1564,N_1113);
and U2250 (N_2250,N_1399,N_1180);
nor U2251 (N_2251,N_1924,N_1283);
nand U2252 (N_2252,N_1797,N_1988);
or U2253 (N_2253,N_1394,N_1499);
nor U2254 (N_2254,N_1804,N_1565);
and U2255 (N_2255,N_1069,N_1081);
nand U2256 (N_2256,N_1664,N_1498);
or U2257 (N_2257,N_1530,N_1301);
or U2258 (N_2258,N_1763,N_1756);
nand U2259 (N_2259,N_1778,N_1468);
and U2260 (N_2260,N_1347,N_1645);
and U2261 (N_2261,N_1288,N_1764);
nor U2262 (N_2262,N_1884,N_1878);
nand U2263 (N_2263,N_1807,N_1403);
and U2264 (N_2264,N_1724,N_1120);
and U2265 (N_2265,N_1578,N_1214);
nor U2266 (N_2266,N_1513,N_1719);
nand U2267 (N_2267,N_1121,N_1128);
or U2268 (N_2268,N_1680,N_1562);
xor U2269 (N_2269,N_1594,N_1124);
nand U2270 (N_2270,N_1566,N_1182);
or U2271 (N_2271,N_1484,N_1181);
nand U2272 (N_2272,N_1102,N_1745);
nor U2273 (N_2273,N_1750,N_1732);
or U2274 (N_2274,N_1675,N_1563);
or U2275 (N_2275,N_1512,N_1853);
nand U2276 (N_2276,N_1768,N_1760);
nor U2277 (N_2277,N_1814,N_1297);
or U2278 (N_2278,N_1202,N_1994);
xnor U2279 (N_2279,N_1207,N_1332);
xnor U2280 (N_2280,N_1250,N_1459);
or U2281 (N_2281,N_1030,N_1166);
nand U2282 (N_2282,N_1941,N_1175);
and U2283 (N_2283,N_1861,N_1111);
or U2284 (N_2284,N_1903,N_1695);
nor U2285 (N_2285,N_1039,N_1402);
or U2286 (N_2286,N_1901,N_1273);
nor U2287 (N_2287,N_1348,N_1416);
nor U2288 (N_2288,N_1521,N_1317);
and U2289 (N_2289,N_1244,N_1223);
nand U2290 (N_2290,N_1208,N_1694);
or U2291 (N_2291,N_1511,N_1684);
nand U2292 (N_2292,N_1203,N_1872);
nor U2293 (N_2293,N_1075,N_1567);
nand U2294 (N_2294,N_1011,N_1904);
and U2295 (N_2295,N_1842,N_1587);
nor U2296 (N_2296,N_1935,N_1944);
nand U2297 (N_2297,N_1735,N_1828);
or U2298 (N_2298,N_1643,N_1058);
nor U2299 (N_2299,N_1796,N_1546);
or U2300 (N_2300,N_1779,N_1533);
or U2301 (N_2301,N_1232,N_1400);
and U2302 (N_2302,N_1655,N_1212);
or U2303 (N_2303,N_1350,N_1308);
or U2304 (N_2304,N_1813,N_1368);
nand U2305 (N_2305,N_1607,N_1312);
nand U2306 (N_2306,N_1137,N_1543);
and U2307 (N_2307,N_1892,N_1952);
nor U2308 (N_2308,N_1671,N_1927);
nand U2309 (N_2309,N_1960,N_1780);
or U2310 (N_2310,N_1860,N_1554);
or U2311 (N_2311,N_1806,N_1801);
and U2312 (N_2312,N_1616,N_1542);
nand U2313 (N_2313,N_1784,N_1123);
or U2314 (N_2314,N_1980,N_1050);
and U2315 (N_2315,N_1442,N_1001);
or U2316 (N_2316,N_1552,N_1880);
nand U2317 (N_2317,N_1254,N_1515);
and U2318 (N_2318,N_1095,N_1631);
nor U2319 (N_2319,N_1835,N_1693);
nand U2320 (N_2320,N_1739,N_1435);
nand U2321 (N_2321,N_1973,N_1940);
or U2322 (N_2322,N_1449,N_1440);
nand U2323 (N_2323,N_1489,N_1819);
nand U2324 (N_2324,N_1282,N_1263);
or U2325 (N_2325,N_1781,N_1829);
or U2326 (N_2326,N_1319,N_1052);
nand U2327 (N_2327,N_1729,N_1786);
nor U2328 (N_2328,N_1185,N_1028);
nor U2329 (N_2329,N_1097,N_1479);
and U2330 (N_2330,N_1085,N_1017);
nor U2331 (N_2331,N_1478,N_1803);
nand U2332 (N_2332,N_1754,N_1008);
nand U2333 (N_2333,N_1601,N_1476);
and U2334 (N_2334,N_1032,N_1580);
or U2335 (N_2335,N_1545,N_1791);
or U2336 (N_2336,N_1603,N_1845);
nor U2337 (N_2337,N_1929,N_1225);
or U2338 (N_2338,N_1345,N_1700);
nor U2339 (N_2339,N_1127,N_1641);
and U2340 (N_2340,N_1811,N_1774);
nand U2341 (N_2341,N_1447,N_1384);
nor U2342 (N_2342,N_1229,N_1422);
or U2343 (N_2343,N_1799,N_1293);
nand U2344 (N_2344,N_1240,N_1605);
or U2345 (N_2345,N_1077,N_1335);
nor U2346 (N_2346,N_1792,N_1965);
nor U2347 (N_2347,N_1245,N_1268);
nand U2348 (N_2348,N_1579,N_1170);
or U2349 (N_2349,N_1777,N_1438);
xnor U2350 (N_2350,N_1126,N_1252);
nand U2351 (N_2351,N_1010,N_1276);
nor U2352 (N_2352,N_1691,N_1366);
nor U2353 (N_2353,N_1125,N_1370);
xor U2354 (N_2354,N_1448,N_1298);
or U2355 (N_2355,N_1267,N_1159);
nand U2356 (N_2356,N_1453,N_1238);
nand U2357 (N_2357,N_1776,N_1597);
nand U2358 (N_2358,N_1020,N_1866);
or U2359 (N_2359,N_1140,N_1336);
xor U2360 (N_2360,N_1728,N_1249);
nand U2361 (N_2361,N_1116,N_1682);
and U2362 (N_2362,N_1408,N_1428);
nor U2363 (N_2363,N_1875,N_1107);
and U2364 (N_2364,N_1844,N_1741);
and U2365 (N_2365,N_1045,N_1743);
nand U2366 (N_2366,N_1699,N_1109);
or U2367 (N_2367,N_1387,N_1809);
nor U2368 (N_2368,N_1291,N_1431);
nor U2369 (N_2369,N_1458,N_1733);
nand U2370 (N_2370,N_1193,N_1519);
or U2371 (N_2371,N_1433,N_1286);
or U2372 (N_2372,N_1574,N_1265);
and U2373 (N_2373,N_1156,N_1759);
or U2374 (N_2374,N_1665,N_1475);
nor U2375 (N_2375,N_1454,N_1026);
or U2376 (N_2376,N_1524,N_1917);
nor U2377 (N_2377,N_1393,N_1152);
nor U2378 (N_2378,N_1206,N_1919);
nand U2379 (N_2379,N_1184,N_1257);
nand U2380 (N_2380,N_1443,N_1491);
or U2381 (N_2381,N_1916,N_1925);
or U2382 (N_2382,N_1242,N_1153);
and U2383 (N_2383,N_1361,N_1706);
or U2384 (N_2384,N_1269,N_1698);
nand U2385 (N_2385,N_1285,N_1737);
or U2386 (N_2386,N_1831,N_1272);
or U2387 (N_2387,N_1217,N_1712);
and U2388 (N_2388,N_1419,N_1823);
nor U2389 (N_2389,N_1068,N_1492);
and U2390 (N_2390,N_1349,N_1570);
and U2391 (N_2391,N_1810,N_1337);
nor U2392 (N_2392,N_1968,N_1192);
and U2393 (N_2393,N_1826,N_1975);
nor U2394 (N_2394,N_1867,N_1375);
nor U2395 (N_2395,N_1441,N_1946);
and U2396 (N_2396,N_1734,N_1119);
nor U2397 (N_2397,N_1852,N_1226);
nor U2398 (N_2398,N_1196,N_1302);
nor U2399 (N_2399,N_1986,N_1034);
and U2400 (N_2400,N_1670,N_1266);
and U2401 (N_2401,N_1568,N_1117);
or U2402 (N_2402,N_1549,N_1129);
nor U2403 (N_2403,N_1379,N_1222);
and U2404 (N_2404,N_1930,N_1963);
and U2405 (N_2405,N_1822,N_1685);
nor U2406 (N_2406,N_1094,N_1324);
xor U2407 (N_2407,N_1146,N_1044);
and U2408 (N_2408,N_1850,N_1427);
or U2409 (N_2409,N_1036,N_1057);
xor U2410 (N_2410,N_1271,N_1894);
and U2411 (N_2411,N_1151,N_1730);
nand U2412 (N_2412,N_1035,N_1537);
nor U2413 (N_2413,N_1477,N_1189);
or U2414 (N_2414,N_1864,N_1342);
nor U2415 (N_2415,N_1171,N_1054);
nor U2416 (N_2416,N_1703,N_1663);
nand U2417 (N_2417,N_1830,N_1679);
nand U2418 (N_2418,N_1676,N_1520);
and U2419 (N_2419,N_1628,N_1486);
nand U2420 (N_2420,N_1364,N_1300);
and U2421 (N_2421,N_1490,N_1548);
nor U2422 (N_2422,N_1761,N_1338);
nand U2423 (N_2423,N_1352,N_1066);
or U2424 (N_2424,N_1736,N_1367);
or U2425 (N_2425,N_1258,N_1620);
and U2426 (N_2426,N_1666,N_1406);
or U2427 (N_2427,N_1913,N_1136);
xor U2428 (N_2428,N_1788,N_1496);
or U2429 (N_2429,N_1280,N_1818);
nand U2430 (N_2430,N_1023,N_1654);
and U2431 (N_2431,N_1582,N_1795);
and U2432 (N_2432,N_1195,N_1473);
and U2433 (N_2433,N_1905,N_1243);
or U2434 (N_2434,N_1198,N_1881);
or U2435 (N_2435,N_1460,N_1848);
or U2436 (N_2436,N_1576,N_1931);
or U2437 (N_2437,N_1757,N_1425);
nor U2438 (N_2438,N_1013,N_1325);
nand U2439 (N_2439,N_1622,N_1985);
or U2440 (N_2440,N_1895,N_1785);
nor U2441 (N_2441,N_1583,N_1681);
and U2442 (N_2442,N_1550,N_1410);
nand U2443 (N_2443,N_1495,N_1220);
or U2444 (N_2444,N_1186,N_1648);
nand U2445 (N_2445,N_1758,N_1569);
xor U2446 (N_2446,N_1516,N_1972);
nor U2447 (N_2447,N_1798,N_1012);
or U2448 (N_2448,N_1417,N_1787);
nand U2449 (N_2449,N_1948,N_1423);
and U2450 (N_2450,N_1600,N_1067);
or U2451 (N_2451,N_1310,N_1560);
nor U2452 (N_2452,N_1674,N_1559);
nand U2453 (N_2453,N_1234,N_1640);
or U2454 (N_2454,N_1642,N_1982);
nand U2455 (N_2455,N_1821,N_1723);
and U2456 (N_2456,N_1617,N_1362);
nor U2457 (N_2457,N_1889,N_1660);
or U2458 (N_2458,N_1721,N_1649);
nand U2459 (N_2459,N_1658,N_1899);
nand U2460 (N_2460,N_1411,N_1755);
nand U2461 (N_2461,N_1897,N_1277);
or U2462 (N_2462,N_1481,N_1259);
nor U2463 (N_2463,N_1547,N_1633);
nor U2464 (N_2464,N_1063,N_1770);
nor U2465 (N_2465,N_1720,N_1188);
or U2466 (N_2466,N_1936,N_1456);
nor U2467 (N_2467,N_1386,N_1168);
and U2468 (N_2468,N_1014,N_1162);
or U2469 (N_2469,N_1561,N_1926);
and U2470 (N_2470,N_1838,N_1825);
or U2471 (N_2471,N_1005,N_1847);
nor U2472 (N_2472,N_1178,N_1871);
nor U2473 (N_2473,N_1320,N_1209);
nor U2474 (N_2474,N_1999,N_1144);
nand U2475 (N_2475,N_1708,N_1647);
or U2476 (N_2476,N_1388,N_1531);
nand U2477 (N_2477,N_1702,N_1632);
xor U2478 (N_2478,N_1239,N_1241);
or U2479 (N_2479,N_1722,N_1365);
and U2480 (N_2480,N_1870,N_1305);
nor U2481 (N_2481,N_1635,N_1027);
nand U2482 (N_2482,N_1071,N_1749);
or U2483 (N_2483,N_1451,N_1275);
and U2484 (N_2484,N_1942,N_1815);
nand U2485 (N_2485,N_1287,N_1782);
nor U2486 (N_2486,N_1713,N_1219);
and U2487 (N_2487,N_1042,N_1911);
and U2488 (N_2488,N_1158,N_1957);
nor U2489 (N_2489,N_1888,N_1625);
or U2490 (N_2490,N_1253,N_1462);
and U2491 (N_2491,N_1201,N_1390);
nor U2492 (N_2492,N_1176,N_1284);
nor U2493 (N_2493,N_1992,N_1627);
nand U2494 (N_2494,N_1169,N_1990);
nand U2495 (N_2495,N_1143,N_1615);
nor U2496 (N_2496,N_1586,N_1426);
or U2497 (N_2497,N_1961,N_1078);
and U2498 (N_2498,N_1398,N_1376);
or U2499 (N_2499,N_1863,N_1304);
or U2500 (N_2500,N_1169,N_1788);
or U2501 (N_2501,N_1725,N_1008);
nor U2502 (N_2502,N_1654,N_1060);
or U2503 (N_2503,N_1234,N_1334);
xor U2504 (N_2504,N_1964,N_1059);
nor U2505 (N_2505,N_1304,N_1066);
and U2506 (N_2506,N_1924,N_1242);
nand U2507 (N_2507,N_1121,N_1003);
nand U2508 (N_2508,N_1335,N_1924);
and U2509 (N_2509,N_1880,N_1332);
nand U2510 (N_2510,N_1390,N_1722);
or U2511 (N_2511,N_1874,N_1845);
nor U2512 (N_2512,N_1421,N_1874);
and U2513 (N_2513,N_1774,N_1131);
xnor U2514 (N_2514,N_1857,N_1196);
and U2515 (N_2515,N_1370,N_1205);
nand U2516 (N_2516,N_1933,N_1835);
nor U2517 (N_2517,N_1575,N_1916);
nand U2518 (N_2518,N_1215,N_1236);
nor U2519 (N_2519,N_1279,N_1827);
and U2520 (N_2520,N_1154,N_1617);
nor U2521 (N_2521,N_1599,N_1764);
nand U2522 (N_2522,N_1657,N_1798);
nor U2523 (N_2523,N_1983,N_1131);
nand U2524 (N_2524,N_1027,N_1041);
and U2525 (N_2525,N_1243,N_1197);
and U2526 (N_2526,N_1544,N_1788);
and U2527 (N_2527,N_1976,N_1250);
nand U2528 (N_2528,N_1996,N_1106);
nor U2529 (N_2529,N_1881,N_1497);
and U2530 (N_2530,N_1439,N_1879);
or U2531 (N_2531,N_1179,N_1722);
and U2532 (N_2532,N_1470,N_1390);
nand U2533 (N_2533,N_1470,N_1300);
or U2534 (N_2534,N_1901,N_1381);
nor U2535 (N_2535,N_1825,N_1223);
nand U2536 (N_2536,N_1634,N_1072);
or U2537 (N_2537,N_1504,N_1903);
or U2538 (N_2538,N_1373,N_1789);
nand U2539 (N_2539,N_1172,N_1667);
or U2540 (N_2540,N_1252,N_1629);
or U2541 (N_2541,N_1709,N_1970);
and U2542 (N_2542,N_1343,N_1287);
nor U2543 (N_2543,N_1539,N_1913);
or U2544 (N_2544,N_1735,N_1105);
nand U2545 (N_2545,N_1877,N_1829);
nor U2546 (N_2546,N_1186,N_1177);
and U2547 (N_2547,N_1736,N_1461);
nor U2548 (N_2548,N_1504,N_1435);
and U2549 (N_2549,N_1038,N_1159);
and U2550 (N_2550,N_1984,N_1722);
xnor U2551 (N_2551,N_1705,N_1538);
nand U2552 (N_2552,N_1773,N_1664);
and U2553 (N_2553,N_1018,N_1293);
and U2554 (N_2554,N_1996,N_1389);
nor U2555 (N_2555,N_1711,N_1618);
nor U2556 (N_2556,N_1183,N_1457);
nor U2557 (N_2557,N_1605,N_1301);
nand U2558 (N_2558,N_1694,N_1897);
or U2559 (N_2559,N_1655,N_1867);
nor U2560 (N_2560,N_1371,N_1527);
or U2561 (N_2561,N_1165,N_1496);
nand U2562 (N_2562,N_1830,N_1368);
nand U2563 (N_2563,N_1155,N_1474);
nor U2564 (N_2564,N_1815,N_1335);
or U2565 (N_2565,N_1114,N_1537);
and U2566 (N_2566,N_1968,N_1246);
and U2567 (N_2567,N_1897,N_1338);
nor U2568 (N_2568,N_1299,N_1099);
or U2569 (N_2569,N_1837,N_1487);
and U2570 (N_2570,N_1617,N_1880);
nor U2571 (N_2571,N_1973,N_1355);
or U2572 (N_2572,N_1518,N_1242);
or U2573 (N_2573,N_1875,N_1171);
nor U2574 (N_2574,N_1858,N_1986);
nor U2575 (N_2575,N_1790,N_1848);
nor U2576 (N_2576,N_1692,N_1149);
or U2577 (N_2577,N_1228,N_1037);
nand U2578 (N_2578,N_1287,N_1048);
nand U2579 (N_2579,N_1610,N_1389);
and U2580 (N_2580,N_1148,N_1794);
xnor U2581 (N_2581,N_1139,N_1826);
nor U2582 (N_2582,N_1701,N_1086);
or U2583 (N_2583,N_1891,N_1494);
nand U2584 (N_2584,N_1713,N_1099);
and U2585 (N_2585,N_1922,N_1497);
and U2586 (N_2586,N_1497,N_1825);
nand U2587 (N_2587,N_1668,N_1841);
nor U2588 (N_2588,N_1822,N_1557);
or U2589 (N_2589,N_1870,N_1388);
and U2590 (N_2590,N_1779,N_1980);
and U2591 (N_2591,N_1918,N_1506);
and U2592 (N_2592,N_1418,N_1563);
or U2593 (N_2593,N_1730,N_1716);
nand U2594 (N_2594,N_1766,N_1396);
and U2595 (N_2595,N_1057,N_1031);
nor U2596 (N_2596,N_1749,N_1218);
and U2597 (N_2597,N_1689,N_1414);
nor U2598 (N_2598,N_1814,N_1122);
and U2599 (N_2599,N_1425,N_1728);
nor U2600 (N_2600,N_1183,N_1733);
nor U2601 (N_2601,N_1056,N_1937);
or U2602 (N_2602,N_1617,N_1339);
or U2603 (N_2603,N_1812,N_1563);
nor U2604 (N_2604,N_1431,N_1805);
and U2605 (N_2605,N_1991,N_1052);
and U2606 (N_2606,N_1099,N_1156);
or U2607 (N_2607,N_1149,N_1778);
and U2608 (N_2608,N_1179,N_1434);
and U2609 (N_2609,N_1548,N_1808);
nor U2610 (N_2610,N_1633,N_1631);
or U2611 (N_2611,N_1754,N_1225);
nor U2612 (N_2612,N_1680,N_1561);
and U2613 (N_2613,N_1506,N_1186);
or U2614 (N_2614,N_1577,N_1924);
nor U2615 (N_2615,N_1122,N_1761);
nand U2616 (N_2616,N_1945,N_1404);
nor U2617 (N_2617,N_1127,N_1564);
and U2618 (N_2618,N_1693,N_1632);
nor U2619 (N_2619,N_1834,N_1048);
or U2620 (N_2620,N_1241,N_1467);
nand U2621 (N_2621,N_1070,N_1744);
and U2622 (N_2622,N_1651,N_1973);
nand U2623 (N_2623,N_1325,N_1986);
or U2624 (N_2624,N_1958,N_1985);
or U2625 (N_2625,N_1689,N_1559);
nor U2626 (N_2626,N_1794,N_1062);
or U2627 (N_2627,N_1094,N_1569);
nand U2628 (N_2628,N_1305,N_1405);
and U2629 (N_2629,N_1593,N_1910);
nor U2630 (N_2630,N_1744,N_1392);
nand U2631 (N_2631,N_1456,N_1605);
nand U2632 (N_2632,N_1261,N_1362);
nand U2633 (N_2633,N_1611,N_1053);
nand U2634 (N_2634,N_1953,N_1184);
and U2635 (N_2635,N_1664,N_1198);
nor U2636 (N_2636,N_1195,N_1257);
nor U2637 (N_2637,N_1090,N_1427);
nor U2638 (N_2638,N_1141,N_1846);
and U2639 (N_2639,N_1676,N_1417);
nor U2640 (N_2640,N_1769,N_1094);
nand U2641 (N_2641,N_1259,N_1050);
or U2642 (N_2642,N_1265,N_1868);
or U2643 (N_2643,N_1584,N_1527);
or U2644 (N_2644,N_1156,N_1909);
nand U2645 (N_2645,N_1338,N_1810);
or U2646 (N_2646,N_1911,N_1250);
nor U2647 (N_2647,N_1635,N_1059);
nor U2648 (N_2648,N_1534,N_1370);
nand U2649 (N_2649,N_1398,N_1385);
or U2650 (N_2650,N_1065,N_1221);
nor U2651 (N_2651,N_1592,N_1256);
or U2652 (N_2652,N_1107,N_1918);
nand U2653 (N_2653,N_1640,N_1835);
nand U2654 (N_2654,N_1584,N_1938);
and U2655 (N_2655,N_1424,N_1682);
nand U2656 (N_2656,N_1150,N_1648);
nand U2657 (N_2657,N_1576,N_1033);
and U2658 (N_2658,N_1228,N_1032);
nand U2659 (N_2659,N_1305,N_1573);
or U2660 (N_2660,N_1776,N_1257);
or U2661 (N_2661,N_1528,N_1449);
or U2662 (N_2662,N_1060,N_1264);
nand U2663 (N_2663,N_1301,N_1228);
or U2664 (N_2664,N_1384,N_1305);
nand U2665 (N_2665,N_1301,N_1355);
or U2666 (N_2666,N_1308,N_1196);
and U2667 (N_2667,N_1582,N_1996);
or U2668 (N_2668,N_1714,N_1833);
or U2669 (N_2669,N_1823,N_1603);
nand U2670 (N_2670,N_1491,N_1195);
nand U2671 (N_2671,N_1192,N_1473);
or U2672 (N_2672,N_1493,N_1456);
nand U2673 (N_2673,N_1282,N_1932);
or U2674 (N_2674,N_1416,N_1538);
and U2675 (N_2675,N_1350,N_1420);
and U2676 (N_2676,N_1461,N_1690);
nand U2677 (N_2677,N_1810,N_1305);
or U2678 (N_2678,N_1136,N_1016);
or U2679 (N_2679,N_1004,N_1190);
or U2680 (N_2680,N_1597,N_1591);
or U2681 (N_2681,N_1124,N_1874);
or U2682 (N_2682,N_1537,N_1838);
nor U2683 (N_2683,N_1485,N_1403);
or U2684 (N_2684,N_1762,N_1892);
nor U2685 (N_2685,N_1258,N_1646);
and U2686 (N_2686,N_1962,N_1097);
and U2687 (N_2687,N_1380,N_1359);
nor U2688 (N_2688,N_1267,N_1878);
nand U2689 (N_2689,N_1353,N_1536);
nand U2690 (N_2690,N_1117,N_1791);
and U2691 (N_2691,N_1839,N_1662);
and U2692 (N_2692,N_1797,N_1500);
nand U2693 (N_2693,N_1693,N_1372);
or U2694 (N_2694,N_1532,N_1502);
or U2695 (N_2695,N_1968,N_1100);
nor U2696 (N_2696,N_1428,N_1048);
nor U2697 (N_2697,N_1969,N_1806);
nand U2698 (N_2698,N_1199,N_1221);
and U2699 (N_2699,N_1363,N_1695);
xor U2700 (N_2700,N_1024,N_1432);
nor U2701 (N_2701,N_1196,N_1115);
nand U2702 (N_2702,N_1377,N_1179);
nor U2703 (N_2703,N_1582,N_1367);
or U2704 (N_2704,N_1755,N_1554);
or U2705 (N_2705,N_1535,N_1862);
nor U2706 (N_2706,N_1276,N_1437);
nand U2707 (N_2707,N_1472,N_1603);
nor U2708 (N_2708,N_1732,N_1113);
or U2709 (N_2709,N_1197,N_1185);
or U2710 (N_2710,N_1137,N_1160);
or U2711 (N_2711,N_1715,N_1237);
nand U2712 (N_2712,N_1955,N_1461);
nand U2713 (N_2713,N_1501,N_1928);
nor U2714 (N_2714,N_1241,N_1657);
and U2715 (N_2715,N_1412,N_1467);
or U2716 (N_2716,N_1644,N_1109);
and U2717 (N_2717,N_1865,N_1477);
or U2718 (N_2718,N_1957,N_1329);
or U2719 (N_2719,N_1531,N_1761);
nand U2720 (N_2720,N_1474,N_1728);
nand U2721 (N_2721,N_1861,N_1241);
nor U2722 (N_2722,N_1483,N_1064);
nor U2723 (N_2723,N_1597,N_1066);
and U2724 (N_2724,N_1052,N_1340);
and U2725 (N_2725,N_1609,N_1468);
nor U2726 (N_2726,N_1532,N_1866);
and U2727 (N_2727,N_1246,N_1985);
and U2728 (N_2728,N_1021,N_1778);
and U2729 (N_2729,N_1928,N_1090);
or U2730 (N_2730,N_1898,N_1743);
nand U2731 (N_2731,N_1340,N_1281);
or U2732 (N_2732,N_1090,N_1172);
and U2733 (N_2733,N_1716,N_1423);
nand U2734 (N_2734,N_1735,N_1793);
nand U2735 (N_2735,N_1501,N_1154);
nor U2736 (N_2736,N_1641,N_1476);
and U2737 (N_2737,N_1520,N_1602);
or U2738 (N_2738,N_1165,N_1542);
nand U2739 (N_2739,N_1953,N_1806);
and U2740 (N_2740,N_1905,N_1988);
and U2741 (N_2741,N_1186,N_1999);
nand U2742 (N_2742,N_1652,N_1792);
and U2743 (N_2743,N_1749,N_1544);
nand U2744 (N_2744,N_1819,N_1184);
nor U2745 (N_2745,N_1898,N_1116);
and U2746 (N_2746,N_1084,N_1948);
nor U2747 (N_2747,N_1595,N_1463);
nor U2748 (N_2748,N_1895,N_1581);
or U2749 (N_2749,N_1950,N_1253);
nand U2750 (N_2750,N_1793,N_1715);
or U2751 (N_2751,N_1749,N_1962);
nor U2752 (N_2752,N_1446,N_1436);
or U2753 (N_2753,N_1451,N_1891);
and U2754 (N_2754,N_1367,N_1136);
nor U2755 (N_2755,N_1176,N_1475);
or U2756 (N_2756,N_1445,N_1832);
or U2757 (N_2757,N_1609,N_1483);
or U2758 (N_2758,N_1433,N_1065);
nand U2759 (N_2759,N_1758,N_1890);
nor U2760 (N_2760,N_1866,N_1153);
and U2761 (N_2761,N_1108,N_1094);
nor U2762 (N_2762,N_1187,N_1384);
nor U2763 (N_2763,N_1112,N_1078);
nand U2764 (N_2764,N_1875,N_1847);
nor U2765 (N_2765,N_1609,N_1807);
nand U2766 (N_2766,N_1487,N_1625);
and U2767 (N_2767,N_1048,N_1365);
or U2768 (N_2768,N_1369,N_1889);
or U2769 (N_2769,N_1101,N_1752);
or U2770 (N_2770,N_1051,N_1153);
or U2771 (N_2771,N_1313,N_1121);
or U2772 (N_2772,N_1011,N_1707);
nor U2773 (N_2773,N_1888,N_1216);
nor U2774 (N_2774,N_1446,N_1683);
nand U2775 (N_2775,N_1115,N_1825);
or U2776 (N_2776,N_1913,N_1813);
or U2777 (N_2777,N_1685,N_1382);
nand U2778 (N_2778,N_1545,N_1522);
and U2779 (N_2779,N_1925,N_1622);
xor U2780 (N_2780,N_1861,N_1550);
nand U2781 (N_2781,N_1376,N_1149);
nand U2782 (N_2782,N_1942,N_1241);
nand U2783 (N_2783,N_1892,N_1200);
and U2784 (N_2784,N_1918,N_1586);
nand U2785 (N_2785,N_1190,N_1610);
or U2786 (N_2786,N_1748,N_1374);
nor U2787 (N_2787,N_1258,N_1411);
or U2788 (N_2788,N_1578,N_1167);
nand U2789 (N_2789,N_1279,N_1870);
and U2790 (N_2790,N_1830,N_1290);
nor U2791 (N_2791,N_1055,N_1486);
nor U2792 (N_2792,N_1779,N_1382);
or U2793 (N_2793,N_1085,N_1780);
nor U2794 (N_2794,N_1157,N_1104);
nand U2795 (N_2795,N_1073,N_1079);
and U2796 (N_2796,N_1299,N_1335);
and U2797 (N_2797,N_1230,N_1167);
nand U2798 (N_2798,N_1176,N_1696);
xnor U2799 (N_2799,N_1234,N_1143);
nand U2800 (N_2800,N_1312,N_1181);
nor U2801 (N_2801,N_1183,N_1351);
or U2802 (N_2802,N_1641,N_1554);
and U2803 (N_2803,N_1146,N_1347);
or U2804 (N_2804,N_1601,N_1231);
or U2805 (N_2805,N_1492,N_1965);
or U2806 (N_2806,N_1449,N_1060);
nand U2807 (N_2807,N_1181,N_1733);
or U2808 (N_2808,N_1506,N_1317);
nor U2809 (N_2809,N_1644,N_1149);
nand U2810 (N_2810,N_1290,N_1444);
and U2811 (N_2811,N_1398,N_1770);
and U2812 (N_2812,N_1379,N_1404);
xor U2813 (N_2813,N_1665,N_1361);
xnor U2814 (N_2814,N_1484,N_1405);
and U2815 (N_2815,N_1309,N_1455);
nor U2816 (N_2816,N_1471,N_1319);
and U2817 (N_2817,N_1398,N_1940);
and U2818 (N_2818,N_1025,N_1611);
nand U2819 (N_2819,N_1636,N_1160);
nor U2820 (N_2820,N_1020,N_1849);
or U2821 (N_2821,N_1194,N_1816);
or U2822 (N_2822,N_1985,N_1245);
or U2823 (N_2823,N_1540,N_1509);
and U2824 (N_2824,N_1511,N_1434);
and U2825 (N_2825,N_1575,N_1995);
nor U2826 (N_2826,N_1579,N_1122);
or U2827 (N_2827,N_1273,N_1472);
and U2828 (N_2828,N_1396,N_1421);
nor U2829 (N_2829,N_1989,N_1906);
nor U2830 (N_2830,N_1373,N_1978);
or U2831 (N_2831,N_1741,N_1543);
xor U2832 (N_2832,N_1589,N_1918);
and U2833 (N_2833,N_1743,N_1086);
nor U2834 (N_2834,N_1612,N_1988);
and U2835 (N_2835,N_1881,N_1624);
nor U2836 (N_2836,N_1672,N_1598);
or U2837 (N_2837,N_1352,N_1437);
nor U2838 (N_2838,N_1476,N_1372);
or U2839 (N_2839,N_1933,N_1832);
or U2840 (N_2840,N_1373,N_1853);
nand U2841 (N_2841,N_1819,N_1070);
nor U2842 (N_2842,N_1105,N_1390);
and U2843 (N_2843,N_1878,N_1152);
nand U2844 (N_2844,N_1517,N_1840);
nor U2845 (N_2845,N_1180,N_1268);
or U2846 (N_2846,N_1634,N_1429);
and U2847 (N_2847,N_1544,N_1231);
nand U2848 (N_2848,N_1321,N_1742);
and U2849 (N_2849,N_1147,N_1914);
nand U2850 (N_2850,N_1072,N_1906);
nor U2851 (N_2851,N_1359,N_1580);
nor U2852 (N_2852,N_1085,N_1251);
nor U2853 (N_2853,N_1730,N_1331);
or U2854 (N_2854,N_1927,N_1410);
and U2855 (N_2855,N_1937,N_1327);
or U2856 (N_2856,N_1417,N_1186);
nor U2857 (N_2857,N_1886,N_1418);
nand U2858 (N_2858,N_1172,N_1097);
and U2859 (N_2859,N_1866,N_1393);
nand U2860 (N_2860,N_1941,N_1101);
nand U2861 (N_2861,N_1900,N_1083);
and U2862 (N_2862,N_1311,N_1959);
and U2863 (N_2863,N_1192,N_1171);
and U2864 (N_2864,N_1479,N_1996);
nand U2865 (N_2865,N_1736,N_1518);
or U2866 (N_2866,N_1412,N_1648);
nand U2867 (N_2867,N_1218,N_1959);
nor U2868 (N_2868,N_1798,N_1287);
nand U2869 (N_2869,N_1395,N_1677);
nand U2870 (N_2870,N_1748,N_1450);
nand U2871 (N_2871,N_1883,N_1242);
nand U2872 (N_2872,N_1808,N_1924);
and U2873 (N_2873,N_1322,N_1221);
and U2874 (N_2874,N_1517,N_1810);
nand U2875 (N_2875,N_1260,N_1852);
nand U2876 (N_2876,N_1411,N_1225);
or U2877 (N_2877,N_1496,N_1339);
and U2878 (N_2878,N_1744,N_1430);
nand U2879 (N_2879,N_1705,N_1376);
and U2880 (N_2880,N_1099,N_1792);
or U2881 (N_2881,N_1873,N_1689);
or U2882 (N_2882,N_1946,N_1141);
and U2883 (N_2883,N_1545,N_1692);
and U2884 (N_2884,N_1951,N_1675);
or U2885 (N_2885,N_1108,N_1388);
and U2886 (N_2886,N_1773,N_1234);
and U2887 (N_2887,N_1107,N_1302);
or U2888 (N_2888,N_1909,N_1549);
and U2889 (N_2889,N_1705,N_1809);
and U2890 (N_2890,N_1259,N_1641);
or U2891 (N_2891,N_1914,N_1225);
and U2892 (N_2892,N_1348,N_1487);
or U2893 (N_2893,N_1945,N_1498);
nand U2894 (N_2894,N_1848,N_1516);
xor U2895 (N_2895,N_1066,N_1485);
nor U2896 (N_2896,N_1185,N_1944);
nor U2897 (N_2897,N_1921,N_1381);
nand U2898 (N_2898,N_1878,N_1007);
and U2899 (N_2899,N_1151,N_1238);
and U2900 (N_2900,N_1323,N_1762);
and U2901 (N_2901,N_1252,N_1678);
nand U2902 (N_2902,N_1242,N_1123);
and U2903 (N_2903,N_1054,N_1556);
nand U2904 (N_2904,N_1885,N_1560);
nor U2905 (N_2905,N_1448,N_1325);
nor U2906 (N_2906,N_1947,N_1168);
or U2907 (N_2907,N_1813,N_1789);
or U2908 (N_2908,N_1848,N_1670);
and U2909 (N_2909,N_1812,N_1224);
nor U2910 (N_2910,N_1069,N_1687);
or U2911 (N_2911,N_1868,N_1590);
and U2912 (N_2912,N_1649,N_1821);
and U2913 (N_2913,N_1955,N_1448);
and U2914 (N_2914,N_1990,N_1561);
nand U2915 (N_2915,N_1882,N_1817);
or U2916 (N_2916,N_1842,N_1661);
xor U2917 (N_2917,N_1036,N_1292);
nor U2918 (N_2918,N_1774,N_1887);
nand U2919 (N_2919,N_1024,N_1361);
or U2920 (N_2920,N_1084,N_1930);
nand U2921 (N_2921,N_1633,N_1450);
nand U2922 (N_2922,N_1621,N_1423);
xnor U2923 (N_2923,N_1260,N_1293);
xor U2924 (N_2924,N_1009,N_1890);
or U2925 (N_2925,N_1995,N_1737);
or U2926 (N_2926,N_1127,N_1787);
or U2927 (N_2927,N_1444,N_1044);
or U2928 (N_2928,N_1742,N_1618);
nor U2929 (N_2929,N_1426,N_1348);
xnor U2930 (N_2930,N_1689,N_1429);
and U2931 (N_2931,N_1603,N_1457);
or U2932 (N_2932,N_1341,N_1119);
and U2933 (N_2933,N_1955,N_1816);
or U2934 (N_2934,N_1260,N_1573);
nand U2935 (N_2935,N_1388,N_1445);
nor U2936 (N_2936,N_1163,N_1528);
and U2937 (N_2937,N_1261,N_1606);
nor U2938 (N_2938,N_1335,N_1865);
nand U2939 (N_2939,N_1319,N_1562);
and U2940 (N_2940,N_1333,N_1514);
nor U2941 (N_2941,N_1668,N_1930);
or U2942 (N_2942,N_1538,N_1697);
nand U2943 (N_2943,N_1273,N_1016);
nor U2944 (N_2944,N_1308,N_1618);
or U2945 (N_2945,N_1173,N_1717);
and U2946 (N_2946,N_1508,N_1259);
nor U2947 (N_2947,N_1939,N_1721);
nor U2948 (N_2948,N_1486,N_1383);
and U2949 (N_2949,N_1386,N_1267);
and U2950 (N_2950,N_1716,N_1752);
nor U2951 (N_2951,N_1262,N_1920);
and U2952 (N_2952,N_1207,N_1560);
xnor U2953 (N_2953,N_1926,N_1795);
or U2954 (N_2954,N_1235,N_1344);
xor U2955 (N_2955,N_1580,N_1333);
nor U2956 (N_2956,N_1992,N_1921);
or U2957 (N_2957,N_1676,N_1008);
nand U2958 (N_2958,N_1768,N_1628);
nor U2959 (N_2959,N_1007,N_1628);
nand U2960 (N_2960,N_1001,N_1898);
nand U2961 (N_2961,N_1124,N_1161);
nand U2962 (N_2962,N_1743,N_1339);
nor U2963 (N_2963,N_1411,N_1115);
or U2964 (N_2964,N_1627,N_1106);
nor U2965 (N_2965,N_1190,N_1638);
or U2966 (N_2966,N_1376,N_1255);
or U2967 (N_2967,N_1741,N_1763);
and U2968 (N_2968,N_1604,N_1387);
or U2969 (N_2969,N_1597,N_1318);
xnor U2970 (N_2970,N_1739,N_1529);
nor U2971 (N_2971,N_1961,N_1415);
nand U2972 (N_2972,N_1404,N_1423);
nand U2973 (N_2973,N_1404,N_1849);
or U2974 (N_2974,N_1385,N_1927);
or U2975 (N_2975,N_1312,N_1083);
and U2976 (N_2976,N_1259,N_1091);
nor U2977 (N_2977,N_1684,N_1968);
nor U2978 (N_2978,N_1502,N_1566);
nand U2979 (N_2979,N_1481,N_1844);
and U2980 (N_2980,N_1962,N_1447);
and U2981 (N_2981,N_1737,N_1784);
and U2982 (N_2982,N_1106,N_1372);
or U2983 (N_2983,N_1799,N_1610);
and U2984 (N_2984,N_1982,N_1443);
and U2985 (N_2985,N_1709,N_1169);
xor U2986 (N_2986,N_1850,N_1100);
nor U2987 (N_2987,N_1638,N_1777);
and U2988 (N_2988,N_1103,N_1547);
nand U2989 (N_2989,N_1164,N_1707);
or U2990 (N_2990,N_1517,N_1440);
nor U2991 (N_2991,N_1136,N_1598);
nor U2992 (N_2992,N_1343,N_1635);
and U2993 (N_2993,N_1251,N_1040);
nand U2994 (N_2994,N_1315,N_1634);
nand U2995 (N_2995,N_1668,N_1123);
nor U2996 (N_2996,N_1740,N_1244);
nor U2997 (N_2997,N_1460,N_1217);
nand U2998 (N_2998,N_1326,N_1920);
xnor U2999 (N_2999,N_1884,N_1299);
and U3000 (N_3000,N_2611,N_2039);
and U3001 (N_3001,N_2449,N_2552);
xor U3002 (N_3002,N_2754,N_2704);
and U3003 (N_3003,N_2154,N_2027);
and U3004 (N_3004,N_2346,N_2213);
nor U3005 (N_3005,N_2999,N_2226);
nand U3006 (N_3006,N_2003,N_2814);
or U3007 (N_3007,N_2526,N_2418);
nor U3008 (N_3008,N_2229,N_2730);
and U3009 (N_3009,N_2087,N_2473);
or U3010 (N_3010,N_2403,N_2189);
or U3011 (N_3011,N_2782,N_2273);
or U3012 (N_3012,N_2053,N_2176);
nand U3013 (N_3013,N_2125,N_2139);
nand U3014 (N_3014,N_2873,N_2299);
and U3015 (N_3015,N_2885,N_2543);
nor U3016 (N_3016,N_2155,N_2617);
and U3017 (N_3017,N_2729,N_2641);
or U3018 (N_3018,N_2806,N_2977);
nor U3019 (N_3019,N_2853,N_2815);
and U3020 (N_3020,N_2111,N_2913);
nand U3021 (N_3021,N_2162,N_2973);
or U3022 (N_3022,N_2394,N_2654);
nand U3023 (N_3023,N_2942,N_2374);
nand U3024 (N_3024,N_2514,N_2080);
xor U3025 (N_3025,N_2347,N_2925);
and U3026 (N_3026,N_2276,N_2326);
or U3027 (N_3027,N_2684,N_2257);
nand U3028 (N_3028,N_2601,N_2996);
and U3029 (N_3029,N_2777,N_2470);
and U3030 (N_3030,N_2126,N_2203);
and U3031 (N_3031,N_2673,N_2370);
or U3032 (N_3032,N_2796,N_2043);
nand U3033 (N_3033,N_2421,N_2739);
nor U3034 (N_3034,N_2545,N_2002);
nor U3035 (N_3035,N_2381,N_2854);
nor U3036 (N_3036,N_2635,N_2882);
and U3037 (N_3037,N_2842,N_2696);
nor U3038 (N_3038,N_2931,N_2095);
or U3039 (N_3039,N_2577,N_2303);
or U3040 (N_3040,N_2339,N_2210);
nor U3041 (N_3041,N_2822,N_2305);
and U3042 (N_3042,N_2817,N_2855);
and U3043 (N_3043,N_2352,N_2711);
or U3044 (N_3044,N_2681,N_2513);
nor U3045 (N_3045,N_2900,N_2354);
and U3046 (N_3046,N_2300,N_2254);
or U3047 (N_3047,N_2712,N_2533);
nand U3048 (N_3048,N_2741,N_2389);
nor U3049 (N_3049,N_2546,N_2458);
or U3050 (N_3050,N_2978,N_2109);
and U3051 (N_3051,N_2564,N_2489);
and U3052 (N_3052,N_2117,N_2959);
or U3053 (N_3053,N_2140,N_2851);
xor U3054 (N_3054,N_2350,N_2762);
or U3055 (N_3055,N_2197,N_2048);
or U3056 (N_3056,N_2718,N_2081);
or U3057 (N_3057,N_2523,N_2905);
nor U3058 (N_3058,N_2287,N_2674);
and U3059 (N_3059,N_2809,N_2258);
xor U3060 (N_3060,N_2264,N_2613);
nor U3061 (N_3061,N_2634,N_2773);
and U3062 (N_3062,N_2883,N_2160);
or U3063 (N_3063,N_2726,N_2693);
and U3064 (N_3064,N_2791,N_2450);
nand U3065 (N_3065,N_2093,N_2889);
xor U3066 (N_3066,N_2290,N_2929);
xor U3067 (N_3067,N_2519,N_2636);
nand U3068 (N_3068,N_2887,N_2753);
or U3069 (N_3069,N_2261,N_2844);
or U3070 (N_3070,N_2628,N_2946);
nand U3071 (N_3071,N_2001,N_2823);
or U3072 (N_3072,N_2733,N_2735);
nor U3073 (N_3073,N_2790,N_2721);
or U3074 (N_3074,N_2677,N_2472);
or U3075 (N_3075,N_2541,N_2411);
xor U3076 (N_3076,N_2983,N_2644);
nor U3077 (N_3077,N_2171,N_2255);
and U3078 (N_3078,N_2870,N_2474);
or U3079 (N_3079,N_2625,N_2938);
and U3080 (N_3080,N_2186,N_2420);
nand U3081 (N_3081,N_2172,N_2372);
xnor U3082 (N_3082,N_2914,N_2891);
nand U3083 (N_3083,N_2764,N_2521);
and U3084 (N_3084,N_2920,N_2437);
or U3085 (N_3085,N_2236,N_2344);
and U3086 (N_3086,N_2044,N_2772);
or U3087 (N_3087,N_2133,N_2868);
nor U3088 (N_3088,N_2025,N_2367);
and U3089 (N_3089,N_2046,N_2585);
nor U3090 (N_3090,N_2967,N_2917);
nor U3091 (N_3091,N_2708,N_2743);
or U3092 (N_3092,N_2579,N_2751);
nand U3093 (N_3093,N_2587,N_2981);
and U3094 (N_3094,N_2834,N_2547);
nand U3095 (N_3095,N_2167,N_2380);
nor U3096 (N_3096,N_2132,N_2476);
and U3097 (N_3097,N_2314,N_2063);
nor U3098 (N_3098,N_2205,N_2645);
nor U3099 (N_3099,N_2828,N_2832);
nand U3100 (N_3100,N_2082,N_2329);
or U3101 (N_3101,N_2477,N_2441);
or U3102 (N_3102,N_2831,N_2972);
nor U3103 (N_3103,N_2884,N_2274);
nand U3104 (N_3104,N_2976,N_2272);
and U3105 (N_3105,N_2185,N_2558);
and U3106 (N_3106,N_2121,N_2247);
nor U3107 (N_3107,N_2019,N_2734);
and U3108 (N_3108,N_2280,N_2955);
and U3109 (N_3109,N_2026,N_2237);
nand U3110 (N_3110,N_2880,N_2952);
or U3111 (N_3111,N_2899,N_2294);
or U3112 (N_3112,N_2387,N_2297);
or U3113 (N_3113,N_2997,N_2024);
nand U3114 (N_3114,N_2841,N_2151);
and U3115 (N_3115,N_2710,N_2758);
nor U3116 (N_3116,N_2149,N_2436);
nor U3117 (N_3117,N_2448,N_2402);
nor U3118 (N_3118,N_2124,N_2009);
and U3119 (N_3119,N_2138,N_2217);
nand U3120 (N_3120,N_2793,N_2985);
and U3121 (N_3121,N_2720,N_2847);
nor U3122 (N_3122,N_2505,N_2827);
or U3123 (N_3123,N_2497,N_2843);
nor U3124 (N_3124,N_2097,N_2191);
nand U3125 (N_3125,N_2695,N_2397);
or U3126 (N_3126,N_2567,N_2669);
or U3127 (N_3127,N_2962,N_2866);
nor U3128 (N_3128,N_2006,N_2408);
or U3129 (N_3129,N_2233,N_2609);
nand U3130 (N_3130,N_2618,N_2285);
or U3131 (N_3131,N_2047,N_2714);
and U3132 (N_3132,N_2454,N_2845);
nor U3133 (N_3133,N_2283,N_2965);
nand U3134 (N_3134,N_2016,N_2120);
or U3135 (N_3135,N_2115,N_2974);
nor U3136 (N_3136,N_2702,N_2486);
and U3137 (N_3137,N_2624,N_2296);
nor U3138 (N_3138,N_2935,N_2651);
and U3139 (N_3139,N_2990,N_2737);
and U3140 (N_3140,N_2595,N_2023);
nor U3141 (N_3141,N_2901,N_2622);
nand U3142 (N_3142,N_2453,N_2295);
and U3143 (N_3143,N_2788,N_2198);
and U3144 (N_3144,N_2569,N_2986);
or U3145 (N_3145,N_2424,N_2770);
and U3146 (N_3146,N_2159,N_2746);
xor U3147 (N_3147,N_2879,N_2113);
or U3148 (N_3148,N_2196,N_2908);
and U3149 (N_3149,N_2017,N_2621);
and U3150 (N_3150,N_2602,N_2607);
and U3151 (N_3151,N_2419,N_2361);
xor U3152 (N_3152,N_2086,N_2452);
and U3153 (N_3153,N_2110,N_2660);
and U3154 (N_3154,N_2262,N_2923);
and U3155 (N_3155,N_2148,N_2244);
nor U3156 (N_3156,N_2656,N_2059);
nor U3157 (N_3157,N_2667,N_2414);
nand U3158 (N_3158,N_2922,N_2833);
nor U3159 (N_3159,N_2032,N_2071);
or U3160 (N_3160,N_2020,N_2340);
or U3161 (N_3161,N_2243,N_2386);
and U3162 (N_3162,N_2252,N_2157);
xor U3163 (N_3163,N_2242,N_2096);
or U3164 (N_3164,N_2164,N_2932);
nor U3165 (N_3165,N_2649,N_2859);
or U3166 (N_3166,N_2948,N_2941);
nand U3167 (N_3167,N_2640,N_2648);
or U3168 (N_3168,N_2878,N_2936);
nand U3169 (N_3169,N_2482,N_2874);
and U3170 (N_3170,N_2553,N_2073);
xnor U3171 (N_3171,N_2334,N_2180);
and U3172 (N_3172,N_2371,N_2015);
or U3173 (N_3173,N_2864,N_2666);
nand U3174 (N_3174,N_2422,N_2218);
nand U3175 (N_3175,N_2562,N_2256);
nor U3176 (N_3176,N_2775,N_2322);
or U3177 (N_3177,N_2129,N_2893);
and U3178 (N_3178,N_2778,N_2119);
nand U3179 (N_3179,N_2443,N_2240);
nand U3180 (N_3180,N_2438,N_2811);
and U3181 (N_3181,N_2503,N_2090);
nand U3182 (N_3182,N_2916,N_2982);
nand U3183 (N_3183,N_2603,N_2532);
nand U3184 (N_3184,N_2592,N_2173);
and U3185 (N_3185,N_2200,N_2079);
nor U3186 (N_3186,N_2434,N_2789);
and U3187 (N_3187,N_2783,N_2105);
and U3188 (N_3188,N_2596,N_2423);
nor U3189 (N_3189,N_2781,N_2805);
nor U3190 (N_3190,N_2060,N_2816);
nor U3191 (N_3191,N_2131,N_2451);
nor U3192 (N_3192,N_2890,N_2515);
or U3193 (N_3193,N_2467,N_2930);
or U3194 (N_3194,N_2857,N_2707);
nand U3195 (N_3195,N_2051,N_2643);
or U3196 (N_3196,N_2747,N_2584);
nand U3197 (N_3197,N_2267,N_2561);
and U3198 (N_3198,N_2638,N_2062);
xor U3199 (N_3199,N_2038,N_2008);
nand U3200 (N_3200,N_2271,N_2365);
and U3201 (N_3201,N_2012,N_2306);
or U3202 (N_3202,N_2685,N_2837);
nand U3203 (N_3203,N_2825,N_2359);
nand U3204 (N_3204,N_2301,N_2033);
and U3205 (N_3205,N_2089,N_2413);
nor U3206 (N_3206,N_2657,N_2494);
nand U3207 (N_3207,N_2442,N_2336);
nor U3208 (N_3208,N_2934,N_2289);
and U3209 (N_3209,N_2535,N_2995);
or U3210 (N_3210,N_2668,N_2462);
nand U3211 (N_3211,N_2337,N_2376);
or U3212 (N_3212,N_2915,N_2277);
or U3213 (N_3213,N_2502,N_2223);
or U3214 (N_3214,N_2642,N_2803);
nand U3215 (N_3215,N_2591,N_2970);
nor U3216 (N_3216,N_2439,N_2364);
or U3217 (N_3217,N_2518,N_2516);
nor U3218 (N_3218,N_2328,N_2507);
nand U3219 (N_3219,N_2911,N_2130);
and U3220 (N_3220,N_2571,N_2722);
nor U3221 (N_3221,N_2145,N_2818);
nor U3222 (N_3222,N_2760,N_2598);
and U3223 (N_3223,N_2190,N_2937);
or U3224 (N_3224,N_2147,N_2517);
or U3225 (N_3225,N_2949,N_2211);
xnor U3226 (N_3226,N_2275,N_2128);
nor U3227 (N_3227,N_2534,N_2320);
xnor U3228 (N_3228,N_2589,N_2572);
and U3229 (N_3229,N_2608,N_2875);
or U3230 (N_3230,N_2716,N_2475);
nand U3231 (N_3231,N_2207,N_2583);
and U3232 (N_3232,N_2045,N_2631);
and U3233 (N_3233,N_2075,N_2975);
nand U3234 (N_3234,N_2425,N_2315);
or U3235 (N_3235,N_2780,N_2091);
nor U3236 (N_3236,N_2542,N_2539);
and U3237 (N_3237,N_2049,N_2860);
nand U3238 (N_3238,N_2525,N_2293);
nand U3239 (N_3239,N_2377,N_2566);
nor U3240 (N_3240,N_2663,N_2785);
nand U3241 (N_3241,N_2819,N_2600);
nor U3242 (N_3242,N_2554,N_2193);
and U3243 (N_3243,N_2756,N_2779);
or U3244 (N_3244,N_2736,N_2989);
or U3245 (N_3245,N_2114,N_2557);
or U3246 (N_3246,N_2118,N_2510);
nor U3247 (N_3247,N_2065,N_2444);
or U3248 (N_3248,N_2056,N_2360);
nand U3249 (N_3249,N_2500,N_2383);
nand U3250 (N_3250,N_2378,N_2688);
and U3251 (N_3251,N_2606,N_2508);
or U3252 (N_3252,N_2745,N_2070);
or U3253 (N_3253,N_2944,N_2616);
nand U3254 (N_3254,N_2083,N_2991);
nor U3255 (N_3255,N_2215,N_2013);
nor U3256 (N_3256,N_2872,N_2431);
nand U3257 (N_3257,N_2835,N_2445);
and U3258 (N_3258,N_2103,N_2522);
or U3259 (N_3259,N_2856,N_2895);
nor U3260 (N_3260,N_2061,N_2417);
or U3261 (N_3261,N_2268,N_2259);
or U3262 (N_3262,N_2331,N_2232);
nor U3263 (N_3263,N_2035,N_2491);
nor U3264 (N_3264,N_2228,N_2031);
and U3265 (N_3265,N_2776,N_2665);
nor U3266 (N_3266,N_2774,N_2456);
or U3267 (N_3267,N_2529,N_2664);
nor U3268 (N_3268,N_2281,N_2787);
nand U3269 (N_3269,N_2342,N_2187);
or U3270 (N_3270,N_2655,N_2993);
or U3271 (N_3271,N_2188,N_2333);
or U3272 (N_3272,N_2610,N_2963);
nor U3273 (N_3273,N_2440,N_2661);
nor U3274 (N_3274,N_2725,N_2980);
or U3275 (N_3275,N_2036,N_2836);
nor U3276 (N_3276,N_2538,N_2573);
nand U3277 (N_3277,N_2165,N_2263);
and U3278 (N_3278,N_2927,N_2672);
or U3279 (N_3279,N_2194,N_2094);
or U3280 (N_3280,N_2840,N_2266);
nor U3281 (N_3281,N_2216,N_2021);
nand U3282 (N_3282,N_2581,N_2169);
or U3283 (N_3283,N_2799,N_2740);
or U3284 (N_3284,N_2919,N_2954);
and U3285 (N_3285,N_2548,N_2204);
nor U3286 (N_3286,N_2988,N_2495);
and U3287 (N_3287,N_2501,N_2310);
nand U3288 (N_3288,N_2338,N_2697);
and U3289 (N_3289,N_2260,N_2373);
nand U3290 (N_3290,N_2706,N_2463);
and U3291 (N_3291,N_2028,N_2633);
nand U3292 (N_3292,N_2906,N_2368);
nand U3293 (N_3293,N_2316,N_2152);
nand U3294 (N_3294,N_2029,N_2951);
and U3295 (N_3295,N_2487,N_2245);
and U3296 (N_3296,N_2166,N_2862);
nor U3297 (N_3297,N_2100,N_2749);
nor U3298 (N_3298,N_2101,N_2112);
or U3299 (N_3299,N_2619,N_2590);
and U3300 (N_3300,N_2018,N_2848);
nor U3301 (N_3301,N_2992,N_2488);
nand U3302 (N_3302,N_2278,N_2605);
and U3303 (N_3303,N_2357,N_2536);
nand U3304 (N_3304,N_2863,N_2135);
nand U3305 (N_3305,N_2593,N_2699);
and U3306 (N_3306,N_2466,N_2395);
xnor U3307 (N_3307,N_2750,N_2524);
nor U3308 (N_3308,N_2356,N_2332);
and U3309 (N_3309,N_2231,N_2994);
nand U3310 (N_3310,N_2464,N_2947);
and U3311 (N_3311,N_2484,N_2158);
and U3312 (N_3312,N_2427,N_2682);
nand U3313 (N_3313,N_2678,N_2446);
nor U3314 (N_3314,N_2037,N_2074);
and U3315 (N_3315,N_2940,N_2214);
and U3316 (N_3316,N_2182,N_2390);
nor U3317 (N_3317,N_2400,N_2544);
nor U3318 (N_3318,N_2212,N_2597);
nor U3319 (N_3319,N_2604,N_2580);
or U3320 (N_3320,N_2909,N_2286);
nor U3321 (N_3321,N_2703,N_2221);
xnor U3322 (N_3322,N_2784,N_2924);
nor U3323 (N_3323,N_2348,N_2404);
or U3324 (N_3324,N_2050,N_2738);
nand U3325 (N_3325,N_2309,N_2201);
nor U3326 (N_3326,N_2318,N_2826);
nor U3327 (N_3327,N_2143,N_2195);
nand U3328 (N_3328,N_2964,N_2072);
and U3329 (N_3329,N_2767,N_2399);
nor U3330 (N_3330,N_2810,N_2582);
xnor U3331 (N_3331,N_2123,N_2362);
or U3332 (N_3332,N_2284,N_2904);
or U3333 (N_3333,N_2493,N_2181);
nand U3334 (N_3334,N_2483,N_2858);
and U3335 (N_3335,N_2183,N_2253);
nor U3336 (N_3336,N_2366,N_2620);
or U3337 (N_3337,N_2998,N_2385);
nand U3338 (N_3338,N_2069,N_2692);
and U3339 (N_3339,N_2680,N_2479);
nand U3340 (N_3340,N_2468,N_2892);
xnor U3341 (N_3341,N_2108,N_2269);
nand U3342 (N_3342,N_2407,N_2715);
nor U3343 (N_3343,N_2499,N_2005);
xor U3344 (N_3344,N_2798,N_2304);
nand U3345 (N_3345,N_2004,N_2064);
and U3346 (N_3346,N_2588,N_2921);
and U3347 (N_3347,N_2757,N_2179);
nor U3348 (N_3348,N_2560,N_2849);
nand U3349 (N_3349,N_2653,N_2926);
or U3350 (N_3350,N_2540,N_2933);
or U3351 (N_3351,N_2961,N_2144);
xor U3352 (N_3352,N_2612,N_2877);
nand U3353 (N_3353,N_2632,N_2786);
nand U3354 (N_3354,N_2650,N_2957);
nand U3355 (N_3355,N_2349,N_2405);
nand U3356 (N_3356,N_2675,N_2391);
nand U3357 (N_3357,N_2637,N_2690);
and U3358 (N_3358,N_2670,N_2496);
nand U3359 (N_3359,N_2614,N_2700);
nand U3360 (N_3360,N_2457,N_2969);
nor U3361 (N_3361,N_2960,N_2351);
or U3362 (N_3362,N_2490,N_2327);
or U3363 (N_3363,N_2698,N_2241);
nand U3364 (N_3364,N_2945,N_2694);
nor U3365 (N_3365,N_2898,N_2078);
nor U3366 (N_3366,N_2709,N_2506);
nor U3367 (N_3367,N_2184,N_2279);
or U3368 (N_3368,N_2528,N_2683);
nand U3369 (N_3369,N_2410,N_2918);
and U3370 (N_3370,N_2717,N_2902);
nand U3371 (N_3371,N_2801,N_2852);
and U3372 (N_3372,N_2471,N_2549);
nor U3373 (N_3373,N_2341,N_2246);
or U3374 (N_3374,N_2098,N_2409);
or U3375 (N_3375,N_2104,N_2759);
and U3376 (N_3376,N_2122,N_2550);
nor U3377 (N_3377,N_2850,N_2401);
or U3378 (N_3378,N_2379,N_2939);
nor U3379 (N_3379,N_2428,N_2594);
nor U3380 (N_3380,N_2235,N_2578);
xnor U3381 (N_3381,N_2896,N_2984);
nand U3382 (N_3382,N_2888,N_2447);
xnor U3383 (N_3383,N_2979,N_2092);
nand U3384 (N_3384,N_2742,N_2755);
nand U3385 (N_3385,N_2792,N_2102);
or U3386 (N_3386,N_2459,N_2153);
nor U3387 (N_3387,N_2586,N_2599);
and U3388 (N_3388,N_2812,N_2199);
nand U3389 (N_3389,N_2363,N_2055);
nor U3390 (N_3390,N_2088,N_2659);
or U3391 (N_3391,N_2876,N_2416);
and U3392 (N_3392,N_2384,N_2686);
and U3393 (N_3393,N_2432,N_2292);
and U3394 (N_3394,N_2839,N_2343);
and U3395 (N_3395,N_2239,N_2627);
nor U3396 (N_3396,N_2498,N_2950);
and U3397 (N_3397,N_2137,N_2830);
and U3398 (N_3398,N_2724,N_2768);
nand U3399 (N_3399,N_2308,N_2054);
or U3400 (N_3400,N_2392,N_2156);
nand U3401 (N_3401,N_2527,N_2202);
or U3402 (N_3402,N_2034,N_2250);
nor U3403 (N_3403,N_2412,N_2085);
nor U3404 (N_3404,N_2106,N_2107);
nand U3405 (N_3405,N_2763,N_2794);
or U3406 (N_3406,N_2270,N_2556);
or U3407 (N_3407,N_2396,N_2469);
or U3408 (N_3408,N_2248,N_2219);
and U3409 (N_3409,N_2282,N_2040);
and U3410 (N_3410,N_2537,N_2465);
and U3411 (N_3411,N_2829,N_2509);
and U3412 (N_3412,N_2208,N_2689);
or U3413 (N_3413,N_2455,N_2615);
nand U3414 (N_3414,N_2429,N_2355);
and U3415 (N_3415,N_2011,N_2192);
or U3416 (N_3416,N_2209,N_2388);
and U3417 (N_3417,N_2705,N_2142);
and U3418 (N_3418,N_2291,N_2353);
and U3419 (N_3419,N_2886,N_2220);
xnor U3420 (N_3420,N_2807,N_2136);
nor U3421 (N_3421,N_2485,N_2430);
and U3422 (N_3422,N_2719,N_2058);
xor U3423 (N_3423,N_2393,N_2570);
or U3424 (N_3424,N_2771,N_2288);
nand U3425 (N_3425,N_2067,N_2820);
nand U3426 (N_3426,N_2630,N_2555);
or U3427 (N_3427,N_2249,N_2802);
or U3428 (N_3428,N_2956,N_2953);
nand U3429 (N_3429,N_2141,N_2731);
nor U3430 (N_3430,N_2865,N_2066);
and U3431 (N_3431,N_2382,N_2821);
nor U3432 (N_3432,N_2795,N_2701);
nor U3433 (N_3433,N_2575,N_2766);
nor U3434 (N_3434,N_2307,N_2134);
nor U3435 (N_3435,N_2869,N_2230);
nand U3436 (N_3436,N_2912,N_2530);
and U3437 (N_3437,N_2433,N_2175);
nand U3438 (N_3438,N_2317,N_2168);
or U3439 (N_3439,N_2007,N_2728);
nor U3440 (N_3440,N_2894,N_2077);
nor U3441 (N_3441,N_2146,N_2068);
nor U3442 (N_3442,N_2178,N_2658);
and U3443 (N_3443,N_2576,N_2398);
and U3444 (N_3444,N_2769,N_2732);
nor U3445 (N_3445,N_2662,N_2568);
nand U3446 (N_3446,N_2478,N_2224);
nor U3447 (N_3447,N_2161,N_2052);
nand U3448 (N_3448,N_2808,N_2225);
or U3449 (N_3449,N_2313,N_2679);
or U3450 (N_3450,N_2713,N_2626);
nor U3451 (N_3451,N_2520,N_2639);
nor U3452 (N_3452,N_2461,N_2369);
nor U3453 (N_3453,N_2966,N_2312);
nand U3454 (N_3454,N_2752,N_2723);
nor U3455 (N_3455,N_2030,N_2127);
or U3456 (N_3456,N_2968,N_2943);
or U3457 (N_3457,N_2415,N_2174);
or U3458 (N_3458,N_2765,N_2492);
nor U3459 (N_3459,N_2907,N_2335);
or U3460 (N_3460,N_2000,N_2406);
or U3461 (N_3461,N_2170,N_2623);
and U3462 (N_3462,N_2084,N_2116);
nand U3463 (N_3463,N_2345,N_2227);
nand U3464 (N_3464,N_2551,N_2647);
nor U3465 (N_3465,N_2206,N_2234);
nor U3466 (N_3466,N_2512,N_2238);
and U3467 (N_3467,N_2676,N_2251);
nor U3468 (N_3468,N_2330,N_2559);
nand U3469 (N_3469,N_2744,N_2426);
nand U3470 (N_3470,N_2629,N_2324);
nand U3471 (N_3471,N_2177,N_2041);
and U3472 (N_3472,N_2504,N_2323);
nor U3473 (N_3473,N_2910,N_2076);
and U3474 (N_3474,N_2846,N_2563);
or U3475 (N_3475,N_2797,N_2321);
and U3476 (N_3476,N_2903,N_2867);
or U3477 (N_3477,N_2480,N_2687);
and U3478 (N_3478,N_2265,N_2010);
nor U3479 (N_3479,N_2971,N_2531);
and U3480 (N_3480,N_2565,N_2574);
and U3481 (N_3481,N_2824,N_2057);
nand U3482 (N_3482,N_2319,N_2800);
and U3483 (N_3483,N_2646,N_2358);
or U3484 (N_3484,N_2099,N_2014);
nor U3485 (N_3485,N_2042,N_2897);
nor U3486 (N_3486,N_2861,N_2222);
nor U3487 (N_3487,N_2481,N_2881);
nor U3488 (N_3488,N_2150,N_2813);
or U3489 (N_3489,N_2671,N_2511);
or U3490 (N_3490,N_2748,N_2460);
and U3491 (N_3491,N_2325,N_2435);
nor U3492 (N_3492,N_2163,N_2987);
nand U3493 (N_3493,N_2928,N_2761);
and U3494 (N_3494,N_2375,N_2311);
and U3495 (N_3495,N_2958,N_2022);
or U3496 (N_3496,N_2727,N_2298);
nand U3497 (N_3497,N_2691,N_2302);
or U3498 (N_3498,N_2838,N_2804);
and U3499 (N_3499,N_2871,N_2652);
nand U3500 (N_3500,N_2858,N_2315);
nor U3501 (N_3501,N_2199,N_2587);
or U3502 (N_3502,N_2996,N_2695);
nand U3503 (N_3503,N_2170,N_2125);
or U3504 (N_3504,N_2189,N_2240);
nor U3505 (N_3505,N_2764,N_2999);
and U3506 (N_3506,N_2046,N_2030);
nand U3507 (N_3507,N_2996,N_2556);
xnor U3508 (N_3508,N_2168,N_2380);
nor U3509 (N_3509,N_2636,N_2483);
nand U3510 (N_3510,N_2373,N_2302);
nand U3511 (N_3511,N_2435,N_2491);
nand U3512 (N_3512,N_2593,N_2748);
or U3513 (N_3513,N_2796,N_2736);
xor U3514 (N_3514,N_2145,N_2527);
or U3515 (N_3515,N_2161,N_2358);
nor U3516 (N_3516,N_2659,N_2003);
nand U3517 (N_3517,N_2687,N_2725);
or U3518 (N_3518,N_2496,N_2947);
or U3519 (N_3519,N_2276,N_2791);
or U3520 (N_3520,N_2573,N_2747);
nand U3521 (N_3521,N_2402,N_2134);
and U3522 (N_3522,N_2954,N_2093);
and U3523 (N_3523,N_2438,N_2817);
or U3524 (N_3524,N_2545,N_2801);
nor U3525 (N_3525,N_2563,N_2295);
nand U3526 (N_3526,N_2409,N_2381);
and U3527 (N_3527,N_2515,N_2260);
and U3528 (N_3528,N_2611,N_2514);
and U3529 (N_3529,N_2724,N_2003);
or U3530 (N_3530,N_2573,N_2252);
and U3531 (N_3531,N_2872,N_2149);
or U3532 (N_3532,N_2894,N_2263);
nand U3533 (N_3533,N_2185,N_2695);
nand U3534 (N_3534,N_2401,N_2766);
nand U3535 (N_3535,N_2937,N_2027);
nand U3536 (N_3536,N_2840,N_2906);
nand U3537 (N_3537,N_2355,N_2845);
nor U3538 (N_3538,N_2683,N_2547);
or U3539 (N_3539,N_2068,N_2665);
nor U3540 (N_3540,N_2851,N_2272);
nand U3541 (N_3541,N_2294,N_2638);
and U3542 (N_3542,N_2082,N_2132);
and U3543 (N_3543,N_2798,N_2007);
or U3544 (N_3544,N_2869,N_2830);
nor U3545 (N_3545,N_2805,N_2653);
or U3546 (N_3546,N_2215,N_2417);
nor U3547 (N_3547,N_2181,N_2189);
or U3548 (N_3548,N_2630,N_2418);
and U3549 (N_3549,N_2499,N_2891);
and U3550 (N_3550,N_2676,N_2057);
xor U3551 (N_3551,N_2417,N_2336);
nor U3552 (N_3552,N_2326,N_2979);
and U3553 (N_3553,N_2251,N_2308);
nand U3554 (N_3554,N_2484,N_2695);
nor U3555 (N_3555,N_2132,N_2490);
nand U3556 (N_3556,N_2278,N_2759);
and U3557 (N_3557,N_2719,N_2993);
or U3558 (N_3558,N_2407,N_2378);
or U3559 (N_3559,N_2283,N_2232);
nor U3560 (N_3560,N_2903,N_2007);
and U3561 (N_3561,N_2037,N_2368);
and U3562 (N_3562,N_2470,N_2422);
and U3563 (N_3563,N_2654,N_2416);
or U3564 (N_3564,N_2287,N_2015);
or U3565 (N_3565,N_2350,N_2487);
or U3566 (N_3566,N_2150,N_2241);
nand U3567 (N_3567,N_2672,N_2454);
nor U3568 (N_3568,N_2317,N_2701);
and U3569 (N_3569,N_2712,N_2587);
nor U3570 (N_3570,N_2645,N_2711);
and U3571 (N_3571,N_2028,N_2602);
and U3572 (N_3572,N_2301,N_2282);
nor U3573 (N_3573,N_2737,N_2330);
nor U3574 (N_3574,N_2939,N_2100);
or U3575 (N_3575,N_2866,N_2562);
and U3576 (N_3576,N_2373,N_2308);
or U3577 (N_3577,N_2133,N_2614);
nor U3578 (N_3578,N_2672,N_2391);
or U3579 (N_3579,N_2452,N_2157);
nor U3580 (N_3580,N_2185,N_2154);
or U3581 (N_3581,N_2203,N_2711);
and U3582 (N_3582,N_2100,N_2917);
or U3583 (N_3583,N_2996,N_2374);
and U3584 (N_3584,N_2367,N_2976);
or U3585 (N_3585,N_2357,N_2493);
xor U3586 (N_3586,N_2778,N_2802);
and U3587 (N_3587,N_2479,N_2696);
or U3588 (N_3588,N_2583,N_2159);
nand U3589 (N_3589,N_2304,N_2739);
and U3590 (N_3590,N_2364,N_2374);
nor U3591 (N_3591,N_2354,N_2515);
or U3592 (N_3592,N_2066,N_2896);
nand U3593 (N_3593,N_2105,N_2367);
nor U3594 (N_3594,N_2328,N_2900);
and U3595 (N_3595,N_2222,N_2492);
or U3596 (N_3596,N_2945,N_2425);
nand U3597 (N_3597,N_2986,N_2515);
nand U3598 (N_3598,N_2337,N_2416);
or U3599 (N_3599,N_2445,N_2158);
and U3600 (N_3600,N_2604,N_2879);
and U3601 (N_3601,N_2061,N_2442);
nand U3602 (N_3602,N_2295,N_2289);
nor U3603 (N_3603,N_2955,N_2136);
or U3604 (N_3604,N_2818,N_2345);
nor U3605 (N_3605,N_2822,N_2964);
and U3606 (N_3606,N_2936,N_2671);
xnor U3607 (N_3607,N_2992,N_2335);
nor U3608 (N_3608,N_2187,N_2765);
nor U3609 (N_3609,N_2320,N_2817);
nand U3610 (N_3610,N_2911,N_2003);
or U3611 (N_3611,N_2325,N_2251);
nor U3612 (N_3612,N_2440,N_2133);
and U3613 (N_3613,N_2960,N_2383);
and U3614 (N_3614,N_2638,N_2750);
or U3615 (N_3615,N_2300,N_2048);
nor U3616 (N_3616,N_2344,N_2112);
or U3617 (N_3617,N_2837,N_2393);
nor U3618 (N_3618,N_2467,N_2010);
nand U3619 (N_3619,N_2408,N_2610);
and U3620 (N_3620,N_2572,N_2397);
or U3621 (N_3621,N_2919,N_2569);
or U3622 (N_3622,N_2031,N_2134);
nor U3623 (N_3623,N_2242,N_2982);
nand U3624 (N_3624,N_2366,N_2910);
nand U3625 (N_3625,N_2797,N_2012);
or U3626 (N_3626,N_2512,N_2421);
nor U3627 (N_3627,N_2207,N_2764);
nand U3628 (N_3628,N_2542,N_2274);
nor U3629 (N_3629,N_2209,N_2706);
and U3630 (N_3630,N_2134,N_2802);
and U3631 (N_3631,N_2715,N_2579);
nor U3632 (N_3632,N_2402,N_2374);
nand U3633 (N_3633,N_2695,N_2626);
nand U3634 (N_3634,N_2876,N_2408);
and U3635 (N_3635,N_2120,N_2917);
nor U3636 (N_3636,N_2027,N_2314);
nand U3637 (N_3637,N_2550,N_2690);
and U3638 (N_3638,N_2990,N_2586);
and U3639 (N_3639,N_2810,N_2711);
nand U3640 (N_3640,N_2650,N_2688);
and U3641 (N_3641,N_2068,N_2142);
nor U3642 (N_3642,N_2118,N_2821);
and U3643 (N_3643,N_2205,N_2093);
or U3644 (N_3644,N_2428,N_2878);
nand U3645 (N_3645,N_2189,N_2885);
nor U3646 (N_3646,N_2360,N_2819);
nand U3647 (N_3647,N_2107,N_2156);
nor U3648 (N_3648,N_2726,N_2893);
nor U3649 (N_3649,N_2458,N_2325);
and U3650 (N_3650,N_2365,N_2075);
and U3651 (N_3651,N_2287,N_2099);
nor U3652 (N_3652,N_2227,N_2771);
or U3653 (N_3653,N_2789,N_2043);
nand U3654 (N_3654,N_2602,N_2837);
or U3655 (N_3655,N_2535,N_2408);
nor U3656 (N_3656,N_2278,N_2358);
nand U3657 (N_3657,N_2163,N_2240);
xor U3658 (N_3658,N_2956,N_2458);
and U3659 (N_3659,N_2671,N_2309);
or U3660 (N_3660,N_2722,N_2397);
and U3661 (N_3661,N_2091,N_2541);
and U3662 (N_3662,N_2892,N_2755);
nor U3663 (N_3663,N_2962,N_2223);
or U3664 (N_3664,N_2268,N_2630);
or U3665 (N_3665,N_2204,N_2111);
or U3666 (N_3666,N_2021,N_2324);
nor U3667 (N_3667,N_2516,N_2072);
nor U3668 (N_3668,N_2209,N_2905);
xor U3669 (N_3669,N_2621,N_2486);
or U3670 (N_3670,N_2568,N_2475);
and U3671 (N_3671,N_2205,N_2749);
and U3672 (N_3672,N_2720,N_2505);
nor U3673 (N_3673,N_2723,N_2961);
nor U3674 (N_3674,N_2271,N_2692);
nor U3675 (N_3675,N_2639,N_2277);
nand U3676 (N_3676,N_2609,N_2348);
nor U3677 (N_3677,N_2017,N_2674);
and U3678 (N_3678,N_2155,N_2502);
and U3679 (N_3679,N_2213,N_2998);
and U3680 (N_3680,N_2327,N_2044);
nor U3681 (N_3681,N_2290,N_2784);
and U3682 (N_3682,N_2106,N_2363);
or U3683 (N_3683,N_2457,N_2356);
nor U3684 (N_3684,N_2792,N_2244);
nor U3685 (N_3685,N_2388,N_2843);
nand U3686 (N_3686,N_2018,N_2133);
and U3687 (N_3687,N_2257,N_2484);
nor U3688 (N_3688,N_2745,N_2375);
nand U3689 (N_3689,N_2973,N_2767);
nor U3690 (N_3690,N_2843,N_2287);
nor U3691 (N_3691,N_2640,N_2651);
nand U3692 (N_3692,N_2872,N_2732);
nor U3693 (N_3693,N_2409,N_2454);
nand U3694 (N_3694,N_2639,N_2986);
or U3695 (N_3695,N_2219,N_2978);
nor U3696 (N_3696,N_2343,N_2873);
and U3697 (N_3697,N_2053,N_2054);
nor U3698 (N_3698,N_2737,N_2025);
or U3699 (N_3699,N_2967,N_2248);
nand U3700 (N_3700,N_2979,N_2635);
nand U3701 (N_3701,N_2727,N_2974);
xnor U3702 (N_3702,N_2017,N_2185);
or U3703 (N_3703,N_2506,N_2275);
or U3704 (N_3704,N_2351,N_2157);
or U3705 (N_3705,N_2718,N_2179);
or U3706 (N_3706,N_2845,N_2689);
or U3707 (N_3707,N_2737,N_2881);
and U3708 (N_3708,N_2707,N_2905);
and U3709 (N_3709,N_2828,N_2005);
nand U3710 (N_3710,N_2257,N_2681);
and U3711 (N_3711,N_2172,N_2133);
and U3712 (N_3712,N_2113,N_2001);
and U3713 (N_3713,N_2857,N_2632);
nor U3714 (N_3714,N_2046,N_2941);
or U3715 (N_3715,N_2142,N_2642);
and U3716 (N_3716,N_2933,N_2743);
nor U3717 (N_3717,N_2945,N_2964);
nor U3718 (N_3718,N_2675,N_2524);
xnor U3719 (N_3719,N_2282,N_2948);
nor U3720 (N_3720,N_2898,N_2630);
or U3721 (N_3721,N_2003,N_2767);
and U3722 (N_3722,N_2014,N_2498);
or U3723 (N_3723,N_2255,N_2717);
nor U3724 (N_3724,N_2941,N_2171);
nor U3725 (N_3725,N_2173,N_2032);
or U3726 (N_3726,N_2408,N_2683);
nand U3727 (N_3727,N_2386,N_2042);
or U3728 (N_3728,N_2730,N_2526);
nand U3729 (N_3729,N_2430,N_2811);
or U3730 (N_3730,N_2422,N_2030);
nand U3731 (N_3731,N_2681,N_2935);
nor U3732 (N_3732,N_2697,N_2541);
or U3733 (N_3733,N_2568,N_2873);
or U3734 (N_3734,N_2574,N_2757);
nor U3735 (N_3735,N_2535,N_2949);
and U3736 (N_3736,N_2599,N_2138);
nor U3737 (N_3737,N_2440,N_2764);
and U3738 (N_3738,N_2237,N_2044);
nand U3739 (N_3739,N_2686,N_2615);
nand U3740 (N_3740,N_2810,N_2302);
and U3741 (N_3741,N_2101,N_2904);
or U3742 (N_3742,N_2264,N_2532);
nand U3743 (N_3743,N_2007,N_2649);
or U3744 (N_3744,N_2525,N_2042);
nand U3745 (N_3745,N_2242,N_2792);
nor U3746 (N_3746,N_2144,N_2182);
and U3747 (N_3747,N_2053,N_2761);
and U3748 (N_3748,N_2351,N_2194);
and U3749 (N_3749,N_2041,N_2479);
and U3750 (N_3750,N_2438,N_2395);
or U3751 (N_3751,N_2555,N_2713);
nor U3752 (N_3752,N_2654,N_2681);
nor U3753 (N_3753,N_2131,N_2791);
or U3754 (N_3754,N_2991,N_2164);
and U3755 (N_3755,N_2110,N_2511);
nor U3756 (N_3756,N_2534,N_2495);
nor U3757 (N_3757,N_2260,N_2533);
nor U3758 (N_3758,N_2958,N_2162);
nor U3759 (N_3759,N_2244,N_2460);
nand U3760 (N_3760,N_2753,N_2740);
xnor U3761 (N_3761,N_2079,N_2855);
nor U3762 (N_3762,N_2760,N_2243);
nor U3763 (N_3763,N_2456,N_2261);
nor U3764 (N_3764,N_2213,N_2926);
nor U3765 (N_3765,N_2438,N_2974);
and U3766 (N_3766,N_2694,N_2843);
and U3767 (N_3767,N_2363,N_2309);
or U3768 (N_3768,N_2400,N_2659);
xor U3769 (N_3769,N_2233,N_2603);
or U3770 (N_3770,N_2138,N_2330);
and U3771 (N_3771,N_2886,N_2723);
nor U3772 (N_3772,N_2871,N_2336);
or U3773 (N_3773,N_2887,N_2114);
or U3774 (N_3774,N_2241,N_2456);
nand U3775 (N_3775,N_2186,N_2699);
and U3776 (N_3776,N_2000,N_2207);
nand U3777 (N_3777,N_2232,N_2569);
or U3778 (N_3778,N_2579,N_2742);
xor U3779 (N_3779,N_2258,N_2686);
or U3780 (N_3780,N_2038,N_2325);
and U3781 (N_3781,N_2013,N_2413);
nand U3782 (N_3782,N_2986,N_2243);
and U3783 (N_3783,N_2522,N_2851);
nand U3784 (N_3784,N_2699,N_2194);
or U3785 (N_3785,N_2707,N_2429);
or U3786 (N_3786,N_2684,N_2792);
nor U3787 (N_3787,N_2887,N_2594);
nor U3788 (N_3788,N_2332,N_2295);
or U3789 (N_3789,N_2787,N_2960);
nor U3790 (N_3790,N_2335,N_2785);
and U3791 (N_3791,N_2036,N_2493);
or U3792 (N_3792,N_2914,N_2540);
nor U3793 (N_3793,N_2630,N_2746);
and U3794 (N_3794,N_2919,N_2430);
or U3795 (N_3795,N_2034,N_2591);
and U3796 (N_3796,N_2593,N_2979);
and U3797 (N_3797,N_2966,N_2631);
or U3798 (N_3798,N_2239,N_2341);
nor U3799 (N_3799,N_2578,N_2776);
or U3800 (N_3800,N_2215,N_2605);
nor U3801 (N_3801,N_2289,N_2524);
and U3802 (N_3802,N_2110,N_2349);
nand U3803 (N_3803,N_2305,N_2071);
or U3804 (N_3804,N_2476,N_2410);
and U3805 (N_3805,N_2749,N_2936);
nor U3806 (N_3806,N_2609,N_2121);
and U3807 (N_3807,N_2058,N_2891);
nor U3808 (N_3808,N_2227,N_2789);
and U3809 (N_3809,N_2151,N_2983);
and U3810 (N_3810,N_2538,N_2955);
nor U3811 (N_3811,N_2950,N_2336);
nor U3812 (N_3812,N_2980,N_2047);
xor U3813 (N_3813,N_2684,N_2723);
nor U3814 (N_3814,N_2856,N_2027);
xor U3815 (N_3815,N_2192,N_2937);
nand U3816 (N_3816,N_2981,N_2284);
nor U3817 (N_3817,N_2622,N_2342);
nand U3818 (N_3818,N_2427,N_2552);
nand U3819 (N_3819,N_2465,N_2435);
nor U3820 (N_3820,N_2045,N_2704);
and U3821 (N_3821,N_2543,N_2089);
nand U3822 (N_3822,N_2055,N_2485);
and U3823 (N_3823,N_2870,N_2096);
and U3824 (N_3824,N_2663,N_2307);
or U3825 (N_3825,N_2528,N_2020);
nor U3826 (N_3826,N_2121,N_2388);
nand U3827 (N_3827,N_2450,N_2232);
and U3828 (N_3828,N_2397,N_2729);
nand U3829 (N_3829,N_2637,N_2609);
and U3830 (N_3830,N_2679,N_2548);
and U3831 (N_3831,N_2601,N_2004);
and U3832 (N_3832,N_2782,N_2385);
nor U3833 (N_3833,N_2729,N_2975);
and U3834 (N_3834,N_2224,N_2688);
xor U3835 (N_3835,N_2286,N_2504);
nor U3836 (N_3836,N_2721,N_2991);
or U3837 (N_3837,N_2977,N_2209);
nand U3838 (N_3838,N_2310,N_2376);
nand U3839 (N_3839,N_2368,N_2789);
nor U3840 (N_3840,N_2831,N_2042);
or U3841 (N_3841,N_2311,N_2229);
nand U3842 (N_3842,N_2274,N_2449);
nand U3843 (N_3843,N_2782,N_2017);
and U3844 (N_3844,N_2734,N_2078);
nand U3845 (N_3845,N_2904,N_2937);
nor U3846 (N_3846,N_2981,N_2074);
or U3847 (N_3847,N_2980,N_2763);
or U3848 (N_3848,N_2664,N_2061);
and U3849 (N_3849,N_2890,N_2454);
or U3850 (N_3850,N_2842,N_2330);
and U3851 (N_3851,N_2767,N_2883);
or U3852 (N_3852,N_2078,N_2433);
and U3853 (N_3853,N_2897,N_2261);
xnor U3854 (N_3854,N_2633,N_2018);
nand U3855 (N_3855,N_2886,N_2787);
or U3856 (N_3856,N_2888,N_2303);
xor U3857 (N_3857,N_2951,N_2909);
xor U3858 (N_3858,N_2898,N_2462);
and U3859 (N_3859,N_2801,N_2756);
nor U3860 (N_3860,N_2547,N_2687);
and U3861 (N_3861,N_2055,N_2626);
or U3862 (N_3862,N_2486,N_2666);
and U3863 (N_3863,N_2097,N_2617);
or U3864 (N_3864,N_2403,N_2491);
or U3865 (N_3865,N_2700,N_2733);
or U3866 (N_3866,N_2155,N_2284);
nand U3867 (N_3867,N_2435,N_2920);
or U3868 (N_3868,N_2876,N_2607);
and U3869 (N_3869,N_2125,N_2888);
nand U3870 (N_3870,N_2390,N_2482);
or U3871 (N_3871,N_2108,N_2357);
nor U3872 (N_3872,N_2228,N_2212);
nand U3873 (N_3873,N_2670,N_2080);
nor U3874 (N_3874,N_2731,N_2425);
or U3875 (N_3875,N_2906,N_2690);
nor U3876 (N_3876,N_2501,N_2772);
nor U3877 (N_3877,N_2030,N_2344);
xor U3878 (N_3878,N_2944,N_2000);
or U3879 (N_3879,N_2627,N_2461);
nor U3880 (N_3880,N_2172,N_2313);
or U3881 (N_3881,N_2695,N_2147);
nor U3882 (N_3882,N_2412,N_2148);
or U3883 (N_3883,N_2602,N_2758);
and U3884 (N_3884,N_2244,N_2968);
nor U3885 (N_3885,N_2700,N_2616);
nand U3886 (N_3886,N_2306,N_2687);
nor U3887 (N_3887,N_2646,N_2709);
or U3888 (N_3888,N_2486,N_2780);
nand U3889 (N_3889,N_2735,N_2670);
nor U3890 (N_3890,N_2866,N_2178);
xor U3891 (N_3891,N_2194,N_2204);
nor U3892 (N_3892,N_2053,N_2516);
and U3893 (N_3893,N_2095,N_2366);
or U3894 (N_3894,N_2968,N_2069);
and U3895 (N_3895,N_2739,N_2931);
or U3896 (N_3896,N_2331,N_2235);
and U3897 (N_3897,N_2184,N_2023);
nor U3898 (N_3898,N_2825,N_2032);
and U3899 (N_3899,N_2710,N_2793);
nand U3900 (N_3900,N_2796,N_2717);
or U3901 (N_3901,N_2603,N_2802);
and U3902 (N_3902,N_2639,N_2040);
nor U3903 (N_3903,N_2254,N_2064);
nor U3904 (N_3904,N_2559,N_2947);
and U3905 (N_3905,N_2436,N_2629);
nor U3906 (N_3906,N_2986,N_2766);
and U3907 (N_3907,N_2230,N_2003);
and U3908 (N_3908,N_2761,N_2158);
xor U3909 (N_3909,N_2128,N_2473);
or U3910 (N_3910,N_2795,N_2956);
or U3911 (N_3911,N_2370,N_2891);
and U3912 (N_3912,N_2782,N_2812);
nand U3913 (N_3913,N_2980,N_2020);
and U3914 (N_3914,N_2021,N_2988);
nand U3915 (N_3915,N_2875,N_2582);
nor U3916 (N_3916,N_2208,N_2787);
nand U3917 (N_3917,N_2811,N_2813);
or U3918 (N_3918,N_2274,N_2083);
or U3919 (N_3919,N_2723,N_2419);
nand U3920 (N_3920,N_2130,N_2786);
or U3921 (N_3921,N_2118,N_2043);
or U3922 (N_3922,N_2089,N_2574);
or U3923 (N_3923,N_2140,N_2202);
and U3924 (N_3924,N_2150,N_2066);
and U3925 (N_3925,N_2528,N_2687);
and U3926 (N_3926,N_2672,N_2605);
or U3927 (N_3927,N_2251,N_2039);
and U3928 (N_3928,N_2740,N_2207);
and U3929 (N_3929,N_2907,N_2231);
or U3930 (N_3930,N_2368,N_2815);
or U3931 (N_3931,N_2211,N_2777);
or U3932 (N_3932,N_2808,N_2993);
and U3933 (N_3933,N_2020,N_2312);
nand U3934 (N_3934,N_2999,N_2321);
or U3935 (N_3935,N_2850,N_2136);
nand U3936 (N_3936,N_2557,N_2689);
nor U3937 (N_3937,N_2213,N_2294);
nand U3938 (N_3938,N_2631,N_2202);
or U3939 (N_3939,N_2627,N_2622);
or U3940 (N_3940,N_2488,N_2427);
and U3941 (N_3941,N_2006,N_2028);
nand U3942 (N_3942,N_2893,N_2892);
or U3943 (N_3943,N_2249,N_2190);
nand U3944 (N_3944,N_2757,N_2463);
nand U3945 (N_3945,N_2634,N_2260);
and U3946 (N_3946,N_2444,N_2217);
and U3947 (N_3947,N_2130,N_2633);
or U3948 (N_3948,N_2661,N_2607);
nor U3949 (N_3949,N_2356,N_2053);
or U3950 (N_3950,N_2045,N_2649);
nand U3951 (N_3951,N_2786,N_2354);
and U3952 (N_3952,N_2030,N_2896);
nand U3953 (N_3953,N_2211,N_2497);
nand U3954 (N_3954,N_2811,N_2070);
nand U3955 (N_3955,N_2486,N_2479);
or U3956 (N_3956,N_2279,N_2171);
nand U3957 (N_3957,N_2382,N_2422);
or U3958 (N_3958,N_2145,N_2333);
nor U3959 (N_3959,N_2728,N_2739);
nor U3960 (N_3960,N_2914,N_2690);
nor U3961 (N_3961,N_2091,N_2479);
nand U3962 (N_3962,N_2588,N_2232);
or U3963 (N_3963,N_2442,N_2165);
or U3964 (N_3964,N_2173,N_2471);
nor U3965 (N_3965,N_2720,N_2365);
and U3966 (N_3966,N_2988,N_2469);
nor U3967 (N_3967,N_2989,N_2139);
nand U3968 (N_3968,N_2069,N_2785);
nand U3969 (N_3969,N_2939,N_2197);
nor U3970 (N_3970,N_2361,N_2260);
and U3971 (N_3971,N_2340,N_2910);
nor U3972 (N_3972,N_2172,N_2946);
and U3973 (N_3973,N_2765,N_2907);
nand U3974 (N_3974,N_2018,N_2311);
nor U3975 (N_3975,N_2861,N_2567);
nand U3976 (N_3976,N_2305,N_2990);
nor U3977 (N_3977,N_2640,N_2451);
or U3978 (N_3978,N_2579,N_2706);
or U3979 (N_3979,N_2259,N_2401);
and U3980 (N_3980,N_2923,N_2033);
nand U3981 (N_3981,N_2846,N_2866);
nand U3982 (N_3982,N_2501,N_2872);
and U3983 (N_3983,N_2774,N_2533);
nand U3984 (N_3984,N_2206,N_2886);
or U3985 (N_3985,N_2233,N_2381);
or U3986 (N_3986,N_2435,N_2713);
and U3987 (N_3987,N_2250,N_2211);
or U3988 (N_3988,N_2686,N_2557);
and U3989 (N_3989,N_2929,N_2398);
nand U3990 (N_3990,N_2002,N_2307);
nand U3991 (N_3991,N_2076,N_2108);
nand U3992 (N_3992,N_2809,N_2423);
nor U3993 (N_3993,N_2054,N_2302);
nor U3994 (N_3994,N_2740,N_2847);
and U3995 (N_3995,N_2447,N_2166);
nand U3996 (N_3996,N_2683,N_2906);
nor U3997 (N_3997,N_2351,N_2437);
nand U3998 (N_3998,N_2326,N_2685);
and U3999 (N_3999,N_2164,N_2535);
nor U4000 (N_4000,N_3041,N_3369);
and U4001 (N_4001,N_3395,N_3518);
nor U4002 (N_4002,N_3329,N_3895);
nor U4003 (N_4003,N_3229,N_3287);
and U4004 (N_4004,N_3015,N_3218);
nand U4005 (N_4005,N_3623,N_3647);
or U4006 (N_4006,N_3602,N_3980);
nor U4007 (N_4007,N_3452,N_3264);
or U4008 (N_4008,N_3413,N_3364);
and U4009 (N_4009,N_3613,N_3976);
nand U4010 (N_4010,N_3078,N_3658);
or U4011 (N_4011,N_3222,N_3012);
and U4012 (N_4012,N_3554,N_3266);
and U4013 (N_4013,N_3180,N_3248);
and U4014 (N_4014,N_3439,N_3774);
and U4015 (N_4015,N_3391,N_3002);
nor U4016 (N_4016,N_3142,N_3922);
and U4017 (N_4017,N_3254,N_3117);
xnor U4018 (N_4018,N_3867,N_3914);
nand U4019 (N_4019,N_3133,N_3838);
nor U4020 (N_4020,N_3455,N_3910);
nor U4021 (N_4021,N_3631,N_3392);
or U4022 (N_4022,N_3597,N_3539);
or U4023 (N_4023,N_3938,N_3058);
nand U4024 (N_4024,N_3127,N_3555);
and U4025 (N_4025,N_3508,N_3782);
and U4026 (N_4026,N_3790,N_3726);
xor U4027 (N_4027,N_3698,N_3188);
nand U4028 (N_4028,N_3183,N_3501);
nor U4029 (N_4029,N_3320,N_3909);
or U4030 (N_4030,N_3925,N_3505);
or U4031 (N_4031,N_3315,N_3869);
nand U4032 (N_4032,N_3594,N_3311);
nand U4033 (N_4033,N_3966,N_3628);
nand U4034 (N_4034,N_3839,N_3020);
or U4035 (N_4035,N_3178,N_3848);
nand U4036 (N_4036,N_3036,N_3171);
nor U4037 (N_4037,N_3521,N_3361);
nor U4038 (N_4038,N_3054,N_3519);
and U4039 (N_4039,N_3177,N_3550);
xor U4040 (N_4040,N_3108,N_3485);
and U4041 (N_4041,N_3932,N_3879);
and U4042 (N_4042,N_3948,N_3131);
nand U4043 (N_4043,N_3414,N_3350);
nor U4044 (N_4044,N_3394,N_3269);
nor U4045 (N_4045,N_3301,N_3008);
and U4046 (N_4046,N_3163,N_3048);
and U4047 (N_4047,N_3368,N_3856);
nand U4048 (N_4048,N_3273,N_3304);
and U4049 (N_4049,N_3622,N_3010);
nor U4050 (N_4050,N_3104,N_3982);
nor U4051 (N_4051,N_3764,N_3215);
nand U4052 (N_4052,N_3242,N_3950);
nand U4053 (N_4053,N_3890,N_3372);
or U4054 (N_4054,N_3478,N_3491);
or U4055 (N_4055,N_3611,N_3748);
and U4056 (N_4056,N_3546,N_3201);
nor U4057 (N_4057,N_3927,N_3003);
and U4058 (N_4058,N_3992,N_3476);
xnor U4059 (N_4059,N_3051,N_3088);
nand U4060 (N_4060,N_3538,N_3044);
nor U4061 (N_4061,N_3668,N_3448);
and U4062 (N_4062,N_3706,N_3154);
and U4063 (N_4063,N_3707,N_3715);
nor U4064 (N_4064,N_3575,N_3302);
nor U4065 (N_4065,N_3007,N_3461);
or U4066 (N_4066,N_3649,N_3576);
nand U4067 (N_4067,N_3028,N_3401);
and U4068 (N_4068,N_3626,N_3703);
and U4069 (N_4069,N_3449,N_3629);
or U4070 (N_4070,N_3990,N_3701);
nand U4071 (N_4071,N_3453,N_3947);
nor U4072 (N_4072,N_3757,N_3915);
or U4073 (N_4073,N_3667,N_3809);
or U4074 (N_4074,N_3637,N_3487);
or U4075 (N_4075,N_3525,N_3109);
and U4076 (N_4076,N_3836,N_3569);
nor U4077 (N_4077,N_3393,N_3591);
and U4078 (N_4078,N_3663,N_3244);
nand U4079 (N_4079,N_3191,N_3516);
nor U4080 (N_4080,N_3016,N_3013);
and U4081 (N_4081,N_3995,N_3573);
nand U4082 (N_4082,N_3110,N_3050);
nand U4083 (N_4083,N_3685,N_3887);
and U4084 (N_4084,N_3857,N_3405);
and U4085 (N_4085,N_3837,N_3428);
or U4086 (N_4086,N_3164,N_3549);
nand U4087 (N_4087,N_3733,N_3736);
nor U4088 (N_4088,N_3833,N_3319);
and U4089 (N_4089,N_3691,N_3831);
nand U4090 (N_4090,N_3195,N_3678);
nand U4091 (N_4091,N_3261,N_3105);
or U4092 (N_4092,N_3472,N_3283);
nor U4093 (N_4093,N_3256,N_3059);
xnor U4094 (N_4094,N_3113,N_3953);
and U4095 (N_4095,N_3221,N_3643);
xor U4096 (N_4096,N_3358,N_3464);
nor U4097 (N_4097,N_3324,N_3237);
nor U4098 (N_4098,N_3123,N_3926);
or U4099 (N_4099,N_3507,N_3719);
nand U4100 (N_4100,N_3822,N_3676);
or U4101 (N_4101,N_3761,N_3470);
and U4102 (N_4102,N_3297,N_3669);
and U4103 (N_4103,N_3704,N_3285);
and U4104 (N_4104,N_3801,N_3959);
xnor U4105 (N_4105,N_3721,N_3042);
xor U4106 (N_4106,N_3483,N_3718);
nor U4107 (N_4107,N_3270,N_3067);
nor U4108 (N_4108,N_3532,N_3427);
nand U4109 (N_4109,N_3381,N_3290);
nor U4110 (N_4110,N_3169,N_3492);
xor U4111 (N_4111,N_3101,N_3349);
and U4112 (N_4112,N_3182,N_3305);
or U4113 (N_4113,N_3714,N_3635);
nand U4114 (N_4114,N_3789,N_3754);
nor U4115 (N_4115,N_3534,N_3403);
nand U4116 (N_4116,N_3217,N_3001);
and U4117 (N_4117,N_3486,N_3328);
nor U4118 (N_4118,N_3321,N_3233);
and U4119 (N_4119,N_3374,N_3974);
nand U4120 (N_4120,N_3306,N_3642);
nor U4121 (N_4121,N_3477,N_3987);
and U4122 (N_4122,N_3230,N_3384);
xnor U4123 (N_4123,N_3093,N_3991);
nor U4124 (N_4124,N_3068,N_3547);
nor U4125 (N_4125,N_3825,N_3921);
nor U4126 (N_4126,N_3167,N_3806);
xnor U4127 (N_4127,N_3904,N_3312);
and U4128 (N_4128,N_3657,N_3097);
or U4129 (N_4129,N_3791,N_3160);
nand U4130 (N_4130,N_3387,N_3794);
nor U4131 (N_4131,N_3636,N_3697);
nand U4132 (N_4132,N_3901,N_3220);
and U4133 (N_4133,N_3677,N_3655);
or U4134 (N_4134,N_3348,N_3046);
nand U4135 (N_4135,N_3600,N_3119);
and U4136 (N_4136,N_3398,N_3713);
nand U4137 (N_4137,N_3265,N_3751);
nand U4138 (N_4138,N_3973,N_3968);
nand U4139 (N_4139,N_3551,N_3080);
nor U4140 (N_4140,N_3605,N_3560);
or U4141 (N_4141,N_3280,N_3434);
and U4142 (N_4142,N_3389,N_3040);
and U4143 (N_4143,N_3043,N_3871);
and U4144 (N_4144,N_3271,N_3337);
nor U4145 (N_4145,N_3943,N_3422);
nand U4146 (N_4146,N_3627,N_3423);
and U4147 (N_4147,N_3488,N_3380);
nand U4148 (N_4148,N_3116,N_3239);
nor U4149 (N_4149,N_3409,N_3883);
or U4150 (N_4150,N_3019,N_3122);
or U4151 (N_4151,N_3245,N_3137);
nand U4152 (N_4152,N_3162,N_3989);
and U4153 (N_4153,N_3797,N_3529);
nand U4154 (N_4154,N_3438,N_3303);
nand U4155 (N_4155,N_3499,N_3341);
nor U4156 (N_4156,N_3695,N_3888);
nor U4157 (N_4157,N_3330,N_3407);
nor U4158 (N_4158,N_3911,N_3143);
or U4159 (N_4159,N_3246,N_3559);
nand U4160 (N_4160,N_3670,N_3199);
and U4161 (N_4161,N_3360,N_3189);
nand U4162 (N_4162,N_3946,N_3225);
and U4163 (N_4163,N_3334,N_3524);
and U4164 (N_4164,N_3813,N_3777);
nor U4165 (N_4165,N_3125,N_3397);
nor U4166 (N_4166,N_3821,N_3996);
and U4167 (N_4167,N_3994,N_3325);
nand U4168 (N_4168,N_3808,N_3640);
and U4169 (N_4169,N_3200,N_3196);
nor U4170 (N_4170,N_3509,N_3582);
and U4171 (N_4171,N_3588,N_3294);
nor U4172 (N_4172,N_3309,N_3069);
and U4173 (N_4173,N_3855,N_3675);
and U4174 (N_4174,N_3033,N_3399);
and U4175 (N_4175,N_3608,N_3557);
nor U4176 (N_4176,N_3683,N_3236);
nor U4177 (N_4177,N_3029,N_3136);
nand U4178 (N_4178,N_3561,N_3999);
nor U4179 (N_4179,N_3945,N_3972);
nand U4180 (N_4180,N_3780,N_3638);
or U4181 (N_4181,N_3111,N_3853);
and U4182 (N_4182,N_3446,N_3209);
or U4183 (N_4183,N_3377,N_3314);
or U4184 (N_4184,N_3696,N_3268);
or U4185 (N_4185,N_3386,N_3146);
and U4186 (N_4186,N_3639,N_3089);
nor U4187 (N_4187,N_3076,N_3690);
or U4188 (N_4188,N_3956,N_3359);
and U4189 (N_4189,N_3371,N_3650);
or U4190 (N_4190,N_3772,N_3936);
and U4191 (N_4191,N_3846,N_3728);
or U4192 (N_4192,N_3278,N_3147);
or U4193 (N_4193,N_3206,N_3984);
nand U4194 (N_4194,N_3882,N_3144);
nand U4195 (N_4195,N_3277,N_3263);
nor U4196 (N_4196,N_3852,N_3416);
nand U4197 (N_4197,N_3625,N_3471);
or U4198 (N_4198,N_3458,N_3231);
or U4199 (N_4199,N_3238,N_3429);
or U4200 (N_4200,N_3584,N_3186);
and U4201 (N_4201,N_3812,N_3443);
and U4202 (N_4202,N_3563,N_3402);
and U4203 (N_4203,N_3845,N_3421);
nor U4204 (N_4204,N_3071,N_3396);
or U4205 (N_4205,N_3942,N_3725);
and U4206 (N_4206,N_3038,N_3975);
nand U4207 (N_4207,N_3954,N_3291);
or U4208 (N_4208,N_3024,N_3679);
nand U4209 (N_4209,N_3579,N_3988);
and U4210 (N_4210,N_3537,N_3343);
nand U4211 (N_4211,N_3333,N_3957);
nor U4212 (N_4212,N_3083,N_3566);
and U4213 (N_4213,N_3811,N_3522);
xnor U4214 (N_4214,N_3426,N_3366);
nand U4215 (N_4215,N_3656,N_3893);
or U4216 (N_4216,N_3260,N_3053);
nor U4217 (N_4217,N_3651,N_3553);
nand U4218 (N_4218,N_3830,N_3479);
and U4219 (N_4219,N_3878,N_3851);
nor U4220 (N_4220,N_3799,N_3150);
nand U4221 (N_4221,N_3198,N_3540);
xor U4222 (N_4222,N_3064,N_3410);
or U4223 (N_4223,N_3376,N_3276);
or U4224 (N_4224,N_3197,N_3899);
nor U4225 (N_4225,N_3565,N_3332);
nand U4226 (N_4226,N_3847,N_3571);
nor U4227 (N_4227,N_3194,N_3624);
and U4228 (N_4228,N_3346,N_3961);
nand U4229 (N_4229,N_3827,N_3365);
nor U4230 (N_4230,N_3710,N_3139);
and U4231 (N_4231,N_3930,N_3460);
or U4232 (N_4232,N_3755,N_3609);
nand U4233 (N_4233,N_3103,N_3440);
and U4234 (N_4234,N_3166,N_3114);
and U4235 (N_4235,N_3275,N_3603);
and U4236 (N_4236,N_3370,N_3606);
and U4237 (N_4237,N_3077,N_3468);
or U4238 (N_4238,N_3288,N_3327);
nand U4239 (N_4239,N_3298,N_3891);
nand U4240 (N_4240,N_3017,N_3185);
and U4241 (N_4241,N_3480,N_3339);
and U4242 (N_4242,N_3192,N_3572);
nand U4243 (N_4243,N_3310,N_3621);
nand U4244 (N_4244,N_3055,N_3255);
and U4245 (N_4245,N_3981,N_3589);
nor U4246 (N_4246,N_3039,N_3929);
xnor U4247 (N_4247,N_3510,N_3208);
nand U4248 (N_4248,N_3214,N_3172);
or U4249 (N_4249,N_3415,N_3660);
or U4250 (N_4250,N_3021,N_3798);
and U4251 (N_4251,N_3768,N_3441);
nand U4252 (N_4252,N_3804,N_3382);
nor U4253 (N_4253,N_3916,N_3620);
nand U4254 (N_4254,N_3466,N_3577);
nand U4255 (N_4255,N_3659,N_3785);
nor U4256 (N_4256,N_3326,N_3430);
or U4257 (N_4257,N_3226,N_3351);
nor U4258 (N_4258,N_3907,N_3528);
nand U4259 (N_4259,N_3556,N_3296);
or U4260 (N_4260,N_3788,N_3086);
nor U4261 (N_4261,N_3065,N_3595);
or U4262 (N_4262,N_3465,N_3749);
nand U4263 (N_4263,N_3235,N_3467);
nor U4264 (N_4264,N_3331,N_3481);
and U4265 (N_4265,N_3026,N_3515);
nor U4266 (N_4266,N_3420,N_3604);
nand U4267 (N_4267,N_3272,N_3340);
and U4268 (N_4268,N_3590,N_3645);
and U4269 (N_4269,N_3031,N_3425);
or U4270 (N_4270,N_3344,N_3740);
or U4271 (N_4271,N_3832,N_3653);
nand U4272 (N_4272,N_3373,N_3781);
or U4273 (N_4273,N_3786,N_3778);
nand U4274 (N_4274,N_3717,N_3875);
or U4275 (N_4275,N_3732,N_3598);
and U4276 (N_4276,N_3082,N_3817);
nand U4277 (N_4277,N_3107,N_3502);
nor U4278 (N_4278,N_3743,N_3601);
or U4279 (N_4279,N_3818,N_3810);
xor U4280 (N_4280,N_3090,N_3843);
nand U4281 (N_4281,N_3709,N_3876);
or U4282 (N_4282,N_3596,N_3874);
xor U4283 (N_4283,N_3543,N_3729);
and U4284 (N_4284,N_3009,N_3952);
or U4285 (N_4285,N_3250,N_3542);
nor U4286 (N_4286,N_3148,N_3129);
nand U4287 (N_4287,N_3977,N_3052);
and U4288 (N_4288,N_3599,N_3099);
nor U4289 (N_4289,N_3496,N_3406);
or U4290 (N_4290,N_3702,N_3944);
and U4291 (N_4291,N_3445,N_3503);
nand U4292 (N_4292,N_3193,N_3955);
and U4293 (N_4293,N_3354,N_3286);
and U4294 (N_4294,N_3390,N_3456);
nor U4295 (N_4295,N_3323,N_3249);
and U4296 (N_4296,N_3993,N_3075);
or U4297 (N_4297,N_3232,N_3828);
or U4298 (N_4298,N_3941,N_3763);
nand U4299 (N_4299,N_3686,N_3849);
xor U4300 (N_4300,N_3512,N_3937);
nand U4301 (N_4301,N_3652,N_3737);
nor U4302 (N_4302,N_3967,N_3451);
nor U4303 (N_4303,N_3877,N_3500);
or U4304 (N_4304,N_3682,N_3687);
nor U4305 (N_4305,N_3979,N_3881);
nand U4306 (N_4306,N_3084,N_3251);
nor U4307 (N_4307,N_3800,N_3473);
or U4308 (N_4308,N_3289,N_3112);
nor U4309 (N_4309,N_3858,N_3152);
nor U4310 (N_4310,N_3868,N_3342);
nor U4311 (N_4311,N_3908,N_3004);
nand U4312 (N_4312,N_3694,N_3617);
nand U4313 (N_4313,N_3661,N_3258);
or U4314 (N_4314,N_3062,N_3023);
or U4315 (N_4315,N_3897,N_3224);
nor U4316 (N_4316,N_3211,N_3523);
nand U4317 (N_4317,N_3493,N_3983);
and U4318 (N_4318,N_3896,N_3353);
and U4319 (N_4319,N_3592,N_3115);
and U4320 (N_4320,N_3066,N_3106);
nand U4321 (N_4321,N_3484,N_3219);
nor U4322 (N_4322,N_3933,N_3664);
or U4323 (N_4323,N_3132,N_3841);
and U4324 (N_4324,N_3204,N_3738);
and U4325 (N_4325,N_3819,N_3262);
nor U4326 (N_4326,N_3355,N_3308);
or U4327 (N_4327,N_3014,N_3648);
or U4328 (N_4328,N_3688,N_3424);
nor U4329 (N_4329,N_3234,N_3917);
nor U4330 (N_4330,N_3151,N_3730);
and U4331 (N_4331,N_3680,N_3437);
nand U4332 (N_4332,N_3000,N_3375);
and U4333 (N_4333,N_3829,N_3367);
nor U4334 (N_4334,N_3165,N_3958);
or U4335 (N_4335,N_3906,N_3767);
nor U4336 (N_4336,N_3784,N_3919);
or U4337 (N_4337,N_3865,N_3247);
and U4338 (N_4338,N_3181,N_3400);
and U4339 (N_4339,N_3918,N_3176);
or U4340 (N_4340,N_3779,N_3844);
or U4341 (N_4341,N_3759,N_3063);
nand U4342 (N_4342,N_3061,N_3792);
and U4343 (N_4343,N_3095,N_3864);
or U4344 (N_4344,N_3712,N_3357);
or U4345 (N_4345,N_3940,N_3227);
and U4346 (N_4346,N_3011,N_3964);
nand U4347 (N_4347,N_3593,N_3535);
nand U4348 (N_4348,N_3920,N_3124);
nand U4349 (N_4349,N_3885,N_3997);
or U4350 (N_4350,N_3570,N_3873);
or U4351 (N_4351,N_3363,N_3533);
and U4352 (N_4352,N_3307,N_3457);
and U4353 (N_4353,N_3923,N_3284);
and U4354 (N_4354,N_3433,N_3121);
nor U4355 (N_4355,N_3274,N_3383);
and U4356 (N_4356,N_3091,N_3120);
and U4357 (N_4357,N_3756,N_3094);
and U4358 (N_4358,N_3037,N_3986);
nor U4359 (N_4359,N_3884,N_3866);
nand U4360 (N_4360,N_3568,N_3074);
nor U4361 (N_4361,N_3385,N_3126);
nand U4362 (N_4362,N_3318,N_3527);
and U4363 (N_4363,N_3970,N_3073);
nor U4364 (N_4364,N_3207,N_3880);
nand U4365 (N_4365,N_3558,N_3985);
xnor U4366 (N_4366,N_3281,N_3722);
and U4367 (N_4367,N_3338,N_3292);
nor U4368 (N_4368,N_3027,N_3860);
nor U4369 (N_4369,N_3795,N_3514);
nand U4370 (N_4370,N_3823,N_3158);
nand U4371 (N_4371,N_3153,N_3734);
nor U4372 (N_4372,N_3689,N_3924);
nor U4373 (N_4373,N_3223,N_3585);
xor U4374 (N_4374,N_3805,N_3892);
nand U4375 (N_4375,N_3861,N_3253);
nand U4376 (N_4376,N_3057,N_3900);
nor U4377 (N_4377,N_3335,N_3969);
nor U4378 (N_4378,N_3267,N_3727);
nand U4379 (N_4379,N_3859,N_3032);
nand U4380 (N_4380,N_3417,N_3870);
and U4381 (N_4381,N_3282,N_3100);
and U4382 (N_4382,N_3674,N_3872);
nor U4383 (N_4383,N_3771,N_3723);
and U4384 (N_4384,N_3419,N_3462);
and U4385 (N_4385,N_3463,N_3459);
or U4386 (N_4386,N_3934,N_3442);
nor U4387 (N_4387,N_3615,N_3854);
and U4388 (N_4388,N_3128,N_3135);
nand U4389 (N_4389,N_3045,N_3436);
nor U4390 (N_4390,N_3336,N_3317);
nor U4391 (N_4391,N_3673,N_3802);
and U4392 (N_4392,N_3513,N_3190);
or U4393 (N_4393,N_3179,N_3741);
and U4394 (N_4394,N_3174,N_3490);
or U4395 (N_4395,N_3241,N_3081);
nor U4396 (N_4396,N_3978,N_3765);
and U4397 (N_4397,N_3641,N_3750);
and U4398 (N_4398,N_3752,N_3257);
nand U4399 (N_4399,N_3431,N_3087);
nor U4400 (N_4400,N_3432,N_3118);
and U4401 (N_4401,N_3787,N_3030);
or U4402 (N_4402,N_3902,N_3184);
xor U4403 (N_4403,N_3156,N_3646);
or U4404 (N_4404,N_3212,N_3935);
and U4405 (N_4405,N_3962,N_3497);
nand U4406 (N_4406,N_3796,N_3047);
and U4407 (N_4407,N_3793,N_3293);
and U4408 (N_4408,N_3141,N_3903);
nor U4409 (N_4409,N_3454,N_3960);
nor U4410 (N_4410,N_3616,N_3739);
or U4411 (N_4411,N_3581,N_3753);
and U4412 (N_4412,N_3654,N_3435);
nor U4413 (N_4413,N_3056,N_3060);
or U4414 (N_4414,N_3963,N_3931);
and U4415 (N_4415,N_3145,N_3913);
nand U4416 (N_4416,N_3049,N_3587);
nand U4417 (N_4417,N_3489,N_3665);
or U4418 (N_4418,N_3295,N_3766);
nand U4419 (N_4419,N_3202,N_3102);
nor U4420 (N_4420,N_3815,N_3834);
or U4421 (N_4421,N_3541,N_3526);
or U4422 (N_4422,N_3092,N_3168);
nor U4423 (N_4423,N_3744,N_3450);
and U4424 (N_4424,N_3520,N_3705);
and U4425 (N_4425,N_3684,N_3134);
and U4426 (N_4426,N_3408,N_3708);
or U4427 (N_4427,N_3322,N_3412);
nand U4428 (N_4428,N_3745,N_3998);
and U4429 (N_4429,N_3418,N_3580);
and U4430 (N_4430,N_3693,N_3758);
or U4431 (N_4431,N_3610,N_3388);
or U4432 (N_4432,N_3530,N_3378);
and U4433 (N_4433,N_3850,N_3018);
nand U4434 (N_4434,N_3700,N_3644);
nand U4435 (N_4435,N_3562,N_3469);
or U4436 (N_4436,N_3379,N_3157);
nor U4437 (N_4437,N_3965,N_3259);
or U4438 (N_4438,N_3612,N_3025);
nor U4439 (N_4439,N_3783,N_3928);
nand U4440 (N_4440,N_3618,N_3474);
xnor U4441 (N_4441,N_3352,N_3130);
and U4442 (N_4442,N_3079,N_3770);
and U4443 (N_4443,N_3711,N_3769);
or U4444 (N_4444,N_3240,N_3475);
and U4445 (N_4445,N_3814,N_3681);
nor U4446 (N_4446,N_3564,N_3005);
nor U4447 (N_4447,N_3699,N_3735);
or U4448 (N_4448,N_3362,N_3567);
nand U4449 (N_4449,N_3724,N_3662);
nand U4450 (N_4450,N_3279,N_3536);
nor U4451 (N_4451,N_3820,N_3159);
or U4452 (N_4452,N_3316,N_3345);
or U4453 (N_4453,N_3213,N_3140);
nand U4454 (N_4454,N_3482,N_3586);
nand U4455 (N_4455,N_3511,N_3760);
nand U4456 (N_4456,N_3889,N_3886);
or U4457 (N_4457,N_3716,N_3096);
and U4458 (N_4458,N_3035,N_3411);
nor U4459 (N_4459,N_3498,N_3149);
nand U4460 (N_4460,N_3632,N_3070);
nand U4461 (N_4461,N_3634,N_3776);
nand U4462 (N_4462,N_3692,N_3347);
nand U4463 (N_4463,N_3228,N_3299);
or U4464 (N_4464,N_3252,N_3614);
or U4465 (N_4465,N_3494,N_3775);
or U4466 (N_4466,N_3578,N_3161);
or U4467 (N_4467,N_3666,N_3444);
nand U4468 (N_4468,N_3006,N_3583);
or U4469 (N_4469,N_3313,N_3672);
nor U4470 (N_4470,N_3742,N_3630);
or U4471 (N_4471,N_3971,N_3155);
or U4472 (N_4472,N_3022,N_3495);
and U4473 (N_4473,N_3731,N_3773);
nand U4474 (N_4474,N_3842,N_3633);
nor U4475 (N_4475,N_3243,N_3720);
xnor U4476 (N_4476,N_3898,N_3506);
and U4477 (N_4477,N_3816,N_3034);
nand U4478 (N_4478,N_3905,N_3531);
and U4479 (N_4479,N_3504,N_3574);
and U4480 (N_4480,N_3517,N_3300);
or U4481 (N_4481,N_3203,N_3671);
nand U4482 (N_4482,N_3072,N_3216);
or U4483 (N_4483,N_3210,N_3173);
nor U4484 (N_4484,N_3762,N_3894);
or U4485 (N_4485,N_3170,N_3619);
or U4486 (N_4486,N_3548,N_3175);
or U4487 (N_4487,N_3746,N_3939);
xor U4488 (N_4488,N_3840,N_3552);
nand U4489 (N_4489,N_3826,N_3607);
or U4490 (N_4490,N_3098,N_3863);
and U4491 (N_4491,N_3949,N_3085);
or U4492 (N_4492,N_3356,N_3205);
nor U4493 (N_4493,N_3187,N_3824);
nand U4494 (N_4494,N_3912,N_3862);
or U4495 (N_4495,N_3747,N_3404);
and U4496 (N_4496,N_3447,N_3951);
and U4497 (N_4497,N_3544,N_3803);
and U4498 (N_4498,N_3138,N_3807);
or U4499 (N_4499,N_3835,N_3545);
or U4500 (N_4500,N_3865,N_3710);
or U4501 (N_4501,N_3654,N_3929);
nor U4502 (N_4502,N_3613,N_3785);
and U4503 (N_4503,N_3043,N_3676);
nand U4504 (N_4504,N_3420,N_3251);
or U4505 (N_4505,N_3698,N_3763);
nand U4506 (N_4506,N_3397,N_3596);
nand U4507 (N_4507,N_3710,N_3905);
and U4508 (N_4508,N_3141,N_3362);
nor U4509 (N_4509,N_3788,N_3446);
and U4510 (N_4510,N_3021,N_3210);
nor U4511 (N_4511,N_3827,N_3147);
nand U4512 (N_4512,N_3496,N_3656);
nand U4513 (N_4513,N_3157,N_3246);
and U4514 (N_4514,N_3272,N_3777);
nor U4515 (N_4515,N_3559,N_3687);
nand U4516 (N_4516,N_3591,N_3317);
or U4517 (N_4517,N_3786,N_3631);
and U4518 (N_4518,N_3563,N_3961);
nand U4519 (N_4519,N_3853,N_3475);
or U4520 (N_4520,N_3566,N_3421);
nor U4521 (N_4521,N_3953,N_3553);
nand U4522 (N_4522,N_3319,N_3800);
nor U4523 (N_4523,N_3691,N_3542);
or U4524 (N_4524,N_3517,N_3768);
or U4525 (N_4525,N_3445,N_3562);
nor U4526 (N_4526,N_3025,N_3458);
nand U4527 (N_4527,N_3284,N_3493);
or U4528 (N_4528,N_3431,N_3537);
and U4529 (N_4529,N_3906,N_3233);
nand U4530 (N_4530,N_3726,N_3040);
nor U4531 (N_4531,N_3991,N_3398);
nand U4532 (N_4532,N_3568,N_3329);
or U4533 (N_4533,N_3786,N_3069);
nor U4534 (N_4534,N_3498,N_3129);
and U4535 (N_4535,N_3301,N_3093);
and U4536 (N_4536,N_3331,N_3018);
and U4537 (N_4537,N_3178,N_3546);
or U4538 (N_4538,N_3014,N_3508);
nor U4539 (N_4539,N_3725,N_3286);
nand U4540 (N_4540,N_3566,N_3486);
nor U4541 (N_4541,N_3265,N_3803);
nand U4542 (N_4542,N_3618,N_3563);
or U4543 (N_4543,N_3740,N_3184);
nand U4544 (N_4544,N_3310,N_3702);
nor U4545 (N_4545,N_3709,N_3112);
and U4546 (N_4546,N_3059,N_3405);
and U4547 (N_4547,N_3867,N_3525);
nor U4548 (N_4548,N_3566,N_3660);
and U4549 (N_4549,N_3852,N_3159);
and U4550 (N_4550,N_3759,N_3566);
or U4551 (N_4551,N_3554,N_3005);
and U4552 (N_4552,N_3302,N_3114);
and U4553 (N_4553,N_3803,N_3501);
nor U4554 (N_4554,N_3440,N_3038);
nor U4555 (N_4555,N_3257,N_3804);
nor U4556 (N_4556,N_3409,N_3236);
nor U4557 (N_4557,N_3511,N_3712);
nor U4558 (N_4558,N_3583,N_3708);
or U4559 (N_4559,N_3935,N_3503);
or U4560 (N_4560,N_3968,N_3684);
and U4561 (N_4561,N_3237,N_3097);
nor U4562 (N_4562,N_3155,N_3236);
or U4563 (N_4563,N_3740,N_3715);
nor U4564 (N_4564,N_3751,N_3339);
nand U4565 (N_4565,N_3196,N_3295);
nor U4566 (N_4566,N_3423,N_3455);
nor U4567 (N_4567,N_3963,N_3002);
nand U4568 (N_4568,N_3638,N_3810);
nor U4569 (N_4569,N_3536,N_3783);
nand U4570 (N_4570,N_3928,N_3788);
and U4571 (N_4571,N_3373,N_3885);
xnor U4572 (N_4572,N_3694,N_3803);
nand U4573 (N_4573,N_3104,N_3893);
or U4574 (N_4574,N_3206,N_3397);
and U4575 (N_4575,N_3755,N_3061);
nor U4576 (N_4576,N_3001,N_3653);
nor U4577 (N_4577,N_3927,N_3025);
nand U4578 (N_4578,N_3591,N_3694);
nand U4579 (N_4579,N_3090,N_3901);
nor U4580 (N_4580,N_3980,N_3873);
nand U4581 (N_4581,N_3570,N_3776);
nor U4582 (N_4582,N_3490,N_3505);
nor U4583 (N_4583,N_3717,N_3735);
or U4584 (N_4584,N_3891,N_3671);
and U4585 (N_4585,N_3142,N_3537);
nand U4586 (N_4586,N_3335,N_3025);
or U4587 (N_4587,N_3169,N_3490);
nor U4588 (N_4588,N_3178,N_3427);
and U4589 (N_4589,N_3713,N_3931);
and U4590 (N_4590,N_3807,N_3487);
and U4591 (N_4591,N_3910,N_3483);
nor U4592 (N_4592,N_3096,N_3514);
nand U4593 (N_4593,N_3455,N_3544);
nand U4594 (N_4594,N_3627,N_3836);
or U4595 (N_4595,N_3947,N_3102);
nand U4596 (N_4596,N_3241,N_3942);
nor U4597 (N_4597,N_3202,N_3192);
or U4598 (N_4598,N_3653,N_3572);
nor U4599 (N_4599,N_3342,N_3260);
nor U4600 (N_4600,N_3963,N_3800);
nor U4601 (N_4601,N_3023,N_3325);
and U4602 (N_4602,N_3883,N_3482);
or U4603 (N_4603,N_3638,N_3975);
or U4604 (N_4604,N_3864,N_3771);
nor U4605 (N_4605,N_3948,N_3198);
nand U4606 (N_4606,N_3311,N_3947);
and U4607 (N_4607,N_3350,N_3273);
nor U4608 (N_4608,N_3380,N_3933);
and U4609 (N_4609,N_3824,N_3458);
and U4610 (N_4610,N_3770,N_3176);
and U4611 (N_4611,N_3960,N_3872);
xor U4612 (N_4612,N_3564,N_3420);
nand U4613 (N_4613,N_3722,N_3256);
or U4614 (N_4614,N_3128,N_3357);
and U4615 (N_4615,N_3313,N_3363);
and U4616 (N_4616,N_3991,N_3540);
or U4617 (N_4617,N_3060,N_3015);
nor U4618 (N_4618,N_3272,N_3264);
or U4619 (N_4619,N_3266,N_3782);
nand U4620 (N_4620,N_3420,N_3216);
and U4621 (N_4621,N_3978,N_3804);
and U4622 (N_4622,N_3655,N_3433);
nor U4623 (N_4623,N_3281,N_3871);
and U4624 (N_4624,N_3685,N_3304);
xor U4625 (N_4625,N_3689,N_3711);
nor U4626 (N_4626,N_3705,N_3535);
and U4627 (N_4627,N_3686,N_3953);
and U4628 (N_4628,N_3739,N_3225);
or U4629 (N_4629,N_3976,N_3831);
and U4630 (N_4630,N_3180,N_3396);
nand U4631 (N_4631,N_3056,N_3765);
or U4632 (N_4632,N_3001,N_3593);
and U4633 (N_4633,N_3920,N_3027);
and U4634 (N_4634,N_3850,N_3278);
nor U4635 (N_4635,N_3103,N_3961);
nor U4636 (N_4636,N_3771,N_3072);
nor U4637 (N_4637,N_3208,N_3351);
nor U4638 (N_4638,N_3072,N_3353);
nor U4639 (N_4639,N_3110,N_3842);
nand U4640 (N_4640,N_3085,N_3253);
or U4641 (N_4641,N_3682,N_3199);
or U4642 (N_4642,N_3012,N_3418);
xor U4643 (N_4643,N_3008,N_3181);
nand U4644 (N_4644,N_3746,N_3590);
or U4645 (N_4645,N_3585,N_3970);
or U4646 (N_4646,N_3484,N_3877);
and U4647 (N_4647,N_3053,N_3718);
nand U4648 (N_4648,N_3751,N_3311);
nor U4649 (N_4649,N_3300,N_3322);
nor U4650 (N_4650,N_3343,N_3885);
nand U4651 (N_4651,N_3054,N_3428);
nand U4652 (N_4652,N_3274,N_3962);
nor U4653 (N_4653,N_3951,N_3136);
xor U4654 (N_4654,N_3157,N_3916);
nor U4655 (N_4655,N_3302,N_3778);
and U4656 (N_4656,N_3832,N_3845);
nand U4657 (N_4657,N_3737,N_3860);
or U4658 (N_4658,N_3799,N_3226);
nand U4659 (N_4659,N_3524,N_3311);
nand U4660 (N_4660,N_3102,N_3291);
nor U4661 (N_4661,N_3335,N_3126);
and U4662 (N_4662,N_3617,N_3757);
and U4663 (N_4663,N_3699,N_3008);
nor U4664 (N_4664,N_3736,N_3645);
and U4665 (N_4665,N_3023,N_3777);
or U4666 (N_4666,N_3233,N_3637);
or U4667 (N_4667,N_3566,N_3528);
nor U4668 (N_4668,N_3928,N_3557);
and U4669 (N_4669,N_3911,N_3346);
and U4670 (N_4670,N_3350,N_3417);
or U4671 (N_4671,N_3779,N_3857);
nand U4672 (N_4672,N_3786,N_3535);
nand U4673 (N_4673,N_3631,N_3461);
nor U4674 (N_4674,N_3921,N_3074);
xnor U4675 (N_4675,N_3214,N_3110);
or U4676 (N_4676,N_3082,N_3233);
or U4677 (N_4677,N_3318,N_3112);
or U4678 (N_4678,N_3236,N_3273);
and U4679 (N_4679,N_3975,N_3522);
or U4680 (N_4680,N_3117,N_3522);
nand U4681 (N_4681,N_3721,N_3844);
nand U4682 (N_4682,N_3644,N_3642);
and U4683 (N_4683,N_3116,N_3089);
nor U4684 (N_4684,N_3143,N_3112);
or U4685 (N_4685,N_3093,N_3871);
and U4686 (N_4686,N_3597,N_3352);
nor U4687 (N_4687,N_3964,N_3017);
and U4688 (N_4688,N_3136,N_3904);
and U4689 (N_4689,N_3567,N_3703);
or U4690 (N_4690,N_3481,N_3678);
nor U4691 (N_4691,N_3016,N_3834);
and U4692 (N_4692,N_3958,N_3555);
or U4693 (N_4693,N_3427,N_3722);
nand U4694 (N_4694,N_3223,N_3028);
nor U4695 (N_4695,N_3598,N_3222);
nand U4696 (N_4696,N_3305,N_3591);
or U4697 (N_4697,N_3114,N_3678);
xor U4698 (N_4698,N_3116,N_3510);
and U4699 (N_4699,N_3153,N_3438);
and U4700 (N_4700,N_3167,N_3673);
nand U4701 (N_4701,N_3196,N_3804);
nand U4702 (N_4702,N_3966,N_3456);
and U4703 (N_4703,N_3974,N_3141);
or U4704 (N_4704,N_3383,N_3826);
or U4705 (N_4705,N_3845,N_3514);
or U4706 (N_4706,N_3616,N_3210);
nor U4707 (N_4707,N_3606,N_3225);
nand U4708 (N_4708,N_3917,N_3349);
nand U4709 (N_4709,N_3660,N_3326);
and U4710 (N_4710,N_3597,N_3033);
xnor U4711 (N_4711,N_3632,N_3556);
or U4712 (N_4712,N_3043,N_3839);
or U4713 (N_4713,N_3465,N_3999);
nor U4714 (N_4714,N_3966,N_3535);
or U4715 (N_4715,N_3734,N_3708);
nor U4716 (N_4716,N_3346,N_3995);
nor U4717 (N_4717,N_3707,N_3349);
and U4718 (N_4718,N_3308,N_3432);
and U4719 (N_4719,N_3615,N_3154);
nor U4720 (N_4720,N_3144,N_3945);
and U4721 (N_4721,N_3363,N_3450);
nand U4722 (N_4722,N_3816,N_3376);
or U4723 (N_4723,N_3904,N_3169);
nor U4724 (N_4724,N_3920,N_3651);
nand U4725 (N_4725,N_3734,N_3239);
nand U4726 (N_4726,N_3763,N_3645);
and U4727 (N_4727,N_3832,N_3192);
or U4728 (N_4728,N_3295,N_3672);
nand U4729 (N_4729,N_3990,N_3782);
nand U4730 (N_4730,N_3099,N_3076);
xor U4731 (N_4731,N_3181,N_3829);
nand U4732 (N_4732,N_3290,N_3376);
and U4733 (N_4733,N_3331,N_3726);
or U4734 (N_4734,N_3644,N_3340);
or U4735 (N_4735,N_3385,N_3065);
nand U4736 (N_4736,N_3189,N_3738);
and U4737 (N_4737,N_3135,N_3379);
nand U4738 (N_4738,N_3553,N_3792);
or U4739 (N_4739,N_3173,N_3768);
nand U4740 (N_4740,N_3445,N_3790);
nor U4741 (N_4741,N_3357,N_3356);
and U4742 (N_4742,N_3389,N_3178);
and U4743 (N_4743,N_3902,N_3082);
nand U4744 (N_4744,N_3796,N_3594);
and U4745 (N_4745,N_3241,N_3460);
or U4746 (N_4746,N_3785,N_3805);
nor U4747 (N_4747,N_3044,N_3759);
and U4748 (N_4748,N_3292,N_3973);
nand U4749 (N_4749,N_3691,N_3963);
nand U4750 (N_4750,N_3408,N_3670);
xnor U4751 (N_4751,N_3490,N_3627);
nor U4752 (N_4752,N_3960,N_3828);
nor U4753 (N_4753,N_3988,N_3486);
nor U4754 (N_4754,N_3291,N_3522);
and U4755 (N_4755,N_3402,N_3926);
and U4756 (N_4756,N_3179,N_3674);
nand U4757 (N_4757,N_3856,N_3727);
or U4758 (N_4758,N_3852,N_3434);
or U4759 (N_4759,N_3151,N_3004);
or U4760 (N_4760,N_3266,N_3532);
xor U4761 (N_4761,N_3459,N_3210);
and U4762 (N_4762,N_3596,N_3169);
or U4763 (N_4763,N_3859,N_3704);
or U4764 (N_4764,N_3286,N_3405);
and U4765 (N_4765,N_3623,N_3701);
or U4766 (N_4766,N_3617,N_3205);
nand U4767 (N_4767,N_3454,N_3707);
and U4768 (N_4768,N_3566,N_3490);
and U4769 (N_4769,N_3469,N_3320);
nor U4770 (N_4770,N_3350,N_3477);
and U4771 (N_4771,N_3248,N_3510);
nor U4772 (N_4772,N_3914,N_3873);
and U4773 (N_4773,N_3974,N_3834);
and U4774 (N_4774,N_3394,N_3865);
and U4775 (N_4775,N_3052,N_3107);
nand U4776 (N_4776,N_3385,N_3028);
nand U4777 (N_4777,N_3952,N_3837);
nand U4778 (N_4778,N_3713,N_3327);
nand U4779 (N_4779,N_3547,N_3405);
nor U4780 (N_4780,N_3976,N_3710);
nand U4781 (N_4781,N_3532,N_3909);
nand U4782 (N_4782,N_3757,N_3690);
and U4783 (N_4783,N_3366,N_3115);
nand U4784 (N_4784,N_3460,N_3243);
or U4785 (N_4785,N_3309,N_3705);
and U4786 (N_4786,N_3014,N_3607);
or U4787 (N_4787,N_3761,N_3957);
nand U4788 (N_4788,N_3984,N_3690);
nand U4789 (N_4789,N_3353,N_3455);
and U4790 (N_4790,N_3895,N_3111);
nand U4791 (N_4791,N_3272,N_3774);
and U4792 (N_4792,N_3610,N_3018);
or U4793 (N_4793,N_3145,N_3380);
and U4794 (N_4794,N_3747,N_3960);
nand U4795 (N_4795,N_3895,N_3632);
nor U4796 (N_4796,N_3740,N_3547);
or U4797 (N_4797,N_3166,N_3794);
or U4798 (N_4798,N_3286,N_3233);
and U4799 (N_4799,N_3844,N_3543);
and U4800 (N_4800,N_3143,N_3102);
and U4801 (N_4801,N_3024,N_3059);
or U4802 (N_4802,N_3395,N_3421);
and U4803 (N_4803,N_3249,N_3948);
and U4804 (N_4804,N_3370,N_3474);
or U4805 (N_4805,N_3904,N_3092);
or U4806 (N_4806,N_3402,N_3585);
nor U4807 (N_4807,N_3172,N_3577);
nand U4808 (N_4808,N_3347,N_3145);
nand U4809 (N_4809,N_3576,N_3263);
and U4810 (N_4810,N_3092,N_3730);
xor U4811 (N_4811,N_3537,N_3781);
or U4812 (N_4812,N_3526,N_3902);
nand U4813 (N_4813,N_3379,N_3064);
nand U4814 (N_4814,N_3446,N_3625);
nand U4815 (N_4815,N_3184,N_3703);
nand U4816 (N_4816,N_3799,N_3555);
nand U4817 (N_4817,N_3914,N_3039);
nand U4818 (N_4818,N_3078,N_3850);
and U4819 (N_4819,N_3380,N_3570);
nand U4820 (N_4820,N_3076,N_3784);
nand U4821 (N_4821,N_3535,N_3954);
or U4822 (N_4822,N_3787,N_3628);
and U4823 (N_4823,N_3332,N_3989);
nor U4824 (N_4824,N_3818,N_3165);
nor U4825 (N_4825,N_3510,N_3672);
nor U4826 (N_4826,N_3527,N_3471);
nor U4827 (N_4827,N_3505,N_3234);
nor U4828 (N_4828,N_3680,N_3660);
nand U4829 (N_4829,N_3685,N_3176);
and U4830 (N_4830,N_3202,N_3248);
nand U4831 (N_4831,N_3755,N_3383);
nand U4832 (N_4832,N_3534,N_3865);
or U4833 (N_4833,N_3200,N_3399);
nor U4834 (N_4834,N_3227,N_3775);
and U4835 (N_4835,N_3476,N_3027);
and U4836 (N_4836,N_3253,N_3395);
and U4837 (N_4837,N_3863,N_3537);
nor U4838 (N_4838,N_3905,N_3295);
or U4839 (N_4839,N_3764,N_3222);
and U4840 (N_4840,N_3407,N_3280);
or U4841 (N_4841,N_3252,N_3712);
nor U4842 (N_4842,N_3438,N_3876);
or U4843 (N_4843,N_3358,N_3290);
and U4844 (N_4844,N_3018,N_3593);
and U4845 (N_4845,N_3087,N_3487);
nand U4846 (N_4846,N_3703,N_3417);
xnor U4847 (N_4847,N_3093,N_3372);
and U4848 (N_4848,N_3892,N_3694);
nand U4849 (N_4849,N_3196,N_3369);
or U4850 (N_4850,N_3081,N_3700);
and U4851 (N_4851,N_3929,N_3470);
nand U4852 (N_4852,N_3438,N_3701);
and U4853 (N_4853,N_3639,N_3565);
nand U4854 (N_4854,N_3969,N_3857);
nand U4855 (N_4855,N_3897,N_3703);
nand U4856 (N_4856,N_3422,N_3742);
and U4857 (N_4857,N_3213,N_3326);
nand U4858 (N_4858,N_3413,N_3273);
or U4859 (N_4859,N_3433,N_3112);
nand U4860 (N_4860,N_3707,N_3946);
and U4861 (N_4861,N_3028,N_3295);
or U4862 (N_4862,N_3496,N_3645);
nand U4863 (N_4863,N_3058,N_3187);
nand U4864 (N_4864,N_3699,N_3253);
nand U4865 (N_4865,N_3859,N_3869);
or U4866 (N_4866,N_3865,N_3365);
or U4867 (N_4867,N_3097,N_3999);
nand U4868 (N_4868,N_3268,N_3003);
and U4869 (N_4869,N_3321,N_3153);
or U4870 (N_4870,N_3420,N_3672);
and U4871 (N_4871,N_3482,N_3091);
and U4872 (N_4872,N_3516,N_3303);
or U4873 (N_4873,N_3954,N_3185);
or U4874 (N_4874,N_3679,N_3935);
or U4875 (N_4875,N_3763,N_3786);
nand U4876 (N_4876,N_3213,N_3918);
nor U4877 (N_4877,N_3363,N_3103);
or U4878 (N_4878,N_3916,N_3181);
nand U4879 (N_4879,N_3151,N_3712);
and U4880 (N_4880,N_3567,N_3971);
nor U4881 (N_4881,N_3352,N_3279);
and U4882 (N_4882,N_3936,N_3002);
or U4883 (N_4883,N_3733,N_3387);
nor U4884 (N_4884,N_3832,N_3928);
or U4885 (N_4885,N_3853,N_3758);
nand U4886 (N_4886,N_3317,N_3051);
nor U4887 (N_4887,N_3235,N_3659);
nand U4888 (N_4888,N_3585,N_3211);
or U4889 (N_4889,N_3165,N_3738);
nor U4890 (N_4890,N_3666,N_3045);
and U4891 (N_4891,N_3722,N_3444);
xor U4892 (N_4892,N_3643,N_3090);
nand U4893 (N_4893,N_3346,N_3416);
or U4894 (N_4894,N_3731,N_3328);
nand U4895 (N_4895,N_3497,N_3383);
nand U4896 (N_4896,N_3171,N_3283);
and U4897 (N_4897,N_3953,N_3361);
nand U4898 (N_4898,N_3598,N_3145);
and U4899 (N_4899,N_3194,N_3873);
nand U4900 (N_4900,N_3041,N_3796);
nor U4901 (N_4901,N_3978,N_3967);
xnor U4902 (N_4902,N_3181,N_3088);
or U4903 (N_4903,N_3830,N_3105);
and U4904 (N_4904,N_3653,N_3708);
nor U4905 (N_4905,N_3620,N_3807);
nand U4906 (N_4906,N_3231,N_3722);
nand U4907 (N_4907,N_3381,N_3023);
nand U4908 (N_4908,N_3142,N_3197);
and U4909 (N_4909,N_3142,N_3980);
nor U4910 (N_4910,N_3754,N_3437);
and U4911 (N_4911,N_3255,N_3689);
or U4912 (N_4912,N_3694,N_3336);
nor U4913 (N_4913,N_3789,N_3225);
and U4914 (N_4914,N_3665,N_3734);
or U4915 (N_4915,N_3273,N_3873);
nor U4916 (N_4916,N_3095,N_3158);
xor U4917 (N_4917,N_3395,N_3676);
or U4918 (N_4918,N_3236,N_3960);
or U4919 (N_4919,N_3025,N_3339);
nor U4920 (N_4920,N_3309,N_3446);
and U4921 (N_4921,N_3062,N_3006);
nor U4922 (N_4922,N_3993,N_3971);
nand U4923 (N_4923,N_3970,N_3972);
nand U4924 (N_4924,N_3408,N_3414);
nor U4925 (N_4925,N_3380,N_3742);
or U4926 (N_4926,N_3071,N_3423);
nor U4927 (N_4927,N_3486,N_3798);
or U4928 (N_4928,N_3302,N_3558);
and U4929 (N_4929,N_3935,N_3865);
nand U4930 (N_4930,N_3584,N_3128);
nor U4931 (N_4931,N_3216,N_3342);
and U4932 (N_4932,N_3999,N_3908);
xor U4933 (N_4933,N_3282,N_3470);
or U4934 (N_4934,N_3905,N_3537);
or U4935 (N_4935,N_3352,N_3184);
and U4936 (N_4936,N_3622,N_3366);
and U4937 (N_4937,N_3093,N_3270);
nor U4938 (N_4938,N_3874,N_3035);
nand U4939 (N_4939,N_3922,N_3757);
nand U4940 (N_4940,N_3857,N_3862);
nor U4941 (N_4941,N_3248,N_3033);
or U4942 (N_4942,N_3293,N_3996);
nand U4943 (N_4943,N_3916,N_3671);
nor U4944 (N_4944,N_3607,N_3368);
nand U4945 (N_4945,N_3687,N_3667);
nand U4946 (N_4946,N_3256,N_3081);
and U4947 (N_4947,N_3750,N_3320);
or U4948 (N_4948,N_3681,N_3864);
nand U4949 (N_4949,N_3296,N_3069);
nand U4950 (N_4950,N_3351,N_3537);
nor U4951 (N_4951,N_3477,N_3033);
and U4952 (N_4952,N_3732,N_3781);
or U4953 (N_4953,N_3646,N_3878);
or U4954 (N_4954,N_3213,N_3268);
or U4955 (N_4955,N_3209,N_3736);
and U4956 (N_4956,N_3418,N_3800);
nor U4957 (N_4957,N_3662,N_3784);
nor U4958 (N_4958,N_3624,N_3094);
nor U4959 (N_4959,N_3436,N_3382);
nor U4960 (N_4960,N_3568,N_3348);
or U4961 (N_4961,N_3809,N_3743);
nand U4962 (N_4962,N_3005,N_3606);
and U4963 (N_4963,N_3952,N_3591);
nand U4964 (N_4964,N_3722,N_3645);
nor U4965 (N_4965,N_3913,N_3469);
nand U4966 (N_4966,N_3098,N_3055);
nand U4967 (N_4967,N_3242,N_3698);
nor U4968 (N_4968,N_3595,N_3822);
or U4969 (N_4969,N_3273,N_3707);
nor U4970 (N_4970,N_3205,N_3909);
nor U4971 (N_4971,N_3238,N_3863);
or U4972 (N_4972,N_3407,N_3729);
nand U4973 (N_4973,N_3275,N_3211);
nand U4974 (N_4974,N_3000,N_3910);
nand U4975 (N_4975,N_3167,N_3971);
and U4976 (N_4976,N_3248,N_3891);
nand U4977 (N_4977,N_3589,N_3287);
nand U4978 (N_4978,N_3304,N_3631);
nor U4979 (N_4979,N_3956,N_3352);
and U4980 (N_4980,N_3343,N_3092);
or U4981 (N_4981,N_3516,N_3143);
or U4982 (N_4982,N_3509,N_3880);
and U4983 (N_4983,N_3134,N_3882);
and U4984 (N_4984,N_3713,N_3595);
and U4985 (N_4985,N_3042,N_3389);
and U4986 (N_4986,N_3823,N_3768);
nand U4987 (N_4987,N_3068,N_3008);
nor U4988 (N_4988,N_3455,N_3411);
nand U4989 (N_4989,N_3330,N_3968);
nor U4990 (N_4990,N_3301,N_3679);
or U4991 (N_4991,N_3199,N_3743);
and U4992 (N_4992,N_3721,N_3401);
nand U4993 (N_4993,N_3338,N_3231);
or U4994 (N_4994,N_3327,N_3952);
or U4995 (N_4995,N_3116,N_3399);
and U4996 (N_4996,N_3056,N_3330);
and U4997 (N_4997,N_3588,N_3478);
nand U4998 (N_4998,N_3876,N_3108);
or U4999 (N_4999,N_3286,N_3113);
and U5000 (N_5000,N_4650,N_4883);
nand U5001 (N_5001,N_4282,N_4734);
nand U5002 (N_5002,N_4008,N_4295);
nor U5003 (N_5003,N_4474,N_4460);
nor U5004 (N_5004,N_4131,N_4330);
or U5005 (N_5005,N_4538,N_4658);
nand U5006 (N_5006,N_4517,N_4497);
nor U5007 (N_5007,N_4750,N_4696);
or U5008 (N_5008,N_4501,N_4686);
and U5009 (N_5009,N_4975,N_4439);
nor U5010 (N_5010,N_4258,N_4444);
or U5011 (N_5011,N_4020,N_4708);
nand U5012 (N_5012,N_4832,N_4056);
nor U5013 (N_5013,N_4300,N_4087);
nor U5014 (N_5014,N_4122,N_4892);
nor U5015 (N_5015,N_4854,N_4745);
or U5016 (N_5016,N_4287,N_4338);
nand U5017 (N_5017,N_4681,N_4978);
xnor U5018 (N_5018,N_4949,N_4553);
and U5019 (N_5019,N_4566,N_4368);
nand U5020 (N_5020,N_4396,N_4414);
nand U5021 (N_5021,N_4349,N_4445);
or U5022 (N_5022,N_4274,N_4625);
or U5023 (N_5023,N_4329,N_4915);
nand U5024 (N_5024,N_4522,N_4134);
nand U5025 (N_5025,N_4255,N_4744);
nand U5026 (N_5026,N_4851,N_4455);
nand U5027 (N_5027,N_4028,N_4470);
or U5028 (N_5028,N_4392,N_4328);
and U5029 (N_5029,N_4977,N_4839);
or U5030 (N_5030,N_4614,N_4551);
nand U5031 (N_5031,N_4194,N_4077);
or U5032 (N_5032,N_4174,N_4072);
nand U5033 (N_5033,N_4270,N_4906);
and U5034 (N_5034,N_4647,N_4506);
or U5035 (N_5035,N_4990,N_4148);
or U5036 (N_5036,N_4342,N_4313);
or U5037 (N_5037,N_4733,N_4714);
nand U5038 (N_5038,N_4905,N_4133);
or U5039 (N_5039,N_4753,N_4026);
nand U5040 (N_5040,N_4556,N_4042);
nand U5041 (N_5041,N_4680,N_4066);
xnor U5042 (N_5042,N_4019,N_4656);
nand U5043 (N_5043,N_4966,N_4081);
or U5044 (N_5044,N_4639,N_4523);
and U5045 (N_5045,N_4128,N_4281);
nand U5046 (N_5046,N_4568,N_4251);
or U5047 (N_5047,N_4849,N_4908);
nand U5048 (N_5048,N_4715,N_4540);
nand U5049 (N_5049,N_4979,N_4557);
nand U5050 (N_5050,N_4651,N_4668);
nor U5051 (N_5051,N_4789,N_4592);
and U5052 (N_5052,N_4593,N_4301);
nand U5053 (N_5053,N_4069,N_4828);
nor U5054 (N_5054,N_4196,N_4292);
and U5055 (N_5055,N_4483,N_4958);
or U5056 (N_5056,N_4306,N_4138);
or U5057 (N_5057,N_4907,N_4935);
nand U5058 (N_5058,N_4494,N_4771);
nand U5059 (N_5059,N_4332,N_4199);
or U5060 (N_5060,N_4456,N_4446);
and U5061 (N_5061,N_4610,N_4272);
nand U5062 (N_5062,N_4297,N_4206);
and U5063 (N_5063,N_4290,N_4805);
and U5064 (N_5064,N_4426,N_4397);
nor U5065 (N_5065,N_4302,N_4182);
or U5066 (N_5066,N_4343,N_4642);
xor U5067 (N_5067,N_4640,N_4660);
nor U5068 (N_5068,N_4067,N_4682);
nor U5069 (N_5069,N_4711,N_4175);
nand U5070 (N_5070,N_4351,N_4560);
or U5071 (N_5071,N_4574,N_4955);
nor U5072 (N_5072,N_4847,N_4068);
and U5073 (N_5073,N_4399,N_4312);
or U5074 (N_5074,N_4146,N_4661);
or U5075 (N_5075,N_4732,N_4524);
or U5076 (N_5076,N_4829,N_4741);
or U5077 (N_5077,N_4794,N_4029);
and U5078 (N_5078,N_4142,N_4369);
nand U5079 (N_5079,N_4362,N_4213);
and U5080 (N_5080,N_4109,N_4018);
nand U5081 (N_5081,N_4846,N_4821);
and U5082 (N_5082,N_4432,N_4289);
and U5083 (N_5083,N_4389,N_4621);
nor U5084 (N_5084,N_4406,N_4463);
nor U5085 (N_5085,N_4939,N_4735);
or U5086 (N_5086,N_4638,N_4319);
nor U5087 (N_5087,N_4273,N_4859);
or U5088 (N_5088,N_4237,N_4981);
and U5089 (N_5089,N_4086,N_4852);
nand U5090 (N_5090,N_4017,N_4836);
and U5091 (N_5091,N_4542,N_4433);
and U5092 (N_5092,N_4713,N_4672);
and U5093 (N_5093,N_4718,N_4361);
nor U5094 (N_5094,N_4486,N_4932);
nand U5095 (N_5095,N_4671,N_4171);
xnor U5096 (N_5096,N_4166,N_4507);
nor U5097 (N_5097,N_4870,N_4132);
nand U5098 (N_5098,N_4189,N_4375);
nand U5099 (N_5099,N_4118,N_4721);
nor U5100 (N_5100,N_4269,N_4936);
nor U5101 (N_5101,N_4223,N_4457);
nand U5102 (N_5102,N_4532,N_4448);
nor U5103 (N_5103,N_4609,N_4280);
or U5104 (N_5104,N_4168,N_4190);
nand U5105 (N_5105,N_4489,N_4944);
nand U5106 (N_5106,N_4675,N_4679);
or U5107 (N_5107,N_4617,N_4451);
and U5108 (N_5108,N_4364,N_4183);
and U5109 (N_5109,N_4726,N_4082);
nor U5110 (N_5110,N_4245,N_4085);
nand U5111 (N_5111,N_4472,N_4394);
or U5112 (N_5112,N_4480,N_4027);
nor U5113 (N_5113,N_4098,N_4074);
nor U5114 (N_5114,N_4985,N_4922);
nand U5115 (N_5115,N_4076,N_4178);
and U5116 (N_5116,N_4150,N_4868);
and U5117 (N_5117,N_4476,N_4716);
nand U5118 (N_5118,N_4965,N_4539);
and U5119 (N_5119,N_4554,N_4136);
nand U5120 (N_5120,N_4752,N_4127);
nand U5121 (N_5121,N_4159,N_4415);
and U5122 (N_5122,N_4673,N_4075);
or U5123 (N_5123,N_4099,N_4222);
and U5124 (N_5124,N_4815,N_4212);
nor U5125 (N_5125,N_4840,N_4144);
nor U5126 (N_5126,N_4482,N_4061);
and U5127 (N_5127,N_4941,N_4348);
or U5128 (N_5128,N_4235,N_4533);
or U5129 (N_5129,N_4408,N_4652);
or U5130 (N_5130,N_4808,N_4124);
nor U5131 (N_5131,N_4937,N_4184);
nor U5132 (N_5132,N_4307,N_4385);
nor U5133 (N_5133,N_4374,N_4210);
nand U5134 (N_5134,N_4107,N_4425);
xnor U5135 (N_5135,N_4736,N_4800);
or U5136 (N_5136,N_4881,N_4767);
or U5137 (N_5137,N_4161,N_4473);
nor U5138 (N_5138,N_4036,N_4565);
nand U5139 (N_5139,N_4856,N_4285);
nand U5140 (N_5140,N_4526,N_4187);
nand U5141 (N_5141,N_4701,N_4830);
nor U5142 (N_5142,N_4125,N_4102);
or U5143 (N_5143,N_4925,N_4106);
and U5144 (N_5144,N_4095,N_4874);
or U5145 (N_5145,N_4275,N_4813);
nor U5146 (N_5146,N_4584,N_4100);
and U5147 (N_5147,N_4663,N_4091);
nand U5148 (N_5148,N_4987,N_4195);
or U5149 (N_5149,N_4126,N_4581);
and U5150 (N_5150,N_4040,N_4308);
and U5151 (N_5151,N_4227,N_4655);
nor U5152 (N_5152,N_4951,N_4059);
nand U5153 (N_5153,N_4751,N_4616);
and U5154 (N_5154,N_4782,N_4685);
and U5155 (N_5155,N_4765,N_4247);
nand U5156 (N_5156,N_4479,N_4717);
nand U5157 (N_5157,N_4645,N_4310);
or U5158 (N_5158,N_4756,N_4683);
nand U5159 (N_5159,N_4676,N_4889);
or U5160 (N_5160,N_4401,N_4305);
and U5161 (N_5161,N_4411,N_4311);
nor U5162 (N_5162,N_4490,N_4968);
nor U5163 (N_5163,N_4427,N_4602);
and U5164 (N_5164,N_4481,N_4780);
nand U5165 (N_5165,N_4153,N_4015);
and U5166 (N_5166,N_4268,N_4535);
xor U5167 (N_5167,N_4694,N_4032);
and U5168 (N_5168,N_4334,N_4705);
and U5169 (N_5169,N_4763,N_4826);
nand U5170 (N_5170,N_4347,N_4594);
and U5171 (N_5171,N_4021,N_4191);
or U5172 (N_5172,N_4790,N_4257);
nor U5173 (N_5173,N_4606,N_4893);
nand U5174 (N_5174,N_4898,N_4240);
nor U5175 (N_5175,N_4097,N_4890);
or U5176 (N_5176,N_4768,N_4366);
and U5177 (N_5177,N_4806,N_4927);
nor U5178 (N_5178,N_4242,N_4909);
nor U5179 (N_5179,N_4510,N_4727);
or U5180 (N_5180,N_4720,N_4811);
nand U5181 (N_5181,N_4033,N_4674);
and U5182 (N_5182,N_4891,N_4271);
nand U5183 (N_5183,N_4279,N_4541);
and U5184 (N_5184,N_4031,N_4046);
and U5185 (N_5185,N_4903,N_4088);
and U5186 (N_5186,N_4452,N_4038);
nand U5187 (N_5187,N_4147,N_4345);
nor U5188 (N_5188,N_4471,N_4410);
or U5189 (N_5189,N_4921,N_4848);
nor U5190 (N_5190,N_4684,N_4405);
and U5191 (N_5191,N_4837,N_4664);
nand U5192 (N_5192,N_4797,N_4207);
nand U5193 (N_5193,N_4591,N_4115);
and U5194 (N_5194,N_4899,N_4559);
nand U5195 (N_5195,N_4587,N_4220);
nand U5196 (N_5196,N_4872,N_4070);
or U5197 (N_5197,N_4895,N_4774);
xnor U5198 (N_5198,N_4502,N_4413);
nand U5199 (N_5199,N_4256,N_4005);
and U5200 (N_5200,N_4969,N_4492);
nor U5201 (N_5201,N_4071,N_4649);
nand U5202 (N_5202,N_4644,N_4824);
nor U5203 (N_5203,N_4162,N_4354);
nor U5204 (N_5204,N_4316,N_4841);
nor U5205 (N_5205,N_4062,N_4704);
and U5206 (N_5206,N_4812,N_4216);
and U5207 (N_5207,N_4450,N_4363);
and U5208 (N_5208,N_4346,N_4509);
or U5209 (N_5209,N_4051,N_4047);
xor U5210 (N_5210,N_4695,N_4322);
nand U5211 (N_5211,N_4145,N_4299);
and U5212 (N_5212,N_4193,N_4853);
nor U5213 (N_5213,N_4700,N_4096);
nor U5214 (N_5214,N_4670,N_4860);
or U5215 (N_5215,N_4615,N_4493);
nor U5216 (N_5216,N_4885,N_4049);
xor U5217 (N_5217,N_4092,N_4180);
nor U5218 (N_5218,N_4887,N_4563);
and U5219 (N_5219,N_4084,N_4155);
and U5220 (N_5220,N_4197,N_4266);
nor U5221 (N_5221,N_4006,N_4417);
nand U5222 (N_5222,N_4972,N_4250);
nand U5223 (N_5223,N_4277,N_4179);
nor U5224 (N_5224,N_4940,N_4192);
nor U5225 (N_5225,N_4231,N_4576);
and U5226 (N_5226,N_4561,N_4697);
nand U5227 (N_5227,N_4983,N_4605);
nand U5228 (N_5228,N_4044,N_4611);
nor U5229 (N_5229,N_4953,N_4123);
nor U5230 (N_5230,N_4436,N_4246);
nor U5231 (N_5231,N_4286,N_4386);
nor U5232 (N_5232,N_4529,N_4573);
nand U5233 (N_5233,N_4357,N_4952);
and U5234 (N_5234,N_4801,N_4208);
nor U5235 (N_5235,N_4788,N_4094);
xor U5236 (N_5236,N_4104,N_4646);
or U5237 (N_5237,N_4588,N_4943);
or U5238 (N_5238,N_4380,N_4988);
or U5239 (N_5239,N_4938,N_4861);
and U5240 (N_5240,N_4064,N_4783);
and U5241 (N_5241,N_4232,N_4263);
or U5242 (N_5242,N_4512,N_4537);
and U5243 (N_5243,N_4011,N_4543);
nor U5244 (N_5244,N_4918,N_4420);
and U5245 (N_5245,N_4278,N_4137);
nor U5246 (N_5246,N_4152,N_4014);
nand U5247 (N_5247,N_4818,N_4467);
or U5248 (N_5248,N_4388,N_4792);
nor U5249 (N_5249,N_4875,N_4117);
or U5250 (N_5250,N_4546,N_4536);
nor U5251 (N_5251,N_4627,N_4461);
nor U5252 (N_5252,N_4570,N_4778);
nand U5253 (N_5253,N_4923,N_4993);
nor U5254 (N_5254,N_4580,N_4202);
nand U5255 (N_5255,N_4234,N_4678);
nor U5256 (N_5256,N_4442,N_4930);
nand U5257 (N_5257,N_4135,N_4498);
nor U5258 (N_5258,N_4749,N_4050);
and U5259 (N_5259,N_4572,N_4484);
xnor U5260 (N_5260,N_4114,N_4379);
or U5261 (N_5261,N_4367,N_4382);
and U5262 (N_5262,N_4920,N_4637);
and U5263 (N_5263,N_4641,N_4666);
nor U5264 (N_5264,N_4912,N_4209);
and U5265 (N_5265,N_4775,N_4113);
nand U5266 (N_5266,N_4186,N_4544);
and U5267 (N_5267,N_4931,N_4283);
or U5268 (N_5268,N_4562,N_4873);
nor U5269 (N_5269,N_4120,N_4986);
nand U5270 (N_5270,N_4996,N_4624);
or U5271 (N_5271,N_4555,N_4667);
and U5272 (N_5272,N_4383,N_4613);
nor U5273 (N_5273,N_4827,N_4514);
nor U5274 (N_5274,N_4239,N_4665);
and U5275 (N_5275,N_4945,N_4995);
nor U5276 (N_5276,N_4904,N_4843);
and U5277 (N_5277,N_4387,N_4934);
and U5278 (N_5278,N_4475,N_4002);
and U5279 (N_5279,N_4948,N_4804);
and U5280 (N_5280,N_4648,N_4897);
or U5281 (N_5281,N_4863,N_4052);
and U5282 (N_5282,N_4518,N_4371);
or U5283 (N_5283,N_4435,N_4946);
nand U5284 (N_5284,N_4787,N_4845);
and U5285 (N_5285,N_4355,N_4200);
nand U5286 (N_5286,N_4933,N_4111);
and U5287 (N_5287,N_4729,N_4377);
and U5288 (N_5288,N_4525,N_4838);
and U5289 (N_5289,N_4400,N_4434);
nor U5290 (N_5290,N_4760,N_4503);
nor U5291 (N_5291,N_4198,N_4950);
nor U5292 (N_5292,N_4217,N_4314);
or U5293 (N_5293,N_4693,N_4016);
nand U5294 (N_5294,N_4723,N_4956);
or U5295 (N_5295,N_4298,N_4236);
and U5296 (N_5296,N_4039,N_4776);
and U5297 (N_5297,N_4037,N_4360);
nand U5298 (N_5298,N_4024,N_4876);
nor U5299 (N_5299,N_4571,N_4449);
or U5300 (N_5300,N_4221,N_4604);
xor U5301 (N_5301,N_4372,N_4073);
nor U5302 (N_5302,N_4112,N_4158);
nand U5303 (N_5303,N_4205,N_4739);
nor U5304 (N_5304,N_4724,N_4228);
and U5305 (N_5305,N_4326,N_4689);
or U5306 (N_5306,N_4970,N_4130);
nand U5307 (N_5307,N_4214,N_4569);
or U5308 (N_5308,N_4317,N_4579);
or U5309 (N_5309,N_4151,N_4916);
or U5310 (N_5310,N_4917,N_4659);
nand U5311 (N_5311,N_4867,N_4176);
nand U5312 (N_5312,N_4600,N_4055);
xor U5313 (N_5313,N_4984,N_4786);
or U5314 (N_5314,N_4842,N_4156);
nand U5315 (N_5315,N_4878,N_4902);
nor U5316 (N_5316,N_4201,N_4438);
nand U5317 (N_5317,N_4203,N_4687);
nor U5318 (N_5318,N_4105,N_4248);
nand U5319 (N_5319,N_4034,N_4798);
nand U5320 (N_5320,N_4582,N_4982);
nand U5321 (N_5321,N_4742,N_4358);
nand U5322 (N_5322,N_4880,N_4487);
nand U5323 (N_5323,N_4063,N_4743);
and U5324 (N_5324,N_4947,N_4858);
nand U5325 (N_5325,N_4141,N_4333);
nand U5326 (N_5326,N_4423,N_4003);
nand U5327 (N_5327,N_4900,N_4381);
or U5328 (N_5328,N_4241,N_4636);
nor U5329 (N_5329,N_4350,N_4294);
and U5330 (N_5330,N_4747,N_4690);
and U5331 (N_5331,N_4337,N_4807);
nand U5332 (N_5332,N_4352,N_4353);
nand U5333 (N_5333,N_4719,N_4419);
or U5334 (N_5334,N_4772,N_4816);
or U5335 (N_5335,N_4833,N_4548);
or U5336 (N_5336,N_4012,N_4601);
and U5337 (N_5337,N_4390,N_4458);
nor U5338 (N_5338,N_4160,N_4459);
nand U5339 (N_5339,N_4971,N_4991);
nand U5340 (N_5340,N_4500,N_4722);
and U5341 (N_5341,N_4809,N_4595);
or U5342 (N_5342,N_4619,N_4929);
xor U5343 (N_5343,N_4564,N_4825);
nor U5344 (N_5344,N_4211,N_4740);
or U5345 (N_5345,N_4478,N_4440);
nand U5346 (N_5346,N_4657,N_4737);
nand U5347 (N_5347,N_4276,N_4688);
nand U5348 (N_5348,N_4129,N_4181);
xnor U5349 (N_5349,N_4079,N_4709);
or U5350 (N_5350,N_4730,N_4428);
nor U5351 (N_5351,N_4669,N_4376);
nor U5352 (N_5352,N_4989,N_4850);
or U5353 (N_5353,N_4831,N_4957);
or U5354 (N_5354,N_4586,N_4528);
nor U5355 (N_5355,N_4154,N_4901);
nor U5356 (N_5356,N_4520,N_4629);
nor U5357 (N_5357,N_4254,N_4928);
xor U5358 (N_5358,N_4465,N_4779);
or U5359 (N_5359,N_4866,N_4877);
nand U5360 (N_5360,N_4335,N_4499);
or U5361 (N_5361,N_4626,N_4777);
and U5362 (N_5362,N_4703,N_4662);
nor U5363 (N_5363,N_4409,N_4612);
nor U5364 (N_5364,N_4384,N_4393);
nand U5365 (N_5365,N_4149,N_4578);
or U5366 (N_5366,N_4942,N_4924);
nand U5367 (N_5367,N_4226,N_4090);
and U5368 (N_5368,N_4163,N_4177);
or U5369 (N_5369,N_4549,N_4598);
and U5370 (N_5370,N_4157,N_4023);
nor U5371 (N_5371,N_4233,N_4992);
nand U5372 (N_5372,N_4653,N_4770);
nand U5373 (N_5373,N_4819,N_4359);
nand U5374 (N_5374,N_4185,N_4910);
nand U5375 (N_5375,N_4976,N_4505);
nand U5376 (N_5376,N_4119,N_4599);
and U5377 (N_5377,N_4677,N_4284);
or U5378 (N_5378,N_4835,N_4974);
nor U5379 (N_5379,N_4395,N_4496);
nand U5380 (N_5380,N_4253,N_4583);
nand U5381 (N_5381,N_4712,N_4632);
nand U5382 (N_5382,N_4622,N_4628);
xnor U5383 (N_5383,N_4911,N_4103);
or U5384 (N_5384,N_4834,N_4441);
and U5385 (N_5385,N_4304,N_4643);
or U5386 (N_5386,N_4058,N_4437);
nand U5387 (N_5387,N_4785,N_4485);
nor U5388 (N_5388,N_4962,N_4378);
nor U5389 (N_5389,N_4630,N_4699);
or U5390 (N_5390,N_4980,N_4864);
nand U5391 (N_5391,N_4238,N_4855);
or U5392 (N_5392,N_4025,N_4759);
or U5393 (N_5393,N_4080,N_4754);
and U5394 (N_5394,N_4823,N_4963);
and U5395 (N_5395,N_4914,N_4001);
nor U5396 (N_5396,N_4865,N_4139);
and U5397 (N_5397,N_4443,N_4429);
nor U5398 (N_5398,N_4309,N_4654);
nand U5399 (N_5399,N_4623,N_4165);
or U5400 (N_5400,N_4803,N_4101);
or U5401 (N_5401,N_4999,N_4204);
nor U5402 (N_5402,N_4344,N_4324);
or U5403 (N_5403,N_4416,N_4164);
or U5404 (N_5404,N_4022,N_4820);
nor U5405 (N_5405,N_4466,N_4994);
nor U5406 (N_5406,N_4009,N_4692);
nor U5407 (N_5407,N_4547,N_4534);
or U5408 (N_5408,N_4244,N_4634);
and U5409 (N_5409,N_4464,N_4884);
or U5410 (N_5410,N_4065,N_4590);
nand U5411 (N_5411,N_4597,N_4869);
nor U5412 (N_5412,N_4545,N_4575);
nand U5413 (N_5413,N_4267,N_4320);
or U5414 (N_5414,N_4093,N_4926);
nor U5415 (N_5415,N_4030,N_4894);
nand U5416 (N_5416,N_4495,N_4356);
and U5417 (N_5417,N_4973,N_4173);
or U5418 (N_5418,N_4249,N_4243);
and U5419 (N_5419,N_4550,N_4871);
nor U5420 (N_5420,N_4391,N_4725);
and U5421 (N_5421,N_4262,N_4886);
or U5422 (N_5422,N_4757,N_4817);
and U5423 (N_5423,N_4230,N_4219);
nand U5424 (N_5424,N_4516,N_4331);
nor U5425 (N_5425,N_4013,N_4961);
and U5426 (N_5426,N_4424,N_4519);
nand U5427 (N_5427,N_4511,N_4288);
nor U5428 (N_5428,N_4585,N_4796);
and U5429 (N_5429,N_4919,N_4967);
nand U5430 (N_5430,N_4421,N_4000);
nand U5431 (N_5431,N_4748,N_4755);
or U5432 (N_5432,N_4608,N_4477);
and U5433 (N_5433,N_4618,N_4293);
or U5434 (N_5434,N_4218,N_4089);
and U5435 (N_5435,N_4888,N_4043);
or U5436 (N_5436,N_4766,N_4710);
nor U5437 (N_5437,N_4252,N_4761);
or U5438 (N_5438,N_4083,N_4121);
nor U5439 (N_5439,N_4321,N_4862);
nand U5440 (N_5440,N_4224,N_4373);
nand U5441 (N_5441,N_4795,N_4110);
and U5442 (N_5442,N_4462,N_4140);
and U5443 (N_5443,N_4521,N_4589);
or U5444 (N_5444,N_4167,N_4530);
or U5445 (N_5445,N_4323,N_4422);
and U5446 (N_5446,N_4215,N_4527);
and U5447 (N_5447,N_4259,N_4265);
nor U5448 (N_5448,N_4170,N_4997);
nand U5449 (N_5449,N_4508,N_4053);
and U5450 (N_5450,N_4291,N_4341);
and U5451 (N_5451,N_4635,N_4447);
nor U5452 (N_5452,N_4764,N_4698);
or U5453 (N_5453,N_4488,N_4454);
or U5454 (N_5454,N_4882,N_4407);
and U5455 (N_5455,N_4007,N_4781);
nand U5456 (N_5456,N_4116,N_4060);
and U5457 (N_5457,N_4225,N_4793);
or U5458 (N_5458,N_4738,N_4260);
nand U5459 (N_5459,N_4004,N_4339);
and U5460 (N_5460,N_4453,N_4577);
nand U5461 (N_5461,N_4998,N_4229);
or U5462 (N_5462,N_4491,N_4964);
nor U5463 (N_5463,N_4296,N_4504);
or U5464 (N_5464,N_4045,N_4327);
nor U5465 (N_5465,N_4325,N_4762);
or U5466 (N_5466,N_4412,N_4603);
nor U5467 (N_5467,N_4814,N_4702);
nor U5468 (N_5468,N_4607,N_4143);
or U5469 (N_5469,N_4879,N_4303);
nand U5470 (N_5470,N_4896,N_4552);
or U5471 (N_5471,N_4728,N_4041);
nor U5472 (N_5472,N_4048,N_4010);
nor U5473 (N_5473,N_4468,N_4773);
and U5474 (N_5474,N_4431,N_4959);
xnor U5475 (N_5475,N_4315,N_4172);
or U5476 (N_5476,N_4822,N_4264);
nand U5477 (N_5477,N_4336,N_4913);
xnor U5478 (N_5478,N_4261,N_4418);
and U5479 (N_5479,N_4960,N_4746);
nor U5480 (N_5480,N_4078,N_4398);
and U5481 (N_5481,N_4402,N_4515);
or U5482 (N_5482,N_4810,N_4188);
and U5483 (N_5483,N_4567,N_4731);
and U5484 (N_5484,N_4469,N_4631);
nor U5485 (N_5485,N_4857,N_4707);
nor U5486 (N_5486,N_4370,N_4620);
and U5487 (N_5487,N_4035,N_4802);
or U5488 (N_5488,N_4531,N_4169);
or U5489 (N_5489,N_4633,N_4784);
and U5490 (N_5490,N_4365,N_4054);
and U5491 (N_5491,N_4844,N_4791);
nand U5492 (N_5492,N_4691,N_4799);
nand U5493 (N_5493,N_4769,N_4758);
or U5494 (N_5494,N_4596,N_4108);
nand U5495 (N_5495,N_4318,N_4954);
and U5496 (N_5496,N_4513,N_4430);
and U5497 (N_5497,N_4057,N_4404);
nor U5498 (N_5498,N_4340,N_4706);
and U5499 (N_5499,N_4403,N_4558);
or U5500 (N_5500,N_4135,N_4506);
nand U5501 (N_5501,N_4097,N_4689);
nand U5502 (N_5502,N_4468,N_4177);
or U5503 (N_5503,N_4610,N_4845);
xor U5504 (N_5504,N_4343,N_4930);
nor U5505 (N_5505,N_4575,N_4335);
or U5506 (N_5506,N_4657,N_4669);
and U5507 (N_5507,N_4313,N_4445);
and U5508 (N_5508,N_4321,N_4612);
or U5509 (N_5509,N_4267,N_4107);
or U5510 (N_5510,N_4717,N_4776);
and U5511 (N_5511,N_4661,N_4927);
or U5512 (N_5512,N_4955,N_4858);
or U5513 (N_5513,N_4100,N_4866);
nand U5514 (N_5514,N_4644,N_4892);
and U5515 (N_5515,N_4700,N_4457);
or U5516 (N_5516,N_4619,N_4748);
and U5517 (N_5517,N_4360,N_4944);
and U5518 (N_5518,N_4909,N_4865);
nand U5519 (N_5519,N_4631,N_4365);
nor U5520 (N_5520,N_4095,N_4890);
nand U5521 (N_5521,N_4533,N_4972);
or U5522 (N_5522,N_4845,N_4311);
and U5523 (N_5523,N_4588,N_4673);
nand U5524 (N_5524,N_4463,N_4582);
or U5525 (N_5525,N_4743,N_4704);
or U5526 (N_5526,N_4226,N_4548);
or U5527 (N_5527,N_4203,N_4374);
nor U5528 (N_5528,N_4308,N_4428);
and U5529 (N_5529,N_4286,N_4501);
nor U5530 (N_5530,N_4570,N_4994);
or U5531 (N_5531,N_4005,N_4699);
nor U5532 (N_5532,N_4195,N_4393);
nor U5533 (N_5533,N_4105,N_4522);
nand U5534 (N_5534,N_4088,N_4833);
nand U5535 (N_5535,N_4036,N_4393);
or U5536 (N_5536,N_4876,N_4124);
nand U5537 (N_5537,N_4739,N_4126);
and U5538 (N_5538,N_4608,N_4837);
nor U5539 (N_5539,N_4571,N_4480);
nor U5540 (N_5540,N_4304,N_4586);
nor U5541 (N_5541,N_4404,N_4555);
nor U5542 (N_5542,N_4666,N_4639);
nor U5543 (N_5543,N_4823,N_4504);
nor U5544 (N_5544,N_4125,N_4533);
or U5545 (N_5545,N_4311,N_4550);
nor U5546 (N_5546,N_4403,N_4711);
and U5547 (N_5547,N_4637,N_4592);
and U5548 (N_5548,N_4095,N_4360);
or U5549 (N_5549,N_4538,N_4379);
nand U5550 (N_5550,N_4585,N_4091);
and U5551 (N_5551,N_4370,N_4042);
and U5552 (N_5552,N_4977,N_4358);
nand U5553 (N_5553,N_4224,N_4209);
nor U5554 (N_5554,N_4183,N_4124);
xor U5555 (N_5555,N_4153,N_4097);
or U5556 (N_5556,N_4653,N_4550);
nor U5557 (N_5557,N_4796,N_4705);
nand U5558 (N_5558,N_4934,N_4514);
nand U5559 (N_5559,N_4551,N_4975);
and U5560 (N_5560,N_4770,N_4585);
and U5561 (N_5561,N_4311,N_4431);
and U5562 (N_5562,N_4579,N_4861);
xnor U5563 (N_5563,N_4197,N_4876);
or U5564 (N_5564,N_4822,N_4578);
nand U5565 (N_5565,N_4742,N_4613);
nand U5566 (N_5566,N_4856,N_4600);
or U5567 (N_5567,N_4615,N_4048);
or U5568 (N_5568,N_4389,N_4540);
nand U5569 (N_5569,N_4222,N_4130);
nor U5570 (N_5570,N_4354,N_4487);
or U5571 (N_5571,N_4417,N_4404);
and U5572 (N_5572,N_4037,N_4960);
nor U5573 (N_5573,N_4695,N_4841);
nand U5574 (N_5574,N_4152,N_4651);
or U5575 (N_5575,N_4845,N_4196);
nand U5576 (N_5576,N_4047,N_4826);
and U5577 (N_5577,N_4817,N_4418);
nand U5578 (N_5578,N_4949,N_4989);
or U5579 (N_5579,N_4947,N_4927);
nor U5580 (N_5580,N_4978,N_4199);
or U5581 (N_5581,N_4830,N_4048);
nor U5582 (N_5582,N_4857,N_4209);
and U5583 (N_5583,N_4716,N_4339);
nor U5584 (N_5584,N_4590,N_4863);
or U5585 (N_5585,N_4386,N_4274);
nand U5586 (N_5586,N_4454,N_4194);
or U5587 (N_5587,N_4075,N_4821);
nand U5588 (N_5588,N_4410,N_4718);
nor U5589 (N_5589,N_4259,N_4075);
nand U5590 (N_5590,N_4096,N_4552);
nor U5591 (N_5591,N_4488,N_4037);
or U5592 (N_5592,N_4484,N_4777);
nand U5593 (N_5593,N_4823,N_4972);
or U5594 (N_5594,N_4017,N_4021);
nand U5595 (N_5595,N_4699,N_4979);
and U5596 (N_5596,N_4776,N_4549);
nand U5597 (N_5597,N_4028,N_4528);
nand U5598 (N_5598,N_4278,N_4054);
and U5599 (N_5599,N_4637,N_4386);
nand U5600 (N_5600,N_4864,N_4708);
nor U5601 (N_5601,N_4459,N_4238);
and U5602 (N_5602,N_4917,N_4262);
and U5603 (N_5603,N_4262,N_4656);
nand U5604 (N_5604,N_4692,N_4170);
nand U5605 (N_5605,N_4710,N_4173);
xnor U5606 (N_5606,N_4659,N_4069);
nand U5607 (N_5607,N_4101,N_4635);
nor U5608 (N_5608,N_4806,N_4333);
nand U5609 (N_5609,N_4938,N_4063);
nor U5610 (N_5610,N_4010,N_4353);
nand U5611 (N_5611,N_4629,N_4823);
xnor U5612 (N_5612,N_4471,N_4396);
or U5613 (N_5613,N_4172,N_4893);
and U5614 (N_5614,N_4317,N_4101);
and U5615 (N_5615,N_4151,N_4098);
or U5616 (N_5616,N_4069,N_4284);
nor U5617 (N_5617,N_4012,N_4071);
nor U5618 (N_5618,N_4071,N_4025);
or U5619 (N_5619,N_4297,N_4120);
nand U5620 (N_5620,N_4843,N_4416);
xnor U5621 (N_5621,N_4088,N_4406);
and U5622 (N_5622,N_4757,N_4069);
xnor U5623 (N_5623,N_4317,N_4485);
or U5624 (N_5624,N_4080,N_4108);
nand U5625 (N_5625,N_4398,N_4582);
or U5626 (N_5626,N_4540,N_4768);
or U5627 (N_5627,N_4680,N_4365);
or U5628 (N_5628,N_4395,N_4471);
and U5629 (N_5629,N_4184,N_4725);
nor U5630 (N_5630,N_4064,N_4315);
nand U5631 (N_5631,N_4532,N_4615);
nor U5632 (N_5632,N_4492,N_4641);
and U5633 (N_5633,N_4316,N_4697);
nor U5634 (N_5634,N_4787,N_4321);
and U5635 (N_5635,N_4334,N_4907);
or U5636 (N_5636,N_4128,N_4332);
and U5637 (N_5637,N_4667,N_4009);
or U5638 (N_5638,N_4213,N_4230);
nor U5639 (N_5639,N_4640,N_4568);
nand U5640 (N_5640,N_4102,N_4219);
xor U5641 (N_5641,N_4105,N_4983);
or U5642 (N_5642,N_4298,N_4579);
nor U5643 (N_5643,N_4481,N_4604);
or U5644 (N_5644,N_4380,N_4688);
or U5645 (N_5645,N_4917,N_4312);
and U5646 (N_5646,N_4450,N_4271);
or U5647 (N_5647,N_4324,N_4034);
nand U5648 (N_5648,N_4401,N_4377);
and U5649 (N_5649,N_4424,N_4103);
nor U5650 (N_5650,N_4063,N_4147);
xor U5651 (N_5651,N_4160,N_4885);
nor U5652 (N_5652,N_4726,N_4483);
and U5653 (N_5653,N_4336,N_4170);
and U5654 (N_5654,N_4436,N_4252);
or U5655 (N_5655,N_4001,N_4806);
and U5656 (N_5656,N_4619,N_4241);
nand U5657 (N_5657,N_4984,N_4787);
nor U5658 (N_5658,N_4918,N_4368);
xnor U5659 (N_5659,N_4314,N_4570);
and U5660 (N_5660,N_4005,N_4997);
or U5661 (N_5661,N_4536,N_4881);
nand U5662 (N_5662,N_4499,N_4905);
nand U5663 (N_5663,N_4422,N_4072);
nand U5664 (N_5664,N_4153,N_4735);
nor U5665 (N_5665,N_4843,N_4845);
or U5666 (N_5666,N_4326,N_4710);
and U5667 (N_5667,N_4288,N_4296);
and U5668 (N_5668,N_4445,N_4161);
nand U5669 (N_5669,N_4853,N_4160);
nand U5670 (N_5670,N_4117,N_4676);
and U5671 (N_5671,N_4935,N_4855);
nor U5672 (N_5672,N_4859,N_4942);
nor U5673 (N_5673,N_4267,N_4272);
and U5674 (N_5674,N_4898,N_4906);
or U5675 (N_5675,N_4302,N_4650);
and U5676 (N_5676,N_4737,N_4064);
or U5677 (N_5677,N_4046,N_4689);
nor U5678 (N_5678,N_4832,N_4187);
nor U5679 (N_5679,N_4913,N_4717);
and U5680 (N_5680,N_4172,N_4699);
and U5681 (N_5681,N_4794,N_4404);
nor U5682 (N_5682,N_4759,N_4076);
and U5683 (N_5683,N_4396,N_4817);
or U5684 (N_5684,N_4438,N_4094);
nand U5685 (N_5685,N_4274,N_4473);
and U5686 (N_5686,N_4162,N_4061);
and U5687 (N_5687,N_4928,N_4267);
nor U5688 (N_5688,N_4663,N_4871);
or U5689 (N_5689,N_4739,N_4961);
nand U5690 (N_5690,N_4472,N_4258);
and U5691 (N_5691,N_4812,N_4447);
nand U5692 (N_5692,N_4968,N_4149);
nor U5693 (N_5693,N_4360,N_4119);
or U5694 (N_5694,N_4982,N_4940);
and U5695 (N_5695,N_4611,N_4853);
nor U5696 (N_5696,N_4518,N_4731);
or U5697 (N_5697,N_4112,N_4725);
or U5698 (N_5698,N_4862,N_4890);
and U5699 (N_5699,N_4863,N_4346);
nand U5700 (N_5700,N_4178,N_4292);
nand U5701 (N_5701,N_4155,N_4426);
or U5702 (N_5702,N_4919,N_4063);
and U5703 (N_5703,N_4840,N_4972);
or U5704 (N_5704,N_4106,N_4439);
or U5705 (N_5705,N_4994,N_4364);
and U5706 (N_5706,N_4963,N_4956);
nand U5707 (N_5707,N_4482,N_4744);
nor U5708 (N_5708,N_4837,N_4062);
nor U5709 (N_5709,N_4174,N_4311);
or U5710 (N_5710,N_4637,N_4340);
nor U5711 (N_5711,N_4724,N_4783);
nor U5712 (N_5712,N_4086,N_4975);
and U5713 (N_5713,N_4106,N_4550);
and U5714 (N_5714,N_4910,N_4092);
and U5715 (N_5715,N_4012,N_4715);
or U5716 (N_5716,N_4095,N_4877);
nand U5717 (N_5717,N_4159,N_4588);
or U5718 (N_5718,N_4229,N_4469);
or U5719 (N_5719,N_4704,N_4945);
or U5720 (N_5720,N_4762,N_4656);
or U5721 (N_5721,N_4125,N_4397);
nand U5722 (N_5722,N_4340,N_4468);
nand U5723 (N_5723,N_4747,N_4336);
nor U5724 (N_5724,N_4710,N_4972);
nor U5725 (N_5725,N_4981,N_4906);
nor U5726 (N_5726,N_4395,N_4986);
nor U5727 (N_5727,N_4081,N_4177);
or U5728 (N_5728,N_4805,N_4364);
or U5729 (N_5729,N_4999,N_4285);
nand U5730 (N_5730,N_4123,N_4896);
or U5731 (N_5731,N_4990,N_4203);
or U5732 (N_5732,N_4901,N_4701);
nor U5733 (N_5733,N_4948,N_4955);
nand U5734 (N_5734,N_4847,N_4944);
or U5735 (N_5735,N_4848,N_4871);
and U5736 (N_5736,N_4154,N_4739);
nor U5737 (N_5737,N_4862,N_4037);
nor U5738 (N_5738,N_4261,N_4776);
nand U5739 (N_5739,N_4087,N_4441);
nor U5740 (N_5740,N_4513,N_4230);
or U5741 (N_5741,N_4315,N_4124);
nor U5742 (N_5742,N_4728,N_4510);
nor U5743 (N_5743,N_4575,N_4227);
and U5744 (N_5744,N_4740,N_4272);
nand U5745 (N_5745,N_4432,N_4254);
nor U5746 (N_5746,N_4546,N_4790);
nand U5747 (N_5747,N_4139,N_4040);
nand U5748 (N_5748,N_4563,N_4255);
nor U5749 (N_5749,N_4605,N_4640);
and U5750 (N_5750,N_4358,N_4411);
nor U5751 (N_5751,N_4499,N_4234);
and U5752 (N_5752,N_4004,N_4599);
and U5753 (N_5753,N_4312,N_4239);
nor U5754 (N_5754,N_4157,N_4237);
nand U5755 (N_5755,N_4979,N_4929);
and U5756 (N_5756,N_4829,N_4422);
nand U5757 (N_5757,N_4226,N_4198);
nor U5758 (N_5758,N_4453,N_4360);
and U5759 (N_5759,N_4503,N_4951);
nand U5760 (N_5760,N_4816,N_4908);
nand U5761 (N_5761,N_4348,N_4966);
nand U5762 (N_5762,N_4823,N_4403);
nor U5763 (N_5763,N_4021,N_4105);
nand U5764 (N_5764,N_4075,N_4596);
nor U5765 (N_5765,N_4093,N_4891);
nand U5766 (N_5766,N_4139,N_4137);
nor U5767 (N_5767,N_4017,N_4343);
nor U5768 (N_5768,N_4907,N_4095);
nand U5769 (N_5769,N_4812,N_4571);
or U5770 (N_5770,N_4258,N_4318);
nand U5771 (N_5771,N_4299,N_4704);
or U5772 (N_5772,N_4531,N_4972);
and U5773 (N_5773,N_4747,N_4549);
or U5774 (N_5774,N_4188,N_4280);
nor U5775 (N_5775,N_4300,N_4466);
nand U5776 (N_5776,N_4920,N_4118);
nor U5777 (N_5777,N_4890,N_4541);
and U5778 (N_5778,N_4666,N_4262);
and U5779 (N_5779,N_4956,N_4265);
and U5780 (N_5780,N_4543,N_4269);
nor U5781 (N_5781,N_4281,N_4750);
nand U5782 (N_5782,N_4894,N_4795);
or U5783 (N_5783,N_4415,N_4946);
nand U5784 (N_5784,N_4895,N_4313);
and U5785 (N_5785,N_4498,N_4281);
nand U5786 (N_5786,N_4253,N_4561);
nand U5787 (N_5787,N_4572,N_4478);
nand U5788 (N_5788,N_4120,N_4716);
nor U5789 (N_5789,N_4381,N_4004);
nand U5790 (N_5790,N_4606,N_4037);
or U5791 (N_5791,N_4061,N_4371);
or U5792 (N_5792,N_4471,N_4450);
and U5793 (N_5793,N_4845,N_4147);
or U5794 (N_5794,N_4348,N_4157);
nand U5795 (N_5795,N_4332,N_4162);
nand U5796 (N_5796,N_4447,N_4275);
nor U5797 (N_5797,N_4488,N_4844);
or U5798 (N_5798,N_4695,N_4079);
and U5799 (N_5799,N_4641,N_4357);
and U5800 (N_5800,N_4576,N_4195);
and U5801 (N_5801,N_4413,N_4806);
nand U5802 (N_5802,N_4292,N_4184);
and U5803 (N_5803,N_4922,N_4915);
nand U5804 (N_5804,N_4226,N_4565);
and U5805 (N_5805,N_4657,N_4871);
and U5806 (N_5806,N_4885,N_4264);
nor U5807 (N_5807,N_4994,N_4265);
nand U5808 (N_5808,N_4579,N_4726);
and U5809 (N_5809,N_4688,N_4137);
or U5810 (N_5810,N_4661,N_4411);
nor U5811 (N_5811,N_4399,N_4580);
nand U5812 (N_5812,N_4907,N_4969);
or U5813 (N_5813,N_4762,N_4563);
and U5814 (N_5814,N_4890,N_4850);
or U5815 (N_5815,N_4426,N_4709);
nor U5816 (N_5816,N_4586,N_4300);
nor U5817 (N_5817,N_4346,N_4292);
or U5818 (N_5818,N_4220,N_4050);
and U5819 (N_5819,N_4827,N_4485);
nor U5820 (N_5820,N_4117,N_4942);
and U5821 (N_5821,N_4304,N_4431);
nor U5822 (N_5822,N_4735,N_4824);
nor U5823 (N_5823,N_4555,N_4820);
and U5824 (N_5824,N_4440,N_4383);
nand U5825 (N_5825,N_4772,N_4208);
nor U5826 (N_5826,N_4918,N_4529);
nor U5827 (N_5827,N_4860,N_4754);
and U5828 (N_5828,N_4308,N_4301);
and U5829 (N_5829,N_4676,N_4069);
or U5830 (N_5830,N_4796,N_4828);
nor U5831 (N_5831,N_4867,N_4746);
nand U5832 (N_5832,N_4712,N_4746);
nor U5833 (N_5833,N_4177,N_4941);
nand U5834 (N_5834,N_4053,N_4622);
and U5835 (N_5835,N_4163,N_4994);
or U5836 (N_5836,N_4465,N_4706);
or U5837 (N_5837,N_4099,N_4045);
nand U5838 (N_5838,N_4095,N_4864);
or U5839 (N_5839,N_4279,N_4186);
nand U5840 (N_5840,N_4167,N_4042);
nand U5841 (N_5841,N_4075,N_4704);
or U5842 (N_5842,N_4652,N_4467);
and U5843 (N_5843,N_4534,N_4191);
nor U5844 (N_5844,N_4361,N_4385);
nand U5845 (N_5845,N_4114,N_4721);
and U5846 (N_5846,N_4668,N_4466);
nand U5847 (N_5847,N_4325,N_4495);
or U5848 (N_5848,N_4920,N_4287);
nor U5849 (N_5849,N_4041,N_4742);
or U5850 (N_5850,N_4376,N_4196);
or U5851 (N_5851,N_4660,N_4037);
nor U5852 (N_5852,N_4783,N_4599);
and U5853 (N_5853,N_4628,N_4485);
and U5854 (N_5854,N_4376,N_4113);
or U5855 (N_5855,N_4475,N_4724);
or U5856 (N_5856,N_4026,N_4458);
xor U5857 (N_5857,N_4397,N_4216);
nand U5858 (N_5858,N_4989,N_4262);
nand U5859 (N_5859,N_4834,N_4493);
nand U5860 (N_5860,N_4968,N_4878);
or U5861 (N_5861,N_4879,N_4556);
xor U5862 (N_5862,N_4892,N_4788);
nor U5863 (N_5863,N_4867,N_4208);
nand U5864 (N_5864,N_4066,N_4179);
nor U5865 (N_5865,N_4326,N_4310);
or U5866 (N_5866,N_4815,N_4884);
and U5867 (N_5867,N_4042,N_4471);
nand U5868 (N_5868,N_4610,N_4293);
and U5869 (N_5869,N_4061,N_4401);
nand U5870 (N_5870,N_4019,N_4000);
nand U5871 (N_5871,N_4827,N_4188);
or U5872 (N_5872,N_4974,N_4563);
nand U5873 (N_5873,N_4098,N_4284);
or U5874 (N_5874,N_4502,N_4934);
nand U5875 (N_5875,N_4372,N_4386);
and U5876 (N_5876,N_4259,N_4593);
and U5877 (N_5877,N_4707,N_4114);
or U5878 (N_5878,N_4461,N_4744);
or U5879 (N_5879,N_4535,N_4704);
and U5880 (N_5880,N_4429,N_4594);
or U5881 (N_5881,N_4017,N_4608);
nor U5882 (N_5882,N_4477,N_4971);
or U5883 (N_5883,N_4154,N_4403);
nand U5884 (N_5884,N_4623,N_4092);
nand U5885 (N_5885,N_4199,N_4936);
and U5886 (N_5886,N_4673,N_4234);
and U5887 (N_5887,N_4967,N_4463);
and U5888 (N_5888,N_4918,N_4430);
and U5889 (N_5889,N_4248,N_4496);
nor U5890 (N_5890,N_4345,N_4172);
and U5891 (N_5891,N_4830,N_4079);
nand U5892 (N_5892,N_4205,N_4231);
nand U5893 (N_5893,N_4398,N_4069);
and U5894 (N_5894,N_4568,N_4807);
and U5895 (N_5895,N_4865,N_4432);
and U5896 (N_5896,N_4056,N_4121);
nand U5897 (N_5897,N_4894,N_4160);
xnor U5898 (N_5898,N_4796,N_4449);
and U5899 (N_5899,N_4352,N_4695);
or U5900 (N_5900,N_4017,N_4066);
xor U5901 (N_5901,N_4631,N_4885);
and U5902 (N_5902,N_4409,N_4470);
or U5903 (N_5903,N_4164,N_4992);
or U5904 (N_5904,N_4752,N_4837);
nand U5905 (N_5905,N_4228,N_4594);
nand U5906 (N_5906,N_4563,N_4571);
or U5907 (N_5907,N_4606,N_4764);
or U5908 (N_5908,N_4613,N_4337);
nor U5909 (N_5909,N_4899,N_4631);
nor U5910 (N_5910,N_4826,N_4676);
and U5911 (N_5911,N_4715,N_4189);
or U5912 (N_5912,N_4305,N_4039);
or U5913 (N_5913,N_4124,N_4607);
nand U5914 (N_5914,N_4156,N_4244);
or U5915 (N_5915,N_4460,N_4121);
and U5916 (N_5916,N_4076,N_4223);
and U5917 (N_5917,N_4519,N_4353);
nor U5918 (N_5918,N_4714,N_4940);
nor U5919 (N_5919,N_4641,N_4700);
nand U5920 (N_5920,N_4984,N_4292);
and U5921 (N_5921,N_4931,N_4471);
nor U5922 (N_5922,N_4710,N_4667);
or U5923 (N_5923,N_4616,N_4290);
or U5924 (N_5924,N_4945,N_4431);
or U5925 (N_5925,N_4507,N_4834);
or U5926 (N_5926,N_4969,N_4123);
nand U5927 (N_5927,N_4498,N_4126);
nand U5928 (N_5928,N_4452,N_4580);
or U5929 (N_5929,N_4260,N_4580);
and U5930 (N_5930,N_4262,N_4241);
nand U5931 (N_5931,N_4342,N_4670);
and U5932 (N_5932,N_4014,N_4493);
nand U5933 (N_5933,N_4043,N_4823);
or U5934 (N_5934,N_4919,N_4471);
or U5935 (N_5935,N_4956,N_4004);
or U5936 (N_5936,N_4274,N_4812);
nor U5937 (N_5937,N_4553,N_4970);
nor U5938 (N_5938,N_4025,N_4973);
or U5939 (N_5939,N_4824,N_4713);
or U5940 (N_5940,N_4756,N_4025);
nor U5941 (N_5941,N_4398,N_4730);
nor U5942 (N_5942,N_4193,N_4788);
nand U5943 (N_5943,N_4555,N_4387);
and U5944 (N_5944,N_4075,N_4314);
nor U5945 (N_5945,N_4142,N_4551);
nor U5946 (N_5946,N_4346,N_4672);
and U5947 (N_5947,N_4921,N_4624);
or U5948 (N_5948,N_4790,N_4247);
nor U5949 (N_5949,N_4427,N_4399);
nand U5950 (N_5950,N_4155,N_4252);
nand U5951 (N_5951,N_4644,N_4176);
nand U5952 (N_5952,N_4301,N_4313);
nand U5953 (N_5953,N_4609,N_4581);
nor U5954 (N_5954,N_4666,N_4903);
nor U5955 (N_5955,N_4871,N_4690);
and U5956 (N_5956,N_4958,N_4073);
or U5957 (N_5957,N_4911,N_4286);
nand U5958 (N_5958,N_4850,N_4416);
nor U5959 (N_5959,N_4359,N_4705);
nor U5960 (N_5960,N_4040,N_4476);
nand U5961 (N_5961,N_4341,N_4902);
xor U5962 (N_5962,N_4093,N_4876);
or U5963 (N_5963,N_4613,N_4095);
or U5964 (N_5964,N_4497,N_4006);
and U5965 (N_5965,N_4772,N_4992);
and U5966 (N_5966,N_4847,N_4098);
nor U5967 (N_5967,N_4696,N_4644);
and U5968 (N_5968,N_4779,N_4607);
and U5969 (N_5969,N_4893,N_4397);
nor U5970 (N_5970,N_4877,N_4017);
nand U5971 (N_5971,N_4537,N_4652);
or U5972 (N_5972,N_4212,N_4906);
and U5973 (N_5973,N_4017,N_4316);
nand U5974 (N_5974,N_4130,N_4191);
nand U5975 (N_5975,N_4718,N_4878);
and U5976 (N_5976,N_4512,N_4520);
and U5977 (N_5977,N_4916,N_4220);
or U5978 (N_5978,N_4472,N_4974);
and U5979 (N_5979,N_4104,N_4014);
and U5980 (N_5980,N_4963,N_4103);
nand U5981 (N_5981,N_4618,N_4830);
or U5982 (N_5982,N_4508,N_4423);
or U5983 (N_5983,N_4139,N_4427);
and U5984 (N_5984,N_4373,N_4581);
nand U5985 (N_5985,N_4089,N_4903);
and U5986 (N_5986,N_4769,N_4309);
nor U5987 (N_5987,N_4845,N_4222);
and U5988 (N_5988,N_4989,N_4823);
nand U5989 (N_5989,N_4945,N_4446);
nand U5990 (N_5990,N_4268,N_4428);
nor U5991 (N_5991,N_4765,N_4110);
or U5992 (N_5992,N_4348,N_4690);
nor U5993 (N_5993,N_4702,N_4729);
and U5994 (N_5994,N_4135,N_4245);
nand U5995 (N_5995,N_4398,N_4634);
and U5996 (N_5996,N_4400,N_4910);
or U5997 (N_5997,N_4493,N_4094);
nor U5998 (N_5998,N_4114,N_4741);
and U5999 (N_5999,N_4754,N_4135);
or U6000 (N_6000,N_5962,N_5096);
nor U6001 (N_6001,N_5467,N_5732);
nor U6002 (N_6002,N_5813,N_5206);
nand U6003 (N_6003,N_5090,N_5597);
and U6004 (N_6004,N_5110,N_5295);
and U6005 (N_6005,N_5001,N_5869);
and U6006 (N_6006,N_5060,N_5863);
nor U6007 (N_6007,N_5140,N_5483);
nor U6008 (N_6008,N_5851,N_5526);
nor U6009 (N_6009,N_5783,N_5364);
nand U6010 (N_6010,N_5893,N_5336);
xor U6011 (N_6011,N_5472,N_5025);
or U6012 (N_6012,N_5022,N_5565);
and U6013 (N_6013,N_5587,N_5917);
and U6014 (N_6014,N_5256,N_5285);
and U6015 (N_6015,N_5533,N_5991);
and U6016 (N_6016,N_5082,N_5099);
or U6017 (N_6017,N_5998,N_5320);
nand U6018 (N_6018,N_5612,N_5963);
or U6019 (N_6019,N_5831,N_5866);
nor U6020 (N_6020,N_5194,N_5355);
nand U6021 (N_6021,N_5409,N_5663);
and U6022 (N_6022,N_5633,N_5094);
or U6023 (N_6023,N_5154,N_5836);
and U6024 (N_6024,N_5574,N_5267);
or U6025 (N_6025,N_5529,N_5404);
and U6026 (N_6026,N_5426,N_5322);
nor U6027 (N_6027,N_5546,N_5468);
or U6028 (N_6028,N_5938,N_5568);
xor U6029 (N_6029,N_5266,N_5715);
or U6030 (N_6030,N_5375,N_5013);
and U6031 (N_6031,N_5536,N_5006);
nand U6032 (N_6032,N_5593,N_5272);
or U6033 (N_6033,N_5173,N_5770);
nand U6034 (N_6034,N_5990,N_5009);
and U6035 (N_6035,N_5844,N_5523);
nand U6036 (N_6036,N_5245,N_5981);
or U6037 (N_6037,N_5498,N_5682);
or U6038 (N_6038,N_5262,N_5307);
and U6039 (N_6039,N_5547,N_5763);
nand U6040 (N_6040,N_5043,N_5445);
and U6041 (N_6041,N_5065,N_5932);
or U6042 (N_6042,N_5578,N_5122);
and U6043 (N_6043,N_5775,N_5632);
or U6044 (N_6044,N_5270,N_5771);
nand U6045 (N_6045,N_5497,N_5857);
nor U6046 (N_6046,N_5135,N_5902);
or U6047 (N_6047,N_5897,N_5802);
or U6048 (N_6048,N_5238,N_5361);
and U6049 (N_6049,N_5779,N_5579);
nor U6050 (N_6050,N_5225,N_5325);
nand U6051 (N_6051,N_5005,N_5200);
and U6052 (N_6052,N_5317,N_5172);
nor U6053 (N_6053,N_5474,N_5431);
and U6054 (N_6054,N_5812,N_5539);
nor U6055 (N_6055,N_5644,N_5714);
or U6056 (N_6056,N_5552,N_5477);
and U6057 (N_6057,N_5166,N_5427);
and U6058 (N_6058,N_5324,N_5672);
or U6059 (N_6059,N_5739,N_5174);
and U6060 (N_6060,N_5856,N_5374);
nor U6061 (N_6061,N_5789,N_5725);
and U6062 (N_6062,N_5089,N_5456);
nand U6063 (N_6063,N_5551,N_5074);
nand U6064 (N_6064,N_5638,N_5058);
nor U6065 (N_6065,N_5260,N_5649);
nand U6066 (N_6066,N_5391,N_5156);
and U6067 (N_6067,N_5636,N_5011);
nor U6068 (N_6068,N_5274,N_5124);
nor U6069 (N_6069,N_5599,N_5846);
nor U6070 (N_6070,N_5750,N_5507);
or U6071 (N_6071,N_5244,N_5128);
nand U6072 (N_6072,N_5449,N_5240);
or U6073 (N_6073,N_5460,N_5713);
and U6074 (N_6074,N_5101,N_5019);
nor U6075 (N_6075,N_5378,N_5177);
nor U6076 (N_6076,N_5561,N_5567);
nor U6077 (N_6077,N_5222,N_5872);
nor U6078 (N_6078,N_5120,N_5050);
and U6079 (N_6079,N_5386,N_5114);
and U6080 (N_6080,N_5247,N_5424);
and U6081 (N_6081,N_5509,N_5948);
nand U6082 (N_6082,N_5545,N_5937);
nor U6083 (N_6083,N_5898,N_5335);
or U6084 (N_6084,N_5916,N_5326);
nor U6085 (N_6085,N_5493,N_5440);
nand U6086 (N_6086,N_5150,N_5740);
nor U6087 (N_6087,N_5622,N_5719);
and U6088 (N_6088,N_5093,N_5112);
or U6089 (N_6089,N_5959,N_5736);
nand U6090 (N_6090,N_5127,N_5070);
or U6091 (N_6091,N_5115,N_5575);
nor U6092 (N_6092,N_5145,N_5010);
nand U6093 (N_6093,N_5626,N_5590);
nand U6094 (N_6094,N_5665,N_5473);
nand U6095 (N_6095,N_5417,N_5936);
or U6096 (N_6096,N_5447,N_5707);
and U6097 (N_6097,N_5218,N_5454);
or U6098 (N_6098,N_5464,N_5870);
nand U6099 (N_6099,N_5211,N_5492);
and U6100 (N_6100,N_5275,N_5268);
or U6101 (N_6101,N_5412,N_5406);
nor U6102 (N_6102,N_5394,N_5571);
or U6103 (N_6103,N_5624,N_5996);
nor U6104 (N_6104,N_5223,N_5372);
and U6105 (N_6105,N_5731,N_5923);
nor U6106 (N_6106,N_5791,N_5603);
nor U6107 (N_6107,N_5380,N_5111);
nor U6108 (N_6108,N_5634,N_5453);
nand U6109 (N_6109,N_5388,N_5861);
nor U6110 (N_6110,N_5138,N_5490);
xnor U6111 (N_6111,N_5535,N_5919);
nor U6112 (N_6112,N_5697,N_5778);
and U6113 (N_6113,N_5982,N_5927);
and U6114 (N_6114,N_5642,N_5729);
or U6115 (N_6115,N_5879,N_5903);
or U6116 (N_6116,N_5169,N_5734);
or U6117 (N_6117,N_5284,N_5541);
and U6118 (N_6118,N_5198,N_5524);
nor U6119 (N_6119,N_5085,N_5834);
nor U6120 (N_6120,N_5422,N_5349);
nand U6121 (N_6121,N_5181,N_5853);
nand U6122 (N_6122,N_5153,N_5976);
or U6123 (N_6123,N_5365,N_5305);
nor U6124 (N_6124,N_5168,N_5155);
nand U6125 (N_6125,N_5604,N_5024);
or U6126 (N_6126,N_5465,N_5691);
and U6127 (N_6127,N_5721,N_5411);
or U6128 (N_6128,N_5443,N_5588);
and U6129 (N_6129,N_5469,N_5584);
or U6130 (N_6130,N_5766,N_5558);
or U6131 (N_6131,N_5659,N_5647);
and U6132 (N_6132,N_5795,N_5532);
or U6133 (N_6133,N_5147,N_5999);
nor U6134 (N_6134,N_5435,N_5038);
or U6135 (N_6135,N_5773,N_5381);
or U6136 (N_6136,N_5143,N_5723);
or U6137 (N_6137,N_5989,N_5265);
nand U6138 (N_6138,N_5727,N_5818);
nor U6139 (N_6139,N_5918,N_5737);
nand U6140 (N_6140,N_5602,N_5966);
and U6141 (N_6141,N_5967,N_5031);
nor U6142 (N_6142,N_5926,N_5652);
xnor U6143 (N_6143,N_5163,N_5913);
nor U6144 (N_6144,N_5514,N_5690);
and U6145 (N_6145,N_5207,N_5296);
nor U6146 (N_6146,N_5014,N_5048);
or U6147 (N_6147,N_5582,N_5606);
nand U6148 (N_6148,N_5432,N_5824);
xnor U6149 (N_6149,N_5214,N_5939);
nand U6150 (N_6150,N_5975,N_5032);
nand U6151 (N_6151,N_5290,N_5041);
and U6152 (N_6152,N_5392,N_5993);
or U6153 (N_6153,N_5909,N_5685);
and U6154 (N_6154,N_5052,N_5291);
or U6155 (N_6155,N_5534,N_5935);
and U6156 (N_6156,N_5092,N_5072);
nor U6157 (N_6157,N_5666,N_5186);
and U6158 (N_6158,N_5889,N_5835);
xor U6159 (N_6159,N_5189,N_5623);
xor U6160 (N_6160,N_5000,N_5873);
and U6161 (N_6161,N_5984,N_5688);
nor U6162 (N_6162,N_5363,N_5928);
and U6163 (N_6163,N_5312,N_5907);
nor U6164 (N_6164,N_5765,N_5769);
nand U6165 (N_6165,N_5202,N_5680);
nor U6166 (N_6166,N_5040,N_5797);
or U6167 (N_6167,N_5661,N_5875);
and U6168 (N_6168,N_5613,N_5689);
or U6169 (N_6169,N_5656,N_5653);
nor U6170 (N_6170,N_5641,N_5243);
or U6171 (N_6171,N_5973,N_5615);
and U6172 (N_6172,N_5977,N_5420);
nor U6173 (N_6173,N_5607,N_5030);
and U6174 (N_6174,N_5330,N_5985);
nand U6175 (N_6175,N_5357,N_5231);
nand U6176 (N_6176,N_5746,N_5847);
and U6177 (N_6177,N_5530,N_5100);
nor U6178 (N_6178,N_5717,N_5308);
nand U6179 (N_6179,N_5953,N_5187);
nor U6180 (N_6180,N_5199,N_5777);
nand U6181 (N_6181,N_5829,N_5944);
or U6182 (N_6182,N_5792,N_5743);
and U6183 (N_6183,N_5811,N_5033);
or U6184 (N_6184,N_5280,N_5159);
and U6185 (N_6185,N_5531,N_5063);
nand U6186 (N_6186,N_5877,N_5113);
nand U6187 (N_6187,N_5356,N_5387);
or U6188 (N_6188,N_5608,N_5970);
or U6189 (N_6189,N_5807,N_5658);
and U6190 (N_6190,N_5430,N_5854);
and U6191 (N_6191,N_5876,N_5886);
nand U6192 (N_6192,N_5091,N_5620);
or U6193 (N_6193,N_5964,N_5995);
or U6194 (N_6194,N_5972,N_5855);
nor U6195 (N_6195,N_5466,N_5496);
nor U6196 (N_6196,N_5793,N_5782);
or U6197 (N_6197,N_5068,N_5720);
or U6198 (N_6198,N_5784,N_5828);
nor U6199 (N_6199,N_5814,N_5358);
and U6200 (N_6200,N_5583,N_5158);
or U6201 (N_6201,N_5895,N_5415);
nor U6202 (N_6202,N_5816,N_5131);
or U6203 (N_6203,N_5436,N_5328);
nand U6204 (N_6204,N_5752,N_5376);
nand U6205 (N_6205,N_5596,N_5728);
and U6206 (N_6206,N_5294,N_5637);
and U6207 (N_6207,N_5152,N_5373);
and U6208 (N_6208,N_5401,N_5076);
xnor U6209 (N_6209,N_5912,N_5359);
nand U6210 (N_6210,N_5452,N_5544);
and U6211 (N_6211,N_5179,N_5306);
or U6212 (N_6212,N_5180,N_5286);
nand U6213 (N_6213,N_5055,N_5045);
or U6214 (N_6214,N_5852,N_5360);
or U6215 (N_6215,N_5416,N_5762);
and U6216 (N_6216,N_5744,N_5188);
nand U6217 (N_6217,N_5883,N_5119);
and U6218 (N_6218,N_5446,N_5162);
nand U6219 (N_6219,N_5887,N_5192);
or U6220 (N_6220,N_5276,N_5566);
nand U6221 (N_6221,N_5017,N_5670);
nor U6222 (N_6222,N_5340,N_5781);
nand U6223 (N_6223,N_5134,N_5758);
nor U6224 (N_6224,N_5350,N_5301);
and U6225 (N_6225,N_5573,N_5269);
and U6226 (N_6226,N_5890,N_5801);
and U6227 (N_6227,N_5149,N_5339);
nor U6228 (N_6228,N_5865,N_5144);
nor U6229 (N_6229,N_5711,N_5683);
and U6230 (N_6230,N_5064,N_5337);
nand U6231 (N_6231,N_5354,N_5292);
nor U6232 (N_6232,N_5705,N_5920);
nand U6233 (N_6233,N_5706,N_5675);
and U6234 (N_6234,N_5319,N_5095);
nand U6235 (N_6235,N_5018,N_5263);
or U6236 (N_6236,N_5020,N_5968);
and U6237 (N_6237,N_5930,N_5600);
nor U6238 (N_6238,N_5800,N_5756);
or U6239 (N_6239,N_5794,N_5616);
nor U6240 (N_6240,N_5511,N_5686);
or U6241 (N_6241,N_5004,N_5423);
and U6242 (N_6242,N_5694,N_5772);
nor U6243 (N_6243,N_5560,N_5235);
nor U6244 (N_6244,N_5505,N_5542);
nand U6245 (N_6245,N_5517,N_5441);
and U6246 (N_6246,N_5334,N_5488);
nand U6247 (N_6247,N_5830,N_5742);
nand U6248 (N_6248,N_5046,N_5471);
and U6249 (N_6249,N_5790,N_5146);
and U6250 (N_6250,N_5674,N_5611);
or U6251 (N_6251,N_5704,N_5513);
or U6252 (N_6252,N_5595,N_5780);
nor U6253 (N_6253,N_5673,N_5651);
and U6254 (N_6254,N_5321,N_5826);
nand U6255 (N_6255,N_5549,N_5681);
nand U6256 (N_6256,N_5804,N_5958);
nor U6257 (N_6257,N_5080,N_5139);
or U6258 (N_6258,N_5457,N_5589);
nor U6259 (N_6259,N_5298,N_5051);
and U6260 (N_6260,N_5304,N_5132);
nand U6261 (N_6261,N_5580,N_5382);
nand U6262 (N_6262,N_5842,N_5104);
or U6263 (N_6263,N_5859,N_5947);
nor U6264 (N_6264,N_5548,N_5979);
nand U6265 (N_6265,N_5160,N_5397);
and U6266 (N_6266,N_5252,N_5323);
or U6267 (N_6267,N_5103,N_5191);
and U6268 (N_6268,N_5282,N_5485);
or U6269 (N_6269,N_5433,N_5904);
nor U6270 (N_6270,N_5209,N_5369);
nand U6271 (N_6271,N_5664,N_5525);
or U6272 (N_6272,N_5988,N_5712);
nor U6273 (N_6273,N_5254,N_5345);
nor U6274 (N_6274,N_5987,N_5822);
or U6275 (N_6275,N_5757,N_5677);
nor U6276 (N_6276,N_5234,N_5858);
nor U6277 (N_6277,N_5843,N_5475);
nor U6278 (N_6278,N_5484,N_5760);
or U6279 (N_6279,N_5874,N_5621);
nand U6280 (N_6280,N_5910,N_5253);
nand U6281 (N_6281,N_5605,N_5283);
nor U6282 (N_6282,N_5461,N_5724);
nor U6283 (N_6283,N_5562,N_5178);
and U6284 (N_6284,N_5839,N_5954);
nand U6285 (N_6285,N_5796,N_5049);
nand U6286 (N_6286,N_5059,N_5402);
and U6287 (N_6287,N_5219,N_5277);
or U6288 (N_6288,N_5880,N_5487);
or U6289 (N_6289,N_5442,N_5479);
nor U6290 (N_6290,N_5217,N_5311);
nand U6291 (N_6291,N_5184,N_5810);
xor U6292 (N_6292,N_5012,N_5825);
nor U6293 (N_6293,N_5761,N_5577);
nor U6294 (N_6294,N_5494,N_5891);
and U6295 (N_6295,N_5171,N_5458);
nor U6296 (N_6296,N_5210,N_5510);
and U6297 (N_6297,N_5429,N_5300);
or U6298 (N_6298,N_5899,N_5331);
or U6299 (N_6299,N_5808,N_5687);
and U6300 (N_6300,N_5237,N_5806);
nand U6301 (N_6301,N_5655,N_5662);
nor U6302 (N_6302,N_5271,N_5933);
or U6303 (N_6303,N_5708,N_5462);
and U6304 (N_6304,N_5543,N_5915);
nand U6305 (N_6305,N_5035,N_5288);
and U6306 (N_6306,N_5820,N_5819);
and U6307 (N_6307,N_5341,N_5116);
nor U6308 (N_6308,N_5701,N_5229);
and U6309 (N_6309,N_5516,N_5259);
xor U6310 (N_6310,N_5125,N_5213);
nand U6311 (N_6311,N_5108,N_5126);
and U6312 (N_6312,N_5097,N_5654);
and U6313 (N_6313,N_5141,N_5313);
or U6314 (N_6314,N_5678,N_5056);
xnor U6315 (N_6315,N_5619,N_5258);
or U6316 (N_6316,N_5508,N_5618);
xor U6317 (N_6317,N_5684,N_5894);
and U6318 (N_6318,N_5609,N_5502);
and U6319 (N_6319,N_5645,N_5515);
nand U6320 (N_6320,N_5550,N_5992);
and U6321 (N_6321,N_5368,N_5695);
and U6322 (N_6322,N_5246,N_5047);
or U6323 (N_6323,N_5648,N_5592);
or U6324 (N_6324,N_5570,N_5241);
nand U6325 (N_6325,N_5137,N_5860);
nor U6326 (N_6326,N_5956,N_5118);
and U6327 (N_6327,N_5418,N_5183);
and U6328 (N_6328,N_5817,N_5730);
nor U6329 (N_6329,N_5521,N_5053);
nor U6330 (N_6330,N_5370,N_5581);
or U6331 (N_6331,N_5946,N_5986);
nor U6332 (N_6332,N_5278,N_5204);
and U6333 (N_6333,N_5226,N_5212);
xnor U6334 (N_6334,N_5084,N_5832);
nor U6335 (N_6335,N_5671,N_5400);
or U6336 (N_6336,N_5302,N_5315);
and U6337 (N_6337,N_5230,N_5557);
nand U6338 (N_6338,N_5338,N_5698);
and U6339 (N_6339,N_5190,N_5242);
or U6340 (N_6340,N_5668,N_5625);
xnor U6341 (N_6341,N_5841,N_5945);
nor U6342 (N_6342,N_5699,N_5702);
nand U6343 (N_6343,N_5827,N_5983);
nor U6344 (N_6344,N_5438,N_5747);
nor U6345 (N_6345,N_5735,N_5385);
nor U6346 (N_6346,N_5520,N_5384);
nand U6347 (N_6347,N_5940,N_5905);
nand U6348 (N_6348,N_5078,N_5563);
nand U6349 (N_6349,N_5840,N_5161);
or U6350 (N_6350,N_5297,N_5850);
or U6351 (N_6351,N_5054,N_5220);
and U6352 (N_6352,N_5726,N_5885);
and U6353 (N_6353,N_5167,N_5251);
nor U6354 (N_6354,N_5925,N_5203);
nor U6355 (N_6355,N_5518,N_5506);
nor U6356 (N_6356,N_5617,N_5088);
or U6357 (N_6357,N_5281,N_5569);
nor U6358 (N_6358,N_5553,N_5598);
or U6359 (N_6359,N_5540,N_5318);
nor U6360 (N_6360,N_5929,N_5884);
xnor U6361 (N_6361,N_5117,N_5196);
nor U6362 (N_6362,N_5439,N_5257);
or U6363 (N_6363,N_5700,N_5503);
nor U6364 (N_6364,N_5785,N_5057);
and U6365 (N_6365,N_5738,N_5414);
nand U6366 (N_6366,N_5419,N_5428);
or U6367 (N_6367,N_5451,N_5455);
or U6368 (N_6368,N_5942,N_5881);
and U6369 (N_6369,N_5748,N_5718);
nand U6370 (N_6370,N_5314,N_5722);
nor U6371 (N_6371,N_5639,N_5333);
or U6372 (N_6372,N_5878,N_5007);
nor U6373 (N_6373,N_5955,N_5036);
nor U6374 (N_6374,N_5037,N_5175);
xnor U6375 (N_6375,N_5931,N_5197);
and U6376 (N_6376,N_5862,N_5774);
or U6377 (N_6377,N_5823,N_5629);
or U6378 (N_6378,N_5585,N_5768);
and U6379 (N_6379,N_5061,N_5239);
nor U6380 (N_6380,N_5151,N_5463);
nor U6381 (N_6381,N_5555,N_5342);
and U6382 (N_6382,N_5407,N_5969);
and U6383 (N_6383,N_5798,N_5486);
nor U6384 (N_6384,N_5289,N_5805);
or U6385 (N_6385,N_5495,N_5398);
or U6386 (N_6386,N_5709,N_5105);
or U6387 (N_6387,N_5892,N_5107);
nand U6388 (N_6388,N_5299,N_5522);
nor U6389 (N_6389,N_5273,N_5667);
nand U6390 (N_6390,N_5236,N_5248);
and U6391 (N_6391,N_5799,N_5170);
and U6392 (N_6392,N_5952,N_5941);
and U6393 (N_6393,N_5086,N_5023);
xnor U6394 (N_6394,N_5512,N_5650);
nor U6395 (N_6395,N_5176,N_5751);
nand U6396 (N_6396,N_5227,N_5759);
and U6397 (N_6397,N_5003,N_5303);
and U6398 (N_6398,N_5233,N_5501);
nand U6399 (N_6399,N_5838,N_5077);
nor U6400 (N_6400,N_5193,N_5316);
nand U6401 (N_6401,N_5142,N_5293);
or U6402 (N_6402,N_5249,N_5343);
nor U6403 (N_6403,N_5755,N_5106);
nor U6404 (N_6404,N_5255,N_5997);
or U6405 (N_6405,N_5848,N_5026);
or U6406 (N_6406,N_5911,N_5205);
nand U6407 (N_6407,N_5327,N_5310);
nor U6408 (N_6408,N_5410,N_5332);
and U6409 (N_6409,N_5833,N_5027);
and U6410 (N_6410,N_5102,N_5039);
or U6411 (N_6411,N_5676,N_5062);
nor U6412 (N_6412,N_5377,N_5924);
nor U6413 (N_6413,N_5733,N_5346);
nand U6414 (N_6414,N_5906,N_5066);
nand U6415 (N_6415,N_5390,N_5123);
and U6416 (N_6416,N_5264,N_5071);
nor U6417 (N_6417,N_5628,N_5971);
and U6418 (N_6418,N_5476,N_5950);
and U6419 (N_6419,N_5867,N_5081);
and U6420 (N_6420,N_5434,N_5185);
nor U6421 (N_6421,N_5900,N_5934);
or U6422 (N_6422,N_5538,N_5660);
and U6423 (N_6423,N_5627,N_5978);
nor U6424 (N_6424,N_5643,N_5367);
nand U6425 (N_6425,N_5129,N_5396);
nor U6426 (N_6426,N_5073,N_5362);
nand U6427 (N_6427,N_5015,N_5136);
nand U6428 (N_6428,N_5745,N_5692);
nand U6429 (N_6429,N_5527,N_5657);
and U6430 (N_6430,N_5366,N_5504);
xor U6431 (N_6431,N_5753,N_5949);
nor U6432 (N_6432,N_5164,N_5554);
or U6433 (N_6433,N_5425,N_5868);
or U6434 (N_6434,N_5821,N_5403);
and U6435 (N_6435,N_5922,N_5448);
nor U6436 (N_6436,N_5901,N_5491);
nand U6437 (N_6437,N_5499,N_5352);
nor U6438 (N_6438,N_5980,N_5351);
or U6439 (N_6439,N_5576,N_5437);
nand U6440 (N_6440,N_5635,N_5408);
and U6441 (N_6441,N_5087,N_5849);
or U6442 (N_6442,N_5130,N_5481);
and U6443 (N_6443,N_5882,N_5016);
nand U6444 (N_6444,N_5764,N_5480);
nand U6445 (N_6445,N_5109,N_5710);
and U6446 (N_6446,N_5888,N_5845);
nor U6447 (N_6447,N_5224,N_5703);
nand U6448 (N_6448,N_5482,N_5208);
and U6449 (N_6449,N_5896,N_5148);
and U6450 (N_6450,N_5421,N_5250);
and U6451 (N_6451,N_5749,N_5261);
or U6452 (N_6452,N_5914,N_5559);
nor U6453 (N_6453,N_5478,N_5610);
or U6454 (N_6454,N_5353,N_5519);
nor U6455 (N_6455,N_5572,N_5837);
nor U6456 (N_6456,N_5537,N_5067);
and U6457 (N_6457,N_5994,N_5069);
nand U6458 (N_6458,N_5098,N_5871);
or U6459 (N_6459,N_5528,N_5961);
and U6460 (N_6460,N_5008,N_5028);
and U6461 (N_6461,N_5329,N_5309);
nand U6462 (N_6462,N_5614,N_5631);
and U6463 (N_6463,N_5044,N_5232);
nor U6464 (N_6464,N_5383,N_5075);
xnor U6465 (N_6465,N_5201,N_5564);
or U6466 (N_6466,N_5002,N_5228);
or U6467 (N_6467,N_5405,N_5450);
nor U6468 (N_6468,N_5221,N_5741);
nor U6469 (N_6469,N_5630,N_5974);
nand U6470 (N_6470,N_5786,N_5029);
or U6471 (N_6471,N_5470,N_5815);
nand U6472 (N_6472,N_5646,N_5347);
or U6473 (N_6473,N_5165,N_5556);
nor U6474 (N_6474,N_5157,N_5586);
or U6475 (N_6475,N_5444,N_5803);
nor U6476 (N_6476,N_5601,N_5379);
and U6477 (N_6477,N_5216,N_5413);
nand U6478 (N_6478,N_5034,N_5787);
nand U6479 (N_6479,N_5182,N_5348);
nor U6480 (N_6480,N_5669,N_5640);
or U6481 (N_6481,N_5951,N_5594);
and U6482 (N_6482,N_5121,N_5921);
or U6483 (N_6483,N_5776,N_5943);
nand U6484 (N_6484,N_5960,N_5788);
nor U6485 (N_6485,N_5279,N_5399);
and U6486 (N_6486,N_5489,N_5767);
or U6487 (N_6487,N_5908,N_5864);
nor U6488 (N_6488,N_5754,N_5395);
nand U6489 (N_6489,N_5679,N_5965);
nor U6490 (N_6490,N_5389,N_5693);
and U6491 (N_6491,N_5079,N_5393);
nand U6492 (N_6492,N_5215,N_5716);
and U6493 (N_6493,N_5083,N_5021);
or U6494 (N_6494,N_5500,N_5042);
nor U6495 (N_6495,N_5344,N_5459);
nand U6496 (N_6496,N_5195,N_5371);
nor U6497 (N_6497,N_5809,N_5133);
nand U6498 (N_6498,N_5591,N_5957);
nand U6499 (N_6499,N_5696,N_5287);
xnor U6500 (N_6500,N_5428,N_5680);
nor U6501 (N_6501,N_5828,N_5862);
and U6502 (N_6502,N_5373,N_5254);
nand U6503 (N_6503,N_5465,N_5283);
or U6504 (N_6504,N_5241,N_5208);
or U6505 (N_6505,N_5854,N_5398);
nand U6506 (N_6506,N_5173,N_5714);
and U6507 (N_6507,N_5662,N_5407);
nand U6508 (N_6508,N_5723,N_5148);
nand U6509 (N_6509,N_5309,N_5727);
and U6510 (N_6510,N_5357,N_5788);
or U6511 (N_6511,N_5139,N_5097);
nand U6512 (N_6512,N_5338,N_5629);
and U6513 (N_6513,N_5595,N_5739);
and U6514 (N_6514,N_5882,N_5015);
nor U6515 (N_6515,N_5373,N_5037);
or U6516 (N_6516,N_5374,N_5027);
and U6517 (N_6517,N_5144,N_5103);
and U6518 (N_6518,N_5131,N_5721);
or U6519 (N_6519,N_5145,N_5155);
or U6520 (N_6520,N_5188,N_5216);
or U6521 (N_6521,N_5818,N_5824);
nand U6522 (N_6522,N_5087,N_5735);
nor U6523 (N_6523,N_5799,N_5776);
nand U6524 (N_6524,N_5510,N_5085);
or U6525 (N_6525,N_5355,N_5962);
nand U6526 (N_6526,N_5003,N_5379);
or U6527 (N_6527,N_5613,N_5185);
or U6528 (N_6528,N_5278,N_5369);
nor U6529 (N_6529,N_5654,N_5031);
and U6530 (N_6530,N_5648,N_5215);
or U6531 (N_6531,N_5731,N_5065);
or U6532 (N_6532,N_5640,N_5570);
or U6533 (N_6533,N_5905,N_5948);
nor U6534 (N_6534,N_5402,N_5131);
and U6535 (N_6535,N_5627,N_5209);
and U6536 (N_6536,N_5407,N_5022);
nand U6537 (N_6537,N_5182,N_5898);
and U6538 (N_6538,N_5999,N_5909);
and U6539 (N_6539,N_5446,N_5409);
and U6540 (N_6540,N_5540,N_5197);
nand U6541 (N_6541,N_5247,N_5097);
nor U6542 (N_6542,N_5500,N_5398);
nand U6543 (N_6543,N_5495,N_5117);
or U6544 (N_6544,N_5893,N_5375);
or U6545 (N_6545,N_5355,N_5113);
and U6546 (N_6546,N_5967,N_5095);
nand U6547 (N_6547,N_5488,N_5975);
nand U6548 (N_6548,N_5927,N_5769);
nor U6549 (N_6549,N_5799,N_5178);
or U6550 (N_6550,N_5728,N_5696);
and U6551 (N_6551,N_5913,N_5885);
or U6552 (N_6552,N_5918,N_5067);
or U6553 (N_6553,N_5143,N_5885);
nand U6554 (N_6554,N_5958,N_5591);
and U6555 (N_6555,N_5531,N_5913);
xnor U6556 (N_6556,N_5145,N_5454);
and U6557 (N_6557,N_5355,N_5937);
nor U6558 (N_6558,N_5529,N_5708);
and U6559 (N_6559,N_5116,N_5724);
nand U6560 (N_6560,N_5148,N_5545);
or U6561 (N_6561,N_5095,N_5286);
or U6562 (N_6562,N_5350,N_5017);
and U6563 (N_6563,N_5384,N_5756);
or U6564 (N_6564,N_5409,N_5928);
nand U6565 (N_6565,N_5119,N_5024);
and U6566 (N_6566,N_5311,N_5919);
nand U6567 (N_6567,N_5010,N_5132);
and U6568 (N_6568,N_5645,N_5241);
or U6569 (N_6569,N_5796,N_5331);
and U6570 (N_6570,N_5964,N_5080);
or U6571 (N_6571,N_5819,N_5771);
or U6572 (N_6572,N_5207,N_5330);
or U6573 (N_6573,N_5299,N_5147);
nand U6574 (N_6574,N_5273,N_5343);
nand U6575 (N_6575,N_5613,N_5023);
nand U6576 (N_6576,N_5726,N_5514);
or U6577 (N_6577,N_5237,N_5622);
and U6578 (N_6578,N_5315,N_5955);
nor U6579 (N_6579,N_5863,N_5188);
and U6580 (N_6580,N_5091,N_5380);
nand U6581 (N_6581,N_5286,N_5970);
nand U6582 (N_6582,N_5311,N_5041);
and U6583 (N_6583,N_5046,N_5958);
nand U6584 (N_6584,N_5441,N_5209);
and U6585 (N_6585,N_5236,N_5844);
and U6586 (N_6586,N_5249,N_5138);
nor U6587 (N_6587,N_5785,N_5560);
nand U6588 (N_6588,N_5093,N_5685);
or U6589 (N_6589,N_5333,N_5741);
and U6590 (N_6590,N_5879,N_5109);
and U6591 (N_6591,N_5892,N_5967);
nand U6592 (N_6592,N_5776,N_5179);
nand U6593 (N_6593,N_5407,N_5994);
and U6594 (N_6594,N_5439,N_5913);
nor U6595 (N_6595,N_5374,N_5485);
nand U6596 (N_6596,N_5726,N_5047);
or U6597 (N_6597,N_5679,N_5193);
nand U6598 (N_6598,N_5509,N_5546);
or U6599 (N_6599,N_5227,N_5274);
nor U6600 (N_6600,N_5812,N_5059);
and U6601 (N_6601,N_5394,N_5554);
nand U6602 (N_6602,N_5396,N_5861);
and U6603 (N_6603,N_5766,N_5933);
nand U6604 (N_6604,N_5965,N_5126);
nor U6605 (N_6605,N_5765,N_5080);
nand U6606 (N_6606,N_5015,N_5657);
nand U6607 (N_6607,N_5861,N_5865);
and U6608 (N_6608,N_5646,N_5186);
nor U6609 (N_6609,N_5215,N_5822);
nor U6610 (N_6610,N_5775,N_5793);
or U6611 (N_6611,N_5615,N_5579);
nor U6612 (N_6612,N_5097,N_5404);
xnor U6613 (N_6613,N_5915,N_5064);
or U6614 (N_6614,N_5583,N_5453);
and U6615 (N_6615,N_5782,N_5867);
nand U6616 (N_6616,N_5497,N_5773);
or U6617 (N_6617,N_5951,N_5278);
and U6618 (N_6618,N_5623,N_5279);
nor U6619 (N_6619,N_5692,N_5650);
nor U6620 (N_6620,N_5374,N_5385);
and U6621 (N_6621,N_5926,N_5454);
and U6622 (N_6622,N_5279,N_5250);
and U6623 (N_6623,N_5227,N_5771);
and U6624 (N_6624,N_5938,N_5529);
nand U6625 (N_6625,N_5727,N_5659);
and U6626 (N_6626,N_5009,N_5358);
or U6627 (N_6627,N_5281,N_5261);
nor U6628 (N_6628,N_5575,N_5655);
or U6629 (N_6629,N_5952,N_5239);
xor U6630 (N_6630,N_5100,N_5378);
nand U6631 (N_6631,N_5408,N_5714);
nand U6632 (N_6632,N_5313,N_5478);
and U6633 (N_6633,N_5046,N_5686);
nor U6634 (N_6634,N_5117,N_5534);
nor U6635 (N_6635,N_5361,N_5281);
and U6636 (N_6636,N_5737,N_5711);
nand U6637 (N_6637,N_5664,N_5276);
or U6638 (N_6638,N_5462,N_5518);
or U6639 (N_6639,N_5861,N_5115);
or U6640 (N_6640,N_5936,N_5113);
and U6641 (N_6641,N_5013,N_5424);
and U6642 (N_6642,N_5937,N_5542);
nor U6643 (N_6643,N_5872,N_5290);
nand U6644 (N_6644,N_5364,N_5696);
nor U6645 (N_6645,N_5832,N_5248);
nor U6646 (N_6646,N_5678,N_5602);
and U6647 (N_6647,N_5363,N_5533);
nor U6648 (N_6648,N_5235,N_5523);
nand U6649 (N_6649,N_5299,N_5617);
nand U6650 (N_6650,N_5265,N_5547);
nand U6651 (N_6651,N_5524,N_5151);
nor U6652 (N_6652,N_5099,N_5220);
and U6653 (N_6653,N_5936,N_5007);
nand U6654 (N_6654,N_5889,N_5132);
nand U6655 (N_6655,N_5513,N_5157);
nor U6656 (N_6656,N_5543,N_5669);
and U6657 (N_6657,N_5224,N_5001);
nor U6658 (N_6658,N_5086,N_5601);
and U6659 (N_6659,N_5919,N_5541);
nand U6660 (N_6660,N_5995,N_5399);
nor U6661 (N_6661,N_5332,N_5894);
xor U6662 (N_6662,N_5549,N_5599);
or U6663 (N_6663,N_5173,N_5722);
nor U6664 (N_6664,N_5488,N_5154);
or U6665 (N_6665,N_5352,N_5097);
nor U6666 (N_6666,N_5616,N_5908);
xnor U6667 (N_6667,N_5366,N_5699);
or U6668 (N_6668,N_5626,N_5644);
nor U6669 (N_6669,N_5816,N_5504);
and U6670 (N_6670,N_5324,N_5071);
or U6671 (N_6671,N_5178,N_5297);
or U6672 (N_6672,N_5756,N_5481);
and U6673 (N_6673,N_5026,N_5386);
nor U6674 (N_6674,N_5708,N_5936);
nand U6675 (N_6675,N_5872,N_5879);
nand U6676 (N_6676,N_5910,N_5331);
and U6677 (N_6677,N_5778,N_5096);
and U6678 (N_6678,N_5357,N_5198);
nor U6679 (N_6679,N_5022,N_5530);
nand U6680 (N_6680,N_5479,N_5434);
nand U6681 (N_6681,N_5367,N_5206);
nor U6682 (N_6682,N_5890,N_5443);
or U6683 (N_6683,N_5590,N_5505);
or U6684 (N_6684,N_5350,N_5360);
nand U6685 (N_6685,N_5146,N_5228);
nand U6686 (N_6686,N_5606,N_5511);
nand U6687 (N_6687,N_5917,N_5893);
nor U6688 (N_6688,N_5843,N_5063);
or U6689 (N_6689,N_5336,N_5419);
nor U6690 (N_6690,N_5441,N_5526);
and U6691 (N_6691,N_5522,N_5587);
or U6692 (N_6692,N_5156,N_5533);
or U6693 (N_6693,N_5732,N_5017);
nand U6694 (N_6694,N_5110,N_5453);
nand U6695 (N_6695,N_5554,N_5962);
xnor U6696 (N_6696,N_5734,N_5905);
nand U6697 (N_6697,N_5671,N_5052);
or U6698 (N_6698,N_5243,N_5004);
and U6699 (N_6699,N_5235,N_5814);
and U6700 (N_6700,N_5146,N_5898);
or U6701 (N_6701,N_5284,N_5772);
nor U6702 (N_6702,N_5145,N_5150);
nand U6703 (N_6703,N_5347,N_5440);
nor U6704 (N_6704,N_5167,N_5276);
nor U6705 (N_6705,N_5911,N_5530);
nand U6706 (N_6706,N_5523,N_5732);
and U6707 (N_6707,N_5283,N_5607);
nor U6708 (N_6708,N_5993,N_5790);
nand U6709 (N_6709,N_5068,N_5965);
nor U6710 (N_6710,N_5757,N_5121);
and U6711 (N_6711,N_5578,N_5388);
xor U6712 (N_6712,N_5384,N_5067);
nor U6713 (N_6713,N_5792,N_5064);
nand U6714 (N_6714,N_5838,N_5336);
nand U6715 (N_6715,N_5011,N_5746);
and U6716 (N_6716,N_5576,N_5058);
nor U6717 (N_6717,N_5364,N_5531);
or U6718 (N_6718,N_5832,N_5540);
and U6719 (N_6719,N_5312,N_5040);
nand U6720 (N_6720,N_5226,N_5461);
nand U6721 (N_6721,N_5849,N_5713);
nand U6722 (N_6722,N_5019,N_5798);
nand U6723 (N_6723,N_5177,N_5801);
nand U6724 (N_6724,N_5322,N_5861);
and U6725 (N_6725,N_5375,N_5705);
or U6726 (N_6726,N_5986,N_5866);
nand U6727 (N_6727,N_5415,N_5671);
and U6728 (N_6728,N_5563,N_5787);
xnor U6729 (N_6729,N_5743,N_5204);
and U6730 (N_6730,N_5594,N_5798);
nor U6731 (N_6731,N_5383,N_5139);
nand U6732 (N_6732,N_5110,N_5777);
nand U6733 (N_6733,N_5897,N_5508);
or U6734 (N_6734,N_5307,N_5799);
nand U6735 (N_6735,N_5844,N_5144);
nor U6736 (N_6736,N_5428,N_5450);
nand U6737 (N_6737,N_5931,N_5528);
nor U6738 (N_6738,N_5604,N_5453);
nor U6739 (N_6739,N_5913,N_5125);
nor U6740 (N_6740,N_5663,N_5730);
nor U6741 (N_6741,N_5927,N_5491);
nand U6742 (N_6742,N_5144,N_5203);
nor U6743 (N_6743,N_5415,N_5770);
nor U6744 (N_6744,N_5853,N_5261);
or U6745 (N_6745,N_5232,N_5618);
nor U6746 (N_6746,N_5832,N_5289);
nand U6747 (N_6747,N_5793,N_5426);
and U6748 (N_6748,N_5529,N_5379);
nand U6749 (N_6749,N_5121,N_5491);
and U6750 (N_6750,N_5162,N_5479);
nor U6751 (N_6751,N_5480,N_5242);
and U6752 (N_6752,N_5818,N_5113);
nand U6753 (N_6753,N_5945,N_5214);
or U6754 (N_6754,N_5824,N_5542);
nand U6755 (N_6755,N_5509,N_5934);
nand U6756 (N_6756,N_5260,N_5450);
xor U6757 (N_6757,N_5590,N_5922);
and U6758 (N_6758,N_5709,N_5670);
nor U6759 (N_6759,N_5048,N_5712);
or U6760 (N_6760,N_5391,N_5060);
and U6761 (N_6761,N_5284,N_5420);
or U6762 (N_6762,N_5186,N_5016);
nand U6763 (N_6763,N_5130,N_5192);
and U6764 (N_6764,N_5935,N_5099);
nand U6765 (N_6765,N_5551,N_5092);
nand U6766 (N_6766,N_5352,N_5257);
nand U6767 (N_6767,N_5224,N_5145);
xnor U6768 (N_6768,N_5745,N_5273);
and U6769 (N_6769,N_5100,N_5788);
nor U6770 (N_6770,N_5361,N_5171);
nand U6771 (N_6771,N_5041,N_5872);
nor U6772 (N_6772,N_5052,N_5488);
or U6773 (N_6773,N_5916,N_5353);
nor U6774 (N_6774,N_5192,N_5641);
nand U6775 (N_6775,N_5973,N_5514);
nor U6776 (N_6776,N_5297,N_5703);
and U6777 (N_6777,N_5757,N_5961);
nor U6778 (N_6778,N_5347,N_5549);
or U6779 (N_6779,N_5533,N_5443);
or U6780 (N_6780,N_5125,N_5569);
nor U6781 (N_6781,N_5602,N_5868);
and U6782 (N_6782,N_5715,N_5897);
nand U6783 (N_6783,N_5687,N_5508);
nor U6784 (N_6784,N_5891,N_5856);
nor U6785 (N_6785,N_5329,N_5805);
and U6786 (N_6786,N_5598,N_5685);
nand U6787 (N_6787,N_5699,N_5811);
and U6788 (N_6788,N_5546,N_5251);
xnor U6789 (N_6789,N_5230,N_5766);
nor U6790 (N_6790,N_5212,N_5303);
and U6791 (N_6791,N_5853,N_5019);
and U6792 (N_6792,N_5193,N_5966);
or U6793 (N_6793,N_5749,N_5307);
nand U6794 (N_6794,N_5129,N_5158);
or U6795 (N_6795,N_5139,N_5544);
nand U6796 (N_6796,N_5538,N_5072);
nor U6797 (N_6797,N_5443,N_5824);
nand U6798 (N_6798,N_5616,N_5569);
or U6799 (N_6799,N_5614,N_5540);
and U6800 (N_6800,N_5254,N_5718);
and U6801 (N_6801,N_5591,N_5491);
nand U6802 (N_6802,N_5023,N_5537);
or U6803 (N_6803,N_5563,N_5608);
or U6804 (N_6804,N_5630,N_5461);
nand U6805 (N_6805,N_5308,N_5704);
nand U6806 (N_6806,N_5091,N_5800);
nor U6807 (N_6807,N_5772,N_5050);
nand U6808 (N_6808,N_5403,N_5802);
and U6809 (N_6809,N_5067,N_5543);
or U6810 (N_6810,N_5688,N_5501);
xnor U6811 (N_6811,N_5816,N_5083);
nor U6812 (N_6812,N_5303,N_5200);
nand U6813 (N_6813,N_5987,N_5694);
and U6814 (N_6814,N_5879,N_5993);
nand U6815 (N_6815,N_5818,N_5323);
and U6816 (N_6816,N_5710,N_5177);
or U6817 (N_6817,N_5397,N_5450);
nor U6818 (N_6818,N_5826,N_5634);
nor U6819 (N_6819,N_5403,N_5274);
and U6820 (N_6820,N_5354,N_5502);
nor U6821 (N_6821,N_5177,N_5302);
nand U6822 (N_6822,N_5827,N_5357);
or U6823 (N_6823,N_5663,N_5010);
nor U6824 (N_6824,N_5838,N_5707);
or U6825 (N_6825,N_5846,N_5440);
nor U6826 (N_6826,N_5819,N_5066);
or U6827 (N_6827,N_5619,N_5215);
or U6828 (N_6828,N_5276,N_5734);
nor U6829 (N_6829,N_5881,N_5321);
nor U6830 (N_6830,N_5944,N_5396);
or U6831 (N_6831,N_5124,N_5230);
and U6832 (N_6832,N_5635,N_5227);
or U6833 (N_6833,N_5279,N_5912);
or U6834 (N_6834,N_5252,N_5731);
nand U6835 (N_6835,N_5886,N_5085);
nor U6836 (N_6836,N_5636,N_5219);
nor U6837 (N_6837,N_5713,N_5440);
and U6838 (N_6838,N_5422,N_5955);
and U6839 (N_6839,N_5851,N_5892);
nand U6840 (N_6840,N_5886,N_5303);
or U6841 (N_6841,N_5530,N_5496);
and U6842 (N_6842,N_5568,N_5227);
nand U6843 (N_6843,N_5253,N_5537);
and U6844 (N_6844,N_5526,N_5978);
nor U6845 (N_6845,N_5253,N_5613);
nor U6846 (N_6846,N_5574,N_5067);
nor U6847 (N_6847,N_5142,N_5641);
nor U6848 (N_6848,N_5615,N_5949);
or U6849 (N_6849,N_5199,N_5864);
or U6850 (N_6850,N_5737,N_5578);
nand U6851 (N_6851,N_5128,N_5846);
or U6852 (N_6852,N_5494,N_5787);
or U6853 (N_6853,N_5770,N_5019);
nor U6854 (N_6854,N_5170,N_5975);
nand U6855 (N_6855,N_5234,N_5801);
or U6856 (N_6856,N_5529,N_5754);
and U6857 (N_6857,N_5659,N_5471);
nand U6858 (N_6858,N_5586,N_5014);
or U6859 (N_6859,N_5536,N_5432);
or U6860 (N_6860,N_5074,N_5242);
nor U6861 (N_6861,N_5392,N_5920);
and U6862 (N_6862,N_5516,N_5473);
and U6863 (N_6863,N_5554,N_5742);
nand U6864 (N_6864,N_5218,N_5898);
or U6865 (N_6865,N_5923,N_5811);
nor U6866 (N_6866,N_5188,N_5415);
nor U6867 (N_6867,N_5222,N_5674);
nand U6868 (N_6868,N_5882,N_5944);
nor U6869 (N_6869,N_5109,N_5073);
nand U6870 (N_6870,N_5236,N_5615);
and U6871 (N_6871,N_5313,N_5489);
nor U6872 (N_6872,N_5449,N_5002);
or U6873 (N_6873,N_5303,N_5744);
nand U6874 (N_6874,N_5915,N_5996);
or U6875 (N_6875,N_5488,N_5207);
nor U6876 (N_6876,N_5552,N_5330);
or U6877 (N_6877,N_5411,N_5654);
or U6878 (N_6878,N_5493,N_5522);
or U6879 (N_6879,N_5663,N_5918);
nand U6880 (N_6880,N_5023,N_5498);
or U6881 (N_6881,N_5649,N_5987);
or U6882 (N_6882,N_5481,N_5385);
nand U6883 (N_6883,N_5985,N_5196);
and U6884 (N_6884,N_5878,N_5432);
or U6885 (N_6885,N_5058,N_5321);
or U6886 (N_6886,N_5697,N_5737);
or U6887 (N_6887,N_5540,N_5830);
and U6888 (N_6888,N_5217,N_5305);
and U6889 (N_6889,N_5180,N_5447);
and U6890 (N_6890,N_5012,N_5133);
nand U6891 (N_6891,N_5164,N_5237);
or U6892 (N_6892,N_5543,N_5044);
and U6893 (N_6893,N_5920,N_5495);
and U6894 (N_6894,N_5746,N_5953);
or U6895 (N_6895,N_5466,N_5688);
nor U6896 (N_6896,N_5805,N_5471);
and U6897 (N_6897,N_5351,N_5744);
or U6898 (N_6898,N_5936,N_5264);
or U6899 (N_6899,N_5100,N_5230);
and U6900 (N_6900,N_5363,N_5126);
or U6901 (N_6901,N_5538,N_5588);
nor U6902 (N_6902,N_5335,N_5151);
and U6903 (N_6903,N_5629,N_5877);
nor U6904 (N_6904,N_5270,N_5506);
or U6905 (N_6905,N_5102,N_5448);
nand U6906 (N_6906,N_5925,N_5391);
nor U6907 (N_6907,N_5524,N_5848);
or U6908 (N_6908,N_5918,N_5573);
or U6909 (N_6909,N_5095,N_5676);
nand U6910 (N_6910,N_5172,N_5782);
nand U6911 (N_6911,N_5289,N_5637);
nor U6912 (N_6912,N_5995,N_5229);
nor U6913 (N_6913,N_5383,N_5945);
nor U6914 (N_6914,N_5874,N_5659);
xor U6915 (N_6915,N_5182,N_5585);
nor U6916 (N_6916,N_5655,N_5145);
nand U6917 (N_6917,N_5015,N_5600);
and U6918 (N_6918,N_5101,N_5255);
and U6919 (N_6919,N_5065,N_5393);
nand U6920 (N_6920,N_5629,N_5517);
nor U6921 (N_6921,N_5713,N_5986);
nand U6922 (N_6922,N_5347,N_5489);
or U6923 (N_6923,N_5857,N_5384);
nor U6924 (N_6924,N_5454,N_5734);
or U6925 (N_6925,N_5468,N_5209);
and U6926 (N_6926,N_5207,N_5760);
nor U6927 (N_6927,N_5049,N_5152);
and U6928 (N_6928,N_5912,N_5072);
nand U6929 (N_6929,N_5253,N_5776);
or U6930 (N_6930,N_5701,N_5894);
nand U6931 (N_6931,N_5745,N_5960);
nand U6932 (N_6932,N_5450,N_5906);
and U6933 (N_6933,N_5644,N_5715);
nand U6934 (N_6934,N_5746,N_5726);
nor U6935 (N_6935,N_5580,N_5277);
nand U6936 (N_6936,N_5520,N_5531);
nand U6937 (N_6937,N_5786,N_5038);
xor U6938 (N_6938,N_5503,N_5607);
or U6939 (N_6939,N_5177,N_5719);
and U6940 (N_6940,N_5917,N_5421);
and U6941 (N_6941,N_5762,N_5472);
nor U6942 (N_6942,N_5708,N_5423);
or U6943 (N_6943,N_5217,N_5868);
nor U6944 (N_6944,N_5578,N_5817);
and U6945 (N_6945,N_5954,N_5081);
or U6946 (N_6946,N_5770,N_5667);
nand U6947 (N_6947,N_5389,N_5683);
or U6948 (N_6948,N_5366,N_5871);
nor U6949 (N_6949,N_5533,N_5661);
nand U6950 (N_6950,N_5742,N_5864);
or U6951 (N_6951,N_5700,N_5279);
nor U6952 (N_6952,N_5735,N_5289);
and U6953 (N_6953,N_5709,N_5200);
nor U6954 (N_6954,N_5545,N_5827);
nor U6955 (N_6955,N_5053,N_5963);
nand U6956 (N_6956,N_5444,N_5724);
nor U6957 (N_6957,N_5118,N_5130);
or U6958 (N_6958,N_5562,N_5945);
nor U6959 (N_6959,N_5384,N_5494);
nand U6960 (N_6960,N_5977,N_5417);
xnor U6961 (N_6961,N_5430,N_5335);
nor U6962 (N_6962,N_5057,N_5231);
nor U6963 (N_6963,N_5058,N_5057);
or U6964 (N_6964,N_5787,N_5504);
nor U6965 (N_6965,N_5954,N_5252);
and U6966 (N_6966,N_5881,N_5955);
or U6967 (N_6967,N_5021,N_5060);
nor U6968 (N_6968,N_5717,N_5584);
and U6969 (N_6969,N_5715,N_5769);
or U6970 (N_6970,N_5315,N_5446);
or U6971 (N_6971,N_5152,N_5133);
and U6972 (N_6972,N_5076,N_5354);
nand U6973 (N_6973,N_5635,N_5588);
and U6974 (N_6974,N_5338,N_5371);
nor U6975 (N_6975,N_5127,N_5779);
or U6976 (N_6976,N_5393,N_5129);
and U6977 (N_6977,N_5324,N_5705);
nand U6978 (N_6978,N_5848,N_5106);
or U6979 (N_6979,N_5156,N_5962);
and U6980 (N_6980,N_5263,N_5977);
and U6981 (N_6981,N_5570,N_5882);
or U6982 (N_6982,N_5858,N_5231);
nor U6983 (N_6983,N_5172,N_5242);
and U6984 (N_6984,N_5282,N_5178);
and U6985 (N_6985,N_5264,N_5656);
nand U6986 (N_6986,N_5034,N_5832);
nor U6987 (N_6987,N_5215,N_5889);
and U6988 (N_6988,N_5273,N_5212);
or U6989 (N_6989,N_5968,N_5686);
and U6990 (N_6990,N_5418,N_5088);
xor U6991 (N_6991,N_5747,N_5744);
xnor U6992 (N_6992,N_5413,N_5992);
and U6993 (N_6993,N_5242,N_5483);
and U6994 (N_6994,N_5440,N_5067);
nor U6995 (N_6995,N_5714,N_5945);
and U6996 (N_6996,N_5113,N_5926);
or U6997 (N_6997,N_5806,N_5811);
or U6998 (N_6998,N_5847,N_5314);
nor U6999 (N_6999,N_5069,N_5805);
and U7000 (N_7000,N_6525,N_6568);
and U7001 (N_7001,N_6010,N_6433);
nand U7002 (N_7002,N_6660,N_6695);
or U7003 (N_7003,N_6925,N_6295);
and U7004 (N_7004,N_6019,N_6068);
and U7005 (N_7005,N_6641,N_6228);
nor U7006 (N_7006,N_6968,N_6986);
nor U7007 (N_7007,N_6051,N_6537);
nor U7008 (N_7008,N_6678,N_6953);
or U7009 (N_7009,N_6382,N_6574);
nand U7010 (N_7010,N_6099,N_6948);
nor U7011 (N_7011,N_6963,N_6760);
nor U7012 (N_7012,N_6244,N_6455);
or U7013 (N_7013,N_6006,N_6701);
nor U7014 (N_7014,N_6539,N_6045);
and U7015 (N_7015,N_6161,N_6384);
and U7016 (N_7016,N_6825,N_6487);
nor U7017 (N_7017,N_6728,N_6935);
or U7018 (N_7018,N_6704,N_6470);
or U7019 (N_7019,N_6600,N_6037);
nor U7020 (N_7020,N_6330,N_6196);
nand U7021 (N_7021,N_6282,N_6867);
nor U7022 (N_7022,N_6849,N_6916);
nand U7023 (N_7023,N_6338,N_6503);
nand U7024 (N_7024,N_6100,N_6693);
nor U7025 (N_7025,N_6608,N_6709);
nand U7026 (N_7026,N_6359,N_6680);
nand U7027 (N_7027,N_6234,N_6242);
or U7028 (N_7028,N_6522,N_6665);
or U7029 (N_7029,N_6349,N_6092);
and U7030 (N_7030,N_6872,N_6500);
nor U7031 (N_7031,N_6418,N_6869);
and U7032 (N_7032,N_6602,N_6669);
and U7033 (N_7033,N_6812,N_6401);
nand U7034 (N_7034,N_6261,N_6969);
nand U7035 (N_7035,N_6572,N_6447);
and U7036 (N_7036,N_6094,N_6932);
or U7037 (N_7037,N_6906,N_6259);
and U7038 (N_7038,N_6769,N_6508);
and U7039 (N_7039,N_6210,N_6553);
xnor U7040 (N_7040,N_6482,N_6144);
or U7041 (N_7041,N_6276,N_6610);
and U7042 (N_7042,N_6871,N_6675);
or U7043 (N_7043,N_6900,N_6979);
and U7044 (N_7044,N_6150,N_6644);
nor U7045 (N_7045,N_6035,N_6926);
or U7046 (N_7046,N_6718,N_6442);
nand U7047 (N_7047,N_6931,N_6791);
and U7048 (N_7048,N_6342,N_6227);
and U7049 (N_7049,N_6648,N_6097);
or U7050 (N_7050,N_6598,N_6505);
nand U7051 (N_7051,N_6381,N_6657);
xnor U7052 (N_7052,N_6663,N_6185);
and U7053 (N_7053,N_6400,N_6393);
or U7054 (N_7054,N_6914,N_6011);
or U7055 (N_7055,N_6782,N_6107);
nand U7056 (N_7056,N_6681,N_6434);
nor U7057 (N_7057,N_6885,N_6367);
nand U7058 (N_7058,N_6403,N_6766);
nand U7059 (N_7059,N_6621,N_6959);
nand U7060 (N_7060,N_6886,N_6221);
or U7061 (N_7061,N_6938,N_6375);
nand U7062 (N_7062,N_6694,N_6379);
or U7063 (N_7063,N_6217,N_6805);
nor U7064 (N_7064,N_6225,N_6910);
and U7065 (N_7065,N_6806,N_6875);
or U7066 (N_7066,N_6363,N_6889);
nor U7067 (N_7067,N_6873,N_6304);
and U7068 (N_7068,N_6321,N_6030);
nand U7069 (N_7069,N_6267,N_6745);
or U7070 (N_7070,N_6836,N_6499);
or U7071 (N_7071,N_6588,N_6133);
and U7072 (N_7072,N_6322,N_6200);
nand U7073 (N_7073,N_6488,N_6879);
or U7074 (N_7074,N_6802,N_6104);
nand U7075 (N_7075,N_6902,N_6898);
or U7076 (N_7076,N_6016,N_6230);
nand U7077 (N_7077,N_6524,N_6826);
or U7078 (N_7078,N_6843,N_6646);
or U7079 (N_7079,N_6049,N_6586);
and U7080 (N_7080,N_6765,N_6197);
nor U7081 (N_7081,N_6854,N_6479);
or U7082 (N_7082,N_6702,N_6134);
and U7083 (N_7083,N_6776,N_6619);
and U7084 (N_7084,N_6033,N_6967);
nand U7085 (N_7085,N_6192,N_6801);
or U7086 (N_7086,N_6461,N_6733);
and U7087 (N_7087,N_6611,N_6477);
and U7088 (N_7088,N_6135,N_6048);
nand U7089 (N_7089,N_6478,N_6369);
and U7090 (N_7090,N_6091,N_6002);
and U7091 (N_7091,N_6506,N_6893);
and U7092 (N_7092,N_6399,N_6162);
nand U7093 (N_7093,N_6157,N_6392);
or U7094 (N_7094,N_6268,N_6587);
nand U7095 (N_7095,N_6951,N_6909);
nand U7096 (N_7096,N_6457,N_6089);
and U7097 (N_7097,N_6545,N_6884);
and U7098 (N_7098,N_6058,N_6489);
or U7099 (N_7099,N_6652,N_6748);
nor U7100 (N_7100,N_6352,N_6140);
nor U7101 (N_7101,N_6582,N_6204);
and U7102 (N_7102,N_6744,N_6655);
nand U7103 (N_7103,N_6296,N_6087);
or U7104 (N_7104,N_6905,N_6737);
or U7105 (N_7105,N_6570,N_6216);
or U7106 (N_7106,N_6146,N_6281);
nand U7107 (N_7107,N_6565,N_6618);
nand U7108 (N_7108,N_6376,N_6449);
nor U7109 (N_7109,N_6891,N_6160);
or U7110 (N_7110,N_6992,N_6111);
and U7111 (N_7111,N_6387,N_6284);
nand U7112 (N_7112,N_6336,N_6498);
nor U7113 (N_7113,N_6725,N_6650);
and U7114 (N_7114,N_6394,N_6763);
and U7115 (N_7115,N_6086,N_6341);
xor U7116 (N_7116,N_6550,N_6260);
and U7117 (N_7117,N_6638,N_6429);
nor U7118 (N_7118,N_6520,N_6647);
nor U7119 (N_7119,N_6291,N_6184);
nor U7120 (N_7120,N_6922,N_6332);
nor U7121 (N_7121,N_6700,N_6233);
and U7122 (N_7122,N_6036,N_6406);
nand U7123 (N_7123,N_6278,N_6437);
nand U7124 (N_7124,N_6417,N_6989);
nand U7125 (N_7125,N_6159,N_6164);
and U7126 (N_7126,N_6542,N_6633);
or U7127 (N_7127,N_6031,N_6102);
or U7128 (N_7128,N_6947,N_6309);
or U7129 (N_7129,N_6209,N_6121);
or U7130 (N_7130,N_6328,N_6380);
nor U7131 (N_7131,N_6564,N_6552);
nor U7132 (N_7132,N_6991,N_6569);
and U7133 (N_7133,N_6915,N_6356);
xnor U7134 (N_7134,N_6696,N_6592);
or U7135 (N_7135,N_6028,N_6013);
and U7136 (N_7136,N_6466,N_6684);
nand U7137 (N_7137,N_6787,N_6865);
nor U7138 (N_7138,N_6088,N_6327);
nand U7139 (N_7139,N_6710,N_6176);
and U7140 (N_7140,N_6739,N_6138);
or U7141 (N_7141,N_6115,N_6612);
nand U7142 (N_7142,N_6651,N_6667);
nor U7143 (N_7143,N_6292,N_6168);
and U7144 (N_7144,N_6324,N_6180);
nor U7145 (N_7145,N_6976,N_6985);
nand U7146 (N_7146,N_6844,N_6531);
and U7147 (N_7147,N_6590,N_6966);
and U7148 (N_7148,N_6368,N_6679);
or U7149 (N_7149,N_6015,N_6713);
nand U7150 (N_7150,N_6562,N_6474);
nand U7151 (N_7151,N_6307,N_6639);
nor U7152 (N_7152,N_6853,N_6996);
nor U7153 (N_7153,N_6751,N_6946);
or U7154 (N_7154,N_6269,N_6012);
nor U7155 (N_7155,N_6476,N_6485);
nand U7156 (N_7156,N_6211,N_6313);
or U7157 (N_7157,N_6014,N_6720);
nor U7158 (N_7158,N_6212,N_6156);
nand U7159 (N_7159,N_6017,N_6558);
and U7160 (N_7160,N_6344,N_6768);
nand U7161 (N_7161,N_6821,N_6214);
or U7162 (N_7162,N_6544,N_6730);
or U7163 (N_7163,N_6056,N_6927);
or U7164 (N_7164,N_6264,N_6706);
nand U7165 (N_7165,N_6365,N_6753);
nand U7166 (N_7166,N_6990,N_6983);
or U7167 (N_7167,N_6073,N_6833);
or U7168 (N_7168,N_6472,N_6205);
or U7169 (N_7169,N_6874,N_6984);
nand U7170 (N_7170,N_6691,N_6166);
nand U7171 (N_7171,N_6517,N_6756);
nor U7172 (N_7172,N_6391,N_6141);
nor U7173 (N_7173,N_6960,N_6090);
nand U7174 (N_7174,N_6154,N_6395);
nand U7175 (N_7175,N_6734,N_6779);
and U7176 (N_7176,N_6813,N_6436);
nand U7177 (N_7177,N_6731,N_6145);
or U7178 (N_7178,N_6546,N_6270);
and U7179 (N_7179,N_6320,N_6512);
nand U7180 (N_7180,N_6523,N_6593);
nand U7181 (N_7181,N_6762,N_6740);
nor U7182 (N_7182,N_6232,N_6754);
nand U7183 (N_7183,N_6152,N_6428);
or U7184 (N_7184,N_6290,N_6082);
or U7185 (N_7185,N_6604,N_6054);
and U7186 (N_7186,N_6974,N_6005);
nor U7187 (N_7187,N_6065,N_6982);
nand U7188 (N_7188,N_6323,N_6777);
or U7189 (N_7189,N_6183,N_6122);
nand U7190 (N_7190,N_6548,N_6796);
nand U7191 (N_7191,N_6131,N_6841);
nor U7192 (N_7192,N_6599,N_6607);
and U7193 (N_7193,N_6852,N_6919);
and U7194 (N_7194,N_6024,N_6827);
nor U7195 (N_7195,N_6075,N_6415);
and U7196 (N_7196,N_6147,N_6697);
nand U7197 (N_7197,N_6772,N_6585);
or U7198 (N_7198,N_6070,N_6993);
and U7199 (N_7199,N_6003,N_6924);
nor U7200 (N_7200,N_6312,N_6819);
and U7201 (N_7201,N_6943,N_6396);
nand U7202 (N_7202,N_6920,N_6007);
nor U7203 (N_7203,N_6761,N_6830);
or U7204 (N_7204,N_6882,N_6239);
xnor U7205 (N_7205,N_6723,N_6972);
xnor U7206 (N_7206,N_6591,N_6021);
nand U7207 (N_7207,N_6858,N_6468);
and U7208 (N_7208,N_6664,N_6334);
nor U7209 (N_7209,N_6559,N_6117);
nand U7210 (N_7210,N_6294,N_6462);
nand U7211 (N_7211,N_6452,N_6136);
nor U7212 (N_7212,N_6224,N_6677);
nor U7213 (N_7213,N_6179,N_6653);
and U7214 (N_7214,N_6670,N_6249);
nand U7215 (N_7215,N_6529,N_6305);
nand U7216 (N_7216,N_6783,N_6957);
or U7217 (N_7217,N_6189,N_6308);
or U7218 (N_7218,N_6518,N_6596);
nand U7219 (N_7219,N_6818,N_6556);
and U7220 (N_7220,N_6732,N_6850);
nand U7221 (N_7221,N_6894,N_6041);
and U7222 (N_7222,N_6186,N_6536);
nor U7223 (N_7223,N_6315,N_6325);
or U7224 (N_7224,N_6888,N_6866);
nand U7225 (N_7225,N_6692,N_6130);
nand U7226 (N_7226,N_6250,N_6551);
or U7227 (N_7227,N_6347,N_6288);
or U7228 (N_7228,N_6842,N_6208);
and U7229 (N_7229,N_6977,N_6907);
nand U7230 (N_7230,N_6809,N_6816);
nand U7231 (N_7231,N_6540,N_6000);
nand U7232 (N_7232,N_6273,N_6170);
or U7233 (N_7233,N_6335,N_6213);
nand U7234 (N_7234,N_6659,N_6950);
and U7235 (N_7235,N_6061,N_6034);
nor U7236 (N_7236,N_6630,N_6254);
and U7237 (N_7237,N_6439,N_6839);
nor U7238 (N_7238,N_6686,N_6509);
or U7239 (N_7239,N_6738,N_6481);
or U7240 (N_7240,N_6158,N_6543);
nand U7241 (N_7241,N_6222,N_6794);
nor U7242 (N_7242,N_6774,N_6823);
nor U7243 (N_7243,N_6052,N_6246);
nor U7244 (N_7244,N_6820,N_6174);
xor U7245 (N_7245,N_6257,N_6845);
nor U7246 (N_7246,N_6661,N_6649);
or U7247 (N_7247,N_6420,N_6412);
nand U7248 (N_7248,N_6719,N_6642);
and U7249 (N_7249,N_6377,N_6448);
nand U7250 (N_7250,N_6705,N_6248);
nor U7251 (N_7251,N_6609,N_6383);
nand U7252 (N_7252,N_6666,N_6980);
nand U7253 (N_7253,N_6673,N_6658);
nor U7254 (N_7254,N_6863,N_6502);
nand U7255 (N_7255,N_6237,N_6577);
or U7256 (N_7256,N_6057,N_6617);
nand U7257 (N_7257,N_6044,N_6188);
nor U7258 (N_7258,N_6530,N_6634);
or U7259 (N_7259,N_6716,N_6202);
or U7260 (N_7260,N_6746,N_6859);
and U7261 (N_7261,N_6930,N_6450);
or U7262 (N_7262,N_6654,N_6469);
or U7263 (N_7263,N_6625,N_6419);
nor U7264 (N_7264,N_6635,N_6864);
or U7265 (N_7265,N_6566,N_6573);
or U7266 (N_7266,N_6965,N_6085);
nand U7267 (N_7267,N_6274,N_6535);
and U7268 (N_7268,N_6119,N_6781);
or U7269 (N_7269,N_6042,N_6892);
and U7270 (N_7270,N_6435,N_6899);
or U7271 (N_7271,N_6632,N_6263);
and U7272 (N_7272,N_6703,N_6473);
and U7273 (N_7273,N_6171,N_6912);
nand U7274 (N_7274,N_6143,N_6835);
nand U7275 (N_7275,N_6672,N_6631);
nor U7276 (N_7276,N_6364,N_6329);
or U7277 (N_7277,N_6516,N_6219);
nand U7278 (N_7278,N_6124,N_6637);
nor U7279 (N_7279,N_6949,N_6220);
and U7280 (N_7280,N_6408,N_6062);
and U7281 (N_7281,N_6771,N_6757);
and U7282 (N_7282,N_6173,N_6767);
and U7283 (N_7283,N_6443,N_6741);
and U7284 (N_7284,N_6319,N_6626);
or U7285 (N_7285,N_6717,N_6624);
or U7286 (N_7286,N_6354,N_6575);
and U7287 (N_7287,N_6108,N_6605);
or U7288 (N_7288,N_6265,N_6764);
nand U7289 (N_7289,N_6861,N_6331);
and U7290 (N_7290,N_6008,N_6759);
and U7291 (N_7291,N_6998,N_6151);
or U7292 (N_7292,N_6149,N_6814);
nand U7293 (N_7293,N_6606,N_6358);
nand U7294 (N_7294,N_6676,N_6390);
nor U7295 (N_7295,N_6125,N_6528);
or U7296 (N_7296,N_6576,N_6807);
nand U7297 (N_7297,N_6510,N_6193);
or U7298 (N_7298,N_6629,N_6688);
nor U7299 (N_7299,N_6431,N_6169);
or U7300 (N_7300,N_6563,N_6962);
nand U7301 (N_7301,N_6275,N_6067);
and U7302 (N_7302,N_6009,N_6775);
or U7303 (N_7303,N_6685,N_6580);
nor U7304 (N_7304,N_6451,N_6640);
and U7305 (N_7305,N_6317,N_6083);
or U7306 (N_7306,N_6271,N_6355);
nand U7307 (N_7307,N_6229,N_6050);
nor U7308 (N_7308,N_6623,N_6620);
or U7309 (N_7309,N_6043,N_6627);
and U7310 (N_7310,N_6194,N_6215);
and U7311 (N_7311,N_6421,N_6360);
and U7312 (N_7312,N_6897,N_6303);
nand U7313 (N_7313,N_6832,N_6126);
and U7314 (N_7314,N_6300,N_6887);
or U7315 (N_7315,N_6615,N_6554);
and U7316 (N_7316,N_6750,N_6671);
nand U7317 (N_7317,N_6792,N_6973);
nand U7318 (N_7318,N_6484,N_6252);
nand U7319 (N_7319,N_6311,N_6103);
or U7320 (N_7320,N_6595,N_6128);
nor U7321 (N_7321,N_6815,N_6432);
or U7322 (N_7322,N_6862,N_6857);
nor U7323 (N_7323,N_6256,N_6579);
or U7324 (N_7324,N_6662,N_6714);
nor U7325 (N_7325,N_6971,N_6939);
xor U7326 (N_7326,N_6808,N_6253);
nand U7327 (N_7327,N_6371,N_6077);
and U7328 (N_7328,N_6454,N_6942);
nand U7329 (N_7329,N_6430,N_6870);
and U7330 (N_7330,N_6306,N_6023);
or U7331 (N_7331,N_6527,N_6109);
nand U7332 (N_7332,N_6172,N_6243);
or U7333 (N_7333,N_6824,N_6712);
or U7334 (N_7334,N_6690,N_6464);
and U7335 (N_7335,N_6567,N_6093);
nor U7336 (N_7336,N_6722,N_6118);
nor U7337 (N_7337,N_6409,N_6046);
nand U7338 (N_7338,N_6682,N_6726);
or U7339 (N_7339,N_6601,N_6445);
nand U7340 (N_7340,N_6923,N_6940);
xor U7341 (N_7341,N_6496,N_6645);
nand U7342 (N_7342,N_6287,N_6533);
or U7343 (N_7343,N_6803,N_6201);
nor U7344 (N_7344,N_6238,N_6933);
or U7345 (N_7345,N_6860,N_6001);
nand U7346 (N_7346,N_6397,N_6416);
and U7347 (N_7347,N_6438,N_6203);
or U7348 (N_7348,N_6069,N_6055);
nor U7349 (N_7349,N_6786,N_6778);
or U7350 (N_7350,N_6426,N_6074);
or U7351 (N_7351,N_6137,N_6280);
or U7352 (N_7352,N_6095,N_6106);
nand U7353 (N_7353,N_6471,N_6921);
or U7354 (N_7354,N_6708,N_6155);
or U7355 (N_7355,N_6080,N_6538);
nor U7356 (N_7356,N_6483,N_6956);
and U7357 (N_7357,N_6402,N_6828);
nor U7358 (N_7358,N_6285,N_6797);
xor U7359 (N_7359,N_6277,N_6316);
and U7360 (N_7360,N_6486,N_6878);
nor U7361 (N_7361,N_6195,N_6495);
nor U7362 (N_7362,N_6715,N_6903);
nand U7363 (N_7363,N_6883,N_6851);
nand U7364 (N_7364,N_6079,N_6848);
nor U7365 (N_7365,N_6343,N_6027);
and U7366 (N_7366,N_6683,N_6594);
nand U7367 (N_7367,N_6339,N_6289);
or U7368 (N_7368,N_6752,N_6226);
or U7369 (N_7369,N_6597,N_6876);
nor U7370 (N_7370,N_6978,N_6521);
or U7371 (N_7371,N_6385,N_6504);
nor U7372 (N_7372,N_6139,N_6440);
and U7373 (N_7373,N_6346,N_6223);
and U7374 (N_7374,N_6492,N_6191);
nor U7375 (N_7375,N_6829,N_6999);
and U7376 (N_7376,N_6788,N_6881);
nor U7377 (N_7377,N_6114,N_6785);
nor U7378 (N_7378,N_6297,N_6370);
nand U7379 (N_7379,N_6362,N_6326);
nand U7380 (N_7380,N_6299,N_6795);
nand U7381 (N_7381,N_6283,N_6129);
nor U7382 (N_7382,N_6236,N_6386);
and U7383 (N_7383,N_6707,N_6231);
nor U7384 (N_7384,N_6987,N_6961);
and U7385 (N_7385,N_6410,N_6467);
and U7386 (N_7386,N_6736,N_6822);
or U7387 (N_7387,N_6072,N_6560);
nand U7388 (N_7388,N_6148,N_6494);
or U7389 (N_7389,N_6798,N_6020);
nor U7390 (N_7390,N_6847,N_6446);
nor U7391 (N_7391,N_6441,N_6954);
and U7392 (N_7392,N_6272,N_6724);
and U7393 (N_7393,N_6241,N_6318);
or U7394 (N_7394,N_6081,N_6247);
nand U7395 (N_7395,N_6643,N_6742);
nand U7396 (N_7396,N_6064,N_6404);
and U7397 (N_7397,N_6532,N_6994);
nand U7398 (N_7398,N_6444,N_6571);
nor U7399 (N_7399,N_6561,N_6749);
and U7400 (N_7400,N_6491,N_6165);
nor U7401 (N_7401,N_6868,N_6790);
nand U7402 (N_7402,N_6747,N_6423);
nor U7403 (N_7403,N_6817,N_6413);
nor U7404 (N_7404,N_6908,N_6970);
and U7405 (N_7405,N_6955,N_6727);
nor U7406 (N_7406,N_6856,N_6799);
and U7407 (N_7407,N_6837,N_6918);
and U7408 (N_7408,N_6698,N_6711);
and U7409 (N_7409,N_6589,N_6032);
xor U7410 (N_7410,N_6901,N_6458);
and U7411 (N_7411,N_6941,N_6934);
and U7412 (N_7412,N_6078,N_6997);
nor U7413 (N_7413,N_6917,N_6025);
or U7414 (N_7414,N_6350,N_6463);
nor U7415 (N_7415,N_6071,N_6846);
nand U7416 (N_7416,N_6348,N_6958);
and U7417 (N_7417,N_6286,N_6513);
and U7418 (N_7418,N_6279,N_6040);
nor U7419 (N_7419,N_6301,N_6182);
nand U7420 (N_7420,N_6519,N_6337);
nor U7421 (N_7421,N_6101,N_6110);
nand U7422 (N_7422,N_6699,N_6378);
nand U7423 (N_7423,N_6583,N_6789);
and U7424 (N_7424,N_6944,N_6459);
nand U7425 (N_7425,N_6310,N_6340);
nor U7426 (N_7426,N_6541,N_6407);
nor U7427 (N_7427,N_6557,N_6112);
or U7428 (N_7428,N_6784,N_6361);
nor U7429 (N_7429,N_6314,N_6258);
or U7430 (N_7430,N_6113,N_6333);
and U7431 (N_7431,N_6026,N_6167);
and U7432 (N_7432,N_6004,N_6255);
and U7433 (N_7433,N_6142,N_6936);
and U7434 (N_7434,N_6465,N_6127);
nand U7435 (N_7435,N_6811,N_6584);
nand U7436 (N_7436,N_6995,N_6218);
and U7437 (N_7437,N_6187,N_6614);
nor U7438 (N_7438,N_6913,N_6411);
nor U7439 (N_7439,N_6029,N_6181);
and U7440 (N_7440,N_6177,N_6603);
nor U7441 (N_7441,N_6235,N_6293);
or U7442 (N_7442,N_6534,N_6022);
or U7443 (N_7443,N_6514,N_6059);
nand U7444 (N_7444,N_6163,N_6735);
or U7445 (N_7445,N_6628,N_6302);
and U7446 (N_7446,N_6613,N_6427);
and U7447 (N_7447,N_6501,N_6493);
nand U7448 (N_7448,N_6855,N_6578);
and U7449 (N_7449,N_6929,N_6687);
nor U7450 (N_7450,N_6729,N_6928);
nor U7451 (N_7451,N_6890,N_6199);
nor U7452 (N_7452,N_6780,N_6262);
nor U7453 (N_7453,N_6840,N_6758);
and U7454 (N_7454,N_6988,N_6123);
and U7455 (N_7455,N_6689,N_6904);
or U7456 (N_7456,N_6098,N_6425);
nand U7457 (N_7457,N_6810,N_6060);
nor U7458 (N_7458,N_6911,N_6206);
and U7459 (N_7459,N_6132,N_6945);
nand U7460 (N_7460,N_6793,N_6674);
or U7461 (N_7461,N_6207,N_6018);
nand U7462 (N_7462,N_6834,N_6076);
or U7463 (N_7463,N_6668,N_6804);
nor U7464 (N_7464,N_6066,N_6116);
nand U7465 (N_7465,N_6047,N_6581);
and U7466 (N_7466,N_6743,N_6721);
nand U7467 (N_7467,N_6063,N_6480);
or U7468 (N_7468,N_6831,N_6053);
nand U7469 (N_7469,N_6547,N_6374);
or U7470 (N_7470,N_6039,N_6120);
or U7471 (N_7471,N_6975,N_6896);
nor U7472 (N_7472,N_6389,N_6251);
or U7473 (N_7473,N_6880,N_6245);
nor U7474 (N_7474,N_6198,N_6981);
and U7475 (N_7475,N_6388,N_6298);
xnor U7476 (N_7476,N_6175,N_6096);
and U7477 (N_7477,N_6460,N_6515);
or U7478 (N_7478,N_6345,N_6105);
nor U7479 (N_7479,N_6084,N_6456);
or U7480 (N_7480,N_6838,N_6497);
nand U7481 (N_7481,N_6190,N_6895);
nor U7482 (N_7482,N_6616,N_6398);
or U7483 (N_7483,N_6351,N_6656);
nor U7484 (N_7484,N_6357,N_6964);
nor U7485 (N_7485,N_6555,N_6372);
nand U7486 (N_7486,N_6240,N_6636);
or U7487 (N_7487,N_6266,N_6937);
nand U7488 (N_7488,N_6414,N_6622);
and U7489 (N_7489,N_6424,N_6405);
nor U7490 (N_7490,N_6153,N_6507);
or U7491 (N_7491,N_6038,N_6422);
and U7492 (N_7492,N_6952,N_6366);
or U7493 (N_7493,N_6773,N_6490);
and U7494 (N_7494,N_6755,N_6453);
and U7495 (N_7495,N_6800,N_6178);
or U7496 (N_7496,N_6353,N_6877);
nor U7497 (N_7497,N_6475,N_6373);
nor U7498 (N_7498,N_6549,N_6770);
or U7499 (N_7499,N_6511,N_6526);
nand U7500 (N_7500,N_6890,N_6196);
or U7501 (N_7501,N_6916,N_6346);
nand U7502 (N_7502,N_6708,N_6892);
or U7503 (N_7503,N_6415,N_6926);
and U7504 (N_7504,N_6751,N_6800);
nor U7505 (N_7505,N_6010,N_6230);
nor U7506 (N_7506,N_6065,N_6706);
and U7507 (N_7507,N_6613,N_6486);
nand U7508 (N_7508,N_6578,N_6045);
nand U7509 (N_7509,N_6771,N_6792);
and U7510 (N_7510,N_6726,N_6101);
nand U7511 (N_7511,N_6514,N_6100);
or U7512 (N_7512,N_6172,N_6517);
and U7513 (N_7513,N_6355,N_6433);
and U7514 (N_7514,N_6407,N_6216);
or U7515 (N_7515,N_6596,N_6908);
or U7516 (N_7516,N_6481,N_6420);
nand U7517 (N_7517,N_6034,N_6560);
or U7518 (N_7518,N_6571,N_6386);
or U7519 (N_7519,N_6901,N_6386);
nor U7520 (N_7520,N_6549,N_6324);
nor U7521 (N_7521,N_6209,N_6923);
and U7522 (N_7522,N_6620,N_6414);
and U7523 (N_7523,N_6442,N_6938);
or U7524 (N_7524,N_6175,N_6662);
xnor U7525 (N_7525,N_6075,N_6676);
xor U7526 (N_7526,N_6243,N_6360);
and U7527 (N_7527,N_6461,N_6164);
nand U7528 (N_7528,N_6848,N_6043);
or U7529 (N_7529,N_6570,N_6281);
or U7530 (N_7530,N_6052,N_6399);
nor U7531 (N_7531,N_6328,N_6071);
and U7532 (N_7532,N_6063,N_6363);
nor U7533 (N_7533,N_6184,N_6222);
nand U7534 (N_7534,N_6254,N_6055);
xnor U7535 (N_7535,N_6367,N_6547);
or U7536 (N_7536,N_6385,N_6186);
nor U7537 (N_7537,N_6668,N_6057);
nand U7538 (N_7538,N_6734,N_6882);
or U7539 (N_7539,N_6080,N_6240);
or U7540 (N_7540,N_6738,N_6562);
or U7541 (N_7541,N_6562,N_6553);
or U7542 (N_7542,N_6578,N_6707);
and U7543 (N_7543,N_6859,N_6782);
or U7544 (N_7544,N_6125,N_6919);
nand U7545 (N_7545,N_6612,N_6026);
and U7546 (N_7546,N_6966,N_6818);
and U7547 (N_7547,N_6334,N_6238);
and U7548 (N_7548,N_6568,N_6498);
nor U7549 (N_7549,N_6725,N_6105);
or U7550 (N_7550,N_6258,N_6149);
and U7551 (N_7551,N_6218,N_6700);
nor U7552 (N_7552,N_6747,N_6296);
nor U7553 (N_7553,N_6134,N_6107);
or U7554 (N_7554,N_6338,N_6326);
nand U7555 (N_7555,N_6269,N_6992);
nand U7556 (N_7556,N_6847,N_6844);
nor U7557 (N_7557,N_6322,N_6416);
or U7558 (N_7558,N_6136,N_6486);
or U7559 (N_7559,N_6912,N_6523);
nor U7560 (N_7560,N_6599,N_6155);
or U7561 (N_7561,N_6964,N_6721);
or U7562 (N_7562,N_6115,N_6753);
nand U7563 (N_7563,N_6461,N_6090);
nor U7564 (N_7564,N_6943,N_6916);
nand U7565 (N_7565,N_6374,N_6230);
or U7566 (N_7566,N_6382,N_6119);
and U7567 (N_7567,N_6458,N_6544);
nor U7568 (N_7568,N_6262,N_6263);
nor U7569 (N_7569,N_6581,N_6220);
nor U7570 (N_7570,N_6579,N_6490);
nand U7571 (N_7571,N_6703,N_6426);
nand U7572 (N_7572,N_6204,N_6024);
or U7573 (N_7573,N_6049,N_6328);
and U7574 (N_7574,N_6183,N_6536);
xor U7575 (N_7575,N_6191,N_6530);
nand U7576 (N_7576,N_6619,N_6671);
nor U7577 (N_7577,N_6568,N_6435);
nand U7578 (N_7578,N_6729,N_6174);
nand U7579 (N_7579,N_6733,N_6463);
and U7580 (N_7580,N_6199,N_6577);
or U7581 (N_7581,N_6446,N_6113);
nor U7582 (N_7582,N_6896,N_6564);
nand U7583 (N_7583,N_6840,N_6810);
nand U7584 (N_7584,N_6969,N_6855);
nor U7585 (N_7585,N_6521,N_6111);
and U7586 (N_7586,N_6732,N_6907);
or U7587 (N_7587,N_6699,N_6448);
and U7588 (N_7588,N_6044,N_6768);
and U7589 (N_7589,N_6167,N_6793);
and U7590 (N_7590,N_6691,N_6082);
or U7591 (N_7591,N_6305,N_6892);
and U7592 (N_7592,N_6635,N_6116);
or U7593 (N_7593,N_6036,N_6658);
nor U7594 (N_7594,N_6313,N_6591);
nor U7595 (N_7595,N_6881,N_6801);
nor U7596 (N_7596,N_6884,N_6095);
or U7597 (N_7597,N_6377,N_6093);
nor U7598 (N_7598,N_6159,N_6336);
or U7599 (N_7599,N_6245,N_6154);
nor U7600 (N_7600,N_6013,N_6365);
nor U7601 (N_7601,N_6333,N_6649);
and U7602 (N_7602,N_6660,N_6676);
nand U7603 (N_7603,N_6246,N_6522);
nand U7604 (N_7604,N_6848,N_6711);
nor U7605 (N_7605,N_6051,N_6743);
or U7606 (N_7606,N_6015,N_6434);
or U7607 (N_7607,N_6095,N_6792);
and U7608 (N_7608,N_6558,N_6418);
nand U7609 (N_7609,N_6942,N_6664);
and U7610 (N_7610,N_6114,N_6106);
nor U7611 (N_7611,N_6454,N_6583);
nor U7612 (N_7612,N_6315,N_6408);
nor U7613 (N_7613,N_6625,N_6889);
nand U7614 (N_7614,N_6187,N_6522);
nand U7615 (N_7615,N_6087,N_6689);
and U7616 (N_7616,N_6790,N_6681);
and U7617 (N_7617,N_6127,N_6501);
and U7618 (N_7618,N_6857,N_6668);
nor U7619 (N_7619,N_6624,N_6365);
and U7620 (N_7620,N_6446,N_6343);
nor U7621 (N_7621,N_6827,N_6465);
nand U7622 (N_7622,N_6852,N_6204);
nand U7623 (N_7623,N_6668,N_6569);
and U7624 (N_7624,N_6827,N_6336);
and U7625 (N_7625,N_6459,N_6376);
nor U7626 (N_7626,N_6991,N_6318);
and U7627 (N_7627,N_6300,N_6637);
nand U7628 (N_7628,N_6093,N_6354);
nand U7629 (N_7629,N_6096,N_6057);
or U7630 (N_7630,N_6656,N_6677);
or U7631 (N_7631,N_6569,N_6391);
nor U7632 (N_7632,N_6188,N_6070);
or U7633 (N_7633,N_6818,N_6432);
nor U7634 (N_7634,N_6935,N_6154);
nor U7635 (N_7635,N_6381,N_6804);
or U7636 (N_7636,N_6645,N_6063);
or U7637 (N_7637,N_6438,N_6875);
and U7638 (N_7638,N_6559,N_6829);
xor U7639 (N_7639,N_6321,N_6527);
nor U7640 (N_7640,N_6413,N_6810);
nor U7641 (N_7641,N_6118,N_6971);
and U7642 (N_7642,N_6067,N_6812);
and U7643 (N_7643,N_6161,N_6335);
nand U7644 (N_7644,N_6843,N_6280);
and U7645 (N_7645,N_6385,N_6573);
or U7646 (N_7646,N_6095,N_6829);
and U7647 (N_7647,N_6054,N_6773);
nor U7648 (N_7648,N_6259,N_6317);
and U7649 (N_7649,N_6087,N_6114);
and U7650 (N_7650,N_6575,N_6155);
or U7651 (N_7651,N_6771,N_6015);
or U7652 (N_7652,N_6171,N_6631);
nor U7653 (N_7653,N_6134,N_6381);
or U7654 (N_7654,N_6396,N_6558);
nor U7655 (N_7655,N_6265,N_6641);
and U7656 (N_7656,N_6970,N_6318);
nor U7657 (N_7657,N_6006,N_6178);
or U7658 (N_7658,N_6203,N_6979);
and U7659 (N_7659,N_6804,N_6742);
and U7660 (N_7660,N_6465,N_6651);
nor U7661 (N_7661,N_6583,N_6098);
nor U7662 (N_7662,N_6363,N_6521);
nand U7663 (N_7663,N_6646,N_6290);
and U7664 (N_7664,N_6016,N_6883);
nor U7665 (N_7665,N_6616,N_6599);
or U7666 (N_7666,N_6114,N_6094);
or U7667 (N_7667,N_6285,N_6978);
nand U7668 (N_7668,N_6671,N_6085);
nor U7669 (N_7669,N_6949,N_6710);
or U7670 (N_7670,N_6810,N_6886);
nor U7671 (N_7671,N_6371,N_6994);
and U7672 (N_7672,N_6734,N_6314);
nand U7673 (N_7673,N_6373,N_6119);
nand U7674 (N_7674,N_6275,N_6286);
nand U7675 (N_7675,N_6181,N_6921);
or U7676 (N_7676,N_6734,N_6460);
nand U7677 (N_7677,N_6892,N_6386);
and U7678 (N_7678,N_6837,N_6242);
and U7679 (N_7679,N_6428,N_6949);
nor U7680 (N_7680,N_6950,N_6159);
or U7681 (N_7681,N_6956,N_6189);
nand U7682 (N_7682,N_6276,N_6200);
nand U7683 (N_7683,N_6560,N_6896);
or U7684 (N_7684,N_6845,N_6031);
and U7685 (N_7685,N_6860,N_6811);
and U7686 (N_7686,N_6164,N_6291);
or U7687 (N_7687,N_6759,N_6221);
nand U7688 (N_7688,N_6319,N_6632);
nor U7689 (N_7689,N_6484,N_6940);
and U7690 (N_7690,N_6603,N_6412);
or U7691 (N_7691,N_6927,N_6550);
or U7692 (N_7692,N_6596,N_6205);
or U7693 (N_7693,N_6410,N_6514);
xor U7694 (N_7694,N_6385,N_6285);
or U7695 (N_7695,N_6245,N_6012);
nor U7696 (N_7696,N_6947,N_6592);
and U7697 (N_7697,N_6926,N_6856);
or U7698 (N_7698,N_6956,N_6800);
xor U7699 (N_7699,N_6467,N_6976);
nand U7700 (N_7700,N_6243,N_6079);
nand U7701 (N_7701,N_6002,N_6256);
or U7702 (N_7702,N_6254,N_6887);
nor U7703 (N_7703,N_6545,N_6607);
nand U7704 (N_7704,N_6418,N_6766);
or U7705 (N_7705,N_6446,N_6541);
nand U7706 (N_7706,N_6345,N_6223);
nand U7707 (N_7707,N_6397,N_6265);
and U7708 (N_7708,N_6311,N_6452);
xnor U7709 (N_7709,N_6133,N_6139);
or U7710 (N_7710,N_6768,N_6636);
nand U7711 (N_7711,N_6294,N_6183);
or U7712 (N_7712,N_6209,N_6126);
nor U7713 (N_7713,N_6610,N_6489);
nor U7714 (N_7714,N_6835,N_6710);
nor U7715 (N_7715,N_6313,N_6859);
nor U7716 (N_7716,N_6137,N_6953);
and U7717 (N_7717,N_6268,N_6738);
or U7718 (N_7718,N_6889,N_6647);
nor U7719 (N_7719,N_6704,N_6821);
or U7720 (N_7720,N_6130,N_6422);
xor U7721 (N_7721,N_6801,N_6808);
or U7722 (N_7722,N_6998,N_6574);
nor U7723 (N_7723,N_6269,N_6460);
or U7724 (N_7724,N_6691,N_6863);
and U7725 (N_7725,N_6635,N_6744);
nor U7726 (N_7726,N_6980,N_6683);
or U7727 (N_7727,N_6211,N_6936);
and U7728 (N_7728,N_6851,N_6098);
nand U7729 (N_7729,N_6835,N_6724);
xnor U7730 (N_7730,N_6260,N_6186);
and U7731 (N_7731,N_6771,N_6006);
or U7732 (N_7732,N_6075,N_6877);
nor U7733 (N_7733,N_6842,N_6978);
nand U7734 (N_7734,N_6991,N_6591);
and U7735 (N_7735,N_6105,N_6027);
or U7736 (N_7736,N_6808,N_6014);
and U7737 (N_7737,N_6895,N_6777);
nand U7738 (N_7738,N_6313,N_6626);
or U7739 (N_7739,N_6831,N_6181);
nand U7740 (N_7740,N_6120,N_6077);
or U7741 (N_7741,N_6318,N_6055);
xor U7742 (N_7742,N_6817,N_6474);
nand U7743 (N_7743,N_6519,N_6159);
nand U7744 (N_7744,N_6669,N_6006);
and U7745 (N_7745,N_6085,N_6971);
and U7746 (N_7746,N_6047,N_6956);
or U7747 (N_7747,N_6498,N_6591);
nand U7748 (N_7748,N_6667,N_6692);
nand U7749 (N_7749,N_6810,N_6235);
or U7750 (N_7750,N_6315,N_6267);
nand U7751 (N_7751,N_6286,N_6460);
and U7752 (N_7752,N_6808,N_6335);
and U7753 (N_7753,N_6289,N_6830);
nor U7754 (N_7754,N_6395,N_6619);
or U7755 (N_7755,N_6433,N_6603);
and U7756 (N_7756,N_6857,N_6548);
nor U7757 (N_7757,N_6034,N_6620);
nor U7758 (N_7758,N_6525,N_6546);
nor U7759 (N_7759,N_6300,N_6022);
nand U7760 (N_7760,N_6036,N_6594);
nor U7761 (N_7761,N_6782,N_6096);
or U7762 (N_7762,N_6630,N_6266);
or U7763 (N_7763,N_6479,N_6602);
nor U7764 (N_7764,N_6214,N_6258);
and U7765 (N_7765,N_6030,N_6331);
or U7766 (N_7766,N_6197,N_6037);
nand U7767 (N_7767,N_6799,N_6301);
or U7768 (N_7768,N_6102,N_6403);
nor U7769 (N_7769,N_6819,N_6489);
xnor U7770 (N_7770,N_6748,N_6448);
nand U7771 (N_7771,N_6947,N_6967);
or U7772 (N_7772,N_6798,N_6482);
and U7773 (N_7773,N_6488,N_6261);
and U7774 (N_7774,N_6915,N_6512);
or U7775 (N_7775,N_6400,N_6484);
and U7776 (N_7776,N_6477,N_6665);
or U7777 (N_7777,N_6432,N_6373);
nor U7778 (N_7778,N_6823,N_6849);
nand U7779 (N_7779,N_6210,N_6319);
and U7780 (N_7780,N_6730,N_6124);
nand U7781 (N_7781,N_6841,N_6056);
nor U7782 (N_7782,N_6831,N_6433);
nand U7783 (N_7783,N_6691,N_6858);
and U7784 (N_7784,N_6583,N_6353);
nand U7785 (N_7785,N_6262,N_6337);
nand U7786 (N_7786,N_6323,N_6628);
nand U7787 (N_7787,N_6096,N_6768);
nor U7788 (N_7788,N_6515,N_6278);
nor U7789 (N_7789,N_6721,N_6228);
or U7790 (N_7790,N_6196,N_6245);
nor U7791 (N_7791,N_6252,N_6090);
nor U7792 (N_7792,N_6584,N_6902);
and U7793 (N_7793,N_6401,N_6640);
or U7794 (N_7794,N_6968,N_6020);
and U7795 (N_7795,N_6264,N_6907);
nand U7796 (N_7796,N_6077,N_6197);
and U7797 (N_7797,N_6933,N_6250);
nand U7798 (N_7798,N_6550,N_6123);
and U7799 (N_7799,N_6750,N_6981);
and U7800 (N_7800,N_6914,N_6466);
nor U7801 (N_7801,N_6350,N_6103);
nor U7802 (N_7802,N_6010,N_6245);
nor U7803 (N_7803,N_6240,N_6126);
or U7804 (N_7804,N_6232,N_6984);
nor U7805 (N_7805,N_6289,N_6058);
or U7806 (N_7806,N_6585,N_6105);
nor U7807 (N_7807,N_6005,N_6133);
or U7808 (N_7808,N_6522,N_6358);
nand U7809 (N_7809,N_6297,N_6870);
nand U7810 (N_7810,N_6319,N_6334);
nor U7811 (N_7811,N_6122,N_6937);
nor U7812 (N_7812,N_6761,N_6516);
and U7813 (N_7813,N_6657,N_6240);
nand U7814 (N_7814,N_6266,N_6599);
nor U7815 (N_7815,N_6206,N_6140);
or U7816 (N_7816,N_6205,N_6755);
and U7817 (N_7817,N_6429,N_6992);
nand U7818 (N_7818,N_6421,N_6661);
and U7819 (N_7819,N_6163,N_6886);
and U7820 (N_7820,N_6093,N_6110);
and U7821 (N_7821,N_6214,N_6361);
nand U7822 (N_7822,N_6717,N_6258);
or U7823 (N_7823,N_6342,N_6836);
nand U7824 (N_7824,N_6787,N_6956);
nand U7825 (N_7825,N_6045,N_6280);
nor U7826 (N_7826,N_6782,N_6245);
or U7827 (N_7827,N_6703,N_6954);
nand U7828 (N_7828,N_6583,N_6075);
and U7829 (N_7829,N_6883,N_6630);
nor U7830 (N_7830,N_6230,N_6235);
and U7831 (N_7831,N_6972,N_6006);
or U7832 (N_7832,N_6274,N_6329);
nor U7833 (N_7833,N_6794,N_6312);
or U7834 (N_7834,N_6564,N_6112);
and U7835 (N_7835,N_6242,N_6011);
nor U7836 (N_7836,N_6067,N_6596);
or U7837 (N_7837,N_6338,N_6537);
and U7838 (N_7838,N_6952,N_6564);
nand U7839 (N_7839,N_6017,N_6944);
xor U7840 (N_7840,N_6310,N_6583);
or U7841 (N_7841,N_6114,N_6048);
nand U7842 (N_7842,N_6855,N_6963);
and U7843 (N_7843,N_6583,N_6671);
nand U7844 (N_7844,N_6640,N_6544);
or U7845 (N_7845,N_6568,N_6009);
or U7846 (N_7846,N_6988,N_6114);
and U7847 (N_7847,N_6007,N_6334);
nand U7848 (N_7848,N_6283,N_6625);
or U7849 (N_7849,N_6600,N_6383);
or U7850 (N_7850,N_6659,N_6123);
nand U7851 (N_7851,N_6081,N_6781);
and U7852 (N_7852,N_6040,N_6668);
or U7853 (N_7853,N_6052,N_6033);
nand U7854 (N_7854,N_6438,N_6656);
or U7855 (N_7855,N_6310,N_6419);
or U7856 (N_7856,N_6591,N_6343);
and U7857 (N_7857,N_6025,N_6222);
nor U7858 (N_7858,N_6351,N_6932);
and U7859 (N_7859,N_6616,N_6536);
nor U7860 (N_7860,N_6546,N_6093);
or U7861 (N_7861,N_6029,N_6659);
nor U7862 (N_7862,N_6275,N_6881);
and U7863 (N_7863,N_6989,N_6570);
and U7864 (N_7864,N_6856,N_6776);
nor U7865 (N_7865,N_6934,N_6664);
nor U7866 (N_7866,N_6398,N_6375);
and U7867 (N_7867,N_6380,N_6391);
nand U7868 (N_7868,N_6829,N_6158);
nand U7869 (N_7869,N_6938,N_6098);
nand U7870 (N_7870,N_6176,N_6198);
nand U7871 (N_7871,N_6774,N_6621);
or U7872 (N_7872,N_6885,N_6979);
nand U7873 (N_7873,N_6319,N_6173);
and U7874 (N_7874,N_6910,N_6177);
xor U7875 (N_7875,N_6401,N_6839);
nand U7876 (N_7876,N_6560,N_6918);
or U7877 (N_7877,N_6396,N_6557);
and U7878 (N_7878,N_6318,N_6319);
and U7879 (N_7879,N_6146,N_6364);
nand U7880 (N_7880,N_6465,N_6216);
nor U7881 (N_7881,N_6356,N_6467);
and U7882 (N_7882,N_6525,N_6518);
nor U7883 (N_7883,N_6052,N_6709);
or U7884 (N_7884,N_6106,N_6667);
and U7885 (N_7885,N_6240,N_6802);
and U7886 (N_7886,N_6519,N_6600);
or U7887 (N_7887,N_6551,N_6785);
or U7888 (N_7888,N_6061,N_6073);
and U7889 (N_7889,N_6284,N_6575);
or U7890 (N_7890,N_6612,N_6491);
or U7891 (N_7891,N_6922,N_6197);
xnor U7892 (N_7892,N_6254,N_6875);
nand U7893 (N_7893,N_6402,N_6072);
or U7894 (N_7894,N_6812,N_6627);
and U7895 (N_7895,N_6926,N_6256);
and U7896 (N_7896,N_6219,N_6167);
nand U7897 (N_7897,N_6613,N_6810);
and U7898 (N_7898,N_6656,N_6356);
or U7899 (N_7899,N_6299,N_6629);
nor U7900 (N_7900,N_6312,N_6430);
nand U7901 (N_7901,N_6498,N_6788);
or U7902 (N_7902,N_6415,N_6421);
nor U7903 (N_7903,N_6792,N_6459);
or U7904 (N_7904,N_6434,N_6376);
or U7905 (N_7905,N_6374,N_6447);
or U7906 (N_7906,N_6618,N_6454);
nor U7907 (N_7907,N_6368,N_6663);
nand U7908 (N_7908,N_6378,N_6389);
nor U7909 (N_7909,N_6019,N_6676);
nor U7910 (N_7910,N_6220,N_6112);
nor U7911 (N_7911,N_6241,N_6642);
or U7912 (N_7912,N_6875,N_6240);
xnor U7913 (N_7913,N_6946,N_6087);
and U7914 (N_7914,N_6228,N_6499);
and U7915 (N_7915,N_6754,N_6239);
and U7916 (N_7916,N_6541,N_6821);
nand U7917 (N_7917,N_6936,N_6976);
nor U7918 (N_7918,N_6481,N_6169);
nor U7919 (N_7919,N_6474,N_6624);
or U7920 (N_7920,N_6174,N_6469);
and U7921 (N_7921,N_6541,N_6334);
nor U7922 (N_7922,N_6587,N_6223);
and U7923 (N_7923,N_6932,N_6159);
nand U7924 (N_7924,N_6849,N_6903);
nand U7925 (N_7925,N_6330,N_6465);
or U7926 (N_7926,N_6616,N_6786);
and U7927 (N_7927,N_6106,N_6658);
and U7928 (N_7928,N_6583,N_6922);
and U7929 (N_7929,N_6585,N_6333);
nor U7930 (N_7930,N_6684,N_6745);
or U7931 (N_7931,N_6349,N_6702);
or U7932 (N_7932,N_6785,N_6666);
and U7933 (N_7933,N_6118,N_6283);
or U7934 (N_7934,N_6509,N_6431);
nand U7935 (N_7935,N_6010,N_6714);
and U7936 (N_7936,N_6357,N_6599);
nand U7937 (N_7937,N_6080,N_6060);
nand U7938 (N_7938,N_6403,N_6995);
and U7939 (N_7939,N_6072,N_6533);
and U7940 (N_7940,N_6074,N_6505);
and U7941 (N_7941,N_6656,N_6564);
nor U7942 (N_7942,N_6141,N_6774);
and U7943 (N_7943,N_6328,N_6366);
and U7944 (N_7944,N_6722,N_6314);
and U7945 (N_7945,N_6969,N_6748);
nor U7946 (N_7946,N_6527,N_6961);
or U7947 (N_7947,N_6097,N_6868);
and U7948 (N_7948,N_6268,N_6864);
nor U7949 (N_7949,N_6543,N_6024);
nand U7950 (N_7950,N_6004,N_6580);
and U7951 (N_7951,N_6492,N_6792);
nor U7952 (N_7952,N_6641,N_6231);
nor U7953 (N_7953,N_6317,N_6544);
nand U7954 (N_7954,N_6411,N_6954);
nor U7955 (N_7955,N_6343,N_6388);
or U7956 (N_7956,N_6041,N_6034);
and U7957 (N_7957,N_6395,N_6310);
and U7958 (N_7958,N_6855,N_6664);
nand U7959 (N_7959,N_6551,N_6610);
and U7960 (N_7960,N_6771,N_6800);
nand U7961 (N_7961,N_6802,N_6232);
nor U7962 (N_7962,N_6027,N_6759);
nor U7963 (N_7963,N_6584,N_6176);
or U7964 (N_7964,N_6430,N_6585);
nand U7965 (N_7965,N_6265,N_6015);
nor U7966 (N_7966,N_6100,N_6716);
nor U7967 (N_7967,N_6680,N_6784);
nand U7968 (N_7968,N_6091,N_6213);
nand U7969 (N_7969,N_6671,N_6220);
nor U7970 (N_7970,N_6871,N_6460);
nand U7971 (N_7971,N_6169,N_6017);
and U7972 (N_7972,N_6447,N_6347);
and U7973 (N_7973,N_6001,N_6443);
nand U7974 (N_7974,N_6385,N_6897);
or U7975 (N_7975,N_6778,N_6822);
or U7976 (N_7976,N_6983,N_6825);
nand U7977 (N_7977,N_6512,N_6829);
nor U7978 (N_7978,N_6881,N_6223);
and U7979 (N_7979,N_6243,N_6456);
nand U7980 (N_7980,N_6973,N_6689);
and U7981 (N_7981,N_6075,N_6034);
nor U7982 (N_7982,N_6562,N_6498);
nor U7983 (N_7983,N_6298,N_6561);
and U7984 (N_7984,N_6325,N_6885);
or U7985 (N_7985,N_6873,N_6693);
or U7986 (N_7986,N_6911,N_6950);
or U7987 (N_7987,N_6689,N_6111);
nand U7988 (N_7988,N_6259,N_6737);
nand U7989 (N_7989,N_6386,N_6003);
nand U7990 (N_7990,N_6282,N_6309);
and U7991 (N_7991,N_6722,N_6389);
and U7992 (N_7992,N_6715,N_6287);
nor U7993 (N_7993,N_6650,N_6784);
nor U7994 (N_7994,N_6252,N_6716);
nand U7995 (N_7995,N_6325,N_6617);
and U7996 (N_7996,N_6915,N_6637);
xor U7997 (N_7997,N_6975,N_6579);
nand U7998 (N_7998,N_6607,N_6831);
nor U7999 (N_7999,N_6028,N_6678);
nor U8000 (N_8000,N_7679,N_7884);
nand U8001 (N_8001,N_7661,N_7330);
or U8002 (N_8002,N_7920,N_7638);
nor U8003 (N_8003,N_7111,N_7314);
or U8004 (N_8004,N_7722,N_7366);
nand U8005 (N_8005,N_7121,N_7467);
nand U8006 (N_8006,N_7685,N_7200);
nand U8007 (N_8007,N_7151,N_7234);
nor U8008 (N_8008,N_7014,N_7710);
or U8009 (N_8009,N_7952,N_7687);
nor U8010 (N_8010,N_7201,N_7398);
or U8011 (N_8011,N_7339,N_7630);
nand U8012 (N_8012,N_7831,N_7423);
nor U8013 (N_8013,N_7525,N_7532);
nand U8014 (N_8014,N_7108,N_7391);
and U8015 (N_8015,N_7678,N_7642);
or U8016 (N_8016,N_7723,N_7916);
nand U8017 (N_8017,N_7349,N_7477);
and U8018 (N_8018,N_7033,N_7341);
nand U8019 (N_8019,N_7793,N_7371);
nor U8020 (N_8020,N_7965,N_7148);
nor U8021 (N_8021,N_7269,N_7196);
or U8022 (N_8022,N_7316,N_7376);
and U8023 (N_8023,N_7069,N_7951);
and U8024 (N_8024,N_7641,N_7946);
nand U8025 (N_8025,N_7870,N_7759);
nor U8026 (N_8026,N_7807,N_7984);
and U8027 (N_8027,N_7011,N_7394);
nor U8028 (N_8028,N_7516,N_7767);
nor U8029 (N_8029,N_7898,N_7303);
nand U8030 (N_8030,N_7610,N_7425);
xnor U8031 (N_8031,N_7671,N_7526);
nand U8032 (N_8032,N_7194,N_7023);
and U8033 (N_8033,N_7596,N_7067);
or U8034 (N_8034,N_7748,N_7862);
nor U8035 (N_8035,N_7060,N_7044);
nor U8036 (N_8036,N_7189,N_7064);
or U8037 (N_8037,N_7774,N_7853);
nor U8038 (N_8038,N_7321,N_7607);
nor U8039 (N_8039,N_7876,N_7606);
or U8040 (N_8040,N_7505,N_7833);
nor U8041 (N_8041,N_7185,N_7739);
or U8042 (N_8042,N_7806,N_7318);
nand U8043 (N_8043,N_7496,N_7810);
and U8044 (N_8044,N_7438,N_7115);
or U8045 (N_8045,N_7621,N_7620);
and U8046 (N_8046,N_7789,N_7363);
and U8047 (N_8047,N_7122,N_7094);
or U8048 (N_8048,N_7420,N_7074);
nor U8049 (N_8049,N_7514,N_7930);
and U8050 (N_8050,N_7478,N_7821);
xnor U8051 (N_8051,N_7163,N_7940);
or U8052 (N_8052,N_7971,N_7721);
nor U8053 (N_8053,N_7399,N_7994);
or U8054 (N_8054,N_7493,N_7003);
or U8055 (N_8055,N_7714,N_7113);
or U8056 (N_8056,N_7960,N_7646);
or U8057 (N_8057,N_7838,N_7312);
xor U8058 (N_8058,N_7707,N_7640);
nand U8059 (N_8059,N_7127,N_7028);
nand U8060 (N_8060,N_7764,N_7631);
nor U8061 (N_8061,N_7665,N_7315);
or U8062 (N_8062,N_7842,N_7024);
nor U8063 (N_8063,N_7490,N_7791);
nor U8064 (N_8064,N_7273,N_7563);
nand U8065 (N_8065,N_7928,N_7480);
or U8066 (N_8066,N_7095,N_7265);
nor U8067 (N_8067,N_7468,N_7908);
or U8068 (N_8068,N_7763,N_7183);
nand U8069 (N_8069,N_7174,N_7677);
or U8070 (N_8070,N_7123,N_7998);
or U8071 (N_8071,N_7531,N_7547);
or U8072 (N_8072,N_7608,N_7843);
and U8073 (N_8073,N_7344,N_7465);
nor U8074 (N_8074,N_7832,N_7818);
nor U8075 (N_8075,N_7839,N_7229);
nor U8076 (N_8076,N_7230,N_7849);
and U8077 (N_8077,N_7829,N_7102);
nor U8078 (N_8078,N_7755,N_7356);
nor U8079 (N_8079,N_7790,N_7348);
nand U8080 (N_8080,N_7456,N_7879);
or U8081 (N_8081,N_7997,N_7735);
or U8082 (N_8082,N_7084,N_7373);
nand U8083 (N_8083,N_7886,N_7482);
and U8084 (N_8084,N_7006,N_7851);
nor U8085 (N_8085,N_7651,N_7897);
nand U8086 (N_8086,N_7645,N_7912);
or U8087 (N_8087,N_7624,N_7180);
or U8088 (N_8088,N_7100,N_7057);
nor U8089 (N_8089,N_7938,N_7383);
and U8090 (N_8090,N_7561,N_7082);
and U8091 (N_8091,N_7684,N_7860);
xor U8092 (N_8092,N_7519,N_7937);
and U8093 (N_8093,N_7109,N_7125);
nand U8094 (N_8094,N_7333,N_7177);
and U8095 (N_8095,N_7439,N_7720);
or U8096 (N_8096,N_7513,N_7257);
nor U8097 (N_8097,N_7548,N_7901);
nand U8098 (N_8098,N_7087,N_7129);
and U8099 (N_8099,N_7429,N_7051);
nor U8100 (N_8100,N_7116,N_7184);
nor U8101 (N_8101,N_7156,N_7291);
nand U8102 (N_8102,N_7107,N_7594);
nor U8103 (N_8103,N_7076,N_7599);
and U8104 (N_8104,N_7390,N_7800);
and U8105 (N_8105,N_7411,N_7470);
and U8106 (N_8106,N_7988,N_7784);
xor U8107 (N_8107,N_7292,N_7696);
xnor U8108 (N_8108,N_7702,N_7388);
nand U8109 (N_8109,N_7947,N_7981);
and U8110 (N_8110,N_7535,N_7559);
or U8111 (N_8111,N_7214,N_7276);
nor U8112 (N_8112,N_7086,N_7452);
and U8113 (N_8113,N_7463,N_7917);
or U8114 (N_8114,N_7217,N_7541);
nor U8115 (N_8115,N_7048,N_7885);
nor U8116 (N_8116,N_7828,N_7091);
or U8117 (N_8117,N_7002,N_7805);
or U8118 (N_8118,N_7726,N_7811);
nor U8119 (N_8119,N_7018,N_7445);
nand U8120 (N_8120,N_7932,N_7106);
or U8121 (N_8121,N_7248,N_7085);
nand U8122 (N_8122,N_7733,N_7058);
nand U8123 (N_8123,N_7978,N_7695);
nand U8124 (N_8124,N_7309,N_7042);
nor U8125 (N_8125,N_7814,N_7510);
or U8126 (N_8126,N_7258,N_7244);
or U8127 (N_8127,N_7138,N_7637);
and U8128 (N_8128,N_7492,N_7841);
or U8129 (N_8129,N_7499,N_7246);
nand U8130 (N_8130,N_7374,N_7626);
or U8131 (N_8131,N_7577,N_7537);
and U8132 (N_8132,N_7893,N_7158);
and U8133 (N_8133,N_7145,N_7591);
or U8134 (N_8134,N_7495,N_7632);
nor U8135 (N_8135,N_7511,N_7779);
nand U8136 (N_8136,N_7694,N_7558);
nor U8137 (N_8137,N_7169,N_7046);
and U8138 (N_8138,N_7536,N_7416);
or U8139 (N_8139,N_7012,N_7055);
nor U8140 (N_8140,N_7080,N_7555);
nor U8141 (N_8141,N_7458,N_7355);
and U8142 (N_8142,N_7802,N_7208);
nor U8143 (N_8143,N_7777,N_7697);
or U8144 (N_8144,N_7215,N_7137);
and U8145 (N_8145,N_7279,N_7464);
nand U8146 (N_8146,N_7290,N_7858);
nor U8147 (N_8147,N_7845,N_7995);
nor U8148 (N_8148,N_7284,N_7350);
or U8149 (N_8149,N_7422,N_7775);
and U8150 (N_8150,N_7240,N_7052);
nor U8151 (N_8151,N_7899,N_7220);
and U8152 (N_8152,N_7746,N_7538);
nand U8153 (N_8153,N_7877,N_7408);
and U8154 (N_8154,N_7396,N_7530);
nand U8155 (N_8155,N_7954,N_7799);
or U8156 (N_8156,N_7262,N_7083);
nor U8157 (N_8157,N_7990,N_7668);
or U8158 (N_8158,N_7529,N_7583);
or U8159 (N_8159,N_7955,N_7099);
or U8160 (N_8160,N_7706,N_7238);
or U8161 (N_8161,N_7323,N_7313);
and U8162 (N_8162,N_7424,N_7427);
nor U8163 (N_8163,N_7079,N_7268);
or U8164 (N_8164,N_7415,N_7073);
and U8165 (N_8165,N_7562,N_7762);
and U8166 (N_8166,N_7534,N_7343);
nand U8167 (N_8167,N_7816,N_7331);
or U8168 (N_8168,N_7022,N_7689);
nand U8169 (N_8169,N_7466,N_7801);
and U8170 (N_8170,N_7013,N_7050);
or U8171 (N_8171,N_7370,N_7662);
nor U8172 (N_8172,N_7546,N_7628);
nor U8173 (N_8173,N_7878,N_7512);
or U8174 (N_8174,N_7487,N_7068);
or U8175 (N_8175,N_7911,N_7092);
and U8176 (N_8176,N_7426,N_7400);
or U8177 (N_8177,N_7629,N_7406);
or U8178 (N_8178,N_7745,N_7327);
or U8179 (N_8179,N_7325,N_7719);
nand U8180 (N_8180,N_7656,N_7486);
nor U8181 (N_8181,N_7543,N_7704);
or U8182 (N_8182,N_7354,N_7923);
and U8183 (N_8183,N_7874,N_7592);
and U8184 (N_8184,N_7900,N_7840);
or U8185 (N_8185,N_7652,N_7259);
or U8186 (N_8186,N_7368,N_7700);
or U8187 (N_8187,N_7680,N_7165);
xnor U8188 (N_8188,N_7672,N_7634);
nor U8189 (N_8189,N_7854,N_7134);
nor U8190 (N_8190,N_7667,N_7617);
nand U8191 (N_8191,N_7302,N_7317);
nand U8192 (N_8192,N_7141,N_7359);
nor U8193 (N_8193,N_7020,N_7176);
nor U8194 (N_8194,N_7025,N_7773);
nand U8195 (N_8195,N_7578,N_7585);
nor U8196 (N_8196,N_7692,N_7703);
and U8197 (N_8197,N_7670,N_7682);
or U8198 (N_8198,N_7360,N_7345);
and U8199 (N_8199,N_7454,N_7298);
nand U8200 (N_8200,N_7734,N_7250);
and U8201 (N_8201,N_7280,N_7117);
or U8202 (N_8202,N_7401,N_7895);
and U8203 (N_8203,N_7889,N_7168);
or U8204 (N_8204,N_7334,N_7286);
and U8205 (N_8205,N_7455,N_7421);
nor U8206 (N_8206,N_7358,N_7846);
and U8207 (N_8207,N_7970,N_7035);
or U8208 (N_8208,N_7139,N_7342);
and U8209 (N_8209,N_7150,N_7673);
nor U8210 (N_8210,N_7847,N_7750);
and U8211 (N_8211,N_7474,N_7757);
and U8212 (N_8212,N_7962,N_7479);
and U8213 (N_8213,N_7504,N_7500);
nand U8214 (N_8214,N_7224,N_7237);
xnor U8215 (N_8215,N_7281,N_7489);
nor U8216 (N_8216,N_7007,N_7882);
nor U8217 (N_8217,N_7943,N_7709);
and U8218 (N_8218,N_7506,N_7812);
or U8219 (N_8219,N_7987,N_7484);
or U8220 (N_8220,N_7872,N_7666);
or U8221 (N_8221,N_7731,N_7471);
or U8222 (N_8222,N_7235,N_7112);
nand U8223 (N_8223,N_7077,N_7999);
nand U8224 (N_8224,N_7300,N_7868);
nor U8225 (N_8225,N_7199,N_7655);
or U8226 (N_8226,N_7473,N_7991);
and U8227 (N_8227,N_7647,N_7730);
or U8228 (N_8228,N_7549,N_7728);
nand U8229 (N_8229,N_7915,N_7865);
and U8230 (N_8230,N_7232,N_7507);
nor U8231 (N_8231,N_7924,N_7407);
nor U8232 (N_8232,N_7649,N_7557);
and U8233 (N_8233,N_7310,N_7712);
and U8234 (N_8234,N_7968,N_7888);
nand U8235 (N_8235,N_7605,N_7434);
nor U8236 (N_8236,N_7785,N_7144);
and U8237 (N_8237,N_7554,N_7056);
or U8238 (N_8238,N_7335,N_7034);
and U8239 (N_8239,N_7338,N_7732);
or U8240 (N_8240,N_7294,N_7372);
nor U8241 (N_8241,N_7615,N_7743);
and U8242 (N_8242,N_7552,N_7902);
nor U8243 (N_8243,N_7922,N_7296);
and U8244 (N_8244,N_7869,N_7336);
nor U8245 (N_8245,N_7616,N_7071);
or U8246 (N_8246,N_7119,N_7756);
nand U8247 (N_8247,N_7809,N_7942);
nor U8248 (N_8248,N_7206,N_7567);
nor U8249 (N_8249,N_7090,N_7825);
nand U8250 (N_8250,N_7494,N_7436);
or U8251 (N_8251,N_7197,N_7983);
nor U8252 (N_8252,N_7708,N_7740);
or U8253 (N_8253,N_7992,N_7266);
nor U8254 (N_8254,N_7193,N_7173);
nor U8255 (N_8255,N_7190,N_7367);
and U8256 (N_8256,N_7040,N_7658);
nand U8257 (N_8257,N_7765,N_7794);
nand U8258 (N_8258,N_7239,N_7653);
nand U8259 (N_8259,N_7819,N_7379);
and U8260 (N_8260,N_7243,N_7446);
or U8261 (N_8261,N_7021,N_7130);
or U8262 (N_8262,N_7103,N_7627);
nand U8263 (N_8263,N_7580,N_7227);
or U8264 (N_8264,N_7760,N_7573);
or U8265 (N_8265,N_7016,N_7319);
or U8266 (N_8266,N_7837,N_7956);
or U8267 (N_8267,N_7167,N_7636);
and U8268 (N_8268,N_7982,N_7412);
or U8269 (N_8269,N_7228,N_7170);
and U8270 (N_8270,N_7075,N_7146);
xor U8271 (N_8271,N_7587,N_7875);
nand U8272 (N_8272,N_7469,N_7518);
or U8273 (N_8273,N_7392,N_7676);
and U8274 (N_8274,N_7282,N_7261);
nor U8275 (N_8275,N_7958,N_7972);
and U8276 (N_8276,N_7934,N_7861);
or U8277 (N_8277,N_7311,N_7571);
or U8278 (N_8278,N_7826,N_7718);
and U8279 (N_8279,N_7569,N_7797);
nor U8280 (N_8280,N_7772,N_7769);
and U8281 (N_8281,N_7254,N_7517);
xor U8282 (N_8282,N_7045,N_7980);
or U8283 (N_8283,N_7669,N_7009);
or U8284 (N_8284,N_7919,N_7114);
or U8285 (N_8285,N_7498,N_7950);
or U8286 (N_8286,N_7110,N_7699);
and U8287 (N_8287,N_7149,N_7223);
nand U8288 (N_8288,N_7365,N_7568);
and U8289 (N_8289,N_7017,N_7979);
nand U8290 (N_8290,N_7043,N_7945);
nand U8291 (N_8291,N_7225,N_7140);
or U8292 (N_8292,N_7483,N_7857);
and U8293 (N_8293,N_7332,N_7172);
and U8294 (N_8294,N_7859,N_7786);
and U8295 (N_8295,N_7126,N_7715);
nor U8296 (N_8296,N_7595,N_7804);
or U8297 (N_8297,N_7939,N_7242);
nand U8298 (N_8298,N_7509,N_7289);
and U8299 (N_8299,N_7864,N_7202);
nor U8300 (N_8300,N_7966,N_7540);
and U8301 (N_8301,N_7059,N_7560);
or U8302 (N_8302,N_7996,N_7211);
nand U8303 (N_8303,N_7570,N_7346);
and U8304 (N_8304,N_7161,N_7941);
or U8305 (N_8305,N_7575,N_7787);
nand U8306 (N_8306,N_7503,N_7328);
nand U8307 (N_8307,N_7263,N_7910);
and U8308 (N_8308,N_7593,N_7221);
xor U8309 (N_8309,N_7926,N_7041);
or U8310 (N_8310,N_7191,N_7418);
and U8311 (N_8311,N_7096,N_7815);
and U8312 (N_8312,N_7929,N_7004);
and U8313 (N_8313,N_7397,N_7528);
nand U8314 (N_8314,N_7822,N_7729);
nand U8315 (N_8315,N_7551,N_7681);
nand U8316 (N_8316,N_7836,N_7625);
nor U8317 (N_8317,N_7753,N_7586);
or U8318 (N_8318,N_7308,N_7476);
xor U8319 (N_8319,N_7295,N_7959);
and U8320 (N_8320,N_7175,N_7188);
or U8321 (N_8321,N_7848,N_7808);
or U8322 (N_8322,N_7351,N_7038);
or U8323 (N_8323,N_7347,N_7824);
nand U8324 (N_8324,N_7460,N_7431);
and U8325 (N_8325,N_7181,N_7545);
and U8326 (N_8326,N_7449,N_7241);
nor U8327 (N_8327,N_7036,N_7001);
nand U8328 (N_8328,N_7906,N_7880);
nor U8329 (N_8329,N_7604,N_7236);
nor U8330 (N_8330,N_7914,N_7362);
and U8331 (N_8331,N_7780,N_7887);
and U8332 (N_8332,N_7603,N_7131);
and U8333 (N_8333,N_7522,N_7896);
nor U8334 (N_8334,N_7993,N_7264);
nand U8335 (N_8335,N_7985,N_7711);
xor U8336 (N_8336,N_7093,N_7231);
and U8337 (N_8337,N_7781,N_7904);
or U8338 (N_8338,N_7986,N_7834);
nor U8339 (N_8339,N_7737,N_7270);
nor U8340 (N_8340,N_7701,N_7648);
and U8341 (N_8341,N_7192,N_7142);
and U8342 (N_8342,N_7053,N_7299);
nand U8343 (N_8343,N_7222,N_7967);
nor U8344 (N_8344,N_7247,N_7873);
and U8345 (N_8345,N_7623,N_7271);
and U8346 (N_8346,N_7933,N_7143);
nor U8347 (N_8347,N_7584,N_7524);
or U8348 (N_8348,N_7612,N_7579);
or U8349 (N_8349,N_7566,N_7961);
or U8350 (N_8350,N_7783,N_7520);
and U8351 (N_8351,N_7830,N_7639);
or U8352 (N_8352,N_7207,N_7778);
nand U8353 (N_8353,N_7361,N_7384);
nor U8354 (N_8354,N_7622,N_7159);
xor U8355 (N_8355,N_7657,N_7686);
and U8356 (N_8356,N_7798,N_7754);
and U8357 (N_8357,N_7963,N_7251);
nand U8358 (N_8358,N_7909,N_7049);
and U8359 (N_8359,N_7758,N_7061);
or U8360 (N_8360,N_7442,N_7633);
or U8361 (N_8361,N_7891,N_7405);
or U8362 (N_8362,N_7213,N_7813);
nand U8363 (N_8363,N_7660,N_7019);
xnor U8364 (N_8364,N_7031,N_7752);
and U8365 (N_8365,N_7154,N_7501);
nand U8366 (N_8366,N_7380,N_7650);
and U8367 (N_8367,N_7964,N_7936);
or U8368 (N_8368,N_7457,N_7433);
nor U8369 (N_8369,N_7957,N_7913);
nor U8370 (N_8370,N_7435,N_7437);
and U8371 (N_8371,N_7850,N_7856);
and U8372 (N_8372,N_7413,N_7508);
nand U8373 (N_8373,N_7609,N_7205);
and U8374 (N_8374,N_7226,N_7588);
and U8375 (N_8375,N_7428,N_7741);
nand U8376 (N_8376,N_7324,N_7385);
or U8377 (N_8377,N_7133,N_7550);
nor U8378 (N_8378,N_7817,N_7152);
or U8379 (N_8379,N_7287,N_7441);
and U8380 (N_8380,N_7182,N_7523);
or U8381 (N_8381,N_7304,N_7481);
and U8382 (N_8382,N_7749,N_7611);
or U8383 (N_8383,N_7403,N_7256);
or U8384 (N_8384,N_7120,N_7472);
nand U8385 (N_8385,N_7005,N_7892);
nand U8386 (N_8386,N_7944,N_7101);
and U8387 (N_8387,N_7614,N_7921);
and U8388 (N_8388,N_7179,N_7063);
nor U8389 (N_8389,N_7782,N_7104);
nor U8390 (N_8390,N_7147,N_7098);
or U8391 (N_8391,N_7015,N_7485);
nor U8392 (N_8392,N_7770,N_7212);
or U8393 (N_8393,N_7301,N_7565);
xor U8394 (N_8394,N_7275,N_7274);
nor U8395 (N_8395,N_7448,N_7553);
nor U8396 (N_8396,N_7440,N_7564);
or U8397 (N_8397,N_7105,N_7124);
and U8398 (N_8398,N_7589,N_7432);
xor U8399 (N_8399,N_7417,N_7977);
or U8400 (N_8400,N_7187,N_7717);
or U8401 (N_8401,N_7277,N_7855);
or U8402 (N_8402,N_7576,N_7690);
or U8403 (N_8403,N_7903,N_7307);
nand U8404 (N_8404,N_7881,N_7157);
xnor U8405 (N_8405,N_7725,N_7894);
nand U8406 (N_8406,N_7674,N_7698);
and U8407 (N_8407,N_7796,N_7572);
nand U8408 (N_8408,N_7210,N_7382);
or U8409 (N_8409,N_7032,N_7613);
nor U8410 (N_8410,N_7381,N_7948);
and U8411 (N_8411,N_7026,N_7683);
or U8412 (N_8412,N_7393,N_7663);
nor U8413 (N_8413,N_7527,N_7402);
nor U8414 (N_8414,N_7047,N_7713);
nor U8415 (N_8415,N_7744,N_7820);
nand U8416 (N_8416,N_7975,N_7218);
nor U8417 (N_8417,N_7203,N_7724);
or U8418 (N_8418,N_7377,N_7705);
nor U8419 (N_8419,N_7443,N_7675);
nand U8420 (N_8420,N_7027,N_7643);
nor U8421 (N_8421,N_7386,N_7453);
nand U8422 (N_8422,N_7375,N_7931);
or U8423 (N_8423,N_7883,N_7581);
or U8424 (N_8424,N_7539,N_7409);
nand U8425 (N_8425,N_7867,N_7267);
nand U8426 (N_8426,N_7204,N_7556);
nand U8427 (N_8427,N_7688,N_7160);
nor U8428 (N_8428,N_7444,N_7450);
nor U8429 (N_8429,N_7000,N_7166);
nand U8430 (N_8430,N_7601,N_7488);
or U8431 (N_8431,N_7272,N_7742);
nand U8432 (N_8432,N_7835,N_7369);
nand U8433 (N_8433,N_7866,N_7378);
or U8434 (N_8434,N_7574,N_7771);
nand U8435 (N_8435,N_7738,N_7404);
xor U8436 (N_8436,N_7618,N_7788);
or U8437 (N_8437,N_7430,N_7419);
nor U8438 (N_8438,N_7907,N_7515);
nand U8439 (N_8439,N_7364,N_7890);
nand U8440 (N_8440,N_7598,N_7927);
nor U8441 (N_8441,N_7054,N_7953);
nand U8442 (N_8442,N_7654,N_7497);
xor U8443 (N_8443,N_7322,N_7844);
and U8444 (N_8444,N_7337,N_7326);
nor U8445 (N_8445,N_7297,N_7039);
nor U8446 (N_8446,N_7072,N_7340);
nor U8447 (N_8447,N_7255,N_7153);
nand U8448 (N_8448,N_7245,N_7475);
nor U8449 (N_8449,N_7065,N_7974);
and U8450 (N_8450,N_7164,N_7823);
or U8451 (N_8451,N_7644,N_7357);
or U8452 (N_8452,N_7078,N_7447);
nand U8453 (N_8453,N_7097,N_7353);
or U8454 (N_8454,N_7410,N_7219);
and U8455 (N_8455,N_7293,N_7542);
nor U8456 (N_8456,N_7795,N_7602);
or U8457 (N_8457,N_7521,N_7155);
nor U8458 (N_8458,N_7260,N_7935);
nand U8459 (N_8459,N_7306,N_7088);
or U8460 (N_8460,N_7597,N_7305);
nand U8461 (N_8461,N_7544,N_7389);
and U8462 (N_8462,N_7582,N_7209);
nand U8463 (N_8463,N_7969,N_7252);
or U8464 (N_8464,N_7253,N_7491);
nand U8465 (N_8465,N_7352,N_7462);
and U8466 (N_8466,N_7030,N_7288);
nand U8467 (N_8467,N_7776,N_7329);
nand U8468 (N_8468,N_7852,N_7089);
nor U8469 (N_8469,N_7905,N_7233);
nor U8470 (N_8470,N_7395,N_7716);
xor U8471 (N_8471,N_7761,N_7925);
or U8472 (N_8472,N_7635,N_7693);
nor U8473 (N_8473,N_7081,N_7451);
nand U8474 (N_8474,N_7070,N_7195);
nand U8475 (N_8475,N_7727,N_7136);
nand U8476 (N_8476,N_7803,N_7128);
nor U8477 (N_8477,N_7502,N_7863);
nand U8478 (N_8478,N_7171,N_7029);
or U8479 (N_8479,N_7216,N_7198);
and U8480 (N_8480,N_7766,N_7973);
nor U8481 (N_8481,N_7008,N_7600);
nand U8482 (N_8482,N_7010,N_7949);
nor U8483 (N_8483,N_7871,N_7320);
nand U8484 (N_8484,N_7414,N_7736);
and U8485 (N_8485,N_7619,N_7178);
and U8486 (N_8486,N_7118,N_7461);
or U8487 (N_8487,N_7459,N_7249);
and U8488 (N_8488,N_7283,N_7989);
and U8489 (N_8489,N_7918,N_7691);
or U8490 (N_8490,N_7387,N_7037);
xor U8491 (N_8491,N_7135,N_7827);
nand U8492 (N_8492,N_7186,N_7659);
or U8493 (N_8493,N_7747,N_7285);
and U8494 (N_8494,N_7768,N_7751);
nor U8495 (N_8495,N_7792,N_7533);
and U8496 (N_8496,N_7062,N_7132);
nor U8497 (N_8497,N_7590,N_7162);
nor U8498 (N_8498,N_7664,N_7278);
nand U8499 (N_8499,N_7066,N_7976);
nor U8500 (N_8500,N_7055,N_7001);
or U8501 (N_8501,N_7764,N_7634);
nand U8502 (N_8502,N_7868,N_7311);
and U8503 (N_8503,N_7875,N_7575);
or U8504 (N_8504,N_7677,N_7147);
or U8505 (N_8505,N_7228,N_7099);
nor U8506 (N_8506,N_7659,N_7395);
nand U8507 (N_8507,N_7081,N_7116);
and U8508 (N_8508,N_7540,N_7982);
and U8509 (N_8509,N_7145,N_7238);
nor U8510 (N_8510,N_7397,N_7312);
and U8511 (N_8511,N_7776,N_7863);
nand U8512 (N_8512,N_7375,N_7016);
nand U8513 (N_8513,N_7965,N_7418);
or U8514 (N_8514,N_7197,N_7781);
nor U8515 (N_8515,N_7353,N_7759);
nor U8516 (N_8516,N_7925,N_7189);
nand U8517 (N_8517,N_7239,N_7536);
nor U8518 (N_8518,N_7613,N_7015);
nor U8519 (N_8519,N_7022,N_7017);
and U8520 (N_8520,N_7202,N_7303);
nand U8521 (N_8521,N_7866,N_7137);
nand U8522 (N_8522,N_7306,N_7424);
nand U8523 (N_8523,N_7937,N_7878);
or U8524 (N_8524,N_7905,N_7247);
and U8525 (N_8525,N_7155,N_7284);
nor U8526 (N_8526,N_7591,N_7405);
and U8527 (N_8527,N_7502,N_7675);
nor U8528 (N_8528,N_7786,N_7783);
or U8529 (N_8529,N_7998,N_7562);
or U8530 (N_8530,N_7986,N_7623);
or U8531 (N_8531,N_7354,N_7950);
nand U8532 (N_8532,N_7174,N_7964);
xnor U8533 (N_8533,N_7348,N_7803);
nand U8534 (N_8534,N_7391,N_7560);
and U8535 (N_8535,N_7423,N_7853);
or U8536 (N_8536,N_7191,N_7373);
nor U8537 (N_8537,N_7804,N_7598);
nor U8538 (N_8538,N_7659,N_7008);
and U8539 (N_8539,N_7608,N_7170);
nor U8540 (N_8540,N_7497,N_7106);
and U8541 (N_8541,N_7338,N_7762);
or U8542 (N_8542,N_7736,N_7381);
nor U8543 (N_8543,N_7421,N_7548);
and U8544 (N_8544,N_7006,N_7521);
nor U8545 (N_8545,N_7624,N_7247);
nand U8546 (N_8546,N_7066,N_7448);
and U8547 (N_8547,N_7733,N_7631);
xnor U8548 (N_8548,N_7704,N_7387);
and U8549 (N_8549,N_7972,N_7089);
and U8550 (N_8550,N_7923,N_7015);
nor U8551 (N_8551,N_7084,N_7361);
nand U8552 (N_8552,N_7690,N_7342);
nand U8553 (N_8553,N_7230,N_7036);
or U8554 (N_8554,N_7676,N_7791);
and U8555 (N_8555,N_7070,N_7107);
nor U8556 (N_8556,N_7017,N_7352);
nor U8557 (N_8557,N_7858,N_7639);
and U8558 (N_8558,N_7310,N_7559);
or U8559 (N_8559,N_7463,N_7962);
nand U8560 (N_8560,N_7284,N_7153);
nand U8561 (N_8561,N_7986,N_7609);
nand U8562 (N_8562,N_7459,N_7124);
or U8563 (N_8563,N_7856,N_7198);
and U8564 (N_8564,N_7602,N_7976);
nor U8565 (N_8565,N_7305,N_7716);
nor U8566 (N_8566,N_7095,N_7345);
nor U8567 (N_8567,N_7965,N_7442);
or U8568 (N_8568,N_7617,N_7724);
xor U8569 (N_8569,N_7979,N_7577);
nand U8570 (N_8570,N_7497,N_7329);
and U8571 (N_8571,N_7395,N_7443);
or U8572 (N_8572,N_7607,N_7767);
nor U8573 (N_8573,N_7871,N_7851);
nor U8574 (N_8574,N_7383,N_7895);
nand U8575 (N_8575,N_7493,N_7976);
and U8576 (N_8576,N_7925,N_7889);
or U8577 (N_8577,N_7925,N_7292);
nand U8578 (N_8578,N_7672,N_7096);
nand U8579 (N_8579,N_7653,N_7055);
and U8580 (N_8580,N_7728,N_7797);
nor U8581 (N_8581,N_7012,N_7575);
nand U8582 (N_8582,N_7486,N_7047);
and U8583 (N_8583,N_7371,N_7324);
nand U8584 (N_8584,N_7711,N_7921);
and U8585 (N_8585,N_7092,N_7170);
nand U8586 (N_8586,N_7675,N_7056);
nand U8587 (N_8587,N_7972,N_7878);
nand U8588 (N_8588,N_7369,N_7687);
or U8589 (N_8589,N_7357,N_7799);
and U8590 (N_8590,N_7725,N_7401);
or U8591 (N_8591,N_7090,N_7489);
and U8592 (N_8592,N_7949,N_7637);
and U8593 (N_8593,N_7103,N_7631);
nand U8594 (N_8594,N_7499,N_7102);
nand U8595 (N_8595,N_7538,N_7395);
or U8596 (N_8596,N_7027,N_7733);
nand U8597 (N_8597,N_7610,N_7173);
nand U8598 (N_8598,N_7327,N_7286);
nor U8599 (N_8599,N_7719,N_7352);
xnor U8600 (N_8600,N_7209,N_7867);
and U8601 (N_8601,N_7101,N_7673);
and U8602 (N_8602,N_7748,N_7137);
nor U8603 (N_8603,N_7888,N_7705);
and U8604 (N_8604,N_7662,N_7977);
nor U8605 (N_8605,N_7874,N_7113);
xnor U8606 (N_8606,N_7824,N_7820);
nand U8607 (N_8607,N_7289,N_7532);
nand U8608 (N_8608,N_7362,N_7864);
or U8609 (N_8609,N_7050,N_7805);
nand U8610 (N_8610,N_7624,N_7352);
nand U8611 (N_8611,N_7735,N_7854);
nand U8612 (N_8612,N_7283,N_7856);
and U8613 (N_8613,N_7671,N_7686);
and U8614 (N_8614,N_7485,N_7906);
nand U8615 (N_8615,N_7173,N_7444);
xnor U8616 (N_8616,N_7871,N_7315);
nand U8617 (N_8617,N_7728,N_7826);
nor U8618 (N_8618,N_7317,N_7038);
or U8619 (N_8619,N_7115,N_7498);
and U8620 (N_8620,N_7952,N_7526);
nand U8621 (N_8621,N_7301,N_7830);
nor U8622 (N_8622,N_7895,N_7045);
nor U8623 (N_8623,N_7682,N_7667);
or U8624 (N_8624,N_7089,N_7275);
or U8625 (N_8625,N_7393,N_7673);
nor U8626 (N_8626,N_7984,N_7129);
and U8627 (N_8627,N_7315,N_7148);
nand U8628 (N_8628,N_7922,N_7899);
and U8629 (N_8629,N_7192,N_7527);
and U8630 (N_8630,N_7753,N_7420);
nor U8631 (N_8631,N_7726,N_7273);
and U8632 (N_8632,N_7673,N_7890);
and U8633 (N_8633,N_7278,N_7616);
and U8634 (N_8634,N_7725,N_7939);
nand U8635 (N_8635,N_7897,N_7954);
or U8636 (N_8636,N_7018,N_7276);
and U8637 (N_8637,N_7130,N_7370);
nor U8638 (N_8638,N_7738,N_7791);
and U8639 (N_8639,N_7659,N_7310);
or U8640 (N_8640,N_7097,N_7005);
and U8641 (N_8641,N_7932,N_7677);
nand U8642 (N_8642,N_7928,N_7336);
or U8643 (N_8643,N_7598,N_7666);
nor U8644 (N_8644,N_7593,N_7560);
or U8645 (N_8645,N_7969,N_7235);
or U8646 (N_8646,N_7290,N_7705);
or U8647 (N_8647,N_7550,N_7241);
or U8648 (N_8648,N_7494,N_7068);
or U8649 (N_8649,N_7108,N_7258);
and U8650 (N_8650,N_7376,N_7260);
and U8651 (N_8651,N_7410,N_7537);
xor U8652 (N_8652,N_7254,N_7084);
nor U8653 (N_8653,N_7734,N_7723);
nor U8654 (N_8654,N_7726,N_7482);
and U8655 (N_8655,N_7123,N_7163);
and U8656 (N_8656,N_7498,N_7563);
nand U8657 (N_8657,N_7663,N_7062);
and U8658 (N_8658,N_7373,N_7689);
nor U8659 (N_8659,N_7210,N_7560);
and U8660 (N_8660,N_7336,N_7442);
or U8661 (N_8661,N_7209,N_7227);
nor U8662 (N_8662,N_7678,N_7102);
nand U8663 (N_8663,N_7357,N_7559);
nand U8664 (N_8664,N_7890,N_7594);
nand U8665 (N_8665,N_7065,N_7962);
and U8666 (N_8666,N_7395,N_7834);
and U8667 (N_8667,N_7161,N_7791);
or U8668 (N_8668,N_7208,N_7331);
and U8669 (N_8669,N_7598,N_7989);
and U8670 (N_8670,N_7990,N_7551);
and U8671 (N_8671,N_7723,N_7761);
and U8672 (N_8672,N_7139,N_7545);
or U8673 (N_8673,N_7936,N_7318);
or U8674 (N_8674,N_7982,N_7604);
and U8675 (N_8675,N_7481,N_7073);
and U8676 (N_8676,N_7925,N_7583);
nor U8677 (N_8677,N_7284,N_7778);
or U8678 (N_8678,N_7129,N_7619);
nand U8679 (N_8679,N_7373,N_7348);
nand U8680 (N_8680,N_7821,N_7237);
and U8681 (N_8681,N_7412,N_7491);
nor U8682 (N_8682,N_7577,N_7339);
nor U8683 (N_8683,N_7495,N_7480);
and U8684 (N_8684,N_7999,N_7792);
or U8685 (N_8685,N_7713,N_7340);
xor U8686 (N_8686,N_7269,N_7534);
and U8687 (N_8687,N_7523,N_7379);
and U8688 (N_8688,N_7246,N_7668);
or U8689 (N_8689,N_7309,N_7336);
or U8690 (N_8690,N_7300,N_7023);
nor U8691 (N_8691,N_7076,N_7519);
and U8692 (N_8692,N_7141,N_7842);
nor U8693 (N_8693,N_7781,N_7438);
nor U8694 (N_8694,N_7723,N_7898);
and U8695 (N_8695,N_7560,N_7368);
nand U8696 (N_8696,N_7094,N_7715);
and U8697 (N_8697,N_7633,N_7302);
nand U8698 (N_8698,N_7509,N_7393);
nand U8699 (N_8699,N_7159,N_7724);
nor U8700 (N_8700,N_7854,N_7821);
nand U8701 (N_8701,N_7675,N_7258);
nand U8702 (N_8702,N_7465,N_7907);
nor U8703 (N_8703,N_7643,N_7901);
or U8704 (N_8704,N_7962,N_7207);
nand U8705 (N_8705,N_7986,N_7115);
nand U8706 (N_8706,N_7918,N_7422);
and U8707 (N_8707,N_7285,N_7370);
nor U8708 (N_8708,N_7410,N_7763);
nand U8709 (N_8709,N_7970,N_7541);
nand U8710 (N_8710,N_7892,N_7209);
or U8711 (N_8711,N_7958,N_7395);
and U8712 (N_8712,N_7918,N_7223);
nor U8713 (N_8713,N_7000,N_7052);
nor U8714 (N_8714,N_7753,N_7340);
or U8715 (N_8715,N_7531,N_7003);
nand U8716 (N_8716,N_7598,N_7322);
nand U8717 (N_8717,N_7177,N_7322);
or U8718 (N_8718,N_7562,N_7398);
and U8719 (N_8719,N_7361,N_7992);
nand U8720 (N_8720,N_7136,N_7847);
and U8721 (N_8721,N_7480,N_7397);
nand U8722 (N_8722,N_7770,N_7415);
or U8723 (N_8723,N_7756,N_7924);
nand U8724 (N_8724,N_7124,N_7504);
and U8725 (N_8725,N_7352,N_7818);
or U8726 (N_8726,N_7901,N_7877);
nand U8727 (N_8727,N_7053,N_7146);
nor U8728 (N_8728,N_7874,N_7562);
nor U8729 (N_8729,N_7037,N_7179);
nor U8730 (N_8730,N_7374,N_7831);
nand U8731 (N_8731,N_7339,N_7506);
and U8732 (N_8732,N_7332,N_7816);
or U8733 (N_8733,N_7207,N_7774);
or U8734 (N_8734,N_7917,N_7280);
or U8735 (N_8735,N_7671,N_7085);
or U8736 (N_8736,N_7616,N_7340);
and U8737 (N_8737,N_7842,N_7282);
nand U8738 (N_8738,N_7135,N_7005);
or U8739 (N_8739,N_7882,N_7153);
nor U8740 (N_8740,N_7887,N_7200);
and U8741 (N_8741,N_7320,N_7565);
nor U8742 (N_8742,N_7488,N_7698);
or U8743 (N_8743,N_7991,N_7515);
and U8744 (N_8744,N_7879,N_7340);
and U8745 (N_8745,N_7089,N_7823);
nor U8746 (N_8746,N_7348,N_7991);
or U8747 (N_8747,N_7301,N_7963);
and U8748 (N_8748,N_7687,N_7292);
or U8749 (N_8749,N_7690,N_7753);
or U8750 (N_8750,N_7252,N_7469);
and U8751 (N_8751,N_7105,N_7760);
nor U8752 (N_8752,N_7376,N_7803);
nand U8753 (N_8753,N_7930,N_7184);
xor U8754 (N_8754,N_7344,N_7875);
or U8755 (N_8755,N_7859,N_7089);
or U8756 (N_8756,N_7501,N_7081);
nand U8757 (N_8757,N_7444,N_7342);
and U8758 (N_8758,N_7560,N_7696);
nor U8759 (N_8759,N_7721,N_7965);
and U8760 (N_8760,N_7294,N_7478);
or U8761 (N_8761,N_7470,N_7493);
nand U8762 (N_8762,N_7195,N_7079);
or U8763 (N_8763,N_7572,N_7259);
or U8764 (N_8764,N_7915,N_7059);
and U8765 (N_8765,N_7879,N_7955);
nor U8766 (N_8766,N_7542,N_7712);
nor U8767 (N_8767,N_7882,N_7559);
nor U8768 (N_8768,N_7555,N_7192);
and U8769 (N_8769,N_7804,N_7971);
nor U8770 (N_8770,N_7267,N_7649);
nor U8771 (N_8771,N_7024,N_7056);
or U8772 (N_8772,N_7148,N_7273);
nand U8773 (N_8773,N_7013,N_7212);
and U8774 (N_8774,N_7295,N_7677);
and U8775 (N_8775,N_7177,N_7077);
or U8776 (N_8776,N_7056,N_7470);
or U8777 (N_8777,N_7085,N_7923);
nand U8778 (N_8778,N_7670,N_7196);
nand U8779 (N_8779,N_7016,N_7258);
nand U8780 (N_8780,N_7626,N_7957);
and U8781 (N_8781,N_7573,N_7915);
nor U8782 (N_8782,N_7004,N_7878);
nor U8783 (N_8783,N_7220,N_7026);
and U8784 (N_8784,N_7923,N_7344);
and U8785 (N_8785,N_7637,N_7877);
nand U8786 (N_8786,N_7291,N_7703);
nand U8787 (N_8787,N_7798,N_7111);
nor U8788 (N_8788,N_7435,N_7026);
nor U8789 (N_8789,N_7527,N_7537);
and U8790 (N_8790,N_7397,N_7203);
or U8791 (N_8791,N_7259,N_7339);
and U8792 (N_8792,N_7984,N_7531);
or U8793 (N_8793,N_7679,N_7663);
nor U8794 (N_8794,N_7102,N_7316);
or U8795 (N_8795,N_7668,N_7114);
or U8796 (N_8796,N_7482,N_7619);
nand U8797 (N_8797,N_7972,N_7763);
nor U8798 (N_8798,N_7128,N_7780);
nor U8799 (N_8799,N_7233,N_7081);
or U8800 (N_8800,N_7744,N_7320);
or U8801 (N_8801,N_7185,N_7133);
or U8802 (N_8802,N_7885,N_7472);
and U8803 (N_8803,N_7875,N_7213);
and U8804 (N_8804,N_7229,N_7233);
nor U8805 (N_8805,N_7697,N_7854);
nand U8806 (N_8806,N_7354,N_7867);
and U8807 (N_8807,N_7341,N_7859);
xor U8808 (N_8808,N_7639,N_7519);
nor U8809 (N_8809,N_7890,N_7765);
nor U8810 (N_8810,N_7390,N_7197);
nand U8811 (N_8811,N_7752,N_7595);
or U8812 (N_8812,N_7919,N_7821);
and U8813 (N_8813,N_7268,N_7252);
and U8814 (N_8814,N_7103,N_7188);
nand U8815 (N_8815,N_7529,N_7223);
nor U8816 (N_8816,N_7230,N_7897);
or U8817 (N_8817,N_7433,N_7211);
nand U8818 (N_8818,N_7090,N_7653);
or U8819 (N_8819,N_7871,N_7920);
nand U8820 (N_8820,N_7253,N_7051);
nand U8821 (N_8821,N_7268,N_7804);
nand U8822 (N_8822,N_7768,N_7525);
nor U8823 (N_8823,N_7246,N_7532);
or U8824 (N_8824,N_7323,N_7639);
nor U8825 (N_8825,N_7540,N_7128);
or U8826 (N_8826,N_7034,N_7368);
nand U8827 (N_8827,N_7540,N_7969);
and U8828 (N_8828,N_7935,N_7147);
nor U8829 (N_8829,N_7423,N_7899);
nor U8830 (N_8830,N_7018,N_7645);
and U8831 (N_8831,N_7016,N_7751);
nand U8832 (N_8832,N_7157,N_7788);
or U8833 (N_8833,N_7446,N_7598);
nand U8834 (N_8834,N_7002,N_7391);
and U8835 (N_8835,N_7019,N_7831);
and U8836 (N_8836,N_7608,N_7676);
or U8837 (N_8837,N_7033,N_7718);
nor U8838 (N_8838,N_7505,N_7988);
nor U8839 (N_8839,N_7846,N_7500);
nand U8840 (N_8840,N_7702,N_7094);
nand U8841 (N_8841,N_7246,N_7322);
nand U8842 (N_8842,N_7701,N_7170);
nor U8843 (N_8843,N_7077,N_7600);
nand U8844 (N_8844,N_7204,N_7029);
and U8845 (N_8845,N_7552,N_7399);
or U8846 (N_8846,N_7466,N_7479);
nor U8847 (N_8847,N_7087,N_7295);
and U8848 (N_8848,N_7477,N_7064);
xor U8849 (N_8849,N_7707,N_7506);
xnor U8850 (N_8850,N_7263,N_7914);
or U8851 (N_8851,N_7100,N_7318);
or U8852 (N_8852,N_7838,N_7823);
and U8853 (N_8853,N_7880,N_7573);
nand U8854 (N_8854,N_7030,N_7630);
nand U8855 (N_8855,N_7571,N_7964);
or U8856 (N_8856,N_7509,N_7024);
and U8857 (N_8857,N_7669,N_7664);
nor U8858 (N_8858,N_7928,N_7459);
nand U8859 (N_8859,N_7140,N_7354);
xnor U8860 (N_8860,N_7859,N_7595);
nor U8861 (N_8861,N_7270,N_7701);
nor U8862 (N_8862,N_7095,N_7403);
nor U8863 (N_8863,N_7540,N_7407);
nand U8864 (N_8864,N_7958,N_7330);
nor U8865 (N_8865,N_7432,N_7419);
nor U8866 (N_8866,N_7595,N_7597);
nor U8867 (N_8867,N_7970,N_7939);
nor U8868 (N_8868,N_7106,N_7866);
and U8869 (N_8869,N_7120,N_7125);
nand U8870 (N_8870,N_7735,N_7805);
and U8871 (N_8871,N_7902,N_7960);
or U8872 (N_8872,N_7294,N_7286);
xor U8873 (N_8873,N_7169,N_7076);
and U8874 (N_8874,N_7702,N_7809);
nor U8875 (N_8875,N_7289,N_7775);
or U8876 (N_8876,N_7353,N_7755);
nor U8877 (N_8877,N_7472,N_7953);
or U8878 (N_8878,N_7860,N_7359);
or U8879 (N_8879,N_7020,N_7066);
or U8880 (N_8880,N_7291,N_7396);
and U8881 (N_8881,N_7106,N_7911);
nand U8882 (N_8882,N_7318,N_7370);
nor U8883 (N_8883,N_7758,N_7942);
nand U8884 (N_8884,N_7265,N_7267);
nand U8885 (N_8885,N_7561,N_7734);
nand U8886 (N_8886,N_7012,N_7659);
and U8887 (N_8887,N_7774,N_7854);
and U8888 (N_8888,N_7800,N_7066);
nand U8889 (N_8889,N_7884,N_7713);
and U8890 (N_8890,N_7100,N_7957);
and U8891 (N_8891,N_7449,N_7963);
nor U8892 (N_8892,N_7826,N_7594);
or U8893 (N_8893,N_7226,N_7455);
xor U8894 (N_8894,N_7114,N_7157);
or U8895 (N_8895,N_7427,N_7729);
nand U8896 (N_8896,N_7020,N_7499);
nor U8897 (N_8897,N_7101,N_7154);
nor U8898 (N_8898,N_7497,N_7425);
or U8899 (N_8899,N_7066,N_7412);
or U8900 (N_8900,N_7474,N_7414);
nor U8901 (N_8901,N_7518,N_7762);
nand U8902 (N_8902,N_7697,N_7698);
or U8903 (N_8903,N_7439,N_7328);
nand U8904 (N_8904,N_7872,N_7486);
and U8905 (N_8905,N_7321,N_7160);
or U8906 (N_8906,N_7861,N_7165);
nor U8907 (N_8907,N_7305,N_7429);
nand U8908 (N_8908,N_7742,N_7387);
nor U8909 (N_8909,N_7234,N_7913);
nor U8910 (N_8910,N_7743,N_7511);
nor U8911 (N_8911,N_7944,N_7844);
or U8912 (N_8912,N_7856,N_7145);
and U8913 (N_8913,N_7450,N_7283);
nor U8914 (N_8914,N_7487,N_7349);
or U8915 (N_8915,N_7769,N_7228);
and U8916 (N_8916,N_7565,N_7055);
xor U8917 (N_8917,N_7302,N_7162);
nor U8918 (N_8918,N_7004,N_7747);
or U8919 (N_8919,N_7134,N_7465);
and U8920 (N_8920,N_7523,N_7510);
nor U8921 (N_8921,N_7153,N_7034);
or U8922 (N_8922,N_7867,N_7770);
nor U8923 (N_8923,N_7354,N_7402);
nor U8924 (N_8924,N_7333,N_7538);
and U8925 (N_8925,N_7295,N_7514);
or U8926 (N_8926,N_7768,N_7354);
nand U8927 (N_8927,N_7013,N_7934);
and U8928 (N_8928,N_7408,N_7257);
and U8929 (N_8929,N_7710,N_7082);
nand U8930 (N_8930,N_7737,N_7117);
nand U8931 (N_8931,N_7659,N_7964);
or U8932 (N_8932,N_7629,N_7086);
and U8933 (N_8933,N_7389,N_7929);
and U8934 (N_8934,N_7502,N_7390);
and U8935 (N_8935,N_7286,N_7415);
nand U8936 (N_8936,N_7981,N_7138);
nand U8937 (N_8937,N_7525,N_7198);
nand U8938 (N_8938,N_7851,N_7760);
nor U8939 (N_8939,N_7714,N_7896);
or U8940 (N_8940,N_7987,N_7986);
and U8941 (N_8941,N_7040,N_7462);
nor U8942 (N_8942,N_7623,N_7410);
and U8943 (N_8943,N_7396,N_7511);
nand U8944 (N_8944,N_7949,N_7910);
nor U8945 (N_8945,N_7172,N_7095);
or U8946 (N_8946,N_7146,N_7259);
nand U8947 (N_8947,N_7647,N_7002);
or U8948 (N_8948,N_7694,N_7242);
and U8949 (N_8949,N_7372,N_7030);
or U8950 (N_8950,N_7047,N_7722);
or U8951 (N_8951,N_7742,N_7049);
and U8952 (N_8952,N_7296,N_7728);
nor U8953 (N_8953,N_7437,N_7062);
nand U8954 (N_8954,N_7451,N_7679);
nand U8955 (N_8955,N_7611,N_7279);
nor U8956 (N_8956,N_7097,N_7819);
and U8957 (N_8957,N_7196,N_7798);
nand U8958 (N_8958,N_7454,N_7371);
nand U8959 (N_8959,N_7221,N_7597);
nand U8960 (N_8960,N_7892,N_7980);
or U8961 (N_8961,N_7282,N_7921);
and U8962 (N_8962,N_7086,N_7449);
nor U8963 (N_8963,N_7645,N_7024);
and U8964 (N_8964,N_7802,N_7271);
nand U8965 (N_8965,N_7550,N_7042);
and U8966 (N_8966,N_7396,N_7580);
and U8967 (N_8967,N_7811,N_7209);
nand U8968 (N_8968,N_7503,N_7691);
or U8969 (N_8969,N_7518,N_7939);
nand U8970 (N_8970,N_7155,N_7539);
nand U8971 (N_8971,N_7411,N_7883);
nand U8972 (N_8972,N_7949,N_7475);
nand U8973 (N_8973,N_7374,N_7200);
nand U8974 (N_8974,N_7098,N_7271);
nand U8975 (N_8975,N_7570,N_7496);
and U8976 (N_8976,N_7565,N_7776);
and U8977 (N_8977,N_7534,N_7037);
xor U8978 (N_8978,N_7075,N_7096);
nor U8979 (N_8979,N_7323,N_7959);
nand U8980 (N_8980,N_7920,N_7466);
or U8981 (N_8981,N_7260,N_7135);
or U8982 (N_8982,N_7691,N_7304);
nand U8983 (N_8983,N_7666,N_7788);
or U8984 (N_8984,N_7296,N_7300);
nand U8985 (N_8985,N_7586,N_7730);
nor U8986 (N_8986,N_7376,N_7091);
and U8987 (N_8987,N_7622,N_7505);
or U8988 (N_8988,N_7106,N_7860);
or U8989 (N_8989,N_7938,N_7320);
nor U8990 (N_8990,N_7656,N_7563);
nand U8991 (N_8991,N_7252,N_7344);
and U8992 (N_8992,N_7589,N_7612);
and U8993 (N_8993,N_7298,N_7080);
nor U8994 (N_8994,N_7636,N_7866);
nor U8995 (N_8995,N_7676,N_7850);
nand U8996 (N_8996,N_7838,N_7156);
nor U8997 (N_8997,N_7157,N_7250);
or U8998 (N_8998,N_7642,N_7619);
and U8999 (N_8999,N_7987,N_7614);
or U9000 (N_9000,N_8240,N_8599);
xor U9001 (N_9001,N_8590,N_8508);
nand U9002 (N_9002,N_8418,N_8193);
and U9003 (N_9003,N_8271,N_8930);
nor U9004 (N_9004,N_8473,N_8184);
nor U9005 (N_9005,N_8293,N_8007);
xnor U9006 (N_9006,N_8361,N_8402);
or U9007 (N_9007,N_8167,N_8298);
nand U9008 (N_9008,N_8991,N_8660);
and U9009 (N_9009,N_8666,N_8090);
nand U9010 (N_9010,N_8408,N_8559);
xor U9011 (N_9011,N_8905,N_8828);
and U9012 (N_9012,N_8430,N_8646);
nor U9013 (N_9013,N_8683,N_8453);
nand U9014 (N_9014,N_8377,N_8650);
nor U9015 (N_9015,N_8403,N_8292);
or U9016 (N_9016,N_8416,N_8482);
or U9017 (N_9017,N_8871,N_8522);
nand U9018 (N_9018,N_8615,N_8637);
and U9019 (N_9019,N_8994,N_8182);
and U9020 (N_9020,N_8220,N_8424);
or U9021 (N_9021,N_8004,N_8947);
nand U9022 (N_9022,N_8788,N_8808);
and U9023 (N_9023,N_8100,N_8885);
or U9024 (N_9024,N_8996,N_8357);
or U9025 (N_9025,N_8029,N_8728);
nor U9026 (N_9026,N_8502,N_8688);
nand U9027 (N_9027,N_8407,N_8276);
nor U9028 (N_9028,N_8720,N_8254);
nor U9029 (N_9029,N_8513,N_8595);
nor U9030 (N_9030,N_8343,N_8040);
and U9031 (N_9031,N_8474,N_8296);
nand U9032 (N_9032,N_8777,N_8133);
nor U9033 (N_9033,N_8366,N_8297);
and U9034 (N_9034,N_8907,N_8232);
nand U9035 (N_9035,N_8628,N_8631);
nor U9036 (N_9036,N_8701,N_8739);
nor U9037 (N_9037,N_8484,N_8710);
and U9038 (N_9038,N_8510,N_8097);
and U9039 (N_9039,N_8951,N_8116);
and U9040 (N_9040,N_8517,N_8176);
and U9041 (N_9041,N_8083,N_8899);
nand U9042 (N_9042,N_8341,N_8845);
and U9043 (N_9043,N_8851,N_8051);
nor U9044 (N_9044,N_8855,N_8241);
or U9045 (N_9045,N_8867,N_8455);
or U9046 (N_9046,N_8505,N_8702);
nor U9047 (N_9047,N_8694,N_8793);
nand U9048 (N_9048,N_8955,N_8149);
nor U9049 (N_9049,N_8993,N_8865);
nand U9050 (N_9050,N_8212,N_8016);
or U9051 (N_9051,N_8236,N_8529);
nand U9052 (N_9052,N_8388,N_8620);
nand U9053 (N_9053,N_8132,N_8437);
or U9054 (N_9054,N_8331,N_8148);
nand U9055 (N_9055,N_8030,N_8180);
nor U9056 (N_9056,N_8814,N_8449);
or U9057 (N_9057,N_8527,N_8381);
nand U9058 (N_9058,N_8909,N_8669);
nand U9059 (N_9059,N_8718,N_8161);
nor U9060 (N_9060,N_8937,N_8759);
nor U9061 (N_9061,N_8664,N_8813);
nor U9062 (N_9062,N_8695,N_8948);
and U9063 (N_9063,N_8018,N_8890);
and U9064 (N_9064,N_8638,N_8641);
or U9065 (N_9065,N_8052,N_8848);
nor U9066 (N_9066,N_8112,N_8099);
nor U9067 (N_9067,N_8802,N_8945);
nor U9068 (N_9068,N_8355,N_8903);
xnor U9069 (N_9069,N_8102,N_8612);
and U9070 (N_9070,N_8094,N_8479);
nor U9071 (N_9071,N_8395,N_8401);
or U9072 (N_9072,N_8724,N_8847);
nand U9073 (N_9073,N_8226,N_8396);
nand U9074 (N_9074,N_8995,N_8797);
or U9075 (N_9075,N_8498,N_8390);
or U9076 (N_9076,N_8764,N_8481);
nand U9077 (N_9077,N_8858,N_8359);
nand U9078 (N_9078,N_8901,N_8539);
and U9079 (N_9079,N_8031,N_8274);
or U9080 (N_9080,N_8105,N_8339);
nor U9081 (N_9081,N_8487,N_8335);
or U9082 (N_9082,N_8749,N_8585);
or U9083 (N_9083,N_8574,N_8217);
nor U9084 (N_9084,N_8801,N_8383);
nor U9085 (N_9085,N_8597,N_8668);
nor U9086 (N_9086,N_8268,N_8711);
and U9087 (N_9087,N_8602,N_8070);
or U9088 (N_9088,N_8556,N_8932);
nand U9089 (N_9089,N_8535,N_8003);
and U9090 (N_9090,N_8613,N_8944);
and U9091 (N_9091,N_8439,N_8767);
or U9092 (N_9092,N_8647,N_8223);
and U9093 (N_9093,N_8192,N_8067);
nor U9094 (N_9094,N_8392,N_8850);
or U9095 (N_9095,N_8821,N_8013);
nand U9096 (N_9096,N_8674,N_8935);
or U9097 (N_9097,N_8338,N_8074);
nor U9098 (N_9098,N_8607,N_8233);
and U9099 (N_9099,N_8404,N_8410);
or U9100 (N_9100,N_8549,N_8216);
nand U9101 (N_9101,N_8747,N_8555);
nand U9102 (N_9102,N_8194,N_8164);
nor U9103 (N_9103,N_8732,N_8389);
nor U9104 (N_9104,N_8805,N_8347);
or U9105 (N_9105,N_8433,N_8405);
and U9106 (N_9106,N_8921,N_8480);
nor U9107 (N_9107,N_8780,N_8111);
and U9108 (N_9108,N_8277,N_8280);
nor U9109 (N_9109,N_8447,N_8746);
or U9110 (N_9110,N_8979,N_8326);
or U9111 (N_9111,N_8726,N_8492);
and U9112 (N_9112,N_8987,N_8920);
and U9113 (N_9113,N_8459,N_8436);
nor U9114 (N_9114,N_8551,N_8796);
or U9115 (N_9115,N_8308,N_8472);
nand U9116 (N_9116,N_8735,N_8380);
nand U9117 (N_9117,N_8126,N_8393);
nand U9118 (N_9118,N_8106,N_8352);
or U9119 (N_9119,N_8970,N_8147);
nand U9120 (N_9120,N_8261,N_8521);
or U9121 (N_9121,N_8137,N_8428);
nor U9122 (N_9122,N_8143,N_8060);
and U9123 (N_9123,N_8744,N_8755);
nor U9124 (N_9124,N_8731,N_8622);
nand U9125 (N_9125,N_8019,N_8619);
nand U9126 (N_9126,N_8832,N_8058);
nor U9127 (N_9127,N_8643,N_8470);
or U9128 (N_9128,N_8697,N_8307);
nand U9129 (N_9129,N_8231,N_8376);
nor U9130 (N_9130,N_8375,N_8868);
nand U9131 (N_9131,N_8659,N_8134);
nand U9132 (N_9132,N_8294,N_8005);
nor U9133 (N_9133,N_8038,N_8128);
or U9134 (N_9134,N_8152,N_8188);
nor U9135 (N_9135,N_8080,N_8036);
nand U9136 (N_9136,N_8454,N_8896);
or U9137 (N_9137,N_8497,N_8491);
or U9138 (N_9138,N_8975,N_8642);
nor U9139 (N_9139,N_8639,N_8982);
and U9140 (N_9140,N_8600,N_8601);
nand U9141 (N_9141,N_8964,N_8566);
and U9142 (N_9142,N_8222,N_8709);
nand U9143 (N_9143,N_8197,N_8931);
and U9144 (N_9144,N_8438,N_8371);
nand U9145 (N_9145,N_8495,N_8630);
xnor U9146 (N_9146,N_8221,N_8026);
or U9147 (N_9147,N_8696,N_8089);
nor U9148 (N_9148,N_8278,N_8892);
or U9149 (N_9149,N_8373,N_8940);
nor U9150 (N_9150,N_8800,N_8101);
and U9151 (N_9151,N_8649,N_8690);
nor U9152 (N_9152,N_8968,N_8795);
or U9153 (N_9153,N_8394,N_8174);
nand U9154 (N_9154,N_8611,N_8916);
nand U9155 (N_9155,N_8758,N_8195);
nand U9156 (N_9156,N_8969,N_8900);
nor U9157 (N_9157,N_8183,N_8568);
nor U9158 (N_9158,N_8206,N_8385);
xnor U9159 (N_9159,N_8209,N_8750);
or U9160 (N_9160,N_8238,N_8006);
nand U9161 (N_9161,N_8440,N_8291);
nor U9162 (N_9162,N_8519,N_8977);
nor U9163 (N_9163,N_8071,N_8730);
nand U9164 (N_9164,N_8525,N_8055);
nand U9165 (N_9165,N_8880,N_8422);
nand U9166 (N_9166,N_8882,N_8235);
or U9167 (N_9167,N_8580,N_8604);
or U9168 (N_9168,N_8789,N_8023);
and U9169 (N_9169,N_8540,N_8243);
nand U9170 (N_9170,N_8378,N_8360);
nor U9171 (N_9171,N_8651,N_8837);
or U9172 (N_9172,N_8504,N_8906);
or U9173 (N_9173,N_8489,N_8565);
nand U9174 (N_9174,N_8486,N_8442);
nand U9175 (N_9175,N_8374,N_8324);
nand U9176 (N_9176,N_8445,N_8873);
nand U9177 (N_9177,N_8707,N_8908);
nor U9178 (N_9178,N_8173,N_8088);
nand U9179 (N_9179,N_8768,N_8985);
nand U9180 (N_9180,N_8869,N_8782);
nand U9181 (N_9181,N_8085,N_8009);
nor U9182 (N_9182,N_8548,N_8520);
or U9183 (N_9183,N_8358,N_8369);
and U9184 (N_9184,N_8725,N_8349);
and U9185 (N_9185,N_8362,N_8398);
and U9186 (N_9186,N_8939,N_8172);
nor U9187 (N_9187,N_8461,N_8002);
nor U9188 (N_9188,N_8765,N_8826);
nand U9189 (N_9189,N_8998,N_8049);
nor U9190 (N_9190,N_8984,N_8082);
nor U9191 (N_9191,N_8772,N_8363);
and U9192 (N_9192,N_8084,N_8992);
or U9193 (N_9193,N_8273,N_8384);
nand U9194 (N_9194,N_8550,N_8345);
nor U9195 (N_9195,N_8840,N_8287);
nor U9196 (N_9196,N_8511,N_8046);
or U9197 (N_9197,N_8564,N_8693);
or U9198 (N_9198,N_8553,N_8965);
nand U9199 (N_9199,N_8317,N_8420);
or U9200 (N_9200,N_8427,N_8458);
nand U9201 (N_9201,N_8861,N_8000);
nor U9202 (N_9202,N_8898,N_8591);
and U9203 (N_9203,N_8823,N_8501);
nand U9204 (N_9204,N_8295,N_8207);
nor U9205 (N_9205,N_8645,N_8952);
and U9206 (N_9206,N_8265,N_8419);
xor U9207 (N_9207,N_8914,N_8835);
and U9208 (N_9208,N_8579,N_8048);
or U9209 (N_9209,N_8211,N_8136);
or U9210 (N_9210,N_8703,N_8213);
or U9211 (N_9211,N_8925,N_8170);
nand U9212 (N_9212,N_8811,N_8103);
or U9213 (N_9213,N_8592,N_8652);
nor U9214 (N_9214,N_8350,N_8258);
or U9215 (N_9215,N_8215,N_8729);
and U9216 (N_9216,N_8839,N_8733);
nor U9217 (N_9217,N_8857,N_8853);
xor U9218 (N_9218,N_8605,N_8583);
or U9219 (N_9219,N_8682,N_8678);
or U9220 (N_9220,N_8762,N_8446);
nand U9221 (N_9221,N_8340,N_8575);
nor U9222 (N_9222,N_8704,N_8648);
nor U9223 (N_9223,N_8904,N_8842);
or U9224 (N_9224,N_8299,N_8059);
or U9225 (N_9225,N_8242,N_8791);
or U9226 (N_9226,N_8949,N_8547);
nand U9227 (N_9227,N_8889,N_8809);
nor U9228 (N_9228,N_8305,N_8999);
nand U9229 (N_9229,N_8098,N_8011);
or U9230 (N_9230,N_8056,N_8434);
nor U9231 (N_9231,N_8027,N_8836);
nand U9232 (N_9232,N_8596,N_8981);
nor U9233 (N_9233,N_8748,N_8593);
nor U9234 (N_9234,N_8015,N_8175);
or U9235 (N_9235,N_8165,N_8320);
or U9236 (N_9236,N_8962,N_8045);
and U9237 (N_9237,N_8692,N_8391);
and U9238 (N_9238,N_8166,N_8816);
and U9239 (N_9239,N_8849,N_8569);
and U9240 (N_9240,N_8301,N_8737);
or U9241 (N_9241,N_8246,N_8856);
and U9242 (N_9242,N_8494,N_8950);
or U9243 (N_9243,N_8064,N_8629);
nand U9244 (N_9244,N_8928,N_8270);
and U9245 (N_9245,N_8541,N_8264);
and U9246 (N_9246,N_8493,N_8160);
or U9247 (N_9247,N_8918,N_8657);
nand U9248 (N_9248,N_8879,N_8198);
nor U9249 (N_9249,N_8656,N_8050);
and U9250 (N_9250,N_8843,N_8512);
and U9251 (N_9251,N_8237,N_8081);
and U9252 (N_9252,N_8065,N_8411);
nand U9253 (N_9253,N_8191,N_8854);
and U9254 (N_9254,N_8584,N_8423);
or U9255 (N_9255,N_8974,N_8108);
nand U9256 (N_9256,N_8382,N_8488);
and U9257 (N_9257,N_8719,N_8431);
or U9258 (N_9258,N_8284,N_8676);
nor U9259 (N_9259,N_8039,N_8344);
or U9260 (N_9260,N_8911,N_8766);
nand U9261 (N_9261,N_8538,N_8205);
or U9262 (N_9262,N_8478,N_8151);
nor U9263 (N_9263,N_8888,N_8761);
or U9264 (N_9264,N_8379,N_8288);
and U9265 (N_9265,N_8956,N_8386);
or U9266 (N_9266,N_8496,N_8154);
xnor U9267 (N_9267,N_8255,N_8125);
xnor U9268 (N_9268,N_8533,N_8753);
or U9269 (N_9269,N_8210,N_8545);
nor U9270 (N_9270,N_8721,N_8763);
xor U9271 (N_9271,N_8989,N_8587);
nor U9272 (N_9272,N_8069,N_8670);
or U9273 (N_9273,N_8554,N_8655);
and U9274 (N_9274,N_8485,N_8367);
nand U9275 (N_9275,N_8150,N_8230);
and U9276 (N_9276,N_8713,N_8515);
or U9277 (N_9277,N_8966,N_8037);
and U9278 (N_9278,N_8714,N_8186);
or U9279 (N_9279,N_8897,N_8745);
nand U9280 (N_9280,N_8567,N_8572);
or U9281 (N_9281,N_8891,N_8783);
or U9282 (N_9282,N_8671,N_8285);
nand U9283 (N_9283,N_8021,N_8435);
or U9284 (N_9284,N_8503,N_8010);
nand U9285 (N_9285,N_8353,N_8068);
and U9286 (N_9286,N_8778,N_8129);
and U9287 (N_9287,N_8627,N_8922);
nand U9288 (N_9288,N_8862,N_8887);
nor U9289 (N_9289,N_8552,N_8421);
or U9290 (N_9290,N_8610,N_8603);
and U9291 (N_9291,N_8980,N_8316);
nor U9292 (N_9292,N_8119,N_8972);
xor U9293 (N_9293,N_8681,N_8444);
nor U9294 (N_9294,N_8414,N_8799);
nor U9295 (N_9295,N_8325,N_8516);
or U9296 (N_9296,N_8528,N_8586);
or U9297 (N_9297,N_8819,N_8181);
nor U9298 (N_9298,N_8001,N_8121);
nor U9299 (N_9299,N_8523,N_8787);
or U9300 (N_9300,N_8432,N_8115);
and U9301 (N_9301,N_8267,N_8754);
or U9302 (N_9302,N_8177,N_8881);
or U9303 (N_9303,N_8912,N_8322);
and U9304 (N_9304,N_8087,N_8334);
or U9305 (N_9305,N_8477,N_8524);
nand U9306 (N_9306,N_8760,N_8262);
or U9307 (N_9307,N_8229,N_8289);
xor U9308 (N_9308,N_8008,N_8626);
nor U9309 (N_9309,N_8044,N_8179);
nor U9310 (N_9310,N_8467,N_8667);
and U9311 (N_9311,N_8448,N_8282);
xor U9312 (N_9312,N_8661,N_8224);
and U9313 (N_9313,N_8594,N_8104);
nor U9314 (N_9314,N_8852,N_8012);
and U9315 (N_9315,N_8537,N_8323);
nand U9316 (N_9316,N_8025,N_8020);
nor U9317 (N_9317,N_8915,N_8573);
and U9318 (N_9318,N_8943,N_8752);
nor U9319 (N_9319,N_8412,N_8877);
nor U9320 (N_9320,N_8239,N_8792);
nor U9321 (N_9321,N_8946,N_8490);
and U9322 (N_9322,N_8319,N_8506);
nand U9323 (N_9323,N_8874,N_8140);
or U9324 (N_9324,N_8689,N_8751);
nor U9325 (N_9325,N_8091,N_8256);
nand U9326 (N_9326,N_8700,N_8919);
nor U9327 (N_9327,N_8634,N_8368);
nand U9328 (N_9328,N_8893,N_8558);
and U9329 (N_9329,N_8153,N_8960);
xor U9330 (N_9330,N_8543,N_8685);
and U9331 (N_9331,N_8644,N_8786);
nand U9332 (N_9332,N_8576,N_8953);
and U9333 (N_9333,N_8159,N_8844);
and U9334 (N_9334,N_8677,N_8640);
nand U9335 (N_9335,N_8321,N_8456);
or U9336 (N_9336,N_8252,N_8327);
or U9337 (N_9337,N_8757,N_8924);
nand U9338 (N_9338,N_8557,N_8475);
or U9339 (N_9339,N_8973,N_8526);
nor U9340 (N_9340,N_8364,N_8356);
and U9341 (N_9341,N_8859,N_8534);
xor U9342 (N_9342,N_8654,N_8077);
nor U9343 (N_9343,N_8986,N_8328);
nand U9344 (N_9344,N_8346,N_8304);
or U9345 (N_9345,N_8976,N_8958);
nor U9346 (N_9346,N_8544,N_8712);
nor U9347 (N_9347,N_8387,N_8846);
and U9348 (N_9348,N_8219,N_8114);
or U9349 (N_9349,N_8397,N_8571);
or U9350 (N_9350,N_8313,N_8281);
or U9351 (N_9351,N_8833,N_8738);
and U9352 (N_9352,N_8124,N_8468);
nand U9353 (N_9353,N_8260,N_8022);
or U9354 (N_9354,N_8417,N_8997);
nand U9355 (N_9355,N_8781,N_8532);
or U9356 (N_9356,N_8279,N_8708);
or U9357 (N_9357,N_8365,N_8451);
or U9358 (N_9358,N_8466,N_8635);
and U9359 (N_9359,N_8530,N_8079);
or U9360 (N_9360,N_8804,N_8109);
nand U9361 (N_9361,N_8618,N_8450);
nand U9362 (N_9362,N_8818,N_8830);
and U9363 (N_9363,N_8415,N_8033);
or U9364 (N_9364,N_8257,N_8190);
and U9365 (N_9365,N_8370,N_8163);
and U9366 (N_9366,N_8872,N_8465);
and U9367 (N_9367,N_8822,N_8196);
and U9368 (N_9368,N_8300,N_8658);
and U9369 (N_9369,N_8158,N_8971);
nand U9370 (N_9370,N_8110,N_8686);
and U9371 (N_9371,N_8679,N_8913);
nor U9372 (N_9372,N_8776,N_8810);
or U9373 (N_9373,N_8563,N_8863);
nand U9374 (N_9374,N_8135,N_8333);
nor U9375 (N_9375,N_8978,N_8028);
and U9376 (N_9376,N_8756,N_8820);
or U9377 (N_9377,N_8086,N_8815);
nor U9378 (N_9378,N_8131,N_8312);
nand U9379 (N_9379,N_8722,N_8169);
nor U9380 (N_9380,N_8988,N_8024);
or U9381 (N_9381,N_8959,N_8866);
xnor U9382 (N_9382,N_8043,N_8118);
xnor U9383 (N_9383,N_8259,N_8878);
nor U9384 (N_9384,N_8336,N_8471);
and U9385 (N_9385,N_8253,N_8306);
and U9386 (N_9386,N_8251,N_8199);
nor U9387 (N_9387,N_8561,N_8577);
nor U9388 (N_9388,N_8933,N_8066);
nand U9389 (N_9389,N_8775,N_8400);
nand U9390 (N_9390,N_8203,N_8041);
nand U9391 (N_9391,N_8684,N_8806);
and U9392 (N_9392,N_8354,N_8653);
xnor U9393 (N_9393,N_8884,N_8589);
or U9394 (N_9394,N_8636,N_8189);
nor U9395 (N_9395,N_8794,N_8588);
and U9396 (N_9396,N_8507,N_8204);
nand U9397 (N_9397,N_8691,N_8936);
nand U9398 (N_9398,N_8162,N_8263);
nand U9399 (N_9399,N_8269,N_8123);
nor U9400 (N_9400,N_8406,N_8734);
nand U9401 (N_9401,N_8286,N_8606);
and U9402 (N_9402,N_8314,N_8441);
nand U9403 (N_9403,N_8598,N_8141);
nor U9404 (N_9404,N_8146,N_8742);
nor U9405 (N_9405,N_8054,N_8145);
or U9406 (N_9406,N_8624,N_8185);
or U9407 (N_9407,N_8807,N_8035);
nand U9408 (N_9408,N_8680,N_8926);
and U9409 (N_9409,N_8075,N_8138);
nor U9410 (N_9410,N_8838,N_8225);
nor U9411 (N_9411,N_8894,N_8303);
nand U9412 (N_9412,N_8784,N_8860);
nor U9413 (N_9413,N_8117,N_8014);
and U9414 (N_9414,N_8127,N_8078);
xnor U9415 (N_9415,N_8774,N_8429);
or U9416 (N_9416,N_8723,N_8332);
nand U9417 (N_9417,N_8063,N_8883);
and U9418 (N_9418,N_8275,N_8923);
nand U9419 (N_9419,N_8500,N_8168);
nor U9420 (N_9420,N_8057,N_8740);
and U9421 (N_9421,N_8803,N_8247);
nand U9422 (N_9422,N_8156,N_8426);
or U9423 (N_9423,N_8076,N_8318);
nand U9424 (N_9424,N_8743,N_8462);
or U9425 (N_9425,N_8917,N_8902);
or U9426 (N_9426,N_8157,N_8248);
and U9427 (N_9427,N_8827,N_8581);
nor U9428 (N_9428,N_8250,N_8770);
nand U9429 (N_9429,N_8929,N_8570);
xor U9430 (N_9430,N_8798,N_8130);
and U9431 (N_9431,N_8113,N_8351);
or U9432 (N_9432,N_8413,N_8609);
nor U9433 (N_9433,N_8214,N_8372);
xor U9434 (N_9434,N_8608,N_8201);
nand U9435 (N_9435,N_8245,N_8073);
or U9436 (N_9436,N_8032,N_8452);
and U9437 (N_9437,N_8687,N_8266);
nand U9438 (N_9438,N_8895,N_8632);
nor U9439 (N_9439,N_8499,N_8773);
or U9440 (N_9440,N_8715,N_8560);
or U9441 (N_9441,N_8736,N_8825);
nor U9442 (N_9442,N_8107,N_8769);
nand U9443 (N_9443,N_8348,N_8483);
or U9444 (N_9444,N_8463,N_8227);
and U9445 (N_9445,N_8812,N_8460);
nand U9446 (N_9446,N_8249,N_8941);
and U9447 (N_9447,N_8942,N_8092);
nor U9448 (N_9448,N_8817,N_8717);
nand U9449 (N_9449,N_8623,N_8272);
xnor U9450 (N_9450,N_8072,N_8824);
or U9451 (N_9451,N_8672,N_8934);
or U9452 (N_9452,N_8673,N_8518);
nand U9453 (N_9453,N_8834,N_8228);
nand U9454 (N_9454,N_8476,N_8315);
or U9455 (N_9455,N_8662,N_8562);
nor U9456 (N_9456,N_8208,N_8716);
nand U9457 (N_9457,N_8663,N_8457);
and U9458 (N_9458,N_8200,N_8542);
or U9459 (N_9459,N_8509,N_8536);
and U9460 (N_9460,N_8042,N_8531);
nand U9461 (N_9461,N_8699,N_8234);
nor U9462 (N_9462,N_8990,N_8957);
nand U9463 (N_9463,N_8309,N_8047);
nor U9464 (N_9464,N_8425,N_8514);
nor U9465 (N_9465,N_8120,N_8954);
nor U9466 (N_9466,N_8705,N_8096);
or U9467 (N_9467,N_8927,N_8464);
nand U9468 (N_9468,N_8142,N_8017);
and U9469 (N_9469,N_8876,N_8144);
nor U9470 (N_9470,N_8139,N_8779);
xor U9471 (N_9471,N_8469,N_8337);
and U9472 (N_9472,N_8062,N_8155);
nor U9473 (N_9473,N_8617,N_8342);
nand U9474 (N_9474,N_8831,N_8399);
or U9475 (N_9475,N_8616,N_8790);
nand U9476 (N_9476,N_8967,N_8741);
nand U9477 (N_9477,N_8171,N_8983);
xor U9478 (N_9478,N_8938,N_8244);
or U9479 (N_9479,N_8910,N_8675);
and U9480 (N_9480,N_8122,N_8665);
or U9481 (N_9481,N_8283,N_8625);
nand U9482 (N_9482,N_8302,N_8582);
nand U9483 (N_9483,N_8329,N_8785);
nand U9484 (N_9484,N_8886,N_8095);
and U9485 (N_9485,N_8870,N_8409);
nor U9486 (N_9486,N_8218,N_8202);
nor U9487 (N_9487,N_8614,N_8034);
and U9488 (N_9488,N_8963,N_8875);
nand U9489 (N_9489,N_8310,N_8053);
xor U9490 (N_9490,N_8829,N_8706);
nor U9491 (N_9491,N_8061,N_8578);
or U9492 (N_9492,N_8178,N_8864);
or U9493 (N_9493,N_8093,N_8771);
nand U9494 (N_9494,N_8621,N_8443);
and U9495 (N_9495,N_8961,N_8841);
or U9496 (N_9496,N_8546,N_8311);
and U9497 (N_9497,N_8330,N_8633);
nor U9498 (N_9498,N_8187,N_8698);
nand U9499 (N_9499,N_8290,N_8727);
nor U9500 (N_9500,N_8153,N_8085);
or U9501 (N_9501,N_8043,N_8790);
or U9502 (N_9502,N_8657,N_8350);
or U9503 (N_9503,N_8887,N_8717);
or U9504 (N_9504,N_8518,N_8199);
and U9505 (N_9505,N_8967,N_8676);
nand U9506 (N_9506,N_8800,N_8535);
xor U9507 (N_9507,N_8006,N_8214);
and U9508 (N_9508,N_8518,N_8037);
nand U9509 (N_9509,N_8182,N_8532);
and U9510 (N_9510,N_8291,N_8520);
or U9511 (N_9511,N_8199,N_8885);
and U9512 (N_9512,N_8986,N_8176);
or U9513 (N_9513,N_8315,N_8413);
nand U9514 (N_9514,N_8669,N_8668);
nand U9515 (N_9515,N_8445,N_8137);
nor U9516 (N_9516,N_8677,N_8837);
or U9517 (N_9517,N_8815,N_8740);
nand U9518 (N_9518,N_8850,N_8070);
nand U9519 (N_9519,N_8016,N_8177);
nand U9520 (N_9520,N_8866,N_8558);
and U9521 (N_9521,N_8436,N_8198);
and U9522 (N_9522,N_8668,N_8418);
nor U9523 (N_9523,N_8994,N_8774);
nor U9524 (N_9524,N_8059,N_8581);
or U9525 (N_9525,N_8136,N_8720);
and U9526 (N_9526,N_8326,N_8516);
xnor U9527 (N_9527,N_8899,N_8141);
nor U9528 (N_9528,N_8438,N_8018);
or U9529 (N_9529,N_8860,N_8234);
and U9530 (N_9530,N_8100,N_8127);
nor U9531 (N_9531,N_8507,N_8552);
or U9532 (N_9532,N_8895,N_8189);
or U9533 (N_9533,N_8612,N_8454);
nor U9534 (N_9534,N_8618,N_8318);
and U9535 (N_9535,N_8916,N_8176);
or U9536 (N_9536,N_8208,N_8350);
nor U9537 (N_9537,N_8044,N_8355);
and U9538 (N_9538,N_8462,N_8303);
or U9539 (N_9539,N_8399,N_8312);
nor U9540 (N_9540,N_8746,N_8717);
nand U9541 (N_9541,N_8403,N_8596);
nor U9542 (N_9542,N_8522,N_8925);
and U9543 (N_9543,N_8368,N_8009);
nand U9544 (N_9544,N_8204,N_8889);
and U9545 (N_9545,N_8482,N_8002);
nand U9546 (N_9546,N_8117,N_8265);
or U9547 (N_9547,N_8475,N_8838);
nor U9548 (N_9548,N_8816,N_8574);
or U9549 (N_9549,N_8560,N_8514);
nor U9550 (N_9550,N_8930,N_8255);
nand U9551 (N_9551,N_8465,N_8123);
and U9552 (N_9552,N_8547,N_8666);
and U9553 (N_9553,N_8748,N_8502);
nor U9554 (N_9554,N_8935,N_8739);
and U9555 (N_9555,N_8640,N_8790);
nand U9556 (N_9556,N_8399,N_8045);
nand U9557 (N_9557,N_8821,N_8321);
nand U9558 (N_9558,N_8158,N_8841);
nand U9559 (N_9559,N_8999,N_8629);
and U9560 (N_9560,N_8197,N_8880);
nor U9561 (N_9561,N_8491,N_8121);
or U9562 (N_9562,N_8759,N_8225);
nand U9563 (N_9563,N_8677,N_8446);
or U9564 (N_9564,N_8054,N_8059);
or U9565 (N_9565,N_8735,N_8007);
or U9566 (N_9566,N_8149,N_8816);
nand U9567 (N_9567,N_8486,N_8168);
nand U9568 (N_9568,N_8862,N_8985);
nand U9569 (N_9569,N_8752,N_8634);
or U9570 (N_9570,N_8187,N_8437);
or U9571 (N_9571,N_8630,N_8646);
nor U9572 (N_9572,N_8711,N_8792);
or U9573 (N_9573,N_8438,N_8127);
and U9574 (N_9574,N_8072,N_8219);
nor U9575 (N_9575,N_8591,N_8996);
and U9576 (N_9576,N_8859,N_8502);
nand U9577 (N_9577,N_8708,N_8617);
xor U9578 (N_9578,N_8518,N_8364);
nor U9579 (N_9579,N_8754,N_8905);
or U9580 (N_9580,N_8272,N_8685);
nor U9581 (N_9581,N_8095,N_8638);
and U9582 (N_9582,N_8951,N_8779);
and U9583 (N_9583,N_8064,N_8335);
nand U9584 (N_9584,N_8486,N_8070);
and U9585 (N_9585,N_8685,N_8132);
nor U9586 (N_9586,N_8946,N_8264);
nor U9587 (N_9587,N_8544,N_8736);
and U9588 (N_9588,N_8281,N_8023);
and U9589 (N_9589,N_8748,N_8981);
nand U9590 (N_9590,N_8344,N_8963);
nand U9591 (N_9591,N_8826,N_8315);
nand U9592 (N_9592,N_8450,N_8355);
nor U9593 (N_9593,N_8218,N_8142);
nand U9594 (N_9594,N_8425,N_8393);
or U9595 (N_9595,N_8867,N_8616);
nand U9596 (N_9596,N_8290,N_8685);
nand U9597 (N_9597,N_8542,N_8403);
nand U9598 (N_9598,N_8602,N_8523);
and U9599 (N_9599,N_8742,N_8000);
or U9600 (N_9600,N_8109,N_8919);
nand U9601 (N_9601,N_8634,N_8719);
nand U9602 (N_9602,N_8034,N_8571);
nand U9603 (N_9603,N_8712,N_8886);
nand U9604 (N_9604,N_8016,N_8584);
nor U9605 (N_9605,N_8179,N_8555);
nand U9606 (N_9606,N_8747,N_8376);
nand U9607 (N_9607,N_8915,N_8484);
nor U9608 (N_9608,N_8634,N_8465);
and U9609 (N_9609,N_8167,N_8983);
nor U9610 (N_9610,N_8194,N_8844);
and U9611 (N_9611,N_8351,N_8216);
and U9612 (N_9612,N_8652,N_8886);
and U9613 (N_9613,N_8525,N_8719);
nor U9614 (N_9614,N_8152,N_8919);
nor U9615 (N_9615,N_8980,N_8199);
nand U9616 (N_9616,N_8092,N_8016);
nor U9617 (N_9617,N_8925,N_8744);
nand U9618 (N_9618,N_8024,N_8184);
and U9619 (N_9619,N_8926,N_8739);
or U9620 (N_9620,N_8573,N_8574);
and U9621 (N_9621,N_8411,N_8599);
or U9622 (N_9622,N_8928,N_8733);
nor U9623 (N_9623,N_8208,N_8475);
or U9624 (N_9624,N_8647,N_8032);
or U9625 (N_9625,N_8299,N_8100);
nand U9626 (N_9626,N_8775,N_8230);
nand U9627 (N_9627,N_8639,N_8316);
or U9628 (N_9628,N_8822,N_8040);
nor U9629 (N_9629,N_8434,N_8670);
nor U9630 (N_9630,N_8719,N_8334);
nand U9631 (N_9631,N_8370,N_8271);
and U9632 (N_9632,N_8588,N_8688);
nand U9633 (N_9633,N_8467,N_8452);
and U9634 (N_9634,N_8913,N_8663);
and U9635 (N_9635,N_8149,N_8586);
and U9636 (N_9636,N_8949,N_8182);
nor U9637 (N_9637,N_8848,N_8093);
nand U9638 (N_9638,N_8135,N_8707);
nand U9639 (N_9639,N_8568,N_8826);
nor U9640 (N_9640,N_8016,N_8961);
or U9641 (N_9641,N_8289,N_8767);
and U9642 (N_9642,N_8822,N_8682);
nand U9643 (N_9643,N_8248,N_8481);
nand U9644 (N_9644,N_8743,N_8242);
and U9645 (N_9645,N_8827,N_8057);
nor U9646 (N_9646,N_8480,N_8924);
nand U9647 (N_9647,N_8584,N_8633);
or U9648 (N_9648,N_8501,N_8170);
nor U9649 (N_9649,N_8163,N_8752);
nor U9650 (N_9650,N_8208,N_8773);
or U9651 (N_9651,N_8925,N_8516);
nand U9652 (N_9652,N_8831,N_8083);
xor U9653 (N_9653,N_8293,N_8289);
nand U9654 (N_9654,N_8964,N_8677);
and U9655 (N_9655,N_8677,N_8733);
and U9656 (N_9656,N_8255,N_8548);
nand U9657 (N_9657,N_8816,N_8514);
or U9658 (N_9658,N_8123,N_8291);
nand U9659 (N_9659,N_8371,N_8963);
or U9660 (N_9660,N_8916,N_8876);
nand U9661 (N_9661,N_8776,N_8223);
or U9662 (N_9662,N_8906,N_8389);
or U9663 (N_9663,N_8762,N_8295);
nand U9664 (N_9664,N_8268,N_8677);
or U9665 (N_9665,N_8509,N_8318);
or U9666 (N_9666,N_8117,N_8884);
and U9667 (N_9667,N_8992,N_8281);
or U9668 (N_9668,N_8241,N_8885);
nor U9669 (N_9669,N_8947,N_8046);
and U9670 (N_9670,N_8105,N_8810);
nor U9671 (N_9671,N_8563,N_8097);
xnor U9672 (N_9672,N_8427,N_8464);
xnor U9673 (N_9673,N_8614,N_8216);
nor U9674 (N_9674,N_8463,N_8206);
nand U9675 (N_9675,N_8334,N_8713);
nand U9676 (N_9676,N_8528,N_8494);
nand U9677 (N_9677,N_8777,N_8796);
nor U9678 (N_9678,N_8541,N_8297);
or U9679 (N_9679,N_8239,N_8307);
and U9680 (N_9680,N_8423,N_8530);
nor U9681 (N_9681,N_8506,N_8501);
or U9682 (N_9682,N_8026,N_8679);
nand U9683 (N_9683,N_8411,N_8372);
and U9684 (N_9684,N_8231,N_8624);
and U9685 (N_9685,N_8785,N_8624);
or U9686 (N_9686,N_8733,N_8565);
nor U9687 (N_9687,N_8609,N_8353);
and U9688 (N_9688,N_8714,N_8388);
nor U9689 (N_9689,N_8588,N_8797);
nor U9690 (N_9690,N_8878,N_8832);
or U9691 (N_9691,N_8392,N_8662);
nand U9692 (N_9692,N_8504,N_8657);
nor U9693 (N_9693,N_8077,N_8281);
nor U9694 (N_9694,N_8277,N_8456);
and U9695 (N_9695,N_8252,N_8790);
nor U9696 (N_9696,N_8200,N_8428);
or U9697 (N_9697,N_8692,N_8485);
nand U9698 (N_9698,N_8807,N_8513);
and U9699 (N_9699,N_8610,N_8235);
nor U9700 (N_9700,N_8386,N_8079);
nand U9701 (N_9701,N_8325,N_8588);
or U9702 (N_9702,N_8528,N_8705);
and U9703 (N_9703,N_8576,N_8527);
or U9704 (N_9704,N_8569,N_8713);
nor U9705 (N_9705,N_8791,N_8275);
or U9706 (N_9706,N_8191,N_8375);
or U9707 (N_9707,N_8245,N_8583);
or U9708 (N_9708,N_8707,N_8627);
or U9709 (N_9709,N_8445,N_8018);
or U9710 (N_9710,N_8726,N_8796);
nor U9711 (N_9711,N_8652,N_8849);
or U9712 (N_9712,N_8466,N_8320);
nand U9713 (N_9713,N_8315,N_8211);
nor U9714 (N_9714,N_8721,N_8117);
nand U9715 (N_9715,N_8835,N_8175);
nand U9716 (N_9716,N_8757,N_8190);
and U9717 (N_9717,N_8594,N_8959);
nor U9718 (N_9718,N_8022,N_8822);
nand U9719 (N_9719,N_8517,N_8856);
or U9720 (N_9720,N_8855,N_8381);
nor U9721 (N_9721,N_8960,N_8753);
nor U9722 (N_9722,N_8574,N_8534);
and U9723 (N_9723,N_8246,N_8853);
nor U9724 (N_9724,N_8873,N_8219);
or U9725 (N_9725,N_8100,N_8141);
or U9726 (N_9726,N_8909,N_8953);
nand U9727 (N_9727,N_8664,N_8773);
nand U9728 (N_9728,N_8684,N_8950);
nand U9729 (N_9729,N_8369,N_8440);
or U9730 (N_9730,N_8676,N_8105);
or U9731 (N_9731,N_8969,N_8718);
nor U9732 (N_9732,N_8955,N_8845);
or U9733 (N_9733,N_8372,N_8524);
nor U9734 (N_9734,N_8531,N_8134);
nand U9735 (N_9735,N_8740,N_8312);
nand U9736 (N_9736,N_8891,N_8610);
or U9737 (N_9737,N_8283,N_8589);
nand U9738 (N_9738,N_8529,N_8353);
nor U9739 (N_9739,N_8129,N_8761);
and U9740 (N_9740,N_8999,N_8464);
or U9741 (N_9741,N_8539,N_8088);
or U9742 (N_9742,N_8247,N_8889);
nand U9743 (N_9743,N_8503,N_8682);
or U9744 (N_9744,N_8626,N_8110);
nand U9745 (N_9745,N_8913,N_8733);
or U9746 (N_9746,N_8402,N_8176);
nand U9747 (N_9747,N_8892,N_8380);
and U9748 (N_9748,N_8976,N_8591);
nand U9749 (N_9749,N_8686,N_8218);
or U9750 (N_9750,N_8612,N_8208);
xnor U9751 (N_9751,N_8503,N_8006);
nand U9752 (N_9752,N_8692,N_8908);
nand U9753 (N_9753,N_8262,N_8198);
nor U9754 (N_9754,N_8124,N_8001);
nor U9755 (N_9755,N_8568,N_8134);
and U9756 (N_9756,N_8854,N_8751);
nor U9757 (N_9757,N_8420,N_8081);
nand U9758 (N_9758,N_8163,N_8230);
nor U9759 (N_9759,N_8538,N_8931);
nand U9760 (N_9760,N_8941,N_8623);
and U9761 (N_9761,N_8150,N_8295);
nand U9762 (N_9762,N_8364,N_8922);
nand U9763 (N_9763,N_8410,N_8536);
or U9764 (N_9764,N_8932,N_8050);
and U9765 (N_9765,N_8692,N_8801);
nor U9766 (N_9766,N_8261,N_8288);
nor U9767 (N_9767,N_8642,N_8202);
nor U9768 (N_9768,N_8901,N_8208);
nor U9769 (N_9769,N_8968,N_8356);
nand U9770 (N_9770,N_8864,N_8049);
nor U9771 (N_9771,N_8935,N_8830);
xor U9772 (N_9772,N_8956,N_8309);
or U9773 (N_9773,N_8672,N_8152);
nand U9774 (N_9774,N_8603,N_8711);
or U9775 (N_9775,N_8222,N_8588);
or U9776 (N_9776,N_8028,N_8318);
or U9777 (N_9777,N_8302,N_8523);
nand U9778 (N_9778,N_8447,N_8170);
and U9779 (N_9779,N_8535,N_8338);
nand U9780 (N_9780,N_8726,N_8246);
and U9781 (N_9781,N_8607,N_8642);
and U9782 (N_9782,N_8540,N_8405);
xor U9783 (N_9783,N_8507,N_8087);
nand U9784 (N_9784,N_8984,N_8193);
nor U9785 (N_9785,N_8367,N_8658);
nand U9786 (N_9786,N_8913,N_8446);
and U9787 (N_9787,N_8445,N_8945);
nor U9788 (N_9788,N_8475,N_8860);
or U9789 (N_9789,N_8140,N_8813);
or U9790 (N_9790,N_8530,N_8025);
or U9791 (N_9791,N_8180,N_8190);
nand U9792 (N_9792,N_8150,N_8028);
nand U9793 (N_9793,N_8058,N_8143);
and U9794 (N_9794,N_8236,N_8370);
or U9795 (N_9795,N_8335,N_8621);
and U9796 (N_9796,N_8766,N_8448);
and U9797 (N_9797,N_8169,N_8778);
nor U9798 (N_9798,N_8557,N_8602);
or U9799 (N_9799,N_8956,N_8172);
or U9800 (N_9800,N_8440,N_8277);
nor U9801 (N_9801,N_8775,N_8385);
and U9802 (N_9802,N_8766,N_8412);
nor U9803 (N_9803,N_8498,N_8962);
nand U9804 (N_9804,N_8804,N_8986);
nor U9805 (N_9805,N_8322,N_8248);
xnor U9806 (N_9806,N_8380,N_8647);
and U9807 (N_9807,N_8496,N_8456);
nor U9808 (N_9808,N_8224,N_8080);
or U9809 (N_9809,N_8736,N_8328);
or U9810 (N_9810,N_8193,N_8211);
or U9811 (N_9811,N_8038,N_8814);
nand U9812 (N_9812,N_8167,N_8407);
nand U9813 (N_9813,N_8347,N_8947);
and U9814 (N_9814,N_8239,N_8544);
and U9815 (N_9815,N_8123,N_8826);
or U9816 (N_9816,N_8990,N_8566);
or U9817 (N_9817,N_8994,N_8470);
nor U9818 (N_9818,N_8736,N_8822);
or U9819 (N_9819,N_8521,N_8468);
and U9820 (N_9820,N_8357,N_8900);
and U9821 (N_9821,N_8537,N_8207);
or U9822 (N_9822,N_8079,N_8347);
nor U9823 (N_9823,N_8868,N_8072);
and U9824 (N_9824,N_8947,N_8736);
or U9825 (N_9825,N_8650,N_8936);
nor U9826 (N_9826,N_8153,N_8517);
and U9827 (N_9827,N_8575,N_8093);
nor U9828 (N_9828,N_8169,N_8319);
and U9829 (N_9829,N_8133,N_8063);
nor U9830 (N_9830,N_8555,N_8775);
nand U9831 (N_9831,N_8438,N_8313);
or U9832 (N_9832,N_8376,N_8698);
or U9833 (N_9833,N_8496,N_8165);
or U9834 (N_9834,N_8307,N_8149);
and U9835 (N_9835,N_8197,N_8894);
nand U9836 (N_9836,N_8933,N_8931);
or U9837 (N_9837,N_8624,N_8675);
and U9838 (N_9838,N_8845,N_8462);
nor U9839 (N_9839,N_8672,N_8254);
and U9840 (N_9840,N_8561,N_8430);
nand U9841 (N_9841,N_8677,N_8364);
nand U9842 (N_9842,N_8456,N_8898);
nor U9843 (N_9843,N_8074,N_8867);
or U9844 (N_9844,N_8090,N_8496);
or U9845 (N_9845,N_8622,N_8514);
and U9846 (N_9846,N_8030,N_8324);
nand U9847 (N_9847,N_8095,N_8250);
or U9848 (N_9848,N_8614,N_8217);
nor U9849 (N_9849,N_8440,N_8573);
and U9850 (N_9850,N_8098,N_8018);
or U9851 (N_9851,N_8608,N_8158);
or U9852 (N_9852,N_8038,N_8921);
nand U9853 (N_9853,N_8977,N_8940);
and U9854 (N_9854,N_8198,N_8777);
or U9855 (N_9855,N_8108,N_8091);
nor U9856 (N_9856,N_8822,N_8429);
and U9857 (N_9857,N_8058,N_8648);
nor U9858 (N_9858,N_8334,N_8738);
nand U9859 (N_9859,N_8002,N_8208);
nor U9860 (N_9860,N_8640,N_8920);
and U9861 (N_9861,N_8792,N_8503);
or U9862 (N_9862,N_8696,N_8929);
and U9863 (N_9863,N_8408,N_8304);
and U9864 (N_9864,N_8643,N_8625);
and U9865 (N_9865,N_8326,N_8588);
or U9866 (N_9866,N_8703,N_8055);
nor U9867 (N_9867,N_8695,N_8865);
or U9868 (N_9868,N_8015,N_8655);
and U9869 (N_9869,N_8493,N_8709);
and U9870 (N_9870,N_8904,N_8367);
nand U9871 (N_9871,N_8706,N_8392);
nand U9872 (N_9872,N_8550,N_8412);
nand U9873 (N_9873,N_8596,N_8801);
or U9874 (N_9874,N_8724,N_8958);
nand U9875 (N_9875,N_8077,N_8832);
nor U9876 (N_9876,N_8582,N_8711);
and U9877 (N_9877,N_8978,N_8137);
or U9878 (N_9878,N_8537,N_8278);
and U9879 (N_9879,N_8036,N_8902);
nor U9880 (N_9880,N_8028,N_8086);
and U9881 (N_9881,N_8041,N_8194);
nor U9882 (N_9882,N_8952,N_8600);
nor U9883 (N_9883,N_8006,N_8406);
and U9884 (N_9884,N_8704,N_8596);
or U9885 (N_9885,N_8343,N_8731);
nor U9886 (N_9886,N_8847,N_8785);
and U9887 (N_9887,N_8024,N_8180);
and U9888 (N_9888,N_8745,N_8207);
nor U9889 (N_9889,N_8345,N_8491);
nor U9890 (N_9890,N_8019,N_8668);
nand U9891 (N_9891,N_8582,N_8976);
or U9892 (N_9892,N_8368,N_8848);
nor U9893 (N_9893,N_8233,N_8187);
nor U9894 (N_9894,N_8465,N_8247);
nor U9895 (N_9895,N_8504,N_8170);
and U9896 (N_9896,N_8942,N_8833);
nand U9897 (N_9897,N_8481,N_8225);
or U9898 (N_9898,N_8557,N_8626);
nand U9899 (N_9899,N_8722,N_8314);
nor U9900 (N_9900,N_8667,N_8147);
or U9901 (N_9901,N_8438,N_8584);
and U9902 (N_9902,N_8513,N_8738);
or U9903 (N_9903,N_8142,N_8257);
nor U9904 (N_9904,N_8825,N_8007);
xnor U9905 (N_9905,N_8716,N_8595);
nor U9906 (N_9906,N_8061,N_8863);
and U9907 (N_9907,N_8355,N_8593);
nand U9908 (N_9908,N_8082,N_8685);
nor U9909 (N_9909,N_8033,N_8598);
or U9910 (N_9910,N_8740,N_8692);
or U9911 (N_9911,N_8861,N_8953);
nand U9912 (N_9912,N_8698,N_8070);
or U9913 (N_9913,N_8728,N_8010);
or U9914 (N_9914,N_8818,N_8367);
and U9915 (N_9915,N_8000,N_8817);
or U9916 (N_9916,N_8270,N_8723);
and U9917 (N_9917,N_8471,N_8582);
and U9918 (N_9918,N_8042,N_8357);
nand U9919 (N_9919,N_8277,N_8621);
nor U9920 (N_9920,N_8872,N_8819);
xnor U9921 (N_9921,N_8824,N_8606);
nand U9922 (N_9922,N_8883,N_8738);
nand U9923 (N_9923,N_8443,N_8023);
or U9924 (N_9924,N_8031,N_8345);
and U9925 (N_9925,N_8553,N_8412);
nand U9926 (N_9926,N_8978,N_8098);
or U9927 (N_9927,N_8451,N_8734);
and U9928 (N_9928,N_8306,N_8568);
or U9929 (N_9929,N_8484,N_8308);
nand U9930 (N_9930,N_8776,N_8807);
and U9931 (N_9931,N_8187,N_8724);
nor U9932 (N_9932,N_8612,N_8277);
and U9933 (N_9933,N_8852,N_8179);
nand U9934 (N_9934,N_8128,N_8363);
nor U9935 (N_9935,N_8379,N_8329);
or U9936 (N_9936,N_8237,N_8402);
or U9937 (N_9937,N_8318,N_8264);
nor U9938 (N_9938,N_8125,N_8718);
nor U9939 (N_9939,N_8867,N_8487);
and U9940 (N_9940,N_8184,N_8310);
nand U9941 (N_9941,N_8216,N_8035);
nor U9942 (N_9942,N_8513,N_8439);
or U9943 (N_9943,N_8341,N_8972);
xor U9944 (N_9944,N_8179,N_8939);
or U9945 (N_9945,N_8155,N_8402);
or U9946 (N_9946,N_8857,N_8788);
and U9947 (N_9947,N_8452,N_8403);
nand U9948 (N_9948,N_8330,N_8870);
nand U9949 (N_9949,N_8720,N_8548);
or U9950 (N_9950,N_8209,N_8108);
and U9951 (N_9951,N_8881,N_8612);
and U9952 (N_9952,N_8041,N_8413);
or U9953 (N_9953,N_8373,N_8410);
or U9954 (N_9954,N_8520,N_8076);
and U9955 (N_9955,N_8882,N_8241);
or U9956 (N_9956,N_8939,N_8987);
nand U9957 (N_9957,N_8208,N_8699);
nand U9958 (N_9958,N_8288,N_8052);
nor U9959 (N_9959,N_8662,N_8256);
and U9960 (N_9960,N_8282,N_8663);
nand U9961 (N_9961,N_8854,N_8661);
nand U9962 (N_9962,N_8617,N_8058);
nand U9963 (N_9963,N_8992,N_8922);
and U9964 (N_9964,N_8987,N_8146);
nand U9965 (N_9965,N_8158,N_8357);
nor U9966 (N_9966,N_8052,N_8570);
nand U9967 (N_9967,N_8273,N_8387);
and U9968 (N_9968,N_8325,N_8075);
or U9969 (N_9969,N_8083,N_8714);
and U9970 (N_9970,N_8723,N_8527);
nor U9971 (N_9971,N_8829,N_8541);
or U9972 (N_9972,N_8140,N_8223);
or U9973 (N_9973,N_8257,N_8963);
and U9974 (N_9974,N_8781,N_8616);
nor U9975 (N_9975,N_8368,N_8044);
or U9976 (N_9976,N_8407,N_8110);
and U9977 (N_9977,N_8948,N_8708);
and U9978 (N_9978,N_8276,N_8476);
nor U9979 (N_9979,N_8672,N_8892);
and U9980 (N_9980,N_8110,N_8475);
nor U9981 (N_9981,N_8167,N_8426);
and U9982 (N_9982,N_8033,N_8278);
and U9983 (N_9983,N_8129,N_8681);
or U9984 (N_9984,N_8898,N_8515);
or U9985 (N_9985,N_8337,N_8141);
nand U9986 (N_9986,N_8908,N_8558);
or U9987 (N_9987,N_8377,N_8769);
and U9988 (N_9988,N_8804,N_8405);
nand U9989 (N_9989,N_8463,N_8074);
nand U9990 (N_9990,N_8708,N_8997);
and U9991 (N_9991,N_8551,N_8852);
nor U9992 (N_9992,N_8564,N_8316);
or U9993 (N_9993,N_8579,N_8059);
and U9994 (N_9994,N_8779,N_8399);
nand U9995 (N_9995,N_8087,N_8564);
nand U9996 (N_9996,N_8201,N_8896);
or U9997 (N_9997,N_8918,N_8695);
and U9998 (N_9998,N_8844,N_8677);
or U9999 (N_9999,N_8305,N_8795);
or UO_0 (O_0,N_9191,N_9701);
nand UO_1 (O_1,N_9034,N_9427);
or UO_2 (O_2,N_9370,N_9496);
and UO_3 (O_3,N_9605,N_9838);
nand UO_4 (O_4,N_9021,N_9631);
and UO_5 (O_5,N_9644,N_9065);
nand UO_6 (O_6,N_9033,N_9176);
nand UO_7 (O_7,N_9294,N_9092);
and UO_8 (O_8,N_9352,N_9994);
nand UO_9 (O_9,N_9369,N_9190);
or UO_10 (O_10,N_9666,N_9948);
and UO_11 (O_11,N_9878,N_9936);
and UO_12 (O_12,N_9080,N_9226);
nand UO_13 (O_13,N_9035,N_9603);
or UO_14 (O_14,N_9965,N_9517);
nand UO_15 (O_15,N_9562,N_9625);
nand UO_16 (O_16,N_9251,N_9183);
and UO_17 (O_17,N_9101,N_9070);
and UO_18 (O_18,N_9103,N_9995);
nand UO_19 (O_19,N_9503,N_9127);
nor UO_20 (O_20,N_9683,N_9163);
or UO_21 (O_21,N_9632,N_9102);
nor UO_22 (O_22,N_9753,N_9032);
or UO_23 (O_23,N_9794,N_9716);
nor UO_24 (O_24,N_9312,N_9570);
nand UO_25 (O_25,N_9292,N_9615);
or UO_26 (O_26,N_9260,N_9330);
nor UO_27 (O_27,N_9720,N_9690);
or UO_28 (O_28,N_9182,N_9610);
or UO_29 (O_29,N_9271,N_9469);
or UO_30 (O_30,N_9588,N_9111);
and UO_31 (O_31,N_9449,N_9923);
and UO_32 (O_32,N_9265,N_9998);
nand UO_33 (O_33,N_9803,N_9952);
and UO_34 (O_34,N_9184,N_9314);
nand UO_35 (O_35,N_9808,N_9036);
nand UO_36 (O_36,N_9408,N_9212);
and UO_37 (O_37,N_9456,N_9406);
and UO_38 (O_38,N_9595,N_9253);
nand UO_39 (O_39,N_9795,N_9098);
and UO_40 (O_40,N_9419,N_9366);
nor UO_41 (O_41,N_9889,N_9596);
nand UO_42 (O_42,N_9641,N_9692);
and UO_43 (O_43,N_9852,N_9219);
nor UO_44 (O_44,N_9992,N_9295);
nand UO_45 (O_45,N_9160,N_9914);
or UO_46 (O_46,N_9071,N_9122);
nor UO_47 (O_47,N_9417,N_9428);
nor UO_48 (O_48,N_9360,N_9131);
or UO_49 (O_49,N_9583,N_9050);
and UO_50 (O_50,N_9693,N_9713);
and UO_51 (O_51,N_9470,N_9984);
or UO_52 (O_52,N_9083,N_9677);
and UO_53 (O_53,N_9565,N_9578);
nand UO_54 (O_54,N_9442,N_9281);
nand UO_55 (O_55,N_9947,N_9572);
nand UO_56 (O_56,N_9571,N_9133);
xnor UO_57 (O_57,N_9434,N_9349);
or UO_58 (O_58,N_9240,N_9973);
and UO_59 (O_59,N_9095,N_9254);
or UO_60 (O_60,N_9397,N_9563);
or UO_61 (O_61,N_9079,N_9384);
and UO_62 (O_62,N_9877,N_9961);
and UO_63 (O_63,N_9532,N_9574);
or UO_64 (O_64,N_9773,N_9308);
nor UO_65 (O_65,N_9680,N_9958);
or UO_66 (O_66,N_9120,N_9669);
and UO_67 (O_67,N_9144,N_9275);
nand UO_68 (O_68,N_9403,N_9657);
and UO_69 (O_69,N_9484,N_9388);
nand UO_70 (O_70,N_9185,N_9293);
nor UO_71 (O_71,N_9582,N_9402);
nor UO_72 (O_72,N_9202,N_9862);
and UO_73 (O_73,N_9387,N_9904);
nand UO_74 (O_74,N_9223,N_9609);
and UO_75 (O_75,N_9674,N_9554);
nor UO_76 (O_76,N_9522,N_9157);
xnor UO_77 (O_77,N_9300,N_9941);
nor UO_78 (O_78,N_9161,N_9651);
and UO_79 (O_79,N_9526,N_9474);
nor UO_80 (O_80,N_9166,N_9718);
nor UO_81 (O_81,N_9617,N_9247);
or UO_82 (O_82,N_9301,N_9780);
or UO_83 (O_83,N_9118,N_9316);
nor UO_84 (O_84,N_9946,N_9222);
or UO_85 (O_85,N_9749,N_9857);
nor UO_86 (O_86,N_9933,N_9438);
or UO_87 (O_87,N_9029,N_9497);
nor UO_88 (O_88,N_9062,N_9956);
xor UO_89 (O_89,N_9466,N_9949);
and UO_90 (O_90,N_9139,N_9900);
or UO_91 (O_91,N_9709,N_9685);
nor UO_92 (O_92,N_9146,N_9698);
nor UO_93 (O_93,N_9473,N_9898);
nor UO_94 (O_94,N_9269,N_9988);
nand UO_95 (O_95,N_9348,N_9210);
nor UO_96 (O_96,N_9879,N_9054);
and UO_97 (O_97,N_9648,N_9010);
and UO_98 (O_98,N_9766,N_9723);
nor UO_99 (O_99,N_9228,N_9204);
nand UO_100 (O_100,N_9699,N_9924);
nor UO_101 (O_101,N_9359,N_9209);
and UO_102 (O_102,N_9052,N_9856);
or UO_103 (O_103,N_9962,N_9302);
and UO_104 (O_104,N_9180,N_9845);
or UO_105 (O_105,N_9041,N_9687);
xnor UO_106 (O_106,N_9665,N_9194);
and UO_107 (O_107,N_9884,N_9654);
nor UO_108 (O_108,N_9091,N_9076);
nor UO_109 (O_109,N_9827,N_9934);
or UO_110 (O_110,N_9471,N_9192);
or UO_111 (O_111,N_9058,N_9530);
nor UO_112 (O_112,N_9660,N_9072);
or UO_113 (O_113,N_9886,N_9964);
and UO_114 (O_114,N_9016,N_9206);
or UO_115 (O_115,N_9493,N_9407);
nor UO_116 (O_116,N_9842,N_9587);
and UO_117 (O_117,N_9391,N_9805);
nand UO_118 (O_118,N_9444,N_9601);
nor UO_119 (O_119,N_9918,N_9899);
nor UO_120 (O_120,N_9511,N_9024);
and UO_121 (O_121,N_9216,N_9800);
and UO_122 (O_122,N_9325,N_9756);
nand UO_123 (O_123,N_9013,N_9682);
nor UO_124 (O_124,N_9329,N_9611);
nand UO_125 (O_125,N_9145,N_9979);
or UO_126 (O_126,N_9436,N_9358);
nand UO_127 (O_127,N_9480,N_9980);
nor UO_128 (O_128,N_9376,N_9170);
and UO_129 (O_129,N_9327,N_9414);
nor UO_130 (O_130,N_9761,N_9671);
and UO_131 (O_131,N_9439,N_9015);
nor UO_132 (O_132,N_9785,N_9652);
nand UO_133 (O_133,N_9782,N_9108);
nor UO_134 (O_134,N_9106,N_9575);
or UO_135 (O_135,N_9126,N_9999);
and UO_136 (O_136,N_9321,N_9598);
nand UO_137 (O_137,N_9492,N_9765);
nor UO_138 (O_138,N_9132,N_9375);
or UO_139 (O_139,N_9819,N_9241);
nor UO_140 (O_140,N_9549,N_9435);
nand UO_141 (O_141,N_9513,N_9931);
nor UO_142 (O_142,N_9121,N_9337);
or UO_143 (O_143,N_9688,N_9515);
nor UO_144 (O_144,N_9287,N_9479);
nor UO_145 (O_145,N_9861,N_9940);
and UO_146 (O_146,N_9916,N_9172);
and UO_147 (O_147,N_9786,N_9211);
or UO_148 (O_148,N_9335,N_9848);
xnor UO_149 (O_149,N_9084,N_9535);
nor UO_150 (O_150,N_9813,N_9158);
nor UO_151 (O_151,N_9623,N_9594);
or UO_152 (O_152,N_9303,N_9835);
or UO_153 (O_153,N_9987,N_9356);
and UO_154 (O_154,N_9930,N_9451);
and UO_155 (O_155,N_9364,N_9097);
nand UO_156 (O_156,N_9905,N_9985);
nand UO_157 (O_157,N_9396,N_9638);
and UO_158 (O_158,N_9664,N_9087);
and UO_159 (O_159,N_9890,N_9917);
and UO_160 (O_160,N_9876,N_9558);
and UO_161 (O_161,N_9841,N_9981);
nor UO_162 (O_162,N_9307,N_9067);
or UO_163 (O_163,N_9804,N_9656);
and UO_164 (O_164,N_9536,N_9353);
and UO_165 (O_165,N_9873,N_9854);
nor UO_166 (O_166,N_9839,N_9745);
or UO_167 (O_167,N_9799,N_9051);
nor UO_168 (O_168,N_9510,N_9775);
nor UO_169 (O_169,N_9802,N_9430);
or UO_170 (O_170,N_9239,N_9467);
nor UO_171 (O_171,N_9735,N_9201);
nand UO_172 (O_172,N_9672,N_9538);
nand UO_173 (O_173,N_9568,N_9566);
nor UO_174 (O_174,N_9268,N_9663);
nand UO_175 (O_175,N_9093,N_9494);
nor UO_176 (O_176,N_9231,N_9728);
or UO_177 (O_177,N_9791,N_9009);
or UO_178 (O_178,N_9870,N_9772);
nand UO_179 (O_179,N_9897,N_9249);
nor UO_180 (O_180,N_9319,N_9027);
nor UO_181 (O_181,N_9825,N_9342);
nand UO_182 (O_182,N_9367,N_9730);
nand UO_183 (O_183,N_9806,N_9282);
or UO_184 (O_184,N_9628,N_9077);
nor UO_185 (O_185,N_9746,N_9218);
and UO_186 (O_186,N_9278,N_9291);
xnor UO_187 (O_187,N_9913,N_9908);
and UO_188 (O_188,N_9432,N_9846);
nand UO_189 (O_189,N_9661,N_9590);
nand UO_190 (O_190,N_9708,N_9831);
nor UO_191 (O_191,N_9602,N_9004);
nand UO_192 (O_192,N_9450,N_9844);
nand UO_193 (O_193,N_9372,N_9483);
nand UO_194 (O_194,N_9863,N_9382);
nor UO_195 (O_195,N_9090,N_9237);
or UO_196 (O_196,N_9039,N_9548);
nand UO_197 (O_197,N_9637,N_9017);
or UO_198 (O_198,N_9885,N_9107);
or UO_199 (O_199,N_9750,N_9350);
nand UO_200 (O_200,N_9042,N_9893);
and UO_201 (O_201,N_9954,N_9619);
nand UO_202 (O_202,N_9950,N_9109);
nor UO_203 (O_203,N_9686,N_9203);
and UO_204 (O_204,N_9576,N_9362);
nand UO_205 (O_205,N_9630,N_9116);
nor UO_206 (O_206,N_9714,N_9264);
nor UO_207 (O_207,N_9640,N_9970);
or UO_208 (O_208,N_9986,N_9380);
nand UO_209 (O_209,N_9817,N_9412);
or UO_210 (O_210,N_9585,N_9464);
nor UO_211 (O_211,N_9213,N_9901);
nor UO_212 (O_212,N_9943,N_9816);
and UO_213 (O_213,N_9922,N_9604);
or UO_214 (O_214,N_9023,N_9200);
and UO_215 (O_215,N_9164,N_9512);
or UO_216 (O_216,N_9853,N_9082);
nor UO_217 (O_217,N_9233,N_9919);
nand UO_218 (O_218,N_9821,N_9323);
or UO_219 (O_219,N_9612,N_9500);
nor UO_220 (O_220,N_9289,N_9215);
nor UO_221 (O_221,N_9276,N_9855);
xnor UO_222 (O_222,N_9894,N_9724);
or UO_223 (O_223,N_9059,N_9755);
xor UO_224 (O_224,N_9525,N_9710);
and UO_225 (O_225,N_9220,N_9426);
nor UO_226 (O_226,N_9818,N_9485);
and UO_227 (O_227,N_9341,N_9501);
nand UO_228 (O_228,N_9207,N_9658);
or UO_229 (O_229,N_9338,N_9151);
and UO_230 (O_230,N_9232,N_9543);
nor UO_231 (O_231,N_9504,N_9860);
nand UO_232 (O_232,N_9912,N_9198);
or UO_233 (O_233,N_9704,N_9368);
and UO_234 (O_234,N_9993,N_9395);
nand UO_235 (O_235,N_9085,N_9398);
or UO_236 (O_236,N_9977,N_9060);
nor UO_237 (O_237,N_9836,N_9519);
or UO_238 (O_238,N_9553,N_9586);
or UO_239 (O_239,N_9221,N_9138);
or UO_240 (O_240,N_9920,N_9463);
and UO_241 (O_241,N_9381,N_9425);
and UO_242 (O_242,N_9357,N_9458);
nand UO_243 (O_243,N_9557,N_9673);
nand UO_244 (O_244,N_9874,N_9064);
and UO_245 (O_245,N_9932,N_9618);
nand UO_246 (O_246,N_9047,N_9270);
or UO_247 (O_247,N_9489,N_9326);
nand UO_248 (O_248,N_9925,N_9740);
and UO_249 (O_249,N_9162,N_9697);
and UO_250 (O_250,N_9778,N_9331);
nor UO_251 (O_251,N_9787,N_9696);
nand UO_252 (O_252,N_9334,N_9681);
or UO_253 (O_253,N_9404,N_9354);
nor UO_254 (O_254,N_9320,N_9476);
and UO_255 (O_255,N_9005,N_9142);
nor UO_256 (O_256,N_9472,N_9869);
nand UO_257 (O_257,N_9227,N_9297);
nand UO_258 (O_258,N_9647,N_9482);
and UO_259 (O_259,N_9872,N_9643);
and UO_260 (O_260,N_9929,N_9187);
nand UO_261 (O_261,N_9012,N_9189);
nand UO_262 (O_262,N_9502,N_9002);
and UO_263 (O_263,N_9383,N_9056);
nand UO_264 (O_264,N_9678,N_9174);
nor UO_265 (O_265,N_9305,N_9840);
and UO_266 (O_266,N_9847,N_9823);
and UO_267 (O_267,N_9256,N_9437);
and UO_268 (O_268,N_9006,N_9891);
nand UO_269 (O_269,N_9117,N_9655);
nand UO_270 (O_270,N_9234,N_9545);
nand UO_271 (O_271,N_9712,N_9089);
xnor UO_272 (O_272,N_9737,N_9812);
and UO_273 (O_273,N_9937,N_9754);
nand UO_274 (O_274,N_9971,N_9031);
and UO_275 (O_275,N_9974,N_9266);
and UO_276 (O_276,N_9246,N_9094);
and UO_277 (O_277,N_9405,N_9834);
nand UO_278 (O_278,N_9255,N_9523);
nor UO_279 (O_279,N_9286,N_9217);
and UO_280 (O_280,N_9277,N_9938);
or UO_281 (O_281,N_9000,N_9273);
nand UO_282 (O_282,N_9882,N_9399);
or UO_283 (O_283,N_9487,N_9379);
nor UO_284 (O_284,N_9274,N_9679);
and UO_285 (O_285,N_9026,N_9053);
nand UO_286 (O_286,N_9634,N_9758);
or UO_287 (O_287,N_9762,N_9784);
nor UO_288 (O_288,N_9252,N_9491);
or UO_289 (O_289,N_9556,N_9564);
and UO_290 (O_290,N_9942,N_9957);
and UO_291 (O_291,N_9747,N_9881);
nand UO_292 (O_292,N_9968,N_9073);
nor UO_293 (O_293,N_9769,N_9099);
and UO_294 (O_294,N_9789,N_9140);
nand UO_295 (O_295,N_9114,N_9205);
nor UO_296 (O_296,N_9150,N_9478);
nor UO_297 (O_297,N_9991,N_9078);
and UO_298 (O_298,N_9007,N_9443);
or UO_299 (O_299,N_9774,N_9048);
or UO_300 (O_300,N_9363,N_9907);
and UO_301 (O_301,N_9744,N_9296);
and UO_302 (O_302,N_9310,N_9129);
nand UO_303 (O_303,N_9707,N_9465);
or UO_304 (O_304,N_9257,N_9810);
nand UO_305 (O_305,N_9577,N_9959);
nor UO_306 (O_306,N_9365,N_9344);
or UO_307 (O_307,N_9020,N_9229);
and UO_308 (O_308,N_9284,N_9178);
or UO_309 (O_309,N_9990,N_9175);
and UO_310 (O_310,N_9389,N_9156);
and UO_311 (O_311,N_9155,N_9371);
and UO_312 (O_312,N_9540,N_9824);
nor UO_313 (O_313,N_9025,N_9448);
or UO_314 (O_314,N_9018,N_9431);
nor UO_315 (O_315,N_9668,N_9168);
or UO_316 (O_316,N_9546,N_9694);
nor UO_317 (O_317,N_9797,N_9411);
and UO_318 (O_318,N_9261,N_9136);
nand UO_319 (O_319,N_9703,N_9475);
nand UO_320 (O_320,N_9460,N_9119);
nand UO_321 (O_321,N_9983,N_9315);
nand UO_322 (O_322,N_9298,N_9199);
and UO_323 (O_323,N_9373,N_9851);
nand UO_324 (O_324,N_9953,N_9629);
nor UO_325 (O_325,N_9626,N_9488);
and UO_326 (O_326,N_9345,N_9801);
and UO_327 (O_327,N_9244,N_9960);
nor UO_328 (O_328,N_9892,N_9462);
and UO_329 (O_329,N_9921,N_9705);
nor UO_330 (O_330,N_9793,N_9250);
or UO_331 (O_331,N_9110,N_9997);
nand UO_332 (O_332,N_9498,N_9534);
nor UO_333 (O_333,N_9642,N_9911);
nand UO_334 (O_334,N_9416,N_9123);
and UO_335 (O_335,N_9509,N_9858);
and UO_336 (O_336,N_9676,N_9299);
nand UO_337 (O_337,N_9547,N_9649);
or UO_338 (O_338,N_9792,N_9646);
and UO_339 (O_339,N_9495,N_9457);
and UO_340 (O_340,N_9400,N_9468);
nor UO_341 (O_341,N_9560,N_9717);
or UO_342 (O_342,N_9508,N_9455);
nand UO_343 (O_343,N_9752,N_9607);
nand UO_344 (O_344,N_9165,N_9499);
nor UO_345 (O_345,N_9763,N_9624);
xnor UO_346 (O_346,N_9700,N_9173);
nor UO_347 (O_347,N_9001,N_9639);
or UO_348 (O_348,N_9620,N_9441);
nor UO_349 (O_349,N_9347,N_9969);
or UO_350 (O_350,N_9055,N_9181);
nand UO_351 (O_351,N_9063,N_9768);
nand UO_352 (O_352,N_9328,N_9506);
or UO_353 (O_353,N_9850,N_9137);
nor UO_354 (O_354,N_9689,N_9423);
xor UO_355 (O_355,N_9248,N_9928);
and UO_356 (O_356,N_9514,N_9230);
nand UO_357 (O_357,N_9600,N_9706);
or UO_358 (O_358,N_9224,N_9552);
nand UO_359 (O_359,N_9195,N_9777);
nand UO_360 (O_360,N_9392,N_9606);
nor UO_361 (O_361,N_9135,N_9684);
or UO_362 (O_362,N_9650,N_9627);
and UO_363 (O_363,N_9608,N_9616);
or UO_364 (O_364,N_9104,N_9242);
nor UO_365 (O_365,N_9011,N_9822);
or UO_366 (O_366,N_9544,N_9521);
or UO_367 (O_367,N_9887,N_9081);
or UO_368 (O_368,N_9243,N_9046);
or UO_369 (O_369,N_9972,N_9729);
nand UO_370 (O_370,N_9662,N_9074);
nand UO_371 (O_371,N_9446,N_9236);
and UO_372 (O_372,N_9670,N_9262);
and UO_373 (O_373,N_9340,N_9169);
nand UO_374 (O_374,N_9429,N_9490);
or UO_375 (O_375,N_9037,N_9711);
nor UO_376 (O_376,N_9313,N_9505);
nand UO_377 (O_377,N_9306,N_9811);
nor UO_378 (O_378,N_9967,N_9263);
nand UO_379 (O_379,N_9691,N_9378);
nand UO_380 (O_380,N_9829,N_9336);
or UO_381 (O_381,N_9896,N_9332);
or UO_382 (O_382,N_9868,N_9069);
or UO_383 (O_383,N_9760,N_9580);
and UO_384 (O_384,N_9105,N_9951);
nor UO_385 (O_385,N_9826,N_9776);
nor UO_386 (O_386,N_9134,N_9541);
or UO_387 (O_387,N_9751,N_9045);
nand UO_388 (O_388,N_9413,N_9767);
nand UO_389 (O_389,N_9113,N_9757);
or UO_390 (O_390,N_9177,N_9783);
or UO_391 (O_391,N_9154,N_9726);
or UO_392 (O_392,N_9420,N_9272);
nand UO_393 (O_393,N_9927,N_9849);
or UO_394 (O_394,N_9725,N_9238);
nor UO_395 (O_395,N_9235,N_9440);
nor UO_396 (O_396,N_9280,N_9736);
nor UO_397 (O_397,N_9770,N_9741);
nand UO_398 (O_398,N_9516,N_9267);
and UO_399 (O_399,N_9393,N_9288);
nor UO_400 (O_400,N_9507,N_9339);
nand UO_401 (O_401,N_9978,N_9153);
and UO_402 (O_402,N_9865,N_9112);
nor UO_403 (O_403,N_9559,N_9635);
and UO_404 (O_404,N_9815,N_9318);
or UO_405 (O_405,N_9567,N_9355);
nand UO_406 (O_406,N_9721,N_9551);
nand UO_407 (O_407,N_9022,N_9867);
nand UO_408 (O_408,N_9410,N_9481);
and UO_409 (O_409,N_9324,N_9186);
or UO_410 (O_410,N_9401,N_9982);
or UO_411 (O_411,N_9732,N_9152);
nor UO_412 (O_412,N_9903,N_9592);
nor UO_413 (O_413,N_9415,N_9915);
or UO_414 (O_414,N_9528,N_9086);
nand UO_415 (O_415,N_9279,N_9167);
nor UO_416 (O_416,N_9066,N_9814);
or UO_417 (O_417,N_9864,N_9390);
nand UO_418 (O_418,N_9179,N_9290);
nor UO_419 (O_419,N_9374,N_9584);
or UO_420 (O_420,N_9727,N_9361);
nand UO_421 (O_421,N_9148,N_9667);
nor UO_422 (O_422,N_9833,N_9028);
nand UO_423 (O_423,N_9910,N_9040);
nand UO_424 (O_424,N_9597,N_9068);
nor UO_425 (O_425,N_9593,N_9542);
nand UO_426 (O_426,N_9963,N_9386);
nand UO_427 (O_427,N_9880,N_9895);
nand UO_428 (O_428,N_9645,N_9790);
and UO_429 (O_429,N_9976,N_9731);
or UO_430 (O_430,N_9581,N_9820);
nor UO_431 (O_431,N_9115,N_9124);
and UO_432 (O_432,N_9520,N_9061);
or UO_433 (O_433,N_9527,N_9722);
nand UO_434 (O_434,N_9322,N_9871);
nand UO_435 (O_435,N_9285,N_9343);
and UO_436 (O_436,N_9225,N_9809);
nor UO_437 (O_437,N_9533,N_9569);
nand UO_438 (O_438,N_9377,N_9738);
nor UO_439 (O_439,N_9599,N_9614);
nor UO_440 (O_440,N_9418,N_9424);
nor UO_441 (O_441,N_9188,N_9579);
nor UO_442 (O_442,N_9734,N_9130);
and UO_443 (O_443,N_9748,N_9333);
nor UO_444 (O_444,N_9659,N_9771);
or UO_445 (O_445,N_9259,N_9989);
nand UO_446 (O_446,N_9171,N_9926);
or UO_447 (O_447,N_9633,N_9351);
nor UO_448 (O_448,N_9003,N_9945);
or UO_449 (O_449,N_9208,N_9796);
nor UO_450 (O_450,N_9902,N_9043);
or UO_451 (O_451,N_9573,N_9125);
nand UO_452 (O_452,N_9524,N_9019);
and UO_453 (O_453,N_9589,N_9621);
nor UO_454 (O_454,N_9014,N_9453);
nor UO_455 (O_455,N_9883,N_9258);
and UO_456 (O_456,N_9739,N_9433);
or UO_457 (O_457,N_9008,N_9038);
xor UO_458 (O_458,N_9779,N_9311);
and UO_459 (O_459,N_9719,N_9075);
nor UO_460 (O_460,N_9159,N_9452);
and UO_461 (O_461,N_9539,N_9445);
or UO_462 (O_462,N_9394,N_9309);
or UO_463 (O_463,N_9447,N_9781);
or UO_464 (O_464,N_9715,N_9422);
nor UO_465 (O_465,N_9830,N_9030);
nand UO_466 (O_466,N_9975,N_9866);
nor UO_467 (O_467,N_9197,N_9875);
and UO_468 (O_468,N_9550,N_9764);
nand UO_469 (O_469,N_9385,N_9828);
nand UO_470 (O_470,N_9807,N_9409);
nor UO_471 (O_471,N_9837,N_9622);
and UO_472 (O_472,N_9935,N_9088);
nor UO_473 (O_473,N_9459,N_9100);
and UO_474 (O_474,N_9049,N_9695);
nor UO_475 (O_475,N_9702,N_9461);
or UO_476 (O_476,N_9555,N_9317);
or UO_477 (O_477,N_9653,N_9955);
nand UO_478 (O_478,N_9057,N_9743);
or UO_479 (O_479,N_9888,N_9304);
nor UO_480 (O_480,N_9733,N_9788);
and UO_481 (O_481,N_9798,N_9939);
or UO_482 (O_482,N_9193,N_9044);
and UO_483 (O_483,N_9486,N_9141);
and UO_484 (O_484,N_9128,N_9477);
or UO_485 (O_485,N_9245,N_9147);
nand UO_486 (O_486,N_9421,N_9832);
or UO_487 (O_487,N_9613,N_9529);
and UO_488 (O_488,N_9759,N_9346);
and UO_489 (O_489,N_9859,N_9944);
and UO_490 (O_490,N_9906,N_9454);
and UO_491 (O_491,N_9537,N_9196);
and UO_492 (O_492,N_9283,N_9909);
and UO_493 (O_493,N_9843,N_9966);
or UO_494 (O_494,N_9742,N_9518);
nor UO_495 (O_495,N_9143,N_9531);
and UO_496 (O_496,N_9636,N_9096);
and UO_497 (O_497,N_9675,N_9561);
nor UO_498 (O_498,N_9214,N_9149);
or UO_499 (O_499,N_9996,N_9591);
nor UO_500 (O_500,N_9677,N_9518);
and UO_501 (O_501,N_9797,N_9871);
and UO_502 (O_502,N_9128,N_9241);
nor UO_503 (O_503,N_9118,N_9549);
xor UO_504 (O_504,N_9406,N_9659);
and UO_505 (O_505,N_9917,N_9483);
nand UO_506 (O_506,N_9397,N_9966);
nor UO_507 (O_507,N_9397,N_9240);
nand UO_508 (O_508,N_9099,N_9515);
nand UO_509 (O_509,N_9014,N_9121);
and UO_510 (O_510,N_9702,N_9701);
nand UO_511 (O_511,N_9930,N_9261);
nand UO_512 (O_512,N_9577,N_9415);
and UO_513 (O_513,N_9339,N_9189);
nor UO_514 (O_514,N_9261,N_9009);
nand UO_515 (O_515,N_9686,N_9052);
nand UO_516 (O_516,N_9085,N_9463);
nor UO_517 (O_517,N_9930,N_9934);
nand UO_518 (O_518,N_9186,N_9784);
nand UO_519 (O_519,N_9002,N_9847);
nor UO_520 (O_520,N_9337,N_9622);
or UO_521 (O_521,N_9958,N_9174);
or UO_522 (O_522,N_9460,N_9290);
and UO_523 (O_523,N_9514,N_9648);
nand UO_524 (O_524,N_9568,N_9104);
nand UO_525 (O_525,N_9222,N_9367);
and UO_526 (O_526,N_9307,N_9374);
and UO_527 (O_527,N_9938,N_9295);
nand UO_528 (O_528,N_9158,N_9778);
and UO_529 (O_529,N_9365,N_9691);
or UO_530 (O_530,N_9111,N_9530);
and UO_531 (O_531,N_9037,N_9549);
nand UO_532 (O_532,N_9434,N_9071);
or UO_533 (O_533,N_9636,N_9359);
nand UO_534 (O_534,N_9854,N_9989);
nand UO_535 (O_535,N_9634,N_9074);
or UO_536 (O_536,N_9821,N_9969);
nor UO_537 (O_537,N_9656,N_9445);
nor UO_538 (O_538,N_9930,N_9839);
nor UO_539 (O_539,N_9129,N_9022);
or UO_540 (O_540,N_9320,N_9108);
or UO_541 (O_541,N_9209,N_9940);
and UO_542 (O_542,N_9125,N_9355);
nand UO_543 (O_543,N_9021,N_9155);
and UO_544 (O_544,N_9743,N_9641);
or UO_545 (O_545,N_9962,N_9742);
and UO_546 (O_546,N_9486,N_9400);
nand UO_547 (O_547,N_9628,N_9117);
nor UO_548 (O_548,N_9581,N_9001);
and UO_549 (O_549,N_9814,N_9617);
or UO_550 (O_550,N_9714,N_9672);
nand UO_551 (O_551,N_9817,N_9333);
nand UO_552 (O_552,N_9075,N_9345);
nor UO_553 (O_553,N_9080,N_9023);
nor UO_554 (O_554,N_9238,N_9762);
or UO_555 (O_555,N_9964,N_9877);
nor UO_556 (O_556,N_9845,N_9388);
and UO_557 (O_557,N_9457,N_9182);
nand UO_558 (O_558,N_9772,N_9019);
or UO_559 (O_559,N_9821,N_9971);
nand UO_560 (O_560,N_9358,N_9674);
nor UO_561 (O_561,N_9346,N_9386);
nor UO_562 (O_562,N_9295,N_9521);
or UO_563 (O_563,N_9524,N_9675);
and UO_564 (O_564,N_9556,N_9975);
or UO_565 (O_565,N_9324,N_9260);
and UO_566 (O_566,N_9604,N_9100);
nand UO_567 (O_567,N_9376,N_9309);
xor UO_568 (O_568,N_9860,N_9492);
nand UO_569 (O_569,N_9218,N_9012);
nand UO_570 (O_570,N_9489,N_9784);
or UO_571 (O_571,N_9336,N_9638);
or UO_572 (O_572,N_9377,N_9710);
and UO_573 (O_573,N_9835,N_9378);
nor UO_574 (O_574,N_9725,N_9269);
or UO_575 (O_575,N_9647,N_9184);
or UO_576 (O_576,N_9238,N_9426);
and UO_577 (O_577,N_9759,N_9094);
nor UO_578 (O_578,N_9472,N_9286);
and UO_579 (O_579,N_9051,N_9435);
nand UO_580 (O_580,N_9703,N_9633);
nor UO_581 (O_581,N_9381,N_9361);
and UO_582 (O_582,N_9486,N_9444);
xnor UO_583 (O_583,N_9074,N_9928);
and UO_584 (O_584,N_9099,N_9282);
nor UO_585 (O_585,N_9265,N_9216);
and UO_586 (O_586,N_9072,N_9519);
nand UO_587 (O_587,N_9919,N_9780);
nor UO_588 (O_588,N_9236,N_9960);
and UO_589 (O_589,N_9031,N_9128);
and UO_590 (O_590,N_9472,N_9510);
or UO_591 (O_591,N_9693,N_9633);
and UO_592 (O_592,N_9433,N_9878);
or UO_593 (O_593,N_9277,N_9825);
or UO_594 (O_594,N_9629,N_9213);
nor UO_595 (O_595,N_9777,N_9674);
nand UO_596 (O_596,N_9974,N_9269);
and UO_597 (O_597,N_9850,N_9271);
or UO_598 (O_598,N_9090,N_9803);
or UO_599 (O_599,N_9426,N_9977);
and UO_600 (O_600,N_9216,N_9789);
and UO_601 (O_601,N_9494,N_9881);
nor UO_602 (O_602,N_9830,N_9702);
nor UO_603 (O_603,N_9703,N_9710);
nor UO_604 (O_604,N_9633,N_9262);
nand UO_605 (O_605,N_9208,N_9143);
nor UO_606 (O_606,N_9479,N_9682);
nor UO_607 (O_607,N_9355,N_9661);
and UO_608 (O_608,N_9475,N_9335);
and UO_609 (O_609,N_9861,N_9176);
or UO_610 (O_610,N_9651,N_9396);
or UO_611 (O_611,N_9128,N_9744);
and UO_612 (O_612,N_9342,N_9127);
nor UO_613 (O_613,N_9464,N_9325);
nor UO_614 (O_614,N_9974,N_9658);
nor UO_615 (O_615,N_9673,N_9092);
nand UO_616 (O_616,N_9674,N_9789);
or UO_617 (O_617,N_9103,N_9176);
nand UO_618 (O_618,N_9933,N_9899);
nand UO_619 (O_619,N_9149,N_9017);
and UO_620 (O_620,N_9879,N_9175);
nand UO_621 (O_621,N_9962,N_9622);
nor UO_622 (O_622,N_9768,N_9184);
nand UO_623 (O_623,N_9882,N_9317);
nor UO_624 (O_624,N_9484,N_9324);
nor UO_625 (O_625,N_9975,N_9385);
and UO_626 (O_626,N_9087,N_9099);
nand UO_627 (O_627,N_9539,N_9101);
or UO_628 (O_628,N_9092,N_9052);
nand UO_629 (O_629,N_9369,N_9883);
or UO_630 (O_630,N_9501,N_9957);
nor UO_631 (O_631,N_9552,N_9818);
or UO_632 (O_632,N_9628,N_9107);
and UO_633 (O_633,N_9639,N_9431);
nor UO_634 (O_634,N_9771,N_9498);
and UO_635 (O_635,N_9866,N_9864);
nand UO_636 (O_636,N_9831,N_9673);
nor UO_637 (O_637,N_9109,N_9175);
and UO_638 (O_638,N_9367,N_9123);
nand UO_639 (O_639,N_9160,N_9232);
and UO_640 (O_640,N_9346,N_9293);
xor UO_641 (O_641,N_9202,N_9151);
nand UO_642 (O_642,N_9083,N_9511);
nand UO_643 (O_643,N_9153,N_9042);
and UO_644 (O_644,N_9870,N_9495);
nand UO_645 (O_645,N_9112,N_9324);
nor UO_646 (O_646,N_9917,N_9181);
nand UO_647 (O_647,N_9153,N_9968);
nor UO_648 (O_648,N_9537,N_9097);
nand UO_649 (O_649,N_9758,N_9467);
nand UO_650 (O_650,N_9624,N_9315);
nor UO_651 (O_651,N_9935,N_9276);
or UO_652 (O_652,N_9393,N_9149);
xor UO_653 (O_653,N_9624,N_9718);
nor UO_654 (O_654,N_9224,N_9859);
and UO_655 (O_655,N_9410,N_9051);
xor UO_656 (O_656,N_9180,N_9040);
or UO_657 (O_657,N_9057,N_9089);
nor UO_658 (O_658,N_9610,N_9037);
and UO_659 (O_659,N_9439,N_9676);
or UO_660 (O_660,N_9019,N_9103);
or UO_661 (O_661,N_9474,N_9088);
nand UO_662 (O_662,N_9099,N_9104);
xor UO_663 (O_663,N_9763,N_9890);
nor UO_664 (O_664,N_9332,N_9395);
nand UO_665 (O_665,N_9687,N_9185);
or UO_666 (O_666,N_9705,N_9252);
nor UO_667 (O_667,N_9160,N_9826);
nor UO_668 (O_668,N_9844,N_9309);
or UO_669 (O_669,N_9858,N_9584);
xor UO_670 (O_670,N_9448,N_9592);
nor UO_671 (O_671,N_9807,N_9026);
nor UO_672 (O_672,N_9737,N_9137);
nor UO_673 (O_673,N_9248,N_9547);
nor UO_674 (O_674,N_9845,N_9264);
nor UO_675 (O_675,N_9368,N_9881);
nor UO_676 (O_676,N_9264,N_9205);
nor UO_677 (O_677,N_9381,N_9095);
nand UO_678 (O_678,N_9554,N_9180);
nor UO_679 (O_679,N_9892,N_9026);
and UO_680 (O_680,N_9028,N_9084);
and UO_681 (O_681,N_9960,N_9261);
nand UO_682 (O_682,N_9905,N_9868);
nor UO_683 (O_683,N_9022,N_9989);
and UO_684 (O_684,N_9287,N_9763);
nand UO_685 (O_685,N_9444,N_9369);
nand UO_686 (O_686,N_9484,N_9336);
nand UO_687 (O_687,N_9381,N_9956);
xor UO_688 (O_688,N_9905,N_9736);
or UO_689 (O_689,N_9598,N_9430);
nor UO_690 (O_690,N_9516,N_9719);
nand UO_691 (O_691,N_9410,N_9257);
nand UO_692 (O_692,N_9601,N_9267);
nor UO_693 (O_693,N_9089,N_9410);
and UO_694 (O_694,N_9862,N_9169);
nand UO_695 (O_695,N_9918,N_9828);
or UO_696 (O_696,N_9438,N_9618);
nand UO_697 (O_697,N_9416,N_9069);
and UO_698 (O_698,N_9305,N_9093);
and UO_699 (O_699,N_9515,N_9125);
nand UO_700 (O_700,N_9408,N_9480);
or UO_701 (O_701,N_9918,N_9879);
or UO_702 (O_702,N_9636,N_9089);
or UO_703 (O_703,N_9227,N_9435);
and UO_704 (O_704,N_9192,N_9113);
nor UO_705 (O_705,N_9102,N_9095);
nor UO_706 (O_706,N_9688,N_9095);
nor UO_707 (O_707,N_9427,N_9001);
nor UO_708 (O_708,N_9840,N_9709);
and UO_709 (O_709,N_9248,N_9936);
nand UO_710 (O_710,N_9672,N_9811);
and UO_711 (O_711,N_9369,N_9905);
and UO_712 (O_712,N_9667,N_9708);
and UO_713 (O_713,N_9499,N_9808);
nor UO_714 (O_714,N_9374,N_9611);
nand UO_715 (O_715,N_9997,N_9193);
and UO_716 (O_716,N_9584,N_9928);
nor UO_717 (O_717,N_9900,N_9661);
nand UO_718 (O_718,N_9697,N_9246);
nor UO_719 (O_719,N_9104,N_9834);
nor UO_720 (O_720,N_9998,N_9900);
nand UO_721 (O_721,N_9883,N_9545);
nand UO_722 (O_722,N_9512,N_9554);
nand UO_723 (O_723,N_9485,N_9074);
and UO_724 (O_724,N_9429,N_9702);
nand UO_725 (O_725,N_9412,N_9516);
and UO_726 (O_726,N_9487,N_9991);
and UO_727 (O_727,N_9047,N_9279);
nand UO_728 (O_728,N_9399,N_9823);
and UO_729 (O_729,N_9068,N_9429);
and UO_730 (O_730,N_9974,N_9591);
or UO_731 (O_731,N_9955,N_9791);
nand UO_732 (O_732,N_9386,N_9334);
or UO_733 (O_733,N_9202,N_9440);
nor UO_734 (O_734,N_9242,N_9634);
and UO_735 (O_735,N_9446,N_9498);
or UO_736 (O_736,N_9387,N_9053);
nor UO_737 (O_737,N_9616,N_9994);
nor UO_738 (O_738,N_9819,N_9185);
or UO_739 (O_739,N_9851,N_9683);
nor UO_740 (O_740,N_9462,N_9408);
nand UO_741 (O_741,N_9823,N_9323);
nor UO_742 (O_742,N_9081,N_9201);
and UO_743 (O_743,N_9637,N_9563);
or UO_744 (O_744,N_9129,N_9815);
nor UO_745 (O_745,N_9311,N_9306);
nand UO_746 (O_746,N_9044,N_9054);
or UO_747 (O_747,N_9672,N_9240);
or UO_748 (O_748,N_9571,N_9667);
nor UO_749 (O_749,N_9934,N_9570);
or UO_750 (O_750,N_9912,N_9275);
nand UO_751 (O_751,N_9982,N_9462);
nor UO_752 (O_752,N_9181,N_9855);
xnor UO_753 (O_753,N_9501,N_9387);
and UO_754 (O_754,N_9756,N_9766);
nor UO_755 (O_755,N_9408,N_9907);
nor UO_756 (O_756,N_9071,N_9460);
and UO_757 (O_757,N_9781,N_9111);
nand UO_758 (O_758,N_9348,N_9901);
and UO_759 (O_759,N_9756,N_9206);
nor UO_760 (O_760,N_9389,N_9338);
or UO_761 (O_761,N_9139,N_9582);
and UO_762 (O_762,N_9310,N_9009);
or UO_763 (O_763,N_9855,N_9409);
nor UO_764 (O_764,N_9223,N_9688);
and UO_765 (O_765,N_9883,N_9428);
nor UO_766 (O_766,N_9288,N_9315);
nand UO_767 (O_767,N_9192,N_9521);
or UO_768 (O_768,N_9646,N_9690);
or UO_769 (O_769,N_9676,N_9026);
nand UO_770 (O_770,N_9582,N_9824);
and UO_771 (O_771,N_9321,N_9361);
and UO_772 (O_772,N_9273,N_9795);
and UO_773 (O_773,N_9840,N_9696);
nor UO_774 (O_774,N_9431,N_9610);
nor UO_775 (O_775,N_9168,N_9947);
or UO_776 (O_776,N_9119,N_9204);
or UO_777 (O_777,N_9514,N_9212);
nand UO_778 (O_778,N_9268,N_9113);
or UO_779 (O_779,N_9504,N_9600);
and UO_780 (O_780,N_9310,N_9967);
and UO_781 (O_781,N_9085,N_9243);
nand UO_782 (O_782,N_9199,N_9413);
nor UO_783 (O_783,N_9365,N_9018);
and UO_784 (O_784,N_9770,N_9570);
nand UO_785 (O_785,N_9720,N_9809);
nand UO_786 (O_786,N_9053,N_9413);
nor UO_787 (O_787,N_9193,N_9847);
or UO_788 (O_788,N_9510,N_9452);
nand UO_789 (O_789,N_9568,N_9299);
nand UO_790 (O_790,N_9996,N_9237);
nor UO_791 (O_791,N_9143,N_9373);
or UO_792 (O_792,N_9611,N_9294);
nand UO_793 (O_793,N_9345,N_9446);
and UO_794 (O_794,N_9124,N_9514);
nor UO_795 (O_795,N_9641,N_9844);
or UO_796 (O_796,N_9291,N_9247);
nand UO_797 (O_797,N_9439,N_9317);
nand UO_798 (O_798,N_9170,N_9893);
or UO_799 (O_799,N_9819,N_9092);
nor UO_800 (O_800,N_9405,N_9970);
nor UO_801 (O_801,N_9698,N_9951);
nand UO_802 (O_802,N_9651,N_9594);
or UO_803 (O_803,N_9215,N_9966);
xnor UO_804 (O_804,N_9859,N_9370);
nand UO_805 (O_805,N_9546,N_9299);
nor UO_806 (O_806,N_9181,N_9861);
and UO_807 (O_807,N_9373,N_9282);
and UO_808 (O_808,N_9567,N_9298);
nand UO_809 (O_809,N_9945,N_9976);
nand UO_810 (O_810,N_9955,N_9169);
and UO_811 (O_811,N_9426,N_9244);
or UO_812 (O_812,N_9751,N_9033);
nand UO_813 (O_813,N_9061,N_9624);
nand UO_814 (O_814,N_9827,N_9416);
and UO_815 (O_815,N_9946,N_9293);
or UO_816 (O_816,N_9004,N_9838);
nand UO_817 (O_817,N_9207,N_9384);
nor UO_818 (O_818,N_9482,N_9612);
nand UO_819 (O_819,N_9252,N_9444);
nor UO_820 (O_820,N_9264,N_9879);
nand UO_821 (O_821,N_9183,N_9874);
nor UO_822 (O_822,N_9411,N_9423);
nor UO_823 (O_823,N_9517,N_9922);
and UO_824 (O_824,N_9526,N_9382);
nand UO_825 (O_825,N_9093,N_9510);
and UO_826 (O_826,N_9678,N_9799);
nor UO_827 (O_827,N_9643,N_9736);
xnor UO_828 (O_828,N_9688,N_9972);
and UO_829 (O_829,N_9783,N_9314);
nor UO_830 (O_830,N_9269,N_9597);
nand UO_831 (O_831,N_9529,N_9165);
nand UO_832 (O_832,N_9031,N_9111);
or UO_833 (O_833,N_9961,N_9163);
and UO_834 (O_834,N_9632,N_9579);
and UO_835 (O_835,N_9818,N_9946);
and UO_836 (O_836,N_9576,N_9298);
or UO_837 (O_837,N_9145,N_9983);
nand UO_838 (O_838,N_9507,N_9553);
or UO_839 (O_839,N_9317,N_9075);
or UO_840 (O_840,N_9195,N_9240);
nand UO_841 (O_841,N_9045,N_9294);
and UO_842 (O_842,N_9430,N_9768);
nand UO_843 (O_843,N_9002,N_9152);
xor UO_844 (O_844,N_9362,N_9133);
nor UO_845 (O_845,N_9684,N_9037);
and UO_846 (O_846,N_9311,N_9742);
and UO_847 (O_847,N_9891,N_9472);
nor UO_848 (O_848,N_9153,N_9213);
or UO_849 (O_849,N_9177,N_9087);
nor UO_850 (O_850,N_9378,N_9376);
and UO_851 (O_851,N_9644,N_9671);
nor UO_852 (O_852,N_9985,N_9656);
nor UO_853 (O_853,N_9390,N_9714);
nand UO_854 (O_854,N_9756,N_9029);
or UO_855 (O_855,N_9641,N_9638);
or UO_856 (O_856,N_9117,N_9081);
xnor UO_857 (O_857,N_9928,N_9683);
nor UO_858 (O_858,N_9796,N_9933);
and UO_859 (O_859,N_9806,N_9628);
or UO_860 (O_860,N_9785,N_9707);
nand UO_861 (O_861,N_9913,N_9338);
nand UO_862 (O_862,N_9156,N_9916);
and UO_863 (O_863,N_9847,N_9875);
nor UO_864 (O_864,N_9856,N_9672);
or UO_865 (O_865,N_9760,N_9182);
or UO_866 (O_866,N_9149,N_9026);
and UO_867 (O_867,N_9311,N_9485);
or UO_868 (O_868,N_9919,N_9950);
and UO_869 (O_869,N_9966,N_9806);
or UO_870 (O_870,N_9130,N_9673);
or UO_871 (O_871,N_9630,N_9889);
nand UO_872 (O_872,N_9368,N_9739);
or UO_873 (O_873,N_9327,N_9196);
nand UO_874 (O_874,N_9180,N_9176);
nand UO_875 (O_875,N_9420,N_9488);
and UO_876 (O_876,N_9135,N_9645);
nor UO_877 (O_877,N_9610,N_9562);
nand UO_878 (O_878,N_9177,N_9103);
and UO_879 (O_879,N_9840,N_9665);
or UO_880 (O_880,N_9831,N_9981);
nand UO_881 (O_881,N_9252,N_9365);
and UO_882 (O_882,N_9613,N_9528);
or UO_883 (O_883,N_9573,N_9389);
xor UO_884 (O_884,N_9819,N_9475);
nand UO_885 (O_885,N_9677,N_9816);
xnor UO_886 (O_886,N_9012,N_9758);
and UO_887 (O_887,N_9548,N_9385);
nand UO_888 (O_888,N_9900,N_9358);
and UO_889 (O_889,N_9524,N_9573);
nor UO_890 (O_890,N_9735,N_9322);
and UO_891 (O_891,N_9129,N_9590);
nor UO_892 (O_892,N_9077,N_9156);
nor UO_893 (O_893,N_9507,N_9748);
nor UO_894 (O_894,N_9061,N_9486);
nand UO_895 (O_895,N_9113,N_9194);
or UO_896 (O_896,N_9281,N_9090);
and UO_897 (O_897,N_9432,N_9377);
nand UO_898 (O_898,N_9964,N_9676);
or UO_899 (O_899,N_9521,N_9686);
and UO_900 (O_900,N_9481,N_9019);
and UO_901 (O_901,N_9373,N_9593);
and UO_902 (O_902,N_9583,N_9222);
or UO_903 (O_903,N_9825,N_9586);
and UO_904 (O_904,N_9035,N_9103);
nand UO_905 (O_905,N_9587,N_9510);
or UO_906 (O_906,N_9750,N_9572);
and UO_907 (O_907,N_9811,N_9797);
nor UO_908 (O_908,N_9178,N_9314);
nand UO_909 (O_909,N_9900,N_9651);
or UO_910 (O_910,N_9178,N_9166);
nor UO_911 (O_911,N_9912,N_9574);
and UO_912 (O_912,N_9997,N_9833);
nor UO_913 (O_913,N_9753,N_9512);
nand UO_914 (O_914,N_9507,N_9047);
or UO_915 (O_915,N_9241,N_9939);
nor UO_916 (O_916,N_9950,N_9517);
nor UO_917 (O_917,N_9436,N_9029);
nor UO_918 (O_918,N_9704,N_9281);
nor UO_919 (O_919,N_9668,N_9719);
nor UO_920 (O_920,N_9497,N_9400);
nor UO_921 (O_921,N_9141,N_9785);
and UO_922 (O_922,N_9844,N_9308);
or UO_923 (O_923,N_9197,N_9387);
or UO_924 (O_924,N_9296,N_9382);
or UO_925 (O_925,N_9002,N_9770);
and UO_926 (O_926,N_9343,N_9695);
or UO_927 (O_927,N_9072,N_9493);
nor UO_928 (O_928,N_9634,N_9144);
nand UO_929 (O_929,N_9163,N_9531);
and UO_930 (O_930,N_9620,N_9972);
nand UO_931 (O_931,N_9033,N_9127);
or UO_932 (O_932,N_9023,N_9631);
or UO_933 (O_933,N_9374,N_9930);
nand UO_934 (O_934,N_9180,N_9254);
nand UO_935 (O_935,N_9704,N_9280);
and UO_936 (O_936,N_9050,N_9434);
nand UO_937 (O_937,N_9650,N_9708);
and UO_938 (O_938,N_9745,N_9692);
nor UO_939 (O_939,N_9617,N_9116);
nor UO_940 (O_940,N_9702,N_9963);
nor UO_941 (O_941,N_9923,N_9348);
nor UO_942 (O_942,N_9546,N_9480);
nand UO_943 (O_943,N_9699,N_9205);
and UO_944 (O_944,N_9856,N_9663);
or UO_945 (O_945,N_9673,N_9065);
or UO_946 (O_946,N_9844,N_9505);
or UO_947 (O_947,N_9577,N_9535);
nor UO_948 (O_948,N_9293,N_9636);
nand UO_949 (O_949,N_9729,N_9960);
nand UO_950 (O_950,N_9622,N_9277);
and UO_951 (O_951,N_9168,N_9602);
or UO_952 (O_952,N_9876,N_9696);
nor UO_953 (O_953,N_9133,N_9265);
and UO_954 (O_954,N_9242,N_9584);
and UO_955 (O_955,N_9011,N_9680);
or UO_956 (O_956,N_9913,N_9053);
and UO_957 (O_957,N_9162,N_9948);
and UO_958 (O_958,N_9708,N_9365);
or UO_959 (O_959,N_9251,N_9853);
or UO_960 (O_960,N_9231,N_9482);
or UO_961 (O_961,N_9535,N_9369);
nand UO_962 (O_962,N_9159,N_9451);
and UO_963 (O_963,N_9134,N_9871);
nor UO_964 (O_964,N_9427,N_9502);
nand UO_965 (O_965,N_9065,N_9559);
and UO_966 (O_966,N_9663,N_9189);
or UO_967 (O_967,N_9489,N_9314);
nor UO_968 (O_968,N_9920,N_9330);
nand UO_969 (O_969,N_9712,N_9921);
or UO_970 (O_970,N_9946,N_9379);
or UO_971 (O_971,N_9395,N_9936);
and UO_972 (O_972,N_9601,N_9459);
nand UO_973 (O_973,N_9100,N_9494);
or UO_974 (O_974,N_9553,N_9873);
or UO_975 (O_975,N_9683,N_9231);
nand UO_976 (O_976,N_9597,N_9136);
nor UO_977 (O_977,N_9993,N_9481);
nand UO_978 (O_978,N_9998,N_9185);
nand UO_979 (O_979,N_9362,N_9155);
nor UO_980 (O_980,N_9436,N_9557);
and UO_981 (O_981,N_9124,N_9642);
or UO_982 (O_982,N_9551,N_9871);
nor UO_983 (O_983,N_9628,N_9453);
xnor UO_984 (O_984,N_9350,N_9732);
nor UO_985 (O_985,N_9038,N_9472);
and UO_986 (O_986,N_9429,N_9910);
or UO_987 (O_987,N_9045,N_9108);
nand UO_988 (O_988,N_9768,N_9612);
nand UO_989 (O_989,N_9185,N_9358);
and UO_990 (O_990,N_9376,N_9513);
or UO_991 (O_991,N_9290,N_9680);
nand UO_992 (O_992,N_9870,N_9584);
or UO_993 (O_993,N_9838,N_9280);
and UO_994 (O_994,N_9083,N_9843);
nand UO_995 (O_995,N_9589,N_9067);
and UO_996 (O_996,N_9164,N_9067);
nand UO_997 (O_997,N_9888,N_9915);
nor UO_998 (O_998,N_9374,N_9112);
nand UO_999 (O_999,N_9430,N_9246);
or UO_1000 (O_1000,N_9365,N_9109);
nand UO_1001 (O_1001,N_9242,N_9676);
nand UO_1002 (O_1002,N_9136,N_9856);
and UO_1003 (O_1003,N_9047,N_9990);
or UO_1004 (O_1004,N_9031,N_9424);
nand UO_1005 (O_1005,N_9797,N_9732);
nor UO_1006 (O_1006,N_9152,N_9633);
nor UO_1007 (O_1007,N_9586,N_9000);
and UO_1008 (O_1008,N_9416,N_9295);
and UO_1009 (O_1009,N_9590,N_9152);
nor UO_1010 (O_1010,N_9859,N_9317);
nand UO_1011 (O_1011,N_9246,N_9422);
and UO_1012 (O_1012,N_9425,N_9705);
or UO_1013 (O_1013,N_9961,N_9982);
and UO_1014 (O_1014,N_9745,N_9630);
nand UO_1015 (O_1015,N_9329,N_9243);
and UO_1016 (O_1016,N_9786,N_9644);
or UO_1017 (O_1017,N_9552,N_9063);
nor UO_1018 (O_1018,N_9399,N_9053);
or UO_1019 (O_1019,N_9089,N_9326);
xnor UO_1020 (O_1020,N_9762,N_9533);
nor UO_1021 (O_1021,N_9780,N_9847);
or UO_1022 (O_1022,N_9998,N_9027);
or UO_1023 (O_1023,N_9998,N_9337);
and UO_1024 (O_1024,N_9975,N_9809);
nand UO_1025 (O_1025,N_9339,N_9433);
or UO_1026 (O_1026,N_9925,N_9985);
nand UO_1027 (O_1027,N_9295,N_9757);
or UO_1028 (O_1028,N_9150,N_9952);
nor UO_1029 (O_1029,N_9846,N_9761);
and UO_1030 (O_1030,N_9629,N_9507);
nor UO_1031 (O_1031,N_9348,N_9360);
nor UO_1032 (O_1032,N_9575,N_9076);
nor UO_1033 (O_1033,N_9700,N_9395);
nor UO_1034 (O_1034,N_9104,N_9856);
nor UO_1035 (O_1035,N_9202,N_9384);
and UO_1036 (O_1036,N_9306,N_9527);
nor UO_1037 (O_1037,N_9463,N_9723);
and UO_1038 (O_1038,N_9822,N_9374);
or UO_1039 (O_1039,N_9271,N_9706);
or UO_1040 (O_1040,N_9416,N_9585);
nand UO_1041 (O_1041,N_9830,N_9087);
nand UO_1042 (O_1042,N_9790,N_9110);
or UO_1043 (O_1043,N_9411,N_9730);
and UO_1044 (O_1044,N_9535,N_9179);
or UO_1045 (O_1045,N_9113,N_9927);
or UO_1046 (O_1046,N_9801,N_9249);
nand UO_1047 (O_1047,N_9501,N_9262);
nor UO_1048 (O_1048,N_9284,N_9816);
nand UO_1049 (O_1049,N_9954,N_9521);
nor UO_1050 (O_1050,N_9221,N_9438);
or UO_1051 (O_1051,N_9226,N_9065);
nand UO_1052 (O_1052,N_9324,N_9705);
or UO_1053 (O_1053,N_9247,N_9661);
nand UO_1054 (O_1054,N_9178,N_9388);
nor UO_1055 (O_1055,N_9658,N_9139);
nand UO_1056 (O_1056,N_9016,N_9790);
or UO_1057 (O_1057,N_9874,N_9923);
nand UO_1058 (O_1058,N_9963,N_9043);
xor UO_1059 (O_1059,N_9219,N_9751);
and UO_1060 (O_1060,N_9152,N_9389);
nor UO_1061 (O_1061,N_9442,N_9269);
and UO_1062 (O_1062,N_9450,N_9043);
nor UO_1063 (O_1063,N_9526,N_9289);
nand UO_1064 (O_1064,N_9826,N_9224);
nand UO_1065 (O_1065,N_9579,N_9545);
or UO_1066 (O_1066,N_9391,N_9437);
or UO_1067 (O_1067,N_9111,N_9170);
nand UO_1068 (O_1068,N_9786,N_9413);
xnor UO_1069 (O_1069,N_9965,N_9778);
and UO_1070 (O_1070,N_9505,N_9139);
or UO_1071 (O_1071,N_9724,N_9672);
or UO_1072 (O_1072,N_9907,N_9746);
and UO_1073 (O_1073,N_9331,N_9081);
and UO_1074 (O_1074,N_9625,N_9181);
nor UO_1075 (O_1075,N_9965,N_9369);
or UO_1076 (O_1076,N_9097,N_9564);
and UO_1077 (O_1077,N_9655,N_9791);
and UO_1078 (O_1078,N_9521,N_9871);
nand UO_1079 (O_1079,N_9687,N_9451);
nand UO_1080 (O_1080,N_9129,N_9364);
nand UO_1081 (O_1081,N_9977,N_9152);
nor UO_1082 (O_1082,N_9827,N_9819);
and UO_1083 (O_1083,N_9764,N_9300);
or UO_1084 (O_1084,N_9888,N_9162);
or UO_1085 (O_1085,N_9688,N_9954);
nand UO_1086 (O_1086,N_9761,N_9453);
and UO_1087 (O_1087,N_9268,N_9951);
nor UO_1088 (O_1088,N_9754,N_9203);
and UO_1089 (O_1089,N_9276,N_9319);
nor UO_1090 (O_1090,N_9660,N_9472);
or UO_1091 (O_1091,N_9441,N_9818);
or UO_1092 (O_1092,N_9963,N_9790);
nand UO_1093 (O_1093,N_9948,N_9077);
and UO_1094 (O_1094,N_9164,N_9014);
nor UO_1095 (O_1095,N_9164,N_9801);
or UO_1096 (O_1096,N_9105,N_9559);
nor UO_1097 (O_1097,N_9856,N_9524);
nor UO_1098 (O_1098,N_9264,N_9039);
nand UO_1099 (O_1099,N_9325,N_9349);
or UO_1100 (O_1100,N_9893,N_9008);
nor UO_1101 (O_1101,N_9739,N_9913);
nor UO_1102 (O_1102,N_9519,N_9000);
nand UO_1103 (O_1103,N_9421,N_9632);
nand UO_1104 (O_1104,N_9634,N_9173);
nand UO_1105 (O_1105,N_9556,N_9885);
xnor UO_1106 (O_1106,N_9698,N_9235);
nand UO_1107 (O_1107,N_9438,N_9653);
and UO_1108 (O_1108,N_9443,N_9936);
and UO_1109 (O_1109,N_9513,N_9109);
xor UO_1110 (O_1110,N_9849,N_9934);
and UO_1111 (O_1111,N_9663,N_9087);
nand UO_1112 (O_1112,N_9156,N_9942);
nand UO_1113 (O_1113,N_9365,N_9480);
nor UO_1114 (O_1114,N_9198,N_9380);
nand UO_1115 (O_1115,N_9314,N_9880);
xnor UO_1116 (O_1116,N_9284,N_9601);
and UO_1117 (O_1117,N_9640,N_9559);
nand UO_1118 (O_1118,N_9196,N_9611);
nor UO_1119 (O_1119,N_9442,N_9538);
or UO_1120 (O_1120,N_9281,N_9071);
xnor UO_1121 (O_1121,N_9566,N_9643);
nor UO_1122 (O_1122,N_9671,N_9686);
nand UO_1123 (O_1123,N_9860,N_9410);
nor UO_1124 (O_1124,N_9988,N_9896);
and UO_1125 (O_1125,N_9903,N_9044);
and UO_1126 (O_1126,N_9195,N_9735);
nor UO_1127 (O_1127,N_9266,N_9328);
and UO_1128 (O_1128,N_9592,N_9503);
and UO_1129 (O_1129,N_9424,N_9357);
and UO_1130 (O_1130,N_9529,N_9885);
or UO_1131 (O_1131,N_9074,N_9775);
nand UO_1132 (O_1132,N_9757,N_9996);
nand UO_1133 (O_1133,N_9786,N_9252);
nor UO_1134 (O_1134,N_9553,N_9185);
or UO_1135 (O_1135,N_9782,N_9881);
or UO_1136 (O_1136,N_9700,N_9619);
and UO_1137 (O_1137,N_9693,N_9406);
or UO_1138 (O_1138,N_9934,N_9118);
nand UO_1139 (O_1139,N_9075,N_9351);
nor UO_1140 (O_1140,N_9875,N_9391);
nand UO_1141 (O_1141,N_9978,N_9376);
nand UO_1142 (O_1142,N_9893,N_9489);
nand UO_1143 (O_1143,N_9857,N_9586);
or UO_1144 (O_1144,N_9884,N_9525);
or UO_1145 (O_1145,N_9322,N_9320);
or UO_1146 (O_1146,N_9414,N_9087);
xnor UO_1147 (O_1147,N_9398,N_9266);
nand UO_1148 (O_1148,N_9632,N_9027);
or UO_1149 (O_1149,N_9250,N_9116);
nand UO_1150 (O_1150,N_9175,N_9852);
xor UO_1151 (O_1151,N_9510,N_9682);
or UO_1152 (O_1152,N_9718,N_9746);
and UO_1153 (O_1153,N_9391,N_9450);
nand UO_1154 (O_1154,N_9399,N_9484);
or UO_1155 (O_1155,N_9074,N_9331);
and UO_1156 (O_1156,N_9125,N_9778);
nand UO_1157 (O_1157,N_9151,N_9609);
and UO_1158 (O_1158,N_9152,N_9432);
or UO_1159 (O_1159,N_9183,N_9950);
and UO_1160 (O_1160,N_9399,N_9410);
or UO_1161 (O_1161,N_9071,N_9833);
nor UO_1162 (O_1162,N_9980,N_9632);
nor UO_1163 (O_1163,N_9686,N_9246);
or UO_1164 (O_1164,N_9916,N_9805);
nand UO_1165 (O_1165,N_9138,N_9067);
and UO_1166 (O_1166,N_9385,N_9749);
and UO_1167 (O_1167,N_9406,N_9462);
and UO_1168 (O_1168,N_9799,N_9912);
and UO_1169 (O_1169,N_9904,N_9848);
or UO_1170 (O_1170,N_9141,N_9530);
nor UO_1171 (O_1171,N_9593,N_9889);
nand UO_1172 (O_1172,N_9491,N_9012);
and UO_1173 (O_1173,N_9968,N_9766);
nand UO_1174 (O_1174,N_9620,N_9301);
nor UO_1175 (O_1175,N_9906,N_9880);
nand UO_1176 (O_1176,N_9450,N_9761);
nor UO_1177 (O_1177,N_9315,N_9523);
nand UO_1178 (O_1178,N_9594,N_9109);
nand UO_1179 (O_1179,N_9982,N_9252);
nor UO_1180 (O_1180,N_9557,N_9096);
and UO_1181 (O_1181,N_9150,N_9960);
nor UO_1182 (O_1182,N_9361,N_9396);
and UO_1183 (O_1183,N_9320,N_9514);
nand UO_1184 (O_1184,N_9342,N_9224);
nand UO_1185 (O_1185,N_9950,N_9298);
xor UO_1186 (O_1186,N_9104,N_9972);
and UO_1187 (O_1187,N_9199,N_9843);
or UO_1188 (O_1188,N_9900,N_9251);
or UO_1189 (O_1189,N_9219,N_9534);
and UO_1190 (O_1190,N_9222,N_9584);
and UO_1191 (O_1191,N_9116,N_9512);
or UO_1192 (O_1192,N_9397,N_9855);
nand UO_1193 (O_1193,N_9089,N_9481);
nand UO_1194 (O_1194,N_9072,N_9327);
nand UO_1195 (O_1195,N_9103,N_9282);
nand UO_1196 (O_1196,N_9212,N_9226);
nor UO_1197 (O_1197,N_9263,N_9176);
and UO_1198 (O_1198,N_9271,N_9987);
and UO_1199 (O_1199,N_9133,N_9832);
nand UO_1200 (O_1200,N_9217,N_9421);
nand UO_1201 (O_1201,N_9633,N_9648);
or UO_1202 (O_1202,N_9096,N_9245);
or UO_1203 (O_1203,N_9134,N_9153);
or UO_1204 (O_1204,N_9867,N_9547);
and UO_1205 (O_1205,N_9655,N_9047);
and UO_1206 (O_1206,N_9826,N_9728);
xor UO_1207 (O_1207,N_9978,N_9861);
and UO_1208 (O_1208,N_9029,N_9469);
nand UO_1209 (O_1209,N_9255,N_9787);
nor UO_1210 (O_1210,N_9645,N_9566);
or UO_1211 (O_1211,N_9375,N_9957);
nor UO_1212 (O_1212,N_9718,N_9084);
or UO_1213 (O_1213,N_9304,N_9183);
and UO_1214 (O_1214,N_9270,N_9340);
nand UO_1215 (O_1215,N_9459,N_9796);
nor UO_1216 (O_1216,N_9586,N_9584);
nand UO_1217 (O_1217,N_9291,N_9594);
nor UO_1218 (O_1218,N_9481,N_9976);
and UO_1219 (O_1219,N_9806,N_9640);
nor UO_1220 (O_1220,N_9803,N_9882);
or UO_1221 (O_1221,N_9411,N_9955);
nor UO_1222 (O_1222,N_9097,N_9768);
and UO_1223 (O_1223,N_9639,N_9592);
or UO_1224 (O_1224,N_9019,N_9538);
or UO_1225 (O_1225,N_9309,N_9835);
and UO_1226 (O_1226,N_9404,N_9258);
nor UO_1227 (O_1227,N_9418,N_9118);
or UO_1228 (O_1228,N_9742,N_9975);
and UO_1229 (O_1229,N_9630,N_9817);
nand UO_1230 (O_1230,N_9434,N_9380);
and UO_1231 (O_1231,N_9999,N_9820);
and UO_1232 (O_1232,N_9190,N_9677);
nand UO_1233 (O_1233,N_9316,N_9530);
or UO_1234 (O_1234,N_9302,N_9590);
nand UO_1235 (O_1235,N_9982,N_9219);
xnor UO_1236 (O_1236,N_9143,N_9352);
and UO_1237 (O_1237,N_9841,N_9708);
or UO_1238 (O_1238,N_9117,N_9260);
or UO_1239 (O_1239,N_9368,N_9632);
or UO_1240 (O_1240,N_9753,N_9483);
nor UO_1241 (O_1241,N_9591,N_9226);
nand UO_1242 (O_1242,N_9045,N_9560);
and UO_1243 (O_1243,N_9105,N_9503);
nand UO_1244 (O_1244,N_9753,N_9607);
or UO_1245 (O_1245,N_9794,N_9254);
or UO_1246 (O_1246,N_9878,N_9594);
and UO_1247 (O_1247,N_9700,N_9720);
and UO_1248 (O_1248,N_9929,N_9325);
or UO_1249 (O_1249,N_9718,N_9523);
nand UO_1250 (O_1250,N_9088,N_9810);
and UO_1251 (O_1251,N_9704,N_9858);
nand UO_1252 (O_1252,N_9883,N_9789);
or UO_1253 (O_1253,N_9889,N_9937);
or UO_1254 (O_1254,N_9615,N_9734);
or UO_1255 (O_1255,N_9062,N_9736);
and UO_1256 (O_1256,N_9819,N_9336);
and UO_1257 (O_1257,N_9384,N_9403);
and UO_1258 (O_1258,N_9922,N_9228);
or UO_1259 (O_1259,N_9234,N_9544);
nor UO_1260 (O_1260,N_9378,N_9166);
and UO_1261 (O_1261,N_9466,N_9118);
or UO_1262 (O_1262,N_9366,N_9192);
nor UO_1263 (O_1263,N_9195,N_9447);
nor UO_1264 (O_1264,N_9879,N_9442);
and UO_1265 (O_1265,N_9390,N_9960);
and UO_1266 (O_1266,N_9506,N_9724);
and UO_1267 (O_1267,N_9710,N_9206);
nor UO_1268 (O_1268,N_9232,N_9009);
and UO_1269 (O_1269,N_9905,N_9213);
and UO_1270 (O_1270,N_9879,N_9850);
nor UO_1271 (O_1271,N_9644,N_9313);
and UO_1272 (O_1272,N_9251,N_9420);
nand UO_1273 (O_1273,N_9052,N_9945);
or UO_1274 (O_1274,N_9854,N_9506);
or UO_1275 (O_1275,N_9081,N_9456);
and UO_1276 (O_1276,N_9782,N_9943);
xnor UO_1277 (O_1277,N_9715,N_9603);
and UO_1278 (O_1278,N_9091,N_9084);
and UO_1279 (O_1279,N_9523,N_9448);
or UO_1280 (O_1280,N_9342,N_9307);
or UO_1281 (O_1281,N_9173,N_9243);
and UO_1282 (O_1282,N_9253,N_9665);
and UO_1283 (O_1283,N_9696,N_9014);
or UO_1284 (O_1284,N_9112,N_9959);
or UO_1285 (O_1285,N_9953,N_9660);
or UO_1286 (O_1286,N_9508,N_9744);
nor UO_1287 (O_1287,N_9289,N_9355);
nand UO_1288 (O_1288,N_9233,N_9885);
nor UO_1289 (O_1289,N_9958,N_9280);
or UO_1290 (O_1290,N_9270,N_9244);
nand UO_1291 (O_1291,N_9239,N_9254);
or UO_1292 (O_1292,N_9352,N_9978);
nand UO_1293 (O_1293,N_9081,N_9202);
nand UO_1294 (O_1294,N_9780,N_9665);
nor UO_1295 (O_1295,N_9665,N_9548);
nand UO_1296 (O_1296,N_9408,N_9985);
or UO_1297 (O_1297,N_9121,N_9260);
nor UO_1298 (O_1298,N_9198,N_9197);
nor UO_1299 (O_1299,N_9325,N_9291);
and UO_1300 (O_1300,N_9630,N_9765);
and UO_1301 (O_1301,N_9571,N_9580);
and UO_1302 (O_1302,N_9711,N_9668);
or UO_1303 (O_1303,N_9070,N_9295);
nor UO_1304 (O_1304,N_9903,N_9030);
and UO_1305 (O_1305,N_9639,N_9841);
or UO_1306 (O_1306,N_9598,N_9608);
and UO_1307 (O_1307,N_9890,N_9219);
nor UO_1308 (O_1308,N_9179,N_9493);
nand UO_1309 (O_1309,N_9243,N_9854);
nand UO_1310 (O_1310,N_9392,N_9045);
nand UO_1311 (O_1311,N_9360,N_9233);
nor UO_1312 (O_1312,N_9685,N_9989);
nand UO_1313 (O_1313,N_9249,N_9313);
nand UO_1314 (O_1314,N_9020,N_9957);
and UO_1315 (O_1315,N_9822,N_9507);
or UO_1316 (O_1316,N_9912,N_9311);
or UO_1317 (O_1317,N_9142,N_9977);
nand UO_1318 (O_1318,N_9355,N_9371);
nor UO_1319 (O_1319,N_9706,N_9922);
nand UO_1320 (O_1320,N_9304,N_9263);
nand UO_1321 (O_1321,N_9003,N_9083);
and UO_1322 (O_1322,N_9191,N_9897);
or UO_1323 (O_1323,N_9907,N_9853);
nand UO_1324 (O_1324,N_9567,N_9934);
nand UO_1325 (O_1325,N_9253,N_9190);
nand UO_1326 (O_1326,N_9242,N_9450);
and UO_1327 (O_1327,N_9004,N_9499);
nor UO_1328 (O_1328,N_9317,N_9246);
nor UO_1329 (O_1329,N_9010,N_9472);
and UO_1330 (O_1330,N_9398,N_9516);
and UO_1331 (O_1331,N_9113,N_9234);
or UO_1332 (O_1332,N_9842,N_9279);
and UO_1333 (O_1333,N_9040,N_9287);
or UO_1334 (O_1334,N_9059,N_9215);
and UO_1335 (O_1335,N_9768,N_9209);
or UO_1336 (O_1336,N_9998,N_9681);
and UO_1337 (O_1337,N_9183,N_9829);
and UO_1338 (O_1338,N_9045,N_9065);
and UO_1339 (O_1339,N_9589,N_9985);
and UO_1340 (O_1340,N_9282,N_9789);
nor UO_1341 (O_1341,N_9081,N_9570);
and UO_1342 (O_1342,N_9486,N_9642);
nor UO_1343 (O_1343,N_9200,N_9385);
nand UO_1344 (O_1344,N_9544,N_9937);
nor UO_1345 (O_1345,N_9298,N_9319);
or UO_1346 (O_1346,N_9028,N_9193);
nand UO_1347 (O_1347,N_9776,N_9405);
or UO_1348 (O_1348,N_9481,N_9458);
and UO_1349 (O_1349,N_9432,N_9931);
xnor UO_1350 (O_1350,N_9855,N_9904);
or UO_1351 (O_1351,N_9521,N_9241);
or UO_1352 (O_1352,N_9887,N_9949);
nor UO_1353 (O_1353,N_9361,N_9448);
nor UO_1354 (O_1354,N_9019,N_9339);
and UO_1355 (O_1355,N_9921,N_9566);
and UO_1356 (O_1356,N_9793,N_9233);
and UO_1357 (O_1357,N_9630,N_9152);
nand UO_1358 (O_1358,N_9402,N_9866);
and UO_1359 (O_1359,N_9976,N_9640);
or UO_1360 (O_1360,N_9349,N_9922);
nand UO_1361 (O_1361,N_9150,N_9637);
nand UO_1362 (O_1362,N_9714,N_9341);
nor UO_1363 (O_1363,N_9081,N_9227);
or UO_1364 (O_1364,N_9624,N_9673);
and UO_1365 (O_1365,N_9623,N_9426);
nor UO_1366 (O_1366,N_9687,N_9530);
or UO_1367 (O_1367,N_9778,N_9163);
nand UO_1368 (O_1368,N_9663,N_9180);
nor UO_1369 (O_1369,N_9208,N_9114);
nand UO_1370 (O_1370,N_9301,N_9805);
or UO_1371 (O_1371,N_9632,N_9935);
and UO_1372 (O_1372,N_9804,N_9310);
nand UO_1373 (O_1373,N_9879,N_9301);
or UO_1374 (O_1374,N_9408,N_9440);
nand UO_1375 (O_1375,N_9071,N_9817);
and UO_1376 (O_1376,N_9698,N_9154);
nand UO_1377 (O_1377,N_9583,N_9997);
and UO_1378 (O_1378,N_9803,N_9380);
nand UO_1379 (O_1379,N_9652,N_9178);
and UO_1380 (O_1380,N_9736,N_9642);
nand UO_1381 (O_1381,N_9944,N_9305);
nand UO_1382 (O_1382,N_9162,N_9315);
nor UO_1383 (O_1383,N_9052,N_9677);
and UO_1384 (O_1384,N_9407,N_9361);
and UO_1385 (O_1385,N_9747,N_9493);
nor UO_1386 (O_1386,N_9842,N_9290);
nand UO_1387 (O_1387,N_9499,N_9758);
nand UO_1388 (O_1388,N_9319,N_9975);
or UO_1389 (O_1389,N_9875,N_9577);
and UO_1390 (O_1390,N_9883,N_9161);
or UO_1391 (O_1391,N_9549,N_9335);
nor UO_1392 (O_1392,N_9516,N_9173);
or UO_1393 (O_1393,N_9498,N_9024);
or UO_1394 (O_1394,N_9630,N_9587);
or UO_1395 (O_1395,N_9915,N_9218);
or UO_1396 (O_1396,N_9928,N_9081);
nand UO_1397 (O_1397,N_9888,N_9555);
or UO_1398 (O_1398,N_9434,N_9617);
and UO_1399 (O_1399,N_9297,N_9512);
nor UO_1400 (O_1400,N_9407,N_9143);
or UO_1401 (O_1401,N_9551,N_9996);
or UO_1402 (O_1402,N_9521,N_9614);
and UO_1403 (O_1403,N_9752,N_9779);
nand UO_1404 (O_1404,N_9734,N_9839);
nand UO_1405 (O_1405,N_9196,N_9341);
and UO_1406 (O_1406,N_9748,N_9220);
and UO_1407 (O_1407,N_9487,N_9846);
or UO_1408 (O_1408,N_9601,N_9235);
and UO_1409 (O_1409,N_9856,N_9144);
and UO_1410 (O_1410,N_9832,N_9854);
and UO_1411 (O_1411,N_9481,N_9580);
nand UO_1412 (O_1412,N_9855,N_9514);
and UO_1413 (O_1413,N_9253,N_9031);
or UO_1414 (O_1414,N_9058,N_9407);
or UO_1415 (O_1415,N_9689,N_9894);
nor UO_1416 (O_1416,N_9948,N_9961);
or UO_1417 (O_1417,N_9589,N_9765);
xnor UO_1418 (O_1418,N_9874,N_9162);
nand UO_1419 (O_1419,N_9144,N_9459);
and UO_1420 (O_1420,N_9913,N_9825);
or UO_1421 (O_1421,N_9057,N_9704);
and UO_1422 (O_1422,N_9502,N_9833);
nor UO_1423 (O_1423,N_9777,N_9328);
and UO_1424 (O_1424,N_9028,N_9962);
nor UO_1425 (O_1425,N_9767,N_9542);
nand UO_1426 (O_1426,N_9145,N_9544);
and UO_1427 (O_1427,N_9426,N_9388);
or UO_1428 (O_1428,N_9940,N_9467);
and UO_1429 (O_1429,N_9468,N_9309);
nand UO_1430 (O_1430,N_9529,N_9522);
nand UO_1431 (O_1431,N_9875,N_9242);
and UO_1432 (O_1432,N_9085,N_9334);
nor UO_1433 (O_1433,N_9140,N_9830);
nand UO_1434 (O_1434,N_9475,N_9723);
or UO_1435 (O_1435,N_9893,N_9424);
nor UO_1436 (O_1436,N_9934,N_9766);
and UO_1437 (O_1437,N_9777,N_9248);
nand UO_1438 (O_1438,N_9274,N_9887);
nand UO_1439 (O_1439,N_9334,N_9351);
or UO_1440 (O_1440,N_9362,N_9759);
nand UO_1441 (O_1441,N_9663,N_9786);
and UO_1442 (O_1442,N_9071,N_9925);
nor UO_1443 (O_1443,N_9136,N_9596);
or UO_1444 (O_1444,N_9808,N_9631);
nand UO_1445 (O_1445,N_9051,N_9810);
and UO_1446 (O_1446,N_9591,N_9869);
nor UO_1447 (O_1447,N_9897,N_9013);
nor UO_1448 (O_1448,N_9859,N_9049);
nand UO_1449 (O_1449,N_9828,N_9783);
nand UO_1450 (O_1450,N_9738,N_9067);
nor UO_1451 (O_1451,N_9911,N_9927);
nand UO_1452 (O_1452,N_9144,N_9306);
and UO_1453 (O_1453,N_9082,N_9417);
or UO_1454 (O_1454,N_9736,N_9401);
or UO_1455 (O_1455,N_9421,N_9298);
or UO_1456 (O_1456,N_9934,N_9936);
or UO_1457 (O_1457,N_9470,N_9136);
nand UO_1458 (O_1458,N_9628,N_9330);
and UO_1459 (O_1459,N_9840,N_9450);
and UO_1460 (O_1460,N_9157,N_9658);
and UO_1461 (O_1461,N_9464,N_9941);
and UO_1462 (O_1462,N_9615,N_9303);
and UO_1463 (O_1463,N_9899,N_9494);
and UO_1464 (O_1464,N_9380,N_9160);
nor UO_1465 (O_1465,N_9040,N_9435);
nor UO_1466 (O_1466,N_9670,N_9942);
nand UO_1467 (O_1467,N_9004,N_9355);
or UO_1468 (O_1468,N_9049,N_9922);
nor UO_1469 (O_1469,N_9184,N_9858);
and UO_1470 (O_1470,N_9047,N_9898);
and UO_1471 (O_1471,N_9262,N_9597);
or UO_1472 (O_1472,N_9003,N_9028);
and UO_1473 (O_1473,N_9225,N_9932);
and UO_1474 (O_1474,N_9044,N_9784);
and UO_1475 (O_1475,N_9037,N_9106);
nor UO_1476 (O_1476,N_9459,N_9496);
nand UO_1477 (O_1477,N_9225,N_9566);
nand UO_1478 (O_1478,N_9428,N_9538);
or UO_1479 (O_1479,N_9268,N_9537);
and UO_1480 (O_1480,N_9531,N_9168);
or UO_1481 (O_1481,N_9610,N_9531);
and UO_1482 (O_1482,N_9372,N_9404);
nand UO_1483 (O_1483,N_9498,N_9793);
nor UO_1484 (O_1484,N_9543,N_9848);
or UO_1485 (O_1485,N_9936,N_9733);
nor UO_1486 (O_1486,N_9195,N_9892);
nor UO_1487 (O_1487,N_9401,N_9009);
and UO_1488 (O_1488,N_9115,N_9716);
nor UO_1489 (O_1489,N_9344,N_9581);
nor UO_1490 (O_1490,N_9803,N_9135);
nor UO_1491 (O_1491,N_9185,N_9495);
and UO_1492 (O_1492,N_9721,N_9834);
or UO_1493 (O_1493,N_9330,N_9068);
or UO_1494 (O_1494,N_9178,N_9960);
and UO_1495 (O_1495,N_9369,N_9122);
and UO_1496 (O_1496,N_9499,N_9959);
nand UO_1497 (O_1497,N_9599,N_9625);
nand UO_1498 (O_1498,N_9118,N_9006);
or UO_1499 (O_1499,N_9021,N_9922);
endmodule