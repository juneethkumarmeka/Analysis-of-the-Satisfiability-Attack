module basic_1500_15000_2000_3_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10028,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10043,N_10044,N_10045,N_10047,N_10048,N_10049,N_10051,N_10052,N_10053,N_10054,N_10056,N_10057,N_10058,N_10059,N_10061,N_10062,N_10063,N_10064,N_10065,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10075,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10086,N_10087,N_10089,N_10091,N_10092,N_10093,N_10094,N_10095,N_10097,N_10098,N_10099,N_10100,N_10101,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10111,N_10112,N_10113,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10143,N_10144,N_10146,N_10147,N_10148,N_10149,N_10151,N_10152,N_10153,N_10155,N_10156,N_10157,N_10158,N_10159,N_10161,N_10162,N_10163,N_10164,N_10166,N_10167,N_10168,N_10172,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10231,N_10232,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10241,N_10243,N_10244,N_10245,N_10246,N_10248,N_10249,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10278,N_10279,N_10280,N_10281,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10310,N_10312,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10322,N_10325,N_10326,N_10327,N_10328,N_10329,N_10332,N_10333,N_10334,N_10337,N_10338,N_10339,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10353,N_10354,N_10355,N_10357,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10367,N_10368,N_10369,N_10370,N_10373,N_10374,N_10375,N_10376,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10406,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10429,N_10430,N_10431,N_10433,N_10434,N_10438,N_10439,N_10440,N_10444,N_10445,N_10446,N_10448,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10505,N_10506,N_10507,N_10509,N_10510,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10529,N_10530,N_10531,N_10532,N_10534,N_10536,N_10537,N_10538,N_10539,N_10540,N_10543,N_10545,N_10546,N_10547,N_10548,N_10549,N_10551,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10562,N_10563,N_10564,N_10568,N_10570,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10597,N_10598,N_10600,N_10601,N_10602,N_10604,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10625,N_10626,N_10628,N_10629,N_10631,N_10632,N_10633,N_10635,N_10637,N_10639,N_10640,N_10641,N_10644,N_10646,N_10647,N_10648,N_10649,N_10650,N_10652,N_10653,N_10654,N_10655,N_10656,N_10658,N_10659,N_10660,N_10661,N_10664,N_10665,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10675,N_10676,N_10677,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10693,N_10694,N_10696,N_10697,N_10698,N_10699,N_10701,N_10702,N_10703,N_10704,N_10705,N_10707,N_10708,N_10710,N_10713,N_10715,N_10718,N_10719,N_10720,N_10726,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10736,N_10737,N_10738,N_10739,N_10740,N_10742,N_10745,N_10746,N_10747,N_10748,N_10749,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10767,N_10768,N_10769,N_10772,N_10773,N_10775,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10791,N_10792,N_10796,N_10797,N_10798,N_10799,N_10801,N_10802,N_10803,N_10804,N_10805,N_10807,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10838,N_10839,N_10841,N_10842,N_10843,N_10845,N_10846,N_10847,N_10848,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10865,N_10866,N_10869,N_10870,N_10875,N_10877,N_10878,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10889,N_10890,N_10891,N_10892,N_10894,N_10895,N_10897,N_10898,N_10899,N_10900,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10910,N_10912,N_10913,N_10914,N_10915,N_10916,N_10919,N_10920,N_10921,N_10924,N_10926,N_10927,N_10928,N_10930,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10952,N_10953,N_10954,N_10957,N_10958,N_10960,N_10962,N_10964,N_10966,N_10967,N_10969,N_10970,N_10971,N_10972,N_10973,N_10975,N_10977,N_10978,N_10980,N_10981,N_10982,N_10983,N_10986,N_10988,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11015,N_11016,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11026,N_11027,N_11029,N_11030,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11040,N_11041,N_11042,N_11043,N_11044,N_11046,N_11047,N_11048,N_11049,N_11051,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11066,N_11067,N_11069,N_11070,N_11071,N_11073,N_11075,N_11076,N_11077,N_11079,N_11080,N_11082,N_11083,N_11084,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11093,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11102,N_11103,N_11105,N_11107,N_11109,N_11110,N_11111,N_11112,N_11113,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11124,N_11125,N_11126,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11146,N_11147,N_11148,N_11150,N_11151,N_11152,N_11153,N_11154,N_11156,N_11157,N_11158,N_11159,N_11161,N_11162,N_11165,N_11166,N_11167,N_11168,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11200,N_11201,N_11205,N_11206,N_11207,N_11208,N_11209,N_11212,N_11214,N_11215,N_11216,N_11218,N_11219,N_11220,N_11222,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11243,N_11244,N_11246,N_11247,N_11248,N_11250,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11259,N_11265,N_11266,N_11267,N_11269,N_11270,N_11271,N_11274,N_11275,N_11277,N_11278,N_11279,N_11281,N_11282,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11309,N_11310,N_11312,N_11313,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11328,N_11329,N_11330,N_11331,N_11332,N_11337,N_11338,N_11339,N_11340,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11366,N_11368,N_11370,N_11371,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11382,N_11383,N_11384,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11397,N_11398,N_11399,N_11401,N_11402,N_11403,N_11404,N_11406,N_11407,N_11408,N_11409,N_11412,N_11414,N_11415,N_11416,N_11417,N_11418,N_11420,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11430,N_11433,N_11434,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11446,N_11448,N_11449,N_11450,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11487,N_11489,N_11490,N_11491,N_11492,N_11493,N_11495,N_11498,N_11499,N_11500,N_11502,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11517,N_11518,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11529,N_11530,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11543,N_11544,N_11547,N_11548,N_11549,N_11550,N_11551,N_11553,N_11554,N_11557,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11575,N_11576,N_11577,N_11578,N_11579,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11599,N_11601,N_11602,N_11603,N_11605,N_11606,N_11607,N_11608,N_11610,N_11613,N_11615,N_11616,N_11618,N_11619,N_11620,N_11622,N_11623,N_11625,N_11627,N_11629,N_11630,N_11631,N_11632,N_11634,N_11637,N_11638,N_11639,N_11640,N_11642,N_11643,N_11644,N_11645,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11663,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11682,N_11683,N_11687,N_11688,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11704,N_11705,N_11706,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11718,N_11719,N_11721,N_11722,N_11723,N_11724,N_11726,N_11727,N_11728,N_11730,N_11731,N_11732,N_11733,N_11736,N_11737,N_11738,N_11739,N_11740,N_11742,N_11744,N_11745,N_11746,N_11747,N_11748,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11761,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11784,N_11785,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11825,N_11826,N_11828,N_11830,N_11831,N_11832,N_11833,N_11834,N_11836,N_11837,N_11839,N_11840,N_11841,N_11843,N_11844,N_11846,N_11847,N_11848,N_11850,N_11851,N_11852,N_11854,N_11855,N_11856,N_11857,N_11859,N_11862,N_11863,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11872,N_11873,N_11874,N_11876,N_11877,N_11878,N_11879,N_11880,N_11882,N_11883,N_11884,N_11885,N_11887,N_11888,N_11889,N_11891,N_11892,N_11893,N_11894,N_11895,N_11897,N_11898,N_11899,N_11900,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11912,N_11913,N_11915,N_11916,N_11917,N_11919,N_11920,N_11921,N_11922,N_11924,N_11926,N_11927,N_11929,N_11930,N_11931,N_11932,N_11933,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11950,N_11953,N_11954,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11972,N_11974,N_11975,N_11976,N_11977,N_11978,N_11980,N_11981,N_11982,N_11984,N_11985,N_11986,N_11987,N_11989,N_11990,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_12000,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12010,N_12012,N_12013,N_12014,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12047,N_12048,N_12050,N_12051,N_12052,N_12054,N_12055,N_12056,N_12057,N_12058,N_12060,N_12061,N_12062,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12071,N_12072,N_12073,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12104,N_12105,N_12106,N_12107,N_12108,N_12110,N_12111,N_12112,N_12113,N_12115,N_12118,N_12119,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12134,N_12135,N_12136,N_12137,N_12138,N_12140,N_12141,N_12142,N_12145,N_12146,N_12147,N_12148,N_12150,N_12151,N_12153,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12162,N_12163,N_12164,N_12165,N_12166,N_12168,N_12169,N_12170,N_12172,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12185,N_12187,N_12189,N_12190,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12212,N_12213,N_12214,N_12216,N_12218,N_12219,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12233,N_12234,N_12235,N_12236,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12245,N_12246,N_12248,N_12249,N_12252,N_12254,N_12255,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12269,N_12270,N_12271,N_12272,N_12273,N_12275,N_12276,N_12277,N_12278,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12300,N_12301,N_12303,N_12304,N_12306,N_12307,N_12308,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12322,N_12323,N_12324,N_12325,N_12326,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12339,N_12340,N_12341,N_12343,N_12344,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12366,N_12367,N_12368,N_12369,N_12371,N_12372,N_12373,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12388,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12402,N_12405,N_12406,N_12407,N_12408,N_12409,N_12411,N_12412,N_12413,N_12414,N_12416,N_12417,N_12418,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12441,N_12442,N_12445,N_12446,N_12447,N_12448,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12457,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12466,N_12467,N_12468,N_12469,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12493,N_12494,N_12495,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12515,N_12516,N_12517,N_12518,N_12519,N_12521,N_12522,N_12524,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12570,N_12571,N_12572,N_12573,N_12574,N_12576,N_12577,N_12578,N_12579,N_12580,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12595,N_12596,N_12597,N_12599,N_12600,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12609,N_12610,N_12611,N_12612,N_12614,N_12616,N_12617,N_12618,N_12619,N_12621,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12632,N_12633,N_12634,N_12635,N_12636,N_12638,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12658,N_12659,N_12662,N_12663,N_12664,N_12666,N_12667,N_12668,N_12669,N_12671,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12690,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12700,N_12701,N_12702,N_12703,N_12704,N_12706,N_12707,N_12708,N_12710,N_12711,N_12712,N_12713,N_12714,N_12716,N_12717,N_12719,N_12720,N_12721,N_12722,N_12723,N_12725,N_12726,N_12727,N_12728,N_12729,N_12731,N_12732,N_12733,N_12734,N_12735,N_12737,N_12738,N_12739,N_12741,N_12742,N_12743,N_12744,N_12745,N_12749,N_12750,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12771,N_12772,N_12773,N_12774,N_12775,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12791,N_12793,N_12795,N_12796,N_12798,N_12800,N_12801,N_12803,N_12805,N_12806,N_12807,N_12809,N_12810,N_12812,N_12814,N_12815,N_12817,N_12819,N_12820,N_12822,N_12823,N_12824,N_12826,N_12827,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12853,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12864,N_12865,N_12866,N_12869,N_12870,N_12871,N_12872,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12888,N_12890,N_12891,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12906,N_12907,N_12909,N_12910,N_12911,N_12912,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12943,N_12945,N_12946,N_12947,N_12948,N_12950,N_12951,N_12953,N_12954,N_12955,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12985,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13008,N_13009,N_13010,N_13011,N_13012,N_13014,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13023,N_13024,N_13025,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13043,N_13044,N_13045,N_13046,N_13047,N_13049,N_13050,N_13051,N_13052,N_13054,N_13057,N_13058,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13068,N_13069,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13083,N_13084,N_13085,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13101,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13118,N_13119,N_13123,N_13124,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13144,N_13145,N_13146,N_13147,N_13148,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13177,N_13178,N_13179,N_13180,N_13181,N_13183,N_13184,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13205,N_13206,N_13207,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13219,N_13221,N_13222,N_13223,N_13224,N_13225,N_13227,N_13228,N_13229,N_13230,N_13231,N_13233,N_13234,N_13235,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13247,N_13249,N_13250,N_13251,N_13252,N_13253,N_13255,N_13256,N_13257,N_13258,N_13259,N_13261,N_13262,N_13263,N_13264,N_13265,N_13267,N_13268,N_13269,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13332,N_13333,N_13334,N_13336,N_13337,N_13338,N_13339,N_13340,N_13342,N_13343,N_13344,N_13345,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13367,N_13368,N_13369,N_13371,N_13372,N_13373,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13382,N_13383,N_13384,N_13385,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13396,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13406,N_13407,N_13409,N_13411,N_13412,N_13413,N_13414,N_13415,N_13417,N_13418,N_13419,N_13420,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13440,N_13441,N_13444,N_13445,N_13446,N_13448,N_13449,N_13450,N_13452,N_13453,N_13454,N_13455,N_13456,N_13458,N_13459,N_13460,N_13461,N_13462,N_13465,N_13466,N_13467,N_13468,N_13469,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13485,N_13486,N_13487,N_13488,N_13489,N_13492,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13504,N_13505,N_13506,N_13507,N_13508,N_13511,N_13512,N_13513,N_13514,N_13515,N_13517,N_13518,N_13519,N_13521,N_13522,N_13523,N_13524,N_13525,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13563,N_13565,N_13566,N_13567,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13578,N_13579,N_13580,N_13581,N_13582,N_13584,N_13585,N_13586,N_13588,N_13589,N_13590,N_13591,N_13592,N_13594,N_13595,N_13596,N_13597,N_13598,N_13600,N_13601,N_13603,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13618,N_13619,N_13621,N_13622,N_13623,N_13624,N_13625,N_13627,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13640,N_13641,N_13642,N_13643,N_13645,N_13646,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13665,N_13667,N_13668,N_13669,N_13670,N_13671,N_13673,N_13674,N_13675,N_13677,N_13678,N_13679,N_13681,N_13682,N_13683,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13704,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13724,N_13725,N_13726,N_13727,N_13729,N_13730,N_13731,N_13732,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13741,N_13742,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13751,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13775,N_13776,N_13777,N_13778,N_13779,N_13781,N_13782,N_13784,N_13787,N_13788,N_13789,N_13790,N_13795,N_13797,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13833,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13873,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13884,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13902,N_13903,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13938,N_13941,N_13944,N_13945,N_13946,N_13948,N_13949,N_13951,N_13952,N_13953,N_13954,N_13955,N_13957,N_13958,N_13959,N_13960,N_13961,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13975,N_13976,N_13979,N_13980,N_13981,N_13983,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13997,N_13998,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14037,N_14038,N_14039,N_14041,N_14042,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14053,N_14054,N_14055,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14084,N_14085,N_14087,N_14088,N_14089,N_14091,N_14092,N_14093,N_14094,N_14095,N_14097,N_14098,N_14099,N_14100,N_14102,N_14104,N_14105,N_14106,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14122,N_14123,N_14124,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14134,N_14135,N_14137,N_14138,N_14139,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14152,N_14153,N_14154,N_14156,N_14158,N_14159,N_14160,N_14162,N_14163,N_14165,N_14167,N_14168,N_14169,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14190,N_14191,N_14192,N_14193,N_14194,N_14196,N_14197,N_14198,N_14199,N_14202,N_14203,N_14204,N_14205,N_14206,N_14208,N_14209,N_14212,N_14214,N_14215,N_14216,N_14217,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14229,N_14231,N_14232,N_14234,N_14235,N_14236,N_14237,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14264,N_14265,N_14266,N_14267,N_14268,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14297,N_14298,N_14299,N_14300,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14319,N_14320,N_14322,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14340,N_14342,N_14344,N_14345,N_14346,N_14348,N_14350,N_14351,N_14352,N_14353,N_14355,N_14356,N_14357,N_14358,N_14360,N_14361,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14375,N_14378,N_14379,N_14380,N_14382,N_14383,N_14384,N_14385,N_14387,N_14388,N_14389,N_14390,N_14392,N_14394,N_14395,N_14396,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14408,N_14409,N_14410,N_14411,N_14415,N_14417,N_14418,N_14420,N_14421,N_14422,N_14424,N_14425,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14435,N_14436,N_14437,N_14438,N_14440,N_14441,N_14442,N_14443,N_14444,N_14446,N_14447,N_14448,N_14449,N_14450,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14475,N_14477,N_14478,N_14479,N_14480,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14490,N_14491,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14505,N_14506,N_14507,N_14508,N_14510,N_14511,N_14512,N_14514,N_14515,N_14516,N_14518,N_14519,N_14520,N_14521,N_14523,N_14524,N_14527,N_14528,N_14529,N_14531,N_14532,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14544,N_14545,N_14546,N_14547,N_14549,N_14550,N_14551,N_14552,N_14555,N_14557,N_14558,N_14560,N_14561,N_14562,N_14563,N_14564,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14580,N_14581,N_14582,N_14583,N_14585,N_14586,N_14587,N_14588,N_14590,N_14591,N_14592,N_14593,N_14594,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14604,N_14606,N_14608,N_14612,N_14614,N_14615,N_14616,N_14617,N_14619,N_14620,N_14622,N_14623,N_14624,N_14625,N_14627,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14640,N_14641,N_14642,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14661,N_14662,N_14663,N_14664,N_14665,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14697,N_14698,N_14699,N_14701,N_14702,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14723,N_14725,N_14726,N_14727,N_14728,N_14730,N_14731,N_14732,N_14736,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14746,N_14747,N_14748,N_14749,N_14750,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14763,N_14764,N_14766,N_14767,N_14768,N_14769,N_14771,N_14772,N_14774,N_14775,N_14776,N_14777,N_14778,N_14780,N_14781,N_14784,N_14785,N_14786,N_14787,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14800,N_14802,N_14803,N_14804,N_14805,N_14807,N_14808,N_14810,N_14812,N_14813,N_14814,N_14815,N_14817,N_14818,N_14819,N_14820,N_14822,N_14823,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14859,N_14860,N_14861,N_14862,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14889,N_14893,N_14894,N_14895,N_14896,N_14897,N_14899,N_14900,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14915,N_14917,N_14918,N_14919,N_14920,N_14922,N_14923,N_14924,N_14925,N_14927,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14941,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14963,N_14966,N_14967,N_14968,N_14970,N_14971,N_14972,N_14973,N_14974,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14987,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14998,N_14999;
nand U0 (N_0,In_368,In_1299);
and U1 (N_1,In_1472,In_1195);
and U2 (N_2,In_881,In_1263);
nand U3 (N_3,In_596,In_450);
nor U4 (N_4,In_411,In_696);
nor U5 (N_5,In_901,In_11);
nand U6 (N_6,In_962,In_331);
or U7 (N_7,In_367,In_8);
or U8 (N_8,In_1421,In_1175);
and U9 (N_9,In_1016,In_258);
or U10 (N_10,In_1058,In_268);
or U11 (N_11,In_1145,In_1433);
nor U12 (N_12,In_888,In_1193);
nor U13 (N_13,In_657,In_92);
or U14 (N_14,In_146,In_666);
nor U15 (N_15,In_417,In_1300);
nand U16 (N_16,In_366,In_1325);
nand U17 (N_17,In_727,In_987);
or U18 (N_18,In_1252,In_1108);
nor U19 (N_19,In_694,In_446);
and U20 (N_20,In_336,In_909);
nor U21 (N_21,In_734,In_209);
or U22 (N_22,In_1120,In_1114);
or U23 (N_23,In_916,In_170);
and U24 (N_24,In_1345,In_489);
and U25 (N_25,In_354,In_976);
nor U26 (N_26,In_830,In_798);
and U27 (N_27,In_862,In_461);
and U28 (N_28,In_1453,In_1071);
or U29 (N_29,In_1329,In_1042);
nand U30 (N_30,In_244,In_444);
nand U31 (N_31,In_1467,In_374);
and U32 (N_32,In_608,In_826);
and U33 (N_33,In_1021,In_555);
and U34 (N_34,In_751,In_955);
nor U35 (N_35,In_676,In_1069);
and U36 (N_36,In_186,In_1428);
nor U37 (N_37,In_169,In_409);
nand U38 (N_38,In_514,In_31);
nor U39 (N_39,In_451,In_587);
or U40 (N_40,In_1171,In_1064);
or U41 (N_41,In_398,In_853);
and U42 (N_42,In_564,In_590);
or U43 (N_43,In_669,In_150);
or U44 (N_44,In_757,In_262);
nand U45 (N_45,In_1310,In_1356);
nor U46 (N_46,In_742,In_1457);
and U47 (N_47,In_57,In_800);
or U48 (N_48,In_1386,In_1471);
nor U49 (N_49,In_245,In_1400);
nor U50 (N_50,In_20,In_1311);
and U51 (N_51,In_414,In_545);
or U52 (N_52,In_1292,In_12);
nor U53 (N_53,In_377,In_1103);
xor U54 (N_54,In_869,In_1125);
and U55 (N_55,In_852,In_740);
and U56 (N_56,In_323,In_988);
nand U57 (N_57,In_1167,In_726);
or U58 (N_58,In_22,In_598);
nor U59 (N_59,In_519,In_36);
and U60 (N_60,In_1346,In_1331);
or U61 (N_61,In_548,In_282);
nand U62 (N_62,In_54,In_1146);
nor U63 (N_63,In_343,In_206);
and U64 (N_64,In_148,In_1289);
and U65 (N_65,In_176,In_1404);
nor U66 (N_66,In_375,In_1025);
and U67 (N_67,In_860,In_1131);
nand U68 (N_68,In_878,In_194);
and U69 (N_69,In_369,In_765);
or U70 (N_70,In_1051,In_1391);
nor U71 (N_71,In_920,In_455);
or U72 (N_72,In_307,In_229);
or U73 (N_73,In_1054,In_153);
nand U74 (N_74,In_1451,In_1220);
or U75 (N_75,In_132,In_15);
nand U76 (N_76,In_1455,In_1168);
nor U77 (N_77,In_864,In_953);
nor U78 (N_78,In_359,In_149);
nor U79 (N_79,In_609,In_1026);
nand U80 (N_80,In_1281,In_661);
and U81 (N_81,In_944,In_567);
nor U82 (N_82,In_168,In_9);
or U83 (N_83,In_1319,In_1340);
nand U84 (N_84,In_356,In_1199);
nand U85 (N_85,In_554,In_958);
nand U86 (N_86,In_1095,In_139);
and U87 (N_87,In_213,In_1094);
nand U88 (N_88,In_810,In_982);
nand U89 (N_89,In_1041,In_1437);
or U90 (N_90,In_775,In_321);
or U91 (N_91,In_113,In_741);
and U92 (N_92,In_175,In_328);
or U93 (N_93,In_314,In_882);
nor U94 (N_94,In_1154,In_685);
nor U95 (N_95,In_755,In_479);
nand U96 (N_96,In_1466,In_1138);
nand U97 (N_97,In_1242,In_349);
and U98 (N_98,In_1362,In_951);
nor U99 (N_99,In_1334,In_1382);
nand U100 (N_100,In_1302,In_1275);
xor U101 (N_101,In_612,In_1491);
or U102 (N_102,In_611,In_434);
or U103 (N_103,In_1269,In_1012);
or U104 (N_104,In_14,In_1076);
or U105 (N_105,In_752,In_1218);
nand U106 (N_106,In_884,In_309);
or U107 (N_107,In_64,In_88);
or U108 (N_108,In_797,In_140);
nand U109 (N_109,In_185,In_838);
or U110 (N_110,In_575,In_1248);
nand U111 (N_111,In_68,In_265);
nand U112 (N_112,In_412,In_805);
nor U113 (N_113,In_906,In_1232);
or U114 (N_114,In_501,In_698);
nand U115 (N_115,In_1082,In_1412);
nor U116 (N_116,In_957,In_943);
xnor U117 (N_117,In_1383,In_678);
and U118 (N_118,In_541,In_1436);
nor U119 (N_119,In_561,In_753);
and U120 (N_120,In_1009,In_792);
nand U121 (N_121,In_303,In_342);
and U122 (N_122,In_1407,In_457);
nor U123 (N_123,In_1169,In_254);
nand U124 (N_124,In_941,In_983);
nor U125 (N_125,In_680,In_115);
or U126 (N_126,In_815,In_1372);
nand U127 (N_127,In_527,In_1161);
nand U128 (N_128,In_1489,In_1014);
nand U129 (N_129,In_263,In_344);
or U130 (N_130,In_1185,In_1264);
and U131 (N_131,In_1036,In_423);
or U132 (N_132,In_106,In_538);
and U133 (N_133,In_580,In_1483);
or U134 (N_134,In_225,In_1461);
or U135 (N_135,In_723,In_513);
nor U136 (N_136,In_1124,In_191);
nor U137 (N_137,In_1115,In_1398);
or U138 (N_138,In_1477,In_19);
or U139 (N_139,In_719,In_1074);
or U140 (N_140,In_189,In_78);
nor U141 (N_141,In_380,In_159);
or U142 (N_142,In_310,In_1011);
xor U143 (N_143,In_1271,In_438);
or U144 (N_144,In_890,In_1367);
nor U145 (N_145,In_854,In_1376);
nand U146 (N_146,In_870,In_529);
nand U147 (N_147,In_280,In_136);
or U148 (N_148,In_1484,In_100);
or U149 (N_149,In_1177,In_634);
or U150 (N_150,In_134,In_1142);
and U151 (N_151,In_181,In_682);
and U152 (N_152,In_493,In_103);
nor U153 (N_153,In_537,In_1465);
xnor U154 (N_154,In_949,In_56);
and U155 (N_155,In_362,In_326);
and U156 (N_156,In_327,In_840);
nand U157 (N_157,In_706,In_1452);
nand U158 (N_158,In_404,In_565);
nand U159 (N_159,In_77,In_468);
nor U160 (N_160,In_1239,In_295);
or U161 (N_161,In_1005,In_872);
and U162 (N_162,In_1134,In_264);
or U163 (N_163,In_37,In_745);
and U164 (N_164,In_1401,In_1265);
and U165 (N_165,In_614,In_316);
or U166 (N_166,In_464,In_760);
nor U167 (N_167,In_1364,In_87);
nand U168 (N_168,In_1022,In_10);
nor U169 (N_169,In_668,In_621);
and U170 (N_170,In_602,In_251);
or U171 (N_171,In_27,In_399);
nor U172 (N_172,In_1377,In_702);
nor U173 (N_173,In_663,In_298);
or U174 (N_174,In_764,In_892);
nor U175 (N_175,In_533,In_1308);
or U176 (N_176,In_1415,In_1130);
nand U177 (N_177,In_17,In_562);
or U178 (N_178,In_63,In_686);
nor U179 (N_179,In_849,In_595);
and U180 (N_180,In_93,In_273);
or U181 (N_181,In_1083,In_281);
nand U182 (N_182,In_214,In_1090);
or U183 (N_183,In_1221,In_467);
or U184 (N_184,In_1055,In_114);
or U185 (N_185,In_341,In_794);
nor U186 (N_186,In_492,In_1040);
or U187 (N_187,In_1222,In_1203);
or U188 (N_188,In_712,In_420);
or U189 (N_189,In_248,In_837);
or U190 (N_190,In_144,In_233);
nand U191 (N_191,In_137,In_1183);
or U192 (N_192,In_1062,In_154);
and U193 (N_193,In_1053,In_692);
and U194 (N_194,In_659,In_459);
or U195 (N_195,In_845,In_488);
nor U196 (N_196,In_1430,In_1347);
and U197 (N_197,In_121,In_728);
and U198 (N_198,In_230,In_1385);
nand U199 (N_199,In_203,In_453);
nor U200 (N_200,In_53,In_118);
nand U201 (N_201,In_439,In_346);
nor U202 (N_202,In_672,In_689);
nand U203 (N_203,In_900,In_60);
and U204 (N_204,In_816,In_1318);
nor U205 (N_205,In_131,In_629);
nor U206 (N_206,In_1337,In_709);
or U207 (N_207,In_861,In_44);
and U208 (N_208,In_631,In_1313);
nand U209 (N_209,In_1333,In_526);
and U210 (N_210,In_543,In_610);
nor U211 (N_211,In_1384,In_990);
nand U212 (N_212,In_572,In_517);
and U213 (N_213,In_1282,In_644);
or U214 (N_214,In_828,In_831);
and U215 (N_215,In_142,In_774);
or U216 (N_216,In_1482,In_939);
nand U217 (N_217,In_556,In_1335);
or U218 (N_218,In_600,In_1112);
nand U219 (N_219,In_1342,In_1093);
nand U220 (N_220,In_41,In_656);
or U221 (N_221,In_1240,In_1078);
and U222 (N_222,In_1170,In_1411);
or U223 (N_223,In_94,In_454);
and U224 (N_224,In_1439,In_1245);
and U225 (N_225,In_211,In_445);
nand U226 (N_226,In_748,In_277);
or U227 (N_227,In_559,In_242);
or U228 (N_228,In_851,In_524);
nor U229 (N_229,In_2,In_337);
nand U230 (N_230,In_866,In_1044);
nand U231 (N_231,In_1061,In_355);
and U232 (N_232,In_1419,In_1119);
nand U233 (N_233,In_1314,In_1387);
nand U234 (N_234,In_1268,In_972);
nor U235 (N_235,In_832,In_1460);
and U236 (N_236,In_437,In_822);
or U237 (N_237,In_1226,In_880);
nand U238 (N_238,In_95,In_1438);
and U239 (N_239,In_827,In_911);
or U240 (N_240,In_1309,In_950);
xnor U241 (N_241,In_675,In_1293);
and U242 (N_242,In_1420,In_397);
and U243 (N_243,In_835,In_440);
and U244 (N_244,In_592,In_141);
or U245 (N_245,In_531,In_642);
nor U246 (N_246,In_758,In_490);
nand U247 (N_247,In_1068,In_690);
and U248 (N_248,In_1374,In_569);
or U249 (N_249,In_253,In_491);
nand U250 (N_250,In_246,In_138);
and U251 (N_251,In_604,In_583);
nand U252 (N_252,In_1323,In_1075);
and U253 (N_253,In_704,In_1086);
xor U254 (N_254,In_782,In_681);
or U255 (N_255,In_1139,In_918);
xnor U256 (N_256,In_744,In_30);
nor U257 (N_257,In_97,In_516);
nand U258 (N_258,In_1305,In_1250);
nor U259 (N_259,In_945,In_58);
and U260 (N_260,In_160,In_495);
nand U261 (N_261,In_735,In_46);
or U262 (N_262,In_407,In_234);
and U263 (N_263,In_802,In_883);
and U264 (N_264,In_166,In_59);
nand U265 (N_265,In_301,In_1454);
nor U266 (N_266,In_979,In_868);
and U267 (N_267,In_1135,In_535);
nand U268 (N_268,In_1351,In_895);
or U269 (N_269,In_410,In_578);
nor U270 (N_270,In_499,In_980);
nor U271 (N_271,In_504,In_266);
and U272 (N_272,In_549,In_1180);
nor U273 (N_273,In_1380,In_750);
nor U274 (N_274,In_429,In_1288);
and U275 (N_275,In_904,In_430);
nand U276 (N_276,In_197,In_640);
or U277 (N_277,In_1246,In_776);
and U278 (N_278,In_550,In_1088);
or U279 (N_279,In_799,In_353);
or U280 (N_280,In_222,In_1072);
and U281 (N_281,In_1298,In_617);
or U282 (N_282,In_1444,In_844);
nand U283 (N_283,In_620,In_974);
nand U284 (N_284,In_730,In_1096);
and U285 (N_285,In_1033,In_238);
nand U286 (N_286,In_985,In_174);
nand U287 (N_287,In_1262,In_171);
or U288 (N_288,In_391,In_1225);
nor U289 (N_289,In_1441,In_848);
xor U290 (N_290,In_385,In_1432);
or U291 (N_291,In_452,In_469);
and U292 (N_292,In_1190,In_584);
or U293 (N_293,In_806,In_542);
nand U294 (N_294,In_319,In_127);
nor U295 (N_295,In_585,In_1092);
or U296 (N_296,In_302,In_956);
xor U297 (N_297,In_1105,In_485);
nand U298 (N_298,In_1067,In_571);
nor U299 (N_299,In_563,In_111);
nand U300 (N_300,In_1132,In_1089);
or U301 (N_301,In_279,In_789);
nor U302 (N_302,In_903,In_219);
nor U303 (N_303,In_915,In_1098);
nand U304 (N_304,In_1000,In_227);
or U305 (N_305,In_35,In_294);
or U306 (N_306,In_1402,In_787);
nand U307 (N_307,In_1109,In_352);
nor U308 (N_308,In_967,In_4);
nand U309 (N_309,In_732,In_306);
nor U310 (N_310,In_1279,In_102);
nand U311 (N_311,In_418,In_1081);
nand U312 (N_312,In_1417,In_403);
nand U313 (N_313,In_922,In_259);
nand U314 (N_314,In_347,In_1297);
and U315 (N_315,In_660,In_812);
nor U316 (N_316,In_162,In_632);
nand U317 (N_317,In_1390,In_1409);
and U318 (N_318,In_52,In_66);
and U319 (N_319,In_196,In_76);
and U320 (N_320,In_885,In_975);
xnor U321 (N_321,In_547,In_643);
xnor U322 (N_322,In_1456,In_978);
nand U323 (N_323,In_893,In_551);
nand U324 (N_324,In_345,In_1446);
nor U325 (N_325,In_670,In_1215);
and U326 (N_326,In_923,In_215);
nand U327 (N_327,In_1003,In_1247);
nor U328 (N_328,In_729,In_1429);
and U329 (N_329,In_593,In_1328);
and U330 (N_330,In_1237,In_1179);
and U331 (N_331,In_599,In_1206);
nand U332 (N_332,In_158,In_338);
or U333 (N_333,In_1148,In_190);
and U334 (N_334,In_473,In_803);
nand U335 (N_335,In_993,In_299);
nand U336 (N_336,In_536,In_766);
or U337 (N_337,In_581,In_465);
and U338 (N_338,In_528,In_1326);
nor U339 (N_339,In_981,In_1201);
nor U340 (N_340,In_1307,In_1200);
and U341 (N_341,In_151,In_1060);
nand U342 (N_342,In_574,In_1359);
nand U343 (N_343,In_261,In_708);
or U344 (N_344,In_21,In_636);
or U345 (N_345,In_715,In_13);
nand U346 (N_346,In_1316,In_220);
or U347 (N_347,In_164,In_1235);
and U348 (N_348,In_1272,In_223);
or U349 (N_349,In_395,In_1143);
nand U350 (N_350,In_1371,In_769);
and U351 (N_351,In_1306,In_520);
or U352 (N_352,In_98,In_873);
nor U353 (N_353,In_684,In_1283);
nor U354 (N_354,In_267,In_24);
and U355 (N_355,In_809,In_1207);
nand U356 (N_356,In_1488,In_616);
nor U357 (N_357,In_1178,In_1123);
nand U358 (N_358,In_1233,In_921);
nand U359 (N_359,In_255,In_436);
nor U360 (N_360,In_655,In_201);
nand U361 (N_361,In_879,In_1485);
and U362 (N_362,In_784,In_1211);
and U363 (N_363,In_503,In_829);
and U364 (N_364,In_699,In_927);
nor U365 (N_365,In_1181,In_458);
nand U366 (N_366,In_272,In_557);
nand U367 (N_367,In_147,In_322);
and U368 (N_368,In_1370,In_311);
or U369 (N_369,In_1274,In_725);
or U370 (N_370,In_1286,In_1153);
or U371 (N_371,In_1015,In_433);
nand U372 (N_372,In_721,In_521);
nor U373 (N_373,In_204,In_867);
and U374 (N_374,In_930,In_496);
nor U375 (N_375,In_1449,In_304);
or U376 (N_376,In_1295,In_1365);
nor U377 (N_377,In_701,In_731);
xnor U378 (N_378,In_217,In_188);
nand U379 (N_379,In_475,In_472);
or U380 (N_380,In_363,In_773);
nand U381 (N_381,In_615,In_746);
nand U382 (N_382,In_1107,In_1353);
and U383 (N_383,In_308,In_713);
nor U384 (N_384,In_441,In_416);
nor U385 (N_385,In_252,In_449);
nand U386 (N_386,In_1192,In_662);
and U387 (N_387,In_257,In_406);
nand U388 (N_388,In_388,In_1373);
and U389 (N_389,In_105,In_202);
nand U390 (N_390,In_1118,In_1017);
nor U391 (N_391,In_1378,In_325);
and U392 (N_392,In_540,In_633);
nor U393 (N_393,In_163,In_591);
nor U394 (N_394,In_1358,In_839);
and U395 (N_395,In_1254,In_84);
nor U396 (N_396,In_928,In_618);
nor U397 (N_397,In_959,In_130);
or U398 (N_398,In_874,In_1128);
or U399 (N_399,In_1410,In_460);
nor U400 (N_400,In_498,In_560);
or U401 (N_401,In_435,In_1251);
nand U402 (N_402,In_1037,In_1198);
nor U403 (N_403,In_899,In_1341);
or U404 (N_404,In_332,In_1445);
nor U405 (N_405,In_534,In_51);
nor U406 (N_406,In_249,In_1487);
nand U407 (N_407,In_1270,In_40);
or U408 (N_408,In_525,In_819);
nor U409 (N_409,In_796,In_1209);
nand U410 (N_410,In_378,In_350);
xnor U411 (N_411,In_484,In_221);
and U412 (N_412,In_1234,In_1219);
nand U413 (N_413,In_365,In_296);
and U414 (N_414,In_964,In_47);
nor U415 (N_415,In_754,In_1052);
and U416 (N_416,In_80,In_90);
nand U417 (N_417,In_929,In_108);
and U418 (N_418,In_711,In_320);
nand U419 (N_419,In_1322,In_70);
nand U420 (N_420,In_1375,In_1097);
nand U421 (N_421,In_200,In_863);
or U422 (N_422,In_952,In_891);
nor U423 (N_423,In_1266,In_339);
nor U424 (N_424,In_1186,In_1324);
or U425 (N_425,In_278,In_1008);
nand U426 (N_426,In_691,In_518);
nor U427 (N_427,In_318,In_335);
or U428 (N_428,In_392,In_700);
nor U429 (N_429,In_1238,In_481);
nand U430 (N_430,In_447,In_371);
or U431 (N_431,In_1202,In_625);
and U432 (N_432,In_1137,In_99);
and U433 (N_433,In_1413,In_1013);
or U434 (N_434,In_1227,In_487);
nor U435 (N_435,In_3,In_1480);
and U436 (N_436,In_61,In_961);
nand U437 (N_437,In_419,In_413);
or U438 (N_438,In_733,In_50);
or U439 (N_439,In_156,In_1468);
and U440 (N_440,In_271,In_476);
and U441 (N_441,In_442,In_79);
nand U442 (N_442,In_207,In_333);
nor U443 (N_443,In_1006,In_530);
nand U444 (N_444,In_954,In_167);
and U445 (N_445,In_1057,In_767);
and U446 (N_446,In_135,In_1073);
nand U447 (N_447,In_897,In_522);
or U448 (N_448,In_783,In_1427);
nor U449 (N_449,In_1287,In_1267);
and U450 (N_450,In_1194,In_1164);
nor U451 (N_451,In_1448,In_1213);
xor U452 (N_452,In_348,In_817);
and U453 (N_453,In_814,In_1059);
and U454 (N_454,In_1163,In_788);
or U455 (N_455,In_850,In_428);
or U456 (N_456,In_208,In_1414);
nor U457 (N_457,In_1047,In_1406);
or U458 (N_458,In_924,In_1197);
or U459 (N_459,In_86,In_1027);
nand U460 (N_460,In_1490,In_1043);
nor U461 (N_461,In_1160,In_358);
and U462 (N_462,In_177,In_1223);
and U463 (N_463,In_1244,In_432);
or U464 (N_464,In_1001,In_902);
nand U465 (N_465,In_107,In_1050);
nand U466 (N_466,In_821,In_558);
and U467 (N_467,In_269,In_737);
nand U468 (N_468,In_1129,In_500);
nand U469 (N_469,In_693,In_1379);
nor U470 (N_470,In_855,In_1034);
nor U471 (N_471,In_422,In_183);
nand U472 (N_472,In_1478,In_566);
or U473 (N_473,In_771,In_1110);
nand U474 (N_474,In_1399,In_1277);
or U475 (N_475,In_973,In_101);
nor U476 (N_476,In_1361,In_421);
or U477 (N_477,In_67,In_651);
nor U478 (N_478,In_1049,In_1315);
nand U479 (N_479,In_372,In_184);
nand U480 (N_480,In_456,In_1204);
and U481 (N_481,In_1162,In_749);
or U482 (N_482,In_1470,In_576);
and U483 (N_483,In_1273,In_72);
nand U484 (N_484,In_589,In_770);
or U485 (N_485,In_544,In_1463);
nor U486 (N_486,In_415,In_931);
and U487 (N_487,In_486,In_568);
nand U488 (N_488,In_334,In_1352);
and U489 (N_489,In_23,In_842);
nand U490 (N_490,In_586,In_1228);
and U491 (N_491,In_739,In_934);
and U492 (N_492,In_224,In_1394);
nor U493 (N_493,In_478,In_1156);
and U494 (N_494,In_1187,In_29);
nor U495 (N_495,In_1366,In_1462);
nor U496 (N_496,In_626,In_989);
xnor U497 (N_497,In_1320,In_619);
nand U498 (N_498,In_1294,In_286);
nor U499 (N_499,In_28,In_1431);
nand U500 (N_500,In_293,In_1440);
and U501 (N_501,In_638,In_1127);
or U502 (N_502,In_243,In_871);
or U503 (N_503,In_1403,In_1113);
nor U504 (N_504,In_155,In_971);
nor U505 (N_505,In_126,In_1158);
nor U506 (N_506,In_1492,In_426);
and U507 (N_507,In_793,In_1327);
nor U508 (N_508,In_205,In_913);
and U509 (N_509,In_1165,In_718);
nand U510 (N_510,In_820,In_289);
and U511 (N_511,In_960,In_1317);
nor U512 (N_512,In_1241,In_824);
nor U513 (N_513,In_42,In_1172);
nand U514 (N_514,In_1066,In_919);
and U515 (N_515,In_502,In_1424);
nor U516 (N_516,In_361,In_38);
and U517 (N_517,In_808,In_511);
or U518 (N_518,In_1,In_1261);
nand U519 (N_519,In_933,In_373);
nand U520 (N_520,In_1304,In_313);
nand U521 (N_521,In_1063,In_187);
and U522 (N_522,In_664,In_1018);
and U523 (N_523,In_297,In_290);
nand U524 (N_524,In_427,In_665);
nand U525 (N_525,In_603,In_179);
nor U526 (N_526,In_762,In_932);
or U527 (N_527,In_1099,In_998);
or U528 (N_528,In_116,In_1070);
and U529 (N_529,In_1450,In_1296);
xnor U530 (N_530,In_1236,In_81);
xor U531 (N_531,In_573,In_687);
nor U532 (N_532,In_143,In_165);
or U533 (N_533,In_1348,In_570);
or U534 (N_534,In_779,In_43);
nand U535 (N_535,In_198,In_1497);
nand U536 (N_536,In_1343,In_351);
and U537 (N_537,In_210,In_546);
or U538 (N_538,In_1212,In_75);
nor U539 (N_539,In_1141,In_791);
or U540 (N_540,In_1435,In_1496);
nor U541 (N_541,In_925,In_761);
or U542 (N_542,In_722,In_940);
or U543 (N_543,In_288,In_1031);
nor U544 (N_544,In_477,In_1077);
nand U545 (N_545,In_1479,In_1464);
or U546 (N_546,In_705,In_1389);
and U547 (N_547,In_256,In_1368);
and U548 (N_548,In_82,In_1344);
nand U549 (N_549,In_1303,In_1349);
or U550 (N_550,In_785,In_247);
and U551 (N_551,In_195,In_597);
nand U552 (N_552,In_1408,In_1208);
nor U553 (N_553,In_697,In_654);
nand U554 (N_554,In_635,In_1140);
or U555 (N_555,In_646,In_966);
nor U556 (N_556,In_1056,In_917);
or U557 (N_557,In_898,In_1473);
or U558 (N_558,In_1144,In_340);
nand U559 (N_559,In_1363,In_1280);
or U560 (N_560,In_482,In_25);
and U561 (N_561,In_470,In_284);
nor U562 (N_562,In_905,In_628);
and U563 (N_563,In_1257,In_1019);
and U564 (N_564,In_1229,In_688);
and U565 (N_565,In_552,In_780);
nand U566 (N_566,In_579,In_1182);
or U567 (N_567,In_497,In_292);
and U568 (N_568,In_1106,In_1100);
nor U569 (N_569,In_389,In_886);
nor U570 (N_570,In_120,In_1116);
nand U571 (N_571,In_965,In_1330);
nand U572 (N_572,In_178,In_846);
nor U573 (N_573,In_33,In_1126);
nor U574 (N_574,In_157,In_1216);
or U575 (N_575,In_471,In_970);
nand U576 (N_576,In_601,In_1243);
and U577 (N_577,In_237,In_239);
and U578 (N_578,In_1495,In_1149);
nor U579 (N_579,In_630,In_1024);
nand U580 (N_580,In_807,In_324);
xor U581 (N_581,In_1290,In_641);
or U582 (N_582,In_627,In_1360);
xnor U583 (N_583,In_1249,In_1085);
nand U584 (N_584,In_448,In_1499);
or U585 (N_585,In_0,In_720);
xor U586 (N_586,In_510,In_1121);
nor U587 (N_587,In_508,In_804);
nand U588 (N_588,In_876,In_813);
or U589 (N_589,In_858,In_55);
nor U590 (N_590,In_1032,In_6);
or U591 (N_591,In_26,In_836);
and U592 (N_592,In_1189,In_647);
and U593 (N_593,In_91,In_1080);
or U594 (N_594,In_1357,In_390);
or U595 (N_595,In_241,In_1338);
nand U596 (N_596,In_1312,In_505);
and U597 (N_597,In_673,In_607);
and U598 (N_598,In_291,In_747);
nor U599 (N_599,In_652,In_859);
or U600 (N_600,In_1259,In_48);
nand U601 (N_601,In_235,In_1028);
or U602 (N_602,In_1191,In_1423);
nand U603 (N_603,In_786,In_7);
and U604 (N_604,In_963,In_283);
nor U605 (N_605,In_128,In_1395);
nor U606 (N_606,In_129,In_62);
nand U607 (N_607,In_1102,In_795);
nor U608 (N_608,In_405,In_152);
nand U609 (N_609,In_969,In_736);
and U610 (N_610,In_763,In_710);
nand U611 (N_611,In_594,In_650);
and U612 (N_612,In_49,In_637);
nor U613 (N_613,In_507,In_653);
nand U614 (N_614,In_1147,In_123);
nand U615 (N_615,In_1205,In_1459);
nand U616 (N_616,In_360,In_825);
or U617 (N_617,In_667,In_639);
nand U618 (N_618,In_122,In_1231);
or U619 (N_619,In_942,In_717);
or U620 (N_620,In_1002,In_577);
nand U621 (N_621,In_425,In_270);
nand U622 (N_622,In_1458,In_218);
nand U623 (N_623,In_977,In_992);
and U624 (N_624,In_1101,In_240);
and U625 (N_625,In_658,In_401);
nor U626 (N_626,In_707,In_996);
nor U627 (N_627,In_777,In_379);
and U628 (N_628,In_494,In_889);
nor U629 (N_629,In_73,In_236);
nor U630 (N_630,In_624,In_384);
and U631 (N_631,In_305,In_1210);
and U632 (N_632,In_1336,In_1481);
nand U633 (N_633,In_865,In_1151);
xnor U634 (N_634,In_104,In_212);
nor U635 (N_635,In_1498,In_1166);
nand U636 (N_636,In_1048,In_843);
and U637 (N_637,In_997,In_679);
and U638 (N_638,In_1157,In_926);
nand U639 (N_639,In_908,In_1442);
or U640 (N_640,In_588,In_216);
or U641 (N_641,In_1029,In_877);
and U642 (N_642,In_984,In_1393);
or U643 (N_643,In_1426,In_509);
and U644 (N_644,In_553,In_110);
nand U645 (N_645,In_790,In_645);
nand U646 (N_646,In_1104,In_462);
or U647 (N_647,In_300,In_85);
nor U648 (N_648,In_1045,In_1174);
nor U649 (N_649,In_875,In_781);
and U650 (N_650,In_370,In_124);
and U651 (N_651,In_109,In_1184);
nor U652 (N_652,In_910,In_677);
and U653 (N_653,In_1278,In_995);
and U654 (N_654,In_759,In_1493);
nor U655 (N_655,In_330,In_887);
nand U656 (N_656,In_938,In_1476);
nand U657 (N_657,In_1217,In_613);
nor U658 (N_658,In_1007,In_329);
nor U659 (N_659,In_65,In_649);
or U660 (N_660,In_1291,In_947);
nand U661 (N_661,In_1079,In_801);
nor U662 (N_662,In_1010,In_1494);
or U663 (N_663,In_1369,In_671);
or U664 (N_664,In_1035,In_936);
nand U665 (N_665,In_1224,In_1396);
and U666 (N_666,In_145,In_1117);
nor U667 (N_667,In_285,In_443);
nor U668 (N_668,In_466,In_45);
xor U669 (N_669,In_703,In_1475);
nor U670 (N_670,In_1388,In_622);
and U671 (N_671,In_1416,In_431);
or U672 (N_672,In_1111,In_935);
nand U673 (N_673,In_182,In_1260);
and U674 (N_674,In_393,In_1133);
nand U675 (N_675,In_228,In_381);
and U676 (N_676,In_512,In_34);
nand U677 (N_677,In_716,In_376);
xor U678 (N_678,In_383,In_480);
nor U679 (N_679,In_1443,In_387);
or U680 (N_680,In_1136,In_991);
or U681 (N_681,In_582,In_364);
nand U682 (N_682,In_133,In_173);
nand U683 (N_683,In_1196,In_1087);
or U684 (N_684,In_896,In_192);
nand U685 (N_685,In_172,In_231);
or U686 (N_686,In_18,In_312);
and U687 (N_687,In_772,In_1301);
nand U688 (N_688,In_968,In_1332);
nand U689 (N_689,In_743,In_994);
nor U690 (N_690,In_674,In_1230);
nand U691 (N_691,In_1046,In_180);
nand U692 (N_692,In_1405,In_1425);
nand U693 (N_693,In_1422,In_408);
xnor U694 (N_694,In_382,In_226);
nor U695 (N_695,In_1253,In_250);
or U696 (N_696,In_778,In_357);
and U697 (N_697,In_424,In_1122);
and U698 (N_698,In_1038,In_1214);
or U699 (N_699,In_83,In_1020);
nand U700 (N_700,In_948,In_857);
nand U701 (N_701,In_1039,In_914);
nand U702 (N_702,In_1447,In_539);
and U703 (N_703,In_32,In_287);
and U704 (N_704,In_386,In_894);
nand U705 (N_705,In_161,In_1486);
nand U706 (N_706,In_1355,In_260);
or U707 (N_707,In_199,In_818);
nor U708 (N_708,In_402,In_986);
nand U709 (N_709,In_847,In_125);
nand U710 (N_710,In_1474,In_1284);
nor U711 (N_711,In_756,In_276);
nand U712 (N_712,In_834,In_193);
nand U713 (N_713,In_119,In_1084);
or U714 (N_714,In_474,In_695);
nor U715 (N_715,In_1004,In_714);
or U716 (N_716,In_907,In_811);
or U717 (N_717,In_1258,In_275);
nand U718 (N_718,In_1023,In_1065);
nor U719 (N_719,In_1339,In_396);
and U720 (N_720,In_463,In_823);
and U721 (N_721,In_1397,In_1256);
nand U722 (N_722,In_1392,In_1276);
and U723 (N_723,In_1150,In_112);
nand U724 (N_724,In_738,In_39);
nand U725 (N_725,In_1434,In_89);
nor U726 (N_726,In_1091,In_1350);
and U727 (N_727,In_606,In_1469);
nand U728 (N_728,In_1188,In_523);
nor U729 (N_729,In_946,In_605);
and U730 (N_730,In_506,In_1381);
and U731 (N_731,In_394,In_483);
nor U732 (N_732,In_515,In_724);
or U733 (N_733,In_1152,In_232);
and U734 (N_734,In_5,In_841);
nor U735 (N_735,In_999,In_532);
and U736 (N_736,In_912,In_1321);
nand U737 (N_737,In_274,In_117);
nand U738 (N_738,In_96,In_1030);
and U739 (N_739,In_1176,In_71);
and U740 (N_740,In_937,In_1159);
and U741 (N_741,In_1255,In_74);
or U742 (N_742,In_315,In_1354);
nor U743 (N_743,In_856,In_1285);
nand U744 (N_744,In_1418,In_683);
nor U745 (N_745,In_623,In_768);
nor U746 (N_746,In_1173,In_69);
or U747 (N_747,In_1155,In_317);
nand U748 (N_748,In_400,In_648);
or U749 (N_749,In_833,In_16);
or U750 (N_750,In_1222,In_1303);
and U751 (N_751,In_1391,In_1478);
nand U752 (N_752,In_930,In_294);
nor U753 (N_753,In_1132,In_1044);
nand U754 (N_754,In_43,In_1194);
and U755 (N_755,In_811,In_1274);
or U756 (N_756,In_81,In_1090);
nand U757 (N_757,In_26,In_1047);
or U758 (N_758,In_931,In_260);
nand U759 (N_759,In_39,In_419);
and U760 (N_760,In_592,In_954);
or U761 (N_761,In_1033,In_1462);
nand U762 (N_762,In_23,In_40);
nor U763 (N_763,In_1200,In_1351);
and U764 (N_764,In_60,In_1192);
and U765 (N_765,In_432,In_421);
nand U766 (N_766,In_856,In_1043);
and U767 (N_767,In_986,In_1231);
or U768 (N_768,In_1114,In_215);
nand U769 (N_769,In_631,In_1248);
nand U770 (N_770,In_162,In_363);
nor U771 (N_771,In_1347,In_479);
xor U772 (N_772,In_558,In_1380);
and U773 (N_773,In_502,In_253);
and U774 (N_774,In_799,In_637);
nand U775 (N_775,In_1288,In_1331);
nor U776 (N_776,In_501,In_1397);
nand U777 (N_777,In_693,In_414);
nor U778 (N_778,In_1001,In_280);
and U779 (N_779,In_30,In_54);
and U780 (N_780,In_785,In_1326);
and U781 (N_781,In_1344,In_757);
nand U782 (N_782,In_4,In_904);
nand U783 (N_783,In_70,In_426);
and U784 (N_784,In_591,In_303);
or U785 (N_785,In_1015,In_1377);
nor U786 (N_786,In_1094,In_504);
or U787 (N_787,In_218,In_1000);
xnor U788 (N_788,In_758,In_1415);
nor U789 (N_789,In_65,In_853);
nor U790 (N_790,In_254,In_672);
and U791 (N_791,In_194,In_1056);
and U792 (N_792,In_306,In_1029);
nand U793 (N_793,In_174,In_649);
nor U794 (N_794,In_1274,In_1360);
nor U795 (N_795,In_78,In_990);
or U796 (N_796,In_1420,In_675);
xnor U797 (N_797,In_501,In_519);
or U798 (N_798,In_823,In_1364);
nand U799 (N_799,In_1197,In_506);
and U800 (N_800,In_254,In_947);
nand U801 (N_801,In_596,In_431);
and U802 (N_802,In_82,In_600);
nand U803 (N_803,In_1207,In_40);
nor U804 (N_804,In_1079,In_1489);
or U805 (N_805,In_1417,In_588);
nand U806 (N_806,In_45,In_741);
and U807 (N_807,In_1235,In_1073);
nor U808 (N_808,In_79,In_441);
nor U809 (N_809,In_579,In_1419);
nor U810 (N_810,In_109,In_982);
and U811 (N_811,In_1127,In_602);
or U812 (N_812,In_776,In_304);
nor U813 (N_813,In_1025,In_474);
nand U814 (N_814,In_893,In_1062);
nand U815 (N_815,In_1366,In_329);
or U816 (N_816,In_1209,In_315);
nand U817 (N_817,In_1318,In_624);
nor U818 (N_818,In_1214,In_1329);
xnor U819 (N_819,In_512,In_1484);
nor U820 (N_820,In_915,In_326);
nor U821 (N_821,In_286,In_789);
nand U822 (N_822,In_273,In_32);
xor U823 (N_823,In_942,In_741);
or U824 (N_824,In_1230,In_1207);
nand U825 (N_825,In_831,In_887);
and U826 (N_826,In_656,In_1397);
nand U827 (N_827,In_96,In_157);
nand U828 (N_828,In_1211,In_1259);
nand U829 (N_829,In_328,In_1324);
or U830 (N_830,In_364,In_1302);
nand U831 (N_831,In_1324,In_424);
or U832 (N_832,In_564,In_1072);
nor U833 (N_833,In_359,In_206);
or U834 (N_834,In_1211,In_605);
nor U835 (N_835,In_860,In_450);
nor U836 (N_836,In_156,In_746);
nand U837 (N_837,In_47,In_494);
or U838 (N_838,In_983,In_234);
nand U839 (N_839,In_109,In_1074);
nor U840 (N_840,In_1173,In_761);
or U841 (N_841,In_628,In_1276);
or U842 (N_842,In_101,In_528);
or U843 (N_843,In_508,In_678);
or U844 (N_844,In_976,In_165);
nor U845 (N_845,In_334,In_115);
nand U846 (N_846,In_895,In_945);
nor U847 (N_847,In_1349,In_8);
or U848 (N_848,In_298,In_1324);
or U849 (N_849,In_473,In_1248);
and U850 (N_850,In_712,In_79);
or U851 (N_851,In_108,In_757);
or U852 (N_852,In_633,In_1203);
and U853 (N_853,In_1435,In_670);
and U854 (N_854,In_196,In_712);
xnor U855 (N_855,In_1441,In_1190);
nand U856 (N_856,In_175,In_33);
nor U857 (N_857,In_1178,In_1194);
nand U858 (N_858,In_786,In_674);
nand U859 (N_859,In_1204,In_1135);
nor U860 (N_860,In_1255,In_36);
nand U861 (N_861,In_1154,In_600);
and U862 (N_862,In_503,In_237);
and U863 (N_863,In_144,In_72);
nand U864 (N_864,In_1241,In_783);
or U865 (N_865,In_1031,In_713);
and U866 (N_866,In_800,In_1272);
nand U867 (N_867,In_1337,In_710);
nor U868 (N_868,In_1419,In_1063);
nor U869 (N_869,In_688,In_730);
nand U870 (N_870,In_1343,In_1449);
or U871 (N_871,In_1223,In_640);
and U872 (N_872,In_608,In_1455);
and U873 (N_873,In_1492,In_1010);
nand U874 (N_874,In_787,In_504);
or U875 (N_875,In_709,In_1389);
nor U876 (N_876,In_1026,In_432);
or U877 (N_877,In_890,In_1449);
or U878 (N_878,In_1387,In_184);
nand U879 (N_879,In_1004,In_1050);
and U880 (N_880,In_106,In_846);
or U881 (N_881,In_915,In_1301);
nor U882 (N_882,In_812,In_1116);
nand U883 (N_883,In_81,In_71);
nor U884 (N_884,In_112,In_32);
nor U885 (N_885,In_243,In_767);
nand U886 (N_886,In_1475,In_718);
and U887 (N_887,In_209,In_1388);
or U888 (N_888,In_8,In_197);
nand U889 (N_889,In_164,In_1113);
nand U890 (N_890,In_1093,In_520);
nand U891 (N_891,In_82,In_276);
or U892 (N_892,In_317,In_1083);
nand U893 (N_893,In_699,In_21);
or U894 (N_894,In_239,In_33);
or U895 (N_895,In_942,In_836);
nand U896 (N_896,In_960,In_1327);
or U897 (N_897,In_491,In_1386);
xnor U898 (N_898,In_1023,In_270);
or U899 (N_899,In_738,In_43);
or U900 (N_900,In_917,In_1451);
nand U901 (N_901,In_699,In_1430);
nor U902 (N_902,In_396,In_131);
nand U903 (N_903,In_144,In_881);
nor U904 (N_904,In_175,In_1176);
xor U905 (N_905,In_647,In_1128);
or U906 (N_906,In_618,In_1061);
nor U907 (N_907,In_670,In_464);
nand U908 (N_908,In_417,In_1003);
nand U909 (N_909,In_699,In_554);
nor U910 (N_910,In_709,In_1082);
nor U911 (N_911,In_812,In_621);
nand U912 (N_912,In_118,In_1314);
or U913 (N_913,In_865,In_956);
or U914 (N_914,In_48,In_823);
nor U915 (N_915,In_124,In_1155);
or U916 (N_916,In_1069,In_415);
and U917 (N_917,In_102,In_1404);
or U918 (N_918,In_852,In_261);
nand U919 (N_919,In_277,In_160);
xor U920 (N_920,In_826,In_1442);
nand U921 (N_921,In_988,In_511);
nand U922 (N_922,In_428,In_889);
and U923 (N_923,In_333,In_632);
nor U924 (N_924,In_255,In_1079);
or U925 (N_925,In_627,In_810);
nand U926 (N_926,In_1239,In_28);
nor U927 (N_927,In_407,In_224);
or U928 (N_928,In_1045,In_1425);
and U929 (N_929,In_977,In_625);
or U930 (N_930,In_1193,In_606);
and U931 (N_931,In_1077,In_1417);
and U932 (N_932,In_1020,In_1255);
and U933 (N_933,In_1090,In_17);
nor U934 (N_934,In_274,In_1010);
nor U935 (N_935,In_530,In_1036);
or U936 (N_936,In_213,In_1136);
and U937 (N_937,In_274,In_338);
xor U938 (N_938,In_1321,In_1043);
and U939 (N_939,In_1019,In_164);
or U940 (N_940,In_248,In_681);
and U941 (N_941,In_627,In_915);
nor U942 (N_942,In_254,In_125);
or U943 (N_943,In_799,In_1287);
or U944 (N_944,In_591,In_1382);
nand U945 (N_945,In_199,In_839);
nand U946 (N_946,In_156,In_59);
or U947 (N_947,In_263,In_189);
nor U948 (N_948,In_546,In_1405);
or U949 (N_949,In_747,In_613);
nand U950 (N_950,In_313,In_13);
nand U951 (N_951,In_660,In_861);
and U952 (N_952,In_537,In_419);
and U953 (N_953,In_1286,In_719);
and U954 (N_954,In_373,In_1048);
nand U955 (N_955,In_1343,In_1363);
nor U956 (N_956,In_142,In_577);
nand U957 (N_957,In_647,In_855);
nor U958 (N_958,In_538,In_720);
and U959 (N_959,In_75,In_859);
xnor U960 (N_960,In_54,In_51);
nor U961 (N_961,In_159,In_1321);
nor U962 (N_962,In_1306,In_348);
nand U963 (N_963,In_1135,In_1364);
nand U964 (N_964,In_151,In_1258);
or U965 (N_965,In_1259,In_1404);
nor U966 (N_966,In_652,In_705);
nor U967 (N_967,In_680,In_292);
or U968 (N_968,In_541,In_1024);
or U969 (N_969,In_426,In_1064);
and U970 (N_970,In_630,In_1145);
xor U971 (N_971,In_345,In_14);
xnor U972 (N_972,In_811,In_399);
nor U973 (N_973,In_1376,In_793);
nor U974 (N_974,In_244,In_300);
nand U975 (N_975,In_763,In_887);
or U976 (N_976,In_877,In_109);
or U977 (N_977,In_999,In_1043);
nand U978 (N_978,In_7,In_830);
and U979 (N_979,In_84,In_545);
or U980 (N_980,In_557,In_1055);
nor U981 (N_981,In_710,In_1214);
and U982 (N_982,In_1472,In_675);
nand U983 (N_983,In_991,In_579);
nor U984 (N_984,In_363,In_268);
nand U985 (N_985,In_935,In_393);
xnor U986 (N_986,In_375,In_1133);
or U987 (N_987,In_1052,In_1275);
and U988 (N_988,In_1358,In_231);
or U989 (N_989,In_1010,In_50);
nand U990 (N_990,In_1435,In_281);
nand U991 (N_991,In_941,In_701);
or U992 (N_992,In_715,In_1271);
nor U993 (N_993,In_250,In_1401);
nor U994 (N_994,In_850,In_1412);
nand U995 (N_995,In_792,In_712);
nor U996 (N_996,In_1063,In_676);
nor U997 (N_997,In_447,In_888);
nand U998 (N_998,In_419,In_525);
nor U999 (N_999,In_609,In_734);
xor U1000 (N_1000,In_496,In_1063);
or U1001 (N_1001,In_487,In_854);
nand U1002 (N_1002,In_364,In_1365);
nor U1003 (N_1003,In_650,In_1437);
or U1004 (N_1004,In_446,In_60);
and U1005 (N_1005,In_744,In_48);
nor U1006 (N_1006,In_688,In_501);
nor U1007 (N_1007,In_1351,In_664);
nand U1008 (N_1008,In_1280,In_333);
and U1009 (N_1009,In_113,In_684);
nand U1010 (N_1010,In_1003,In_480);
or U1011 (N_1011,In_1200,In_247);
or U1012 (N_1012,In_1114,In_600);
or U1013 (N_1013,In_1285,In_1320);
nand U1014 (N_1014,In_1491,In_158);
or U1015 (N_1015,In_756,In_1218);
and U1016 (N_1016,In_22,In_554);
and U1017 (N_1017,In_980,In_490);
and U1018 (N_1018,In_268,In_1247);
nand U1019 (N_1019,In_857,In_547);
and U1020 (N_1020,In_362,In_207);
nand U1021 (N_1021,In_127,In_855);
nand U1022 (N_1022,In_956,In_1021);
nor U1023 (N_1023,In_876,In_1215);
or U1024 (N_1024,In_591,In_9);
nand U1025 (N_1025,In_919,In_1255);
nor U1026 (N_1026,In_1384,In_539);
or U1027 (N_1027,In_823,In_142);
nor U1028 (N_1028,In_533,In_874);
or U1029 (N_1029,In_1104,In_1032);
nor U1030 (N_1030,In_284,In_882);
nor U1031 (N_1031,In_1087,In_582);
or U1032 (N_1032,In_725,In_761);
nand U1033 (N_1033,In_846,In_1076);
and U1034 (N_1034,In_1351,In_575);
nor U1035 (N_1035,In_259,In_1466);
nand U1036 (N_1036,In_583,In_286);
or U1037 (N_1037,In_1008,In_582);
nand U1038 (N_1038,In_403,In_46);
nor U1039 (N_1039,In_1206,In_1341);
nand U1040 (N_1040,In_1291,In_973);
nor U1041 (N_1041,In_405,In_650);
nand U1042 (N_1042,In_1412,In_306);
or U1043 (N_1043,In_1266,In_63);
nor U1044 (N_1044,In_882,In_1209);
nand U1045 (N_1045,In_1019,In_1303);
or U1046 (N_1046,In_392,In_1432);
nand U1047 (N_1047,In_236,In_888);
nor U1048 (N_1048,In_944,In_780);
nand U1049 (N_1049,In_906,In_1420);
nor U1050 (N_1050,In_430,In_371);
and U1051 (N_1051,In_1248,In_1211);
and U1052 (N_1052,In_698,In_950);
nor U1053 (N_1053,In_214,In_330);
or U1054 (N_1054,In_836,In_49);
nor U1055 (N_1055,In_287,In_935);
nand U1056 (N_1056,In_19,In_1364);
or U1057 (N_1057,In_1110,In_847);
or U1058 (N_1058,In_139,In_25);
nor U1059 (N_1059,In_1188,In_1373);
nand U1060 (N_1060,In_931,In_118);
or U1061 (N_1061,In_470,In_101);
and U1062 (N_1062,In_1380,In_966);
nand U1063 (N_1063,In_1450,In_428);
and U1064 (N_1064,In_651,In_153);
nand U1065 (N_1065,In_456,In_807);
or U1066 (N_1066,In_1266,In_345);
nand U1067 (N_1067,In_752,In_626);
nor U1068 (N_1068,In_1126,In_672);
or U1069 (N_1069,In_392,In_444);
nor U1070 (N_1070,In_1081,In_295);
or U1071 (N_1071,In_61,In_759);
nor U1072 (N_1072,In_266,In_273);
or U1073 (N_1073,In_1334,In_1118);
and U1074 (N_1074,In_1058,In_766);
and U1075 (N_1075,In_213,In_259);
nor U1076 (N_1076,In_210,In_442);
nand U1077 (N_1077,In_140,In_1459);
or U1078 (N_1078,In_881,In_431);
or U1079 (N_1079,In_377,In_287);
and U1080 (N_1080,In_117,In_249);
nor U1081 (N_1081,In_390,In_1085);
nand U1082 (N_1082,In_223,In_523);
nor U1083 (N_1083,In_980,In_1324);
nor U1084 (N_1084,In_606,In_251);
or U1085 (N_1085,In_66,In_222);
nand U1086 (N_1086,In_676,In_989);
or U1087 (N_1087,In_683,In_1132);
nor U1088 (N_1088,In_1123,In_966);
and U1089 (N_1089,In_243,In_751);
or U1090 (N_1090,In_737,In_491);
nand U1091 (N_1091,In_82,In_941);
or U1092 (N_1092,In_979,In_566);
nand U1093 (N_1093,In_87,In_4);
nor U1094 (N_1094,In_1295,In_259);
and U1095 (N_1095,In_950,In_613);
nand U1096 (N_1096,In_91,In_1302);
and U1097 (N_1097,In_1089,In_705);
nand U1098 (N_1098,In_892,In_274);
nand U1099 (N_1099,In_541,In_962);
nor U1100 (N_1100,In_653,In_681);
or U1101 (N_1101,In_739,In_1322);
nor U1102 (N_1102,In_936,In_41);
and U1103 (N_1103,In_948,In_412);
and U1104 (N_1104,In_458,In_337);
or U1105 (N_1105,In_1449,In_1469);
nand U1106 (N_1106,In_184,In_691);
xnor U1107 (N_1107,In_1092,In_1347);
and U1108 (N_1108,In_729,In_437);
or U1109 (N_1109,In_275,In_410);
nand U1110 (N_1110,In_1230,In_614);
nor U1111 (N_1111,In_635,In_743);
nand U1112 (N_1112,In_1064,In_1225);
nor U1113 (N_1113,In_1474,In_58);
or U1114 (N_1114,In_957,In_123);
or U1115 (N_1115,In_529,In_1424);
nor U1116 (N_1116,In_675,In_1004);
and U1117 (N_1117,In_441,In_1373);
xor U1118 (N_1118,In_232,In_128);
nor U1119 (N_1119,In_523,In_326);
or U1120 (N_1120,In_962,In_219);
nor U1121 (N_1121,In_1173,In_626);
nand U1122 (N_1122,In_977,In_877);
and U1123 (N_1123,In_5,In_282);
and U1124 (N_1124,In_28,In_463);
xor U1125 (N_1125,In_541,In_201);
and U1126 (N_1126,In_1099,In_283);
or U1127 (N_1127,In_685,In_1012);
nor U1128 (N_1128,In_330,In_1225);
and U1129 (N_1129,In_1364,In_1004);
or U1130 (N_1130,In_572,In_550);
nand U1131 (N_1131,In_601,In_1015);
and U1132 (N_1132,In_1037,In_270);
and U1133 (N_1133,In_296,In_1313);
and U1134 (N_1134,In_418,In_990);
and U1135 (N_1135,In_1219,In_816);
nor U1136 (N_1136,In_231,In_1339);
or U1137 (N_1137,In_383,In_178);
nor U1138 (N_1138,In_560,In_1304);
and U1139 (N_1139,In_518,In_1194);
and U1140 (N_1140,In_960,In_878);
nor U1141 (N_1141,In_1030,In_287);
nor U1142 (N_1142,In_551,In_318);
nor U1143 (N_1143,In_1283,In_1127);
and U1144 (N_1144,In_176,In_512);
nand U1145 (N_1145,In_611,In_688);
or U1146 (N_1146,In_12,In_646);
nor U1147 (N_1147,In_189,In_168);
nand U1148 (N_1148,In_294,In_94);
or U1149 (N_1149,In_586,In_921);
or U1150 (N_1150,In_1412,In_1391);
or U1151 (N_1151,In_450,In_228);
nand U1152 (N_1152,In_1188,In_902);
nand U1153 (N_1153,In_768,In_1162);
nand U1154 (N_1154,In_407,In_1090);
nor U1155 (N_1155,In_1495,In_1463);
and U1156 (N_1156,In_869,In_347);
and U1157 (N_1157,In_445,In_98);
and U1158 (N_1158,In_1410,In_887);
nand U1159 (N_1159,In_1066,In_251);
nand U1160 (N_1160,In_590,In_757);
and U1161 (N_1161,In_1376,In_399);
nor U1162 (N_1162,In_1152,In_1162);
and U1163 (N_1163,In_819,In_166);
and U1164 (N_1164,In_1000,In_1268);
or U1165 (N_1165,In_537,In_1356);
nand U1166 (N_1166,In_930,In_777);
or U1167 (N_1167,In_1382,In_1213);
nor U1168 (N_1168,In_917,In_1036);
or U1169 (N_1169,In_235,In_585);
nor U1170 (N_1170,In_44,In_857);
nor U1171 (N_1171,In_310,In_894);
or U1172 (N_1172,In_388,In_513);
and U1173 (N_1173,In_1394,In_168);
or U1174 (N_1174,In_421,In_1493);
nand U1175 (N_1175,In_1209,In_65);
nand U1176 (N_1176,In_742,In_696);
and U1177 (N_1177,In_901,In_704);
nor U1178 (N_1178,In_652,In_515);
and U1179 (N_1179,In_51,In_754);
and U1180 (N_1180,In_765,In_853);
or U1181 (N_1181,In_342,In_639);
and U1182 (N_1182,In_744,In_1406);
xor U1183 (N_1183,In_597,In_638);
or U1184 (N_1184,In_1084,In_1253);
and U1185 (N_1185,In_435,In_1145);
nand U1186 (N_1186,In_476,In_123);
or U1187 (N_1187,In_681,In_1106);
nand U1188 (N_1188,In_984,In_31);
or U1189 (N_1189,In_1473,In_520);
or U1190 (N_1190,In_850,In_1080);
or U1191 (N_1191,In_776,In_1405);
nand U1192 (N_1192,In_109,In_487);
nor U1193 (N_1193,In_41,In_308);
xnor U1194 (N_1194,In_121,In_590);
nor U1195 (N_1195,In_1017,In_329);
or U1196 (N_1196,In_1151,In_964);
or U1197 (N_1197,In_1044,In_164);
or U1198 (N_1198,In_1086,In_853);
nor U1199 (N_1199,In_1379,In_519);
nor U1200 (N_1200,In_24,In_753);
and U1201 (N_1201,In_922,In_394);
nor U1202 (N_1202,In_915,In_1429);
nor U1203 (N_1203,In_851,In_889);
nand U1204 (N_1204,In_471,In_23);
nand U1205 (N_1205,In_1392,In_963);
nand U1206 (N_1206,In_1112,In_989);
nand U1207 (N_1207,In_411,In_109);
nand U1208 (N_1208,In_561,In_581);
and U1209 (N_1209,In_16,In_515);
or U1210 (N_1210,In_367,In_1026);
nor U1211 (N_1211,In_306,In_1334);
nand U1212 (N_1212,In_83,In_385);
or U1213 (N_1213,In_327,In_1054);
or U1214 (N_1214,In_986,In_1281);
and U1215 (N_1215,In_463,In_357);
and U1216 (N_1216,In_1242,In_711);
nand U1217 (N_1217,In_484,In_928);
nand U1218 (N_1218,In_621,In_212);
nand U1219 (N_1219,In_1338,In_831);
or U1220 (N_1220,In_1451,In_570);
nor U1221 (N_1221,In_1033,In_249);
or U1222 (N_1222,In_400,In_602);
or U1223 (N_1223,In_497,In_1032);
nor U1224 (N_1224,In_264,In_733);
nor U1225 (N_1225,In_915,In_1199);
and U1226 (N_1226,In_493,In_1206);
and U1227 (N_1227,In_1355,In_957);
or U1228 (N_1228,In_383,In_481);
nand U1229 (N_1229,In_1462,In_1088);
or U1230 (N_1230,In_16,In_26);
or U1231 (N_1231,In_1442,In_939);
nand U1232 (N_1232,In_591,In_668);
nand U1233 (N_1233,In_110,In_803);
nor U1234 (N_1234,In_1311,In_1419);
or U1235 (N_1235,In_695,In_855);
nand U1236 (N_1236,In_1397,In_264);
and U1237 (N_1237,In_526,In_577);
nand U1238 (N_1238,In_467,In_463);
nand U1239 (N_1239,In_1171,In_157);
nor U1240 (N_1240,In_1362,In_31);
and U1241 (N_1241,In_82,In_333);
and U1242 (N_1242,In_945,In_920);
nand U1243 (N_1243,In_1364,In_631);
nand U1244 (N_1244,In_346,In_1080);
xnor U1245 (N_1245,In_1074,In_507);
nand U1246 (N_1246,In_167,In_1030);
or U1247 (N_1247,In_1400,In_96);
or U1248 (N_1248,In_104,In_1455);
nand U1249 (N_1249,In_110,In_183);
and U1250 (N_1250,In_954,In_991);
nand U1251 (N_1251,In_1008,In_879);
nor U1252 (N_1252,In_339,In_1018);
nand U1253 (N_1253,In_241,In_1347);
nand U1254 (N_1254,In_619,In_637);
or U1255 (N_1255,In_493,In_982);
nand U1256 (N_1256,In_421,In_738);
xnor U1257 (N_1257,In_1104,In_440);
or U1258 (N_1258,In_1186,In_1007);
nor U1259 (N_1259,In_1352,In_594);
nor U1260 (N_1260,In_477,In_116);
and U1261 (N_1261,In_977,In_1445);
or U1262 (N_1262,In_410,In_813);
nand U1263 (N_1263,In_374,In_25);
nor U1264 (N_1264,In_890,In_770);
nand U1265 (N_1265,In_131,In_55);
and U1266 (N_1266,In_1182,In_1150);
or U1267 (N_1267,In_1171,In_364);
nand U1268 (N_1268,In_1410,In_97);
or U1269 (N_1269,In_809,In_972);
nor U1270 (N_1270,In_369,In_241);
xnor U1271 (N_1271,In_316,In_84);
and U1272 (N_1272,In_988,In_186);
nand U1273 (N_1273,In_241,In_1116);
nor U1274 (N_1274,In_899,In_662);
nor U1275 (N_1275,In_950,In_1065);
nor U1276 (N_1276,In_63,In_534);
or U1277 (N_1277,In_1186,In_1046);
and U1278 (N_1278,In_1251,In_1390);
or U1279 (N_1279,In_609,In_39);
and U1280 (N_1280,In_1470,In_442);
nand U1281 (N_1281,In_1402,In_740);
and U1282 (N_1282,In_7,In_550);
or U1283 (N_1283,In_849,In_191);
nand U1284 (N_1284,In_112,In_1194);
nand U1285 (N_1285,In_313,In_1007);
and U1286 (N_1286,In_1232,In_1047);
nand U1287 (N_1287,In_121,In_519);
nor U1288 (N_1288,In_141,In_799);
nand U1289 (N_1289,In_607,In_467);
or U1290 (N_1290,In_735,In_1290);
nor U1291 (N_1291,In_508,In_1303);
and U1292 (N_1292,In_970,In_442);
or U1293 (N_1293,In_75,In_351);
and U1294 (N_1294,In_241,In_126);
nor U1295 (N_1295,In_1184,In_1001);
nor U1296 (N_1296,In_178,In_1093);
and U1297 (N_1297,In_99,In_757);
nand U1298 (N_1298,In_271,In_118);
nand U1299 (N_1299,In_1460,In_1394);
nand U1300 (N_1300,In_723,In_611);
nand U1301 (N_1301,In_326,In_1327);
and U1302 (N_1302,In_1461,In_727);
nor U1303 (N_1303,In_703,In_285);
nor U1304 (N_1304,In_1079,In_369);
or U1305 (N_1305,In_199,In_311);
and U1306 (N_1306,In_114,In_176);
nand U1307 (N_1307,In_1464,In_1416);
nor U1308 (N_1308,In_19,In_11);
nor U1309 (N_1309,In_936,In_850);
and U1310 (N_1310,In_271,In_813);
nor U1311 (N_1311,In_399,In_227);
and U1312 (N_1312,In_479,In_463);
and U1313 (N_1313,In_1469,In_551);
nand U1314 (N_1314,In_1426,In_870);
or U1315 (N_1315,In_448,In_962);
or U1316 (N_1316,In_832,In_1119);
and U1317 (N_1317,In_282,In_1032);
nand U1318 (N_1318,In_606,In_780);
and U1319 (N_1319,In_1273,In_1228);
nor U1320 (N_1320,In_246,In_203);
nand U1321 (N_1321,In_1207,In_528);
nor U1322 (N_1322,In_76,In_1198);
and U1323 (N_1323,In_733,In_471);
nand U1324 (N_1324,In_35,In_794);
nand U1325 (N_1325,In_100,In_1032);
nand U1326 (N_1326,In_577,In_386);
nand U1327 (N_1327,In_1038,In_728);
nand U1328 (N_1328,In_288,In_278);
nand U1329 (N_1329,In_739,In_1272);
and U1330 (N_1330,In_84,In_752);
and U1331 (N_1331,In_127,In_809);
and U1332 (N_1332,In_417,In_690);
nor U1333 (N_1333,In_383,In_693);
nor U1334 (N_1334,In_596,In_320);
and U1335 (N_1335,In_957,In_800);
xor U1336 (N_1336,In_369,In_408);
and U1337 (N_1337,In_345,In_1344);
xor U1338 (N_1338,In_1147,In_971);
xnor U1339 (N_1339,In_1191,In_977);
and U1340 (N_1340,In_611,In_624);
and U1341 (N_1341,In_736,In_1167);
nand U1342 (N_1342,In_872,In_25);
and U1343 (N_1343,In_1025,In_143);
or U1344 (N_1344,In_325,In_114);
nand U1345 (N_1345,In_1349,In_1174);
and U1346 (N_1346,In_669,In_931);
nand U1347 (N_1347,In_1323,In_627);
nand U1348 (N_1348,In_375,In_1275);
nor U1349 (N_1349,In_1245,In_724);
nor U1350 (N_1350,In_247,In_1343);
nand U1351 (N_1351,In_603,In_36);
nor U1352 (N_1352,In_354,In_1457);
nand U1353 (N_1353,In_1083,In_1165);
and U1354 (N_1354,In_1460,In_509);
xnor U1355 (N_1355,In_1402,In_931);
nand U1356 (N_1356,In_419,In_646);
xor U1357 (N_1357,In_390,In_893);
nand U1358 (N_1358,In_608,In_628);
nor U1359 (N_1359,In_792,In_1447);
or U1360 (N_1360,In_1260,In_653);
and U1361 (N_1361,In_69,In_522);
or U1362 (N_1362,In_684,In_1445);
nand U1363 (N_1363,In_1230,In_1373);
nand U1364 (N_1364,In_1164,In_709);
nand U1365 (N_1365,In_1481,In_768);
nor U1366 (N_1366,In_293,In_1397);
nand U1367 (N_1367,In_1133,In_1482);
and U1368 (N_1368,In_809,In_283);
nor U1369 (N_1369,In_453,In_23);
or U1370 (N_1370,In_941,In_994);
nand U1371 (N_1371,In_641,In_706);
nand U1372 (N_1372,In_646,In_380);
and U1373 (N_1373,In_96,In_283);
nand U1374 (N_1374,In_300,In_168);
and U1375 (N_1375,In_12,In_834);
and U1376 (N_1376,In_855,In_339);
or U1377 (N_1377,In_649,In_1222);
nand U1378 (N_1378,In_500,In_93);
or U1379 (N_1379,In_108,In_561);
or U1380 (N_1380,In_50,In_333);
nor U1381 (N_1381,In_1026,In_1380);
or U1382 (N_1382,In_459,In_1317);
or U1383 (N_1383,In_38,In_396);
nor U1384 (N_1384,In_1275,In_529);
nor U1385 (N_1385,In_740,In_1327);
nor U1386 (N_1386,In_52,In_821);
or U1387 (N_1387,In_22,In_369);
and U1388 (N_1388,In_288,In_974);
or U1389 (N_1389,In_376,In_429);
and U1390 (N_1390,In_1144,In_415);
nor U1391 (N_1391,In_55,In_80);
or U1392 (N_1392,In_921,In_1434);
or U1393 (N_1393,In_1480,In_1380);
nand U1394 (N_1394,In_380,In_503);
and U1395 (N_1395,In_1254,In_747);
nand U1396 (N_1396,In_1480,In_685);
and U1397 (N_1397,In_1314,In_1064);
nand U1398 (N_1398,In_1386,In_314);
nand U1399 (N_1399,In_822,In_366);
nor U1400 (N_1400,In_594,In_1292);
nor U1401 (N_1401,In_104,In_718);
nor U1402 (N_1402,In_123,In_211);
or U1403 (N_1403,In_1386,In_848);
nand U1404 (N_1404,In_419,In_721);
nand U1405 (N_1405,In_416,In_1333);
or U1406 (N_1406,In_188,In_10);
nor U1407 (N_1407,In_1016,In_1088);
or U1408 (N_1408,In_1219,In_1098);
and U1409 (N_1409,In_1036,In_509);
xor U1410 (N_1410,In_398,In_854);
nor U1411 (N_1411,In_1246,In_444);
nand U1412 (N_1412,In_1441,In_67);
nand U1413 (N_1413,In_1435,In_1369);
and U1414 (N_1414,In_720,In_417);
nor U1415 (N_1415,In_249,In_94);
and U1416 (N_1416,In_18,In_807);
nand U1417 (N_1417,In_368,In_197);
or U1418 (N_1418,In_305,In_176);
or U1419 (N_1419,In_1025,In_684);
nor U1420 (N_1420,In_580,In_613);
or U1421 (N_1421,In_1067,In_962);
nor U1422 (N_1422,In_322,In_232);
or U1423 (N_1423,In_755,In_416);
nand U1424 (N_1424,In_970,In_1121);
or U1425 (N_1425,In_655,In_871);
nand U1426 (N_1426,In_1499,In_1287);
or U1427 (N_1427,In_565,In_411);
nand U1428 (N_1428,In_1344,In_1278);
or U1429 (N_1429,In_1192,In_197);
and U1430 (N_1430,In_1284,In_608);
nor U1431 (N_1431,In_64,In_1075);
nand U1432 (N_1432,In_676,In_1391);
and U1433 (N_1433,In_215,In_1411);
nor U1434 (N_1434,In_3,In_24);
nand U1435 (N_1435,In_800,In_784);
nand U1436 (N_1436,In_757,In_1456);
nand U1437 (N_1437,In_1023,In_334);
nor U1438 (N_1438,In_1154,In_1014);
nor U1439 (N_1439,In_703,In_462);
and U1440 (N_1440,In_929,In_619);
and U1441 (N_1441,In_373,In_353);
nor U1442 (N_1442,In_206,In_360);
or U1443 (N_1443,In_84,In_1038);
or U1444 (N_1444,In_79,In_1011);
nand U1445 (N_1445,In_471,In_794);
nand U1446 (N_1446,In_1476,In_1359);
nand U1447 (N_1447,In_916,In_1490);
and U1448 (N_1448,In_1175,In_1101);
and U1449 (N_1449,In_1402,In_412);
and U1450 (N_1450,In_880,In_1430);
and U1451 (N_1451,In_1243,In_471);
or U1452 (N_1452,In_549,In_825);
or U1453 (N_1453,In_527,In_834);
nor U1454 (N_1454,In_1198,In_686);
nor U1455 (N_1455,In_164,In_1040);
and U1456 (N_1456,In_1342,In_663);
nand U1457 (N_1457,In_692,In_1010);
nand U1458 (N_1458,In_1239,In_656);
or U1459 (N_1459,In_1261,In_587);
nor U1460 (N_1460,In_127,In_1327);
and U1461 (N_1461,In_993,In_1329);
nor U1462 (N_1462,In_1321,In_624);
nor U1463 (N_1463,In_1246,In_439);
or U1464 (N_1464,In_843,In_788);
nand U1465 (N_1465,In_752,In_1173);
nand U1466 (N_1466,In_1360,In_853);
nor U1467 (N_1467,In_1372,In_1217);
or U1468 (N_1468,In_1033,In_818);
nand U1469 (N_1469,In_1195,In_387);
and U1470 (N_1470,In_899,In_938);
and U1471 (N_1471,In_541,In_1298);
nor U1472 (N_1472,In_1094,In_774);
or U1473 (N_1473,In_93,In_481);
nand U1474 (N_1474,In_560,In_997);
or U1475 (N_1475,In_259,In_708);
nor U1476 (N_1476,In_635,In_828);
nand U1477 (N_1477,In_1409,In_51);
and U1478 (N_1478,In_295,In_1391);
or U1479 (N_1479,In_227,In_649);
or U1480 (N_1480,In_504,In_207);
or U1481 (N_1481,In_773,In_1354);
and U1482 (N_1482,In_81,In_412);
nor U1483 (N_1483,In_1173,In_131);
or U1484 (N_1484,In_701,In_1317);
or U1485 (N_1485,In_1208,In_1377);
or U1486 (N_1486,In_677,In_10);
or U1487 (N_1487,In_1281,In_770);
or U1488 (N_1488,In_979,In_131);
nand U1489 (N_1489,In_694,In_1423);
or U1490 (N_1490,In_1196,In_208);
nand U1491 (N_1491,In_98,In_795);
nor U1492 (N_1492,In_994,In_1123);
and U1493 (N_1493,In_264,In_240);
and U1494 (N_1494,In_105,In_603);
and U1495 (N_1495,In_1178,In_241);
and U1496 (N_1496,In_1222,In_863);
or U1497 (N_1497,In_169,In_401);
or U1498 (N_1498,In_741,In_1309);
or U1499 (N_1499,In_1205,In_1019);
and U1500 (N_1500,In_167,In_887);
and U1501 (N_1501,In_769,In_1238);
and U1502 (N_1502,In_1028,In_241);
or U1503 (N_1503,In_1103,In_1200);
and U1504 (N_1504,In_1071,In_1400);
nor U1505 (N_1505,In_636,In_565);
nand U1506 (N_1506,In_1377,In_1407);
and U1507 (N_1507,In_1376,In_105);
nand U1508 (N_1508,In_101,In_987);
or U1509 (N_1509,In_1381,In_821);
and U1510 (N_1510,In_914,In_1480);
or U1511 (N_1511,In_1202,In_506);
nand U1512 (N_1512,In_971,In_1201);
and U1513 (N_1513,In_244,In_94);
xnor U1514 (N_1514,In_461,In_198);
nand U1515 (N_1515,In_623,In_941);
nor U1516 (N_1516,In_50,In_1230);
nand U1517 (N_1517,In_825,In_622);
nor U1518 (N_1518,In_427,In_199);
nor U1519 (N_1519,In_864,In_116);
nor U1520 (N_1520,In_439,In_413);
and U1521 (N_1521,In_122,In_195);
and U1522 (N_1522,In_340,In_678);
nor U1523 (N_1523,In_786,In_235);
nor U1524 (N_1524,In_754,In_848);
nand U1525 (N_1525,In_123,In_1437);
or U1526 (N_1526,In_475,In_202);
nand U1527 (N_1527,In_372,In_1260);
nor U1528 (N_1528,In_264,In_1325);
nor U1529 (N_1529,In_1336,In_978);
and U1530 (N_1530,In_201,In_1331);
and U1531 (N_1531,In_1158,In_176);
nand U1532 (N_1532,In_1450,In_524);
nand U1533 (N_1533,In_1016,In_1292);
nor U1534 (N_1534,In_106,In_39);
nand U1535 (N_1535,In_421,In_202);
nor U1536 (N_1536,In_722,In_943);
and U1537 (N_1537,In_1255,In_260);
or U1538 (N_1538,In_1051,In_592);
or U1539 (N_1539,In_617,In_385);
or U1540 (N_1540,In_1124,In_888);
nor U1541 (N_1541,In_910,In_485);
nor U1542 (N_1542,In_270,In_1222);
xnor U1543 (N_1543,In_1098,In_954);
and U1544 (N_1544,In_1362,In_1169);
nor U1545 (N_1545,In_1292,In_1132);
and U1546 (N_1546,In_1393,In_1435);
and U1547 (N_1547,In_283,In_1088);
and U1548 (N_1548,In_690,In_266);
nand U1549 (N_1549,In_821,In_487);
nor U1550 (N_1550,In_1327,In_768);
and U1551 (N_1551,In_251,In_1192);
nor U1552 (N_1552,In_754,In_1073);
and U1553 (N_1553,In_444,In_614);
nand U1554 (N_1554,In_796,In_224);
nand U1555 (N_1555,In_941,In_847);
or U1556 (N_1556,In_818,In_710);
nand U1557 (N_1557,In_888,In_1277);
and U1558 (N_1558,In_366,In_20);
nand U1559 (N_1559,In_1490,In_1027);
or U1560 (N_1560,In_840,In_716);
nor U1561 (N_1561,In_155,In_1119);
nand U1562 (N_1562,In_602,In_1477);
nand U1563 (N_1563,In_95,In_1010);
nand U1564 (N_1564,In_75,In_206);
nand U1565 (N_1565,In_260,In_559);
nor U1566 (N_1566,In_710,In_1254);
and U1567 (N_1567,In_1345,In_416);
and U1568 (N_1568,In_1033,In_588);
and U1569 (N_1569,In_1133,In_623);
and U1570 (N_1570,In_301,In_565);
and U1571 (N_1571,In_244,In_1300);
nand U1572 (N_1572,In_537,In_673);
or U1573 (N_1573,In_810,In_351);
nor U1574 (N_1574,In_807,In_288);
or U1575 (N_1575,In_1445,In_902);
nand U1576 (N_1576,In_847,In_593);
nand U1577 (N_1577,In_818,In_1440);
or U1578 (N_1578,In_252,In_385);
nand U1579 (N_1579,In_818,In_1094);
nand U1580 (N_1580,In_1042,In_286);
nor U1581 (N_1581,In_36,In_138);
nand U1582 (N_1582,In_494,In_1448);
nor U1583 (N_1583,In_1188,In_807);
or U1584 (N_1584,In_1123,In_1459);
nor U1585 (N_1585,In_407,In_804);
and U1586 (N_1586,In_1256,In_1277);
nand U1587 (N_1587,In_731,In_102);
nor U1588 (N_1588,In_891,In_18);
nor U1589 (N_1589,In_1299,In_1480);
nand U1590 (N_1590,In_582,In_993);
nand U1591 (N_1591,In_1414,In_1187);
nand U1592 (N_1592,In_317,In_879);
nor U1593 (N_1593,In_1182,In_571);
and U1594 (N_1594,In_695,In_104);
nor U1595 (N_1595,In_70,In_1328);
nor U1596 (N_1596,In_601,In_702);
or U1597 (N_1597,In_1468,In_833);
or U1598 (N_1598,In_837,In_275);
nand U1599 (N_1599,In_1115,In_1162);
nand U1600 (N_1600,In_86,In_410);
nand U1601 (N_1601,In_264,In_29);
nor U1602 (N_1602,In_834,In_318);
and U1603 (N_1603,In_329,In_1355);
and U1604 (N_1604,In_176,In_1399);
nand U1605 (N_1605,In_981,In_226);
or U1606 (N_1606,In_1472,In_1166);
or U1607 (N_1607,In_313,In_505);
nand U1608 (N_1608,In_484,In_1196);
or U1609 (N_1609,In_540,In_1369);
nand U1610 (N_1610,In_398,In_1048);
nor U1611 (N_1611,In_1107,In_47);
or U1612 (N_1612,In_927,In_1101);
and U1613 (N_1613,In_833,In_406);
xor U1614 (N_1614,In_129,In_208);
nand U1615 (N_1615,In_218,In_138);
or U1616 (N_1616,In_1079,In_804);
nand U1617 (N_1617,In_82,In_417);
nand U1618 (N_1618,In_557,In_957);
or U1619 (N_1619,In_543,In_1317);
nand U1620 (N_1620,In_591,In_1109);
nor U1621 (N_1621,In_1110,In_522);
nand U1622 (N_1622,In_366,In_75);
xor U1623 (N_1623,In_424,In_1428);
nor U1624 (N_1624,In_1007,In_305);
and U1625 (N_1625,In_1338,In_30);
or U1626 (N_1626,In_1014,In_591);
nor U1627 (N_1627,In_1470,In_43);
and U1628 (N_1628,In_234,In_459);
and U1629 (N_1629,In_1448,In_553);
and U1630 (N_1630,In_83,In_520);
or U1631 (N_1631,In_1276,In_1480);
and U1632 (N_1632,In_432,In_1038);
or U1633 (N_1633,In_395,In_105);
and U1634 (N_1634,In_1073,In_95);
nor U1635 (N_1635,In_1286,In_1257);
and U1636 (N_1636,In_516,In_382);
and U1637 (N_1637,In_746,In_527);
or U1638 (N_1638,In_480,In_1072);
nor U1639 (N_1639,In_1433,In_565);
or U1640 (N_1640,In_349,In_599);
xnor U1641 (N_1641,In_54,In_1342);
or U1642 (N_1642,In_1056,In_1001);
or U1643 (N_1643,In_960,In_235);
nor U1644 (N_1644,In_789,In_1292);
and U1645 (N_1645,In_1206,In_1329);
or U1646 (N_1646,In_742,In_475);
nand U1647 (N_1647,In_886,In_409);
or U1648 (N_1648,In_348,In_1196);
or U1649 (N_1649,In_705,In_78);
and U1650 (N_1650,In_578,In_1316);
nand U1651 (N_1651,In_1374,In_1479);
or U1652 (N_1652,In_281,In_1348);
and U1653 (N_1653,In_593,In_1409);
nor U1654 (N_1654,In_850,In_827);
nor U1655 (N_1655,In_88,In_194);
or U1656 (N_1656,In_1124,In_21);
or U1657 (N_1657,In_554,In_26);
or U1658 (N_1658,In_1328,In_759);
nor U1659 (N_1659,In_1220,In_985);
nor U1660 (N_1660,In_921,In_532);
or U1661 (N_1661,In_389,In_71);
nand U1662 (N_1662,In_1081,In_1027);
or U1663 (N_1663,In_358,In_590);
or U1664 (N_1664,In_1432,In_863);
or U1665 (N_1665,In_429,In_242);
and U1666 (N_1666,In_415,In_932);
and U1667 (N_1667,In_556,In_490);
or U1668 (N_1668,In_150,In_367);
nand U1669 (N_1669,In_81,In_1467);
nand U1670 (N_1670,In_133,In_712);
nand U1671 (N_1671,In_588,In_1191);
nand U1672 (N_1672,In_1144,In_1105);
and U1673 (N_1673,In_263,In_415);
or U1674 (N_1674,In_385,In_1350);
or U1675 (N_1675,In_778,In_1010);
or U1676 (N_1676,In_1348,In_517);
nand U1677 (N_1677,In_212,In_215);
and U1678 (N_1678,In_978,In_1012);
nand U1679 (N_1679,In_1457,In_443);
and U1680 (N_1680,In_1003,In_613);
nand U1681 (N_1681,In_85,In_3);
and U1682 (N_1682,In_1258,In_377);
and U1683 (N_1683,In_1075,In_217);
nand U1684 (N_1684,In_1441,In_1431);
and U1685 (N_1685,In_901,In_252);
and U1686 (N_1686,In_1499,In_1296);
and U1687 (N_1687,In_388,In_731);
nor U1688 (N_1688,In_677,In_176);
or U1689 (N_1689,In_581,In_972);
and U1690 (N_1690,In_1191,In_1331);
xor U1691 (N_1691,In_423,In_1019);
or U1692 (N_1692,In_506,In_570);
nand U1693 (N_1693,In_1383,In_757);
or U1694 (N_1694,In_367,In_1316);
nand U1695 (N_1695,In_740,In_988);
and U1696 (N_1696,In_1043,In_1077);
and U1697 (N_1697,In_617,In_1220);
and U1698 (N_1698,In_674,In_397);
and U1699 (N_1699,In_591,In_129);
and U1700 (N_1700,In_282,In_1246);
or U1701 (N_1701,In_1207,In_586);
nor U1702 (N_1702,In_740,In_931);
nor U1703 (N_1703,In_146,In_140);
nand U1704 (N_1704,In_1433,In_1168);
nor U1705 (N_1705,In_108,In_1275);
or U1706 (N_1706,In_1391,In_1074);
xnor U1707 (N_1707,In_1396,In_1139);
or U1708 (N_1708,In_1444,In_1432);
nand U1709 (N_1709,In_660,In_125);
nor U1710 (N_1710,In_360,In_837);
nor U1711 (N_1711,In_378,In_631);
or U1712 (N_1712,In_514,In_1468);
nand U1713 (N_1713,In_756,In_1496);
or U1714 (N_1714,In_911,In_312);
nor U1715 (N_1715,In_1198,In_5);
nand U1716 (N_1716,In_1035,In_1342);
nand U1717 (N_1717,In_45,In_967);
and U1718 (N_1718,In_1437,In_1486);
or U1719 (N_1719,In_665,In_1253);
nor U1720 (N_1720,In_41,In_350);
nand U1721 (N_1721,In_1010,In_192);
and U1722 (N_1722,In_793,In_929);
or U1723 (N_1723,In_1342,In_1048);
and U1724 (N_1724,In_277,In_471);
and U1725 (N_1725,In_1168,In_1448);
or U1726 (N_1726,In_1420,In_978);
nor U1727 (N_1727,In_147,In_662);
or U1728 (N_1728,In_969,In_1040);
nand U1729 (N_1729,In_1367,In_420);
nand U1730 (N_1730,In_975,In_1038);
and U1731 (N_1731,In_467,In_1491);
nor U1732 (N_1732,In_701,In_180);
and U1733 (N_1733,In_44,In_1237);
and U1734 (N_1734,In_1356,In_629);
nor U1735 (N_1735,In_684,In_244);
nand U1736 (N_1736,In_84,In_1120);
nor U1737 (N_1737,In_701,In_836);
and U1738 (N_1738,In_485,In_1415);
and U1739 (N_1739,In_1409,In_574);
and U1740 (N_1740,In_441,In_533);
and U1741 (N_1741,In_1480,In_1060);
nand U1742 (N_1742,In_953,In_993);
nor U1743 (N_1743,In_588,In_869);
nor U1744 (N_1744,In_74,In_1095);
or U1745 (N_1745,In_1123,In_1215);
and U1746 (N_1746,In_990,In_579);
xor U1747 (N_1747,In_646,In_96);
and U1748 (N_1748,In_325,In_672);
xor U1749 (N_1749,In_540,In_949);
and U1750 (N_1750,In_56,In_260);
nand U1751 (N_1751,In_570,In_1229);
and U1752 (N_1752,In_639,In_1382);
or U1753 (N_1753,In_470,In_403);
xnor U1754 (N_1754,In_189,In_1000);
nor U1755 (N_1755,In_1357,In_547);
or U1756 (N_1756,In_160,In_396);
and U1757 (N_1757,In_1351,In_158);
and U1758 (N_1758,In_40,In_241);
or U1759 (N_1759,In_585,In_706);
nand U1760 (N_1760,In_536,In_145);
nand U1761 (N_1761,In_1066,In_812);
and U1762 (N_1762,In_1166,In_944);
or U1763 (N_1763,In_801,In_1031);
or U1764 (N_1764,In_431,In_485);
nor U1765 (N_1765,In_1251,In_419);
nor U1766 (N_1766,In_1407,In_661);
nand U1767 (N_1767,In_1173,In_10);
or U1768 (N_1768,In_1341,In_130);
nand U1769 (N_1769,In_573,In_855);
or U1770 (N_1770,In_653,In_775);
and U1771 (N_1771,In_242,In_1449);
or U1772 (N_1772,In_12,In_426);
or U1773 (N_1773,In_1433,In_1065);
nand U1774 (N_1774,In_341,In_428);
nand U1775 (N_1775,In_14,In_29);
or U1776 (N_1776,In_224,In_793);
and U1777 (N_1777,In_692,In_1497);
and U1778 (N_1778,In_1326,In_574);
nor U1779 (N_1779,In_120,In_1329);
or U1780 (N_1780,In_76,In_815);
or U1781 (N_1781,In_1366,In_806);
nand U1782 (N_1782,In_1122,In_903);
nand U1783 (N_1783,In_243,In_1101);
and U1784 (N_1784,In_953,In_1494);
and U1785 (N_1785,In_1295,In_1077);
nor U1786 (N_1786,In_71,In_529);
nor U1787 (N_1787,In_302,In_219);
nor U1788 (N_1788,In_626,In_169);
and U1789 (N_1789,In_174,In_402);
and U1790 (N_1790,In_1122,In_479);
nand U1791 (N_1791,In_35,In_569);
or U1792 (N_1792,In_1101,In_449);
or U1793 (N_1793,In_632,In_666);
nand U1794 (N_1794,In_327,In_338);
xnor U1795 (N_1795,In_381,In_605);
nand U1796 (N_1796,In_1126,In_1052);
nor U1797 (N_1797,In_709,In_579);
nand U1798 (N_1798,In_1320,In_395);
nand U1799 (N_1799,In_159,In_76);
xor U1800 (N_1800,In_736,In_226);
and U1801 (N_1801,In_1419,In_396);
and U1802 (N_1802,In_876,In_1009);
or U1803 (N_1803,In_562,In_1470);
nand U1804 (N_1804,In_190,In_331);
or U1805 (N_1805,In_966,In_860);
or U1806 (N_1806,In_928,In_500);
nand U1807 (N_1807,In_222,In_864);
and U1808 (N_1808,In_1081,In_967);
nand U1809 (N_1809,In_794,In_113);
nor U1810 (N_1810,In_902,In_38);
nor U1811 (N_1811,In_723,In_359);
nand U1812 (N_1812,In_1053,In_1423);
nand U1813 (N_1813,In_1009,In_1040);
xnor U1814 (N_1814,In_1318,In_176);
or U1815 (N_1815,In_138,In_444);
nand U1816 (N_1816,In_731,In_121);
nand U1817 (N_1817,In_1363,In_1080);
or U1818 (N_1818,In_659,In_149);
nor U1819 (N_1819,In_130,In_1033);
nor U1820 (N_1820,In_687,In_1210);
nor U1821 (N_1821,In_1045,In_1407);
or U1822 (N_1822,In_1169,In_200);
nor U1823 (N_1823,In_1023,In_1124);
and U1824 (N_1824,In_458,In_686);
nor U1825 (N_1825,In_215,In_1183);
and U1826 (N_1826,In_226,In_414);
and U1827 (N_1827,In_172,In_1128);
or U1828 (N_1828,In_208,In_1314);
nand U1829 (N_1829,In_323,In_1253);
and U1830 (N_1830,In_253,In_140);
and U1831 (N_1831,In_482,In_1061);
or U1832 (N_1832,In_1104,In_247);
and U1833 (N_1833,In_1224,In_997);
nor U1834 (N_1834,In_13,In_1368);
and U1835 (N_1835,In_1164,In_550);
and U1836 (N_1836,In_181,In_1111);
and U1837 (N_1837,In_736,In_886);
nor U1838 (N_1838,In_831,In_652);
and U1839 (N_1839,In_475,In_1279);
nor U1840 (N_1840,In_1118,In_193);
nand U1841 (N_1841,In_789,In_1127);
nor U1842 (N_1842,In_1494,In_1091);
nor U1843 (N_1843,In_740,In_272);
xnor U1844 (N_1844,In_1228,In_152);
nor U1845 (N_1845,In_1412,In_835);
nor U1846 (N_1846,In_792,In_949);
nor U1847 (N_1847,In_309,In_159);
and U1848 (N_1848,In_283,In_1053);
nor U1849 (N_1849,In_1090,In_140);
nor U1850 (N_1850,In_1311,In_673);
or U1851 (N_1851,In_1458,In_762);
and U1852 (N_1852,In_1174,In_592);
and U1853 (N_1853,In_208,In_166);
nand U1854 (N_1854,In_818,In_344);
nand U1855 (N_1855,In_1327,In_930);
nand U1856 (N_1856,In_8,In_497);
or U1857 (N_1857,In_309,In_993);
nand U1858 (N_1858,In_115,In_546);
or U1859 (N_1859,In_478,In_33);
or U1860 (N_1860,In_1466,In_498);
nor U1861 (N_1861,In_946,In_1186);
nor U1862 (N_1862,In_210,In_924);
nand U1863 (N_1863,In_1180,In_1392);
nand U1864 (N_1864,In_54,In_1159);
nand U1865 (N_1865,In_1316,In_437);
nor U1866 (N_1866,In_1283,In_901);
nor U1867 (N_1867,In_630,In_268);
or U1868 (N_1868,In_1399,In_1166);
nor U1869 (N_1869,In_674,In_56);
and U1870 (N_1870,In_169,In_1419);
nor U1871 (N_1871,In_77,In_804);
xnor U1872 (N_1872,In_884,In_663);
and U1873 (N_1873,In_1147,In_682);
nor U1874 (N_1874,In_1488,In_339);
nor U1875 (N_1875,In_1030,In_678);
nor U1876 (N_1876,In_669,In_792);
and U1877 (N_1877,In_1224,In_893);
or U1878 (N_1878,In_1169,In_733);
nand U1879 (N_1879,In_938,In_145);
and U1880 (N_1880,In_564,In_795);
or U1881 (N_1881,In_200,In_1122);
and U1882 (N_1882,In_1120,In_749);
and U1883 (N_1883,In_1086,In_366);
nor U1884 (N_1884,In_1482,In_571);
nor U1885 (N_1885,In_1450,In_1088);
or U1886 (N_1886,In_775,In_437);
or U1887 (N_1887,In_1177,In_875);
nand U1888 (N_1888,In_1251,In_707);
or U1889 (N_1889,In_1223,In_312);
nand U1890 (N_1890,In_872,In_561);
nor U1891 (N_1891,In_868,In_230);
nand U1892 (N_1892,In_1440,In_637);
and U1893 (N_1893,In_1139,In_1289);
or U1894 (N_1894,In_1334,In_755);
or U1895 (N_1895,In_337,In_335);
xor U1896 (N_1896,In_1273,In_1442);
nor U1897 (N_1897,In_534,In_1258);
nor U1898 (N_1898,In_1289,In_1067);
nand U1899 (N_1899,In_669,In_840);
nand U1900 (N_1900,In_1016,In_630);
and U1901 (N_1901,In_1328,In_1213);
and U1902 (N_1902,In_983,In_1479);
and U1903 (N_1903,In_1226,In_504);
nor U1904 (N_1904,In_1185,In_467);
nor U1905 (N_1905,In_1006,In_458);
or U1906 (N_1906,In_1365,In_577);
or U1907 (N_1907,In_201,In_1189);
or U1908 (N_1908,In_1126,In_856);
or U1909 (N_1909,In_1190,In_86);
nand U1910 (N_1910,In_1273,In_1435);
and U1911 (N_1911,In_414,In_1289);
or U1912 (N_1912,In_587,In_542);
nor U1913 (N_1913,In_665,In_1381);
or U1914 (N_1914,In_345,In_891);
and U1915 (N_1915,In_69,In_555);
or U1916 (N_1916,In_617,In_281);
and U1917 (N_1917,In_175,In_938);
or U1918 (N_1918,In_64,In_1169);
or U1919 (N_1919,In_1202,In_1321);
or U1920 (N_1920,In_1220,In_308);
nand U1921 (N_1921,In_559,In_1160);
nor U1922 (N_1922,In_997,In_947);
xor U1923 (N_1923,In_234,In_1001);
or U1924 (N_1924,In_762,In_591);
nand U1925 (N_1925,In_221,In_222);
and U1926 (N_1926,In_1446,In_482);
or U1927 (N_1927,In_1309,In_747);
nand U1928 (N_1928,In_521,In_1245);
or U1929 (N_1929,In_778,In_482);
nand U1930 (N_1930,In_823,In_832);
nand U1931 (N_1931,In_206,In_577);
and U1932 (N_1932,In_434,In_1340);
nor U1933 (N_1933,In_1306,In_1396);
nor U1934 (N_1934,In_1104,In_565);
or U1935 (N_1935,In_1212,In_952);
or U1936 (N_1936,In_1462,In_1118);
and U1937 (N_1937,In_787,In_613);
or U1938 (N_1938,In_1295,In_1448);
nand U1939 (N_1939,In_1364,In_620);
and U1940 (N_1940,In_1482,In_996);
xnor U1941 (N_1941,In_981,In_425);
nor U1942 (N_1942,In_1012,In_987);
nand U1943 (N_1943,In_142,In_302);
nand U1944 (N_1944,In_1235,In_126);
and U1945 (N_1945,In_109,In_768);
nand U1946 (N_1946,In_782,In_1183);
and U1947 (N_1947,In_1087,In_156);
or U1948 (N_1948,In_934,In_874);
or U1949 (N_1949,In_1337,In_1410);
or U1950 (N_1950,In_441,In_239);
and U1951 (N_1951,In_1160,In_902);
nor U1952 (N_1952,In_521,In_1418);
nor U1953 (N_1953,In_320,In_808);
nor U1954 (N_1954,In_395,In_201);
or U1955 (N_1955,In_882,In_1327);
xor U1956 (N_1956,In_229,In_1383);
nand U1957 (N_1957,In_1092,In_342);
nand U1958 (N_1958,In_578,In_743);
nand U1959 (N_1959,In_698,In_574);
nand U1960 (N_1960,In_55,In_721);
or U1961 (N_1961,In_391,In_435);
and U1962 (N_1962,In_643,In_860);
nand U1963 (N_1963,In_936,In_700);
nand U1964 (N_1964,In_1215,In_535);
or U1965 (N_1965,In_251,In_758);
nor U1966 (N_1966,In_351,In_1335);
and U1967 (N_1967,In_1172,In_621);
or U1968 (N_1968,In_632,In_368);
nor U1969 (N_1969,In_592,In_750);
and U1970 (N_1970,In_1034,In_1313);
nand U1971 (N_1971,In_1197,In_260);
nor U1972 (N_1972,In_441,In_569);
or U1973 (N_1973,In_165,In_239);
or U1974 (N_1974,In_1012,In_893);
or U1975 (N_1975,In_36,In_70);
nor U1976 (N_1976,In_487,In_1322);
or U1977 (N_1977,In_644,In_103);
nand U1978 (N_1978,In_540,In_628);
and U1979 (N_1979,In_718,In_396);
and U1980 (N_1980,In_140,In_1437);
nand U1981 (N_1981,In_937,In_1027);
and U1982 (N_1982,In_791,In_99);
nor U1983 (N_1983,In_597,In_1124);
nor U1984 (N_1984,In_879,In_292);
xnor U1985 (N_1985,In_1495,In_1232);
nand U1986 (N_1986,In_129,In_384);
xnor U1987 (N_1987,In_166,In_382);
and U1988 (N_1988,In_43,In_79);
nor U1989 (N_1989,In_653,In_67);
and U1990 (N_1990,In_416,In_1041);
nor U1991 (N_1991,In_181,In_662);
nand U1992 (N_1992,In_588,In_1442);
nor U1993 (N_1993,In_1130,In_370);
nor U1994 (N_1994,In_327,In_1212);
or U1995 (N_1995,In_942,In_523);
or U1996 (N_1996,In_790,In_1466);
or U1997 (N_1997,In_1351,In_1224);
xor U1998 (N_1998,In_176,In_688);
nand U1999 (N_1999,In_357,In_687);
nand U2000 (N_2000,In_534,In_851);
nand U2001 (N_2001,In_1086,In_1275);
nand U2002 (N_2002,In_19,In_406);
or U2003 (N_2003,In_1496,In_1053);
and U2004 (N_2004,In_719,In_1150);
xor U2005 (N_2005,In_1340,In_751);
and U2006 (N_2006,In_494,In_1478);
xnor U2007 (N_2007,In_237,In_1209);
and U2008 (N_2008,In_621,In_1356);
and U2009 (N_2009,In_586,In_1256);
or U2010 (N_2010,In_691,In_519);
nand U2011 (N_2011,In_597,In_861);
and U2012 (N_2012,In_323,In_939);
and U2013 (N_2013,In_1393,In_1148);
nand U2014 (N_2014,In_1342,In_449);
xnor U2015 (N_2015,In_1029,In_148);
nor U2016 (N_2016,In_1150,In_468);
nand U2017 (N_2017,In_499,In_732);
nor U2018 (N_2018,In_359,In_362);
and U2019 (N_2019,In_4,In_1147);
nand U2020 (N_2020,In_1135,In_322);
nand U2021 (N_2021,In_1301,In_7);
nand U2022 (N_2022,In_721,In_1176);
or U2023 (N_2023,In_1292,In_1097);
and U2024 (N_2024,In_1233,In_615);
nand U2025 (N_2025,In_1203,In_138);
nand U2026 (N_2026,In_128,In_6);
and U2027 (N_2027,In_1311,In_1383);
nand U2028 (N_2028,In_56,In_1499);
or U2029 (N_2029,In_475,In_566);
nand U2030 (N_2030,In_414,In_260);
nand U2031 (N_2031,In_1356,In_1145);
nor U2032 (N_2032,In_565,In_835);
nand U2033 (N_2033,In_866,In_1102);
or U2034 (N_2034,In_1356,In_501);
and U2035 (N_2035,In_1266,In_346);
or U2036 (N_2036,In_1039,In_883);
nand U2037 (N_2037,In_595,In_25);
nand U2038 (N_2038,In_1150,In_929);
nor U2039 (N_2039,In_250,In_440);
or U2040 (N_2040,In_1086,In_1013);
or U2041 (N_2041,In_40,In_1338);
or U2042 (N_2042,In_1069,In_1144);
or U2043 (N_2043,In_351,In_829);
nand U2044 (N_2044,In_810,In_972);
nor U2045 (N_2045,In_205,In_891);
or U2046 (N_2046,In_1324,In_43);
or U2047 (N_2047,In_1436,In_1175);
nor U2048 (N_2048,In_49,In_1091);
nand U2049 (N_2049,In_306,In_112);
nand U2050 (N_2050,In_911,In_1220);
nand U2051 (N_2051,In_111,In_1221);
and U2052 (N_2052,In_1136,In_425);
xnor U2053 (N_2053,In_569,In_97);
nand U2054 (N_2054,In_952,In_501);
and U2055 (N_2055,In_1256,In_1396);
and U2056 (N_2056,In_211,In_787);
and U2057 (N_2057,In_1001,In_480);
or U2058 (N_2058,In_1023,In_847);
or U2059 (N_2059,In_804,In_1158);
nand U2060 (N_2060,In_867,In_1187);
and U2061 (N_2061,In_1217,In_1201);
nor U2062 (N_2062,In_1327,In_643);
and U2063 (N_2063,In_18,In_944);
nand U2064 (N_2064,In_829,In_143);
nor U2065 (N_2065,In_1089,In_387);
nand U2066 (N_2066,In_1272,In_337);
nor U2067 (N_2067,In_725,In_634);
xnor U2068 (N_2068,In_1236,In_327);
nor U2069 (N_2069,In_731,In_406);
or U2070 (N_2070,In_1188,In_578);
and U2071 (N_2071,In_1254,In_1017);
and U2072 (N_2072,In_909,In_19);
or U2073 (N_2073,In_1029,In_804);
nor U2074 (N_2074,In_194,In_866);
nor U2075 (N_2075,In_92,In_55);
and U2076 (N_2076,In_1197,In_130);
nand U2077 (N_2077,In_1195,In_600);
nand U2078 (N_2078,In_175,In_99);
or U2079 (N_2079,In_427,In_180);
or U2080 (N_2080,In_1498,In_1404);
nor U2081 (N_2081,In_1166,In_1236);
and U2082 (N_2082,In_1182,In_249);
and U2083 (N_2083,In_687,In_895);
nor U2084 (N_2084,In_1238,In_601);
or U2085 (N_2085,In_928,In_885);
and U2086 (N_2086,In_334,In_935);
nor U2087 (N_2087,In_488,In_855);
nor U2088 (N_2088,In_1204,In_985);
and U2089 (N_2089,In_379,In_1061);
or U2090 (N_2090,In_343,In_1227);
nand U2091 (N_2091,In_1093,In_1021);
nand U2092 (N_2092,In_429,In_471);
and U2093 (N_2093,In_88,In_304);
nand U2094 (N_2094,In_682,In_591);
nor U2095 (N_2095,In_1190,In_1195);
nand U2096 (N_2096,In_180,In_1419);
nand U2097 (N_2097,In_371,In_179);
and U2098 (N_2098,In_825,In_968);
or U2099 (N_2099,In_1476,In_372);
nand U2100 (N_2100,In_1351,In_208);
or U2101 (N_2101,In_1481,In_1174);
and U2102 (N_2102,In_763,In_550);
nand U2103 (N_2103,In_318,In_321);
nor U2104 (N_2104,In_537,In_1179);
nor U2105 (N_2105,In_1371,In_1291);
nand U2106 (N_2106,In_1305,In_1252);
or U2107 (N_2107,In_76,In_455);
nand U2108 (N_2108,In_911,In_1434);
and U2109 (N_2109,In_1397,In_903);
or U2110 (N_2110,In_811,In_841);
xor U2111 (N_2111,In_632,In_1133);
nor U2112 (N_2112,In_1491,In_959);
nor U2113 (N_2113,In_1042,In_3);
and U2114 (N_2114,In_809,In_25);
or U2115 (N_2115,In_731,In_1488);
and U2116 (N_2116,In_176,In_774);
nand U2117 (N_2117,In_538,In_823);
nand U2118 (N_2118,In_1036,In_489);
nor U2119 (N_2119,In_40,In_696);
and U2120 (N_2120,In_314,In_1398);
and U2121 (N_2121,In_862,In_1352);
nor U2122 (N_2122,In_1207,In_1060);
or U2123 (N_2123,In_647,In_123);
nor U2124 (N_2124,In_785,In_1040);
nand U2125 (N_2125,In_1427,In_220);
and U2126 (N_2126,In_790,In_426);
and U2127 (N_2127,In_120,In_51);
nand U2128 (N_2128,In_1352,In_370);
and U2129 (N_2129,In_742,In_708);
xnor U2130 (N_2130,In_1041,In_957);
nor U2131 (N_2131,In_579,In_225);
nand U2132 (N_2132,In_925,In_1432);
and U2133 (N_2133,In_7,In_654);
and U2134 (N_2134,In_483,In_477);
nand U2135 (N_2135,In_1403,In_791);
or U2136 (N_2136,In_1407,In_554);
nor U2137 (N_2137,In_41,In_1150);
nor U2138 (N_2138,In_870,In_1185);
and U2139 (N_2139,In_785,In_1390);
and U2140 (N_2140,In_698,In_566);
nor U2141 (N_2141,In_233,In_1095);
nor U2142 (N_2142,In_960,In_995);
nand U2143 (N_2143,In_134,In_1024);
and U2144 (N_2144,In_714,In_1387);
or U2145 (N_2145,In_1279,In_978);
nor U2146 (N_2146,In_481,In_1275);
xnor U2147 (N_2147,In_341,In_1145);
or U2148 (N_2148,In_851,In_603);
nor U2149 (N_2149,In_998,In_126);
and U2150 (N_2150,In_1174,In_1250);
nor U2151 (N_2151,In_958,In_45);
nor U2152 (N_2152,In_137,In_921);
or U2153 (N_2153,In_318,In_693);
or U2154 (N_2154,In_698,In_263);
and U2155 (N_2155,In_71,In_109);
nor U2156 (N_2156,In_43,In_1038);
and U2157 (N_2157,In_199,In_1281);
nand U2158 (N_2158,In_106,In_1152);
nor U2159 (N_2159,In_1217,In_1312);
nand U2160 (N_2160,In_614,In_253);
and U2161 (N_2161,In_911,In_517);
nand U2162 (N_2162,In_367,In_296);
and U2163 (N_2163,In_30,In_916);
and U2164 (N_2164,In_827,In_873);
xor U2165 (N_2165,In_598,In_563);
nor U2166 (N_2166,In_441,In_318);
and U2167 (N_2167,In_401,In_1198);
nand U2168 (N_2168,In_607,In_426);
and U2169 (N_2169,In_1348,In_333);
and U2170 (N_2170,In_476,In_1251);
nor U2171 (N_2171,In_1091,In_385);
nor U2172 (N_2172,In_149,In_296);
or U2173 (N_2173,In_666,In_927);
nand U2174 (N_2174,In_646,In_579);
nor U2175 (N_2175,In_524,In_841);
or U2176 (N_2176,In_156,In_1463);
and U2177 (N_2177,In_1249,In_466);
and U2178 (N_2178,In_1260,In_383);
nand U2179 (N_2179,In_729,In_637);
or U2180 (N_2180,In_1402,In_652);
xnor U2181 (N_2181,In_35,In_819);
nand U2182 (N_2182,In_1350,In_1381);
nor U2183 (N_2183,In_592,In_849);
or U2184 (N_2184,In_204,In_863);
or U2185 (N_2185,In_229,In_1209);
and U2186 (N_2186,In_1255,In_1308);
and U2187 (N_2187,In_1041,In_1252);
nor U2188 (N_2188,In_188,In_181);
nand U2189 (N_2189,In_1189,In_839);
nand U2190 (N_2190,In_417,In_537);
and U2191 (N_2191,In_670,In_159);
or U2192 (N_2192,In_292,In_1154);
or U2193 (N_2193,In_814,In_556);
nand U2194 (N_2194,In_1234,In_992);
nor U2195 (N_2195,In_31,In_561);
or U2196 (N_2196,In_1111,In_754);
nand U2197 (N_2197,In_207,In_1374);
and U2198 (N_2198,In_789,In_549);
or U2199 (N_2199,In_703,In_181);
or U2200 (N_2200,In_850,In_343);
nand U2201 (N_2201,In_59,In_951);
xor U2202 (N_2202,In_1461,In_1021);
nand U2203 (N_2203,In_27,In_142);
xnor U2204 (N_2204,In_1446,In_1450);
and U2205 (N_2205,In_583,In_416);
nand U2206 (N_2206,In_924,In_541);
nand U2207 (N_2207,In_1346,In_404);
and U2208 (N_2208,In_57,In_478);
and U2209 (N_2209,In_1057,In_1003);
nand U2210 (N_2210,In_391,In_561);
and U2211 (N_2211,In_1122,In_469);
or U2212 (N_2212,In_1139,In_1108);
nor U2213 (N_2213,In_1230,In_365);
nand U2214 (N_2214,In_171,In_1121);
and U2215 (N_2215,In_843,In_1483);
or U2216 (N_2216,In_1291,In_451);
and U2217 (N_2217,In_1419,In_1267);
nand U2218 (N_2218,In_789,In_67);
and U2219 (N_2219,In_1428,In_1312);
nor U2220 (N_2220,In_519,In_291);
nand U2221 (N_2221,In_173,In_504);
and U2222 (N_2222,In_355,In_39);
or U2223 (N_2223,In_264,In_120);
or U2224 (N_2224,In_726,In_10);
nor U2225 (N_2225,In_435,In_1308);
or U2226 (N_2226,In_1440,In_413);
nand U2227 (N_2227,In_99,In_122);
and U2228 (N_2228,In_665,In_1282);
xor U2229 (N_2229,In_625,In_1419);
nor U2230 (N_2230,In_990,In_122);
and U2231 (N_2231,In_1367,In_785);
xor U2232 (N_2232,In_686,In_226);
or U2233 (N_2233,In_127,In_86);
or U2234 (N_2234,In_510,In_765);
nor U2235 (N_2235,In_496,In_653);
nand U2236 (N_2236,In_54,In_374);
and U2237 (N_2237,In_34,In_1242);
nand U2238 (N_2238,In_272,In_1283);
nand U2239 (N_2239,In_1415,In_1064);
or U2240 (N_2240,In_1224,In_158);
and U2241 (N_2241,In_780,In_1437);
or U2242 (N_2242,In_1400,In_108);
and U2243 (N_2243,In_1142,In_1404);
or U2244 (N_2244,In_756,In_178);
and U2245 (N_2245,In_162,In_155);
and U2246 (N_2246,In_441,In_361);
nor U2247 (N_2247,In_558,In_1427);
and U2248 (N_2248,In_1363,In_607);
nor U2249 (N_2249,In_182,In_12);
and U2250 (N_2250,In_375,In_984);
or U2251 (N_2251,In_449,In_1174);
and U2252 (N_2252,In_37,In_322);
nor U2253 (N_2253,In_640,In_920);
nand U2254 (N_2254,In_548,In_735);
or U2255 (N_2255,In_1155,In_529);
nor U2256 (N_2256,In_160,In_819);
or U2257 (N_2257,In_214,In_1476);
nor U2258 (N_2258,In_623,In_1389);
and U2259 (N_2259,In_882,In_946);
or U2260 (N_2260,In_577,In_665);
or U2261 (N_2261,In_1369,In_1179);
xnor U2262 (N_2262,In_114,In_18);
and U2263 (N_2263,In_1245,In_291);
and U2264 (N_2264,In_353,In_573);
nand U2265 (N_2265,In_48,In_592);
or U2266 (N_2266,In_632,In_1421);
nand U2267 (N_2267,In_276,In_8);
or U2268 (N_2268,In_1301,In_1180);
and U2269 (N_2269,In_973,In_1387);
nor U2270 (N_2270,In_453,In_224);
or U2271 (N_2271,In_90,In_569);
nor U2272 (N_2272,In_540,In_978);
nand U2273 (N_2273,In_1005,In_217);
nand U2274 (N_2274,In_57,In_1058);
nor U2275 (N_2275,In_1403,In_416);
and U2276 (N_2276,In_729,In_1483);
and U2277 (N_2277,In_903,In_689);
nand U2278 (N_2278,In_872,In_991);
and U2279 (N_2279,In_446,In_1322);
and U2280 (N_2280,In_731,In_849);
or U2281 (N_2281,In_996,In_429);
and U2282 (N_2282,In_1015,In_1040);
nor U2283 (N_2283,In_1209,In_1030);
or U2284 (N_2284,In_316,In_988);
nand U2285 (N_2285,In_877,In_25);
or U2286 (N_2286,In_962,In_1212);
nor U2287 (N_2287,In_739,In_1250);
and U2288 (N_2288,In_1377,In_1174);
nand U2289 (N_2289,In_226,In_933);
and U2290 (N_2290,In_12,In_808);
and U2291 (N_2291,In_1370,In_1430);
or U2292 (N_2292,In_490,In_815);
and U2293 (N_2293,In_1434,In_1019);
or U2294 (N_2294,In_271,In_290);
and U2295 (N_2295,In_1379,In_790);
and U2296 (N_2296,In_186,In_614);
or U2297 (N_2297,In_1395,In_387);
nor U2298 (N_2298,In_1487,In_78);
or U2299 (N_2299,In_1111,In_942);
nand U2300 (N_2300,In_1403,In_836);
nand U2301 (N_2301,In_597,In_296);
or U2302 (N_2302,In_1218,In_38);
nand U2303 (N_2303,In_314,In_1266);
and U2304 (N_2304,In_1065,In_938);
and U2305 (N_2305,In_281,In_990);
nand U2306 (N_2306,In_565,In_221);
nor U2307 (N_2307,In_1280,In_768);
and U2308 (N_2308,In_562,In_397);
and U2309 (N_2309,In_1281,In_1135);
nand U2310 (N_2310,In_946,In_49);
nor U2311 (N_2311,In_1069,In_1461);
nand U2312 (N_2312,In_1206,In_375);
or U2313 (N_2313,In_246,In_43);
or U2314 (N_2314,In_657,In_978);
and U2315 (N_2315,In_557,In_860);
or U2316 (N_2316,In_984,In_1276);
nor U2317 (N_2317,In_809,In_1340);
or U2318 (N_2318,In_1187,In_1036);
and U2319 (N_2319,In_131,In_682);
nor U2320 (N_2320,In_807,In_1127);
and U2321 (N_2321,In_153,In_573);
or U2322 (N_2322,In_1489,In_221);
nand U2323 (N_2323,In_572,In_1322);
and U2324 (N_2324,In_792,In_231);
nor U2325 (N_2325,In_203,In_392);
nand U2326 (N_2326,In_181,In_161);
nand U2327 (N_2327,In_1305,In_568);
nor U2328 (N_2328,In_1258,In_721);
nor U2329 (N_2329,In_1116,In_429);
nand U2330 (N_2330,In_180,In_1066);
or U2331 (N_2331,In_163,In_500);
and U2332 (N_2332,In_684,In_1361);
or U2333 (N_2333,In_1168,In_1483);
and U2334 (N_2334,In_1295,In_432);
nor U2335 (N_2335,In_522,In_1150);
or U2336 (N_2336,In_1322,In_733);
xnor U2337 (N_2337,In_980,In_1136);
and U2338 (N_2338,In_227,In_1015);
nor U2339 (N_2339,In_607,In_482);
nor U2340 (N_2340,In_553,In_994);
or U2341 (N_2341,In_426,In_1356);
and U2342 (N_2342,In_1006,In_1162);
and U2343 (N_2343,In_284,In_931);
nor U2344 (N_2344,In_620,In_1150);
or U2345 (N_2345,In_375,In_164);
nor U2346 (N_2346,In_324,In_60);
and U2347 (N_2347,In_53,In_1289);
nand U2348 (N_2348,In_1156,In_683);
nor U2349 (N_2349,In_1185,In_123);
or U2350 (N_2350,In_1227,In_1147);
nand U2351 (N_2351,In_266,In_1168);
nand U2352 (N_2352,In_702,In_689);
nor U2353 (N_2353,In_337,In_1132);
and U2354 (N_2354,In_1378,In_1412);
nor U2355 (N_2355,In_1265,In_724);
nor U2356 (N_2356,In_1347,In_680);
or U2357 (N_2357,In_315,In_1308);
and U2358 (N_2358,In_1025,In_894);
or U2359 (N_2359,In_1469,In_1155);
nand U2360 (N_2360,In_11,In_1395);
nor U2361 (N_2361,In_774,In_850);
nor U2362 (N_2362,In_467,In_506);
nor U2363 (N_2363,In_194,In_492);
or U2364 (N_2364,In_1358,In_1275);
nor U2365 (N_2365,In_670,In_19);
and U2366 (N_2366,In_542,In_537);
or U2367 (N_2367,In_709,In_1118);
nand U2368 (N_2368,In_948,In_81);
and U2369 (N_2369,In_950,In_1316);
nor U2370 (N_2370,In_1314,In_1498);
nand U2371 (N_2371,In_488,In_1253);
or U2372 (N_2372,In_1170,In_371);
nor U2373 (N_2373,In_742,In_1475);
or U2374 (N_2374,In_749,In_47);
and U2375 (N_2375,In_206,In_255);
nor U2376 (N_2376,In_595,In_1183);
nor U2377 (N_2377,In_303,In_244);
nand U2378 (N_2378,In_1110,In_355);
nand U2379 (N_2379,In_1498,In_924);
and U2380 (N_2380,In_1221,In_1296);
and U2381 (N_2381,In_992,In_54);
nand U2382 (N_2382,In_1268,In_81);
and U2383 (N_2383,In_1113,In_726);
nand U2384 (N_2384,In_595,In_690);
or U2385 (N_2385,In_1425,In_771);
or U2386 (N_2386,In_525,In_745);
nor U2387 (N_2387,In_981,In_680);
nor U2388 (N_2388,In_30,In_659);
and U2389 (N_2389,In_853,In_203);
and U2390 (N_2390,In_802,In_538);
nor U2391 (N_2391,In_335,In_102);
nor U2392 (N_2392,In_874,In_1163);
nor U2393 (N_2393,In_453,In_536);
nand U2394 (N_2394,In_26,In_1183);
nand U2395 (N_2395,In_601,In_1326);
and U2396 (N_2396,In_1247,In_308);
and U2397 (N_2397,In_1189,In_627);
and U2398 (N_2398,In_481,In_1340);
or U2399 (N_2399,In_854,In_578);
or U2400 (N_2400,In_197,In_890);
and U2401 (N_2401,In_643,In_1256);
and U2402 (N_2402,In_1355,In_320);
nand U2403 (N_2403,In_1185,In_1472);
nor U2404 (N_2404,In_869,In_1068);
nand U2405 (N_2405,In_864,In_524);
or U2406 (N_2406,In_364,In_949);
nor U2407 (N_2407,In_471,In_1307);
nand U2408 (N_2408,In_921,In_336);
nor U2409 (N_2409,In_53,In_1008);
and U2410 (N_2410,In_171,In_472);
and U2411 (N_2411,In_1347,In_1024);
or U2412 (N_2412,In_1006,In_1118);
and U2413 (N_2413,In_1380,In_738);
nor U2414 (N_2414,In_21,In_1213);
and U2415 (N_2415,In_661,In_1375);
and U2416 (N_2416,In_1196,In_899);
and U2417 (N_2417,In_650,In_391);
nand U2418 (N_2418,In_806,In_849);
nor U2419 (N_2419,In_346,In_955);
nand U2420 (N_2420,In_1289,In_1350);
and U2421 (N_2421,In_1198,In_779);
nand U2422 (N_2422,In_866,In_1297);
nand U2423 (N_2423,In_1342,In_901);
nand U2424 (N_2424,In_841,In_1436);
or U2425 (N_2425,In_41,In_79);
nor U2426 (N_2426,In_717,In_1258);
and U2427 (N_2427,In_1159,In_298);
or U2428 (N_2428,In_1201,In_480);
and U2429 (N_2429,In_233,In_966);
nor U2430 (N_2430,In_1075,In_1228);
or U2431 (N_2431,In_575,In_1309);
and U2432 (N_2432,In_165,In_129);
and U2433 (N_2433,In_661,In_1488);
and U2434 (N_2434,In_1316,In_62);
or U2435 (N_2435,In_457,In_285);
nor U2436 (N_2436,In_675,In_193);
and U2437 (N_2437,In_671,In_961);
and U2438 (N_2438,In_1120,In_1315);
and U2439 (N_2439,In_1427,In_717);
nor U2440 (N_2440,In_543,In_1058);
and U2441 (N_2441,In_585,In_1251);
nand U2442 (N_2442,In_756,In_1492);
nor U2443 (N_2443,In_329,In_146);
or U2444 (N_2444,In_181,In_1272);
nor U2445 (N_2445,In_817,In_635);
and U2446 (N_2446,In_778,In_1221);
nor U2447 (N_2447,In_422,In_130);
or U2448 (N_2448,In_1280,In_893);
or U2449 (N_2449,In_1028,In_268);
nor U2450 (N_2450,In_1187,In_113);
nor U2451 (N_2451,In_1429,In_1499);
or U2452 (N_2452,In_881,In_843);
nor U2453 (N_2453,In_1289,In_69);
or U2454 (N_2454,In_361,In_1049);
or U2455 (N_2455,In_200,In_1340);
and U2456 (N_2456,In_885,In_490);
or U2457 (N_2457,In_1,In_648);
and U2458 (N_2458,In_1069,In_1050);
nor U2459 (N_2459,In_287,In_1210);
nand U2460 (N_2460,In_598,In_324);
or U2461 (N_2461,In_1038,In_833);
and U2462 (N_2462,In_1331,In_37);
or U2463 (N_2463,In_883,In_1286);
or U2464 (N_2464,In_155,In_1402);
nor U2465 (N_2465,In_1420,In_304);
and U2466 (N_2466,In_366,In_927);
or U2467 (N_2467,In_1331,In_38);
nor U2468 (N_2468,In_1426,In_284);
and U2469 (N_2469,In_1160,In_342);
nor U2470 (N_2470,In_260,In_832);
nand U2471 (N_2471,In_273,In_521);
or U2472 (N_2472,In_1336,In_368);
or U2473 (N_2473,In_1355,In_275);
or U2474 (N_2474,In_996,In_220);
nor U2475 (N_2475,In_313,In_229);
or U2476 (N_2476,In_721,In_1447);
nand U2477 (N_2477,In_902,In_381);
nand U2478 (N_2478,In_156,In_622);
nand U2479 (N_2479,In_1247,In_950);
or U2480 (N_2480,In_1012,In_263);
and U2481 (N_2481,In_1422,In_613);
or U2482 (N_2482,In_1273,In_162);
nor U2483 (N_2483,In_373,In_1467);
nor U2484 (N_2484,In_1433,In_1125);
or U2485 (N_2485,In_781,In_1113);
nor U2486 (N_2486,In_1055,In_1162);
nand U2487 (N_2487,In_734,In_780);
nor U2488 (N_2488,In_1254,In_81);
and U2489 (N_2489,In_937,In_892);
or U2490 (N_2490,In_472,In_809);
or U2491 (N_2491,In_978,In_1228);
nand U2492 (N_2492,In_611,In_1038);
and U2493 (N_2493,In_652,In_1084);
nor U2494 (N_2494,In_537,In_299);
nor U2495 (N_2495,In_814,In_141);
and U2496 (N_2496,In_546,In_191);
nor U2497 (N_2497,In_828,In_238);
and U2498 (N_2498,In_1461,In_760);
or U2499 (N_2499,In_1008,In_917);
and U2500 (N_2500,In_973,In_533);
nor U2501 (N_2501,In_13,In_961);
nor U2502 (N_2502,In_1405,In_15);
and U2503 (N_2503,In_395,In_97);
nor U2504 (N_2504,In_8,In_853);
xnor U2505 (N_2505,In_1142,In_448);
nand U2506 (N_2506,In_991,In_1254);
nor U2507 (N_2507,In_937,In_31);
or U2508 (N_2508,In_998,In_513);
xor U2509 (N_2509,In_383,In_948);
xor U2510 (N_2510,In_1008,In_895);
nor U2511 (N_2511,In_1080,In_458);
nor U2512 (N_2512,In_850,In_1071);
or U2513 (N_2513,In_1341,In_414);
or U2514 (N_2514,In_356,In_1480);
nand U2515 (N_2515,In_841,In_45);
and U2516 (N_2516,In_462,In_369);
or U2517 (N_2517,In_1302,In_1455);
and U2518 (N_2518,In_1024,In_1307);
or U2519 (N_2519,In_670,In_833);
and U2520 (N_2520,In_1429,In_536);
nor U2521 (N_2521,In_1276,In_321);
nand U2522 (N_2522,In_944,In_1023);
nand U2523 (N_2523,In_1000,In_22);
or U2524 (N_2524,In_824,In_323);
and U2525 (N_2525,In_1442,In_148);
and U2526 (N_2526,In_183,In_621);
and U2527 (N_2527,In_72,In_315);
nand U2528 (N_2528,In_1265,In_380);
xor U2529 (N_2529,In_504,In_1133);
xor U2530 (N_2530,In_927,In_433);
and U2531 (N_2531,In_660,In_1190);
nand U2532 (N_2532,In_581,In_677);
nor U2533 (N_2533,In_786,In_96);
or U2534 (N_2534,In_1069,In_1217);
nor U2535 (N_2535,In_1380,In_514);
nand U2536 (N_2536,In_885,In_1223);
and U2537 (N_2537,In_87,In_136);
and U2538 (N_2538,In_541,In_1063);
or U2539 (N_2539,In_946,In_204);
and U2540 (N_2540,In_370,In_1028);
nor U2541 (N_2541,In_182,In_1372);
nand U2542 (N_2542,In_381,In_235);
nand U2543 (N_2543,In_842,In_74);
and U2544 (N_2544,In_699,In_1249);
nand U2545 (N_2545,In_1432,In_578);
nor U2546 (N_2546,In_1407,In_399);
or U2547 (N_2547,In_931,In_264);
nand U2548 (N_2548,In_786,In_324);
or U2549 (N_2549,In_1484,In_1489);
nand U2550 (N_2550,In_512,In_1475);
nand U2551 (N_2551,In_1176,In_930);
and U2552 (N_2552,In_17,In_275);
nand U2553 (N_2553,In_1261,In_217);
or U2554 (N_2554,In_89,In_729);
nand U2555 (N_2555,In_913,In_131);
and U2556 (N_2556,In_1315,In_1187);
or U2557 (N_2557,In_1438,In_565);
nor U2558 (N_2558,In_344,In_963);
or U2559 (N_2559,In_1456,In_718);
nand U2560 (N_2560,In_524,In_216);
and U2561 (N_2561,In_790,In_297);
and U2562 (N_2562,In_208,In_1170);
and U2563 (N_2563,In_891,In_35);
nor U2564 (N_2564,In_997,In_639);
nand U2565 (N_2565,In_382,In_658);
nand U2566 (N_2566,In_1318,In_621);
nor U2567 (N_2567,In_26,In_70);
or U2568 (N_2568,In_561,In_774);
and U2569 (N_2569,In_731,In_915);
or U2570 (N_2570,In_1045,In_748);
nor U2571 (N_2571,In_330,In_367);
or U2572 (N_2572,In_644,In_438);
nor U2573 (N_2573,In_1098,In_1206);
nand U2574 (N_2574,In_485,In_577);
nor U2575 (N_2575,In_742,In_784);
nor U2576 (N_2576,In_647,In_1319);
nor U2577 (N_2577,In_76,In_900);
nand U2578 (N_2578,In_1254,In_321);
nor U2579 (N_2579,In_987,In_936);
or U2580 (N_2580,In_1329,In_482);
or U2581 (N_2581,In_482,In_665);
nor U2582 (N_2582,In_986,In_1383);
nand U2583 (N_2583,In_119,In_1270);
nor U2584 (N_2584,In_288,In_833);
and U2585 (N_2585,In_1338,In_542);
nand U2586 (N_2586,In_1299,In_1495);
or U2587 (N_2587,In_208,In_809);
nor U2588 (N_2588,In_273,In_548);
or U2589 (N_2589,In_737,In_53);
nor U2590 (N_2590,In_209,In_546);
and U2591 (N_2591,In_1090,In_821);
and U2592 (N_2592,In_85,In_296);
nor U2593 (N_2593,In_1475,In_1062);
or U2594 (N_2594,In_753,In_1353);
nand U2595 (N_2595,In_461,In_1497);
or U2596 (N_2596,In_10,In_708);
and U2597 (N_2597,In_1152,In_556);
nor U2598 (N_2598,In_962,In_990);
and U2599 (N_2599,In_651,In_275);
or U2600 (N_2600,In_274,In_1123);
and U2601 (N_2601,In_1414,In_1485);
nand U2602 (N_2602,In_1302,In_1072);
nor U2603 (N_2603,In_1176,In_1014);
and U2604 (N_2604,In_1158,In_1020);
nor U2605 (N_2605,In_1147,In_1265);
xor U2606 (N_2606,In_538,In_639);
nor U2607 (N_2607,In_1143,In_502);
and U2608 (N_2608,In_5,In_984);
nand U2609 (N_2609,In_766,In_484);
and U2610 (N_2610,In_1063,In_862);
or U2611 (N_2611,In_686,In_705);
or U2612 (N_2612,In_922,In_731);
nand U2613 (N_2613,In_31,In_840);
or U2614 (N_2614,In_761,In_1239);
nand U2615 (N_2615,In_546,In_1440);
nor U2616 (N_2616,In_280,In_1250);
and U2617 (N_2617,In_541,In_1198);
nand U2618 (N_2618,In_404,In_1228);
nand U2619 (N_2619,In_389,In_172);
or U2620 (N_2620,In_455,In_776);
or U2621 (N_2621,In_1415,In_745);
nor U2622 (N_2622,In_1124,In_301);
nand U2623 (N_2623,In_1378,In_164);
nor U2624 (N_2624,In_1479,In_261);
nor U2625 (N_2625,In_355,In_224);
and U2626 (N_2626,In_297,In_35);
or U2627 (N_2627,In_1395,In_691);
and U2628 (N_2628,In_741,In_1160);
nand U2629 (N_2629,In_566,In_907);
or U2630 (N_2630,In_721,In_415);
nor U2631 (N_2631,In_1162,In_1168);
or U2632 (N_2632,In_1326,In_1405);
nor U2633 (N_2633,In_1421,In_1068);
nor U2634 (N_2634,In_340,In_535);
or U2635 (N_2635,In_1223,In_100);
xor U2636 (N_2636,In_970,In_19);
nand U2637 (N_2637,In_619,In_999);
or U2638 (N_2638,In_786,In_937);
and U2639 (N_2639,In_74,In_315);
nand U2640 (N_2640,In_316,In_262);
nand U2641 (N_2641,In_1417,In_486);
nand U2642 (N_2642,In_1471,In_611);
nor U2643 (N_2643,In_1328,In_813);
nand U2644 (N_2644,In_1153,In_315);
and U2645 (N_2645,In_509,In_348);
nand U2646 (N_2646,In_654,In_328);
or U2647 (N_2647,In_546,In_793);
or U2648 (N_2648,In_1116,In_1375);
nor U2649 (N_2649,In_1196,In_438);
and U2650 (N_2650,In_960,In_860);
nand U2651 (N_2651,In_229,In_1289);
nand U2652 (N_2652,In_888,In_570);
nand U2653 (N_2653,In_1321,In_67);
nor U2654 (N_2654,In_123,In_546);
nand U2655 (N_2655,In_188,In_212);
or U2656 (N_2656,In_899,In_585);
and U2657 (N_2657,In_799,In_226);
nor U2658 (N_2658,In_801,In_961);
and U2659 (N_2659,In_446,In_884);
or U2660 (N_2660,In_1155,In_1005);
nand U2661 (N_2661,In_535,In_481);
nand U2662 (N_2662,In_304,In_747);
nor U2663 (N_2663,In_111,In_832);
nand U2664 (N_2664,In_513,In_272);
or U2665 (N_2665,In_943,In_659);
nor U2666 (N_2666,In_1103,In_1410);
and U2667 (N_2667,In_1425,In_131);
nand U2668 (N_2668,In_175,In_1489);
nor U2669 (N_2669,In_613,In_655);
and U2670 (N_2670,In_1190,In_351);
and U2671 (N_2671,In_289,In_970);
and U2672 (N_2672,In_1266,In_225);
nand U2673 (N_2673,In_984,In_360);
nand U2674 (N_2674,In_1023,In_379);
or U2675 (N_2675,In_507,In_317);
nand U2676 (N_2676,In_1454,In_982);
and U2677 (N_2677,In_471,In_1036);
nand U2678 (N_2678,In_630,In_549);
nand U2679 (N_2679,In_1018,In_808);
or U2680 (N_2680,In_643,In_7);
nand U2681 (N_2681,In_563,In_593);
nor U2682 (N_2682,In_850,In_1191);
or U2683 (N_2683,In_1254,In_218);
nor U2684 (N_2684,In_659,In_11);
nor U2685 (N_2685,In_479,In_714);
and U2686 (N_2686,In_1165,In_895);
or U2687 (N_2687,In_1102,In_412);
nand U2688 (N_2688,In_147,In_1081);
or U2689 (N_2689,In_40,In_1185);
nor U2690 (N_2690,In_631,In_8);
nor U2691 (N_2691,In_1493,In_585);
or U2692 (N_2692,In_792,In_110);
and U2693 (N_2693,In_520,In_1343);
nand U2694 (N_2694,In_810,In_723);
or U2695 (N_2695,In_218,In_1001);
nand U2696 (N_2696,In_162,In_1400);
or U2697 (N_2697,In_476,In_884);
or U2698 (N_2698,In_1132,In_1112);
and U2699 (N_2699,In_1043,In_158);
nand U2700 (N_2700,In_77,In_93);
nand U2701 (N_2701,In_378,In_1440);
nor U2702 (N_2702,In_331,In_305);
nand U2703 (N_2703,In_482,In_437);
nand U2704 (N_2704,In_94,In_175);
nand U2705 (N_2705,In_753,In_1273);
and U2706 (N_2706,In_1308,In_1483);
nor U2707 (N_2707,In_1335,In_22);
nor U2708 (N_2708,In_1056,In_1483);
or U2709 (N_2709,In_1287,In_507);
nor U2710 (N_2710,In_578,In_764);
and U2711 (N_2711,In_1281,In_493);
or U2712 (N_2712,In_1160,In_1017);
or U2713 (N_2713,In_1109,In_455);
nor U2714 (N_2714,In_406,In_1252);
and U2715 (N_2715,In_1273,In_1041);
nand U2716 (N_2716,In_165,In_1326);
nand U2717 (N_2717,In_246,In_895);
nand U2718 (N_2718,In_646,In_1041);
nor U2719 (N_2719,In_1091,In_535);
and U2720 (N_2720,In_146,In_1420);
nor U2721 (N_2721,In_27,In_458);
nor U2722 (N_2722,In_1194,In_548);
nand U2723 (N_2723,In_28,In_147);
and U2724 (N_2724,In_34,In_869);
and U2725 (N_2725,In_806,In_828);
nor U2726 (N_2726,In_816,In_12);
nand U2727 (N_2727,In_1319,In_1214);
or U2728 (N_2728,In_1327,In_648);
nor U2729 (N_2729,In_470,In_960);
or U2730 (N_2730,In_345,In_583);
or U2731 (N_2731,In_513,In_733);
or U2732 (N_2732,In_1045,In_1325);
nand U2733 (N_2733,In_413,In_836);
and U2734 (N_2734,In_856,In_242);
nand U2735 (N_2735,In_279,In_795);
or U2736 (N_2736,In_679,In_1358);
and U2737 (N_2737,In_407,In_857);
and U2738 (N_2738,In_731,In_1251);
and U2739 (N_2739,In_612,In_965);
and U2740 (N_2740,In_989,In_1113);
or U2741 (N_2741,In_762,In_1448);
or U2742 (N_2742,In_1238,In_437);
or U2743 (N_2743,In_235,In_137);
nand U2744 (N_2744,In_471,In_1198);
and U2745 (N_2745,In_1109,In_214);
and U2746 (N_2746,In_59,In_881);
nor U2747 (N_2747,In_273,In_300);
or U2748 (N_2748,In_1080,In_332);
and U2749 (N_2749,In_822,In_781);
nand U2750 (N_2750,In_242,In_738);
nand U2751 (N_2751,In_1232,In_192);
and U2752 (N_2752,In_696,In_1239);
nor U2753 (N_2753,In_813,In_778);
xor U2754 (N_2754,In_83,In_1013);
or U2755 (N_2755,In_1339,In_310);
nor U2756 (N_2756,In_1114,In_559);
or U2757 (N_2757,In_1327,In_1028);
xnor U2758 (N_2758,In_1065,In_1053);
nor U2759 (N_2759,In_640,In_188);
or U2760 (N_2760,In_161,In_1110);
and U2761 (N_2761,In_957,In_703);
nor U2762 (N_2762,In_994,In_712);
or U2763 (N_2763,In_1270,In_1497);
nand U2764 (N_2764,In_156,In_1197);
nor U2765 (N_2765,In_897,In_1494);
nand U2766 (N_2766,In_764,In_470);
nor U2767 (N_2767,In_669,In_925);
nand U2768 (N_2768,In_635,In_783);
nor U2769 (N_2769,In_408,In_935);
nor U2770 (N_2770,In_958,In_942);
nand U2771 (N_2771,In_162,In_486);
or U2772 (N_2772,In_182,In_55);
nor U2773 (N_2773,In_852,In_967);
nor U2774 (N_2774,In_250,In_1034);
nand U2775 (N_2775,In_1166,In_1389);
nand U2776 (N_2776,In_129,In_297);
and U2777 (N_2777,In_1025,In_786);
nor U2778 (N_2778,In_1071,In_1330);
or U2779 (N_2779,In_669,In_311);
nand U2780 (N_2780,In_241,In_428);
nand U2781 (N_2781,In_945,In_1457);
and U2782 (N_2782,In_396,In_645);
nand U2783 (N_2783,In_1099,In_880);
or U2784 (N_2784,In_234,In_31);
nor U2785 (N_2785,In_719,In_1186);
and U2786 (N_2786,In_984,In_773);
nand U2787 (N_2787,In_30,In_493);
and U2788 (N_2788,In_239,In_1021);
or U2789 (N_2789,In_268,In_961);
and U2790 (N_2790,In_623,In_474);
nand U2791 (N_2791,In_418,In_438);
and U2792 (N_2792,In_649,In_577);
nand U2793 (N_2793,In_568,In_348);
or U2794 (N_2794,In_962,In_893);
nor U2795 (N_2795,In_1156,In_690);
and U2796 (N_2796,In_21,In_738);
nand U2797 (N_2797,In_992,In_1272);
nor U2798 (N_2798,In_1167,In_676);
nor U2799 (N_2799,In_1064,In_449);
nor U2800 (N_2800,In_622,In_1115);
or U2801 (N_2801,In_1216,In_1295);
and U2802 (N_2802,In_1129,In_516);
and U2803 (N_2803,In_892,In_25);
nand U2804 (N_2804,In_379,In_1257);
nor U2805 (N_2805,In_211,In_1285);
nor U2806 (N_2806,In_1470,In_1054);
and U2807 (N_2807,In_416,In_1037);
and U2808 (N_2808,In_1448,In_518);
nor U2809 (N_2809,In_492,In_830);
or U2810 (N_2810,In_750,In_890);
or U2811 (N_2811,In_34,In_873);
nand U2812 (N_2812,In_1205,In_145);
nand U2813 (N_2813,In_1379,In_615);
and U2814 (N_2814,In_1198,In_317);
nand U2815 (N_2815,In_1011,In_381);
nor U2816 (N_2816,In_502,In_1289);
and U2817 (N_2817,In_241,In_72);
or U2818 (N_2818,In_387,In_1095);
and U2819 (N_2819,In_790,In_1031);
nor U2820 (N_2820,In_282,In_741);
and U2821 (N_2821,In_994,In_105);
or U2822 (N_2822,In_177,In_1347);
nor U2823 (N_2823,In_240,In_0);
nand U2824 (N_2824,In_256,In_72);
and U2825 (N_2825,In_338,In_1189);
nand U2826 (N_2826,In_612,In_729);
nand U2827 (N_2827,In_770,In_722);
nor U2828 (N_2828,In_803,In_80);
nor U2829 (N_2829,In_536,In_402);
or U2830 (N_2830,In_1377,In_1125);
and U2831 (N_2831,In_1347,In_594);
and U2832 (N_2832,In_225,In_1005);
and U2833 (N_2833,In_1147,In_225);
nand U2834 (N_2834,In_183,In_434);
nor U2835 (N_2835,In_662,In_693);
or U2836 (N_2836,In_37,In_1140);
or U2837 (N_2837,In_63,In_1275);
nor U2838 (N_2838,In_754,In_991);
and U2839 (N_2839,In_935,In_1334);
and U2840 (N_2840,In_502,In_1364);
xor U2841 (N_2841,In_528,In_679);
or U2842 (N_2842,In_740,In_937);
and U2843 (N_2843,In_1159,In_352);
xnor U2844 (N_2844,In_1414,In_464);
or U2845 (N_2845,In_116,In_1069);
nor U2846 (N_2846,In_336,In_381);
and U2847 (N_2847,In_1042,In_910);
and U2848 (N_2848,In_1459,In_578);
nor U2849 (N_2849,In_797,In_843);
and U2850 (N_2850,In_706,In_664);
and U2851 (N_2851,In_957,In_261);
nand U2852 (N_2852,In_1260,In_1019);
or U2853 (N_2853,In_273,In_384);
nor U2854 (N_2854,In_720,In_1041);
nand U2855 (N_2855,In_168,In_1450);
nand U2856 (N_2856,In_1403,In_648);
nand U2857 (N_2857,In_279,In_1352);
or U2858 (N_2858,In_1043,In_649);
nand U2859 (N_2859,In_95,In_845);
and U2860 (N_2860,In_603,In_564);
nor U2861 (N_2861,In_1464,In_355);
and U2862 (N_2862,In_1209,In_1176);
or U2863 (N_2863,In_514,In_906);
and U2864 (N_2864,In_9,In_1362);
and U2865 (N_2865,In_982,In_968);
or U2866 (N_2866,In_46,In_1374);
and U2867 (N_2867,In_1189,In_1001);
nand U2868 (N_2868,In_733,In_1121);
or U2869 (N_2869,In_689,In_652);
nand U2870 (N_2870,In_1234,In_673);
and U2871 (N_2871,In_769,In_1026);
and U2872 (N_2872,In_481,In_643);
or U2873 (N_2873,In_28,In_382);
nand U2874 (N_2874,In_138,In_357);
or U2875 (N_2875,In_669,In_327);
nand U2876 (N_2876,In_865,In_221);
and U2877 (N_2877,In_721,In_75);
nor U2878 (N_2878,In_1485,In_431);
nand U2879 (N_2879,In_579,In_1155);
or U2880 (N_2880,In_1497,In_168);
nor U2881 (N_2881,In_1033,In_341);
nor U2882 (N_2882,In_263,In_434);
nor U2883 (N_2883,In_362,In_991);
nand U2884 (N_2884,In_1494,In_905);
and U2885 (N_2885,In_192,In_87);
nand U2886 (N_2886,In_496,In_59);
and U2887 (N_2887,In_606,In_1197);
or U2888 (N_2888,In_1191,In_363);
xor U2889 (N_2889,In_799,In_306);
or U2890 (N_2890,In_381,In_387);
nand U2891 (N_2891,In_615,In_608);
nor U2892 (N_2892,In_1285,In_651);
nand U2893 (N_2893,In_1255,In_1201);
nor U2894 (N_2894,In_117,In_1409);
nor U2895 (N_2895,In_1136,In_1201);
or U2896 (N_2896,In_844,In_249);
and U2897 (N_2897,In_621,In_996);
nor U2898 (N_2898,In_1432,In_397);
nand U2899 (N_2899,In_32,In_518);
and U2900 (N_2900,In_37,In_417);
or U2901 (N_2901,In_732,In_1151);
nor U2902 (N_2902,In_76,In_443);
and U2903 (N_2903,In_318,In_1231);
and U2904 (N_2904,In_330,In_1052);
or U2905 (N_2905,In_603,In_534);
nand U2906 (N_2906,In_477,In_436);
and U2907 (N_2907,In_542,In_1274);
nor U2908 (N_2908,In_662,In_116);
nor U2909 (N_2909,In_1261,In_611);
nor U2910 (N_2910,In_605,In_1404);
nand U2911 (N_2911,In_1282,In_643);
nand U2912 (N_2912,In_821,In_764);
nor U2913 (N_2913,In_620,In_543);
nor U2914 (N_2914,In_962,In_1216);
and U2915 (N_2915,In_428,In_79);
nor U2916 (N_2916,In_106,In_1480);
nand U2917 (N_2917,In_1024,In_496);
nor U2918 (N_2918,In_1096,In_421);
and U2919 (N_2919,In_1152,In_1183);
nand U2920 (N_2920,In_843,In_502);
nand U2921 (N_2921,In_434,In_443);
nand U2922 (N_2922,In_64,In_296);
nand U2923 (N_2923,In_519,In_1347);
or U2924 (N_2924,In_519,In_540);
nand U2925 (N_2925,In_1167,In_1236);
nor U2926 (N_2926,In_1358,In_749);
nor U2927 (N_2927,In_719,In_1346);
and U2928 (N_2928,In_943,In_238);
nor U2929 (N_2929,In_469,In_441);
and U2930 (N_2930,In_262,In_795);
and U2931 (N_2931,In_1396,In_1109);
nand U2932 (N_2932,In_1161,In_243);
and U2933 (N_2933,In_1465,In_190);
nor U2934 (N_2934,In_695,In_1432);
nand U2935 (N_2935,In_496,In_220);
nor U2936 (N_2936,In_16,In_1427);
and U2937 (N_2937,In_1494,In_801);
or U2938 (N_2938,In_900,In_1289);
and U2939 (N_2939,In_667,In_1046);
and U2940 (N_2940,In_510,In_108);
or U2941 (N_2941,In_99,In_529);
and U2942 (N_2942,In_445,In_1115);
or U2943 (N_2943,In_446,In_930);
nand U2944 (N_2944,In_641,In_1127);
and U2945 (N_2945,In_728,In_192);
or U2946 (N_2946,In_375,In_838);
nor U2947 (N_2947,In_803,In_434);
and U2948 (N_2948,In_126,In_1077);
nor U2949 (N_2949,In_943,In_265);
and U2950 (N_2950,In_659,In_1447);
nor U2951 (N_2951,In_1140,In_569);
nand U2952 (N_2952,In_981,In_202);
nand U2953 (N_2953,In_1232,In_519);
xnor U2954 (N_2954,In_1498,In_167);
and U2955 (N_2955,In_129,In_1322);
xnor U2956 (N_2956,In_1252,In_1137);
nor U2957 (N_2957,In_534,In_677);
nand U2958 (N_2958,In_178,In_22);
nor U2959 (N_2959,In_13,In_540);
nor U2960 (N_2960,In_360,In_1119);
or U2961 (N_2961,In_803,In_358);
xnor U2962 (N_2962,In_1004,In_68);
and U2963 (N_2963,In_971,In_507);
nor U2964 (N_2964,In_46,In_728);
and U2965 (N_2965,In_1155,In_363);
or U2966 (N_2966,In_1010,In_609);
or U2967 (N_2967,In_435,In_1282);
xnor U2968 (N_2968,In_504,In_1228);
and U2969 (N_2969,In_1384,In_853);
nor U2970 (N_2970,In_4,In_888);
nand U2971 (N_2971,In_1368,In_1338);
nand U2972 (N_2972,In_330,In_1441);
and U2973 (N_2973,In_866,In_1139);
or U2974 (N_2974,In_1169,In_1012);
or U2975 (N_2975,In_998,In_94);
or U2976 (N_2976,In_633,In_419);
nand U2977 (N_2977,In_255,In_685);
nand U2978 (N_2978,In_346,In_987);
or U2979 (N_2979,In_1464,In_1407);
nand U2980 (N_2980,In_361,In_875);
and U2981 (N_2981,In_501,In_1455);
or U2982 (N_2982,In_1121,In_299);
nand U2983 (N_2983,In_1191,In_1464);
nand U2984 (N_2984,In_1425,In_952);
nand U2985 (N_2985,In_1394,In_458);
nor U2986 (N_2986,In_876,In_1214);
nor U2987 (N_2987,In_950,In_714);
nand U2988 (N_2988,In_94,In_1052);
nand U2989 (N_2989,In_1148,In_460);
or U2990 (N_2990,In_1147,In_1115);
nand U2991 (N_2991,In_1499,In_324);
and U2992 (N_2992,In_962,In_1284);
and U2993 (N_2993,In_58,In_255);
or U2994 (N_2994,In_242,In_498);
or U2995 (N_2995,In_383,In_819);
and U2996 (N_2996,In_598,In_723);
nor U2997 (N_2997,In_1393,In_1333);
nor U2998 (N_2998,In_1041,In_1246);
nand U2999 (N_2999,In_879,In_1176);
or U3000 (N_3000,In_1062,In_396);
xor U3001 (N_3001,In_576,In_1383);
or U3002 (N_3002,In_483,In_1209);
or U3003 (N_3003,In_1305,In_959);
nor U3004 (N_3004,In_12,In_1002);
nor U3005 (N_3005,In_229,In_1482);
nand U3006 (N_3006,In_443,In_234);
nor U3007 (N_3007,In_68,In_1472);
nand U3008 (N_3008,In_947,In_1184);
nor U3009 (N_3009,In_986,In_666);
nor U3010 (N_3010,In_179,In_864);
nand U3011 (N_3011,In_324,In_1384);
nand U3012 (N_3012,In_404,In_1054);
nor U3013 (N_3013,In_268,In_508);
nor U3014 (N_3014,In_1267,In_1172);
nand U3015 (N_3015,In_884,In_393);
nor U3016 (N_3016,In_59,In_715);
nand U3017 (N_3017,In_200,In_1446);
and U3018 (N_3018,In_952,In_960);
nor U3019 (N_3019,In_666,In_219);
nand U3020 (N_3020,In_286,In_352);
and U3021 (N_3021,In_1287,In_185);
and U3022 (N_3022,In_1256,In_1283);
and U3023 (N_3023,In_1448,In_570);
and U3024 (N_3024,In_764,In_1269);
nor U3025 (N_3025,In_704,In_834);
nand U3026 (N_3026,In_134,In_1175);
nand U3027 (N_3027,In_775,In_920);
nand U3028 (N_3028,In_884,In_930);
nor U3029 (N_3029,In_1323,In_722);
nand U3030 (N_3030,In_107,In_1348);
and U3031 (N_3031,In_49,In_814);
and U3032 (N_3032,In_818,In_1443);
or U3033 (N_3033,In_1148,In_759);
nor U3034 (N_3034,In_1260,In_1078);
or U3035 (N_3035,In_552,In_503);
or U3036 (N_3036,In_118,In_1443);
nor U3037 (N_3037,In_263,In_382);
xor U3038 (N_3038,In_1011,In_705);
and U3039 (N_3039,In_1036,In_406);
and U3040 (N_3040,In_251,In_661);
nand U3041 (N_3041,In_1250,In_1181);
nand U3042 (N_3042,In_819,In_347);
nor U3043 (N_3043,In_0,In_837);
nor U3044 (N_3044,In_541,In_1327);
or U3045 (N_3045,In_762,In_1499);
or U3046 (N_3046,In_1406,In_1157);
nand U3047 (N_3047,In_555,In_743);
or U3048 (N_3048,In_1412,In_872);
nor U3049 (N_3049,In_492,In_1082);
or U3050 (N_3050,In_1047,In_1422);
or U3051 (N_3051,In_630,In_500);
nor U3052 (N_3052,In_281,In_230);
nor U3053 (N_3053,In_294,In_630);
nor U3054 (N_3054,In_547,In_549);
and U3055 (N_3055,In_535,In_1458);
or U3056 (N_3056,In_482,In_1062);
or U3057 (N_3057,In_991,In_740);
nand U3058 (N_3058,In_1022,In_1291);
xor U3059 (N_3059,In_872,In_288);
nor U3060 (N_3060,In_403,In_500);
and U3061 (N_3061,In_942,In_1007);
and U3062 (N_3062,In_175,In_1013);
or U3063 (N_3063,In_998,In_296);
and U3064 (N_3064,In_956,In_1233);
nor U3065 (N_3065,In_1131,In_1022);
nor U3066 (N_3066,In_245,In_150);
nand U3067 (N_3067,In_1075,In_815);
nand U3068 (N_3068,In_241,In_1382);
nor U3069 (N_3069,In_942,In_594);
nand U3070 (N_3070,In_471,In_767);
and U3071 (N_3071,In_801,In_28);
nor U3072 (N_3072,In_1084,In_641);
and U3073 (N_3073,In_1489,In_1452);
and U3074 (N_3074,In_978,In_1260);
or U3075 (N_3075,In_669,In_973);
or U3076 (N_3076,In_282,In_1068);
and U3077 (N_3077,In_345,In_356);
or U3078 (N_3078,In_650,In_86);
nor U3079 (N_3079,In_791,In_57);
nor U3080 (N_3080,In_668,In_1034);
nand U3081 (N_3081,In_1337,In_1019);
or U3082 (N_3082,In_1106,In_1439);
xnor U3083 (N_3083,In_1498,In_1428);
nor U3084 (N_3084,In_752,In_578);
or U3085 (N_3085,In_240,In_787);
nor U3086 (N_3086,In_212,In_1029);
nand U3087 (N_3087,In_315,In_37);
and U3088 (N_3088,In_274,In_875);
or U3089 (N_3089,In_1206,In_882);
and U3090 (N_3090,In_1277,In_834);
and U3091 (N_3091,In_1450,In_445);
or U3092 (N_3092,In_962,In_101);
or U3093 (N_3093,In_168,In_1248);
nor U3094 (N_3094,In_960,In_754);
nor U3095 (N_3095,In_896,In_1368);
nand U3096 (N_3096,In_344,In_45);
and U3097 (N_3097,In_1460,In_884);
nor U3098 (N_3098,In_1329,In_1080);
nand U3099 (N_3099,In_1376,In_441);
and U3100 (N_3100,In_257,In_366);
nand U3101 (N_3101,In_1122,In_1137);
and U3102 (N_3102,In_14,In_105);
xnor U3103 (N_3103,In_382,In_283);
and U3104 (N_3104,In_407,In_10);
nand U3105 (N_3105,In_395,In_761);
nor U3106 (N_3106,In_1074,In_912);
nor U3107 (N_3107,In_1498,In_820);
nand U3108 (N_3108,In_606,In_1356);
nand U3109 (N_3109,In_1322,In_995);
and U3110 (N_3110,In_585,In_1314);
and U3111 (N_3111,In_1359,In_672);
nand U3112 (N_3112,In_1382,In_363);
nor U3113 (N_3113,In_417,In_1481);
or U3114 (N_3114,In_1424,In_930);
or U3115 (N_3115,In_158,In_615);
xnor U3116 (N_3116,In_928,In_645);
nand U3117 (N_3117,In_1466,In_1491);
or U3118 (N_3118,In_1424,In_1212);
and U3119 (N_3119,In_430,In_369);
or U3120 (N_3120,In_1409,In_517);
or U3121 (N_3121,In_345,In_485);
nor U3122 (N_3122,In_1493,In_130);
nand U3123 (N_3123,In_999,In_103);
nor U3124 (N_3124,In_332,In_991);
nor U3125 (N_3125,In_615,In_675);
nand U3126 (N_3126,In_557,In_16);
nand U3127 (N_3127,In_191,In_444);
nor U3128 (N_3128,In_533,In_692);
nand U3129 (N_3129,In_1103,In_705);
nor U3130 (N_3130,In_589,In_99);
nor U3131 (N_3131,In_942,In_530);
nand U3132 (N_3132,In_1057,In_1144);
or U3133 (N_3133,In_3,In_1309);
or U3134 (N_3134,In_911,In_435);
and U3135 (N_3135,In_616,In_120);
nand U3136 (N_3136,In_947,In_1159);
nand U3137 (N_3137,In_368,In_135);
nor U3138 (N_3138,In_606,In_1247);
xor U3139 (N_3139,In_922,In_609);
and U3140 (N_3140,In_507,In_1143);
and U3141 (N_3141,In_965,In_946);
nand U3142 (N_3142,In_891,In_636);
xnor U3143 (N_3143,In_372,In_3);
nand U3144 (N_3144,In_1147,In_930);
nor U3145 (N_3145,In_515,In_1269);
and U3146 (N_3146,In_306,In_692);
nor U3147 (N_3147,In_1215,In_385);
or U3148 (N_3148,In_1110,In_524);
nand U3149 (N_3149,In_890,In_731);
and U3150 (N_3150,In_1460,In_764);
nand U3151 (N_3151,In_535,In_5);
or U3152 (N_3152,In_142,In_461);
and U3153 (N_3153,In_1471,In_1181);
nor U3154 (N_3154,In_26,In_324);
and U3155 (N_3155,In_1332,In_350);
or U3156 (N_3156,In_1007,In_1148);
nand U3157 (N_3157,In_696,In_708);
nand U3158 (N_3158,In_137,In_1000);
and U3159 (N_3159,In_581,In_43);
and U3160 (N_3160,In_1033,In_1173);
and U3161 (N_3161,In_534,In_1352);
or U3162 (N_3162,In_1391,In_1302);
or U3163 (N_3163,In_299,In_1339);
or U3164 (N_3164,In_1225,In_1401);
or U3165 (N_3165,In_1293,In_754);
or U3166 (N_3166,In_81,In_867);
nand U3167 (N_3167,In_899,In_219);
or U3168 (N_3168,In_465,In_553);
and U3169 (N_3169,In_857,In_573);
nand U3170 (N_3170,In_633,In_530);
or U3171 (N_3171,In_1305,In_1307);
nor U3172 (N_3172,In_798,In_643);
nand U3173 (N_3173,In_1441,In_370);
or U3174 (N_3174,In_1485,In_540);
nor U3175 (N_3175,In_1047,In_83);
and U3176 (N_3176,In_809,In_511);
or U3177 (N_3177,In_1280,In_123);
or U3178 (N_3178,In_150,In_59);
nor U3179 (N_3179,In_195,In_836);
and U3180 (N_3180,In_766,In_573);
or U3181 (N_3181,In_1426,In_1139);
nor U3182 (N_3182,In_544,In_224);
nor U3183 (N_3183,In_541,In_990);
or U3184 (N_3184,In_1263,In_273);
nor U3185 (N_3185,In_801,In_914);
nor U3186 (N_3186,In_1177,In_582);
nand U3187 (N_3187,In_342,In_925);
or U3188 (N_3188,In_1284,In_1339);
nand U3189 (N_3189,In_643,In_1028);
nand U3190 (N_3190,In_1107,In_1421);
and U3191 (N_3191,In_1259,In_1096);
and U3192 (N_3192,In_844,In_423);
nand U3193 (N_3193,In_906,In_1096);
nor U3194 (N_3194,In_1475,In_1331);
or U3195 (N_3195,In_1326,In_517);
nor U3196 (N_3196,In_1189,In_109);
or U3197 (N_3197,In_1163,In_107);
and U3198 (N_3198,In_57,In_656);
nor U3199 (N_3199,In_56,In_397);
nor U3200 (N_3200,In_509,In_1417);
nor U3201 (N_3201,In_718,In_866);
or U3202 (N_3202,In_916,In_1370);
nand U3203 (N_3203,In_1363,In_1351);
or U3204 (N_3204,In_486,In_825);
nand U3205 (N_3205,In_290,In_1282);
or U3206 (N_3206,In_1104,In_1060);
xor U3207 (N_3207,In_310,In_217);
nor U3208 (N_3208,In_1179,In_795);
nand U3209 (N_3209,In_948,In_1083);
or U3210 (N_3210,In_169,In_530);
and U3211 (N_3211,In_401,In_1389);
and U3212 (N_3212,In_211,In_643);
nand U3213 (N_3213,In_178,In_1398);
or U3214 (N_3214,In_1229,In_158);
and U3215 (N_3215,In_782,In_1136);
and U3216 (N_3216,In_948,In_872);
nor U3217 (N_3217,In_703,In_568);
nand U3218 (N_3218,In_1443,In_1000);
xnor U3219 (N_3219,In_909,In_520);
nor U3220 (N_3220,In_675,In_340);
or U3221 (N_3221,In_1130,In_580);
and U3222 (N_3222,In_895,In_1360);
and U3223 (N_3223,In_128,In_1327);
and U3224 (N_3224,In_1217,In_75);
or U3225 (N_3225,In_800,In_1118);
nor U3226 (N_3226,In_105,In_580);
or U3227 (N_3227,In_1277,In_846);
or U3228 (N_3228,In_90,In_17);
or U3229 (N_3229,In_594,In_1222);
and U3230 (N_3230,In_1141,In_1489);
nand U3231 (N_3231,In_333,In_918);
and U3232 (N_3232,In_1325,In_576);
nor U3233 (N_3233,In_1440,In_1068);
nor U3234 (N_3234,In_848,In_606);
nand U3235 (N_3235,In_1266,In_628);
and U3236 (N_3236,In_473,In_894);
nor U3237 (N_3237,In_719,In_598);
or U3238 (N_3238,In_259,In_57);
and U3239 (N_3239,In_276,In_227);
nand U3240 (N_3240,In_1445,In_620);
nand U3241 (N_3241,In_84,In_62);
or U3242 (N_3242,In_551,In_1114);
nand U3243 (N_3243,In_1395,In_932);
and U3244 (N_3244,In_694,In_1078);
or U3245 (N_3245,In_1427,In_1091);
nor U3246 (N_3246,In_1432,In_363);
or U3247 (N_3247,In_650,In_208);
nor U3248 (N_3248,In_587,In_106);
and U3249 (N_3249,In_628,In_1208);
and U3250 (N_3250,In_1185,In_1440);
nor U3251 (N_3251,In_986,In_764);
and U3252 (N_3252,In_875,In_997);
or U3253 (N_3253,In_1327,In_142);
and U3254 (N_3254,In_1333,In_1077);
or U3255 (N_3255,In_1267,In_356);
nand U3256 (N_3256,In_343,In_516);
and U3257 (N_3257,In_843,In_1482);
or U3258 (N_3258,In_1041,In_1433);
nor U3259 (N_3259,In_1456,In_10);
or U3260 (N_3260,In_596,In_1047);
nor U3261 (N_3261,In_4,In_640);
nand U3262 (N_3262,In_1081,In_897);
nand U3263 (N_3263,In_406,In_1315);
nand U3264 (N_3264,In_1308,In_1297);
and U3265 (N_3265,In_1231,In_20);
nor U3266 (N_3266,In_215,In_1337);
or U3267 (N_3267,In_594,In_787);
nand U3268 (N_3268,In_750,In_737);
or U3269 (N_3269,In_1019,In_815);
nor U3270 (N_3270,In_271,In_330);
nor U3271 (N_3271,In_1265,In_1261);
nand U3272 (N_3272,In_1266,In_1323);
or U3273 (N_3273,In_662,In_1483);
or U3274 (N_3274,In_63,In_630);
and U3275 (N_3275,In_1135,In_1162);
or U3276 (N_3276,In_660,In_193);
and U3277 (N_3277,In_984,In_309);
nand U3278 (N_3278,In_485,In_1308);
nand U3279 (N_3279,In_1062,In_1261);
and U3280 (N_3280,In_1466,In_734);
nor U3281 (N_3281,In_608,In_939);
nor U3282 (N_3282,In_322,In_939);
and U3283 (N_3283,In_990,In_714);
or U3284 (N_3284,In_770,In_973);
or U3285 (N_3285,In_585,In_1077);
or U3286 (N_3286,In_1113,In_460);
or U3287 (N_3287,In_1132,In_863);
and U3288 (N_3288,In_1047,In_241);
nand U3289 (N_3289,In_1468,In_290);
nor U3290 (N_3290,In_280,In_83);
and U3291 (N_3291,In_782,In_1023);
and U3292 (N_3292,In_457,In_1284);
and U3293 (N_3293,In_1283,In_170);
nor U3294 (N_3294,In_575,In_254);
nand U3295 (N_3295,In_1083,In_909);
and U3296 (N_3296,In_1331,In_758);
or U3297 (N_3297,In_874,In_837);
and U3298 (N_3298,In_827,In_1268);
nor U3299 (N_3299,In_1052,In_56);
or U3300 (N_3300,In_1077,In_858);
nor U3301 (N_3301,In_1225,In_1257);
nand U3302 (N_3302,In_831,In_1495);
and U3303 (N_3303,In_736,In_702);
or U3304 (N_3304,In_761,In_460);
or U3305 (N_3305,In_1321,In_339);
nand U3306 (N_3306,In_1286,In_1178);
or U3307 (N_3307,In_785,In_738);
nand U3308 (N_3308,In_34,In_1110);
or U3309 (N_3309,In_610,In_587);
nor U3310 (N_3310,In_769,In_317);
nand U3311 (N_3311,In_1294,In_104);
nor U3312 (N_3312,In_582,In_797);
or U3313 (N_3313,In_1307,In_587);
nor U3314 (N_3314,In_519,In_851);
and U3315 (N_3315,In_1387,In_484);
or U3316 (N_3316,In_902,In_520);
and U3317 (N_3317,In_1454,In_597);
nand U3318 (N_3318,In_869,In_807);
xor U3319 (N_3319,In_373,In_1492);
nor U3320 (N_3320,In_1477,In_791);
and U3321 (N_3321,In_1240,In_149);
nor U3322 (N_3322,In_1013,In_392);
or U3323 (N_3323,In_714,In_1364);
and U3324 (N_3324,In_1184,In_1157);
and U3325 (N_3325,In_1366,In_1478);
and U3326 (N_3326,In_61,In_1215);
nor U3327 (N_3327,In_1429,In_1281);
xnor U3328 (N_3328,In_897,In_247);
nand U3329 (N_3329,In_1339,In_847);
nand U3330 (N_3330,In_759,In_1485);
nor U3331 (N_3331,In_1395,In_226);
nor U3332 (N_3332,In_951,In_1123);
or U3333 (N_3333,In_1496,In_924);
nand U3334 (N_3334,In_949,In_1444);
and U3335 (N_3335,In_1325,In_124);
and U3336 (N_3336,In_938,In_1201);
nor U3337 (N_3337,In_243,In_170);
or U3338 (N_3338,In_123,In_641);
or U3339 (N_3339,In_117,In_1316);
or U3340 (N_3340,In_1327,In_190);
nand U3341 (N_3341,In_118,In_647);
nor U3342 (N_3342,In_198,In_653);
or U3343 (N_3343,In_1392,In_513);
nand U3344 (N_3344,In_690,In_1247);
and U3345 (N_3345,In_549,In_23);
and U3346 (N_3346,In_573,In_1214);
nor U3347 (N_3347,In_519,In_948);
nor U3348 (N_3348,In_841,In_1069);
nand U3349 (N_3349,In_478,In_286);
and U3350 (N_3350,In_610,In_1269);
nand U3351 (N_3351,In_774,In_316);
and U3352 (N_3352,In_571,In_12);
nand U3353 (N_3353,In_1368,In_1054);
nand U3354 (N_3354,In_1477,In_1133);
nor U3355 (N_3355,In_1175,In_1027);
or U3356 (N_3356,In_872,In_1143);
nor U3357 (N_3357,In_535,In_949);
nor U3358 (N_3358,In_993,In_990);
nand U3359 (N_3359,In_772,In_1127);
nor U3360 (N_3360,In_1285,In_1097);
or U3361 (N_3361,In_1153,In_592);
and U3362 (N_3362,In_930,In_806);
or U3363 (N_3363,In_576,In_431);
nand U3364 (N_3364,In_1313,In_569);
nor U3365 (N_3365,In_647,In_666);
nor U3366 (N_3366,In_1421,In_1263);
nand U3367 (N_3367,In_421,In_700);
nor U3368 (N_3368,In_2,In_1420);
or U3369 (N_3369,In_631,In_1173);
nand U3370 (N_3370,In_1044,In_1090);
nand U3371 (N_3371,In_154,In_1359);
or U3372 (N_3372,In_1160,In_484);
and U3373 (N_3373,In_379,In_163);
nor U3374 (N_3374,In_57,In_1270);
and U3375 (N_3375,In_1029,In_780);
nor U3376 (N_3376,In_769,In_1471);
nand U3377 (N_3377,In_1147,In_1349);
or U3378 (N_3378,In_1480,In_999);
nand U3379 (N_3379,In_510,In_450);
nor U3380 (N_3380,In_1344,In_914);
or U3381 (N_3381,In_443,In_62);
nand U3382 (N_3382,In_1048,In_388);
and U3383 (N_3383,In_11,In_759);
nor U3384 (N_3384,In_651,In_696);
nand U3385 (N_3385,In_467,In_1312);
nor U3386 (N_3386,In_841,In_628);
and U3387 (N_3387,In_307,In_873);
nor U3388 (N_3388,In_299,In_1282);
and U3389 (N_3389,In_613,In_32);
nor U3390 (N_3390,In_494,In_221);
nand U3391 (N_3391,In_491,In_1063);
and U3392 (N_3392,In_1316,In_1188);
and U3393 (N_3393,In_566,In_1423);
nor U3394 (N_3394,In_1405,In_229);
nor U3395 (N_3395,In_319,In_339);
and U3396 (N_3396,In_948,In_138);
or U3397 (N_3397,In_680,In_621);
and U3398 (N_3398,In_1229,In_1185);
or U3399 (N_3399,In_1470,In_1319);
nand U3400 (N_3400,In_458,In_829);
nand U3401 (N_3401,In_625,In_366);
nand U3402 (N_3402,In_1491,In_808);
or U3403 (N_3403,In_1236,In_1324);
nor U3404 (N_3404,In_520,In_86);
or U3405 (N_3405,In_107,In_384);
and U3406 (N_3406,In_1467,In_312);
nand U3407 (N_3407,In_577,In_1179);
nor U3408 (N_3408,In_718,In_555);
nor U3409 (N_3409,In_470,In_418);
and U3410 (N_3410,In_965,In_980);
or U3411 (N_3411,In_414,In_379);
and U3412 (N_3412,In_449,In_116);
or U3413 (N_3413,In_222,In_540);
and U3414 (N_3414,In_596,In_1491);
xor U3415 (N_3415,In_176,In_275);
nor U3416 (N_3416,In_35,In_750);
nor U3417 (N_3417,In_54,In_35);
nand U3418 (N_3418,In_912,In_58);
nand U3419 (N_3419,In_672,In_548);
nor U3420 (N_3420,In_1337,In_1034);
and U3421 (N_3421,In_1050,In_340);
xnor U3422 (N_3422,In_1437,In_822);
or U3423 (N_3423,In_1006,In_738);
and U3424 (N_3424,In_796,In_845);
and U3425 (N_3425,In_51,In_426);
and U3426 (N_3426,In_523,In_1006);
nand U3427 (N_3427,In_866,In_1000);
and U3428 (N_3428,In_1220,In_182);
nor U3429 (N_3429,In_673,In_1173);
and U3430 (N_3430,In_1298,In_1410);
or U3431 (N_3431,In_1111,In_429);
or U3432 (N_3432,In_454,In_144);
and U3433 (N_3433,In_569,In_699);
nor U3434 (N_3434,In_1377,In_1241);
and U3435 (N_3435,In_1095,In_1275);
nand U3436 (N_3436,In_1105,In_1181);
and U3437 (N_3437,In_750,In_577);
and U3438 (N_3438,In_516,In_577);
nor U3439 (N_3439,In_441,In_537);
nand U3440 (N_3440,In_424,In_62);
nor U3441 (N_3441,In_472,In_33);
nor U3442 (N_3442,In_1483,In_991);
nor U3443 (N_3443,In_171,In_1101);
nor U3444 (N_3444,In_543,In_1051);
nor U3445 (N_3445,In_1246,In_572);
nor U3446 (N_3446,In_151,In_855);
or U3447 (N_3447,In_361,In_381);
and U3448 (N_3448,In_357,In_1055);
xnor U3449 (N_3449,In_1413,In_1458);
or U3450 (N_3450,In_529,In_489);
nor U3451 (N_3451,In_1435,In_21);
xnor U3452 (N_3452,In_785,In_98);
or U3453 (N_3453,In_354,In_446);
nand U3454 (N_3454,In_602,In_617);
nor U3455 (N_3455,In_671,In_1436);
nor U3456 (N_3456,In_289,In_907);
nor U3457 (N_3457,In_1201,In_1402);
and U3458 (N_3458,In_1320,In_977);
nor U3459 (N_3459,In_153,In_1397);
and U3460 (N_3460,In_1334,In_833);
nand U3461 (N_3461,In_645,In_1136);
nand U3462 (N_3462,In_70,In_852);
or U3463 (N_3463,In_1337,In_1302);
nand U3464 (N_3464,In_144,In_537);
nor U3465 (N_3465,In_1463,In_581);
and U3466 (N_3466,In_303,In_308);
and U3467 (N_3467,In_920,In_269);
nor U3468 (N_3468,In_264,In_961);
nor U3469 (N_3469,In_777,In_761);
or U3470 (N_3470,In_1471,In_689);
nand U3471 (N_3471,In_825,In_1219);
and U3472 (N_3472,In_739,In_550);
or U3473 (N_3473,In_142,In_1360);
nand U3474 (N_3474,In_698,In_551);
nand U3475 (N_3475,In_437,In_217);
nor U3476 (N_3476,In_436,In_487);
or U3477 (N_3477,In_286,In_1192);
nand U3478 (N_3478,In_861,In_1128);
or U3479 (N_3479,In_1401,In_726);
or U3480 (N_3480,In_669,In_170);
and U3481 (N_3481,In_1337,In_627);
and U3482 (N_3482,In_684,In_1174);
nor U3483 (N_3483,In_982,In_1081);
nand U3484 (N_3484,In_511,In_685);
nor U3485 (N_3485,In_22,In_338);
nor U3486 (N_3486,In_182,In_1197);
nand U3487 (N_3487,In_1463,In_1343);
or U3488 (N_3488,In_408,In_815);
nand U3489 (N_3489,In_910,In_94);
nand U3490 (N_3490,In_1302,In_1443);
nand U3491 (N_3491,In_1009,In_516);
nand U3492 (N_3492,In_1488,In_283);
and U3493 (N_3493,In_221,In_996);
or U3494 (N_3494,In_612,In_1363);
xnor U3495 (N_3495,In_254,In_633);
or U3496 (N_3496,In_476,In_743);
nand U3497 (N_3497,In_684,In_1204);
and U3498 (N_3498,In_1175,In_311);
and U3499 (N_3499,In_609,In_605);
or U3500 (N_3500,In_907,In_1251);
nor U3501 (N_3501,In_1290,In_759);
nand U3502 (N_3502,In_660,In_1245);
nand U3503 (N_3503,In_843,In_435);
and U3504 (N_3504,In_901,In_652);
nand U3505 (N_3505,In_20,In_420);
nor U3506 (N_3506,In_469,In_1483);
or U3507 (N_3507,In_101,In_955);
nor U3508 (N_3508,In_815,In_592);
nor U3509 (N_3509,In_1267,In_482);
or U3510 (N_3510,In_592,In_431);
and U3511 (N_3511,In_256,In_592);
and U3512 (N_3512,In_596,In_479);
xnor U3513 (N_3513,In_779,In_456);
and U3514 (N_3514,In_1129,In_184);
and U3515 (N_3515,In_416,In_178);
nor U3516 (N_3516,In_643,In_824);
nand U3517 (N_3517,In_989,In_116);
nand U3518 (N_3518,In_824,In_1062);
or U3519 (N_3519,In_203,In_891);
and U3520 (N_3520,In_1428,In_1252);
nand U3521 (N_3521,In_179,In_699);
or U3522 (N_3522,In_235,In_1188);
nand U3523 (N_3523,In_1226,In_1235);
and U3524 (N_3524,In_259,In_25);
and U3525 (N_3525,In_461,In_699);
nand U3526 (N_3526,In_971,In_1262);
nand U3527 (N_3527,In_443,In_608);
nor U3528 (N_3528,In_522,In_1194);
nor U3529 (N_3529,In_739,In_1178);
nand U3530 (N_3530,In_269,In_267);
nor U3531 (N_3531,In_1387,In_641);
nand U3532 (N_3532,In_675,In_700);
nand U3533 (N_3533,In_85,In_1377);
or U3534 (N_3534,In_55,In_562);
nor U3535 (N_3535,In_195,In_251);
and U3536 (N_3536,In_190,In_15);
nand U3537 (N_3537,In_917,In_1002);
nand U3538 (N_3538,In_680,In_990);
and U3539 (N_3539,In_1108,In_1493);
nand U3540 (N_3540,In_279,In_1262);
nor U3541 (N_3541,In_1350,In_1354);
nand U3542 (N_3542,In_1199,In_522);
nor U3543 (N_3543,In_672,In_179);
and U3544 (N_3544,In_321,In_334);
and U3545 (N_3545,In_856,In_954);
or U3546 (N_3546,In_466,In_284);
nand U3547 (N_3547,In_1409,In_168);
nor U3548 (N_3548,In_311,In_164);
or U3549 (N_3549,In_11,In_941);
nand U3550 (N_3550,In_421,In_90);
nand U3551 (N_3551,In_336,In_1036);
or U3552 (N_3552,In_1185,In_407);
nand U3553 (N_3553,In_1480,In_764);
nor U3554 (N_3554,In_950,In_627);
nand U3555 (N_3555,In_745,In_333);
and U3556 (N_3556,In_322,In_1454);
or U3557 (N_3557,In_1142,In_409);
nor U3558 (N_3558,In_1327,In_908);
and U3559 (N_3559,In_441,In_11);
nand U3560 (N_3560,In_343,In_156);
nand U3561 (N_3561,In_60,In_943);
and U3562 (N_3562,In_782,In_642);
nor U3563 (N_3563,In_754,In_1179);
nand U3564 (N_3564,In_47,In_1276);
and U3565 (N_3565,In_575,In_909);
and U3566 (N_3566,In_569,In_1445);
and U3567 (N_3567,In_917,In_1018);
or U3568 (N_3568,In_1207,In_997);
nor U3569 (N_3569,In_555,In_1097);
nor U3570 (N_3570,In_130,In_1257);
and U3571 (N_3571,In_549,In_622);
and U3572 (N_3572,In_520,In_1288);
nor U3573 (N_3573,In_116,In_781);
and U3574 (N_3574,In_303,In_462);
and U3575 (N_3575,In_773,In_1050);
nor U3576 (N_3576,In_1197,In_1064);
nand U3577 (N_3577,In_1250,In_828);
and U3578 (N_3578,In_760,In_146);
and U3579 (N_3579,In_738,In_651);
nand U3580 (N_3580,In_1086,In_1244);
nor U3581 (N_3581,In_1057,In_104);
nand U3582 (N_3582,In_31,In_491);
xnor U3583 (N_3583,In_197,In_191);
and U3584 (N_3584,In_1107,In_849);
nand U3585 (N_3585,In_271,In_528);
nand U3586 (N_3586,In_1193,In_1208);
nor U3587 (N_3587,In_875,In_888);
or U3588 (N_3588,In_1102,In_664);
nand U3589 (N_3589,In_949,In_1415);
and U3590 (N_3590,In_776,In_525);
or U3591 (N_3591,In_1459,In_845);
or U3592 (N_3592,In_1054,In_237);
nand U3593 (N_3593,In_1033,In_334);
and U3594 (N_3594,In_1443,In_183);
nor U3595 (N_3595,In_1342,In_745);
and U3596 (N_3596,In_1230,In_1235);
and U3597 (N_3597,In_815,In_1455);
and U3598 (N_3598,In_1217,In_681);
and U3599 (N_3599,In_867,In_1189);
nand U3600 (N_3600,In_26,In_173);
and U3601 (N_3601,In_750,In_235);
and U3602 (N_3602,In_1088,In_481);
and U3603 (N_3603,In_866,In_320);
xor U3604 (N_3604,In_1176,In_43);
nor U3605 (N_3605,In_743,In_970);
and U3606 (N_3606,In_265,In_498);
nor U3607 (N_3607,In_869,In_534);
and U3608 (N_3608,In_230,In_1341);
and U3609 (N_3609,In_587,In_328);
nor U3610 (N_3610,In_174,In_1340);
or U3611 (N_3611,In_991,In_602);
or U3612 (N_3612,In_1254,In_1330);
nor U3613 (N_3613,In_47,In_854);
or U3614 (N_3614,In_1142,In_1151);
nand U3615 (N_3615,In_634,In_1414);
or U3616 (N_3616,In_360,In_1226);
nand U3617 (N_3617,In_308,In_376);
or U3618 (N_3618,In_1461,In_223);
nor U3619 (N_3619,In_90,In_803);
nor U3620 (N_3620,In_556,In_792);
and U3621 (N_3621,In_14,In_388);
and U3622 (N_3622,In_325,In_371);
and U3623 (N_3623,In_1278,In_1219);
and U3624 (N_3624,In_1485,In_48);
or U3625 (N_3625,In_706,In_1353);
and U3626 (N_3626,In_625,In_681);
nand U3627 (N_3627,In_723,In_1399);
or U3628 (N_3628,In_1164,In_1020);
or U3629 (N_3629,In_824,In_622);
nand U3630 (N_3630,In_933,In_1318);
and U3631 (N_3631,In_1361,In_384);
and U3632 (N_3632,In_895,In_1051);
and U3633 (N_3633,In_522,In_281);
nand U3634 (N_3634,In_130,In_197);
or U3635 (N_3635,In_562,In_910);
or U3636 (N_3636,In_477,In_894);
or U3637 (N_3637,In_1261,In_1358);
or U3638 (N_3638,In_867,In_719);
nand U3639 (N_3639,In_399,In_1335);
or U3640 (N_3640,In_1293,In_145);
nor U3641 (N_3641,In_994,In_1058);
or U3642 (N_3642,In_1470,In_1038);
or U3643 (N_3643,In_1427,In_1435);
nand U3644 (N_3644,In_100,In_667);
nor U3645 (N_3645,In_537,In_109);
or U3646 (N_3646,In_665,In_1212);
nor U3647 (N_3647,In_416,In_620);
xor U3648 (N_3648,In_132,In_590);
and U3649 (N_3649,In_1044,In_1361);
nand U3650 (N_3650,In_94,In_521);
nor U3651 (N_3651,In_1389,In_13);
nor U3652 (N_3652,In_1393,In_1426);
nor U3653 (N_3653,In_172,In_182);
nor U3654 (N_3654,In_1204,In_1212);
nor U3655 (N_3655,In_930,In_1498);
nand U3656 (N_3656,In_483,In_827);
and U3657 (N_3657,In_1422,In_199);
and U3658 (N_3658,In_1312,In_1214);
nand U3659 (N_3659,In_480,In_94);
nand U3660 (N_3660,In_1264,In_909);
nor U3661 (N_3661,In_1191,In_1152);
and U3662 (N_3662,In_1076,In_35);
nand U3663 (N_3663,In_1126,In_1207);
nor U3664 (N_3664,In_1286,In_1468);
or U3665 (N_3665,In_1064,In_26);
nand U3666 (N_3666,In_1204,In_1081);
nand U3667 (N_3667,In_960,In_394);
or U3668 (N_3668,In_647,In_136);
nor U3669 (N_3669,In_1419,In_1443);
nor U3670 (N_3670,In_423,In_1158);
and U3671 (N_3671,In_1175,In_1396);
nand U3672 (N_3672,In_161,In_378);
and U3673 (N_3673,In_423,In_175);
and U3674 (N_3674,In_866,In_930);
nand U3675 (N_3675,In_1054,In_530);
and U3676 (N_3676,In_987,In_494);
nand U3677 (N_3677,In_3,In_93);
or U3678 (N_3678,In_432,In_59);
nor U3679 (N_3679,In_881,In_994);
or U3680 (N_3680,In_1400,In_452);
nor U3681 (N_3681,In_1418,In_1179);
or U3682 (N_3682,In_833,In_1267);
nor U3683 (N_3683,In_583,In_559);
and U3684 (N_3684,In_255,In_540);
and U3685 (N_3685,In_885,In_493);
or U3686 (N_3686,In_446,In_458);
nand U3687 (N_3687,In_1011,In_418);
and U3688 (N_3688,In_112,In_291);
or U3689 (N_3689,In_316,In_108);
nor U3690 (N_3690,In_725,In_87);
or U3691 (N_3691,In_72,In_188);
or U3692 (N_3692,In_642,In_18);
or U3693 (N_3693,In_838,In_1305);
or U3694 (N_3694,In_1302,In_1034);
nor U3695 (N_3695,In_572,In_126);
nor U3696 (N_3696,In_31,In_1412);
or U3697 (N_3697,In_948,In_1359);
or U3698 (N_3698,In_1216,In_504);
nand U3699 (N_3699,In_242,In_635);
xor U3700 (N_3700,In_1335,In_48);
and U3701 (N_3701,In_1478,In_539);
nand U3702 (N_3702,In_1441,In_892);
xor U3703 (N_3703,In_991,In_447);
and U3704 (N_3704,In_1065,In_1172);
and U3705 (N_3705,In_1213,In_365);
and U3706 (N_3706,In_36,In_1190);
and U3707 (N_3707,In_715,In_122);
nor U3708 (N_3708,In_169,In_590);
or U3709 (N_3709,In_673,In_454);
or U3710 (N_3710,In_654,In_598);
and U3711 (N_3711,In_831,In_475);
or U3712 (N_3712,In_1047,In_207);
nand U3713 (N_3713,In_1161,In_229);
or U3714 (N_3714,In_394,In_213);
or U3715 (N_3715,In_943,In_151);
nor U3716 (N_3716,In_859,In_146);
xnor U3717 (N_3717,In_744,In_634);
nand U3718 (N_3718,In_1194,In_62);
or U3719 (N_3719,In_1437,In_55);
or U3720 (N_3720,In_1006,In_86);
nor U3721 (N_3721,In_980,In_1046);
nand U3722 (N_3722,In_1071,In_231);
nor U3723 (N_3723,In_31,In_1224);
and U3724 (N_3724,In_868,In_850);
nor U3725 (N_3725,In_1102,In_1100);
nand U3726 (N_3726,In_763,In_643);
and U3727 (N_3727,In_39,In_919);
nand U3728 (N_3728,In_327,In_1492);
and U3729 (N_3729,In_1188,In_625);
and U3730 (N_3730,In_627,In_64);
and U3731 (N_3731,In_673,In_195);
nor U3732 (N_3732,In_1119,In_608);
and U3733 (N_3733,In_1060,In_800);
nor U3734 (N_3734,In_1441,In_1046);
and U3735 (N_3735,In_347,In_108);
nor U3736 (N_3736,In_681,In_1231);
nand U3737 (N_3737,In_535,In_1360);
nand U3738 (N_3738,In_1405,In_386);
and U3739 (N_3739,In_994,In_806);
nor U3740 (N_3740,In_1364,In_491);
and U3741 (N_3741,In_523,In_1031);
nand U3742 (N_3742,In_475,In_693);
nand U3743 (N_3743,In_99,In_1340);
nand U3744 (N_3744,In_315,In_648);
or U3745 (N_3745,In_766,In_724);
nor U3746 (N_3746,In_425,In_1346);
nor U3747 (N_3747,In_530,In_572);
nand U3748 (N_3748,In_96,In_1372);
and U3749 (N_3749,In_461,In_137);
nand U3750 (N_3750,In_563,In_1138);
nand U3751 (N_3751,In_1433,In_632);
and U3752 (N_3752,In_716,In_130);
and U3753 (N_3753,In_635,In_994);
or U3754 (N_3754,In_639,In_550);
and U3755 (N_3755,In_1119,In_1115);
nand U3756 (N_3756,In_1295,In_222);
nand U3757 (N_3757,In_1300,In_618);
nor U3758 (N_3758,In_850,In_1216);
or U3759 (N_3759,In_1321,In_1352);
and U3760 (N_3760,In_171,In_868);
and U3761 (N_3761,In_752,In_252);
nor U3762 (N_3762,In_583,In_1032);
or U3763 (N_3763,In_550,In_866);
nand U3764 (N_3764,In_1445,In_614);
nor U3765 (N_3765,In_816,In_220);
nor U3766 (N_3766,In_640,In_468);
or U3767 (N_3767,In_616,In_645);
nor U3768 (N_3768,In_213,In_41);
nand U3769 (N_3769,In_930,In_121);
or U3770 (N_3770,In_442,In_686);
and U3771 (N_3771,In_1123,In_601);
nor U3772 (N_3772,In_1032,In_1026);
or U3773 (N_3773,In_902,In_564);
and U3774 (N_3774,In_493,In_313);
nand U3775 (N_3775,In_690,In_319);
nand U3776 (N_3776,In_205,In_1189);
and U3777 (N_3777,In_510,In_1475);
nand U3778 (N_3778,In_1041,In_1044);
nand U3779 (N_3779,In_740,In_909);
nor U3780 (N_3780,In_193,In_1321);
and U3781 (N_3781,In_1126,In_157);
or U3782 (N_3782,In_446,In_1015);
or U3783 (N_3783,In_912,In_866);
nand U3784 (N_3784,In_1126,In_186);
and U3785 (N_3785,In_259,In_622);
nor U3786 (N_3786,In_893,In_981);
and U3787 (N_3787,In_908,In_1168);
or U3788 (N_3788,In_1395,In_339);
nand U3789 (N_3789,In_488,In_530);
xnor U3790 (N_3790,In_1368,In_1038);
and U3791 (N_3791,In_1446,In_331);
and U3792 (N_3792,In_1020,In_580);
nand U3793 (N_3793,In_1359,In_552);
nor U3794 (N_3794,In_98,In_1438);
nor U3795 (N_3795,In_266,In_1409);
or U3796 (N_3796,In_1447,In_958);
nand U3797 (N_3797,In_306,In_421);
nor U3798 (N_3798,In_1328,In_853);
nand U3799 (N_3799,In_521,In_926);
and U3800 (N_3800,In_53,In_421);
nor U3801 (N_3801,In_552,In_351);
nor U3802 (N_3802,In_567,In_394);
or U3803 (N_3803,In_307,In_1387);
and U3804 (N_3804,In_807,In_576);
nand U3805 (N_3805,In_78,In_55);
nor U3806 (N_3806,In_721,In_1432);
or U3807 (N_3807,In_892,In_849);
nor U3808 (N_3808,In_1396,In_1227);
nor U3809 (N_3809,In_1104,In_129);
nand U3810 (N_3810,In_872,In_1195);
or U3811 (N_3811,In_115,In_965);
or U3812 (N_3812,In_482,In_1134);
nand U3813 (N_3813,In_1284,In_337);
nand U3814 (N_3814,In_354,In_167);
or U3815 (N_3815,In_606,In_278);
and U3816 (N_3816,In_794,In_1420);
and U3817 (N_3817,In_406,In_706);
xnor U3818 (N_3818,In_287,In_1036);
and U3819 (N_3819,In_1287,In_640);
nor U3820 (N_3820,In_18,In_766);
and U3821 (N_3821,In_1407,In_716);
and U3822 (N_3822,In_38,In_46);
nand U3823 (N_3823,In_298,In_1132);
and U3824 (N_3824,In_1112,In_708);
and U3825 (N_3825,In_345,In_198);
or U3826 (N_3826,In_297,In_628);
nand U3827 (N_3827,In_987,In_487);
xnor U3828 (N_3828,In_697,In_815);
or U3829 (N_3829,In_1420,In_812);
nor U3830 (N_3830,In_1344,In_1450);
and U3831 (N_3831,In_187,In_1453);
nor U3832 (N_3832,In_104,In_1197);
nor U3833 (N_3833,In_733,In_491);
nand U3834 (N_3834,In_1415,In_728);
nor U3835 (N_3835,In_1318,In_1243);
and U3836 (N_3836,In_1323,In_1385);
nor U3837 (N_3837,In_1286,In_1066);
xnor U3838 (N_3838,In_1112,In_78);
nor U3839 (N_3839,In_566,In_605);
nand U3840 (N_3840,In_239,In_873);
and U3841 (N_3841,In_225,In_311);
or U3842 (N_3842,In_978,In_1019);
xnor U3843 (N_3843,In_528,In_977);
nor U3844 (N_3844,In_81,In_48);
nor U3845 (N_3845,In_1494,In_1217);
or U3846 (N_3846,In_412,In_728);
or U3847 (N_3847,In_1096,In_1413);
and U3848 (N_3848,In_1248,In_1233);
nand U3849 (N_3849,In_1477,In_153);
nand U3850 (N_3850,In_831,In_586);
and U3851 (N_3851,In_1318,In_1228);
nor U3852 (N_3852,In_1433,In_224);
nand U3853 (N_3853,In_584,In_423);
and U3854 (N_3854,In_1332,In_756);
nand U3855 (N_3855,In_432,In_1025);
or U3856 (N_3856,In_285,In_1112);
and U3857 (N_3857,In_494,In_794);
nor U3858 (N_3858,In_1392,In_312);
nand U3859 (N_3859,In_294,In_883);
nor U3860 (N_3860,In_1123,In_1015);
and U3861 (N_3861,In_1354,In_561);
nor U3862 (N_3862,In_176,In_198);
or U3863 (N_3863,In_1288,In_1301);
and U3864 (N_3864,In_1237,In_1272);
nor U3865 (N_3865,In_818,In_503);
and U3866 (N_3866,In_189,In_767);
nand U3867 (N_3867,In_595,In_704);
nor U3868 (N_3868,In_1255,In_1478);
or U3869 (N_3869,In_1334,In_1494);
and U3870 (N_3870,In_1293,In_447);
xor U3871 (N_3871,In_288,In_79);
and U3872 (N_3872,In_782,In_1245);
or U3873 (N_3873,In_1182,In_639);
or U3874 (N_3874,In_700,In_1484);
or U3875 (N_3875,In_746,In_765);
nand U3876 (N_3876,In_1261,In_1068);
or U3877 (N_3877,In_1494,In_750);
or U3878 (N_3878,In_506,In_1000);
or U3879 (N_3879,In_1482,In_920);
and U3880 (N_3880,In_1384,In_709);
or U3881 (N_3881,In_1489,In_47);
xnor U3882 (N_3882,In_1108,In_1012);
nand U3883 (N_3883,In_664,In_951);
or U3884 (N_3884,In_1402,In_1308);
and U3885 (N_3885,In_524,In_1305);
nor U3886 (N_3886,In_671,In_1239);
nand U3887 (N_3887,In_1431,In_1002);
nor U3888 (N_3888,In_469,In_971);
or U3889 (N_3889,In_176,In_966);
nand U3890 (N_3890,In_581,In_516);
or U3891 (N_3891,In_519,In_811);
and U3892 (N_3892,In_44,In_65);
and U3893 (N_3893,In_1448,In_1098);
nand U3894 (N_3894,In_367,In_818);
or U3895 (N_3895,In_990,In_1001);
nor U3896 (N_3896,In_1221,In_217);
and U3897 (N_3897,In_461,In_1182);
and U3898 (N_3898,In_419,In_1185);
and U3899 (N_3899,In_1226,In_357);
nor U3900 (N_3900,In_3,In_1050);
nand U3901 (N_3901,In_405,In_980);
and U3902 (N_3902,In_808,In_749);
nand U3903 (N_3903,In_753,In_112);
nand U3904 (N_3904,In_839,In_236);
or U3905 (N_3905,In_1210,In_179);
or U3906 (N_3906,In_1478,In_515);
and U3907 (N_3907,In_1061,In_696);
or U3908 (N_3908,In_786,In_455);
and U3909 (N_3909,In_144,In_704);
nand U3910 (N_3910,In_4,In_199);
nand U3911 (N_3911,In_726,In_44);
nand U3912 (N_3912,In_482,In_287);
and U3913 (N_3913,In_1255,In_447);
nand U3914 (N_3914,In_1268,In_1166);
nor U3915 (N_3915,In_722,In_37);
and U3916 (N_3916,In_1368,In_1328);
xor U3917 (N_3917,In_177,In_892);
nor U3918 (N_3918,In_1168,In_891);
nor U3919 (N_3919,In_344,In_728);
nand U3920 (N_3920,In_26,In_574);
or U3921 (N_3921,In_991,In_144);
and U3922 (N_3922,In_163,In_32);
nand U3923 (N_3923,In_327,In_896);
nor U3924 (N_3924,In_434,In_717);
nand U3925 (N_3925,In_675,In_1302);
or U3926 (N_3926,In_490,In_68);
nor U3927 (N_3927,In_498,In_340);
nor U3928 (N_3928,In_904,In_1385);
and U3929 (N_3929,In_257,In_86);
nand U3930 (N_3930,In_1161,In_561);
nand U3931 (N_3931,In_846,In_322);
and U3932 (N_3932,In_580,In_698);
nand U3933 (N_3933,In_1044,In_902);
and U3934 (N_3934,In_99,In_1191);
and U3935 (N_3935,In_1105,In_742);
nor U3936 (N_3936,In_564,In_757);
xnor U3937 (N_3937,In_116,In_233);
nor U3938 (N_3938,In_1297,In_851);
or U3939 (N_3939,In_1115,In_368);
xnor U3940 (N_3940,In_1358,In_171);
nor U3941 (N_3941,In_1368,In_1084);
nand U3942 (N_3942,In_757,In_1274);
nand U3943 (N_3943,In_1048,In_567);
nand U3944 (N_3944,In_200,In_548);
nor U3945 (N_3945,In_305,In_144);
nor U3946 (N_3946,In_975,In_1413);
nand U3947 (N_3947,In_1028,In_1030);
and U3948 (N_3948,In_1315,In_1458);
or U3949 (N_3949,In_97,In_10);
and U3950 (N_3950,In_912,In_1194);
and U3951 (N_3951,In_1102,In_848);
nor U3952 (N_3952,In_1396,In_678);
nand U3953 (N_3953,In_63,In_855);
nand U3954 (N_3954,In_807,In_887);
nor U3955 (N_3955,In_977,In_1418);
or U3956 (N_3956,In_803,In_867);
or U3957 (N_3957,In_951,In_808);
or U3958 (N_3958,In_947,In_392);
or U3959 (N_3959,In_817,In_1434);
and U3960 (N_3960,In_814,In_66);
and U3961 (N_3961,In_860,In_1448);
nand U3962 (N_3962,In_1132,In_733);
nand U3963 (N_3963,In_1092,In_1441);
or U3964 (N_3964,In_1208,In_730);
or U3965 (N_3965,In_356,In_347);
nor U3966 (N_3966,In_711,In_253);
nor U3967 (N_3967,In_1096,In_146);
nand U3968 (N_3968,In_854,In_1119);
and U3969 (N_3969,In_292,In_348);
nor U3970 (N_3970,In_602,In_871);
nand U3971 (N_3971,In_1320,In_1455);
or U3972 (N_3972,In_405,In_1108);
or U3973 (N_3973,In_1128,In_1001);
nor U3974 (N_3974,In_229,In_454);
nor U3975 (N_3975,In_480,In_366);
and U3976 (N_3976,In_183,In_1130);
and U3977 (N_3977,In_567,In_1262);
or U3978 (N_3978,In_944,In_1134);
and U3979 (N_3979,In_340,In_1067);
nand U3980 (N_3980,In_1147,In_1297);
nand U3981 (N_3981,In_1171,In_875);
and U3982 (N_3982,In_590,In_341);
nor U3983 (N_3983,In_1240,In_674);
or U3984 (N_3984,In_36,In_1433);
nand U3985 (N_3985,In_954,In_1434);
or U3986 (N_3986,In_741,In_325);
or U3987 (N_3987,In_1350,In_493);
or U3988 (N_3988,In_654,In_214);
nor U3989 (N_3989,In_299,In_926);
nand U3990 (N_3990,In_53,In_538);
and U3991 (N_3991,In_412,In_1352);
nand U3992 (N_3992,In_453,In_786);
nand U3993 (N_3993,In_816,In_43);
or U3994 (N_3994,In_1072,In_756);
nand U3995 (N_3995,In_641,In_1285);
or U3996 (N_3996,In_286,In_971);
and U3997 (N_3997,In_614,In_317);
xor U3998 (N_3998,In_1341,In_505);
and U3999 (N_3999,In_739,In_217);
or U4000 (N_4000,In_417,In_191);
nor U4001 (N_4001,In_205,In_40);
xnor U4002 (N_4002,In_193,In_644);
nand U4003 (N_4003,In_126,In_462);
and U4004 (N_4004,In_1048,In_871);
and U4005 (N_4005,In_379,In_48);
or U4006 (N_4006,In_1376,In_755);
or U4007 (N_4007,In_1407,In_222);
and U4008 (N_4008,In_769,In_922);
nor U4009 (N_4009,In_539,In_586);
nor U4010 (N_4010,In_319,In_705);
and U4011 (N_4011,In_928,In_112);
nand U4012 (N_4012,In_1124,In_1194);
or U4013 (N_4013,In_1410,In_129);
nand U4014 (N_4014,In_1393,In_1279);
xnor U4015 (N_4015,In_854,In_244);
nand U4016 (N_4016,In_931,In_28);
and U4017 (N_4017,In_1124,In_877);
nand U4018 (N_4018,In_106,In_1417);
xnor U4019 (N_4019,In_27,In_436);
nor U4020 (N_4020,In_1015,In_783);
or U4021 (N_4021,In_894,In_631);
and U4022 (N_4022,In_382,In_43);
nor U4023 (N_4023,In_184,In_987);
nor U4024 (N_4024,In_674,In_1239);
nor U4025 (N_4025,In_83,In_576);
and U4026 (N_4026,In_345,In_613);
and U4027 (N_4027,In_544,In_1102);
and U4028 (N_4028,In_241,In_198);
nand U4029 (N_4029,In_1460,In_1206);
or U4030 (N_4030,In_217,In_14);
or U4031 (N_4031,In_1060,In_336);
nand U4032 (N_4032,In_574,In_77);
or U4033 (N_4033,In_195,In_1402);
nand U4034 (N_4034,In_584,In_1463);
or U4035 (N_4035,In_970,In_1341);
xnor U4036 (N_4036,In_1096,In_564);
nor U4037 (N_4037,In_626,In_1203);
and U4038 (N_4038,In_620,In_8);
and U4039 (N_4039,In_614,In_506);
and U4040 (N_4040,In_1134,In_224);
or U4041 (N_4041,In_753,In_377);
nor U4042 (N_4042,In_759,In_168);
nor U4043 (N_4043,In_1051,In_632);
and U4044 (N_4044,In_1229,In_503);
nand U4045 (N_4045,In_1122,In_825);
nand U4046 (N_4046,In_397,In_1479);
nand U4047 (N_4047,In_309,In_780);
nor U4048 (N_4048,In_474,In_1478);
and U4049 (N_4049,In_406,In_536);
nor U4050 (N_4050,In_665,In_611);
and U4051 (N_4051,In_129,In_1421);
nor U4052 (N_4052,In_933,In_753);
or U4053 (N_4053,In_1496,In_382);
and U4054 (N_4054,In_413,In_365);
and U4055 (N_4055,In_560,In_761);
or U4056 (N_4056,In_441,In_507);
nor U4057 (N_4057,In_1446,In_172);
nand U4058 (N_4058,In_459,In_314);
nor U4059 (N_4059,In_1406,In_802);
nand U4060 (N_4060,In_173,In_406);
nor U4061 (N_4061,In_663,In_758);
xnor U4062 (N_4062,In_1054,In_1307);
nand U4063 (N_4063,In_200,In_1063);
nor U4064 (N_4064,In_506,In_865);
or U4065 (N_4065,In_1419,In_98);
or U4066 (N_4066,In_978,In_1007);
nor U4067 (N_4067,In_676,In_500);
or U4068 (N_4068,In_1100,In_225);
or U4069 (N_4069,In_1089,In_601);
xnor U4070 (N_4070,In_211,In_584);
nor U4071 (N_4071,In_1094,In_386);
and U4072 (N_4072,In_772,In_359);
or U4073 (N_4073,In_733,In_13);
nand U4074 (N_4074,In_1385,In_745);
and U4075 (N_4075,In_592,In_1126);
and U4076 (N_4076,In_1379,In_1460);
nand U4077 (N_4077,In_1199,In_1062);
nand U4078 (N_4078,In_991,In_235);
xnor U4079 (N_4079,In_156,In_678);
nor U4080 (N_4080,In_580,In_890);
and U4081 (N_4081,In_802,In_315);
nand U4082 (N_4082,In_17,In_1321);
nor U4083 (N_4083,In_636,In_375);
nor U4084 (N_4084,In_668,In_1116);
or U4085 (N_4085,In_269,In_519);
nand U4086 (N_4086,In_828,In_546);
or U4087 (N_4087,In_176,In_1325);
or U4088 (N_4088,In_451,In_1389);
and U4089 (N_4089,In_623,In_257);
nor U4090 (N_4090,In_1132,In_85);
nand U4091 (N_4091,In_1003,In_1105);
and U4092 (N_4092,In_1289,In_875);
or U4093 (N_4093,In_59,In_1057);
nor U4094 (N_4094,In_852,In_1277);
or U4095 (N_4095,In_767,In_673);
or U4096 (N_4096,In_1228,In_117);
nand U4097 (N_4097,In_867,In_338);
nor U4098 (N_4098,In_782,In_783);
nor U4099 (N_4099,In_1145,In_1420);
nor U4100 (N_4100,In_1061,In_613);
and U4101 (N_4101,In_125,In_104);
nand U4102 (N_4102,In_404,In_1319);
xor U4103 (N_4103,In_712,In_1017);
nor U4104 (N_4104,In_708,In_1408);
or U4105 (N_4105,In_291,In_623);
nand U4106 (N_4106,In_780,In_972);
nor U4107 (N_4107,In_1436,In_615);
or U4108 (N_4108,In_622,In_853);
xnor U4109 (N_4109,In_467,In_118);
and U4110 (N_4110,In_416,In_17);
xnor U4111 (N_4111,In_163,In_1493);
nand U4112 (N_4112,In_230,In_989);
and U4113 (N_4113,In_876,In_1187);
nor U4114 (N_4114,In_851,In_917);
nand U4115 (N_4115,In_414,In_139);
nor U4116 (N_4116,In_1360,In_1233);
or U4117 (N_4117,In_40,In_723);
or U4118 (N_4118,In_226,In_1425);
nor U4119 (N_4119,In_803,In_30);
and U4120 (N_4120,In_153,In_1470);
nor U4121 (N_4121,In_505,In_498);
nor U4122 (N_4122,In_1150,In_612);
nor U4123 (N_4123,In_1211,In_267);
or U4124 (N_4124,In_1294,In_650);
or U4125 (N_4125,In_1282,In_1461);
or U4126 (N_4126,In_1155,In_1353);
or U4127 (N_4127,In_1227,In_39);
nor U4128 (N_4128,In_161,In_255);
nor U4129 (N_4129,In_91,In_244);
and U4130 (N_4130,In_482,In_1459);
nand U4131 (N_4131,In_1346,In_664);
and U4132 (N_4132,In_1400,In_1110);
or U4133 (N_4133,In_693,In_1152);
or U4134 (N_4134,In_1383,In_453);
nor U4135 (N_4135,In_911,In_1451);
nand U4136 (N_4136,In_1350,In_663);
or U4137 (N_4137,In_563,In_1476);
or U4138 (N_4138,In_293,In_909);
nand U4139 (N_4139,In_1318,In_249);
and U4140 (N_4140,In_402,In_1231);
nor U4141 (N_4141,In_743,In_615);
and U4142 (N_4142,In_1235,In_465);
or U4143 (N_4143,In_1026,In_195);
and U4144 (N_4144,In_554,In_1115);
and U4145 (N_4145,In_389,In_200);
nor U4146 (N_4146,In_376,In_522);
nand U4147 (N_4147,In_7,In_1140);
and U4148 (N_4148,In_560,In_394);
or U4149 (N_4149,In_627,In_522);
nand U4150 (N_4150,In_959,In_1394);
or U4151 (N_4151,In_897,In_523);
or U4152 (N_4152,In_209,In_1006);
nand U4153 (N_4153,In_839,In_835);
and U4154 (N_4154,In_1276,In_108);
and U4155 (N_4155,In_391,In_390);
and U4156 (N_4156,In_775,In_159);
nand U4157 (N_4157,In_903,In_1497);
xnor U4158 (N_4158,In_329,In_1214);
nor U4159 (N_4159,In_1268,In_1246);
nor U4160 (N_4160,In_1245,In_510);
nor U4161 (N_4161,In_1093,In_1352);
nand U4162 (N_4162,In_1166,In_1237);
or U4163 (N_4163,In_193,In_1231);
nand U4164 (N_4164,In_1246,In_1385);
and U4165 (N_4165,In_30,In_830);
and U4166 (N_4166,In_876,In_834);
nand U4167 (N_4167,In_254,In_774);
or U4168 (N_4168,In_1453,In_64);
nor U4169 (N_4169,In_1131,In_1084);
nor U4170 (N_4170,In_1145,In_1104);
nor U4171 (N_4171,In_1281,In_619);
and U4172 (N_4172,In_295,In_1282);
nand U4173 (N_4173,In_68,In_521);
or U4174 (N_4174,In_749,In_1173);
and U4175 (N_4175,In_189,In_633);
or U4176 (N_4176,In_312,In_943);
nand U4177 (N_4177,In_215,In_433);
nor U4178 (N_4178,In_74,In_817);
or U4179 (N_4179,In_992,In_1072);
or U4180 (N_4180,In_228,In_64);
nor U4181 (N_4181,In_839,In_1150);
nand U4182 (N_4182,In_850,In_373);
nand U4183 (N_4183,In_1261,In_197);
nand U4184 (N_4184,In_1462,In_983);
or U4185 (N_4185,In_340,In_1168);
or U4186 (N_4186,In_1144,In_292);
and U4187 (N_4187,In_404,In_657);
or U4188 (N_4188,In_441,In_302);
nand U4189 (N_4189,In_1206,In_11);
nand U4190 (N_4190,In_503,In_1497);
nand U4191 (N_4191,In_213,In_654);
nor U4192 (N_4192,In_585,In_1162);
nor U4193 (N_4193,In_740,In_29);
and U4194 (N_4194,In_428,In_648);
or U4195 (N_4195,In_1123,In_447);
nand U4196 (N_4196,In_5,In_929);
or U4197 (N_4197,In_492,In_1038);
nand U4198 (N_4198,In_413,In_1096);
or U4199 (N_4199,In_1389,In_507);
nand U4200 (N_4200,In_302,In_696);
and U4201 (N_4201,In_42,In_1033);
or U4202 (N_4202,In_134,In_1162);
xor U4203 (N_4203,In_1185,In_925);
nand U4204 (N_4204,In_895,In_988);
nor U4205 (N_4205,In_1123,In_110);
and U4206 (N_4206,In_214,In_1391);
nor U4207 (N_4207,In_485,In_1352);
or U4208 (N_4208,In_534,In_1276);
and U4209 (N_4209,In_901,In_467);
and U4210 (N_4210,In_1121,In_1429);
nor U4211 (N_4211,In_674,In_1496);
nand U4212 (N_4212,In_545,In_446);
and U4213 (N_4213,In_52,In_633);
nand U4214 (N_4214,In_1024,In_43);
and U4215 (N_4215,In_1260,In_1426);
nor U4216 (N_4216,In_1334,In_987);
xor U4217 (N_4217,In_458,In_1470);
or U4218 (N_4218,In_462,In_646);
nor U4219 (N_4219,In_1339,In_872);
or U4220 (N_4220,In_502,In_1472);
nand U4221 (N_4221,In_997,In_1312);
or U4222 (N_4222,In_247,In_134);
nand U4223 (N_4223,In_767,In_690);
and U4224 (N_4224,In_1409,In_1416);
nor U4225 (N_4225,In_416,In_531);
and U4226 (N_4226,In_1402,In_184);
or U4227 (N_4227,In_616,In_870);
nand U4228 (N_4228,In_1316,In_1024);
nand U4229 (N_4229,In_861,In_1247);
nand U4230 (N_4230,In_184,In_1223);
or U4231 (N_4231,In_1200,In_469);
or U4232 (N_4232,In_803,In_1221);
nand U4233 (N_4233,In_510,In_1127);
nand U4234 (N_4234,In_1400,In_572);
and U4235 (N_4235,In_192,In_592);
or U4236 (N_4236,In_229,In_893);
or U4237 (N_4237,In_290,In_1425);
nor U4238 (N_4238,In_148,In_358);
and U4239 (N_4239,In_127,In_1295);
or U4240 (N_4240,In_1310,In_323);
nand U4241 (N_4241,In_1121,In_964);
nand U4242 (N_4242,In_255,In_705);
nand U4243 (N_4243,In_1188,In_1035);
and U4244 (N_4244,In_805,In_1060);
nand U4245 (N_4245,In_508,In_807);
xor U4246 (N_4246,In_1221,In_1019);
or U4247 (N_4247,In_1399,In_499);
or U4248 (N_4248,In_1371,In_582);
nand U4249 (N_4249,In_889,In_14);
and U4250 (N_4250,In_165,In_530);
or U4251 (N_4251,In_483,In_324);
or U4252 (N_4252,In_48,In_292);
nand U4253 (N_4253,In_1338,In_867);
and U4254 (N_4254,In_1092,In_82);
xnor U4255 (N_4255,In_1083,In_1374);
nand U4256 (N_4256,In_192,In_503);
and U4257 (N_4257,In_1034,In_390);
nand U4258 (N_4258,In_1057,In_300);
or U4259 (N_4259,In_170,In_924);
or U4260 (N_4260,In_449,In_468);
nor U4261 (N_4261,In_563,In_1360);
and U4262 (N_4262,In_1494,In_441);
xnor U4263 (N_4263,In_820,In_52);
and U4264 (N_4264,In_916,In_1186);
or U4265 (N_4265,In_938,In_930);
nand U4266 (N_4266,In_545,In_163);
or U4267 (N_4267,In_1136,In_739);
or U4268 (N_4268,In_1253,In_861);
or U4269 (N_4269,In_1472,In_299);
xor U4270 (N_4270,In_811,In_1032);
or U4271 (N_4271,In_350,In_566);
nand U4272 (N_4272,In_1424,In_1472);
nand U4273 (N_4273,In_261,In_19);
nor U4274 (N_4274,In_71,In_996);
nor U4275 (N_4275,In_1076,In_31);
xnor U4276 (N_4276,In_662,In_1156);
and U4277 (N_4277,In_12,In_1092);
and U4278 (N_4278,In_502,In_543);
nand U4279 (N_4279,In_1282,In_453);
and U4280 (N_4280,In_90,In_729);
or U4281 (N_4281,In_387,In_102);
nor U4282 (N_4282,In_1472,In_404);
or U4283 (N_4283,In_787,In_70);
nand U4284 (N_4284,In_224,In_1445);
or U4285 (N_4285,In_894,In_1276);
and U4286 (N_4286,In_838,In_722);
nand U4287 (N_4287,In_662,In_1278);
or U4288 (N_4288,In_532,In_798);
and U4289 (N_4289,In_836,In_854);
or U4290 (N_4290,In_105,In_1225);
nand U4291 (N_4291,In_172,In_1291);
and U4292 (N_4292,In_1285,In_1383);
nor U4293 (N_4293,In_1115,In_26);
and U4294 (N_4294,In_233,In_1176);
or U4295 (N_4295,In_310,In_689);
or U4296 (N_4296,In_1188,In_81);
or U4297 (N_4297,In_783,In_152);
nor U4298 (N_4298,In_747,In_663);
or U4299 (N_4299,In_147,In_857);
nor U4300 (N_4300,In_1462,In_592);
nor U4301 (N_4301,In_1250,In_459);
and U4302 (N_4302,In_1212,In_106);
nand U4303 (N_4303,In_51,In_1272);
nor U4304 (N_4304,In_697,In_130);
or U4305 (N_4305,In_774,In_1114);
and U4306 (N_4306,In_702,In_1322);
and U4307 (N_4307,In_849,In_744);
and U4308 (N_4308,In_841,In_880);
and U4309 (N_4309,In_666,In_1478);
nor U4310 (N_4310,In_1358,In_206);
and U4311 (N_4311,In_883,In_716);
or U4312 (N_4312,In_1303,In_1400);
nor U4313 (N_4313,In_286,In_1387);
nand U4314 (N_4314,In_549,In_388);
or U4315 (N_4315,In_404,In_241);
or U4316 (N_4316,In_208,In_1305);
or U4317 (N_4317,In_280,In_147);
and U4318 (N_4318,In_1226,In_1178);
or U4319 (N_4319,In_997,In_465);
nand U4320 (N_4320,In_416,In_75);
and U4321 (N_4321,In_1306,In_269);
nand U4322 (N_4322,In_301,In_77);
and U4323 (N_4323,In_953,In_1025);
nand U4324 (N_4324,In_529,In_445);
nor U4325 (N_4325,In_68,In_461);
xnor U4326 (N_4326,In_1363,In_1222);
nor U4327 (N_4327,In_60,In_1412);
and U4328 (N_4328,In_771,In_1431);
nand U4329 (N_4329,In_1403,In_165);
and U4330 (N_4330,In_537,In_178);
nor U4331 (N_4331,In_82,In_248);
and U4332 (N_4332,In_992,In_680);
nand U4333 (N_4333,In_1460,In_629);
nor U4334 (N_4334,In_1004,In_729);
nand U4335 (N_4335,In_1025,In_1188);
nor U4336 (N_4336,In_588,In_239);
nand U4337 (N_4337,In_62,In_520);
nor U4338 (N_4338,In_1453,In_850);
nor U4339 (N_4339,In_967,In_737);
or U4340 (N_4340,In_181,In_628);
nand U4341 (N_4341,In_150,In_872);
nand U4342 (N_4342,In_999,In_947);
nor U4343 (N_4343,In_405,In_219);
and U4344 (N_4344,In_571,In_542);
and U4345 (N_4345,In_23,In_537);
nor U4346 (N_4346,In_1058,In_1224);
nand U4347 (N_4347,In_162,In_336);
or U4348 (N_4348,In_1054,In_219);
xor U4349 (N_4349,In_179,In_623);
nor U4350 (N_4350,In_64,In_1178);
nand U4351 (N_4351,In_136,In_1311);
nor U4352 (N_4352,In_104,In_564);
nor U4353 (N_4353,In_1315,In_362);
and U4354 (N_4354,In_879,In_1414);
nor U4355 (N_4355,In_413,In_1180);
or U4356 (N_4356,In_818,In_179);
nand U4357 (N_4357,In_1331,In_708);
xor U4358 (N_4358,In_1345,In_1008);
nand U4359 (N_4359,In_875,In_1388);
or U4360 (N_4360,In_1101,In_151);
and U4361 (N_4361,In_1042,In_1219);
and U4362 (N_4362,In_562,In_617);
or U4363 (N_4363,In_354,In_162);
nor U4364 (N_4364,In_217,In_1206);
nand U4365 (N_4365,In_143,In_1196);
nand U4366 (N_4366,In_1353,In_1093);
or U4367 (N_4367,In_332,In_377);
nand U4368 (N_4368,In_795,In_415);
nor U4369 (N_4369,In_67,In_743);
or U4370 (N_4370,In_1126,In_59);
and U4371 (N_4371,In_872,In_1368);
xnor U4372 (N_4372,In_494,In_1089);
xnor U4373 (N_4373,In_479,In_77);
nor U4374 (N_4374,In_672,In_1209);
nand U4375 (N_4375,In_456,In_552);
nand U4376 (N_4376,In_238,In_880);
and U4377 (N_4377,In_440,In_569);
nor U4378 (N_4378,In_595,In_1437);
nor U4379 (N_4379,In_1154,In_359);
nand U4380 (N_4380,In_234,In_1022);
or U4381 (N_4381,In_5,In_1477);
nor U4382 (N_4382,In_586,In_762);
nor U4383 (N_4383,In_263,In_1180);
or U4384 (N_4384,In_1225,In_635);
or U4385 (N_4385,In_693,In_861);
or U4386 (N_4386,In_1176,In_983);
or U4387 (N_4387,In_934,In_102);
nor U4388 (N_4388,In_16,In_574);
nand U4389 (N_4389,In_341,In_560);
nor U4390 (N_4390,In_1302,In_1003);
or U4391 (N_4391,In_14,In_843);
and U4392 (N_4392,In_373,In_1365);
nand U4393 (N_4393,In_301,In_196);
or U4394 (N_4394,In_1492,In_1005);
nor U4395 (N_4395,In_1150,In_1190);
nand U4396 (N_4396,In_784,In_841);
and U4397 (N_4397,In_532,In_364);
and U4398 (N_4398,In_944,In_139);
nand U4399 (N_4399,In_758,In_417);
nor U4400 (N_4400,In_1008,In_953);
and U4401 (N_4401,In_1016,In_531);
or U4402 (N_4402,In_905,In_1129);
nor U4403 (N_4403,In_1394,In_361);
nand U4404 (N_4404,In_1028,In_106);
and U4405 (N_4405,In_864,In_466);
nor U4406 (N_4406,In_438,In_1395);
or U4407 (N_4407,In_1308,In_565);
nor U4408 (N_4408,In_488,In_570);
or U4409 (N_4409,In_842,In_1194);
and U4410 (N_4410,In_786,In_1438);
nand U4411 (N_4411,In_556,In_1217);
and U4412 (N_4412,In_1006,In_1391);
nand U4413 (N_4413,In_917,In_642);
nand U4414 (N_4414,In_125,In_1442);
nor U4415 (N_4415,In_1303,In_73);
nand U4416 (N_4416,In_1058,In_203);
nor U4417 (N_4417,In_1169,In_1220);
nand U4418 (N_4418,In_1435,In_654);
and U4419 (N_4419,In_1444,In_304);
nand U4420 (N_4420,In_1365,In_1406);
nand U4421 (N_4421,In_1499,In_77);
nor U4422 (N_4422,In_1164,In_1295);
nand U4423 (N_4423,In_1315,In_813);
nand U4424 (N_4424,In_703,In_865);
nand U4425 (N_4425,In_1381,In_6);
nor U4426 (N_4426,In_1179,In_1276);
and U4427 (N_4427,In_1131,In_1079);
nor U4428 (N_4428,In_187,In_1252);
nor U4429 (N_4429,In_708,In_1182);
nand U4430 (N_4430,In_150,In_491);
and U4431 (N_4431,In_570,In_529);
or U4432 (N_4432,In_673,In_1328);
nor U4433 (N_4433,In_291,In_77);
nor U4434 (N_4434,In_1,In_1314);
or U4435 (N_4435,In_1180,In_129);
and U4436 (N_4436,In_227,In_906);
and U4437 (N_4437,In_1325,In_1326);
nand U4438 (N_4438,In_117,In_1165);
and U4439 (N_4439,In_1471,In_1203);
nand U4440 (N_4440,In_320,In_1216);
nand U4441 (N_4441,In_903,In_1038);
and U4442 (N_4442,In_836,In_205);
nor U4443 (N_4443,In_168,In_880);
nand U4444 (N_4444,In_755,In_1193);
or U4445 (N_4445,In_240,In_530);
nand U4446 (N_4446,In_49,In_478);
nor U4447 (N_4447,In_1109,In_666);
nor U4448 (N_4448,In_363,In_419);
and U4449 (N_4449,In_44,In_14);
nand U4450 (N_4450,In_414,In_612);
and U4451 (N_4451,In_118,In_1283);
or U4452 (N_4452,In_201,In_732);
or U4453 (N_4453,In_1003,In_741);
and U4454 (N_4454,In_47,In_600);
and U4455 (N_4455,In_846,In_490);
nor U4456 (N_4456,In_125,In_751);
and U4457 (N_4457,In_666,In_91);
and U4458 (N_4458,In_243,In_1333);
or U4459 (N_4459,In_670,In_296);
nand U4460 (N_4460,In_417,In_1254);
nand U4461 (N_4461,In_1486,In_1273);
or U4462 (N_4462,In_198,In_139);
nand U4463 (N_4463,In_916,In_733);
and U4464 (N_4464,In_1110,In_357);
and U4465 (N_4465,In_331,In_481);
nand U4466 (N_4466,In_653,In_260);
nor U4467 (N_4467,In_969,In_1073);
or U4468 (N_4468,In_982,In_1371);
nand U4469 (N_4469,In_1325,In_1235);
nand U4470 (N_4470,In_269,In_218);
nor U4471 (N_4471,In_969,In_501);
or U4472 (N_4472,In_833,In_126);
and U4473 (N_4473,In_1022,In_461);
nand U4474 (N_4474,In_911,In_508);
nand U4475 (N_4475,In_1499,In_839);
nor U4476 (N_4476,In_1352,In_672);
and U4477 (N_4477,In_998,In_819);
nand U4478 (N_4478,In_1403,In_71);
xnor U4479 (N_4479,In_298,In_207);
and U4480 (N_4480,In_866,In_326);
and U4481 (N_4481,In_426,In_327);
nor U4482 (N_4482,In_644,In_1291);
nand U4483 (N_4483,In_970,In_536);
nor U4484 (N_4484,In_630,In_1393);
nor U4485 (N_4485,In_117,In_374);
and U4486 (N_4486,In_663,In_378);
or U4487 (N_4487,In_118,In_1451);
and U4488 (N_4488,In_1405,In_347);
nor U4489 (N_4489,In_1112,In_381);
nor U4490 (N_4490,In_1415,In_515);
and U4491 (N_4491,In_86,In_710);
and U4492 (N_4492,In_1250,In_216);
and U4493 (N_4493,In_619,In_447);
xnor U4494 (N_4494,In_132,In_410);
and U4495 (N_4495,In_1248,In_146);
or U4496 (N_4496,In_237,In_948);
nand U4497 (N_4497,In_1479,In_294);
nand U4498 (N_4498,In_73,In_1332);
nor U4499 (N_4499,In_725,In_699);
or U4500 (N_4500,In_308,In_623);
nand U4501 (N_4501,In_923,In_1437);
nor U4502 (N_4502,In_910,In_42);
and U4503 (N_4503,In_1243,In_1141);
or U4504 (N_4504,In_603,In_824);
or U4505 (N_4505,In_725,In_1344);
and U4506 (N_4506,In_1321,In_155);
or U4507 (N_4507,In_1306,In_414);
xnor U4508 (N_4508,In_1406,In_1130);
or U4509 (N_4509,In_125,In_1362);
or U4510 (N_4510,In_464,In_197);
nor U4511 (N_4511,In_933,In_284);
or U4512 (N_4512,In_1084,In_1193);
and U4513 (N_4513,In_1350,In_244);
or U4514 (N_4514,In_988,In_95);
and U4515 (N_4515,In_780,In_81);
and U4516 (N_4516,In_425,In_984);
nand U4517 (N_4517,In_763,In_1375);
nand U4518 (N_4518,In_615,In_1305);
or U4519 (N_4519,In_1092,In_23);
nand U4520 (N_4520,In_1493,In_1281);
or U4521 (N_4521,In_927,In_1216);
nand U4522 (N_4522,In_424,In_122);
xor U4523 (N_4523,In_443,In_304);
nand U4524 (N_4524,In_355,In_409);
nand U4525 (N_4525,In_524,In_644);
and U4526 (N_4526,In_499,In_837);
nor U4527 (N_4527,In_1387,In_138);
xor U4528 (N_4528,In_1319,In_565);
and U4529 (N_4529,In_963,In_220);
and U4530 (N_4530,In_455,In_1191);
and U4531 (N_4531,In_88,In_806);
and U4532 (N_4532,In_1367,In_22);
nor U4533 (N_4533,In_1247,In_694);
and U4534 (N_4534,In_946,In_150);
and U4535 (N_4535,In_968,In_624);
and U4536 (N_4536,In_1381,In_1284);
or U4537 (N_4537,In_1454,In_1375);
nand U4538 (N_4538,In_654,In_1018);
or U4539 (N_4539,In_719,In_618);
or U4540 (N_4540,In_454,In_239);
or U4541 (N_4541,In_960,In_250);
nor U4542 (N_4542,In_525,In_1333);
nand U4543 (N_4543,In_528,In_1405);
nand U4544 (N_4544,In_258,In_807);
nand U4545 (N_4545,In_868,In_690);
nor U4546 (N_4546,In_938,In_1230);
nor U4547 (N_4547,In_776,In_1093);
nor U4548 (N_4548,In_1309,In_1463);
and U4549 (N_4549,In_828,In_981);
nor U4550 (N_4550,In_234,In_985);
or U4551 (N_4551,In_454,In_1315);
xor U4552 (N_4552,In_1353,In_106);
nand U4553 (N_4553,In_678,In_997);
nor U4554 (N_4554,In_1424,In_1360);
nand U4555 (N_4555,In_622,In_95);
and U4556 (N_4556,In_1479,In_1064);
nor U4557 (N_4557,In_609,In_1296);
or U4558 (N_4558,In_1123,In_478);
or U4559 (N_4559,In_1145,In_909);
or U4560 (N_4560,In_932,In_426);
nand U4561 (N_4561,In_786,In_86);
nor U4562 (N_4562,In_1159,In_26);
nor U4563 (N_4563,In_215,In_117);
and U4564 (N_4564,In_1286,In_1360);
or U4565 (N_4565,In_62,In_493);
nor U4566 (N_4566,In_897,In_425);
nor U4567 (N_4567,In_1232,In_1135);
or U4568 (N_4568,In_63,In_945);
xor U4569 (N_4569,In_41,In_1);
and U4570 (N_4570,In_1360,In_359);
nand U4571 (N_4571,In_323,In_845);
or U4572 (N_4572,In_342,In_463);
nand U4573 (N_4573,In_237,In_271);
xnor U4574 (N_4574,In_286,In_779);
or U4575 (N_4575,In_500,In_63);
and U4576 (N_4576,In_160,In_1341);
or U4577 (N_4577,In_296,In_1210);
nor U4578 (N_4578,In_1285,In_755);
nor U4579 (N_4579,In_1427,In_22);
and U4580 (N_4580,In_1054,In_1262);
nand U4581 (N_4581,In_579,In_583);
and U4582 (N_4582,In_1014,In_1340);
nand U4583 (N_4583,In_1223,In_878);
or U4584 (N_4584,In_1194,In_1143);
or U4585 (N_4585,In_1127,In_1383);
nand U4586 (N_4586,In_289,In_823);
nor U4587 (N_4587,In_60,In_194);
or U4588 (N_4588,In_959,In_442);
xor U4589 (N_4589,In_865,In_426);
nand U4590 (N_4590,In_323,In_548);
nor U4591 (N_4591,In_511,In_626);
nor U4592 (N_4592,In_818,In_521);
nor U4593 (N_4593,In_963,In_455);
or U4594 (N_4594,In_146,In_913);
nand U4595 (N_4595,In_1316,In_298);
nor U4596 (N_4596,In_1362,In_1014);
nand U4597 (N_4597,In_1216,In_1143);
and U4598 (N_4598,In_1234,In_210);
nand U4599 (N_4599,In_1113,In_1362);
nor U4600 (N_4600,In_280,In_1217);
and U4601 (N_4601,In_776,In_211);
or U4602 (N_4602,In_566,In_439);
nand U4603 (N_4603,In_572,In_1294);
nor U4604 (N_4604,In_1357,In_796);
or U4605 (N_4605,In_50,In_624);
nand U4606 (N_4606,In_1040,In_307);
or U4607 (N_4607,In_992,In_957);
nand U4608 (N_4608,In_1018,In_55);
nand U4609 (N_4609,In_470,In_106);
nand U4610 (N_4610,In_834,In_1486);
or U4611 (N_4611,In_760,In_468);
and U4612 (N_4612,In_1140,In_161);
nor U4613 (N_4613,In_252,In_1472);
or U4614 (N_4614,In_1245,In_247);
nor U4615 (N_4615,In_1034,In_1224);
and U4616 (N_4616,In_1498,In_1038);
nand U4617 (N_4617,In_777,In_1361);
or U4618 (N_4618,In_1238,In_562);
and U4619 (N_4619,In_970,In_1440);
nor U4620 (N_4620,In_234,In_26);
nand U4621 (N_4621,In_119,In_78);
nor U4622 (N_4622,In_591,In_127);
or U4623 (N_4623,In_470,In_381);
or U4624 (N_4624,In_1170,In_1158);
nand U4625 (N_4625,In_1084,In_147);
nor U4626 (N_4626,In_647,In_409);
nor U4627 (N_4627,In_97,In_1085);
or U4628 (N_4628,In_1489,In_1202);
or U4629 (N_4629,In_1152,In_663);
or U4630 (N_4630,In_124,In_31);
nor U4631 (N_4631,In_30,In_807);
nand U4632 (N_4632,In_246,In_744);
nor U4633 (N_4633,In_1218,In_1258);
nand U4634 (N_4634,In_1265,In_1034);
and U4635 (N_4635,In_608,In_1100);
or U4636 (N_4636,In_320,In_451);
nor U4637 (N_4637,In_547,In_75);
and U4638 (N_4638,In_286,In_696);
nor U4639 (N_4639,In_970,In_885);
nand U4640 (N_4640,In_1463,In_716);
or U4641 (N_4641,In_29,In_846);
nor U4642 (N_4642,In_234,In_1453);
or U4643 (N_4643,In_74,In_204);
nor U4644 (N_4644,In_33,In_7);
nand U4645 (N_4645,In_778,In_523);
or U4646 (N_4646,In_623,In_1190);
or U4647 (N_4647,In_442,In_1196);
nor U4648 (N_4648,In_139,In_167);
nor U4649 (N_4649,In_1246,In_550);
nand U4650 (N_4650,In_351,In_353);
or U4651 (N_4651,In_278,In_520);
nor U4652 (N_4652,In_775,In_1152);
or U4653 (N_4653,In_535,In_1054);
or U4654 (N_4654,In_1040,In_756);
or U4655 (N_4655,In_422,In_1476);
nor U4656 (N_4656,In_104,In_594);
and U4657 (N_4657,In_1122,In_926);
or U4658 (N_4658,In_384,In_938);
and U4659 (N_4659,In_595,In_1178);
nand U4660 (N_4660,In_287,In_863);
nor U4661 (N_4661,In_1375,In_380);
nand U4662 (N_4662,In_1073,In_797);
nand U4663 (N_4663,In_58,In_1038);
or U4664 (N_4664,In_912,In_1256);
nand U4665 (N_4665,In_1420,In_883);
and U4666 (N_4666,In_742,In_73);
nand U4667 (N_4667,In_1365,In_1483);
and U4668 (N_4668,In_219,In_1211);
and U4669 (N_4669,In_545,In_733);
nand U4670 (N_4670,In_651,In_118);
or U4671 (N_4671,In_908,In_52);
and U4672 (N_4672,In_881,In_335);
nor U4673 (N_4673,In_1349,In_1008);
or U4674 (N_4674,In_668,In_187);
nand U4675 (N_4675,In_68,In_1224);
and U4676 (N_4676,In_1371,In_353);
or U4677 (N_4677,In_716,In_486);
xnor U4678 (N_4678,In_1170,In_137);
and U4679 (N_4679,In_658,In_659);
or U4680 (N_4680,In_324,In_552);
nor U4681 (N_4681,In_1352,In_239);
nor U4682 (N_4682,In_311,In_67);
or U4683 (N_4683,In_586,In_618);
or U4684 (N_4684,In_105,In_1445);
nand U4685 (N_4685,In_455,In_229);
nand U4686 (N_4686,In_1243,In_376);
nor U4687 (N_4687,In_931,In_466);
nor U4688 (N_4688,In_241,In_117);
nor U4689 (N_4689,In_1324,In_451);
or U4690 (N_4690,In_893,In_360);
xnor U4691 (N_4691,In_954,In_1311);
or U4692 (N_4692,In_1021,In_1192);
nand U4693 (N_4693,In_94,In_680);
nand U4694 (N_4694,In_269,In_941);
or U4695 (N_4695,In_952,In_1020);
and U4696 (N_4696,In_254,In_1096);
nor U4697 (N_4697,In_902,In_170);
nor U4698 (N_4698,In_758,In_724);
and U4699 (N_4699,In_1258,In_568);
nor U4700 (N_4700,In_308,In_450);
and U4701 (N_4701,In_1391,In_1078);
nor U4702 (N_4702,In_813,In_1423);
nand U4703 (N_4703,In_23,In_1207);
nand U4704 (N_4704,In_683,In_159);
and U4705 (N_4705,In_1483,In_48);
nand U4706 (N_4706,In_672,In_1471);
nand U4707 (N_4707,In_242,In_299);
or U4708 (N_4708,In_311,In_357);
nand U4709 (N_4709,In_595,In_502);
or U4710 (N_4710,In_556,In_292);
nand U4711 (N_4711,In_864,In_705);
or U4712 (N_4712,In_436,In_968);
nand U4713 (N_4713,In_270,In_431);
and U4714 (N_4714,In_1419,In_828);
nand U4715 (N_4715,In_448,In_1017);
and U4716 (N_4716,In_1048,In_1160);
or U4717 (N_4717,In_1330,In_170);
or U4718 (N_4718,In_1050,In_110);
nor U4719 (N_4719,In_1097,In_304);
nand U4720 (N_4720,In_711,In_933);
nand U4721 (N_4721,In_292,In_470);
and U4722 (N_4722,In_1416,In_785);
nor U4723 (N_4723,In_1178,In_744);
nand U4724 (N_4724,In_234,In_1222);
nor U4725 (N_4725,In_438,In_99);
nand U4726 (N_4726,In_71,In_894);
or U4727 (N_4727,In_1347,In_1371);
nand U4728 (N_4728,In_524,In_2);
and U4729 (N_4729,In_730,In_240);
nor U4730 (N_4730,In_1218,In_317);
and U4731 (N_4731,In_1171,In_474);
nand U4732 (N_4732,In_662,In_1358);
nand U4733 (N_4733,In_377,In_350);
nor U4734 (N_4734,In_27,In_1146);
and U4735 (N_4735,In_969,In_715);
and U4736 (N_4736,In_59,In_797);
and U4737 (N_4737,In_761,In_570);
and U4738 (N_4738,In_1233,In_450);
and U4739 (N_4739,In_1326,In_1151);
nand U4740 (N_4740,In_633,In_759);
and U4741 (N_4741,In_683,In_1052);
or U4742 (N_4742,In_503,In_975);
nand U4743 (N_4743,In_1042,In_1370);
xor U4744 (N_4744,In_1101,In_909);
nand U4745 (N_4745,In_463,In_1443);
nand U4746 (N_4746,In_1029,In_1388);
nor U4747 (N_4747,In_1094,In_247);
nor U4748 (N_4748,In_346,In_674);
and U4749 (N_4749,In_1416,In_877);
and U4750 (N_4750,In_1148,In_1313);
nor U4751 (N_4751,In_595,In_1007);
nor U4752 (N_4752,In_705,In_192);
nand U4753 (N_4753,In_367,In_1122);
or U4754 (N_4754,In_1286,In_1405);
nand U4755 (N_4755,In_603,In_252);
nor U4756 (N_4756,In_922,In_703);
nor U4757 (N_4757,In_32,In_413);
nor U4758 (N_4758,In_1064,In_835);
nor U4759 (N_4759,In_532,In_1450);
and U4760 (N_4760,In_1172,In_440);
or U4761 (N_4761,In_1477,In_880);
or U4762 (N_4762,In_389,In_1440);
nand U4763 (N_4763,In_48,In_457);
nand U4764 (N_4764,In_354,In_787);
nand U4765 (N_4765,In_713,In_778);
nand U4766 (N_4766,In_560,In_37);
nor U4767 (N_4767,In_125,In_1260);
nor U4768 (N_4768,In_410,In_1177);
nor U4769 (N_4769,In_1208,In_457);
nor U4770 (N_4770,In_1099,In_1431);
and U4771 (N_4771,In_794,In_597);
or U4772 (N_4772,In_869,In_91);
nand U4773 (N_4773,In_71,In_188);
nor U4774 (N_4774,In_1374,In_650);
nand U4775 (N_4775,In_863,In_761);
or U4776 (N_4776,In_354,In_733);
or U4777 (N_4777,In_890,In_1187);
nor U4778 (N_4778,In_1251,In_389);
and U4779 (N_4779,In_124,In_831);
nor U4780 (N_4780,In_1141,In_533);
and U4781 (N_4781,In_365,In_1030);
and U4782 (N_4782,In_478,In_725);
nor U4783 (N_4783,In_867,In_945);
nand U4784 (N_4784,In_1340,In_1364);
or U4785 (N_4785,In_1046,In_624);
nand U4786 (N_4786,In_287,In_113);
nor U4787 (N_4787,In_568,In_6);
nor U4788 (N_4788,In_740,In_804);
or U4789 (N_4789,In_217,In_297);
or U4790 (N_4790,In_303,In_141);
nand U4791 (N_4791,In_1107,In_741);
and U4792 (N_4792,In_1384,In_357);
or U4793 (N_4793,In_1092,In_674);
xor U4794 (N_4794,In_497,In_1276);
nor U4795 (N_4795,In_296,In_1476);
or U4796 (N_4796,In_19,In_1171);
or U4797 (N_4797,In_308,In_236);
or U4798 (N_4798,In_774,In_556);
nand U4799 (N_4799,In_1400,In_672);
nor U4800 (N_4800,In_761,In_263);
nor U4801 (N_4801,In_630,In_700);
nor U4802 (N_4802,In_663,In_673);
nor U4803 (N_4803,In_1404,In_1052);
nand U4804 (N_4804,In_709,In_212);
nand U4805 (N_4805,In_1342,In_446);
or U4806 (N_4806,In_769,In_458);
or U4807 (N_4807,In_56,In_856);
and U4808 (N_4808,In_993,In_179);
nand U4809 (N_4809,In_549,In_410);
and U4810 (N_4810,In_722,In_409);
xor U4811 (N_4811,In_1039,In_1094);
nor U4812 (N_4812,In_955,In_535);
nor U4813 (N_4813,In_441,In_1356);
nor U4814 (N_4814,In_232,In_639);
nand U4815 (N_4815,In_178,In_922);
or U4816 (N_4816,In_1226,In_1498);
nor U4817 (N_4817,In_1065,In_1277);
and U4818 (N_4818,In_1379,In_89);
xnor U4819 (N_4819,In_605,In_542);
nor U4820 (N_4820,In_1466,In_251);
nor U4821 (N_4821,In_257,In_1152);
nand U4822 (N_4822,In_1467,In_181);
nand U4823 (N_4823,In_695,In_1257);
or U4824 (N_4824,In_1438,In_112);
nand U4825 (N_4825,In_451,In_1091);
nand U4826 (N_4826,In_630,In_124);
or U4827 (N_4827,In_1057,In_1014);
and U4828 (N_4828,In_335,In_627);
nand U4829 (N_4829,In_361,In_1389);
and U4830 (N_4830,In_852,In_345);
or U4831 (N_4831,In_26,In_240);
nor U4832 (N_4832,In_700,In_46);
nand U4833 (N_4833,In_912,In_341);
and U4834 (N_4834,In_1361,In_606);
or U4835 (N_4835,In_243,In_1246);
or U4836 (N_4836,In_790,In_43);
nor U4837 (N_4837,In_516,In_965);
or U4838 (N_4838,In_258,In_507);
nand U4839 (N_4839,In_970,In_760);
and U4840 (N_4840,In_1373,In_959);
nand U4841 (N_4841,In_405,In_160);
or U4842 (N_4842,In_457,In_533);
or U4843 (N_4843,In_656,In_621);
nand U4844 (N_4844,In_290,In_837);
nor U4845 (N_4845,In_803,In_370);
nand U4846 (N_4846,In_902,In_679);
or U4847 (N_4847,In_1094,In_1248);
and U4848 (N_4848,In_812,In_602);
or U4849 (N_4849,In_1432,In_1142);
nor U4850 (N_4850,In_40,In_483);
nand U4851 (N_4851,In_551,In_1029);
and U4852 (N_4852,In_554,In_668);
and U4853 (N_4853,In_1200,In_558);
nor U4854 (N_4854,In_1461,In_1371);
or U4855 (N_4855,In_125,In_990);
or U4856 (N_4856,In_1373,In_1210);
nand U4857 (N_4857,In_521,In_1246);
nand U4858 (N_4858,In_988,In_934);
nor U4859 (N_4859,In_982,In_696);
or U4860 (N_4860,In_1421,In_777);
or U4861 (N_4861,In_58,In_500);
nand U4862 (N_4862,In_1369,In_1350);
or U4863 (N_4863,In_1314,In_563);
and U4864 (N_4864,In_1388,In_512);
nor U4865 (N_4865,In_1414,In_1427);
and U4866 (N_4866,In_663,In_1067);
or U4867 (N_4867,In_941,In_536);
and U4868 (N_4868,In_205,In_416);
or U4869 (N_4869,In_715,In_1157);
nor U4870 (N_4870,In_694,In_954);
or U4871 (N_4871,In_1060,In_549);
nand U4872 (N_4872,In_1006,In_968);
and U4873 (N_4873,In_1138,In_1296);
nor U4874 (N_4874,In_160,In_979);
or U4875 (N_4875,In_348,In_1337);
and U4876 (N_4876,In_305,In_1314);
nand U4877 (N_4877,In_1139,In_818);
or U4878 (N_4878,In_1011,In_224);
nand U4879 (N_4879,In_761,In_1115);
or U4880 (N_4880,In_34,In_234);
or U4881 (N_4881,In_808,In_1467);
and U4882 (N_4882,In_609,In_615);
nor U4883 (N_4883,In_245,In_868);
nor U4884 (N_4884,In_345,In_1343);
xnor U4885 (N_4885,In_957,In_519);
nand U4886 (N_4886,In_1164,In_17);
nor U4887 (N_4887,In_1497,In_1241);
and U4888 (N_4888,In_1239,In_1223);
or U4889 (N_4889,In_258,In_1020);
nand U4890 (N_4890,In_1172,In_1378);
nand U4891 (N_4891,In_1056,In_497);
and U4892 (N_4892,In_711,In_1380);
or U4893 (N_4893,In_1431,In_382);
nand U4894 (N_4894,In_56,In_204);
nand U4895 (N_4895,In_889,In_264);
or U4896 (N_4896,In_1385,In_35);
and U4897 (N_4897,In_787,In_1344);
nand U4898 (N_4898,In_1498,In_793);
nand U4899 (N_4899,In_228,In_655);
xnor U4900 (N_4900,In_134,In_1258);
nor U4901 (N_4901,In_957,In_720);
or U4902 (N_4902,In_23,In_897);
nand U4903 (N_4903,In_827,In_1401);
or U4904 (N_4904,In_646,In_402);
nor U4905 (N_4905,In_688,In_692);
and U4906 (N_4906,In_812,In_1430);
nand U4907 (N_4907,In_49,In_364);
nand U4908 (N_4908,In_814,In_47);
or U4909 (N_4909,In_531,In_701);
or U4910 (N_4910,In_1306,In_834);
or U4911 (N_4911,In_456,In_296);
and U4912 (N_4912,In_828,In_1466);
nor U4913 (N_4913,In_1281,In_973);
and U4914 (N_4914,In_602,In_1284);
nand U4915 (N_4915,In_1297,In_422);
or U4916 (N_4916,In_678,In_1154);
nand U4917 (N_4917,In_1337,In_58);
or U4918 (N_4918,In_1129,In_1057);
nand U4919 (N_4919,In_763,In_938);
nand U4920 (N_4920,In_1061,In_906);
nand U4921 (N_4921,In_810,In_353);
and U4922 (N_4922,In_845,In_692);
nor U4923 (N_4923,In_1205,In_584);
nand U4924 (N_4924,In_919,In_1308);
and U4925 (N_4925,In_357,In_278);
nand U4926 (N_4926,In_531,In_663);
or U4927 (N_4927,In_42,In_1008);
and U4928 (N_4928,In_1195,In_57);
nor U4929 (N_4929,In_279,In_46);
and U4930 (N_4930,In_539,In_288);
nand U4931 (N_4931,In_1069,In_158);
nand U4932 (N_4932,In_1079,In_614);
and U4933 (N_4933,In_664,In_1410);
nand U4934 (N_4934,In_281,In_81);
or U4935 (N_4935,In_1273,In_389);
and U4936 (N_4936,In_517,In_274);
or U4937 (N_4937,In_1364,In_93);
nor U4938 (N_4938,In_358,In_245);
nand U4939 (N_4939,In_1348,In_1273);
nand U4940 (N_4940,In_445,In_1219);
or U4941 (N_4941,In_1486,In_1233);
nor U4942 (N_4942,In_208,In_726);
or U4943 (N_4943,In_691,In_1118);
and U4944 (N_4944,In_813,In_327);
and U4945 (N_4945,In_873,In_900);
and U4946 (N_4946,In_262,In_457);
and U4947 (N_4947,In_1186,In_400);
and U4948 (N_4948,In_724,In_219);
or U4949 (N_4949,In_370,In_638);
nand U4950 (N_4950,In_28,In_612);
nor U4951 (N_4951,In_293,In_1442);
and U4952 (N_4952,In_125,In_979);
or U4953 (N_4953,In_414,In_846);
or U4954 (N_4954,In_123,In_740);
nand U4955 (N_4955,In_471,In_1338);
nand U4956 (N_4956,In_33,In_679);
and U4957 (N_4957,In_362,In_486);
nor U4958 (N_4958,In_756,In_173);
nand U4959 (N_4959,In_442,In_608);
nor U4960 (N_4960,In_1047,In_594);
nand U4961 (N_4961,In_546,In_374);
nand U4962 (N_4962,In_405,In_222);
or U4963 (N_4963,In_683,In_626);
nand U4964 (N_4964,In_136,In_139);
nor U4965 (N_4965,In_1169,In_238);
nor U4966 (N_4966,In_303,In_194);
nor U4967 (N_4967,In_1369,In_252);
nand U4968 (N_4968,In_47,In_183);
nor U4969 (N_4969,In_1240,In_1231);
nand U4970 (N_4970,In_551,In_666);
nand U4971 (N_4971,In_657,In_1192);
and U4972 (N_4972,In_972,In_140);
nand U4973 (N_4973,In_1067,In_1213);
or U4974 (N_4974,In_156,In_1138);
nor U4975 (N_4975,In_767,In_924);
xnor U4976 (N_4976,In_215,In_1204);
nor U4977 (N_4977,In_1289,In_587);
nor U4978 (N_4978,In_277,In_459);
nor U4979 (N_4979,In_634,In_0);
or U4980 (N_4980,In_608,In_500);
nand U4981 (N_4981,In_904,In_7);
and U4982 (N_4982,In_1052,In_201);
nor U4983 (N_4983,In_312,In_747);
nand U4984 (N_4984,In_779,In_1109);
and U4985 (N_4985,In_233,In_910);
or U4986 (N_4986,In_1125,In_841);
nor U4987 (N_4987,In_1432,In_1093);
nand U4988 (N_4988,In_189,In_1347);
nand U4989 (N_4989,In_1474,In_868);
or U4990 (N_4990,In_1096,In_1002);
nand U4991 (N_4991,In_1330,In_941);
xnor U4992 (N_4992,In_1120,In_1498);
and U4993 (N_4993,In_1303,In_1101);
nand U4994 (N_4994,In_1023,In_1289);
or U4995 (N_4995,In_1492,In_856);
and U4996 (N_4996,In_291,In_1203);
nor U4997 (N_4997,In_564,In_671);
nor U4998 (N_4998,In_1043,In_1178);
or U4999 (N_4999,In_398,In_1368);
nor U5000 (N_5000,N_960,N_2912);
nor U5001 (N_5001,N_907,N_2398);
or U5002 (N_5002,N_1593,N_305);
or U5003 (N_5003,N_2000,N_714);
and U5004 (N_5004,N_688,N_2184);
or U5005 (N_5005,N_211,N_2206);
nand U5006 (N_5006,N_1344,N_3240);
nand U5007 (N_5007,N_279,N_4635);
xor U5008 (N_5008,N_3972,N_4099);
nor U5009 (N_5009,N_3469,N_3505);
nor U5010 (N_5010,N_2710,N_4433);
and U5011 (N_5011,N_1499,N_1196);
and U5012 (N_5012,N_85,N_2343);
and U5013 (N_5013,N_940,N_2396);
nand U5014 (N_5014,N_1414,N_4638);
nand U5015 (N_5015,N_2285,N_3233);
or U5016 (N_5016,N_3190,N_1622);
nand U5017 (N_5017,N_3936,N_274);
nand U5018 (N_5018,N_2911,N_3485);
xor U5019 (N_5019,N_932,N_398);
nor U5020 (N_5020,N_1731,N_605);
or U5021 (N_5021,N_2445,N_1819);
nand U5022 (N_5022,N_4487,N_572);
nand U5023 (N_5023,N_1541,N_2957);
and U5024 (N_5024,N_1276,N_3804);
or U5025 (N_5025,N_942,N_1894);
nor U5026 (N_5026,N_4465,N_2501);
nor U5027 (N_5027,N_1476,N_4656);
or U5028 (N_5028,N_2632,N_510);
and U5029 (N_5029,N_2590,N_2741);
or U5030 (N_5030,N_1717,N_3313);
and U5031 (N_5031,N_854,N_4946);
nor U5032 (N_5032,N_1035,N_2769);
nand U5033 (N_5033,N_3203,N_1493);
or U5034 (N_5034,N_4663,N_4291);
nor U5035 (N_5035,N_1034,N_2047);
and U5036 (N_5036,N_2611,N_3929);
nand U5037 (N_5037,N_3149,N_3268);
nand U5038 (N_5038,N_3013,N_1869);
nand U5039 (N_5039,N_570,N_1084);
or U5040 (N_5040,N_338,N_1381);
nand U5041 (N_5041,N_2978,N_3780);
nand U5042 (N_5042,N_1867,N_4050);
or U5043 (N_5043,N_767,N_1413);
or U5044 (N_5044,N_2889,N_242);
nor U5045 (N_5045,N_2132,N_1854);
and U5046 (N_5046,N_2932,N_4300);
or U5047 (N_5047,N_2780,N_23);
nand U5048 (N_5048,N_4799,N_3810);
nand U5049 (N_5049,N_4596,N_2353);
or U5050 (N_5050,N_3223,N_2421);
and U5051 (N_5051,N_756,N_3718);
nand U5052 (N_5052,N_397,N_3974);
or U5053 (N_5053,N_353,N_2458);
xor U5054 (N_5054,N_3993,N_4254);
nand U5055 (N_5055,N_3822,N_1095);
nand U5056 (N_5056,N_1671,N_2467);
and U5057 (N_5057,N_2256,N_1912);
nor U5058 (N_5058,N_2393,N_896);
or U5059 (N_5059,N_4018,N_4074);
nor U5060 (N_5060,N_1324,N_525);
and U5061 (N_5061,N_342,N_2365);
xnor U5062 (N_5062,N_3747,N_562);
or U5063 (N_5063,N_4605,N_1401);
nor U5064 (N_5064,N_3062,N_797);
nand U5065 (N_5065,N_2158,N_3768);
and U5066 (N_5066,N_1159,N_4706);
and U5067 (N_5067,N_3510,N_1432);
and U5068 (N_5068,N_2255,N_1473);
and U5069 (N_5069,N_1467,N_1469);
nand U5070 (N_5070,N_3743,N_1966);
nand U5071 (N_5071,N_1422,N_410);
nand U5072 (N_5072,N_312,N_47);
or U5073 (N_5073,N_3776,N_2919);
nand U5074 (N_5074,N_3658,N_3181);
nand U5075 (N_5075,N_3388,N_108);
nand U5076 (N_5076,N_433,N_2341);
nand U5077 (N_5077,N_3597,N_1524);
and U5078 (N_5078,N_4174,N_2492);
or U5079 (N_5079,N_281,N_3899);
and U5080 (N_5080,N_2950,N_2301);
nor U5081 (N_5081,N_4841,N_4123);
and U5082 (N_5082,N_1345,N_1764);
nor U5083 (N_5083,N_4936,N_3507);
nor U5084 (N_5084,N_101,N_2112);
and U5085 (N_5085,N_2767,N_4741);
nor U5086 (N_5086,N_2007,N_4550);
and U5087 (N_5087,N_114,N_4118);
nand U5088 (N_5088,N_2391,N_3551);
or U5089 (N_5089,N_1069,N_3868);
and U5090 (N_5090,N_2991,N_4827);
nor U5091 (N_5091,N_4774,N_3148);
or U5092 (N_5092,N_2635,N_1694);
xor U5093 (N_5093,N_1817,N_1026);
nor U5094 (N_5094,N_3296,N_2736);
and U5095 (N_5095,N_2,N_2488);
nor U5096 (N_5096,N_841,N_2144);
nor U5097 (N_5097,N_3234,N_4055);
nor U5098 (N_5098,N_2753,N_1691);
or U5099 (N_5099,N_1318,N_3664);
and U5100 (N_5100,N_544,N_2977);
nor U5101 (N_5101,N_1763,N_2961);
or U5102 (N_5102,N_3947,N_591);
nor U5103 (N_5103,N_212,N_2561);
or U5104 (N_5104,N_1204,N_2350);
and U5105 (N_5105,N_4629,N_4366);
nor U5106 (N_5106,N_4928,N_3845);
or U5107 (N_5107,N_1194,N_2495);
and U5108 (N_5108,N_1531,N_2465);
nor U5109 (N_5109,N_2845,N_2665);
nand U5110 (N_5110,N_1279,N_2656);
and U5111 (N_5111,N_457,N_2661);
or U5112 (N_5112,N_1885,N_635);
or U5113 (N_5113,N_294,N_474);
nand U5114 (N_5114,N_939,N_3183);
nor U5115 (N_5115,N_1706,N_4937);
or U5116 (N_5116,N_4302,N_906);
or U5117 (N_5117,N_4468,N_676);
and U5118 (N_5118,N_4283,N_3809);
nand U5119 (N_5119,N_2581,N_1425);
nor U5120 (N_5120,N_1237,N_45);
or U5121 (N_5121,N_1559,N_1769);
or U5122 (N_5122,N_2213,N_1248);
nand U5123 (N_5123,N_1686,N_2096);
nand U5124 (N_5124,N_4747,N_284);
and U5125 (N_5125,N_412,N_3028);
or U5126 (N_5126,N_3905,N_3645);
nand U5127 (N_5127,N_3129,N_4627);
and U5128 (N_5128,N_3123,N_4671);
or U5129 (N_5129,N_1280,N_3343);
nand U5130 (N_5130,N_2062,N_1393);
and U5131 (N_5131,N_636,N_384);
nor U5132 (N_5132,N_4708,N_3686);
or U5133 (N_5133,N_2183,N_371);
and U5134 (N_5134,N_2810,N_3842);
nand U5135 (N_5135,N_1322,N_1709);
nand U5136 (N_5136,N_291,N_4733);
and U5137 (N_5137,N_1915,N_3039);
nor U5138 (N_5138,N_2960,N_4649);
nand U5139 (N_5139,N_1342,N_4617);
and U5140 (N_5140,N_3191,N_3833);
or U5141 (N_5141,N_1234,N_1967);
or U5142 (N_5142,N_2336,N_2615);
or U5143 (N_5143,N_646,N_2123);
nand U5144 (N_5144,N_1098,N_3592);
nand U5145 (N_5145,N_4316,N_566);
nor U5146 (N_5146,N_3133,N_251);
or U5147 (N_5147,N_2828,N_1121);
xnor U5148 (N_5148,N_574,N_1061);
nand U5149 (N_5149,N_3126,N_4453);
xor U5150 (N_5150,N_3187,N_780);
or U5151 (N_5151,N_2815,N_3047);
and U5152 (N_5152,N_4721,N_1019);
nor U5153 (N_5153,N_1562,N_2071);
nor U5154 (N_5154,N_2015,N_2189);
nand U5155 (N_5155,N_1742,N_243);
or U5156 (N_5156,N_1526,N_4507);
nand U5157 (N_5157,N_4492,N_4725);
nor U5158 (N_5158,N_3043,N_3050);
nor U5159 (N_5159,N_4409,N_1264);
and U5160 (N_5160,N_3695,N_2076);
or U5161 (N_5161,N_2918,N_1454);
and U5162 (N_5162,N_4272,N_1002);
or U5163 (N_5163,N_2633,N_3211);
nor U5164 (N_5164,N_186,N_3509);
nand U5165 (N_5165,N_2174,N_130);
and U5166 (N_5166,N_3475,N_3751);
nor U5167 (N_5167,N_4408,N_2239);
or U5168 (N_5168,N_496,N_3871);
nand U5169 (N_5169,N_1336,N_4510);
nand U5170 (N_5170,N_2622,N_2072);
nor U5171 (N_5171,N_2618,N_925);
nand U5172 (N_5172,N_58,N_4621);
xor U5173 (N_5173,N_4204,N_541);
nor U5174 (N_5174,N_4023,N_4684);
nand U5175 (N_5175,N_4518,N_1856);
nor U5176 (N_5176,N_375,N_3142);
or U5177 (N_5177,N_1827,N_4662);
nor U5178 (N_5178,N_4758,N_2716);
and U5179 (N_5179,N_909,N_3113);
or U5180 (N_5180,N_1337,N_1082);
or U5181 (N_5181,N_1387,N_3032);
nor U5182 (N_5182,N_886,N_4543);
nand U5183 (N_5183,N_1305,N_815);
xnor U5184 (N_5184,N_231,N_1704);
nor U5185 (N_5185,N_1652,N_4343);
nand U5186 (N_5186,N_4551,N_1618);
nor U5187 (N_5187,N_2657,N_3634);
or U5188 (N_5188,N_4223,N_824);
or U5189 (N_5189,N_4997,N_666);
or U5190 (N_5190,N_4368,N_3956);
and U5191 (N_5191,N_4083,N_4677);
and U5192 (N_5192,N_4440,N_911);
or U5193 (N_5193,N_97,N_3430);
and U5194 (N_5194,N_3463,N_1110);
or U5195 (N_5195,N_2087,N_3119);
and U5196 (N_5196,N_664,N_2502);
nand U5197 (N_5197,N_340,N_1078);
or U5198 (N_5198,N_3954,N_730);
or U5199 (N_5199,N_3428,N_3449);
nand U5200 (N_5200,N_1053,N_4009);
and U5201 (N_5201,N_1926,N_2326);
and U5202 (N_5202,N_2101,N_1996);
nor U5203 (N_5203,N_787,N_3609);
or U5204 (N_5204,N_4171,N_2329);
xor U5205 (N_5205,N_3086,N_807);
or U5206 (N_5206,N_2140,N_564);
nor U5207 (N_5207,N_2559,N_4398);
nor U5208 (N_5208,N_1537,N_3967);
nor U5209 (N_5209,N_2679,N_3228);
or U5210 (N_5210,N_4712,N_3624);
nand U5211 (N_5211,N_2200,N_2576);
and U5212 (N_5212,N_4734,N_3543);
and U5213 (N_5213,N_1215,N_1358);
nand U5214 (N_5214,N_2510,N_2457);
and U5215 (N_5215,N_3347,N_119);
nand U5216 (N_5216,N_3437,N_4380);
nand U5217 (N_5217,N_3051,N_3474);
nor U5218 (N_5218,N_506,N_1535);
and U5219 (N_5219,N_2781,N_3356);
nor U5220 (N_5220,N_4579,N_1891);
nor U5221 (N_5221,N_4274,N_13);
nor U5222 (N_5222,N_928,N_2658);
nor U5223 (N_5223,N_4867,N_3554);
nand U5224 (N_5224,N_1221,N_4650);
nor U5225 (N_5225,N_3452,N_4845);
nand U5226 (N_5226,N_4698,N_3851);
or U5227 (N_5227,N_3971,N_2592);
and U5228 (N_5228,N_172,N_2821);
nor U5229 (N_5229,N_568,N_3569);
nor U5230 (N_5230,N_2014,N_1605);
and U5231 (N_5231,N_2225,N_249);
and U5232 (N_5232,N_3275,N_3096);
nor U5233 (N_5233,N_2493,N_1573);
or U5234 (N_5234,N_3171,N_3647);
nand U5235 (N_5235,N_4224,N_513);
nor U5236 (N_5236,N_334,N_2727);
or U5237 (N_5237,N_3346,N_4842);
nand U5238 (N_5238,N_4,N_253);
nand U5239 (N_5239,N_148,N_2429);
and U5240 (N_5240,N_2253,N_2652);
nand U5241 (N_5241,N_4732,N_4945);
or U5242 (N_5242,N_4833,N_3828);
nor U5243 (N_5243,N_1792,N_4076);
and U5244 (N_5244,N_2704,N_1649);
and U5245 (N_5245,N_4080,N_3515);
xor U5246 (N_5246,N_764,N_4334);
or U5247 (N_5247,N_3873,N_1338);
nand U5248 (N_5248,N_2166,N_1630);
nor U5249 (N_5249,N_3359,N_2053);
nand U5250 (N_5250,N_3014,N_4971);
nor U5251 (N_5251,N_2690,N_453);
nor U5252 (N_5252,N_3716,N_1346);
xor U5253 (N_5253,N_961,N_4585);
nand U5254 (N_5254,N_2327,N_1602);
nand U5255 (N_5255,N_2317,N_2204);
nor U5256 (N_5256,N_2846,N_2552);
and U5257 (N_5257,N_2032,N_1699);
nand U5258 (N_5258,N_843,N_2411);
nor U5259 (N_5259,N_1989,N_4456);
and U5260 (N_5260,N_3154,N_4989);
nor U5261 (N_5261,N_4546,N_3182);
or U5262 (N_5262,N_1879,N_2039);
nand U5263 (N_5263,N_2049,N_875);
or U5264 (N_5264,N_4121,N_2593);
nor U5265 (N_5265,N_4280,N_1257);
xnor U5266 (N_5266,N_1375,N_163);
nand U5267 (N_5267,N_4960,N_522);
nor U5268 (N_5268,N_1529,N_2582);
or U5269 (N_5269,N_2278,N_1753);
or U5270 (N_5270,N_3710,N_4668);
nand U5271 (N_5271,N_4594,N_4378);
nand U5272 (N_5272,N_3859,N_3079);
and U5273 (N_5273,N_336,N_4476);
and U5274 (N_5274,N_2890,N_1635);
or U5275 (N_5275,N_1456,N_4081);
nor U5276 (N_5276,N_81,N_1673);
or U5277 (N_5277,N_4201,N_1423);
nor U5278 (N_5278,N_1240,N_2004);
or U5279 (N_5279,N_2086,N_885);
and U5280 (N_5280,N_3197,N_2237);
nand U5281 (N_5281,N_1052,N_723);
or U5282 (N_5282,N_1446,N_4643);
nor U5283 (N_5283,N_1849,N_3054);
or U5284 (N_5284,N_516,N_966);
nand U5285 (N_5285,N_1416,N_4069);
nor U5286 (N_5286,N_3403,N_483);
or U5287 (N_5287,N_3641,N_974);
and U5288 (N_5288,N_4640,N_2403);
and U5289 (N_5289,N_3324,N_3982);
nor U5290 (N_5290,N_4979,N_563);
and U5291 (N_5291,N_3961,N_2328);
xnor U5292 (N_5292,N_1255,N_2536);
and U5293 (N_5293,N_1860,N_2963);
and U5294 (N_5294,N_4349,N_2702);
nor U5295 (N_5295,N_1029,N_2740);
nor U5296 (N_5296,N_438,N_549);
or U5297 (N_5297,N_1356,N_341);
nand U5298 (N_5298,N_3254,N_2038);
and U5299 (N_5299,N_2010,N_3843);
and U5300 (N_5300,N_1700,N_1420);
nor U5301 (N_5301,N_3413,N_557);
nor U5302 (N_5302,N_1195,N_761);
and U5303 (N_5303,N_3351,N_2817);
or U5304 (N_5304,N_499,N_48);
nand U5305 (N_5305,N_3965,N_3422);
or U5306 (N_5306,N_4307,N_1654);
nor U5307 (N_5307,N_2532,N_1702);
nor U5308 (N_5308,N_4043,N_704);
or U5309 (N_5309,N_2137,N_4428);
and U5310 (N_5310,N_480,N_624);
nand U5311 (N_5311,N_3849,N_184);
nor U5312 (N_5312,N_2325,N_343);
or U5313 (N_5313,N_4450,N_4026);
nor U5314 (N_5314,N_1486,N_3745);
or U5315 (N_5315,N_3372,N_2527);
nand U5316 (N_5316,N_864,N_1408);
nor U5317 (N_5317,N_834,N_514);
nand U5318 (N_5318,N_112,N_4578);
nor U5319 (N_5319,N_3017,N_103);
nand U5320 (N_5320,N_290,N_4931);
nand U5321 (N_5321,N_4905,N_388);
and U5322 (N_5322,N_1517,N_486);
and U5323 (N_5323,N_1519,N_3375);
and U5324 (N_5324,N_2382,N_2566);
and U5325 (N_5325,N_2178,N_672);
nor U5326 (N_5326,N_140,N_1661);
or U5327 (N_5327,N_4147,N_1656);
and U5328 (N_5328,N_408,N_919);
nand U5329 (N_5329,N_3407,N_804);
or U5330 (N_5330,N_4369,N_1167);
nand U5331 (N_5331,N_3350,N_1211);
or U5332 (N_5332,N_4965,N_3756);
nor U5333 (N_5333,N_1871,N_3328);
nor U5334 (N_5334,N_3015,N_2884);
and U5335 (N_5335,N_4187,N_1491);
nor U5336 (N_5336,N_3753,N_1728);
nor U5337 (N_5337,N_973,N_1983);
or U5338 (N_5338,N_3614,N_645);
and U5339 (N_5339,N_2648,N_2612);
nand U5340 (N_5340,N_2944,N_2190);
nor U5341 (N_5341,N_3629,N_4743);
nor U5342 (N_5342,N_2587,N_4342);
nand U5343 (N_5343,N_759,N_4383);
nor U5344 (N_5344,N_2078,N_1311);
nand U5345 (N_5345,N_1880,N_856);
nand U5346 (N_5346,N_356,N_3262);
or U5347 (N_5347,N_3490,N_4319);
nand U5348 (N_5348,N_2337,N_1334);
and U5349 (N_5349,N_2029,N_4869);
nand U5350 (N_5350,N_2672,N_4815);
and U5351 (N_5351,N_3966,N_2787);
nor U5352 (N_5352,N_3646,N_2079);
and U5353 (N_5353,N_1837,N_2673);
or U5354 (N_5354,N_1489,N_4008);
nand U5355 (N_5355,N_302,N_3491);
nand U5356 (N_5356,N_3701,N_4568);
or U5357 (N_5357,N_2525,N_2820);
or U5358 (N_5358,N_4480,N_1757);
nor U5359 (N_5359,N_3620,N_3057);
nor U5360 (N_5360,N_4687,N_853);
nor U5361 (N_5361,N_1300,N_2866);
nand U5362 (N_5362,N_2496,N_414);
nor U5363 (N_5363,N_2943,N_1760);
nand U5364 (N_5364,N_4388,N_3378);
nand U5365 (N_5365,N_4211,N_1929);
nor U5366 (N_5366,N_4310,N_3406);
nand U5367 (N_5367,N_2872,N_3942);
and U5368 (N_5368,N_321,N_3029);
nand U5369 (N_5369,N_1203,N_2054);
or U5370 (N_5370,N_4589,N_2198);
and U5371 (N_5371,N_2099,N_1538);
nand U5372 (N_5372,N_2934,N_2640);
and U5373 (N_5373,N_4850,N_4049);
nand U5374 (N_5374,N_1758,N_3579);
and U5375 (N_5375,N_2695,N_1340);
or U5376 (N_5376,N_181,N_710);
nor U5377 (N_5377,N_4181,N_4315);
xnor U5378 (N_5378,N_2689,N_1406);
and U5379 (N_5379,N_1917,N_1135);
nor U5380 (N_5380,N_4113,N_4430);
nor U5381 (N_5381,N_4301,N_596);
nand U5382 (N_5382,N_581,N_4048);
and U5383 (N_5383,N_4710,N_2246);
and U5384 (N_5384,N_3145,N_2899);
nor U5385 (N_5385,N_2313,N_2708);
or U5386 (N_5386,N_4271,N_2138);
and U5387 (N_5387,N_3379,N_59);
nor U5388 (N_5388,N_3423,N_3411);
or U5389 (N_5389,N_2725,N_2993);
nor U5390 (N_5390,N_1374,N_1056);
xor U5391 (N_5391,N_3735,N_2916);
or U5392 (N_5392,N_3504,N_3933);
or U5393 (N_5393,N_283,N_2586);
nor U5394 (N_5394,N_4047,N_4017);
and U5395 (N_5395,N_390,N_2284);
nand U5396 (N_5396,N_3415,N_728);
xor U5397 (N_5397,N_3962,N_162);
nand U5398 (N_5398,N_4218,N_123);
xor U5399 (N_5399,N_4875,N_2220);
nand U5400 (N_5400,N_4107,N_944);
nand U5401 (N_5401,N_755,N_3559);
or U5402 (N_5402,N_1665,N_2425);
nand U5403 (N_5403,N_2745,N_1607);
nor U5404 (N_5404,N_871,N_1007);
and U5405 (N_5405,N_4358,N_3177);
or U5406 (N_5406,N_425,N_4179);
nand U5407 (N_5407,N_560,N_1364);
nand U5408 (N_5408,N_2942,N_105);
or U5409 (N_5409,N_3218,N_4679);
or U5410 (N_5410,N_1613,N_2992);
nand U5411 (N_5411,N_794,N_4266);
nand U5412 (N_5412,N_1615,N_1919);
and U5413 (N_5413,N_4004,N_2999);
and U5414 (N_5414,N_3545,N_923);
nor U5415 (N_5415,N_2152,N_3311);
xor U5416 (N_5416,N_372,N_151);
nand U5417 (N_5417,N_879,N_4691);
nor U5418 (N_5418,N_25,N_46);
nand U5419 (N_5419,N_3244,N_838);
and U5420 (N_5420,N_3730,N_392);
nand U5421 (N_5421,N_2830,N_1735);
nand U5422 (N_5422,N_3464,N_4911);
xor U5423 (N_5423,N_4096,N_1944);
and U5424 (N_5424,N_1465,N_4330);
nand U5425 (N_5425,N_1132,N_4292);
nand U5426 (N_5426,N_4950,N_111);
and U5427 (N_5427,N_1916,N_1292);
nand U5428 (N_5428,N_1036,N_3578);
nor U5429 (N_5429,N_3528,N_2876);
nand U5430 (N_5430,N_3713,N_1427);
or U5431 (N_5431,N_1624,N_4309);
and U5432 (N_5432,N_4336,N_2093);
nand U5433 (N_5433,N_232,N_1767);
and U5434 (N_5434,N_2869,N_1904);
and U5435 (N_5435,N_1128,N_1951);
nor U5436 (N_5436,N_1310,N_18);
nor U5437 (N_5437,N_1325,N_3402);
nor U5438 (N_5438,N_2913,N_4769);
nor U5439 (N_5439,N_275,N_2085);
and U5440 (N_5440,N_1554,N_4728);
or U5441 (N_5441,N_3370,N_3018);
or U5442 (N_5442,N_313,N_2895);
and U5443 (N_5443,N_2342,N_4630);
or U5444 (N_5444,N_4007,N_3848);
nand U5445 (N_5445,N_2692,N_3790);
nor U5446 (N_5446,N_1161,N_3793);
and U5447 (N_5447,N_902,N_2676);
nand U5448 (N_5448,N_2937,N_2173);
nand U5449 (N_5449,N_1302,N_2121);
or U5450 (N_5450,N_2797,N_4719);
or U5451 (N_5451,N_850,N_3976);
or U5452 (N_5452,N_3271,N_4759);
and U5453 (N_5453,N_3456,N_4750);
or U5454 (N_5454,N_1227,N_394);
nand U5455 (N_5455,N_1958,N_1129);
or U5456 (N_5456,N_4681,N_4901);
nand U5457 (N_5457,N_4455,N_3317);
or U5458 (N_5458,N_2251,N_1165);
and U5459 (N_5459,N_65,N_117);
or U5460 (N_5460,N_4933,N_1898);
or U5461 (N_5461,N_122,N_3761);
and U5462 (N_5462,N_1164,N_2075);
nand U5463 (N_5463,N_1137,N_191);
and U5464 (N_5464,N_943,N_4874);
nor U5465 (N_5465,N_3535,N_4119);
and U5466 (N_5466,N_2299,N_1126);
nand U5467 (N_5467,N_551,N_2726);
nand U5468 (N_5468,N_4894,N_550);
nor U5469 (N_5469,N_4548,N_3409);
nor U5470 (N_5470,N_2322,N_722);
and U5471 (N_5471,N_3516,N_863);
nand U5472 (N_5472,N_1755,N_2603);
nand U5473 (N_5473,N_362,N_4454);
or U5474 (N_5474,N_4431,N_4611);
nand U5475 (N_5475,N_3721,N_3533);
or U5476 (N_5476,N_1859,N_1587);
nor U5477 (N_5477,N_1960,N_4041);
nor U5478 (N_5478,N_1718,N_3255);
nand U5479 (N_5479,N_2385,N_619);
nand U5480 (N_5480,N_4614,N_3823);
and U5481 (N_5481,N_2435,N_3128);
nor U5482 (N_5482,N_4751,N_2363);
nor U5483 (N_5483,N_2258,N_2777);
and U5484 (N_5484,N_2987,N_4943);
nand U5485 (N_5485,N_1645,N_4192);
and U5486 (N_5486,N_169,N_154);
nor U5487 (N_5487,N_2296,N_2939);
nand U5488 (N_5488,N_796,N_2283);
and U5489 (N_5489,N_1277,N_1968);
nor U5490 (N_5490,N_4622,N_2844);
or U5491 (N_5491,N_1603,N_1044);
or U5492 (N_5492,N_3717,N_2017);
or U5493 (N_5493,N_1550,N_2288);
nand U5494 (N_5494,N_2677,N_4093);
or U5495 (N_5495,N_819,N_245);
or U5496 (N_5496,N_4406,N_344);
or U5497 (N_5497,N_3875,N_1059);
nor U5498 (N_5498,N_3151,N_1511);
and U5499 (N_5499,N_2683,N_1125);
nand U5500 (N_5500,N_3778,N_1555);
or U5501 (N_5501,N_3921,N_3937);
or U5502 (N_5502,N_369,N_3385);
nand U5503 (N_5503,N_3655,N_139);
or U5504 (N_5504,N_3295,N_4983);
nor U5505 (N_5505,N_4131,N_2335);
nand U5506 (N_5506,N_12,N_2444);
nor U5507 (N_5507,N_1313,N_507);
or U5508 (N_5508,N_1016,N_333);
and U5509 (N_5509,N_3907,N_4415);
nor U5510 (N_5510,N_2441,N_4626);
or U5511 (N_5511,N_183,N_489);
or U5512 (N_5512,N_2241,N_268);
and U5513 (N_5513,N_3021,N_1772);
xor U5514 (N_5514,N_1969,N_1395);
and U5515 (N_5515,N_3247,N_2238);
nor U5516 (N_5516,N_262,N_4222);
and U5517 (N_5517,N_2596,N_4318);
and U5518 (N_5518,N_1360,N_2949);
nor U5519 (N_5519,N_3251,N_2813);
or U5520 (N_5520,N_2759,N_360);
nor U5521 (N_5521,N_2623,N_4389);
nand U5522 (N_5522,N_725,N_1579);
nand U5523 (N_5523,N_4959,N_3282);
nor U5524 (N_5524,N_4367,N_2030);
or U5525 (N_5525,N_1014,N_3393);
or U5526 (N_5526,N_2808,N_1858);
nor U5527 (N_5527,N_4072,N_1887);
xnor U5528 (N_5528,N_1890,N_161);
nor U5529 (N_5529,N_2883,N_2020);
nand U5530 (N_5530,N_1546,N_1080);
and U5531 (N_5531,N_4860,N_2426);
or U5532 (N_5532,N_3539,N_1287);
xnor U5533 (N_5533,N_584,N_3118);
nor U5534 (N_5534,N_2698,N_2837);
and U5535 (N_5535,N_49,N_1747);
nand U5536 (N_5536,N_3630,N_504);
nand U5537 (N_5537,N_3769,N_2009);
or U5538 (N_5538,N_2264,N_4124);
nand U5539 (N_5539,N_3940,N_2036);
nand U5540 (N_5540,N_3417,N_617);
or U5541 (N_5541,N_4466,N_1878);
nand U5542 (N_5542,N_39,N_1123);
nor U5543 (N_5543,N_3911,N_1385);
nor U5544 (N_5544,N_2373,N_2712);
nor U5545 (N_5545,N_802,N_1862);
nand U5546 (N_5546,N_309,N_2616);
nor U5547 (N_5547,N_2271,N_2750);
and U5548 (N_5548,N_2369,N_3194);
nor U5549 (N_5549,N_3706,N_1484);
or U5550 (N_5550,N_862,N_175);
nor U5551 (N_5551,N_3134,N_213);
or U5552 (N_5552,N_1543,N_3335);
nor U5553 (N_5553,N_4806,N_196);
nand U5554 (N_5554,N_1807,N_857);
nand U5555 (N_5555,N_921,N_3781);
and U5556 (N_5556,N_4166,N_1533);
and U5557 (N_5557,N_790,N_4951);
and U5558 (N_5558,N_2168,N_1355);
nand U5559 (N_5559,N_2118,N_1662);
xnor U5560 (N_5560,N_2842,N_280);
nor U5561 (N_5561,N_2127,N_2824);
nand U5562 (N_5562,N_4436,N_538);
or U5563 (N_5563,N_3287,N_2768);
nand U5564 (N_5564,N_1687,N_3481);
nor U5565 (N_5565,N_1114,N_4267);
or U5566 (N_5566,N_1657,N_4159);
and U5567 (N_5567,N_2904,N_777);
nand U5568 (N_5568,N_3105,N_752);
and U5569 (N_5569,N_152,N_1291);
and U5570 (N_5570,N_4213,N_4108);
nor U5571 (N_5571,N_1365,N_4537);
or U5572 (N_5572,N_1810,N_731);
and U5573 (N_5573,N_427,N_4694);
nor U5574 (N_5574,N_2286,N_4574);
or U5575 (N_5575,N_331,N_318);
and U5576 (N_5576,N_3665,N_1112);
nor U5577 (N_5577,N_3532,N_2031);
nand U5578 (N_5578,N_2699,N_3836);
nand U5579 (N_5579,N_736,N_1761);
and U5580 (N_5580,N_1874,N_141);
or U5581 (N_5581,N_3957,N_825);
or U5582 (N_5582,N_289,N_604);
and U5583 (N_5583,N_56,N_3900);
nand U5584 (N_5584,N_4857,N_14);
nor U5585 (N_5585,N_40,N_2282);
or U5586 (N_5586,N_2671,N_2227);
and U5587 (N_5587,N_972,N_3323);
nand U5588 (N_5588,N_2356,N_4757);
and U5589 (N_5589,N_3772,N_1506);
nor U5590 (N_5590,N_783,N_200);
or U5591 (N_5591,N_980,N_3038);
nor U5592 (N_5592,N_3636,N_4844);
and U5593 (N_5593,N_1166,N_4985);
and U5594 (N_5594,N_545,N_269);
xnor U5595 (N_5595,N_3293,N_4296);
nor U5596 (N_5596,N_2858,N_4073);
or U5597 (N_5597,N_2498,N_4962);
nor U5598 (N_5598,N_4286,N_2188);
nand U5599 (N_5599,N_1048,N_623);
nand U5600 (N_5600,N_3765,N_2073);
nor U5601 (N_5601,N_659,N_2833);
and U5602 (N_5602,N_1818,N_4900);
nor U5603 (N_5603,N_3952,N_3691);
or U5604 (N_5604,N_3731,N_1189);
nand U5605 (N_5605,N_3130,N_1668);
xnor U5606 (N_5606,N_2314,N_4390);
and U5607 (N_5607,N_4344,N_4033);
nor U5608 (N_5608,N_4526,N_4898);
and U5609 (N_5609,N_490,N_4193);
nor U5610 (N_5610,N_2818,N_4412);
or U5611 (N_5611,N_2194,N_3153);
nand U5612 (N_5612,N_1501,N_1741);
or U5613 (N_5613,N_561,N_3360);
xnor U5614 (N_5614,N_3819,N_216);
nor U5615 (N_5615,N_4221,N_396);
or U5616 (N_5616,N_1928,N_3914);
nand U5617 (N_5617,N_1663,N_2097);
or U5618 (N_5618,N_1066,N_2482);
nand U5619 (N_5619,N_4553,N_772);
nor U5620 (N_5620,N_4419,N_1952);
nor U5621 (N_5621,N_2224,N_3264);
and U5622 (N_5622,N_4020,N_3377);
nand U5623 (N_5623,N_1974,N_1017);
nor U5624 (N_5624,N_4952,N_4233);
nor U5625 (N_5625,N_3818,N_1986);
nand U5626 (N_5626,N_3143,N_3310);
nand U5627 (N_5627,N_2856,N_4499);
nor U5628 (N_5628,N_1470,N_616);
nand U5629 (N_5629,N_1168,N_2643);
nor U5630 (N_5630,N_4981,N_3112);
nand U5631 (N_5631,N_4802,N_818);
nor U5632 (N_5632,N_2312,N_3520);
or U5633 (N_5633,N_3453,N_1238);
nor U5634 (N_5634,N_4354,N_2562);
or U5635 (N_5635,N_2423,N_4458);
nand U5636 (N_5636,N_368,N_1843);
nor U5637 (N_5637,N_4005,N_1680);
nor U5638 (N_5638,N_3684,N_4206);
nand U5639 (N_5639,N_4164,N_1963);
nor U5640 (N_5640,N_1099,N_3557);
or U5641 (N_5641,N_2909,N_179);
or U5642 (N_5642,N_2107,N_2816);
nand U5643 (N_5643,N_1873,N_4689);
or U5644 (N_5644,N_1339,N_985);
and U5645 (N_5645,N_4519,N_2167);
nand U5646 (N_5646,N_1461,N_2785);
and U5647 (N_5647,N_4573,N_2989);
nand U5648 (N_5648,N_4290,N_399);
nor U5649 (N_5649,N_2997,N_2878);
and U5650 (N_5650,N_826,N_4491);
nor U5651 (N_5651,N_3091,N_391);
or U5652 (N_5652,N_1627,N_346);
or U5653 (N_5653,N_1599,N_182);
nor U5654 (N_5654,N_4566,N_1480);
nand U5655 (N_5655,N_3755,N_263);
or U5656 (N_5656,N_478,N_2260);
or U5657 (N_5657,N_1721,N_3380);
and U5658 (N_5658,N_1949,N_1522);
nor U5659 (N_5659,N_4699,N_2066);
and U5660 (N_5660,N_1092,N_1651);
nor U5661 (N_5661,N_4256,N_3839);
nand U5662 (N_5662,N_4328,N_3139);
or U5663 (N_5663,N_4341,N_4794);
and U5664 (N_5664,N_4257,N_4459);
nand U5665 (N_5665,N_115,N_193);
and U5666 (N_5666,N_2799,N_3589);
nand U5667 (N_5667,N_4813,N_1601);
nand U5668 (N_5668,N_4592,N_1319);
nand U5669 (N_5669,N_3173,N_4958);
nor U5670 (N_5670,N_3944,N_4030);
nor U5671 (N_5671,N_2417,N_64);
nand U5672 (N_5672,N_3061,N_984);
and U5673 (N_5673,N_2022,N_3448);
xor U5674 (N_5674,N_611,N_4360);
nor U5675 (N_5675,N_2051,N_15);
and U5676 (N_5676,N_4565,N_1120);
or U5677 (N_5677,N_2257,N_2117);
nor U5678 (N_5678,N_3922,N_1122);
nor U5679 (N_5679,N_3176,N_1252);
or U5680 (N_5680,N_359,N_1836);
and U5681 (N_5681,N_240,N_3362);
nand U5682 (N_5682,N_3752,N_1389);
and U5683 (N_5683,N_1888,N_1284);
nor U5684 (N_5684,N_1188,N_4232);
or U5685 (N_5685,N_4209,N_4685);
or U5686 (N_5686,N_1049,N_2948);
and U5687 (N_5687,N_3482,N_606);
or U5688 (N_5688,N_1430,N_2693);
or U5689 (N_5689,N_4178,N_347);
or U5690 (N_5690,N_4253,N_3263);
nor U5691 (N_5691,N_317,N_435);
nor U5692 (N_5692,N_4146,N_3459);
nor U5693 (N_5693,N_3660,N_3342);
and U5694 (N_5694,N_4667,N_3441);
nand U5695 (N_5695,N_3910,N_4095);
nor U5696 (N_5696,N_136,N_2625);
or U5697 (N_5697,N_1710,N_1206);
nor U5698 (N_5698,N_3888,N_1421);
or U5699 (N_5699,N_1672,N_1833);
and U5700 (N_5700,N_1825,N_68);
xor U5701 (N_5701,N_1527,N_2215);
or U5702 (N_5702,N_1492,N_3103);
nand U5703 (N_5703,N_260,N_1471);
or U5704 (N_5704,N_2011,N_2788);
or U5705 (N_5705,N_4186,N_2794);
nand U5706 (N_5706,N_4243,N_4742);
nand U5707 (N_5707,N_2505,N_2792);
nand U5708 (N_5708,N_607,N_205);
nor U5709 (N_5709,N_4467,N_4683);
and U5710 (N_5710,N_2057,N_247);
nor U5711 (N_5711,N_1326,N_996);
nand U5712 (N_5712,N_4994,N_2428);
or U5713 (N_5713,N_3585,N_4333);
nand U5714 (N_5714,N_4035,N_1214);
nor U5715 (N_5715,N_3639,N_1169);
or U5716 (N_5716,N_1679,N_946);
or U5717 (N_5717,N_1695,N_3705);
nor U5718 (N_5718,N_3527,N_4184);
and U5719 (N_5719,N_1510,N_3110);
nor U5720 (N_5720,N_3626,N_3656);
xor U5721 (N_5721,N_4969,N_2668);
and U5722 (N_5722,N_3987,N_3135);
or U5723 (N_5723,N_2424,N_2068);
nor U5724 (N_5724,N_882,N_2080);
nand U5725 (N_5725,N_2060,N_2214);
nand U5726 (N_5726,N_2361,N_2277);
xor U5727 (N_5727,N_389,N_377);
nor U5728 (N_5728,N_3673,N_637);
nand U5729 (N_5729,N_1906,N_3092);
and U5730 (N_5730,N_1965,N_1544);
nand U5731 (N_5731,N_3283,N_3058);
and U5732 (N_5732,N_4980,N_2751);
nor U5733 (N_5733,N_2402,N_1160);
nor U5734 (N_5734,N_3975,N_4270);
xor U5735 (N_5735,N_4197,N_2406);
and U5736 (N_5736,N_1411,N_2468);
or U5737 (N_5737,N_3146,N_1868);
and U5738 (N_5738,N_3420,N_643);
nor U5739 (N_5739,N_4370,N_2706);
nand U5740 (N_5740,N_1784,N_2715);
and U5741 (N_5741,N_3855,N_2354);
xor U5742 (N_5742,N_367,N_2275);
and U5743 (N_5743,N_3089,N_4588);
and U5744 (N_5744,N_893,N_3261);
and U5745 (N_5745,N_1424,N_1771);
and U5746 (N_5746,N_2516,N_782);
and U5747 (N_5747,N_3298,N_3084);
and U5748 (N_5748,N_4474,N_3573);
or U5749 (N_5749,N_16,N_3120);
and U5750 (N_5750,N_2694,N_2538);
nand U5751 (N_5751,N_2857,N_1495);
and U5752 (N_5752,N_2849,N_1614);
and U5753 (N_5753,N_2442,N_4610);
or U5754 (N_5754,N_1391,N_4481);
nor U5755 (N_5755,N_3959,N_1634);
nor U5756 (N_5756,N_2392,N_2366);
nor U5757 (N_5757,N_4661,N_717);
and U5758 (N_5758,N_2548,N_4893);
or U5759 (N_5759,N_2739,N_1831);
nand U5760 (N_5760,N_4675,N_1127);
nor U5761 (N_5761,N_4002,N_534);
nor U5762 (N_5762,N_3983,N_4422);
nor U5763 (N_5763,N_1134,N_201);
nand U5764 (N_5764,N_3702,N_2854);
and U5765 (N_5765,N_4984,N_3644);
nor U5766 (N_5766,N_1233,N_322);
and U5767 (N_5767,N_3260,N_3410);
nor U5768 (N_5768,N_1520,N_4838);
and U5769 (N_5769,N_7,N_35);
nor U5770 (N_5770,N_4673,N_2059);
and U5771 (N_5771,N_2003,N_2655);
or U5772 (N_5772,N_1530,N_314);
and U5773 (N_5773,N_2383,N_3657);
or U5774 (N_5774,N_2945,N_1734);
and U5775 (N_5775,N_1643,N_2686);
or U5776 (N_5776,N_2801,N_3802);
nand U5777 (N_5777,N_2463,N_4495);
and U5778 (N_5778,N_424,N_2245);
or U5779 (N_5779,N_2547,N_649);
nor U5780 (N_5780,N_3229,N_1043);
xnor U5781 (N_5781,N_443,N_90);
or U5782 (N_5782,N_3085,N_891);
and U5783 (N_5783,N_332,N_4581);
or U5784 (N_5784,N_1925,N_4407);
or U5785 (N_5785,N_436,N_2451);
and U5786 (N_5786,N_2551,N_4167);
and U5787 (N_5787,N_4669,N_3497);
or U5788 (N_5788,N_4508,N_2489);
nand U5789 (N_5789,N_2958,N_555);
nand U5790 (N_5790,N_2554,N_2829);
nor U5791 (N_5791,N_4392,N_1088);
and U5792 (N_5792,N_2564,N_2631);
nor U5793 (N_5793,N_2520,N_4658);
nand U5794 (N_5794,N_660,N_1720);
nor U5795 (N_5795,N_3281,N_404);
and U5796 (N_5796,N_1903,N_2521);
xnor U5797 (N_5797,N_4273,N_670);
and U5798 (N_5798,N_847,N_2474);
nor U5799 (N_5799,N_2292,N_3209);
or U5800 (N_5800,N_386,N_1910);
nand U5801 (N_5801,N_4382,N_2931);
and U5802 (N_5802,N_3694,N_4245);
and U5803 (N_5803,N_2637,N_586);
or U5804 (N_5804,N_3016,N_3408);
or U5805 (N_5805,N_406,N_4834);
and U5806 (N_5806,N_2998,N_4281);
or U5807 (N_5807,N_1299,N_2279);
or U5808 (N_5808,N_2563,N_1131);
or U5809 (N_5809,N_4202,N_1964);
nor U5810 (N_5810,N_3912,N_2181);
or U5811 (N_5811,N_1172,N_2850);
and U5812 (N_5812,N_4264,N_518);
xnor U5813 (N_5813,N_4125,N_1895);
nand U5814 (N_5814,N_1021,N_4331);
nand U5815 (N_5815,N_814,N_1863);
or U5816 (N_5816,N_257,N_1178);
or U5817 (N_5817,N_2549,N_3575);
and U5818 (N_5818,N_613,N_2602);
nand U5819 (N_5819,N_1677,N_3893);
nand U5820 (N_5820,N_4421,N_2212);
or U5821 (N_5821,N_2100,N_2217);
nor U5822 (N_5822,N_3446,N_1115);
nand U5823 (N_5823,N_786,N_4314);
and U5824 (N_5824,N_1434,N_467);
nand U5825 (N_5825,N_3891,N_579);
or U5826 (N_5826,N_1405,N_798);
nor U5827 (N_5827,N_3945,N_1403);
and U5828 (N_5828,N_1813,N_4372);
nand U5829 (N_5829,N_4015,N_3250);
nor U5830 (N_5830,N_1354,N_4228);
and U5831 (N_5831,N_4356,N_4138);
nand U5832 (N_5832,N_4811,N_3265);
nand U5833 (N_5833,N_4282,N_3472);
or U5834 (N_5834,N_2310,N_958);
nand U5835 (N_5835,N_146,N_185);
nor U5836 (N_5836,N_1224,N_4556);
nand U5837 (N_5837,N_1972,N_2834);
or U5838 (N_5838,N_4864,N_63);
xor U5839 (N_5839,N_3447,N_3861);
or U5840 (N_5840,N_3434,N_55);
nand U5841 (N_5841,N_610,N_2139);
or U5842 (N_5842,N_4170,N_1959);
or U5843 (N_5843,N_3919,N_2272);
or U5844 (N_5844,N_1936,N_4540);
and U5845 (N_5845,N_3320,N_1433);
nor U5846 (N_5846,N_4584,N_2814);
nor U5847 (N_5847,N_4570,N_776);
nor U5848 (N_5848,N_2809,N_4926);
nor U5849 (N_5849,N_1223,N_2862);
nor U5850 (N_5850,N_3593,N_1343);
and U5851 (N_5851,N_4500,N_3894);
nand U5852 (N_5852,N_3538,N_3257);
nor U5853 (N_5853,N_1269,N_4022);
or U5854 (N_5854,N_3932,N_4129);
nor U5855 (N_5855,N_4966,N_3164);
nor U5856 (N_5856,N_2806,N_352);
or U5857 (N_5857,N_4284,N_1249);
nor U5858 (N_5858,N_1111,N_839);
and U5859 (N_5859,N_405,N_1620);
nand U5860 (N_5860,N_698,N_2843);
nor U5861 (N_5861,N_1632,N_3432);
nand U5862 (N_5862,N_821,N_701);
and U5863 (N_5863,N_4438,N_4098);
nand U5864 (N_5864,N_2268,N_2208);
and U5865 (N_5865,N_2147,N_4836);
nand U5866 (N_5866,N_4724,N_1273);
and U5867 (N_5867,N_1730,N_1886);
or U5868 (N_5868,N_1198,N_4446);
or U5869 (N_5869,N_2595,N_4880);
or U5870 (N_5870,N_4237,N_4930);
nand U5871 (N_5871,N_1384,N_4961);
nor U5872 (N_5872,N_2133,N_669);
or U5873 (N_5873,N_1568,N_3121);
and U5874 (N_5874,N_4917,N_3185);
nor U5875 (N_5875,N_1953,N_1621);
nand U5876 (N_5876,N_1497,N_393);
nand U5877 (N_5877,N_3941,N_2535);
and U5878 (N_5878,N_3580,N_187);
or U5879 (N_5879,N_1267,N_4249);
or U5880 (N_5880,N_2749,N_757);
nand U5881 (N_5881,N_3897,N_1191);
nand U5882 (N_5882,N_2569,N_53);
or U5883 (N_5883,N_4862,N_1766);
or U5884 (N_5884,N_3588,N_4242);
or U5885 (N_5885,N_264,N_1570);
nand U5886 (N_5886,N_840,N_2907);
nand U5887 (N_5887,N_3245,N_2419);
or U5888 (N_5888,N_3568,N_1816);
nand U5889 (N_5889,N_4820,N_3926);
nand U5890 (N_5890,N_2644,N_4297);
nand U5891 (N_5891,N_2236,N_1777);
and U5892 (N_5892,N_4071,N_4153);
and U5893 (N_5893,N_1504,N_4756);
or U5894 (N_5894,N_4066,N_4824);
nand U5895 (N_5895,N_4522,N_922);
or U5896 (N_5896,N_1847,N_3256);
and U5897 (N_5897,N_779,N_892);
xor U5898 (N_5898,N_1180,N_4177);
or U5899 (N_5899,N_4425,N_2311);
and U5900 (N_5900,N_4199,N_2321);
nor U5901 (N_5901,N_2868,N_3424);
and U5902 (N_5902,N_3786,N_2163);
nor U5903 (N_5903,N_224,N_4554);
nor U5904 (N_5904,N_598,N_1428);
nor U5905 (N_5905,N_4603,N_950);
and U5906 (N_5906,N_3920,N_3759);
or U5907 (N_5907,N_1994,N_4405);
nor U5908 (N_5908,N_3928,N_2742);
or U5909 (N_5909,N_4781,N_3106);
nor U5910 (N_5910,N_2882,N_1445);
nand U5911 (N_5911,N_376,N_4571);
nand U5912 (N_5912,N_4447,N_3027);
and U5913 (N_5913,N_1955,N_2688);
nand U5914 (N_5914,N_2307,N_543);
and U5915 (N_5915,N_878,N_3662);
nor U5916 (N_5916,N_2095,N_3276);
nand U5917 (N_5917,N_271,N_3663);
or U5918 (N_5918,N_460,N_1678);
nor U5919 (N_5919,N_3426,N_3565);
nor U5920 (N_5920,N_4702,N_2567);
and U5921 (N_5921,N_3570,N_1239);
nand U5922 (N_5922,N_463,N_3814);
nor U5923 (N_5923,N_3341,N_3345);
or U5924 (N_5924,N_2761,N_874);
and U5925 (N_5925,N_1236,N_683);
or U5926 (N_5926,N_3095,N_4896);
nand U5927 (N_5927,N_465,N_1558);
nand U5928 (N_5928,N_947,N_2550);
and U5929 (N_5929,N_3652,N_1838);
nor U5930 (N_5930,N_4881,N_1457);
or U5931 (N_5931,N_4766,N_2379);
nand U5932 (N_5932,N_2104,N_3358);
nand U5933 (N_5933,N_1083,N_107);
nor U5934 (N_5934,N_2043,N_2908);
or U5935 (N_5935,N_665,N_3688);
nor U5936 (N_5936,N_1108,N_1023);
nor U5937 (N_5937,N_524,N_1074);
and U5938 (N_5938,N_4285,N_3506);
nand U5939 (N_5939,N_4248,N_2136);
and U5940 (N_5940,N_2455,N_316);
or U5941 (N_5941,N_592,N_2915);
and U5942 (N_5942,N_1412,N_4101);
and U5943 (N_5943,N_1743,N_3239);
and U5944 (N_5944,N_737,N_1136);
and U5945 (N_5945,N_440,N_3450);
nand U5946 (N_5946,N_867,N_3219);
or U5947 (N_5947,N_1565,N_4337);
and U5948 (N_5948,N_4351,N_4745);
and U5949 (N_5949,N_3757,N_3080);
or U5950 (N_5950,N_639,N_501);
nor U5951 (N_5951,N_131,N_2165);
and U5952 (N_5952,N_3999,N_3315);
nand U5953 (N_5953,N_4157,N_4837);
and U5954 (N_5954,N_1481,N_1724);
and U5955 (N_5955,N_3692,N_238);
nor U5956 (N_5956,N_1145,N_4511);
or U5957 (N_5957,N_1357,N_2646);
and U5958 (N_5958,N_2935,N_3846);
nor U5959 (N_5959,N_3995,N_3078);
nand U5960 (N_5960,N_2760,N_4777);
and U5961 (N_5961,N_4940,N_3591);
and U5962 (N_5962,N_2826,N_2334);
and U5963 (N_5963,N_2146,N_2927);
xor U5964 (N_5964,N_533,N_2340);
or U5965 (N_5965,N_380,N_2585);
and U5966 (N_5966,N_2514,N_2629);
nand U5967 (N_5967,N_2624,N_1186);
or U5968 (N_5968,N_351,N_315);
nor U5969 (N_5969,N_1902,N_3290);
or U5970 (N_5970,N_1566,N_4778);
or U5971 (N_5971,N_866,N_3712);
or U5972 (N_5972,N_2177,N_789);
or U5973 (N_5973,N_1426,N_2831);
or U5974 (N_5974,N_2024,N_1485);
nand U5975 (N_5975,N_3221,N_28);
nor U5976 (N_5976,N_3476,N_1193);
or U5977 (N_5977,N_3337,N_477);
or U5978 (N_5978,N_1152,N_2378);
nor U5979 (N_5979,N_3198,N_2110);
nor U5980 (N_5980,N_4800,N_3649);
and U5981 (N_5981,N_1569,N_1512);
xor U5982 (N_5982,N_3333,N_3361);
nand U5983 (N_5983,N_2835,N_770);
or U5984 (N_5984,N_2764,N_4104);
and U5985 (N_5985,N_2323,N_4775);
nand U5986 (N_5986,N_27,N_512);
nor U5987 (N_5987,N_1750,N_1293);
or U5988 (N_5988,N_2302,N_4607);
nand U5989 (N_5989,N_3594,N_1939);
nor U5990 (N_5990,N_4053,N_3838);
and U5991 (N_5991,N_2231,N_774);
nand U5992 (N_5992,N_2270,N_1604);
and U5993 (N_5993,N_729,N_295);
nor U5994 (N_5994,N_199,N_2605);
and U5995 (N_5995,N_4916,N_3292);
or U5996 (N_5996,N_235,N_1435);
and U5997 (N_5997,N_2565,N_3724);
nand U5998 (N_5998,N_276,N_3460);
nand U5999 (N_5999,N_3461,N_937);
nand U6000 (N_6000,N_4180,N_62);
nand U6001 (N_6001,N_3405,N_2791);
and U6002 (N_6002,N_855,N_3704);
and U6003 (N_6003,N_3366,N_1363);
nand U6004 (N_6004,N_832,N_1260);
nor U6005 (N_6005,N_1812,N_349);
nor U6006 (N_6006,N_2647,N_600);
or U6007 (N_6007,N_237,N_3006);
nor U6008 (N_6008,N_3812,N_60);
nand U6009 (N_6009,N_3517,N_4582);
or U6010 (N_6010,N_1918,N_3479);
and U6011 (N_6011,N_4321,N_4039);
and U6012 (N_6012,N_1586,N_2344);
or U6013 (N_6013,N_3100,N_292);
and U6014 (N_6014,N_444,N_2440);
nor U6015 (N_6015,N_4402,N_3596);
nor U6016 (N_6016,N_962,N_325);
nor U6017 (N_6017,N_1674,N_653);
or U6018 (N_6018,N_3782,N_147);
nor U6019 (N_6019,N_4175,N_4934);
or U6020 (N_6020,N_1199,N_4371);
or U6021 (N_6021,N_2148,N_4915);
or U6022 (N_6022,N_3817,N_3374);
nand U6023 (N_6023,N_2412,N_2984);
or U6024 (N_6024,N_4416,N_93);
nand U6025 (N_6025,N_298,N_4657);
or U6026 (N_6026,N_4075,N_1396);
nor U6027 (N_6027,N_1472,N_1201);
and U6028 (N_6028,N_4261,N_1051);
or U6029 (N_6029,N_658,N_1013);
nand U6030 (N_6030,N_1085,N_4173);
and U6031 (N_6031,N_762,N_799);
nor U6032 (N_6032,N_1347,N_4317);
nor U6033 (N_6033,N_2717,N_527);
nor U6034 (N_6034,N_2259,N_2674);
and U6035 (N_6035,N_2263,N_1583);
and U6036 (N_6036,N_4196,N_1317);
nor U6037 (N_6037,N_92,N_3309);
nor U6038 (N_6038,N_1451,N_1245);
nor U6039 (N_6039,N_1528,N_1076);
or U6040 (N_6040,N_2533,N_1071);
nor U6041 (N_6041,N_956,N_4503);
nor U6042 (N_6042,N_1027,N_2626);
nand U6043 (N_6043,N_1025,N_3788);
and U6044 (N_6044,N_2384,N_2026);
nor U6045 (N_6045,N_582,N_3494);
and U6046 (N_6046,N_2867,N_155);
nor U6047 (N_6047,N_128,N_1417);
nand U6048 (N_6048,N_3386,N_991);
or U6049 (N_6049,N_2069,N_1258);
nor U6050 (N_6050,N_4498,N_2273);
and U6051 (N_6051,N_4355,N_986);
nor U6052 (N_6052,N_1946,N_3800);
or U6053 (N_6053,N_2464,N_3304);
or U6054 (N_6054,N_476,N_936);
or U6055 (N_6055,N_998,N_4214);
nor U6056 (N_6056,N_4413,N_4516);
nand U6057 (N_6057,N_976,N_4391);
nand U6058 (N_6058,N_3008,N_1640);
nor U6059 (N_6059,N_1884,N_3700);
or U6060 (N_6060,N_1398,N_1368);
nor U6061 (N_6061,N_2416,N_3623);
nor U6062 (N_6062,N_3404,N_3637);
and U6063 (N_6063,N_4364,N_3035);
nand U6064 (N_6064,N_2397,N_634);
nor U6065 (N_6065,N_1908,N_2627);
nor U6066 (N_6066,N_3220,N_1037);
nand U6067 (N_6067,N_3258,N_964);
nor U6068 (N_6068,N_1462,N_2923);
and U6069 (N_6069,N_1182,N_20);
or U6070 (N_6070,N_3699,N_4191);
and U6071 (N_6071,N_1503,N_1839);
nor U6072 (N_6072,N_2519,N_4060);
nand U6073 (N_6073,N_432,N_1577);
or U6074 (N_6074,N_2113,N_784);
xnor U6075 (N_6075,N_1183,N_3445);
nor U6076 (N_6076,N_1054,N_2303);
nand U6077 (N_6077,N_1975,N_1113);
nor U6078 (N_6078,N_3348,N_1697);
and U6079 (N_6079,N_3167,N_381);
nor U6080 (N_6080,N_2778,N_4918);
and U6081 (N_6081,N_3779,N_2933);
nor U6082 (N_6082,N_3034,N_873);
or U6083 (N_6083,N_2920,N_3950);
nand U6084 (N_6084,N_4814,N_3046);
nor U6085 (N_6085,N_1087,N_981);
and U6086 (N_6086,N_1392,N_2008);
and U6087 (N_6087,N_8,N_3205);
or U6088 (N_6088,N_1639,N_4103);
or U6089 (N_6089,N_3576,N_1961);
nand U6090 (N_6090,N_2436,N_747);
nand U6091 (N_6091,N_1509,N_1923);
xnor U6092 (N_6092,N_3053,N_1815);
or U6093 (N_6093,N_1229,N_4031);
nor U6094 (N_6094,N_1716,N_2023);
nand U6095 (N_6095,N_21,N_4133);
and U6096 (N_6096,N_4609,N_1582);
and U6097 (N_6097,N_3318,N_104);
nor U6098 (N_6098,N_3480,N_3763);
and U6099 (N_6099,N_145,N_2724);
or U6100 (N_6100,N_2490,N_2667);
and U6101 (N_6101,N_3856,N_2300);
nor U6102 (N_6102,N_3853,N_227);
nand U6103 (N_6103,N_4231,N_4532);
or U6104 (N_6104,N_441,N_3090);
nor U6105 (N_6105,N_1719,N_2701);
and U6106 (N_6106,N_3170,N_76);
nand U6107 (N_6107,N_3303,N_1576);
and U6108 (N_6108,N_2143,N_4942);
and U6109 (N_6109,N_109,N_2115);
nand U6110 (N_6110,N_434,N_3729);
nand U6111 (N_6111,N_3132,N_481);
nand U6112 (N_6112,N_2875,N_2291);
nand U6113 (N_6113,N_2111,N_2591);
or U6114 (N_6114,N_4087,N_3147);
nor U6115 (N_6115,N_3796,N_989);
xnor U6116 (N_6116,N_1752,N_4145);
nand U6117 (N_6117,N_2555,N_3454);
and U6118 (N_6118,N_3774,N_1625);
nor U6119 (N_6119,N_4575,N_266);
and U6120 (N_6120,N_915,N_3353);
or U6121 (N_6121,N_673,N_2600);
or U6122 (N_6122,N_3661,N_929);
and U6123 (N_6123,N_2359,N_4634);
and U6124 (N_6124,N_3117,N_1479);
nand U6125 (N_6125,N_509,N_3798);
and U6126 (N_6126,N_373,N_2013);
nor U6127 (N_6127,N_3502,N_576);
and U6128 (N_6128,N_3396,N_225);
and U6129 (N_6129,N_4736,N_740);
nor U6130 (N_6130,N_2798,N_734);
nand U6131 (N_6131,N_835,N_3943);
nor U6132 (N_6132,N_4381,N_706);
and U6133 (N_6133,N_2044,N_628);
or U6134 (N_6134,N_1231,N_4279);
nor U6135 (N_6135,N_2851,N_2229);
or U6136 (N_6136,N_2281,N_1285);
nand U6137 (N_6137,N_1006,N_2558);
nor U6138 (N_6138,N_2407,N_4863);
and U6139 (N_6139,N_3906,N_2475);
and U6140 (N_6140,N_953,N_1353);
nand U6141 (N_6141,N_3427,N_4670);
nor U6142 (N_6142,N_4250,N_3805);
or U6143 (N_6143,N_2659,N_3336);
nand U6144 (N_6144,N_121,N_2979);
or U6145 (N_6145,N_471,N_2719);
or U6146 (N_6146,N_3640,N_1438);
nand U6147 (N_6147,N_1840,N_3742);
nand U6148 (N_6148,N_935,N_4473);
and U6149 (N_6149,N_2332,N_1950);
or U6150 (N_6150,N_3770,N_4659);
nor U6151 (N_6151,N_4276,N_4873);
or U6152 (N_6152,N_4682,N_3994);
nor U6153 (N_6153,N_2471,N_3334);
nor U6154 (N_6154,N_3179,N_2094);
nor U6155 (N_6155,N_1447,N_51);
and U6156 (N_6156,N_3820,N_1140);
nand U6157 (N_6157,N_2386,N_2261);
and U6158 (N_6158,N_1725,N_3915);
nor U6159 (N_6159,N_3160,N_270);
and U6160 (N_6160,N_113,N_3202);
nand U6161 (N_6161,N_2364,N_1696);
or U6162 (N_6162,N_519,N_1118);
nor U6163 (N_6163,N_4737,N_3009);
nand U6164 (N_6164,N_4054,N_3002);
nand U6165 (N_6165,N_1090,N_2083);
nor U6166 (N_6166,N_4625,N_3274);
nor U6167 (N_6167,N_4379,N_2409);
or U6168 (N_6168,N_1441,N_3451);
nand U6169 (N_6169,N_4183,N_1633);
nor U6170 (N_6170,N_498,N_11);
xor U6171 (N_6171,N_2898,N_2210);
or U6172 (N_6172,N_3837,N_2848);
nand U6173 (N_6173,N_4132,N_1055);
nor U6174 (N_6174,N_708,N_1400);
or U6175 (N_6175,N_329,N_1213);
nand U6176 (N_6176,N_3892,N_978);
nor U6177 (N_6177,N_2287,N_2610);
xor U6178 (N_6178,N_4886,N_1588);
nor U6179 (N_6179,N_2812,N_1466);
nor U6180 (N_6180,N_1658,N_4789);
nor U6181 (N_6181,N_4059,N_1350);
or U6182 (N_6182,N_633,N_2233);
nand U6183 (N_6183,N_1957,N_778);
nor U6184 (N_6184,N_204,N_4796);
and U6185 (N_6185,N_748,N_1985);
and U6186 (N_6186,N_963,N_1726);
nor U6187 (N_6187,N_4326,N_2067);
nand U6188 (N_6188,N_387,N_10);
nor U6189 (N_6189,N_4818,N_72);
or U6190 (N_6190,N_1689,N_4822);
and U6191 (N_6191,N_2041,N_4717);
and U6192 (N_6192,N_4967,N_4090);
nor U6193 (N_6193,N_4497,N_4664);
and U6194 (N_6194,N_1796,N_4034);
nor U6195 (N_6195,N_1800,N_3196);
nand U6196 (N_6196,N_3340,N_1592);
nand U6197 (N_6197,N_3397,N_385);
xnor U6198 (N_6198,N_2775,N_1329);
or U6199 (N_6199,N_1521,N_402);
or U6200 (N_6200,N_2783,N_945);
nand U6201 (N_6201,N_4229,N_4996);
and U6202 (N_6202,N_3440,N_400);
nor U6203 (N_6203,N_2381,N_1684);
or U6204 (N_6204,N_727,N_4520);
and U6205 (N_6205,N_894,N_2352);
and U6206 (N_6206,N_4432,N_2265);
nor U6207 (N_6207,N_1042,N_469);
nor U6208 (N_6208,N_73,N_1294);
or U6209 (N_6209,N_1394,N_3563);
nor U6210 (N_6210,N_899,N_30);
nor U6211 (N_6211,N_95,N_2037);
and U6212 (N_6212,N_795,N_2308);
nor U6213 (N_6213,N_4651,N_449);
or U6214 (N_6214,N_1610,N_4924);
or U6215 (N_6215,N_949,N_3969);
or U6216 (N_6216,N_2331,N_1513);
or U6217 (N_6217,N_2172,N_788);
nor U6218 (N_6218,N_3433,N_3065);
nand U6219 (N_6219,N_3267,N_4395);
nand U6220 (N_6220,N_2274,N_500);
nor U6221 (N_6221,N_4070,N_4478);
and U6222 (N_6222,N_2330,N_703);
nand U6223 (N_6223,N_1653,N_1770);
or U6224 (N_6224,N_4361,N_214);
nand U6225 (N_6225,N_1105,N_4552);
nor U6226 (N_6226,N_4420,N_851);
and U6227 (N_6227,N_2929,N_1641);
nand U6228 (N_6228,N_4858,N_3394);
nand U6229 (N_6229,N_2216,N_3081);
nor U6230 (N_6230,N_3467,N_4780);
nand U6231 (N_6231,N_2243,N_3416);
nor U6232 (N_6232,N_99,N_2021);
and U6233 (N_6233,N_1970,N_775);
and U6234 (N_6234,N_1443,N_2388);
nor U6235 (N_6235,N_3314,N_2367);
nor U6236 (N_6236,N_4462,N_1244);
and U6237 (N_6237,N_4134,N_3217);
nand U6238 (N_6238,N_3622,N_1811);
nand U6239 (N_6239,N_2394,N_2804);
nand U6240 (N_6240,N_2295,N_4057);
nand U6241 (N_6241,N_4866,N_4776);
nand U6242 (N_6242,N_1463,N_2180);
and U6243 (N_6243,N_2770,N_1316);
nor U6244 (N_6244,N_3,N_2048);
or U6245 (N_6245,N_2150,N_1556);
or U6246 (N_6246,N_4225,N_1097);
and U6247 (N_6247,N_3550,N_4482);
nand U6248 (N_6248,N_2202,N_2664);
nand U6249 (N_6249,N_1039,N_1367);
nand U6250 (N_6250,N_959,N_2235);
or U6251 (N_6251,N_3012,N_890);
nand U6252 (N_6252,N_4993,N_4404);
and U6253 (N_6253,N_888,N_1314);
or U6254 (N_6254,N_4401,N_4632);
nand U6255 (N_6255,N_2634,N_4693);
nand U6256 (N_6256,N_3400,N_361);
or U6257 (N_6257,N_69,N_1217);
or U6258 (N_6258,N_2319,N_2946);
nor U6259 (N_6259,N_2106,N_256);
nor U6260 (N_6260,N_1289,N_2348);
nor U6261 (N_6261,N_1124,N_831);
and U6262 (N_6262,N_2090,N_2333);
nor U6263 (N_6263,N_2606,N_2447);
or U6264 (N_6264,N_771,N_3075);
and U6265 (N_6265,N_1263,N_900);
and U6266 (N_6266,N_702,N_192);
nor U6267 (N_6267,N_681,N_4642);
nand U6268 (N_6268,N_437,N_3390);
or U6269 (N_6269,N_4067,N_2669);
or U6270 (N_6270,N_1749,N_1834);
or U6271 (N_6271,N_2380,N_4703);
nand U6272 (N_6272,N_3462,N_2207);
nor U6273 (N_6273,N_2847,N_4365);
nand U6274 (N_6274,N_2575,N_3923);
nand U6275 (N_6275,N_4483,N_1516);
or U6276 (N_6276,N_526,N_2840);
nand U6277 (N_6277,N_430,N_3675);
nand U6278 (N_6278,N_3564,N_3518);
and U6279 (N_6279,N_918,N_1383);
and U6280 (N_6280,N_1712,N_3979);
and U6281 (N_6281,N_158,N_171);
xnor U6282 (N_6282,N_3666,N_920);
and U6283 (N_6283,N_3064,N_1778);
or U6284 (N_6284,N_1281,N_4114);
or U6285 (N_6285,N_2422,N_2737);
or U6286 (N_6286,N_3174,N_3094);
nand U6287 (N_6287,N_2731,N_1028);
and U6288 (N_6288,N_1606,N_2776);
and U6289 (N_6289,N_680,N_2653);
nor U6290 (N_6290,N_2155,N_2159);
or U6291 (N_6291,N_685,N_1564);
and U6292 (N_6292,N_195,N_3444);
xnor U6293 (N_6293,N_517,N_1736);
nor U6294 (N_6294,N_3574,N_1882);
or U6295 (N_6295,N_4514,N_699);
nand U6296 (N_6296,N_2405,N_2654);
and U6297 (N_6297,N_4531,N_3988);
and U6298 (N_6298,N_620,N_4890);
nand U6299 (N_6299,N_3500,N_4040);
nor U6300 (N_6300,N_2478,N_255);
or U6301 (N_6301,N_2711,N_3863);
or U6302 (N_6302,N_4618,N_1096);
and U6303 (N_6303,N_3124,N_3600);
nor U6304 (N_6304,N_3627,N_1759);
nor U6305 (N_6305,N_2452,N_2175);
or U6306 (N_6306,N_4149,N_4641);
or U6307 (N_6307,N_4308,N_210);
nand U6308 (N_6308,N_588,N_288);
nand U6309 (N_6309,N_1987,N_3749);
or U6310 (N_6310,N_2714,N_3732);
or U6311 (N_6311,N_134,N_3650);
nand U6312 (N_6312,N_2156,N_2103);
and U6313 (N_6313,N_3418,N_2395);
or U6314 (N_6314,N_3669,N_1241);
or U6315 (N_6315,N_462,N_4189);
nor U6316 (N_6316,N_38,N_4555);
or U6317 (N_6317,N_2758,N_1103);
or U6318 (N_6318,N_2670,N_1942);
and U6319 (N_6319,N_3881,N_3098);
or U6320 (N_6320,N_4889,N_1440);
nor U6321 (N_6321,N_521,N_642);
and U6322 (N_6322,N_4523,N_3189);
nor U6323 (N_6323,N_1372,N_4876);
nand U6324 (N_6324,N_4097,N_4953);
or U6325 (N_6325,N_3207,N_4956);
nand U6326 (N_6326,N_2506,N_765);
nor U6327 (N_6327,N_865,N_75);
nand U6328 (N_6328,N_2838,N_3758);
xor U6329 (N_6329,N_4387,N_355);
and U6330 (N_6330,N_3608,N_1832);
nor U6331 (N_6331,N_4128,N_1740);
and U6332 (N_6332,N_4493,N_4718);
nand U6333 (N_6333,N_738,N_2226);
nand U6334 (N_6334,N_938,N_2583);
nand U6335 (N_6335,N_4763,N_3726);
nor U6336 (N_6336,N_1765,N_3238);
xor U6337 (N_6337,N_472,N_2518);
nand U6338 (N_6338,N_2803,N_3784);
nor U6339 (N_6339,N_3056,N_350);
nor U6340 (N_6340,N_3044,N_2955);
and U6341 (N_6341,N_320,N_1927);
or U6342 (N_6342,N_3628,N_2205);
or U6343 (N_6343,N_2885,N_2924);
and U6344 (N_6344,N_2149,N_2720);
nand U6345 (N_6345,N_4722,N_655);
nand U6346 (N_6346,N_277,N_3069);
nor U6347 (N_6347,N_2619,N_4077);
or U6348 (N_6348,N_1793,N_995);
and U6349 (N_6349,N_2628,N_4839);
nand U6350 (N_6350,N_3037,N_2735);
or U6351 (N_6351,N_265,N_354);
and U6352 (N_6352,N_1222,N_3224);
nor U6353 (N_6353,N_2091,N_1295);
nor U6354 (N_6354,N_718,N_599);
or U6355 (N_6355,N_4696,N_532);
nand U6356 (N_6356,N_4707,N_656);
and U6357 (N_6357,N_2604,N_4140);
nor U6358 (N_6358,N_3373,N_1);
nor U6359 (N_6359,N_4230,N_70);
xor U6360 (N_6360,N_2511,N_37);
or U6361 (N_6361,N_4828,N_1349);
and U6362 (N_6362,N_2990,N_2721);
nand U6363 (N_6363,N_567,N_1179);
nor U6364 (N_6364,N_905,N_1359);
nor U6365 (N_6365,N_470,N_1275);
or U6366 (N_6366,N_1595,N_2347);
or U6367 (N_6367,N_2589,N_1841);
and U6368 (N_6368,N_1616,N_209);
nor U6369 (N_6369,N_2560,N_3567);
nor U6370 (N_6370,N_4779,N_2460);
or U6371 (N_6371,N_812,N_3890);
nand U6372 (N_6372,N_1664,N_4720);
nand U6373 (N_6373,N_466,N_1914);
nand U6374 (N_6374,N_29,N_4788);
xor U6375 (N_6375,N_178,N_2746);
and U6376 (N_6376,N_6,N_3011);
nor U6377 (N_6377,N_2128,N_2196);
nand U6378 (N_6378,N_828,N_4086);
or U6379 (N_6379,N_1081,N_2675);
nor U6380 (N_6380,N_1988,N_4835);
or U6381 (N_6381,N_2450,N_4016);
and U6382 (N_6382,N_3052,N_2052);
nor U6383 (N_6383,N_4783,N_80);
xnor U6384 (N_6384,N_1508,N_306);
nand U6385 (N_6385,N_2968,N_4932);
and U6386 (N_6386,N_4567,N_1872);
nor U6387 (N_6387,N_1209,N_2537);
or U6388 (N_6388,N_4028,N_2608);
nand U6389 (N_6389,N_3331,N_4037);
or U6390 (N_6390,N_668,N_459);
nand U6391 (N_6391,N_173,N_503);
nor U6392 (N_6392,N_36,N_4155);
nand U6393 (N_6393,N_971,N_4359);
nor U6394 (N_6394,N_3719,N_594);
xor U6395 (N_6395,N_4084,N_1612);
xor U6396 (N_6396,N_421,N_988);
nor U6397 (N_6397,N_2201,N_3213);
and U6398 (N_6398,N_3111,N_2360);
nand U6399 (N_6399,N_2903,N_3059);
and U6400 (N_6400,N_4226,N_383);
and U6401 (N_6401,N_4348,N_3076);
nand U6402 (N_6402,N_3231,N_2171);
nor U6403 (N_6403,N_1773,N_4185);
xor U6404 (N_6404,N_407,N_2345);
or U6405 (N_6405,N_3338,N_222);
nand U6406 (N_6406,N_4562,N_2119);
or U6407 (N_6407,N_3486,N_4907);
and U6408 (N_6408,N_4660,N_697);
nor U6409 (N_6409,N_3184,N_1312);
nand U6410 (N_6410,N_2515,N_817);
or U6411 (N_6411,N_2448,N_2620);
nor U6412 (N_6412,N_3246,N_715);
nor U6413 (N_6413,N_3741,N_1732);
nand U6414 (N_6414,N_1032,N_4429);
nand U6415 (N_6415,N_2546,N_2028);
and U6416 (N_6416,N_3156,N_4019);
and U6417 (N_6417,N_4560,N_2871);
nand U6418 (N_6418,N_3201,N_3266);
nand U6419 (N_6419,N_3236,N_3439);
nand U6420 (N_6420,N_3895,N_1722);
nor U6421 (N_6421,N_479,N_3562);
nand U6422 (N_6422,N_4740,N_217);
and U6423 (N_6423,N_2557,N_2940);
nand U6424 (N_6424,N_1038,N_33);
nor U6425 (N_6425,N_3468,N_3082);
or U6426 (N_6426,N_3670,N_2980);
nand U6427 (N_6427,N_1711,N_3777);
and U6428 (N_6428,N_4269,N_3206);
or U6429 (N_6429,N_3243,N_4909);
or U6430 (N_6430,N_712,N_2002);
nor U6431 (N_6431,N_684,N_2240);
or U6432 (N_6432,N_1990,N_3010);
or U6433 (N_6433,N_735,N_4678);
and U6434 (N_6434,N_2088,N_102);
or U6435 (N_6435,N_2568,N_411);
nand U6436 (N_6436,N_1971,N_4829);
and U6437 (N_6437,N_2861,N_2921);
nand U6438 (N_6438,N_638,N_2304);
nor U6439 (N_6439,N_301,N_482);
or U6440 (N_6440,N_515,N_742);
nor U6441 (N_6441,N_931,N_3097);
or U6442 (N_6442,N_464,N_3556);
or U6443 (N_6443,N_4156,N_1956);
and U6444 (N_6444,N_3714,N_3114);
nand U6445 (N_6445,N_785,N_4885);
and U6446 (N_6446,N_4418,N_2485);
and U6447 (N_6447,N_2164,N_849);
nor U6448 (N_6448,N_4338,N_468);
nand U6449 (N_6449,N_4606,N_3767);
nand U6450 (N_6450,N_382,N_4505);
nand U6451 (N_6451,N_2193,N_805);
xnor U6452 (N_6452,N_2389,N_2476);
or U6453 (N_6453,N_1141,N_261);
and U6454 (N_6454,N_1567,N_1738);
nand U6455 (N_6455,N_4215,N_678);
and U6456 (N_6456,N_4115,N_3775);
and U6457 (N_6457,N_4572,N_1532);
and U6458 (N_6458,N_4539,N_887);
nand U6459 (N_6459,N_913,N_1682);
or U6460 (N_6460,N_1623,N_4152);
or U6461 (N_6461,N_2836,N_4288);
and U6462 (N_6462,N_4340,N_4879);
and U6463 (N_6463,N_4987,N_4052);
and U6464 (N_6464,N_3709,N_982);
nand U6465 (N_6465,N_2199,N_4804);
nor U6466 (N_6466,N_3680,N_1176);
or U6467 (N_6467,N_2880,N_4921);
nand U6468 (N_6468,N_2542,N_3939);
nand U6469 (N_6469,N_667,N_4161);
and U6470 (N_6470,N_2754,N_3161);
nand U6471 (N_6471,N_2786,N_220);
nand U6472 (N_6472,N_448,N_1144);
nor U6473 (N_6473,N_3889,N_1327);
nand U6474 (N_6474,N_640,N_1482);
and U6475 (N_6475,N_4927,N_3738);
nand U6476 (N_6476,N_3549,N_2700);
nand U6477 (N_6477,N_2160,N_1271);
nor U6478 (N_6478,N_2800,N_2762);
nand U6479 (N_6479,N_1943,N_3330);
or U6480 (N_6480,N_2186,N_626);
nor U6481 (N_6481,N_2621,N_3740);
or U6482 (N_6482,N_3023,N_1745);
and U6483 (N_6483,N_1619,N_2431);
nand U6484 (N_6484,N_751,N_2045);
nand U6485 (N_6485,N_160,N_1094);
and U6486 (N_6486,N_3791,N_4812);
or U6487 (N_6487,N_1617,N_4964);
or U6488 (N_6488,N_3525,N_3832);
or U6489 (N_6489,N_1794,N_709);
and U6490 (N_6490,N_1776,N_2454);
nor U6491 (N_6491,N_3305,N_4819);
nand U6492 (N_6492,N_1308,N_4599);
and U6493 (N_6493,N_4832,N_1638);
nor U6494 (N_6494,N_1133,N_852);
or U6495 (N_6495,N_3116,N_2477);
and U6496 (N_6496,N_3270,N_1881);
or U6497 (N_6497,N_2779,N_2211);
and U6498 (N_6498,N_1478,N_4252);
and U6499 (N_6499,N_3511,N_285);
nor U6500 (N_6500,N_3301,N_2374);
nor U6501 (N_6501,N_1003,N_4127);
or U6502 (N_6502,N_733,N_3866);
nor U6503 (N_6503,N_1937,N_335);
nor U6504 (N_6504,N_1751,N_4258);
or U6505 (N_6505,N_1729,N_3806);
and U6506 (N_6506,N_4126,N_1060);
and U6507 (N_6507,N_1298,N_569);
nor U6508 (N_6508,N_4293,N_2470);
nand U6509 (N_6509,N_2182,N_3631);
or U6510 (N_6510,N_1388,N_100);
or U6511 (N_6511,N_2294,N_3876);
and U6512 (N_6512,N_3799,N_4219);
and U6513 (N_6513,N_230,N_3632);
nand U6514 (N_6514,N_3241,N_3074);
nor U6515 (N_6515,N_1723,N_3958);
and U6516 (N_6516,N_4488,N_415);
or U6517 (N_6517,N_2154,N_4393);
or U6518 (N_6518,N_2131,N_3960);
or U6519 (N_6519,N_3455,N_769);
and U6520 (N_6520,N_1219,N_4329);
or U6521 (N_6521,N_3087,N_22);
nand U6522 (N_6522,N_773,N_153);
nand U6523 (N_6523,N_3141,N_3431);
or U6524 (N_6524,N_2642,N_3093);
nand U6525 (N_6525,N_2084,N_4753);
or U6526 (N_6526,N_4424,N_2873);
and U6527 (N_6527,N_1998,N_2161);
or U6528 (N_6528,N_1659,N_4345);
xnor U6529 (N_6529,N_2996,N_150);
nand U6530 (N_6530,N_4322,N_4490);
xor U6531 (N_6531,N_78,N_1250);
or U6532 (N_6532,N_1660,N_3115);
and U6533 (N_6533,N_1708,N_4790);
nor U6534 (N_6534,N_4452,N_1611);
and U6535 (N_6535,N_2305,N_1306);
nor U6536 (N_6536,N_845,N_4029);
nor U6537 (N_6537,N_4613,N_3948);
and U6538 (N_6538,N_110,N_2784);
and U6539 (N_6539,N_2324,N_168);
and U6540 (N_6540,N_1041,N_3953);
nor U6541 (N_6541,N_1851,N_4762);
nor U6542 (N_6542,N_3750,N_3615);
nor U6543 (N_6543,N_4711,N_89);
or U6544 (N_6544,N_1386,N_565);
nand U6545 (N_6545,N_2179,N_3371);
nor U6546 (N_6546,N_967,N_547);
nor U6547 (N_6547,N_493,N_3659);
and U6548 (N_6548,N_2930,N_3934);
nor U6549 (N_6549,N_4470,N_4032);
or U6550 (N_6550,N_2744,N_1155);
and U6551 (N_6551,N_1688,N_4558);
and U6552 (N_6552,N_1235,N_4376);
or U6553 (N_6553,N_4448,N_952);
and U6554 (N_6554,N_74,N_1870);
nor U6555 (N_6555,N_4580,N_194);
or U6556 (N_6556,N_4840,N_1626);
nand U6557 (N_6557,N_1089,N_418);
and U6558 (N_6558,N_1429,N_3235);
or U6559 (N_6559,N_2687,N_1139);
and U6560 (N_6560,N_451,N_2748);
nor U6561 (N_6561,N_4854,N_2601);
nor U6562 (N_6562,N_1265,N_132);
nor U6563 (N_6563,N_884,N_1507);
nand U6564 (N_6564,N_1119,N_4972);
nor U6565 (N_6565,N_3369,N_627);
xor U6566 (N_6566,N_1185,N_1181);
nor U6567 (N_6567,N_2938,N_3259);
nand U6568 (N_6568,N_916,N_1572);
xor U6569 (N_6569,N_1288,N_2439);
xor U6570 (N_6570,N_3821,N_1913);
nand U6571 (N_6571,N_2645,N_4882);
or U6572 (N_6572,N_4373,N_3544);
nand U6573 (N_6573,N_3807,N_2040);
and U6574 (N_6574,N_4849,N_395);
or U6575 (N_6575,N_1012,N_1845);
nand U6576 (N_6576,N_3916,N_3395);
nor U6577 (N_6577,N_4731,N_4111);
nand U6578 (N_6578,N_79,N_4012);
and U6579 (N_6579,N_3860,N_3158);
nor U6580 (N_6580,N_868,N_3192);
and U6581 (N_6581,N_711,N_2375);
and U6582 (N_6582,N_1842,N_3604);
or U6583 (N_6583,N_4765,N_4871);
nand U6584 (N_6584,N_96,N_287);
and U6585 (N_6585,N_1628,N_3357);
nand U6586 (N_6586,N_2034,N_4091);
or U6587 (N_6587,N_3571,N_423);
or U6588 (N_6588,N_1707,N_2796);
and U6589 (N_6589,N_1399,N_3883);
xnor U6590 (N_6590,N_3438,N_2681);
nor U6591 (N_6591,N_3489,N_4730);
and U6592 (N_6592,N_4892,N_1924);
nand U6593 (N_6593,N_1001,N_1954);
nor U6594 (N_6594,N_4615,N_159);
and U6595 (N_6595,N_3734,N_3984);
or U6596 (N_6596,N_4200,N_1676);
and U6597 (N_6597,N_4247,N_4198);
or U6598 (N_6598,N_229,N_2947);
xor U6599 (N_6599,N_4709,N_228);
nor U6600 (N_6600,N_3722,N_993);
or U6601 (N_6601,N_4944,N_1590);
or U6602 (N_6602,N_4141,N_3200);
xor U6603 (N_6603,N_1251,N_2556);
nand U6604 (N_6604,N_202,N_4920);
or U6605 (N_6605,N_1116,N_4764);
and U6606 (N_6606,N_4212,N_4461);
and U6607 (N_6607,N_4922,N_1202);
and U6608 (N_6608,N_3466,N_4925);
or U6609 (N_6609,N_833,N_3909);
and U6610 (N_6610,N_1666,N_4652);
nand U6611 (N_6611,N_2599,N_4485);
or U6612 (N_6612,N_3697,N_2680);
nand U6613 (N_6613,N_1629,N_2487);
or U6614 (N_6614,N_4760,N_3617);
nor U6615 (N_6615,N_3547,N_3762);
nor U6616 (N_6616,N_1941,N_165);
nor U6617 (N_6617,N_2896,N_2793);
or U6618 (N_6618,N_4100,N_1575);
and U6619 (N_6619,N_4888,N_450);
nor U6620 (N_6620,N_1597,N_508);
nand U6621 (N_6621,N_3389,N_3887);
nor U6622 (N_6622,N_1230,N_1210);
nand U6623 (N_6623,N_955,N_2362);
nor U6624 (N_6624,N_693,N_3760);
or U6625 (N_6625,N_1008,N_1900);
or U6626 (N_6626,N_2771,N_837);
or U6627 (N_6627,N_4535,N_4062);
and U6628 (N_6628,N_2176,N_3917);
nor U6629 (N_6629,N_4512,N_3381);
nor U6630 (N_6630,N_4471,N_1174);
nor U6631 (N_6631,N_1149,N_2819);
nand U6632 (N_6632,N_883,N_116);
and U6633 (N_6633,N_2928,N_374);
nor U6634 (N_6634,N_721,N_189);
nand U6635 (N_6635,N_1820,N_810);
nand U6636 (N_6636,N_4595,N_914);
and U6637 (N_6637,N_2058,N_3850);
or U6638 (N_6638,N_4645,N_167);
or U6639 (N_6639,N_948,N_2124);
nor U6640 (N_6640,N_1783,N_2976);
or U6641 (N_6641,N_641,N_632);
and U6642 (N_6642,N_1670,N_750);
xnor U6643 (N_6643,N_3297,N_1216);
or U6644 (N_6644,N_2483,N_3042);
and U6645 (N_6645,N_2089,N_4908);
nand U6646 (N_6646,N_1713,N_910);
and U6647 (N_6647,N_2863,N_2427);
nand U6648 (N_6648,N_2580,N_4752);
nor U6649 (N_6649,N_2922,N_4809);
or U6650 (N_6650,N_442,N_2526);
and U6651 (N_6651,N_3827,N_4304);
nor U6652 (N_6652,N_4102,N_1321);
xor U6653 (N_6653,N_1073,N_3553);
and U6654 (N_6654,N_1683,N_3152);
nor U6655 (N_6655,N_2639,N_3526);
and U6656 (N_6656,N_2432,N_2728);
and U6657 (N_6657,N_2953,N_741);
nand U6658 (N_6658,N_3473,N_4165);
or U6659 (N_6659,N_3376,N_2982);
nand U6660 (N_6660,N_3870,N_3540);
or U6661 (N_6661,N_2678,N_4851);
nor U6662 (N_6662,N_889,N_2108);
nor U6663 (N_6663,N_3107,N_2415);
nor U6664 (N_6664,N_1775,N_732);
nand U6665 (N_6665,N_4955,N_2975);
or U6666 (N_6666,N_766,N_297);
nor U6667 (N_6667,N_743,N_2832);
and U6668 (N_6668,N_2666,N_1637);
nand U6669 (N_6669,N_4895,N_1331);
and U6670 (N_6670,N_118,N_4569);
and U6671 (N_6671,N_1005,N_3162);
and U6672 (N_6672,N_1589,N_535);
or U6673 (N_6673,N_1040,N_4092);
or U6674 (N_6674,N_1242,N_1864);
and U6675 (N_6675,N_926,N_1004);
nor U6676 (N_6676,N_3679,N_3172);
nand U6677 (N_6677,N_3099,N_2774);
or U6678 (N_6678,N_2906,N_3072);
nand U6679 (N_6679,N_1278,N_4808);
nand U6680 (N_6680,N_758,N_3789);
or U6681 (N_6681,N_4089,N_4078);
and U6682 (N_6682,N_250,N_2508);
or U6683 (N_6683,N_1899,N_4463);
or U6684 (N_6684,N_603,N_3421);
and U6685 (N_6685,N_2500,N_2481);
nor U6686 (N_6686,N_3980,N_2855);
nor U6687 (N_6687,N_583,N_530);
or U6688 (N_6688,N_4021,N_4220);
and U6689 (N_6689,N_4210,N_4823);
nor U6690 (N_6690,N_3278,N_4639);
nor U6691 (N_6691,N_3896,N_650);
nor U6692 (N_6692,N_278,N_330);
and U6693 (N_6693,N_2531,N_2368);
nor U6694 (N_6694,N_4767,N_4616);
nand U6695 (N_6695,N_1448,N_2660);
or U6696 (N_6696,N_491,N_3443);
and U6697 (N_6697,N_3606,N_686);
or U6698 (N_6698,N_2480,N_3964);
nor U6699 (N_6699,N_1130,N_2722);
and U6700 (N_6700,N_3436,N_705);
or U6701 (N_6701,N_601,N_1207);
nor U6702 (N_6702,N_417,N_3852);
nor U6703 (N_6703,N_2479,N_452);
nand U6704 (N_6704,N_3648,N_2607);
nor U6705 (N_6705,N_2266,N_2614);
or U6706 (N_6706,N_2346,N_1940);
or U6707 (N_6707,N_4506,N_1156);
nor U6708 (N_6708,N_1650,N_1142);
nand U6709 (N_6709,N_662,N_233);
or U6710 (N_6710,N_2747,N_3289);
nor U6711 (N_6711,N_2517,N_4238);
and U6712 (N_6712,N_4715,N_4674);
or U6713 (N_6713,N_422,N_2573);
nand U6714 (N_6714,N_239,N_3854);
nand U6715 (N_6715,N_3465,N_1050);
and U6716 (N_6716,N_2588,N_2859);
or U6717 (N_6717,N_1797,N_3633);
and U6718 (N_6718,N_1801,N_1453);
and U6719 (N_6719,N_1058,N_4998);
or U6720 (N_6720,N_2153,N_1931);
or U6721 (N_6721,N_1536,N_3577);
nand U6722 (N_6722,N_4992,N_1477);
and U6723 (N_6723,N_4312,N_1107);
and U6724 (N_6724,N_4163,N_3685);
or U6725 (N_6725,N_4870,N_3419);
nand U6726 (N_6726,N_3248,N_1578);
nor U6727 (N_6727,N_2061,N_679);
nor U6728 (N_6728,N_3985,N_2893);
nor U6729 (N_6729,N_2881,N_4504);
or U6730 (N_6730,N_1525,N_4109);
and U6731 (N_6731,N_3908,N_4003);
and U6732 (N_6732,N_4729,N_3867);
nand U6733 (N_6733,N_571,N_2042);
and U6734 (N_6734,N_691,N_1853);
or U6735 (N_6735,N_1380,N_324);
nor U6736 (N_6736,N_2755,N_4137);
nand U6737 (N_6737,N_618,N_2376);
and U6738 (N_6738,N_877,N_3387);
and U6739 (N_6739,N_2125,N_4417);
or U6740 (N_6740,N_1973,N_3232);
and U6741 (N_6741,N_4486,N_4919);
and U6742 (N_6742,N_4122,N_143);
nor U6743 (N_6743,N_2966,N_4528);
nand U6744 (N_6744,N_3253,N_3070);
nor U6745 (N_6745,N_2250,N_3088);
nand U6746 (N_6746,N_2636,N_4362);
nand U6747 (N_6747,N_3973,N_2732);
nand U6748 (N_6748,N_4843,N_3901);
and U6749 (N_6749,N_745,N_2597);
or U6750 (N_6750,N_768,N_127);
nor U6751 (N_6751,N_2290,N_2703);
nand U6752 (N_6752,N_2905,N_1212);
nor U6753 (N_6753,N_1826,N_3215);
or U6754 (N_6754,N_4644,N_677);
or U6755 (N_6755,N_1301,N_3840);
or U6756 (N_6756,N_876,N_2387);
nor U6757 (N_6757,N_3978,N_1600);
nand U6758 (N_6758,N_3879,N_1075);
nor U6759 (N_6759,N_4172,N_1861);
and U6760 (N_6760,N_2807,N_1153);
nand U6761 (N_6761,N_1835,N_4978);
and U6762 (N_6762,N_1545,N_1243);
nor U6763 (N_6763,N_3537,N_724);
nand U6764 (N_6764,N_3471,N_4044);
nor U6765 (N_6765,N_622,N_3066);
nor U6766 (N_6766,N_1093,N_593);
or U6767 (N_6767,N_1382,N_1361);
nand U6768 (N_6768,N_3764,N_4923);
and U6769 (N_6769,N_133,N_3783);
or U6770 (N_6770,N_138,N_1274);
or U6771 (N_6771,N_4168,N_4397);
and U6772 (N_6772,N_4335,N_4427);
nor U6773 (N_6773,N_2936,N_2823);
xor U6774 (N_6774,N_4399,N_2981);
nand U6775 (N_6775,N_895,N_4494);
and U6776 (N_6776,N_4457,N_4727);
or U6777 (N_6777,N_1991,N_3355);
nor U6778 (N_6778,N_4410,N_4244);
nor U6779 (N_6779,N_3352,N_3654);
nor U6780 (N_6780,N_700,N_485);
nand U6781 (N_6781,N_3166,N_4036);
nor U6782 (N_6782,N_590,N_2507);
nand U6783 (N_6783,N_4305,N_1808);
and U6784 (N_6784,N_4116,N_4217);
nor U6785 (N_6785,N_4451,N_488);
and U6786 (N_6786,N_3541,N_413);
or U6787 (N_6787,N_1046,N_4275);
nor U6788 (N_6788,N_1866,N_4853);
or U6789 (N_6789,N_1290,N_1714);
or U6790 (N_6790,N_2228,N_1483);
or U6791 (N_6791,N_3746,N_1876);
nor U6792 (N_6792,N_1947,N_1560);
or U6793 (N_6793,N_4716,N_2244);
nor U6794 (N_6794,N_166,N_2504);
nand U6795 (N_6795,N_3195,N_4151);
nor U6796 (N_6796,N_3584,N_2486);
nand U6797 (N_6797,N_1458,N_4529);
and U6798 (N_6798,N_898,N_3773);
or U6799 (N_6799,N_203,N_3531);
or U6800 (N_6800,N_50,N_4906);
and U6801 (N_6801,N_17,N_4013);
or U6802 (N_6802,N_1148,N_267);
nor U6803 (N_6803,N_2473,N_2734);
or U6804 (N_6804,N_2315,N_1642);
nand U6805 (N_6805,N_760,N_4748);
or U6806 (N_6806,N_3299,N_3797);
nand U6807 (N_6807,N_3748,N_749);
and U6808 (N_6808,N_647,N_625);
nand U6809 (N_6809,N_54,N_3325);
nor U6810 (N_6810,N_91,N_1553);
xnor U6811 (N_6811,N_1101,N_3326);
nor U6812 (N_6812,N_2696,N_2267);
and U6813 (N_6813,N_793,N_4190);
nand U6814 (N_6814,N_2309,N_4324);
or U6815 (N_6815,N_2572,N_3036);
and U6816 (N_6816,N_3996,N_739);
and U6817 (N_6817,N_3847,N_3582);
or U6818 (N_6818,N_2766,N_3321);
and U6819 (N_6819,N_2853,N_3552);
or U6820 (N_6820,N_556,N_608);
or U6821 (N_6821,N_1404,N_3878);
nor U6822 (N_6822,N_951,N_2733);
nand U6823 (N_6823,N_3279,N_1262);
nor U6824 (N_6824,N_2318,N_3938);
and U6825 (N_6825,N_4148,N_4770);
and U6826 (N_6826,N_4793,N_2092);
and U6827 (N_6827,N_2685,N_3005);
nor U6828 (N_6828,N_2269,N_461);
and U6829 (N_6829,N_4563,N_2594);
nand U6830 (N_6830,N_695,N_2609);
nand U6831 (N_6831,N_3723,N_2649);
or U6832 (N_6832,N_3618,N_125);
nand U6833 (N_6833,N_1369,N_1584);
and U6834 (N_6834,N_4884,N_4602);
nand U6835 (N_6835,N_3858,N_2114);
nor U6836 (N_6836,N_3616,N_3102);
and U6837 (N_6837,N_528,N_4207);
xor U6838 (N_6838,N_1806,N_3484);
or U6839 (N_6839,N_2491,N_3498);
nand U6840 (N_6840,N_1646,N_1371);
or U6841 (N_6841,N_1828,N_690);
nand U6842 (N_6842,N_1982,N_4914);
and U6843 (N_6843,N_1370,N_1109);
and U6844 (N_6844,N_3693,N_1790);
or U6845 (N_6845,N_2522,N_575);
or U6846 (N_6846,N_836,N_252);
and U6847 (N_6847,N_363,N_3487);
or U6848 (N_6848,N_2956,N_4400);
or U6849 (N_6849,N_4999,N_3307);
and U6850 (N_6850,N_1822,N_9);
nand U6851 (N_6851,N_2074,N_540);
or U6852 (N_6852,N_3602,N_3150);
nand U6853 (N_6853,N_52,N_157);
nand U6854 (N_6854,N_1500,N_1377);
or U6855 (N_6855,N_2055,N_4501);
or U6856 (N_6856,N_3587,N_3744);
or U6857 (N_6857,N_869,N_4586);
or U6858 (N_6858,N_3739,N_1999);
and U6859 (N_6859,N_4278,N_1768);
and U6860 (N_6860,N_4058,N_1175);
nand U6861 (N_6861,N_2122,N_3136);
nor U6862 (N_6862,N_4899,N_3382);
xnor U6863 (N_6863,N_2613,N_2897);
and U6864 (N_6864,N_531,N_82);
and U6865 (N_6865,N_3638,N_2790);
nand U6866 (N_6866,N_2528,N_1581);
nand U6867 (N_6867,N_3068,N_983);
or U6868 (N_6868,N_1911,N_2006);
and U6869 (N_6869,N_4011,N_2247);
nor U6870 (N_6870,N_3946,N_4902);
or U6871 (N_6871,N_3991,N_3514);
and U6872 (N_6872,N_4666,N_1756);
nand U6873 (N_6873,N_3522,N_2584);
and U6874 (N_6874,N_1490,N_4771);
and U6875 (N_6875,N_846,N_4704);
or U6876 (N_6876,N_720,N_3903);
or U6877 (N_6877,N_4676,N_4527);
nand U6878 (N_6878,N_4289,N_3529);
nand U6879 (N_6879,N_4646,N_3771);
nor U6880 (N_6880,N_3222,N_1789);
and U6881 (N_6881,N_3488,N_2446);
nor U6882 (N_6882,N_370,N_2887);
nand U6883 (N_6883,N_3924,N_4807);
xnor U6884 (N_6884,N_3877,N_2063);
nor U6885 (N_6885,N_1795,N_4541);
nand U6886 (N_6886,N_3020,N_4612);
nor U6887 (N_6887,N_1272,N_1259);
nand U6888 (N_6888,N_1984,N_1830);
and U6889 (N_6889,N_1978,N_687);
and U6890 (N_6890,N_3590,N_4182);
nand U6891 (N_6891,N_1824,N_3322);
and U6892 (N_6892,N_791,N_2469);
or U6893 (N_6893,N_4394,N_1024);
or U6894 (N_6894,N_299,N_2234);
and U6895 (N_6895,N_4648,N_3642);
or U6896 (N_6896,N_808,N_3383);
or U6897 (N_6897,N_1703,N_1487);
and U6898 (N_6898,N_188,N_4624);
nor U6899 (N_6899,N_4935,N_3725);
or U6900 (N_6900,N_903,N_3108);
or U6901 (N_6901,N_546,N_4386);
nor U6902 (N_6902,N_692,N_651);
nand U6903 (N_6903,N_4445,N_3831);
or U6904 (N_6904,N_3635,N_1450);
or U6905 (N_6905,N_1631,N_1523);
and U6906 (N_6906,N_2209,N_1009);
nor U6907 (N_6907,N_2988,N_2408);
nand U6908 (N_6908,N_1268,N_1187);
or U6909 (N_6909,N_1496,N_4277);
nor U6910 (N_6910,N_3787,N_3595);
or U6911 (N_6911,N_3963,N_2098);
nand U6912 (N_6912,N_1077,N_1829);
nand U6913 (N_6913,N_4139,N_3653);
nor U6914 (N_6914,N_428,N_323);
nor U6915 (N_6915,N_1228,N_2130);
xnor U6916 (N_6916,N_2795,N_3285);
and U6917 (N_6917,N_1938,N_1897);
nand U6918 (N_6918,N_2370,N_1591);
nand U6919 (N_6919,N_615,N_2404);
nor U6920 (N_6920,N_2019,N_2242);
nand U6921 (N_6921,N_4350,N_1962);
and U6922 (N_6922,N_2018,N_282);
nor U6923 (N_6923,N_4697,N_3216);
nor U6924 (N_6924,N_987,N_1675);
or U6925 (N_6925,N_2901,N_4444);
and U6926 (N_6926,N_3989,N_429);
nand U6927 (N_6927,N_3931,N_1852);
or U6928 (N_6928,N_120,N_234);
nand U6929 (N_6929,N_4085,N_3643);
and U6930 (N_6930,N_1865,N_4374);
xnor U6931 (N_6931,N_4496,N_2663);
nand U6932 (N_6932,N_3521,N_4294);
or U6933 (N_6933,N_446,N_719);
and U6934 (N_6934,N_1907,N_379);
xnor U6935 (N_6935,N_3512,N_1072);
and U6936 (N_6936,N_1855,N_3560);
nand U6937 (N_6937,N_2914,N_2811);
nor U6938 (N_6938,N_4544,N_3001);
nand U6939 (N_6939,N_753,N_3316);
nand U6940 (N_6940,N_3785,N_3155);
and U6941 (N_6941,N_3492,N_2437);
and U6942 (N_6942,N_4976,N_4542);
nand U6943 (N_6943,N_1102,N_1905);
nand U6944 (N_6944,N_4754,N_1809);
nand U6945 (N_6945,N_378,N_3193);
nor U6946 (N_6946,N_1779,N_3030);
nor U6947 (N_6947,N_4887,N_3913);
and U6948 (N_6948,N_4489,N_3041);
nand U6949 (N_6949,N_2970,N_3811);
nor U6950 (N_6950,N_858,N_2320);
and U6951 (N_6951,N_2952,N_3925);
and U6952 (N_6952,N_3586,N_4968);
or U6953 (N_6953,N_4068,N_4130);
nand U6954 (N_6954,N_2534,N_587);
and U6955 (N_6955,N_456,N_2540);
or U6956 (N_6956,N_3003,N_4787);
nand U6957 (N_6957,N_1548,N_106);
nand U6958 (N_6958,N_365,N_4891);
and U6959 (N_6959,N_3902,N_2651);
or U6960 (N_6960,N_4947,N_4320);
and U6961 (N_6961,N_4263,N_3363);
and U6962 (N_6962,N_523,N_273);
xor U6963 (N_6963,N_1883,N_1170);
nand U6964 (N_6964,N_2891,N_3365);
nand U6965 (N_6965,N_1418,N_303);
nor U6966 (N_6966,N_3026,N_4475);
and U6967 (N_6967,N_2730,N_1850);
nor U6968 (N_6968,N_927,N_3534);
nor U6969 (N_6969,N_4327,N_3501);
or U6970 (N_6970,N_348,N_1518);
and U6971 (N_6971,N_3803,N_3835);
nor U6972 (N_6972,N_2789,N_1935);
and U6973 (N_6973,N_979,N_597);
and U6974 (N_6974,N_3997,N_3169);
or U6975 (N_6975,N_4051,N_4561);
nand U6976 (N_6976,N_2297,N_4791);
nor U6977 (N_6977,N_2971,N_2900);
nor U6978 (N_6978,N_4195,N_2414);
nor U6979 (N_6979,N_1561,N_3927);
nor U6980 (N_6980,N_4601,N_1366);
nand U6981 (N_6981,N_648,N_3815);
nand U6982 (N_6982,N_3857,N_4810);
nor U6983 (N_6983,N_2338,N_2877);
or U6984 (N_6984,N_1436,N_1205);
xor U6985 (N_6985,N_1297,N_2513);
or U6986 (N_6986,N_4564,N_2157);
or U6987 (N_6987,N_4502,N_339);
nor U6988 (N_6988,N_1163,N_2443);
nor U6989 (N_6989,N_4234,N_4437);
nand U6990 (N_6990,N_4705,N_2650);
and U6991 (N_6991,N_2081,N_4846);
nand U6992 (N_6992,N_3736,N_2954);
nor U6993 (N_6993,N_2293,N_2713);
nand U6994 (N_6994,N_492,N_4856);
nand U6995 (N_6995,N_3990,N_580);
nor U6996 (N_6996,N_823,N_2162);
nand U6997 (N_6997,N_2459,N_124);
or U6998 (N_6998,N_3483,N_2151);
xor U6999 (N_6999,N_2187,N_941);
and U7000 (N_7000,N_137,N_1256);
or U7001 (N_7001,N_4235,N_4377);
or U7002 (N_7002,N_4957,N_4001);
nand U7003 (N_7003,N_3530,N_1225);
and U7004 (N_7004,N_4608,N_3708);
and U7005 (N_7005,N_4883,N_206);
nor U7006 (N_7006,N_2541,N_2805);
nor U7007 (N_7007,N_3392,N_3272);
or U7008 (N_7008,N_1431,N_2280);
or U7009 (N_7009,N_4545,N_1332);
nor U7010 (N_7010,N_589,N_1762);
nor U7011 (N_7011,N_1254,N_4162);
nor U7012 (N_7012,N_2530,N_1514);
nand U7013 (N_7013,N_409,N_539);
nand U7014 (N_7014,N_1373,N_4973);
and U7015 (N_7015,N_1997,N_2539);
nand U7016 (N_7016,N_2772,N_2630);
and U7017 (N_7017,N_4411,N_1045);
or U7018 (N_7018,N_1468,N_4260);
nand U7019 (N_7019,N_4855,N_2743);
nand U7020 (N_7020,N_2129,N_1352);
and U7021 (N_7021,N_1283,N_548);
nor U7022 (N_7022,N_4472,N_272);
or U7023 (N_7023,N_1992,N_1922);
nand U7024 (N_7024,N_1286,N_326);
or U7025 (N_7025,N_3698,N_3674);
and U7026 (N_7026,N_1636,N_4690);
nand U7027 (N_7027,N_4025,N_4746);
and U7028 (N_7028,N_1893,N_1282);
or U7029 (N_7029,N_4414,N_4559);
nor U7030 (N_7030,N_135,N_484);
nor U7031 (N_7031,N_1091,N_2965);
nand U7032 (N_7032,N_716,N_2617);
nand U7033 (N_7033,N_3503,N_2025);
nand U7034 (N_7034,N_4826,N_2120);
or U7035 (N_7035,N_3269,N_1208);
and U7036 (N_7036,N_2925,N_4735);
nand U7037 (N_7037,N_3844,N_3144);
or U7038 (N_7038,N_4848,N_3682);
nor U7039 (N_7039,N_744,N_307);
and U7040 (N_7040,N_872,N_2973);
nand U7041 (N_7041,N_3898,N_2192);
and U7042 (N_7042,N_174,N_3727);
xor U7043 (N_7043,N_3977,N_803);
or U7044 (N_7044,N_816,N_3625);
nor U7045 (N_7045,N_3813,N_4738);
nand U7046 (N_7046,N_2497,N_924);
or U7047 (N_7047,N_4524,N_164);
nand U7048 (N_7048,N_1158,N_4801);
and U7049 (N_7049,N_3715,N_1309);
and U7050 (N_7050,N_1320,N_4583);
and U7051 (N_7051,N_1303,N_999);
and U7052 (N_7052,N_3458,N_3442);
or U7053 (N_7053,N_1774,N_3681);
and U7054 (N_7054,N_3354,N_2577);
nor U7055 (N_7055,N_2729,N_4637);
or U7056 (N_7056,N_198,N_3138);
nor U7057 (N_7057,N_2738,N_4339);
or U7058 (N_7058,N_965,N_1197);
or U7059 (N_7059,N_3728,N_3073);
or U7060 (N_7060,N_4688,N_2705);
nand U7061 (N_7061,N_3493,N_1889);
or U7062 (N_7062,N_4469,N_2358);
or U7063 (N_7063,N_2420,N_3496);
nand U7064 (N_7064,N_1701,N_4396);
nor U7065 (N_7065,N_957,N_4363);
and U7066 (N_7066,N_4817,N_3412);
or U7067 (N_7067,N_4385,N_1993);
or U7068 (N_7068,N_1502,N_4831);
nand U7069 (N_7069,N_1644,N_57);
nand U7070 (N_7070,N_3055,N_2718);
nand U7071 (N_7071,N_3104,N_4654);
and U7072 (N_7072,N_2339,N_1415);
nor U7073 (N_7073,N_2218,N_630);
or U7074 (N_7074,N_3291,N_671);
and U7075 (N_7075,N_3208,N_1162);
and U7076 (N_7076,N_4208,N_1791);
nor U7077 (N_7077,N_3834,N_1010);
nor U7078 (N_7078,N_537,N_4262);
or U7079 (N_7079,N_416,N_2553);
or U7080 (N_7080,N_1459,N_621);
or U7081 (N_7081,N_3795,N_1000);
nor U7082 (N_7082,N_1932,N_455);
or U7083 (N_7083,N_4904,N_4150);
nand U7084 (N_7084,N_3071,N_3175);
nand U7085 (N_7085,N_2983,N_219);
nand U7086 (N_7086,N_197,N_2410);
nand U7087 (N_7087,N_4298,N_1534);
nor U7088 (N_7088,N_2543,N_2723);
nand U7089 (N_7089,N_3707,N_2472);
and U7090 (N_7090,N_1563,N_3226);
and U7091 (N_7091,N_1341,N_43);
nor U7092 (N_7092,N_149,N_4443);
nor U7093 (N_7093,N_3140,N_3477);
or U7094 (N_7094,N_3880,N_3284);
nand U7095 (N_7095,N_3470,N_3801);
nor U7096 (N_7096,N_4045,N_77);
or U7097 (N_7097,N_420,N_3188);
and U7098 (N_7098,N_26,N_4587);
nor U7099 (N_7099,N_1047,N_3277);
nor U7100 (N_7100,N_2894,N_4723);
nand U7101 (N_7101,N_1410,N_4106);
nor U7102 (N_7102,N_3137,N_1798);
nor U7103 (N_7103,N_1799,N_4194);
and U7104 (N_7104,N_1296,N_2941);
nand U7105 (N_7105,N_44,N_4434);
and U7106 (N_7106,N_1498,N_4515);
nand U7107 (N_7107,N_3519,N_1647);
or U7108 (N_7108,N_1494,N_3157);
nand U7109 (N_7109,N_4346,N_4852);
xnor U7110 (N_7110,N_3368,N_1057);
or U7111 (N_7111,N_4517,N_2262);
and U7112 (N_7112,N_977,N_3884);
nor U7113 (N_7113,N_3398,N_2825);
nor U7114 (N_7114,N_1190,N_904);
nor U7115 (N_7115,N_2390,N_4384);
or U7116 (N_7116,N_4910,N_4216);
nor U7117 (N_7117,N_3294,N_4306);
nor U7118 (N_7118,N_4105,N_2499);
or U7119 (N_7119,N_1981,N_310);
nor U7120 (N_7120,N_88,N_3690);
and U7121 (N_7121,N_992,N_3546);
or U7122 (N_7122,N_1786,N_3508);
nand U7123 (N_7123,N_2545,N_3955);
or U7124 (N_7124,N_1552,N_4577);
and U7125 (N_7125,N_746,N_1455);
or U7126 (N_7126,N_602,N_3273);
and U7127 (N_7127,N_4830,N_3882);
or U7128 (N_7128,N_3067,N_1669);
and U7129 (N_7129,N_1781,N_4449);
or U7130 (N_7130,N_552,N_4597);
nor U7131 (N_7131,N_4713,N_4604);
or U7132 (N_7132,N_1348,N_3621);
nor U7133 (N_7133,N_1220,N_1397);
and U7134 (N_7134,N_5,N_401);
and U7135 (N_7135,N_1515,N_3495);
and U7136 (N_7136,N_1976,N_2860);
and U7137 (N_7137,N_1934,N_3599);
and U7138 (N_7138,N_2962,N_180);
or U7139 (N_7139,N_4598,N_2357);
or U7140 (N_7140,N_3830,N_3612);
nor U7141 (N_7141,N_4154,N_34);
nand U7142 (N_7142,N_3816,N_1580);
nor U7143 (N_7143,N_3312,N_3414);
nand U7144 (N_7144,N_1896,N_4117);
and U7145 (N_7145,N_661,N_3344);
and U7146 (N_7146,N_4265,N_1744);
or U7147 (N_7147,N_2316,N_3165);
or U7148 (N_7148,N_4135,N_4647);
or U7149 (N_7149,N_296,N_4251);
and U7150 (N_7150,N_4299,N_4176);
nand U7151 (N_7151,N_475,N_3872);
nor U7152 (N_7152,N_3025,N_2109);
or U7153 (N_7153,N_1780,N_1979);
nor U7154 (N_7154,N_447,N_652);
nor U7155 (N_7155,N_1805,N_2077);
nand U7156 (N_7156,N_917,N_3004);
nor U7157 (N_7157,N_83,N_4653);
nand U7158 (N_7158,N_4795,N_3019);
nand U7159 (N_7159,N_2579,N_4847);
or U7160 (N_7160,N_511,N_3611);
nor U7161 (N_7161,N_1474,N_3918);
nor U7162 (N_7162,N_2203,N_806);
nand U7163 (N_7163,N_3457,N_319);
nand U7164 (N_7164,N_4000,N_3689);
nor U7165 (N_7165,N_2438,N_4591);
nand U7166 (N_7166,N_2254,N_1551);
nor U7167 (N_7167,N_4024,N_3581);
and U7168 (N_7168,N_4623,N_654);
nor U7169 (N_7169,N_3083,N_98);
nand U7170 (N_7170,N_4259,N_236);
and U7171 (N_7171,N_1787,N_4872);
nand U7172 (N_7172,N_4557,N_3109);
nor U7173 (N_7173,N_2682,N_3677);
or U7174 (N_7174,N_3049,N_609);
nand U7175 (N_7175,N_1698,N_3007);
nand U7176 (N_7176,N_559,N_3555);
and U7177 (N_7177,N_2917,N_2765);
nand U7178 (N_7178,N_3349,N_2782);
nand U7179 (N_7179,N_1802,N_2413);
nor U7180 (N_7180,N_4479,N_259);
or U7181 (N_7181,N_954,N_4236);
nor U7182 (N_7182,N_2134,N_4046);
nor U7183 (N_7183,N_4941,N_4158);
nor U7184 (N_7184,N_2116,N_990);
and U7185 (N_7185,N_2802,N_4912);
nand U7186 (N_7186,N_1138,N_3678);
and U7187 (N_7187,N_4313,N_1930);
and U7188 (N_7188,N_792,N_86);
or U7189 (N_7189,N_2756,N_897);
or U7190 (N_7190,N_3242,N_4772);
and U7191 (N_7191,N_4120,N_2959);
or U7192 (N_7192,N_3302,N_2888);
and U7193 (N_7193,N_2865,N_4530);
or U7194 (N_7194,N_337,N_1402);
xnor U7195 (N_7195,N_2529,N_4576);
and U7196 (N_7196,N_4056,N_3542);
xnor U7197 (N_7197,N_4006,N_494);
and U7198 (N_7198,N_3131,N_1086);
or U7199 (N_7199,N_763,N_4160);
or U7200 (N_7200,N_1157,N_4995);
nand U7201 (N_7201,N_3163,N_2377);
or U7202 (N_7202,N_3063,N_4079);
or U7203 (N_7203,N_908,N_4426);
xor U7204 (N_7204,N_800,N_644);
and U7205 (N_7205,N_811,N_1151);
or U7206 (N_7206,N_1846,N_1065);
nand U7207 (N_7207,N_2951,N_4533);
nor U7208 (N_7208,N_1200,N_1598);
or U7209 (N_7209,N_2433,N_3826);
or U7210 (N_7210,N_3429,N_612);
or U7211 (N_7211,N_4227,N_4939);
xnor U7212 (N_7212,N_2967,N_3829);
and U7213 (N_7213,N_1452,N_2065);
nand U7214 (N_7214,N_244,N_901);
nor U7215 (N_7215,N_1020,N_529);
and U7216 (N_7216,N_2926,N_2219);
or U7217 (N_7217,N_4014,N_2035);
nand U7218 (N_7218,N_1068,N_4042);
or U7219 (N_7219,N_3869,N_84);
or U7220 (N_7220,N_754,N_1030);
and U7221 (N_7221,N_3548,N_536);
and U7222 (N_7222,N_1596,N_4739);
nor U7223 (N_7223,N_1261,N_241);
nor U7224 (N_7224,N_2985,N_2662);
or U7225 (N_7225,N_4672,N_4695);
or U7226 (N_7226,N_1980,N_1226);
xor U7227 (N_7227,N_663,N_3935);
nand U7228 (N_7228,N_4633,N_3300);
nand U7229 (N_7229,N_1608,N_860);
nor U7230 (N_7230,N_1948,N_2752);
nand U7231 (N_7231,N_3237,N_3199);
nor U7232 (N_7232,N_2974,N_4797);
or U7233 (N_7233,N_3667,N_3904);
or U7234 (N_7234,N_4954,N_4442);
nand U7235 (N_7235,N_3561,N_2232);
and U7236 (N_7236,N_2598,N_2453);
and U7237 (N_7237,N_520,N_156);
or U7238 (N_7238,N_2197,N_3022);
or U7239 (N_7239,N_32,N_822);
nor U7240 (N_7240,N_1407,N_2822);
nor U7241 (N_7241,N_1266,N_2418);
and U7242 (N_7242,N_4803,N_3841);
or U7243 (N_7243,N_829,N_682);
and U7244 (N_7244,N_3865,N_2456);
or U7245 (N_7245,N_1018,N_2697);
nor U7246 (N_7246,N_2371,N_969);
and U7247 (N_7247,N_3792,N_2449);
nor U7248 (N_7248,N_3399,N_997);
nand U7249 (N_7249,N_1539,N_4938);
nor U7250 (N_7250,N_2050,N_3970);
nor U7251 (N_7251,N_726,N_1022);
nor U7252 (N_7252,N_1475,N_327);
nand U7253 (N_7253,N_2972,N_1419);
and U7254 (N_7254,N_4082,N_4188);
and U7255 (N_7255,N_1977,N_2056);
nand U7256 (N_7256,N_1104,N_254);
or U7257 (N_7257,N_3766,N_4061);
or U7258 (N_7258,N_3040,N_1315);
nand U7259 (N_7259,N_454,N_3676);
and U7260 (N_7260,N_554,N_3711);
or U7261 (N_7261,N_1814,N_694);
xor U7262 (N_7262,N_3000,N_3308);
nand U7263 (N_7263,N_1173,N_4375);
nor U7264 (N_7264,N_2016,N_4441);
or U7265 (N_7265,N_1892,N_2571);
nor U7266 (N_7266,N_1804,N_1574);
nor U7267 (N_7267,N_2223,N_2763);
xor U7268 (N_7268,N_4110,N_3668);
or U7269 (N_7269,N_3252,N_4761);
xnor U7270 (N_7270,N_1748,N_4094);
xor U7271 (N_7271,N_2105,N_2995);
nor U7272 (N_7272,N_3180,N_1390);
nor U7273 (N_7273,N_345,N_4332);
and U7274 (N_7274,N_713,N_820);
or U7275 (N_7275,N_2709,N_827);
or U7276 (N_7276,N_1875,N_304);
or U7277 (N_7277,N_215,N_2027);
nor U7278 (N_7278,N_2170,N_3874);
or U7279 (N_7279,N_1307,N_3523);
nor U7280 (N_7280,N_1785,N_2544);
nor U7281 (N_7281,N_1933,N_487);
nand U7282 (N_7282,N_1437,N_2773);
nand U7283 (N_7283,N_3288,N_1823);
or U7284 (N_7284,N_4665,N_3339);
or U7285 (N_7285,N_1150,N_403);
and U7286 (N_7286,N_3613,N_1692);
nor U7287 (N_7287,N_502,N_366);
and U7288 (N_7288,N_357,N_1067);
or U7289 (N_7289,N_71,N_848);
or U7290 (N_7290,N_3566,N_208);
nor U7291 (N_7291,N_129,N_2126);
nand U7292 (N_7292,N_4929,N_1746);
nor U7293 (N_7293,N_2142,N_4027);
nor U7294 (N_7294,N_2994,N_1681);
and U7295 (N_7295,N_4484,N_3610);
nor U7296 (N_7296,N_4970,N_4352);
nand U7297 (N_7297,N_1218,N_4547);
xnor U7298 (N_7298,N_4477,N_1803);
nand U7299 (N_7299,N_3951,N_4038);
nand U7300 (N_7300,N_2195,N_4782);
nor U7301 (N_7301,N_300,N_2102);
and U7302 (N_7302,N_4821,N_3364);
and U7303 (N_7303,N_861,N_4805);
nor U7304 (N_7304,N_3204,N_1648);
nand U7305 (N_7305,N_2355,N_1690);
xnor U7306 (N_7306,N_2638,N_3499);
nand U7307 (N_7307,N_2874,N_1323);
and U7308 (N_7308,N_4949,N_4991);
and U7309 (N_7309,N_42,N_3583);
nand U7310 (N_7310,N_3513,N_24);
nand U7311 (N_7311,N_4534,N_2524);
or U7312 (N_7312,N_4240,N_1409);
nor U7313 (N_7313,N_1106,N_585);
nand U7314 (N_7314,N_1184,N_975);
or U7315 (N_7315,N_3045,N_4636);
nand U7316 (N_7316,N_4988,N_4549);
and U7317 (N_7317,N_1015,N_4865);
nor U7318 (N_7318,N_2230,N_1232);
nand U7319 (N_7319,N_2276,N_3930);
nand U7320 (N_7320,N_4977,N_1571);
nor U7321 (N_7321,N_3401,N_3687);
nand U7322 (N_7322,N_2707,N_1328);
nor U7323 (N_7323,N_1330,N_3210);
nand U7324 (N_7324,N_577,N_248);
nand U7325 (N_7325,N_2570,N_1333);
nand U7326 (N_7326,N_4268,N_4403);
and U7327 (N_7327,N_809,N_3048);
and U7328 (N_7328,N_1147,N_2757);
nor U7329 (N_7329,N_1460,N_1031);
and U7330 (N_7330,N_2684,N_3435);
nor U7331 (N_7331,N_126,N_207);
and U7332 (N_7332,N_1247,N_3605);
nand U7333 (N_7333,N_61,N_657);
and U7334 (N_7334,N_4063,N_675);
and U7335 (N_7335,N_2401,N_3306);
and U7336 (N_7336,N_4590,N_2221);
nand U7337 (N_7337,N_1901,N_3754);
and U7338 (N_7338,N_2400,N_1585);
nor U7339 (N_7339,N_1177,N_934);
nand U7340 (N_7340,N_3720,N_1733);
or U7341 (N_7341,N_2641,N_2349);
and U7342 (N_7342,N_842,N_3862);
and U7343 (N_7343,N_1270,N_67);
nand U7344 (N_7344,N_1909,N_4974);
or U7345 (N_7345,N_4655,N_1540);
nand U7346 (N_7346,N_1444,N_4112);
or U7347 (N_7347,N_595,N_2512);
or U7348 (N_7348,N_4878,N_2070);
and U7349 (N_7349,N_1488,N_2892);
nor U7350 (N_7350,N_311,N_142);
or U7351 (N_7351,N_696,N_3733);
or U7352 (N_7352,N_3329,N_3601);
and U7353 (N_7353,N_629,N_4631);
nand U7354 (N_7354,N_1945,N_3672);
or U7355 (N_7355,N_830,N_3033);
and U7356 (N_7356,N_1064,N_4423);
nor U7357 (N_7357,N_431,N_4435);
nand U7358 (N_7358,N_3671,N_3825);
nand U7359 (N_7359,N_2870,N_1378);
nor U7360 (N_7360,N_3737,N_94);
nand U7361 (N_7361,N_2298,N_3607);
nand U7362 (N_7362,N_4990,N_689);
xnor U7363 (N_7363,N_31,N_4088);
nand U7364 (N_7364,N_2191,N_3214);
nand U7365 (N_7365,N_1439,N_1192);
and U7366 (N_7366,N_1449,N_4897);
nor U7367 (N_7367,N_439,N_473);
or U7368 (N_7368,N_4963,N_3186);
nand U7369 (N_7369,N_286,N_3125);
nand U7370 (N_7370,N_3168,N_3332);
and U7371 (N_7371,N_223,N_4353);
nand U7372 (N_7372,N_3127,N_2484);
or U7373 (N_7373,N_4784,N_880);
or U7374 (N_7374,N_1727,N_1442);
and U7375 (N_7375,N_4065,N_631);
or U7376 (N_7376,N_1821,N_4861);
nand U7377 (N_7377,N_176,N_4755);
nor U7378 (N_7378,N_1304,N_1655);
nor U7379 (N_7379,N_2249,N_3824);
or U7380 (N_7380,N_2046,N_859);
nand U7381 (N_7381,N_4203,N_4816);
or U7382 (N_7382,N_3391,N_4239);
or U7383 (N_7383,N_1376,N_844);
nand U7384 (N_7384,N_1782,N_2902);
or U7385 (N_7385,N_1715,N_2248);
nor U7386 (N_7386,N_1011,N_3367);
or U7387 (N_7387,N_1362,N_3225);
or U7388 (N_7388,N_2289,N_614);
and U7389 (N_7389,N_1921,N_218);
and U7390 (N_7390,N_4700,N_1547);
nand U7391 (N_7391,N_1070,N_3864);
nor U7392 (N_7392,N_2351,N_4136);
xnor U7393 (N_7393,N_505,N_2852);
and U7394 (N_7394,N_3703,N_2372);
nand U7395 (N_7395,N_2169,N_3651);
nor U7396 (N_7396,N_3212,N_246);
nor U7397 (N_7397,N_1154,N_41);
and U7398 (N_7398,N_4786,N_542);
and U7399 (N_7399,N_4877,N_4241);
nand U7400 (N_7400,N_2033,N_3981);
and U7401 (N_7401,N_2964,N_1542);
nor U7402 (N_7402,N_2434,N_1557);
nand U7403 (N_7403,N_4975,N_221);
nand U7404 (N_7404,N_2012,N_2222);
and U7405 (N_7405,N_2523,N_497);
nand U7406 (N_7406,N_4323,N_0);
nor U7407 (N_7407,N_558,N_781);
nor U7408 (N_7408,N_2005,N_4311);
nand U7409 (N_7409,N_1754,N_3572);
nand U7410 (N_7410,N_3603,N_1079);
or U7411 (N_7411,N_4726,N_4768);
nor U7412 (N_7412,N_1857,N_1920);
and U7413 (N_7413,N_578,N_2430);
nor U7414 (N_7414,N_4246,N_1464);
and U7415 (N_7415,N_4798,N_4948);
or U7416 (N_7416,N_1379,N_1549);
and U7417 (N_7417,N_3683,N_177);
or U7418 (N_7418,N_3319,N_4460);
nand U7419 (N_7419,N_2574,N_2141);
and U7420 (N_7420,N_2503,N_4680);
and U7421 (N_7421,N_4464,N_1877);
nand U7422 (N_7422,N_2864,N_4859);
nor U7423 (N_7423,N_4692,N_2185);
nor U7424 (N_7424,N_4287,N_3886);
or U7425 (N_7425,N_3478,N_358);
and U7426 (N_7426,N_912,N_2886);
or U7427 (N_7427,N_4347,N_4620);
or U7428 (N_7428,N_4144,N_3230);
nor U7429 (N_7429,N_364,N_2001);
nand U7430 (N_7430,N_1609,N_2910);
or U7431 (N_7431,N_2969,N_4509);
or U7432 (N_7432,N_1505,N_4010);
or U7433 (N_7433,N_4205,N_4303);
or U7434 (N_7434,N_813,N_2578);
nand U7435 (N_7435,N_4600,N_3808);
nand U7436 (N_7436,N_4325,N_2509);
nor U7437 (N_7437,N_328,N_4903);
nor U7438 (N_7438,N_870,N_1705);
or U7439 (N_7439,N_968,N_2461);
or U7440 (N_7440,N_674,N_1253);
nand U7441 (N_7441,N_4439,N_3286);
and U7442 (N_7442,N_445,N_2839);
nand U7443 (N_7443,N_1146,N_2879);
nand U7444 (N_7444,N_1117,N_3986);
or U7445 (N_7445,N_994,N_495);
or U7446 (N_7446,N_293,N_4982);
nor U7447 (N_7447,N_4521,N_4169);
xnor U7448 (N_7448,N_226,N_1063);
nand U7449 (N_7449,N_3327,N_4064);
and U7450 (N_7450,N_4255,N_4295);
xor U7451 (N_7451,N_3949,N_4773);
or U7452 (N_7452,N_3227,N_2466);
or U7453 (N_7453,N_1667,N_4525);
and U7454 (N_7454,N_87,N_3159);
nor U7455 (N_7455,N_170,N_2462);
nor U7456 (N_7456,N_66,N_3696);
and U7457 (N_7457,N_4536,N_2691);
xor U7458 (N_7458,N_2082,N_4619);
nor U7459 (N_7459,N_4628,N_4686);
or U7460 (N_7460,N_4913,N_4701);
nor U7461 (N_7461,N_19,N_308);
and U7462 (N_7462,N_1685,N_2145);
and U7463 (N_7463,N_1143,N_3178);
and U7464 (N_7464,N_4868,N_1848);
nand U7465 (N_7465,N_4785,N_3998);
and U7466 (N_7466,N_3384,N_3536);
nor U7467 (N_7467,N_2135,N_3425);
and U7468 (N_7468,N_3249,N_1995);
nand U7469 (N_7469,N_258,N_4513);
nor U7470 (N_7470,N_1171,N_3794);
nand U7471 (N_7471,N_1100,N_2252);
nor U7472 (N_7472,N_1739,N_933);
and U7473 (N_7473,N_3992,N_3968);
nand U7474 (N_7474,N_4142,N_1335);
nand U7475 (N_7475,N_3077,N_3122);
and U7476 (N_7476,N_190,N_3024);
nor U7477 (N_7477,N_1693,N_3619);
or U7478 (N_7478,N_144,N_4825);
and U7479 (N_7479,N_1594,N_3598);
and U7480 (N_7480,N_2986,N_930);
nor U7481 (N_7481,N_2064,N_3280);
xor U7482 (N_7482,N_707,N_3524);
nand U7483 (N_7483,N_426,N_4593);
or U7484 (N_7484,N_801,N_2841);
or U7485 (N_7485,N_458,N_3885);
nor U7486 (N_7486,N_573,N_4749);
and U7487 (N_7487,N_4538,N_1788);
or U7488 (N_7488,N_1062,N_3558);
nand U7489 (N_7489,N_2494,N_1033);
and U7490 (N_7490,N_4714,N_419);
nor U7491 (N_7491,N_1844,N_2827);
nand U7492 (N_7492,N_2399,N_1351);
nor U7493 (N_7493,N_4986,N_3031);
or U7494 (N_7494,N_553,N_3101);
nor U7495 (N_7495,N_970,N_4744);
nand U7496 (N_7496,N_2306,N_3060);
and U7497 (N_7497,N_4792,N_881);
and U7498 (N_7498,N_1737,N_1246);
and U7499 (N_7499,N_4357,N_4143);
nor U7500 (N_7500,N_1844,N_541);
and U7501 (N_7501,N_2400,N_3026);
xor U7502 (N_7502,N_2272,N_3798);
nor U7503 (N_7503,N_2783,N_1611);
nand U7504 (N_7504,N_1084,N_2742);
nor U7505 (N_7505,N_373,N_16);
nand U7506 (N_7506,N_3713,N_2877);
and U7507 (N_7507,N_4300,N_2516);
nor U7508 (N_7508,N_4516,N_2477);
or U7509 (N_7509,N_704,N_1845);
xor U7510 (N_7510,N_920,N_3449);
or U7511 (N_7511,N_3340,N_4700);
nand U7512 (N_7512,N_1092,N_4423);
nor U7513 (N_7513,N_780,N_233);
and U7514 (N_7514,N_2472,N_4524);
nor U7515 (N_7515,N_4270,N_2590);
and U7516 (N_7516,N_252,N_2131);
or U7517 (N_7517,N_731,N_4760);
or U7518 (N_7518,N_3226,N_2574);
or U7519 (N_7519,N_191,N_2834);
nor U7520 (N_7520,N_630,N_3748);
nand U7521 (N_7521,N_1017,N_3306);
nand U7522 (N_7522,N_1629,N_14);
nand U7523 (N_7523,N_2564,N_3520);
and U7524 (N_7524,N_1472,N_3840);
nor U7525 (N_7525,N_3425,N_3964);
or U7526 (N_7526,N_164,N_2752);
and U7527 (N_7527,N_853,N_4601);
nor U7528 (N_7528,N_3611,N_2078);
and U7529 (N_7529,N_4250,N_3444);
or U7530 (N_7530,N_3287,N_1727);
nand U7531 (N_7531,N_3665,N_3688);
nor U7532 (N_7532,N_477,N_1407);
nand U7533 (N_7533,N_1487,N_2151);
and U7534 (N_7534,N_1721,N_2116);
nand U7535 (N_7535,N_430,N_2513);
and U7536 (N_7536,N_1759,N_260);
nor U7537 (N_7537,N_2196,N_1211);
xnor U7538 (N_7538,N_4777,N_3194);
and U7539 (N_7539,N_2947,N_2225);
xnor U7540 (N_7540,N_4624,N_296);
nand U7541 (N_7541,N_735,N_1638);
and U7542 (N_7542,N_4150,N_2289);
nand U7543 (N_7543,N_2794,N_735);
and U7544 (N_7544,N_3106,N_3596);
nand U7545 (N_7545,N_4017,N_2198);
nor U7546 (N_7546,N_988,N_796);
or U7547 (N_7547,N_3611,N_1046);
nor U7548 (N_7548,N_1179,N_429);
or U7549 (N_7549,N_2731,N_499);
and U7550 (N_7550,N_4661,N_1611);
nor U7551 (N_7551,N_337,N_1820);
or U7552 (N_7552,N_1970,N_2162);
or U7553 (N_7553,N_1862,N_2284);
nor U7554 (N_7554,N_1355,N_4564);
and U7555 (N_7555,N_3925,N_2703);
nand U7556 (N_7556,N_3724,N_668);
nand U7557 (N_7557,N_1418,N_2021);
nor U7558 (N_7558,N_3959,N_3026);
or U7559 (N_7559,N_3031,N_1311);
nand U7560 (N_7560,N_444,N_2988);
xnor U7561 (N_7561,N_1160,N_523);
or U7562 (N_7562,N_2735,N_506);
nor U7563 (N_7563,N_1164,N_2567);
or U7564 (N_7564,N_4729,N_4723);
nor U7565 (N_7565,N_2226,N_2724);
and U7566 (N_7566,N_1856,N_964);
nor U7567 (N_7567,N_1037,N_1922);
or U7568 (N_7568,N_1184,N_2002);
nand U7569 (N_7569,N_2928,N_233);
and U7570 (N_7570,N_1564,N_3354);
nor U7571 (N_7571,N_4209,N_4843);
and U7572 (N_7572,N_2605,N_1339);
or U7573 (N_7573,N_344,N_2108);
nand U7574 (N_7574,N_2601,N_3096);
nor U7575 (N_7575,N_4560,N_2806);
or U7576 (N_7576,N_1309,N_3375);
nor U7577 (N_7577,N_357,N_2873);
and U7578 (N_7578,N_661,N_3260);
nor U7579 (N_7579,N_3378,N_1539);
and U7580 (N_7580,N_2085,N_1462);
or U7581 (N_7581,N_3833,N_4554);
or U7582 (N_7582,N_253,N_2426);
and U7583 (N_7583,N_2556,N_2044);
and U7584 (N_7584,N_4216,N_2724);
xor U7585 (N_7585,N_621,N_3521);
nand U7586 (N_7586,N_4484,N_2980);
or U7587 (N_7587,N_3245,N_2080);
nand U7588 (N_7588,N_732,N_3228);
nor U7589 (N_7589,N_3323,N_1411);
or U7590 (N_7590,N_795,N_4006);
and U7591 (N_7591,N_178,N_882);
or U7592 (N_7592,N_4380,N_3845);
nor U7593 (N_7593,N_1803,N_660);
xnor U7594 (N_7594,N_4653,N_1788);
nor U7595 (N_7595,N_669,N_1905);
nand U7596 (N_7596,N_1971,N_141);
nor U7597 (N_7597,N_4101,N_1477);
nor U7598 (N_7598,N_3398,N_4124);
nand U7599 (N_7599,N_830,N_2497);
and U7600 (N_7600,N_3608,N_1132);
and U7601 (N_7601,N_2465,N_1512);
nand U7602 (N_7602,N_1138,N_2377);
or U7603 (N_7603,N_3959,N_2641);
or U7604 (N_7604,N_2030,N_4124);
nand U7605 (N_7605,N_3292,N_1325);
and U7606 (N_7606,N_1457,N_4734);
or U7607 (N_7607,N_4133,N_3243);
nor U7608 (N_7608,N_200,N_139);
and U7609 (N_7609,N_2591,N_3534);
and U7610 (N_7610,N_3989,N_3195);
xor U7611 (N_7611,N_3526,N_2087);
and U7612 (N_7612,N_2459,N_2411);
or U7613 (N_7613,N_2130,N_4562);
or U7614 (N_7614,N_2043,N_1767);
or U7615 (N_7615,N_3001,N_1583);
nand U7616 (N_7616,N_390,N_1294);
nor U7617 (N_7617,N_3534,N_2706);
nor U7618 (N_7618,N_2316,N_2435);
or U7619 (N_7619,N_2777,N_1240);
and U7620 (N_7620,N_4927,N_2573);
nand U7621 (N_7621,N_4951,N_2254);
nand U7622 (N_7622,N_3514,N_765);
nor U7623 (N_7623,N_4862,N_4757);
xnor U7624 (N_7624,N_128,N_1604);
and U7625 (N_7625,N_4378,N_2856);
nand U7626 (N_7626,N_3582,N_3778);
nor U7627 (N_7627,N_1728,N_3215);
nand U7628 (N_7628,N_1800,N_3235);
nand U7629 (N_7629,N_2377,N_1303);
and U7630 (N_7630,N_2899,N_3249);
xor U7631 (N_7631,N_2844,N_4001);
and U7632 (N_7632,N_2069,N_2649);
nand U7633 (N_7633,N_4554,N_1291);
and U7634 (N_7634,N_2660,N_3340);
nand U7635 (N_7635,N_4190,N_4496);
and U7636 (N_7636,N_3956,N_4661);
nand U7637 (N_7637,N_220,N_3119);
nand U7638 (N_7638,N_1116,N_4322);
xor U7639 (N_7639,N_812,N_2548);
and U7640 (N_7640,N_3083,N_1534);
or U7641 (N_7641,N_610,N_1183);
nand U7642 (N_7642,N_1806,N_4311);
nor U7643 (N_7643,N_606,N_4680);
and U7644 (N_7644,N_3064,N_4233);
nand U7645 (N_7645,N_925,N_4922);
nand U7646 (N_7646,N_149,N_129);
xnor U7647 (N_7647,N_70,N_985);
nor U7648 (N_7648,N_3912,N_4186);
and U7649 (N_7649,N_3133,N_4018);
or U7650 (N_7650,N_4457,N_853);
or U7651 (N_7651,N_2839,N_4894);
and U7652 (N_7652,N_153,N_130);
nor U7653 (N_7653,N_1459,N_2775);
nor U7654 (N_7654,N_1725,N_402);
nand U7655 (N_7655,N_57,N_2664);
and U7656 (N_7656,N_1031,N_4234);
nand U7657 (N_7657,N_4148,N_3404);
nand U7658 (N_7658,N_2713,N_3204);
nor U7659 (N_7659,N_3905,N_3535);
or U7660 (N_7660,N_3919,N_3758);
nand U7661 (N_7661,N_3958,N_921);
nand U7662 (N_7662,N_1009,N_2390);
nand U7663 (N_7663,N_2989,N_3950);
or U7664 (N_7664,N_2914,N_1061);
nor U7665 (N_7665,N_2042,N_4050);
nor U7666 (N_7666,N_2247,N_633);
nor U7667 (N_7667,N_2259,N_1174);
or U7668 (N_7668,N_865,N_396);
nor U7669 (N_7669,N_399,N_3117);
nor U7670 (N_7670,N_4922,N_414);
nand U7671 (N_7671,N_3498,N_597);
nand U7672 (N_7672,N_1645,N_2163);
or U7673 (N_7673,N_4265,N_4714);
or U7674 (N_7674,N_958,N_335);
or U7675 (N_7675,N_798,N_4836);
or U7676 (N_7676,N_1369,N_4629);
nand U7677 (N_7677,N_776,N_2569);
and U7678 (N_7678,N_2653,N_4871);
nand U7679 (N_7679,N_4232,N_3504);
nand U7680 (N_7680,N_2154,N_3309);
nand U7681 (N_7681,N_1025,N_4731);
nor U7682 (N_7682,N_1403,N_1394);
xor U7683 (N_7683,N_4237,N_1323);
nand U7684 (N_7684,N_2975,N_2760);
or U7685 (N_7685,N_2803,N_4969);
or U7686 (N_7686,N_1323,N_1082);
or U7687 (N_7687,N_1948,N_4332);
or U7688 (N_7688,N_4968,N_1835);
or U7689 (N_7689,N_1931,N_816);
or U7690 (N_7690,N_3212,N_1223);
nand U7691 (N_7691,N_4533,N_4119);
or U7692 (N_7692,N_1532,N_4262);
nand U7693 (N_7693,N_2511,N_3233);
or U7694 (N_7694,N_3753,N_4566);
nand U7695 (N_7695,N_618,N_4491);
nor U7696 (N_7696,N_1885,N_68);
nand U7697 (N_7697,N_790,N_2647);
and U7698 (N_7698,N_3545,N_2581);
nand U7699 (N_7699,N_2063,N_1008);
nor U7700 (N_7700,N_4637,N_3749);
nand U7701 (N_7701,N_4897,N_1228);
nor U7702 (N_7702,N_2513,N_3306);
or U7703 (N_7703,N_992,N_1109);
and U7704 (N_7704,N_3861,N_4803);
and U7705 (N_7705,N_2335,N_104);
or U7706 (N_7706,N_2381,N_1186);
and U7707 (N_7707,N_3101,N_3117);
or U7708 (N_7708,N_3830,N_676);
and U7709 (N_7709,N_914,N_3485);
nor U7710 (N_7710,N_3596,N_2241);
nor U7711 (N_7711,N_4332,N_832);
and U7712 (N_7712,N_1781,N_767);
nand U7713 (N_7713,N_2864,N_556);
and U7714 (N_7714,N_1566,N_2687);
nor U7715 (N_7715,N_4233,N_360);
nand U7716 (N_7716,N_3212,N_1170);
and U7717 (N_7717,N_3508,N_2285);
or U7718 (N_7718,N_514,N_1249);
or U7719 (N_7719,N_4916,N_2651);
nand U7720 (N_7720,N_863,N_4847);
and U7721 (N_7721,N_361,N_2858);
nand U7722 (N_7722,N_821,N_1846);
nand U7723 (N_7723,N_4414,N_1032);
or U7724 (N_7724,N_2290,N_2766);
nand U7725 (N_7725,N_1996,N_698);
nor U7726 (N_7726,N_4808,N_2642);
nor U7727 (N_7727,N_2418,N_2164);
or U7728 (N_7728,N_3671,N_4995);
nor U7729 (N_7729,N_2672,N_2054);
and U7730 (N_7730,N_3112,N_3782);
and U7731 (N_7731,N_2308,N_4787);
and U7732 (N_7732,N_4994,N_1056);
or U7733 (N_7733,N_4904,N_2935);
nor U7734 (N_7734,N_4363,N_871);
and U7735 (N_7735,N_3797,N_1705);
nor U7736 (N_7736,N_2897,N_1728);
or U7737 (N_7737,N_4769,N_3342);
and U7738 (N_7738,N_3013,N_2481);
nand U7739 (N_7739,N_4616,N_1351);
nor U7740 (N_7740,N_172,N_3984);
and U7741 (N_7741,N_1246,N_249);
or U7742 (N_7742,N_2540,N_3025);
nand U7743 (N_7743,N_2008,N_4859);
or U7744 (N_7744,N_3728,N_578);
or U7745 (N_7745,N_4837,N_4281);
nor U7746 (N_7746,N_1457,N_1425);
nor U7747 (N_7747,N_170,N_2364);
nand U7748 (N_7748,N_3244,N_4224);
or U7749 (N_7749,N_1752,N_661);
nor U7750 (N_7750,N_1360,N_3963);
nand U7751 (N_7751,N_3819,N_1805);
nor U7752 (N_7752,N_3049,N_4937);
nand U7753 (N_7753,N_4998,N_3139);
and U7754 (N_7754,N_22,N_2006);
or U7755 (N_7755,N_379,N_2568);
and U7756 (N_7756,N_3096,N_1012);
nor U7757 (N_7757,N_969,N_4255);
or U7758 (N_7758,N_3045,N_3338);
nor U7759 (N_7759,N_283,N_1614);
or U7760 (N_7760,N_4290,N_2118);
nor U7761 (N_7761,N_941,N_1607);
nor U7762 (N_7762,N_963,N_984);
nand U7763 (N_7763,N_1964,N_639);
nor U7764 (N_7764,N_919,N_4379);
or U7765 (N_7765,N_2761,N_3583);
or U7766 (N_7766,N_3049,N_2086);
or U7767 (N_7767,N_3524,N_2535);
nor U7768 (N_7768,N_4725,N_793);
nand U7769 (N_7769,N_1176,N_2675);
and U7770 (N_7770,N_1904,N_1114);
and U7771 (N_7771,N_1167,N_4263);
nor U7772 (N_7772,N_1400,N_4448);
nor U7773 (N_7773,N_3475,N_2304);
or U7774 (N_7774,N_2077,N_1582);
or U7775 (N_7775,N_1386,N_2780);
nand U7776 (N_7776,N_1311,N_3050);
nor U7777 (N_7777,N_1230,N_966);
or U7778 (N_7778,N_2192,N_1773);
and U7779 (N_7779,N_3660,N_3811);
nor U7780 (N_7780,N_1003,N_536);
nand U7781 (N_7781,N_4502,N_2283);
or U7782 (N_7782,N_651,N_1332);
and U7783 (N_7783,N_192,N_151);
and U7784 (N_7784,N_2155,N_2480);
or U7785 (N_7785,N_2238,N_3951);
or U7786 (N_7786,N_1125,N_3138);
nand U7787 (N_7787,N_1235,N_1967);
nand U7788 (N_7788,N_20,N_4159);
nand U7789 (N_7789,N_2559,N_2675);
nor U7790 (N_7790,N_535,N_3814);
xor U7791 (N_7791,N_3709,N_1891);
nand U7792 (N_7792,N_1184,N_1051);
nand U7793 (N_7793,N_4840,N_1217);
or U7794 (N_7794,N_987,N_1580);
and U7795 (N_7795,N_4662,N_3979);
nand U7796 (N_7796,N_4587,N_2479);
nand U7797 (N_7797,N_3765,N_1716);
nand U7798 (N_7798,N_1074,N_2799);
nand U7799 (N_7799,N_4166,N_1203);
nor U7800 (N_7800,N_442,N_579);
nor U7801 (N_7801,N_1169,N_2031);
nor U7802 (N_7802,N_2534,N_27);
nand U7803 (N_7803,N_1758,N_1280);
nor U7804 (N_7804,N_1599,N_3884);
and U7805 (N_7805,N_2318,N_2119);
or U7806 (N_7806,N_4752,N_93);
nand U7807 (N_7807,N_842,N_3945);
nor U7808 (N_7808,N_2113,N_2716);
and U7809 (N_7809,N_4057,N_2519);
or U7810 (N_7810,N_4090,N_4151);
and U7811 (N_7811,N_3413,N_221);
nand U7812 (N_7812,N_3407,N_4057);
and U7813 (N_7813,N_26,N_3527);
and U7814 (N_7814,N_1309,N_2628);
or U7815 (N_7815,N_4745,N_1631);
or U7816 (N_7816,N_974,N_3900);
nand U7817 (N_7817,N_4810,N_119);
nand U7818 (N_7818,N_3052,N_3810);
nand U7819 (N_7819,N_1378,N_4566);
nand U7820 (N_7820,N_4956,N_688);
and U7821 (N_7821,N_2305,N_1506);
nand U7822 (N_7822,N_1483,N_1582);
nor U7823 (N_7823,N_2804,N_2997);
xnor U7824 (N_7824,N_3601,N_2274);
and U7825 (N_7825,N_629,N_4265);
nand U7826 (N_7826,N_2580,N_170);
nor U7827 (N_7827,N_2690,N_2047);
nor U7828 (N_7828,N_1642,N_4989);
nand U7829 (N_7829,N_1386,N_1093);
nor U7830 (N_7830,N_2917,N_166);
and U7831 (N_7831,N_4847,N_3699);
or U7832 (N_7832,N_1502,N_2655);
or U7833 (N_7833,N_3766,N_4921);
or U7834 (N_7834,N_537,N_108);
nor U7835 (N_7835,N_1226,N_364);
nor U7836 (N_7836,N_2215,N_4332);
and U7837 (N_7837,N_1293,N_2036);
or U7838 (N_7838,N_4280,N_1740);
nor U7839 (N_7839,N_3707,N_3688);
or U7840 (N_7840,N_4857,N_2077);
and U7841 (N_7841,N_3661,N_3226);
or U7842 (N_7842,N_518,N_4001);
nor U7843 (N_7843,N_340,N_936);
and U7844 (N_7844,N_1418,N_206);
nor U7845 (N_7845,N_3875,N_960);
nor U7846 (N_7846,N_2908,N_4220);
nand U7847 (N_7847,N_3923,N_2343);
nor U7848 (N_7848,N_604,N_3781);
nor U7849 (N_7849,N_3953,N_139);
and U7850 (N_7850,N_3685,N_171);
or U7851 (N_7851,N_1436,N_1141);
nor U7852 (N_7852,N_4676,N_1420);
nand U7853 (N_7853,N_1882,N_2339);
nand U7854 (N_7854,N_4411,N_4598);
nor U7855 (N_7855,N_4087,N_208);
nor U7856 (N_7856,N_1694,N_2674);
nand U7857 (N_7857,N_3470,N_1132);
or U7858 (N_7858,N_799,N_4252);
or U7859 (N_7859,N_4554,N_705);
or U7860 (N_7860,N_1384,N_2384);
nand U7861 (N_7861,N_3235,N_522);
nand U7862 (N_7862,N_293,N_1272);
nor U7863 (N_7863,N_508,N_3079);
or U7864 (N_7864,N_3976,N_3286);
nand U7865 (N_7865,N_303,N_3402);
xor U7866 (N_7866,N_3483,N_1796);
or U7867 (N_7867,N_1153,N_3948);
nand U7868 (N_7868,N_1060,N_2737);
and U7869 (N_7869,N_2764,N_1859);
and U7870 (N_7870,N_1075,N_312);
xnor U7871 (N_7871,N_2018,N_765);
or U7872 (N_7872,N_3897,N_351);
or U7873 (N_7873,N_2144,N_171);
or U7874 (N_7874,N_1813,N_4323);
nand U7875 (N_7875,N_1390,N_1555);
xor U7876 (N_7876,N_3133,N_2116);
or U7877 (N_7877,N_2018,N_3330);
or U7878 (N_7878,N_3190,N_1000);
and U7879 (N_7879,N_3271,N_3435);
and U7880 (N_7880,N_3041,N_481);
or U7881 (N_7881,N_3613,N_539);
nor U7882 (N_7882,N_4892,N_3632);
and U7883 (N_7883,N_2533,N_2357);
nand U7884 (N_7884,N_2461,N_4500);
and U7885 (N_7885,N_660,N_710);
and U7886 (N_7886,N_3924,N_4945);
and U7887 (N_7887,N_1357,N_3343);
xor U7888 (N_7888,N_4882,N_1605);
and U7889 (N_7889,N_620,N_2786);
or U7890 (N_7890,N_298,N_1655);
nor U7891 (N_7891,N_1849,N_1381);
nand U7892 (N_7892,N_4348,N_2437);
nand U7893 (N_7893,N_910,N_4142);
or U7894 (N_7894,N_2567,N_4584);
nor U7895 (N_7895,N_4079,N_2183);
nand U7896 (N_7896,N_150,N_2423);
nand U7897 (N_7897,N_3126,N_4811);
or U7898 (N_7898,N_3761,N_3641);
nor U7899 (N_7899,N_3460,N_3286);
nor U7900 (N_7900,N_2205,N_4053);
nand U7901 (N_7901,N_2766,N_1410);
nand U7902 (N_7902,N_1083,N_243);
nand U7903 (N_7903,N_1705,N_1986);
nor U7904 (N_7904,N_780,N_1798);
nand U7905 (N_7905,N_3910,N_1965);
and U7906 (N_7906,N_4263,N_2299);
nor U7907 (N_7907,N_453,N_3640);
nor U7908 (N_7908,N_299,N_3537);
xnor U7909 (N_7909,N_4614,N_448);
and U7910 (N_7910,N_3460,N_3435);
nand U7911 (N_7911,N_941,N_3199);
or U7912 (N_7912,N_2384,N_4716);
and U7913 (N_7913,N_517,N_4970);
and U7914 (N_7914,N_4946,N_2692);
or U7915 (N_7915,N_793,N_4023);
and U7916 (N_7916,N_3818,N_3414);
or U7917 (N_7917,N_4553,N_4170);
or U7918 (N_7918,N_4353,N_3842);
and U7919 (N_7919,N_2077,N_1489);
nor U7920 (N_7920,N_2472,N_998);
and U7921 (N_7921,N_2797,N_51);
and U7922 (N_7922,N_4081,N_3891);
and U7923 (N_7923,N_641,N_3940);
nor U7924 (N_7924,N_4941,N_1250);
nand U7925 (N_7925,N_2591,N_222);
or U7926 (N_7926,N_422,N_3697);
nand U7927 (N_7927,N_1820,N_2559);
nor U7928 (N_7928,N_4596,N_3744);
and U7929 (N_7929,N_4118,N_1451);
nand U7930 (N_7930,N_359,N_1576);
nor U7931 (N_7931,N_421,N_3116);
nor U7932 (N_7932,N_1434,N_512);
and U7933 (N_7933,N_4851,N_1641);
nand U7934 (N_7934,N_3640,N_2456);
or U7935 (N_7935,N_3937,N_2858);
or U7936 (N_7936,N_3764,N_1419);
nand U7937 (N_7937,N_522,N_2817);
or U7938 (N_7938,N_3459,N_3277);
nor U7939 (N_7939,N_1338,N_4900);
nand U7940 (N_7940,N_421,N_180);
and U7941 (N_7941,N_355,N_3638);
or U7942 (N_7942,N_3456,N_1462);
nand U7943 (N_7943,N_2587,N_2239);
and U7944 (N_7944,N_1736,N_2560);
nand U7945 (N_7945,N_3446,N_145);
or U7946 (N_7946,N_3169,N_4371);
xor U7947 (N_7947,N_2830,N_2337);
nand U7948 (N_7948,N_1434,N_2142);
or U7949 (N_7949,N_4225,N_2145);
or U7950 (N_7950,N_4518,N_4040);
or U7951 (N_7951,N_2764,N_1085);
or U7952 (N_7952,N_4792,N_4266);
nand U7953 (N_7953,N_3108,N_735);
nand U7954 (N_7954,N_2442,N_3009);
or U7955 (N_7955,N_514,N_1359);
or U7956 (N_7956,N_2868,N_4518);
or U7957 (N_7957,N_1251,N_1370);
and U7958 (N_7958,N_3603,N_199);
and U7959 (N_7959,N_4476,N_1702);
nor U7960 (N_7960,N_4906,N_2001);
nand U7961 (N_7961,N_2822,N_4042);
or U7962 (N_7962,N_1583,N_2338);
and U7963 (N_7963,N_4788,N_3610);
nor U7964 (N_7964,N_584,N_4407);
or U7965 (N_7965,N_1599,N_2306);
nand U7966 (N_7966,N_1306,N_625);
nand U7967 (N_7967,N_856,N_1174);
nand U7968 (N_7968,N_1344,N_313);
nor U7969 (N_7969,N_2463,N_1319);
or U7970 (N_7970,N_3150,N_232);
or U7971 (N_7971,N_3720,N_1646);
and U7972 (N_7972,N_4424,N_3640);
nor U7973 (N_7973,N_4879,N_1971);
and U7974 (N_7974,N_1676,N_405);
and U7975 (N_7975,N_4552,N_4241);
or U7976 (N_7976,N_4181,N_252);
nand U7977 (N_7977,N_2676,N_1623);
xor U7978 (N_7978,N_556,N_1137);
nand U7979 (N_7979,N_2553,N_3880);
or U7980 (N_7980,N_59,N_2576);
and U7981 (N_7981,N_469,N_2705);
and U7982 (N_7982,N_2602,N_1524);
nor U7983 (N_7983,N_3807,N_965);
or U7984 (N_7984,N_4804,N_995);
xnor U7985 (N_7985,N_652,N_1244);
nand U7986 (N_7986,N_1983,N_2483);
xor U7987 (N_7987,N_132,N_984);
nand U7988 (N_7988,N_179,N_3224);
or U7989 (N_7989,N_4487,N_266);
or U7990 (N_7990,N_4558,N_1218);
nand U7991 (N_7991,N_238,N_2380);
nor U7992 (N_7992,N_3440,N_3466);
and U7993 (N_7993,N_2310,N_452);
or U7994 (N_7994,N_4299,N_1979);
and U7995 (N_7995,N_4491,N_2399);
or U7996 (N_7996,N_841,N_1824);
or U7997 (N_7997,N_3415,N_926);
xor U7998 (N_7998,N_3612,N_596);
nor U7999 (N_7999,N_1792,N_2855);
nand U8000 (N_8000,N_2984,N_4328);
and U8001 (N_8001,N_1162,N_4494);
nor U8002 (N_8002,N_3984,N_1202);
and U8003 (N_8003,N_3768,N_4702);
or U8004 (N_8004,N_4393,N_4482);
nor U8005 (N_8005,N_1895,N_3987);
and U8006 (N_8006,N_4315,N_1406);
and U8007 (N_8007,N_1357,N_15);
nand U8008 (N_8008,N_875,N_3225);
or U8009 (N_8009,N_3911,N_2418);
or U8010 (N_8010,N_396,N_2263);
or U8011 (N_8011,N_2007,N_3336);
nor U8012 (N_8012,N_542,N_1687);
or U8013 (N_8013,N_2512,N_4630);
xnor U8014 (N_8014,N_3640,N_284);
and U8015 (N_8015,N_2986,N_2946);
nor U8016 (N_8016,N_838,N_783);
nand U8017 (N_8017,N_2030,N_4228);
and U8018 (N_8018,N_626,N_642);
nand U8019 (N_8019,N_554,N_1087);
and U8020 (N_8020,N_486,N_2231);
or U8021 (N_8021,N_3952,N_1833);
or U8022 (N_8022,N_1491,N_1016);
or U8023 (N_8023,N_3973,N_1584);
or U8024 (N_8024,N_1139,N_3463);
nor U8025 (N_8025,N_3811,N_3880);
nand U8026 (N_8026,N_3550,N_4017);
and U8027 (N_8027,N_1447,N_948);
and U8028 (N_8028,N_3763,N_2820);
or U8029 (N_8029,N_3821,N_1667);
or U8030 (N_8030,N_1407,N_675);
nor U8031 (N_8031,N_102,N_1779);
nand U8032 (N_8032,N_563,N_1282);
nand U8033 (N_8033,N_439,N_2710);
and U8034 (N_8034,N_2836,N_481);
nand U8035 (N_8035,N_2981,N_2232);
nor U8036 (N_8036,N_3775,N_267);
nor U8037 (N_8037,N_3923,N_1106);
or U8038 (N_8038,N_3790,N_667);
or U8039 (N_8039,N_2182,N_527);
or U8040 (N_8040,N_1414,N_3744);
nand U8041 (N_8041,N_443,N_976);
nor U8042 (N_8042,N_2828,N_2841);
nor U8043 (N_8043,N_3893,N_2102);
nor U8044 (N_8044,N_98,N_977);
nor U8045 (N_8045,N_2032,N_4566);
and U8046 (N_8046,N_67,N_4920);
and U8047 (N_8047,N_1827,N_2875);
or U8048 (N_8048,N_1811,N_1363);
or U8049 (N_8049,N_1530,N_255);
and U8050 (N_8050,N_3725,N_552);
and U8051 (N_8051,N_2672,N_2742);
nor U8052 (N_8052,N_3146,N_3741);
nor U8053 (N_8053,N_3738,N_852);
nor U8054 (N_8054,N_1685,N_4456);
or U8055 (N_8055,N_861,N_2324);
or U8056 (N_8056,N_504,N_1202);
or U8057 (N_8057,N_3194,N_4183);
and U8058 (N_8058,N_2572,N_1376);
nor U8059 (N_8059,N_2179,N_171);
or U8060 (N_8060,N_627,N_557);
nor U8061 (N_8061,N_192,N_3304);
nand U8062 (N_8062,N_2096,N_3513);
nand U8063 (N_8063,N_3205,N_1858);
or U8064 (N_8064,N_876,N_189);
or U8065 (N_8065,N_868,N_4627);
nor U8066 (N_8066,N_2691,N_899);
nand U8067 (N_8067,N_35,N_4828);
nor U8068 (N_8068,N_2695,N_581);
and U8069 (N_8069,N_52,N_2354);
nand U8070 (N_8070,N_1793,N_4978);
nand U8071 (N_8071,N_3155,N_1151);
nand U8072 (N_8072,N_1345,N_3226);
nand U8073 (N_8073,N_24,N_2085);
nor U8074 (N_8074,N_2581,N_3528);
or U8075 (N_8075,N_3515,N_37);
nor U8076 (N_8076,N_1340,N_2463);
or U8077 (N_8077,N_4909,N_3512);
nor U8078 (N_8078,N_4919,N_3354);
nor U8079 (N_8079,N_1359,N_3522);
nand U8080 (N_8080,N_3694,N_2168);
nand U8081 (N_8081,N_338,N_4480);
nor U8082 (N_8082,N_2286,N_3861);
nand U8083 (N_8083,N_4990,N_1633);
nand U8084 (N_8084,N_669,N_2106);
and U8085 (N_8085,N_3697,N_3325);
nor U8086 (N_8086,N_2611,N_884);
and U8087 (N_8087,N_3237,N_2331);
nor U8088 (N_8088,N_974,N_3805);
and U8089 (N_8089,N_2595,N_4867);
or U8090 (N_8090,N_624,N_2047);
xnor U8091 (N_8091,N_1569,N_2678);
nor U8092 (N_8092,N_1563,N_1061);
and U8093 (N_8093,N_1469,N_1054);
nand U8094 (N_8094,N_1112,N_3278);
xnor U8095 (N_8095,N_3396,N_624);
nor U8096 (N_8096,N_1338,N_2078);
nand U8097 (N_8097,N_4408,N_445);
or U8098 (N_8098,N_278,N_4954);
and U8099 (N_8099,N_4771,N_1462);
and U8100 (N_8100,N_837,N_856);
or U8101 (N_8101,N_2312,N_2419);
nand U8102 (N_8102,N_2463,N_1084);
or U8103 (N_8103,N_769,N_1127);
and U8104 (N_8104,N_3749,N_843);
nand U8105 (N_8105,N_3643,N_3081);
nor U8106 (N_8106,N_242,N_4292);
and U8107 (N_8107,N_4643,N_1714);
nor U8108 (N_8108,N_3075,N_2833);
or U8109 (N_8109,N_2997,N_4130);
or U8110 (N_8110,N_2526,N_234);
nor U8111 (N_8111,N_945,N_1914);
and U8112 (N_8112,N_1407,N_2920);
nor U8113 (N_8113,N_1374,N_3760);
and U8114 (N_8114,N_883,N_2356);
or U8115 (N_8115,N_4567,N_3881);
nor U8116 (N_8116,N_1968,N_3729);
and U8117 (N_8117,N_3806,N_1524);
or U8118 (N_8118,N_395,N_281);
nand U8119 (N_8119,N_3670,N_3039);
and U8120 (N_8120,N_4531,N_578);
nand U8121 (N_8121,N_2743,N_3295);
nor U8122 (N_8122,N_4800,N_1845);
nand U8123 (N_8123,N_1749,N_3575);
and U8124 (N_8124,N_3297,N_4369);
xnor U8125 (N_8125,N_4289,N_3864);
and U8126 (N_8126,N_3233,N_198);
and U8127 (N_8127,N_4426,N_2962);
nand U8128 (N_8128,N_3656,N_144);
nor U8129 (N_8129,N_3775,N_84);
nor U8130 (N_8130,N_506,N_4253);
or U8131 (N_8131,N_1558,N_2020);
nand U8132 (N_8132,N_4539,N_2829);
nor U8133 (N_8133,N_4115,N_1731);
or U8134 (N_8134,N_1082,N_4175);
nand U8135 (N_8135,N_823,N_3710);
nand U8136 (N_8136,N_883,N_3720);
nor U8137 (N_8137,N_191,N_2022);
nor U8138 (N_8138,N_3287,N_3153);
or U8139 (N_8139,N_3711,N_3860);
or U8140 (N_8140,N_2630,N_4553);
and U8141 (N_8141,N_3068,N_4281);
nand U8142 (N_8142,N_3897,N_2122);
and U8143 (N_8143,N_213,N_1523);
nand U8144 (N_8144,N_4339,N_2719);
nand U8145 (N_8145,N_3336,N_1223);
or U8146 (N_8146,N_1422,N_1476);
or U8147 (N_8147,N_3372,N_4555);
nor U8148 (N_8148,N_1698,N_712);
or U8149 (N_8149,N_3209,N_358);
nand U8150 (N_8150,N_3890,N_3649);
nand U8151 (N_8151,N_739,N_2747);
nor U8152 (N_8152,N_603,N_4964);
nor U8153 (N_8153,N_3230,N_4463);
or U8154 (N_8154,N_1132,N_4685);
or U8155 (N_8155,N_3701,N_3860);
nand U8156 (N_8156,N_4215,N_3900);
nand U8157 (N_8157,N_1754,N_2554);
nand U8158 (N_8158,N_2302,N_2660);
and U8159 (N_8159,N_2496,N_321);
and U8160 (N_8160,N_1814,N_4057);
nor U8161 (N_8161,N_997,N_4582);
and U8162 (N_8162,N_1005,N_4332);
xor U8163 (N_8163,N_3000,N_31);
and U8164 (N_8164,N_3888,N_970);
or U8165 (N_8165,N_2576,N_3988);
or U8166 (N_8166,N_1319,N_2577);
nand U8167 (N_8167,N_4403,N_4785);
nor U8168 (N_8168,N_1769,N_3377);
or U8169 (N_8169,N_4866,N_751);
nand U8170 (N_8170,N_3154,N_3336);
nand U8171 (N_8171,N_3353,N_4937);
nand U8172 (N_8172,N_1201,N_2956);
or U8173 (N_8173,N_4551,N_2430);
nand U8174 (N_8174,N_2645,N_814);
nor U8175 (N_8175,N_4186,N_17);
nor U8176 (N_8176,N_399,N_952);
nand U8177 (N_8177,N_3682,N_3024);
or U8178 (N_8178,N_2334,N_1943);
or U8179 (N_8179,N_1351,N_1800);
nor U8180 (N_8180,N_153,N_1951);
nand U8181 (N_8181,N_4580,N_962);
and U8182 (N_8182,N_2683,N_534);
and U8183 (N_8183,N_1740,N_3526);
and U8184 (N_8184,N_4100,N_1757);
nand U8185 (N_8185,N_340,N_835);
or U8186 (N_8186,N_1060,N_4332);
nor U8187 (N_8187,N_343,N_193);
and U8188 (N_8188,N_1081,N_1760);
nand U8189 (N_8189,N_2774,N_4713);
and U8190 (N_8190,N_3349,N_767);
or U8191 (N_8191,N_1904,N_928);
and U8192 (N_8192,N_2931,N_1919);
and U8193 (N_8193,N_1470,N_4505);
nand U8194 (N_8194,N_2484,N_4093);
or U8195 (N_8195,N_4728,N_334);
nand U8196 (N_8196,N_802,N_1788);
nand U8197 (N_8197,N_3608,N_2847);
nand U8198 (N_8198,N_1630,N_3338);
nor U8199 (N_8199,N_2694,N_2630);
nor U8200 (N_8200,N_4934,N_4342);
and U8201 (N_8201,N_3635,N_3208);
nand U8202 (N_8202,N_1667,N_2021);
nor U8203 (N_8203,N_3088,N_478);
nand U8204 (N_8204,N_3745,N_4686);
and U8205 (N_8205,N_414,N_4259);
and U8206 (N_8206,N_110,N_287);
nor U8207 (N_8207,N_2624,N_3604);
nor U8208 (N_8208,N_2231,N_1491);
nor U8209 (N_8209,N_544,N_1415);
nor U8210 (N_8210,N_774,N_2881);
or U8211 (N_8211,N_4354,N_3453);
and U8212 (N_8212,N_3321,N_2793);
nand U8213 (N_8213,N_1436,N_2762);
or U8214 (N_8214,N_4034,N_740);
or U8215 (N_8215,N_312,N_4719);
or U8216 (N_8216,N_600,N_1833);
and U8217 (N_8217,N_1305,N_307);
nand U8218 (N_8218,N_2496,N_2894);
nor U8219 (N_8219,N_1084,N_4905);
and U8220 (N_8220,N_2270,N_390);
and U8221 (N_8221,N_4444,N_279);
nand U8222 (N_8222,N_2702,N_544);
nand U8223 (N_8223,N_3528,N_890);
or U8224 (N_8224,N_1493,N_2334);
or U8225 (N_8225,N_528,N_3737);
and U8226 (N_8226,N_1463,N_729);
or U8227 (N_8227,N_4404,N_3749);
and U8228 (N_8228,N_3770,N_941);
nand U8229 (N_8229,N_1811,N_3845);
or U8230 (N_8230,N_3668,N_877);
nor U8231 (N_8231,N_3640,N_3532);
or U8232 (N_8232,N_309,N_4358);
nand U8233 (N_8233,N_2088,N_1938);
and U8234 (N_8234,N_3491,N_2381);
or U8235 (N_8235,N_1442,N_1201);
nand U8236 (N_8236,N_2583,N_1461);
nor U8237 (N_8237,N_939,N_4320);
and U8238 (N_8238,N_4285,N_1529);
nor U8239 (N_8239,N_1940,N_3492);
and U8240 (N_8240,N_4911,N_2266);
nand U8241 (N_8241,N_3910,N_1675);
and U8242 (N_8242,N_847,N_2728);
nor U8243 (N_8243,N_3490,N_46);
or U8244 (N_8244,N_21,N_999);
nand U8245 (N_8245,N_3506,N_4605);
nor U8246 (N_8246,N_1314,N_1261);
nor U8247 (N_8247,N_1750,N_802);
or U8248 (N_8248,N_4116,N_4745);
nor U8249 (N_8249,N_932,N_4436);
or U8250 (N_8250,N_4039,N_377);
or U8251 (N_8251,N_402,N_867);
nand U8252 (N_8252,N_42,N_322);
nand U8253 (N_8253,N_1463,N_1889);
nor U8254 (N_8254,N_1750,N_2120);
or U8255 (N_8255,N_2238,N_1562);
nand U8256 (N_8256,N_4737,N_558);
and U8257 (N_8257,N_3382,N_1227);
nand U8258 (N_8258,N_4926,N_2887);
nor U8259 (N_8259,N_395,N_1943);
or U8260 (N_8260,N_4085,N_557);
and U8261 (N_8261,N_3362,N_1404);
nand U8262 (N_8262,N_736,N_2818);
nor U8263 (N_8263,N_773,N_1866);
nor U8264 (N_8264,N_2272,N_3484);
or U8265 (N_8265,N_337,N_889);
and U8266 (N_8266,N_4382,N_1328);
and U8267 (N_8267,N_1346,N_4104);
and U8268 (N_8268,N_236,N_325);
nand U8269 (N_8269,N_3514,N_2635);
or U8270 (N_8270,N_2555,N_3975);
nand U8271 (N_8271,N_113,N_2764);
nor U8272 (N_8272,N_1939,N_260);
and U8273 (N_8273,N_3791,N_1327);
nand U8274 (N_8274,N_3743,N_3804);
or U8275 (N_8275,N_4595,N_4787);
nand U8276 (N_8276,N_4179,N_1247);
nand U8277 (N_8277,N_4871,N_3435);
and U8278 (N_8278,N_1464,N_2226);
and U8279 (N_8279,N_3888,N_585);
nand U8280 (N_8280,N_2538,N_3283);
and U8281 (N_8281,N_2812,N_2207);
or U8282 (N_8282,N_1405,N_3309);
and U8283 (N_8283,N_2652,N_4287);
or U8284 (N_8284,N_3036,N_4350);
nor U8285 (N_8285,N_2510,N_3925);
and U8286 (N_8286,N_3640,N_3925);
or U8287 (N_8287,N_333,N_3950);
nand U8288 (N_8288,N_4005,N_1235);
nor U8289 (N_8289,N_2122,N_973);
nand U8290 (N_8290,N_1528,N_186);
and U8291 (N_8291,N_192,N_2811);
nand U8292 (N_8292,N_2058,N_3892);
nor U8293 (N_8293,N_2329,N_4074);
nand U8294 (N_8294,N_2207,N_1278);
nand U8295 (N_8295,N_431,N_1790);
or U8296 (N_8296,N_3325,N_2388);
nand U8297 (N_8297,N_4886,N_3506);
or U8298 (N_8298,N_2167,N_34);
nand U8299 (N_8299,N_4422,N_3519);
nand U8300 (N_8300,N_1548,N_587);
and U8301 (N_8301,N_1560,N_3934);
or U8302 (N_8302,N_1911,N_3708);
nor U8303 (N_8303,N_1601,N_4874);
nand U8304 (N_8304,N_4057,N_1083);
nor U8305 (N_8305,N_503,N_2293);
nor U8306 (N_8306,N_2538,N_4056);
nor U8307 (N_8307,N_1020,N_4912);
nor U8308 (N_8308,N_3209,N_3811);
nand U8309 (N_8309,N_1291,N_4922);
and U8310 (N_8310,N_2860,N_3832);
nor U8311 (N_8311,N_2947,N_240);
nor U8312 (N_8312,N_561,N_1406);
nor U8313 (N_8313,N_3515,N_2879);
and U8314 (N_8314,N_714,N_2664);
and U8315 (N_8315,N_1952,N_4451);
and U8316 (N_8316,N_801,N_695);
nand U8317 (N_8317,N_3591,N_4796);
and U8318 (N_8318,N_2789,N_4538);
and U8319 (N_8319,N_4999,N_993);
nand U8320 (N_8320,N_941,N_339);
nor U8321 (N_8321,N_4316,N_4564);
and U8322 (N_8322,N_3793,N_2342);
nand U8323 (N_8323,N_1158,N_2392);
and U8324 (N_8324,N_3747,N_2044);
nand U8325 (N_8325,N_691,N_4667);
nand U8326 (N_8326,N_4101,N_1525);
and U8327 (N_8327,N_3178,N_1436);
xor U8328 (N_8328,N_358,N_1230);
nor U8329 (N_8329,N_4141,N_848);
or U8330 (N_8330,N_1473,N_3881);
and U8331 (N_8331,N_1108,N_2212);
nor U8332 (N_8332,N_2392,N_4906);
nand U8333 (N_8333,N_3883,N_1345);
or U8334 (N_8334,N_4771,N_3074);
or U8335 (N_8335,N_2351,N_4742);
nor U8336 (N_8336,N_4099,N_315);
or U8337 (N_8337,N_3852,N_4696);
nand U8338 (N_8338,N_446,N_3253);
nand U8339 (N_8339,N_4110,N_2723);
nand U8340 (N_8340,N_1388,N_4146);
nand U8341 (N_8341,N_2980,N_2302);
nand U8342 (N_8342,N_2458,N_2599);
and U8343 (N_8343,N_3698,N_3708);
nand U8344 (N_8344,N_3657,N_4920);
nor U8345 (N_8345,N_4071,N_3651);
and U8346 (N_8346,N_3902,N_1511);
and U8347 (N_8347,N_3627,N_1966);
xor U8348 (N_8348,N_1157,N_3971);
nand U8349 (N_8349,N_3873,N_2967);
or U8350 (N_8350,N_3680,N_3445);
and U8351 (N_8351,N_3550,N_4617);
or U8352 (N_8352,N_512,N_3498);
or U8353 (N_8353,N_2483,N_2254);
and U8354 (N_8354,N_644,N_2962);
nor U8355 (N_8355,N_1710,N_4943);
nor U8356 (N_8356,N_4567,N_4488);
nor U8357 (N_8357,N_2265,N_4034);
and U8358 (N_8358,N_4316,N_1084);
and U8359 (N_8359,N_819,N_4431);
and U8360 (N_8360,N_2181,N_2966);
nand U8361 (N_8361,N_3170,N_208);
or U8362 (N_8362,N_1339,N_1329);
nand U8363 (N_8363,N_373,N_1456);
nor U8364 (N_8364,N_2855,N_4051);
nor U8365 (N_8365,N_3176,N_453);
and U8366 (N_8366,N_3631,N_2569);
or U8367 (N_8367,N_3663,N_3898);
nor U8368 (N_8368,N_1689,N_305);
and U8369 (N_8369,N_875,N_1468);
nor U8370 (N_8370,N_500,N_322);
or U8371 (N_8371,N_3996,N_4563);
and U8372 (N_8372,N_1214,N_3527);
or U8373 (N_8373,N_4290,N_674);
or U8374 (N_8374,N_2202,N_1869);
nand U8375 (N_8375,N_354,N_71);
or U8376 (N_8376,N_230,N_3997);
nand U8377 (N_8377,N_3528,N_1694);
nand U8378 (N_8378,N_4738,N_4097);
nor U8379 (N_8379,N_2953,N_1361);
and U8380 (N_8380,N_4570,N_992);
and U8381 (N_8381,N_1814,N_4008);
or U8382 (N_8382,N_4225,N_2146);
and U8383 (N_8383,N_4172,N_3275);
and U8384 (N_8384,N_2699,N_3333);
and U8385 (N_8385,N_2082,N_2176);
nand U8386 (N_8386,N_1086,N_667);
and U8387 (N_8387,N_1292,N_2023);
nor U8388 (N_8388,N_3827,N_160);
nor U8389 (N_8389,N_340,N_1636);
nor U8390 (N_8390,N_2007,N_1505);
nor U8391 (N_8391,N_3884,N_4663);
or U8392 (N_8392,N_1871,N_1849);
nor U8393 (N_8393,N_736,N_3140);
nor U8394 (N_8394,N_149,N_1460);
and U8395 (N_8395,N_4056,N_1795);
and U8396 (N_8396,N_307,N_1401);
or U8397 (N_8397,N_1262,N_211);
nor U8398 (N_8398,N_1119,N_1606);
or U8399 (N_8399,N_1571,N_2362);
or U8400 (N_8400,N_4510,N_2060);
or U8401 (N_8401,N_1081,N_4679);
nand U8402 (N_8402,N_396,N_3920);
nand U8403 (N_8403,N_3990,N_4159);
and U8404 (N_8404,N_4201,N_27);
xor U8405 (N_8405,N_3552,N_4367);
nand U8406 (N_8406,N_4154,N_4350);
nand U8407 (N_8407,N_1800,N_4667);
nor U8408 (N_8408,N_657,N_3912);
nand U8409 (N_8409,N_2198,N_591);
and U8410 (N_8410,N_3436,N_3020);
or U8411 (N_8411,N_3629,N_4184);
or U8412 (N_8412,N_2523,N_516);
nor U8413 (N_8413,N_229,N_4397);
or U8414 (N_8414,N_852,N_2430);
or U8415 (N_8415,N_4373,N_411);
and U8416 (N_8416,N_75,N_1671);
or U8417 (N_8417,N_4090,N_3561);
and U8418 (N_8418,N_4125,N_4269);
and U8419 (N_8419,N_4504,N_1128);
nor U8420 (N_8420,N_4984,N_786);
nor U8421 (N_8421,N_4199,N_2156);
nor U8422 (N_8422,N_192,N_4928);
nor U8423 (N_8423,N_3469,N_2250);
nand U8424 (N_8424,N_4701,N_4382);
and U8425 (N_8425,N_1177,N_4381);
and U8426 (N_8426,N_1532,N_3523);
or U8427 (N_8427,N_4011,N_157);
or U8428 (N_8428,N_4419,N_2378);
and U8429 (N_8429,N_4785,N_4343);
or U8430 (N_8430,N_4326,N_2882);
and U8431 (N_8431,N_716,N_4573);
nor U8432 (N_8432,N_1361,N_1217);
nand U8433 (N_8433,N_543,N_3949);
or U8434 (N_8434,N_4478,N_995);
and U8435 (N_8435,N_4813,N_4872);
or U8436 (N_8436,N_3087,N_1879);
and U8437 (N_8437,N_630,N_2514);
or U8438 (N_8438,N_430,N_4941);
or U8439 (N_8439,N_1832,N_1079);
nand U8440 (N_8440,N_3678,N_604);
and U8441 (N_8441,N_1619,N_2115);
and U8442 (N_8442,N_930,N_1742);
nand U8443 (N_8443,N_4057,N_782);
nor U8444 (N_8444,N_4776,N_258);
nor U8445 (N_8445,N_4589,N_909);
nor U8446 (N_8446,N_3591,N_2675);
and U8447 (N_8447,N_1163,N_1056);
and U8448 (N_8448,N_3655,N_3665);
nor U8449 (N_8449,N_3487,N_995);
nand U8450 (N_8450,N_1972,N_4772);
nor U8451 (N_8451,N_252,N_2911);
or U8452 (N_8452,N_2367,N_4956);
and U8453 (N_8453,N_3432,N_4541);
and U8454 (N_8454,N_2882,N_2608);
nor U8455 (N_8455,N_4640,N_319);
nor U8456 (N_8456,N_1693,N_516);
nor U8457 (N_8457,N_1836,N_2100);
nand U8458 (N_8458,N_3389,N_4608);
or U8459 (N_8459,N_4464,N_1329);
or U8460 (N_8460,N_1440,N_1076);
nor U8461 (N_8461,N_4428,N_3933);
nor U8462 (N_8462,N_3118,N_3470);
nor U8463 (N_8463,N_1357,N_2710);
or U8464 (N_8464,N_1088,N_2422);
and U8465 (N_8465,N_907,N_4137);
nor U8466 (N_8466,N_2967,N_3882);
nor U8467 (N_8467,N_2758,N_2987);
or U8468 (N_8468,N_789,N_573);
nor U8469 (N_8469,N_3644,N_2080);
and U8470 (N_8470,N_2647,N_4648);
or U8471 (N_8471,N_2796,N_2351);
or U8472 (N_8472,N_2939,N_4408);
and U8473 (N_8473,N_3786,N_308);
nand U8474 (N_8474,N_435,N_509);
or U8475 (N_8475,N_1731,N_1611);
nand U8476 (N_8476,N_4865,N_3929);
nor U8477 (N_8477,N_82,N_1461);
or U8478 (N_8478,N_2374,N_1509);
nor U8479 (N_8479,N_4144,N_2655);
nand U8480 (N_8480,N_2807,N_3419);
nor U8481 (N_8481,N_4911,N_4251);
or U8482 (N_8482,N_1853,N_798);
and U8483 (N_8483,N_1441,N_4553);
or U8484 (N_8484,N_1113,N_1488);
and U8485 (N_8485,N_3164,N_2543);
and U8486 (N_8486,N_3843,N_4413);
nand U8487 (N_8487,N_4183,N_242);
or U8488 (N_8488,N_1416,N_2946);
nor U8489 (N_8489,N_3894,N_3799);
nand U8490 (N_8490,N_4725,N_2844);
nor U8491 (N_8491,N_3842,N_3986);
nand U8492 (N_8492,N_258,N_2559);
or U8493 (N_8493,N_415,N_2912);
nand U8494 (N_8494,N_3920,N_1273);
nand U8495 (N_8495,N_1214,N_1745);
nand U8496 (N_8496,N_1369,N_404);
nand U8497 (N_8497,N_2382,N_4378);
or U8498 (N_8498,N_825,N_1513);
nand U8499 (N_8499,N_3630,N_42);
nand U8500 (N_8500,N_282,N_1637);
nor U8501 (N_8501,N_779,N_4010);
nor U8502 (N_8502,N_4571,N_1479);
or U8503 (N_8503,N_150,N_3663);
nor U8504 (N_8504,N_3485,N_4739);
nand U8505 (N_8505,N_3627,N_4479);
or U8506 (N_8506,N_1939,N_2120);
and U8507 (N_8507,N_1059,N_876);
nor U8508 (N_8508,N_2028,N_2716);
nor U8509 (N_8509,N_4972,N_848);
and U8510 (N_8510,N_806,N_4049);
nor U8511 (N_8511,N_4857,N_2899);
nor U8512 (N_8512,N_3594,N_2159);
nor U8513 (N_8513,N_4836,N_3811);
nor U8514 (N_8514,N_4399,N_4433);
nand U8515 (N_8515,N_1884,N_4602);
and U8516 (N_8516,N_3837,N_494);
and U8517 (N_8517,N_2284,N_1378);
or U8518 (N_8518,N_2644,N_3943);
and U8519 (N_8519,N_2131,N_212);
or U8520 (N_8520,N_1546,N_2838);
and U8521 (N_8521,N_955,N_4340);
nor U8522 (N_8522,N_4957,N_3734);
nand U8523 (N_8523,N_464,N_3121);
nor U8524 (N_8524,N_4109,N_4997);
nand U8525 (N_8525,N_3960,N_4549);
nor U8526 (N_8526,N_413,N_1901);
xnor U8527 (N_8527,N_3962,N_999);
and U8528 (N_8528,N_5,N_1337);
nor U8529 (N_8529,N_3122,N_1313);
or U8530 (N_8530,N_2834,N_2329);
nor U8531 (N_8531,N_888,N_517);
or U8532 (N_8532,N_3961,N_3390);
nor U8533 (N_8533,N_1711,N_870);
nand U8534 (N_8534,N_4636,N_3429);
and U8535 (N_8535,N_4647,N_4455);
nor U8536 (N_8536,N_2798,N_2522);
or U8537 (N_8537,N_4675,N_2599);
and U8538 (N_8538,N_2519,N_4975);
nor U8539 (N_8539,N_2200,N_4660);
and U8540 (N_8540,N_429,N_2286);
nor U8541 (N_8541,N_878,N_81);
nand U8542 (N_8542,N_4337,N_466);
nand U8543 (N_8543,N_2261,N_1036);
nor U8544 (N_8544,N_2391,N_3259);
nor U8545 (N_8545,N_4371,N_1099);
nor U8546 (N_8546,N_3212,N_2615);
nor U8547 (N_8547,N_692,N_2888);
or U8548 (N_8548,N_2655,N_2342);
nor U8549 (N_8549,N_4497,N_2665);
nor U8550 (N_8550,N_4234,N_2880);
nand U8551 (N_8551,N_723,N_1122);
nor U8552 (N_8552,N_672,N_224);
and U8553 (N_8553,N_3713,N_2977);
nor U8554 (N_8554,N_2802,N_3109);
and U8555 (N_8555,N_2206,N_2713);
and U8556 (N_8556,N_712,N_3703);
nor U8557 (N_8557,N_2294,N_4007);
or U8558 (N_8558,N_471,N_3842);
nor U8559 (N_8559,N_379,N_320);
and U8560 (N_8560,N_3106,N_1367);
and U8561 (N_8561,N_4921,N_3764);
nand U8562 (N_8562,N_472,N_4654);
nand U8563 (N_8563,N_4616,N_4968);
and U8564 (N_8564,N_1715,N_1038);
and U8565 (N_8565,N_2221,N_969);
nand U8566 (N_8566,N_3816,N_3858);
or U8567 (N_8567,N_3275,N_318);
nand U8568 (N_8568,N_1459,N_3788);
and U8569 (N_8569,N_4600,N_1630);
or U8570 (N_8570,N_4931,N_4626);
or U8571 (N_8571,N_769,N_835);
nand U8572 (N_8572,N_4340,N_4092);
nor U8573 (N_8573,N_4185,N_4924);
nor U8574 (N_8574,N_3485,N_2603);
or U8575 (N_8575,N_171,N_931);
nand U8576 (N_8576,N_2677,N_4614);
nor U8577 (N_8577,N_3260,N_3126);
or U8578 (N_8578,N_1341,N_3673);
nor U8579 (N_8579,N_46,N_4899);
nand U8580 (N_8580,N_317,N_4641);
nand U8581 (N_8581,N_2246,N_4167);
and U8582 (N_8582,N_4649,N_770);
xor U8583 (N_8583,N_2259,N_3680);
nand U8584 (N_8584,N_556,N_2611);
and U8585 (N_8585,N_2655,N_1256);
or U8586 (N_8586,N_2146,N_2064);
or U8587 (N_8587,N_1935,N_3773);
nor U8588 (N_8588,N_4653,N_1113);
or U8589 (N_8589,N_379,N_3291);
nand U8590 (N_8590,N_254,N_1974);
nor U8591 (N_8591,N_653,N_2148);
nor U8592 (N_8592,N_236,N_3565);
nor U8593 (N_8593,N_4117,N_4248);
nor U8594 (N_8594,N_937,N_2035);
and U8595 (N_8595,N_3489,N_1037);
or U8596 (N_8596,N_2412,N_2244);
or U8597 (N_8597,N_4076,N_3389);
nand U8598 (N_8598,N_2538,N_2275);
nor U8599 (N_8599,N_76,N_2123);
nand U8600 (N_8600,N_433,N_313);
nor U8601 (N_8601,N_3288,N_4738);
nor U8602 (N_8602,N_2517,N_4682);
or U8603 (N_8603,N_2350,N_1370);
or U8604 (N_8604,N_2967,N_1303);
or U8605 (N_8605,N_4251,N_1297);
nor U8606 (N_8606,N_4028,N_3782);
or U8607 (N_8607,N_2692,N_350);
or U8608 (N_8608,N_1586,N_1446);
or U8609 (N_8609,N_2265,N_2670);
nor U8610 (N_8610,N_2313,N_521);
or U8611 (N_8611,N_3274,N_3465);
and U8612 (N_8612,N_941,N_2036);
or U8613 (N_8613,N_400,N_2567);
or U8614 (N_8614,N_2896,N_1955);
or U8615 (N_8615,N_1197,N_1799);
nor U8616 (N_8616,N_3247,N_4846);
and U8617 (N_8617,N_1221,N_426);
and U8618 (N_8618,N_3555,N_3281);
nand U8619 (N_8619,N_1350,N_3535);
nor U8620 (N_8620,N_3216,N_1118);
nand U8621 (N_8621,N_2171,N_4912);
nor U8622 (N_8622,N_2946,N_4342);
and U8623 (N_8623,N_559,N_4769);
and U8624 (N_8624,N_2634,N_256);
nor U8625 (N_8625,N_2921,N_4049);
nand U8626 (N_8626,N_3780,N_1587);
or U8627 (N_8627,N_3354,N_3270);
or U8628 (N_8628,N_2938,N_2134);
nand U8629 (N_8629,N_4382,N_1672);
and U8630 (N_8630,N_1033,N_1244);
and U8631 (N_8631,N_2491,N_4147);
nor U8632 (N_8632,N_424,N_1425);
nand U8633 (N_8633,N_3515,N_798);
or U8634 (N_8634,N_4672,N_1613);
or U8635 (N_8635,N_359,N_3143);
and U8636 (N_8636,N_3580,N_4484);
and U8637 (N_8637,N_2292,N_4390);
or U8638 (N_8638,N_4521,N_2045);
or U8639 (N_8639,N_1279,N_2529);
and U8640 (N_8640,N_904,N_3743);
nand U8641 (N_8641,N_2381,N_1788);
and U8642 (N_8642,N_3839,N_3236);
nor U8643 (N_8643,N_2447,N_1037);
or U8644 (N_8644,N_3379,N_1459);
and U8645 (N_8645,N_1687,N_3812);
xor U8646 (N_8646,N_3191,N_4672);
or U8647 (N_8647,N_1313,N_2988);
nand U8648 (N_8648,N_3479,N_2293);
xor U8649 (N_8649,N_321,N_3718);
or U8650 (N_8650,N_683,N_1496);
nor U8651 (N_8651,N_904,N_4232);
or U8652 (N_8652,N_2193,N_1390);
nand U8653 (N_8653,N_2349,N_511);
and U8654 (N_8654,N_2795,N_104);
xnor U8655 (N_8655,N_1621,N_2645);
or U8656 (N_8656,N_352,N_1156);
and U8657 (N_8657,N_767,N_2845);
nand U8658 (N_8658,N_4935,N_2538);
nand U8659 (N_8659,N_2887,N_359);
and U8660 (N_8660,N_2447,N_4549);
nand U8661 (N_8661,N_2394,N_1478);
nand U8662 (N_8662,N_554,N_2398);
and U8663 (N_8663,N_3539,N_2935);
and U8664 (N_8664,N_820,N_2492);
nand U8665 (N_8665,N_3941,N_1106);
nand U8666 (N_8666,N_246,N_2757);
nand U8667 (N_8667,N_3017,N_4208);
and U8668 (N_8668,N_3481,N_1377);
nand U8669 (N_8669,N_4626,N_770);
and U8670 (N_8670,N_4889,N_41);
or U8671 (N_8671,N_2983,N_3307);
or U8672 (N_8672,N_1651,N_281);
and U8673 (N_8673,N_1410,N_2349);
nor U8674 (N_8674,N_3366,N_3530);
and U8675 (N_8675,N_99,N_3938);
nor U8676 (N_8676,N_2225,N_1726);
nand U8677 (N_8677,N_2750,N_3085);
nor U8678 (N_8678,N_1898,N_2943);
nand U8679 (N_8679,N_3581,N_3310);
or U8680 (N_8680,N_2835,N_3126);
nor U8681 (N_8681,N_4269,N_1235);
or U8682 (N_8682,N_1317,N_1652);
xor U8683 (N_8683,N_3023,N_2907);
and U8684 (N_8684,N_4810,N_3351);
and U8685 (N_8685,N_122,N_3423);
xor U8686 (N_8686,N_2421,N_1296);
nor U8687 (N_8687,N_3401,N_1305);
nor U8688 (N_8688,N_1991,N_4792);
or U8689 (N_8689,N_1294,N_4801);
or U8690 (N_8690,N_3554,N_524);
nor U8691 (N_8691,N_3998,N_1597);
nor U8692 (N_8692,N_3510,N_103);
or U8693 (N_8693,N_3452,N_1127);
nor U8694 (N_8694,N_3730,N_246);
nor U8695 (N_8695,N_1426,N_1366);
and U8696 (N_8696,N_2388,N_4681);
nand U8697 (N_8697,N_4013,N_2641);
or U8698 (N_8698,N_2130,N_188);
or U8699 (N_8699,N_652,N_784);
nor U8700 (N_8700,N_22,N_2065);
or U8701 (N_8701,N_3185,N_2327);
or U8702 (N_8702,N_619,N_679);
and U8703 (N_8703,N_2353,N_1911);
and U8704 (N_8704,N_4973,N_865);
nand U8705 (N_8705,N_3071,N_1778);
nor U8706 (N_8706,N_2896,N_3929);
nor U8707 (N_8707,N_3320,N_4313);
or U8708 (N_8708,N_196,N_312);
or U8709 (N_8709,N_2078,N_464);
or U8710 (N_8710,N_2549,N_4314);
nor U8711 (N_8711,N_2103,N_3174);
or U8712 (N_8712,N_462,N_1316);
nand U8713 (N_8713,N_1288,N_640);
nand U8714 (N_8714,N_1916,N_3056);
and U8715 (N_8715,N_4411,N_537);
nand U8716 (N_8716,N_1171,N_272);
or U8717 (N_8717,N_3473,N_1323);
xnor U8718 (N_8718,N_2952,N_2463);
nor U8719 (N_8719,N_1826,N_1489);
or U8720 (N_8720,N_3402,N_3168);
nor U8721 (N_8721,N_3798,N_1713);
nand U8722 (N_8722,N_3732,N_4255);
and U8723 (N_8723,N_797,N_2097);
or U8724 (N_8724,N_3231,N_1759);
or U8725 (N_8725,N_108,N_4469);
or U8726 (N_8726,N_2135,N_1461);
or U8727 (N_8727,N_4161,N_3948);
or U8728 (N_8728,N_4255,N_1337);
or U8729 (N_8729,N_922,N_3124);
nand U8730 (N_8730,N_3352,N_4030);
and U8731 (N_8731,N_1394,N_3243);
and U8732 (N_8732,N_4874,N_3412);
nor U8733 (N_8733,N_2796,N_4199);
nand U8734 (N_8734,N_3753,N_4735);
or U8735 (N_8735,N_1161,N_2563);
and U8736 (N_8736,N_4501,N_4545);
nand U8737 (N_8737,N_1202,N_706);
nor U8738 (N_8738,N_1282,N_179);
or U8739 (N_8739,N_2896,N_366);
or U8740 (N_8740,N_357,N_3779);
nand U8741 (N_8741,N_2882,N_3425);
and U8742 (N_8742,N_874,N_4376);
and U8743 (N_8743,N_1452,N_3267);
nor U8744 (N_8744,N_1866,N_3802);
nand U8745 (N_8745,N_4898,N_2121);
and U8746 (N_8746,N_1919,N_4340);
nor U8747 (N_8747,N_4962,N_1302);
nand U8748 (N_8748,N_3932,N_3536);
or U8749 (N_8749,N_2178,N_4981);
nor U8750 (N_8750,N_3629,N_645);
or U8751 (N_8751,N_4968,N_104);
nand U8752 (N_8752,N_3787,N_1822);
and U8753 (N_8753,N_1591,N_1728);
nor U8754 (N_8754,N_840,N_3922);
nor U8755 (N_8755,N_142,N_4022);
or U8756 (N_8756,N_2948,N_3561);
nand U8757 (N_8757,N_121,N_2205);
or U8758 (N_8758,N_1444,N_4008);
or U8759 (N_8759,N_2300,N_4913);
nand U8760 (N_8760,N_4093,N_3639);
nor U8761 (N_8761,N_4581,N_2412);
nand U8762 (N_8762,N_4922,N_1276);
or U8763 (N_8763,N_462,N_2486);
and U8764 (N_8764,N_2967,N_1763);
or U8765 (N_8765,N_1198,N_2970);
nand U8766 (N_8766,N_4635,N_4092);
nor U8767 (N_8767,N_3974,N_1005);
nand U8768 (N_8768,N_806,N_2280);
or U8769 (N_8769,N_1885,N_4929);
nor U8770 (N_8770,N_148,N_511);
nand U8771 (N_8771,N_1484,N_4962);
nand U8772 (N_8772,N_2760,N_1274);
nor U8773 (N_8773,N_3962,N_3014);
and U8774 (N_8774,N_732,N_2724);
nor U8775 (N_8775,N_102,N_2261);
or U8776 (N_8776,N_2452,N_4600);
and U8777 (N_8777,N_2948,N_647);
or U8778 (N_8778,N_3973,N_3534);
or U8779 (N_8779,N_1819,N_3248);
nand U8780 (N_8780,N_4364,N_4413);
or U8781 (N_8781,N_760,N_535);
xor U8782 (N_8782,N_4946,N_493);
and U8783 (N_8783,N_4077,N_2699);
and U8784 (N_8784,N_4493,N_3710);
or U8785 (N_8785,N_3230,N_4126);
or U8786 (N_8786,N_3008,N_2062);
xnor U8787 (N_8787,N_4401,N_2397);
and U8788 (N_8788,N_4072,N_4177);
nand U8789 (N_8789,N_4939,N_3234);
xor U8790 (N_8790,N_218,N_920);
nor U8791 (N_8791,N_1555,N_4546);
nand U8792 (N_8792,N_4358,N_2877);
xnor U8793 (N_8793,N_410,N_2046);
and U8794 (N_8794,N_1758,N_1907);
nand U8795 (N_8795,N_186,N_1868);
nor U8796 (N_8796,N_1032,N_4923);
and U8797 (N_8797,N_3796,N_4029);
or U8798 (N_8798,N_2545,N_4635);
and U8799 (N_8799,N_2124,N_1153);
nor U8800 (N_8800,N_2592,N_4208);
nor U8801 (N_8801,N_2537,N_969);
nor U8802 (N_8802,N_3749,N_2263);
and U8803 (N_8803,N_4723,N_1955);
or U8804 (N_8804,N_439,N_337);
nor U8805 (N_8805,N_4564,N_2874);
nand U8806 (N_8806,N_1119,N_623);
nor U8807 (N_8807,N_2864,N_4342);
nand U8808 (N_8808,N_4731,N_467);
nor U8809 (N_8809,N_80,N_2482);
and U8810 (N_8810,N_19,N_1147);
and U8811 (N_8811,N_4135,N_1905);
or U8812 (N_8812,N_4033,N_4069);
nand U8813 (N_8813,N_4630,N_2673);
nor U8814 (N_8814,N_3232,N_426);
and U8815 (N_8815,N_4986,N_3696);
or U8816 (N_8816,N_2950,N_4036);
or U8817 (N_8817,N_1397,N_3477);
nand U8818 (N_8818,N_3389,N_3574);
xor U8819 (N_8819,N_1797,N_2773);
or U8820 (N_8820,N_2779,N_3368);
or U8821 (N_8821,N_220,N_4171);
nand U8822 (N_8822,N_2762,N_287);
nor U8823 (N_8823,N_3036,N_4826);
nand U8824 (N_8824,N_3191,N_842);
nand U8825 (N_8825,N_797,N_3450);
or U8826 (N_8826,N_289,N_4734);
nor U8827 (N_8827,N_4688,N_2611);
or U8828 (N_8828,N_4216,N_3230);
nor U8829 (N_8829,N_1081,N_3317);
and U8830 (N_8830,N_4678,N_541);
and U8831 (N_8831,N_268,N_4847);
or U8832 (N_8832,N_2344,N_1685);
and U8833 (N_8833,N_3680,N_4583);
and U8834 (N_8834,N_1888,N_146);
and U8835 (N_8835,N_2990,N_4686);
nand U8836 (N_8836,N_1400,N_168);
nor U8837 (N_8837,N_3012,N_1731);
or U8838 (N_8838,N_1777,N_3563);
or U8839 (N_8839,N_1946,N_4383);
nand U8840 (N_8840,N_4448,N_1258);
and U8841 (N_8841,N_154,N_1800);
and U8842 (N_8842,N_4527,N_1959);
nand U8843 (N_8843,N_1926,N_1743);
nand U8844 (N_8844,N_1576,N_2164);
or U8845 (N_8845,N_3479,N_4206);
xor U8846 (N_8846,N_3389,N_4117);
nor U8847 (N_8847,N_3788,N_4462);
and U8848 (N_8848,N_4478,N_259);
nor U8849 (N_8849,N_1925,N_4926);
and U8850 (N_8850,N_2831,N_102);
nor U8851 (N_8851,N_173,N_255);
and U8852 (N_8852,N_10,N_3167);
nor U8853 (N_8853,N_2563,N_3126);
and U8854 (N_8854,N_4722,N_2136);
or U8855 (N_8855,N_4056,N_36);
or U8856 (N_8856,N_3078,N_2639);
and U8857 (N_8857,N_2643,N_2591);
nor U8858 (N_8858,N_3479,N_3765);
nand U8859 (N_8859,N_3870,N_2566);
or U8860 (N_8860,N_4910,N_2858);
nand U8861 (N_8861,N_1139,N_4545);
and U8862 (N_8862,N_1165,N_1072);
nor U8863 (N_8863,N_1343,N_4634);
nand U8864 (N_8864,N_4437,N_3726);
and U8865 (N_8865,N_2526,N_2152);
nor U8866 (N_8866,N_2413,N_3508);
or U8867 (N_8867,N_1536,N_1918);
and U8868 (N_8868,N_1661,N_762);
or U8869 (N_8869,N_1275,N_4354);
and U8870 (N_8870,N_2589,N_705);
and U8871 (N_8871,N_4002,N_4235);
xnor U8872 (N_8872,N_3637,N_2737);
and U8873 (N_8873,N_1701,N_4162);
nand U8874 (N_8874,N_3146,N_1610);
and U8875 (N_8875,N_3200,N_2717);
nor U8876 (N_8876,N_1805,N_3560);
nand U8877 (N_8877,N_2196,N_941);
or U8878 (N_8878,N_2766,N_1008);
and U8879 (N_8879,N_3399,N_2652);
nor U8880 (N_8880,N_2879,N_4263);
or U8881 (N_8881,N_3158,N_839);
or U8882 (N_8882,N_2058,N_4725);
nand U8883 (N_8883,N_536,N_1667);
nand U8884 (N_8884,N_1695,N_3084);
nand U8885 (N_8885,N_1192,N_306);
nand U8886 (N_8886,N_4144,N_4192);
and U8887 (N_8887,N_4160,N_1377);
nand U8888 (N_8888,N_1889,N_4868);
and U8889 (N_8889,N_41,N_3803);
or U8890 (N_8890,N_2117,N_4420);
or U8891 (N_8891,N_2684,N_2730);
or U8892 (N_8892,N_2583,N_2595);
nand U8893 (N_8893,N_704,N_1780);
or U8894 (N_8894,N_3790,N_656);
and U8895 (N_8895,N_4344,N_2798);
or U8896 (N_8896,N_4668,N_1092);
or U8897 (N_8897,N_388,N_3813);
and U8898 (N_8898,N_1061,N_3800);
nor U8899 (N_8899,N_1958,N_2719);
and U8900 (N_8900,N_2676,N_157);
xnor U8901 (N_8901,N_3700,N_4705);
and U8902 (N_8902,N_3954,N_2722);
or U8903 (N_8903,N_1016,N_4403);
nand U8904 (N_8904,N_3000,N_4858);
nand U8905 (N_8905,N_2289,N_4460);
nand U8906 (N_8906,N_1559,N_4250);
or U8907 (N_8907,N_3218,N_4084);
nand U8908 (N_8908,N_677,N_3685);
or U8909 (N_8909,N_915,N_2417);
nor U8910 (N_8910,N_4501,N_1933);
nand U8911 (N_8911,N_3726,N_1620);
and U8912 (N_8912,N_1053,N_814);
or U8913 (N_8913,N_1004,N_1405);
nand U8914 (N_8914,N_831,N_1023);
and U8915 (N_8915,N_3149,N_3729);
nand U8916 (N_8916,N_2817,N_2119);
nor U8917 (N_8917,N_2222,N_4659);
nand U8918 (N_8918,N_4051,N_2508);
or U8919 (N_8919,N_1823,N_1216);
or U8920 (N_8920,N_4494,N_1761);
nor U8921 (N_8921,N_4582,N_1426);
and U8922 (N_8922,N_2501,N_901);
nand U8923 (N_8923,N_577,N_1158);
nand U8924 (N_8924,N_1178,N_4516);
nor U8925 (N_8925,N_2835,N_3609);
nand U8926 (N_8926,N_2367,N_374);
nor U8927 (N_8927,N_4083,N_4792);
or U8928 (N_8928,N_4032,N_833);
or U8929 (N_8929,N_971,N_3652);
nor U8930 (N_8930,N_4242,N_4374);
and U8931 (N_8931,N_4081,N_1154);
and U8932 (N_8932,N_4627,N_2615);
or U8933 (N_8933,N_3353,N_4753);
or U8934 (N_8934,N_986,N_2805);
nand U8935 (N_8935,N_3530,N_4155);
nand U8936 (N_8936,N_4448,N_2190);
nand U8937 (N_8937,N_542,N_1690);
or U8938 (N_8938,N_4491,N_2843);
nor U8939 (N_8939,N_2693,N_4398);
or U8940 (N_8940,N_1305,N_3292);
nand U8941 (N_8941,N_1487,N_1628);
nand U8942 (N_8942,N_2661,N_320);
nand U8943 (N_8943,N_1341,N_3570);
or U8944 (N_8944,N_1885,N_2715);
and U8945 (N_8945,N_2749,N_2462);
or U8946 (N_8946,N_3621,N_3607);
and U8947 (N_8947,N_420,N_2681);
or U8948 (N_8948,N_3017,N_4281);
nand U8949 (N_8949,N_4549,N_2081);
nand U8950 (N_8950,N_2572,N_101);
nor U8951 (N_8951,N_997,N_2292);
nand U8952 (N_8952,N_306,N_2292);
and U8953 (N_8953,N_4616,N_3654);
or U8954 (N_8954,N_3804,N_4858);
nand U8955 (N_8955,N_3366,N_1076);
nor U8956 (N_8956,N_4651,N_2246);
nor U8957 (N_8957,N_2727,N_1440);
nor U8958 (N_8958,N_3730,N_278);
or U8959 (N_8959,N_2436,N_989);
nor U8960 (N_8960,N_844,N_4941);
xor U8961 (N_8961,N_1739,N_2002);
and U8962 (N_8962,N_2951,N_2854);
or U8963 (N_8963,N_2160,N_1723);
and U8964 (N_8964,N_1412,N_2856);
and U8965 (N_8965,N_3356,N_2355);
nor U8966 (N_8966,N_2912,N_456);
nor U8967 (N_8967,N_3101,N_2561);
nand U8968 (N_8968,N_1748,N_3079);
and U8969 (N_8969,N_2004,N_3025);
nor U8970 (N_8970,N_1623,N_4147);
nand U8971 (N_8971,N_2744,N_3625);
and U8972 (N_8972,N_455,N_925);
nand U8973 (N_8973,N_2767,N_2291);
or U8974 (N_8974,N_4936,N_4184);
nor U8975 (N_8975,N_4594,N_3619);
and U8976 (N_8976,N_1763,N_2246);
and U8977 (N_8977,N_2017,N_4572);
and U8978 (N_8978,N_1062,N_4578);
nand U8979 (N_8979,N_4722,N_1702);
or U8980 (N_8980,N_4586,N_339);
or U8981 (N_8981,N_690,N_139);
and U8982 (N_8982,N_4957,N_1985);
nor U8983 (N_8983,N_1575,N_4883);
nor U8984 (N_8984,N_1711,N_4667);
nor U8985 (N_8985,N_1242,N_2874);
nor U8986 (N_8986,N_3387,N_3433);
nand U8987 (N_8987,N_264,N_277);
nand U8988 (N_8988,N_2356,N_3653);
or U8989 (N_8989,N_417,N_3531);
nand U8990 (N_8990,N_3687,N_1166);
nor U8991 (N_8991,N_199,N_722);
or U8992 (N_8992,N_3026,N_4750);
nor U8993 (N_8993,N_1172,N_63);
or U8994 (N_8994,N_210,N_2701);
xnor U8995 (N_8995,N_472,N_3567);
nand U8996 (N_8996,N_2684,N_3629);
nor U8997 (N_8997,N_565,N_1807);
nand U8998 (N_8998,N_4774,N_4622);
nor U8999 (N_8999,N_456,N_3105);
nand U9000 (N_9000,N_328,N_4823);
and U9001 (N_9001,N_2892,N_4862);
nor U9002 (N_9002,N_4215,N_2359);
nand U9003 (N_9003,N_2464,N_3139);
nand U9004 (N_9004,N_1238,N_1154);
nand U9005 (N_9005,N_922,N_4476);
nand U9006 (N_9006,N_4535,N_4135);
nor U9007 (N_9007,N_2030,N_1937);
or U9008 (N_9008,N_3354,N_1387);
or U9009 (N_9009,N_431,N_2973);
nor U9010 (N_9010,N_31,N_3328);
nand U9011 (N_9011,N_1782,N_1051);
or U9012 (N_9012,N_2384,N_4818);
nor U9013 (N_9013,N_2323,N_2442);
xor U9014 (N_9014,N_3019,N_1418);
nand U9015 (N_9015,N_2493,N_4341);
nor U9016 (N_9016,N_2931,N_2654);
and U9017 (N_9017,N_2149,N_3486);
or U9018 (N_9018,N_1973,N_1483);
nor U9019 (N_9019,N_4754,N_3957);
nor U9020 (N_9020,N_4779,N_1445);
nor U9021 (N_9021,N_568,N_3315);
and U9022 (N_9022,N_3282,N_1636);
xor U9023 (N_9023,N_878,N_2225);
and U9024 (N_9024,N_3547,N_3916);
nand U9025 (N_9025,N_4105,N_608);
nor U9026 (N_9026,N_4350,N_2920);
nor U9027 (N_9027,N_3559,N_939);
or U9028 (N_9028,N_3920,N_1041);
and U9029 (N_9029,N_3550,N_1429);
or U9030 (N_9030,N_4124,N_374);
or U9031 (N_9031,N_558,N_2036);
xnor U9032 (N_9032,N_222,N_2557);
nand U9033 (N_9033,N_43,N_2807);
nand U9034 (N_9034,N_2766,N_2846);
nor U9035 (N_9035,N_334,N_123);
and U9036 (N_9036,N_3561,N_235);
or U9037 (N_9037,N_2208,N_3743);
and U9038 (N_9038,N_1901,N_2758);
or U9039 (N_9039,N_4836,N_910);
or U9040 (N_9040,N_2379,N_270);
and U9041 (N_9041,N_981,N_2543);
or U9042 (N_9042,N_2482,N_3829);
or U9043 (N_9043,N_3291,N_3732);
nand U9044 (N_9044,N_1944,N_3246);
nor U9045 (N_9045,N_454,N_2974);
nand U9046 (N_9046,N_941,N_4931);
or U9047 (N_9047,N_1460,N_2634);
nand U9048 (N_9048,N_1746,N_3204);
nor U9049 (N_9049,N_4846,N_1999);
nor U9050 (N_9050,N_1518,N_2478);
or U9051 (N_9051,N_2970,N_3879);
and U9052 (N_9052,N_2657,N_82);
xnor U9053 (N_9053,N_1244,N_389);
or U9054 (N_9054,N_4750,N_1469);
xnor U9055 (N_9055,N_4709,N_2761);
or U9056 (N_9056,N_599,N_1295);
nand U9057 (N_9057,N_2174,N_2501);
or U9058 (N_9058,N_2338,N_3700);
xor U9059 (N_9059,N_2839,N_4796);
nor U9060 (N_9060,N_2694,N_3278);
nor U9061 (N_9061,N_969,N_2274);
nor U9062 (N_9062,N_2968,N_240);
nor U9063 (N_9063,N_1854,N_935);
xnor U9064 (N_9064,N_417,N_3504);
nor U9065 (N_9065,N_303,N_3763);
xnor U9066 (N_9066,N_2043,N_1629);
or U9067 (N_9067,N_3382,N_3971);
nor U9068 (N_9068,N_3359,N_1966);
and U9069 (N_9069,N_2605,N_3881);
nand U9070 (N_9070,N_4687,N_2540);
and U9071 (N_9071,N_38,N_1462);
or U9072 (N_9072,N_331,N_3228);
or U9073 (N_9073,N_3728,N_4122);
xor U9074 (N_9074,N_3064,N_1626);
and U9075 (N_9075,N_1098,N_2518);
nand U9076 (N_9076,N_3068,N_1070);
nor U9077 (N_9077,N_2261,N_3243);
nor U9078 (N_9078,N_1915,N_4061);
xnor U9079 (N_9079,N_2848,N_2142);
and U9080 (N_9080,N_1419,N_1501);
nand U9081 (N_9081,N_4760,N_1015);
or U9082 (N_9082,N_983,N_3724);
xnor U9083 (N_9083,N_1966,N_2581);
or U9084 (N_9084,N_3284,N_2962);
nand U9085 (N_9085,N_322,N_2663);
nor U9086 (N_9086,N_3283,N_2539);
nor U9087 (N_9087,N_3777,N_1557);
nor U9088 (N_9088,N_576,N_1757);
nor U9089 (N_9089,N_685,N_2545);
nor U9090 (N_9090,N_1329,N_2541);
and U9091 (N_9091,N_776,N_772);
nor U9092 (N_9092,N_1641,N_4723);
and U9093 (N_9093,N_2224,N_2218);
or U9094 (N_9094,N_912,N_4677);
nand U9095 (N_9095,N_2315,N_4217);
nand U9096 (N_9096,N_1281,N_128);
nor U9097 (N_9097,N_1059,N_770);
nor U9098 (N_9098,N_3492,N_2990);
xnor U9099 (N_9099,N_3363,N_4220);
and U9100 (N_9100,N_155,N_2172);
xor U9101 (N_9101,N_1606,N_77);
or U9102 (N_9102,N_2823,N_1295);
nor U9103 (N_9103,N_2339,N_2675);
and U9104 (N_9104,N_2283,N_1764);
and U9105 (N_9105,N_1039,N_3646);
or U9106 (N_9106,N_1882,N_1054);
nand U9107 (N_9107,N_607,N_4940);
or U9108 (N_9108,N_3706,N_846);
nor U9109 (N_9109,N_3757,N_4454);
nor U9110 (N_9110,N_2318,N_11);
nand U9111 (N_9111,N_4952,N_535);
nand U9112 (N_9112,N_2525,N_1233);
nand U9113 (N_9113,N_3671,N_1580);
and U9114 (N_9114,N_4262,N_253);
nor U9115 (N_9115,N_1075,N_1131);
nor U9116 (N_9116,N_784,N_3488);
or U9117 (N_9117,N_882,N_1220);
nor U9118 (N_9118,N_1038,N_2871);
nand U9119 (N_9119,N_2713,N_3318);
or U9120 (N_9120,N_171,N_3283);
and U9121 (N_9121,N_3220,N_2748);
nand U9122 (N_9122,N_4314,N_202);
and U9123 (N_9123,N_2604,N_890);
or U9124 (N_9124,N_3817,N_471);
or U9125 (N_9125,N_414,N_2751);
xor U9126 (N_9126,N_879,N_3753);
nand U9127 (N_9127,N_3804,N_863);
and U9128 (N_9128,N_3753,N_4534);
and U9129 (N_9129,N_4572,N_4283);
and U9130 (N_9130,N_1458,N_2306);
or U9131 (N_9131,N_1144,N_4133);
and U9132 (N_9132,N_2161,N_4095);
and U9133 (N_9133,N_1227,N_2183);
nand U9134 (N_9134,N_2395,N_1796);
or U9135 (N_9135,N_3237,N_710);
nor U9136 (N_9136,N_2810,N_4253);
nand U9137 (N_9137,N_2054,N_3857);
or U9138 (N_9138,N_3056,N_4755);
nand U9139 (N_9139,N_4870,N_1675);
and U9140 (N_9140,N_269,N_4521);
and U9141 (N_9141,N_3487,N_2617);
nand U9142 (N_9142,N_2016,N_1873);
and U9143 (N_9143,N_3438,N_4592);
nor U9144 (N_9144,N_4284,N_3366);
nand U9145 (N_9145,N_812,N_1910);
and U9146 (N_9146,N_3652,N_2852);
nand U9147 (N_9147,N_569,N_3473);
or U9148 (N_9148,N_1024,N_1525);
nand U9149 (N_9149,N_1577,N_981);
nor U9150 (N_9150,N_2445,N_1330);
or U9151 (N_9151,N_47,N_2673);
and U9152 (N_9152,N_999,N_2568);
or U9153 (N_9153,N_289,N_2313);
xor U9154 (N_9154,N_3278,N_3575);
and U9155 (N_9155,N_3163,N_3743);
or U9156 (N_9156,N_4958,N_2104);
xnor U9157 (N_9157,N_291,N_1614);
or U9158 (N_9158,N_4703,N_1768);
and U9159 (N_9159,N_1419,N_2021);
nand U9160 (N_9160,N_3291,N_4355);
and U9161 (N_9161,N_1107,N_3904);
or U9162 (N_9162,N_3813,N_3521);
nor U9163 (N_9163,N_277,N_541);
or U9164 (N_9164,N_2409,N_1033);
nand U9165 (N_9165,N_3282,N_1977);
nor U9166 (N_9166,N_1235,N_3632);
or U9167 (N_9167,N_3868,N_4311);
nor U9168 (N_9168,N_4331,N_1615);
nand U9169 (N_9169,N_3448,N_3172);
and U9170 (N_9170,N_2340,N_4192);
nand U9171 (N_9171,N_3216,N_3056);
nor U9172 (N_9172,N_1229,N_195);
nor U9173 (N_9173,N_4396,N_3907);
nand U9174 (N_9174,N_858,N_15);
or U9175 (N_9175,N_3366,N_3044);
or U9176 (N_9176,N_3726,N_3007);
xnor U9177 (N_9177,N_2642,N_4809);
or U9178 (N_9178,N_3799,N_2442);
and U9179 (N_9179,N_325,N_1876);
nor U9180 (N_9180,N_4368,N_3671);
nor U9181 (N_9181,N_2327,N_614);
nor U9182 (N_9182,N_2350,N_3378);
nand U9183 (N_9183,N_3003,N_1507);
nor U9184 (N_9184,N_2777,N_3263);
or U9185 (N_9185,N_140,N_1331);
and U9186 (N_9186,N_3225,N_856);
nor U9187 (N_9187,N_3462,N_4346);
and U9188 (N_9188,N_4666,N_3442);
nor U9189 (N_9189,N_805,N_221);
nor U9190 (N_9190,N_4250,N_1295);
nand U9191 (N_9191,N_136,N_1561);
or U9192 (N_9192,N_1575,N_1882);
and U9193 (N_9193,N_1093,N_3381);
nor U9194 (N_9194,N_3900,N_1371);
and U9195 (N_9195,N_4050,N_4614);
nor U9196 (N_9196,N_3956,N_2054);
or U9197 (N_9197,N_4217,N_2603);
nand U9198 (N_9198,N_464,N_2090);
nand U9199 (N_9199,N_4855,N_3678);
nor U9200 (N_9200,N_2407,N_3542);
nor U9201 (N_9201,N_2995,N_3476);
nand U9202 (N_9202,N_1760,N_763);
nand U9203 (N_9203,N_2277,N_2918);
and U9204 (N_9204,N_3130,N_1040);
nand U9205 (N_9205,N_3341,N_999);
nand U9206 (N_9206,N_2730,N_1542);
nor U9207 (N_9207,N_1242,N_4179);
nor U9208 (N_9208,N_1490,N_738);
or U9209 (N_9209,N_3226,N_2743);
and U9210 (N_9210,N_4147,N_4613);
nor U9211 (N_9211,N_451,N_831);
xor U9212 (N_9212,N_2792,N_769);
or U9213 (N_9213,N_1340,N_1558);
and U9214 (N_9214,N_4593,N_4057);
or U9215 (N_9215,N_2229,N_3676);
nor U9216 (N_9216,N_3719,N_3200);
or U9217 (N_9217,N_385,N_4284);
xnor U9218 (N_9218,N_1219,N_895);
nor U9219 (N_9219,N_1435,N_4773);
nor U9220 (N_9220,N_361,N_2105);
and U9221 (N_9221,N_1460,N_3281);
nand U9222 (N_9222,N_1819,N_4350);
or U9223 (N_9223,N_2893,N_3234);
and U9224 (N_9224,N_2033,N_146);
nor U9225 (N_9225,N_1477,N_1165);
and U9226 (N_9226,N_4785,N_4983);
xor U9227 (N_9227,N_902,N_982);
nand U9228 (N_9228,N_2826,N_175);
or U9229 (N_9229,N_1263,N_3752);
nand U9230 (N_9230,N_4171,N_4941);
nor U9231 (N_9231,N_3699,N_1225);
nor U9232 (N_9232,N_534,N_4989);
nor U9233 (N_9233,N_1042,N_3136);
and U9234 (N_9234,N_2811,N_1077);
and U9235 (N_9235,N_4340,N_3469);
or U9236 (N_9236,N_161,N_4857);
and U9237 (N_9237,N_4558,N_4582);
or U9238 (N_9238,N_168,N_4912);
nand U9239 (N_9239,N_74,N_3197);
nand U9240 (N_9240,N_2119,N_1110);
or U9241 (N_9241,N_4379,N_4171);
nor U9242 (N_9242,N_4946,N_2610);
nand U9243 (N_9243,N_2456,N_3336);
nand U9244 (N_9244,N_2968,N_4026);
and U9245 (N_9245,N_862,N_2318);
and U9246 (N_9246,N_1403,N_4506);
nand U9247 (N_9247,N_1256,N_2685);
nor U9248 (N_9248,N_4181,N_270);
or U9249 (N_9249,N_1532,N_3774);
and U9250 (N_9250,N_2151,N_645);
nand U9251 (N_9251,N_1111,N_49);
or U9252 (N_9252,N_109,N_4233);
nor U9253 (N_9253,N_3068,N_4559);
nor U9254 (N_9254,N_1589,N_1050);
nor U9255 (N_9255,N_4488,N_4648);
and U9256 (N_9256,N_563,N_3163);
or U9257 (N_9257,N_2976,N_4620);
nor U9258 (N_9258,N_2266,N_1397);
nand U9259 (N_9259,N_3471,N_1855);
or U9260 (N_9260,N_3520,N_44);
nor U9261 (N_9261,N_2935,N_1817);
nor U9262 (N_9262,N_1803,N_369);
and U9263 (N_9263,N_929,N_742);
nand U9264 (N_9264,N_4402,N_3183);
or U9265 (N_9265,N_1110,N_4228);
and U9266 (N_9266,N_4189,N_2991);
nor U9267 (N_9267,N_867,N_4858);
or U9268 (N_9268,N_533,N_2831);
or U9269 (N_9269,N_233,N_2053);
xnor U9270 (N_9270,N_134,N_2355);
or U9271 (N_9271,N_564,N_556);
nor U9272 (N_9272,N_773,N_1803);
nand U9273 (N_9273,N_1328,N_3205);
nand U9274 (N_9274,N_4119,N_4351);
nor U9275 (N_9275,N_1279,N_4750);
nand U9276 (N_9276,N_1135,N_2495);
nor U9277 (N_9277,N_4555,N_2660);
nor U9278 (N_9278,N_201,N_1735);
or U9279 (N_9279,N_979,N_110);
or U9280 (N_9280,N_4140,N_4462);
and U9281 (N_9281,N_3296,N_453);
or U9282 (N_9282,N_2250,N_3662);
nor U9283 (N_9283,N_2895,N_8);
nor U9284 (N_9284,N_2988,N_4759);
nor U9285 (N_9285,N_1674,N_2737);
nor U9286 (N_9286,N_1186,N_3442);
or U9287 (N_9287,N_1904,N_3329);
nand U9288 (N_9288,N_2943,N_2531);
and U9289 (N_9289,N_1589,N_1885);
and U9290 (N_9290,N_2112,N_3997);
or U9291 (N_9291,N_3471,N_1713);
nor U9292 (N_9292,N_2787,N_2282);
nand U9293 (N_9293,N_1595,N_2302);
or U9294 (N_9294,N_3261,N_149);
nand U9295 (N_9295,N_3433,N_216);
nand U9296 (N_9296,N_2409,N_2312);
and U9297 (N_9297,N_1777,N_205);
or U9298 (N_9298,N_1018,N_2417);
nand U9299 (N_9299,N_3671,N_2822);
nand U9300 (N_9300,N_4393,N_1929);
or U9301 (N_9301,N_3307,N_4510);
or U9302 (N_9302,N_830,N_59);
nor U9303 (N_9303,N_2083,N_3236);
and U9304 (N_9304,N_4825,N_1169);
nor U9305 (N_9305,N_4395,N_423);
nor U9306 (N_9306,N_3216,N_2785);
nor U9307 (N_9307,N_3954,N_3226);
or U9308 (N_9308,N_3637,N_2752);
nor U9309 (N_9309,N_3040,N_423);
nor U9310 (N_9310,N_4049,N_1626);
nand U9311 (N_9311,N_3286,N_3344);
or U9312 (N_9312,N_3104,N_3122);
nor U9313 (N_9313,N_3292,N_4467);
and U9314 (N_9314,N_262,N_1110);
and U9315 (N_9315,N_858,N_3576);
nor U9316 (N_9316,N_4105,N_539);
and U9317 (N_9317,N_1621,N_2323);
or U9318 (N_9318,N_4820,N_2633);
nand U9319 (N_9319,N_2119,N_3261);
nand U9320 (N_9320,N_4119,N_4469);
or U9321 (N_9321,N_4900,N_2886);
or U9322 (N_9322,N_4663,N_1726);
nor U9323 (N_9323,N_918,N_4265);
nand U9324 (N_9324,N_919,N_3816);
nand U9325 (N_9325,N_2717,N_1175);
nand U9326 (N_9326,N_3945,N_3295);
nor U9327 (N_9327,N_143,N_4679);
nor U9328 (N_9328,N_2022,N_3642);
or U9329 (N_9329,N_4335,N_4594);
or U9330 (N_9330,N_653,N_657);
or U9331 (N_9331,N_4571,N_2255);
nor U9332 (N_9332,N_4889,N_1422);
nand U9333 (N_9333,N_4581,N_4295);
nor U9334 (N_9334,N_788,N_1823);
or U9335 (N_9335,N_795,N_3550);
or U9336 (N_9336,N_87,N_3070);
or U9337 (N_9337,N_2263,N_2549);
nand U9338 (N_9338,N_3996,N_4923);
and U9339 (N_9339,N_1902,N_2644);
nor U9340 (N_9340,N_4223,N_3109);
nand U9341 (N_9341,N_3880,N_377);
or U9342 (N_9342,N_1767,N_4422);
nand U9343 (N_9343,N_3925,N_133);
nor U9344 (N_9344,N_2721,N_3834);
nand U9345 (N_9345,N_382,N_1217);
and U9346 (N_9346,N_4780,N_2456);
nor U9347 (N_9347,N_1150,N_1966);
and U9348 (N_9348,N_2770,N_2419);
and U9349 (N_9349,N_4609,N_4405);
and U9350 (N_9350,N_2790,N_3879);
or U9351 (N_9351,N_4539,N_3266);
and U9352 (N_9352,N_544,N_353);
or U9353 (N_9353,N_3416,N_1856);
nand U9354 (N_9354,N_2919,N_329);
or U9355 (N_9355,N_2910,N_1023);
and U9356 (N_9356,N_143,N_1649);
or U9357 (N_9357,N_3515,N_2399);
nand U9358 (N_9358,N_4340,N_2504);
nand U9359 (N_9359,N_2605,N_1495);
or U9360 (N_9360,N_4389,N_4544);
nor U9361 (N_9361,N_3190,N_1952);
and U9362 (N_9362,N_2548,N_1892);
nand U9363 (N_9363,N_805,N_4775);
xor U9364 (N_9364,N_219,N_1727);
and U9365 (N_9365,N_2871,N_3306);
and U9366 (N_9366,N_271,N_503);
nand U9367 (N_9367,N_3906,N_1468);
nand U9368 (N_9368,N_3366,N_1603);
xor U9369 (N_9369,N_1350,N_1450);
nand U9370 (N_9370,N_1940,N_967);
and U9371 (N_9371,N_2947,N_36);
nand U9372 (N_9372,N_4525,N_4607);
or U9373 (N_9373,N_2278,N_2257);
or U9374 (N_9374,N_766,N_322);
nand U9375 (N_9375,N_4763,N_4874);
nor U9376 (N_9376,N_542,N_3847);
or U9377 (N_9377,N_190,N_2082);
xor U9378 (N_9378,N_2623,N_727);
and U9379 (N_9379,N_3748,N_1568);
nor U9380 (N_9380,N_3496,N_3545);
or U9381 (N_9381,N_3732,N_1224);
nor U9382 (N_9382,N_2304,N_2198);
or U9383 (N_9383,N_1270,N_1754);
and U9384 (N_9384,N_3751,N_234);
and U9385 (N_9385,N_2089,N_57);
and U9386 (N_9386,N_2777,N_3201);
and U9387 (N_9387,N_1162,N_2123);
or U9388 (N_9388,N_662,N_4789);
nor U9389 (N_9389,N_4533,N_4072);
or U9390 (N_9390,N_4326,N_810);
and U9391 (N_9391,N_3669,N_4977);
or U9392 (N_9392,N_3707,N_4315);
nand U9393 (N_9393,N_4288,N_2368);
or U9394 (N_9394,N_221,N_4690);
nor U9395 (N_9395,N_3286,N_1391);
nor U9396 (N_9396,N_2039,N_4216);
nand U9397 (N_9397,N_1593,N_3939);
or U9398 (N_9398,N_4525,N_4033);
and U9399 (N_9399,N_1785,N_3382);
or U9400 (N_9400,N_3305,N_3241);
nand U9401 (N_9401,N_4359,N_2831);
and U9402 (N_9402,N_3707,N_1874);
nand U9403 (N_9403,N_2332,N_4040);
and U9404 (N_9404,N_3215,N_269);
nor U9405 (N_9405,N_275,N_72);
nor U9406 (N_9406,N_4168,N_1466);
nor U9407 (N_9407,N_1537,N_4937);
nor U9408 (N_9408,N_3046,N_3307);
nand U9409 (N_9409,N_3726,N_4859);
and U9410 (N_9410,N_3666,N_157);
or U9411 (N_9411,N_4393,N_986);
and U9412 (N_9412,N_1306,N_602);
and U9413 (N_9413,N_2761,N_1669);
nand U9414 (N_9414,N_4524,N_2894);
nor U9415 (N_9415,N_679,N_3811);
nand U9416 (N_9416,N_149,N_1889);
or U9417 (N_9417,N_972,N_2688);
or U9418 (N_9418,N_136,N_177);
or U9419 (N_9419,N_431,N_4947);
nor U9420 (N_9420,N_2426,N_3189);
or U9421 (N_9421,N_4906,N_1406);
and U9422 (N_9422,N_257,N_3821);
and U9423 (N_9423,N_3209,N_669);
or U9424 (N_9424,N_1816,N_4045);
or U9425 (N_9425,N_3917,N_3051);
or U9426 (N_9426,N_1420,N_1195);
nand U9427 (N_9427,N_4227,N_4817);
and U9428 (N_9428,N_886,N_2621);
and U9429 (N_9429,N_4939,N_3856);
and U9430 (N_9430,N_252,N_541);
or U9431 (N_9431,N_1091,N_4316);
nand U9432 (N_9432,N_4603,N_4739);
and U9433 (N_9433,N_4612,N_1636);
nor U9434 (N_9434,N_4993,N_2265);
or U9435 (N_9435,N_2119,N_1962);
or U9436 (N_9436,N_394,N_2631);
and U9437 (N_9437,N_3626,N_2637);
xnor U9438 (N_9438,N_454,N_2952);
or U9439 (N_9439,N_2727,N_3075);
or U9440 (N_9440,N_3524,N_3910);
or U9441 (N_9441,N_3097,N_4817);
nor U9442 (N_9442,N_3376,N_2326);
nand U9443 (N_9443,N_1208,N_1028);
and U9444 (N_9444,N_2585,N_3844);
or U9445 (N_9445,N_4242,N_319);
and U9446 (N_9446,N_4938,N_124);
or U9447 (N_9447,N_206,N_1886);
and U9448 (N_9448,N_4582,N_3921);
nor U9449 (N_9449,N_41,N_830);
or U9450 (N_9450,N_3321,N_2476);
nor U9451 (N_9451,N_4025,N_2607);
nor U9452 (N_9452,N_3121,N_1713);
nand U9453 (N_9453,N_3538,N_2906);
nand U9454 (N_9454,N_4499,N_3411);
or U9455 (N_9455,N_4616,N_3126);
or U9456 (N_9456,N_4058,N_1827);
and U9457 (N_9457,N_2345,N_4422);
nand U9458 (N_9458,N_2066,N_761);
or U9459 (N_9459,N_4469,N_2308);
xnor U9460 (N_9460,N_3495,N_4428);
nand U9461 (N_9461,N_3901,N_4433);
or U9462 (N_9462,N_4660,N_4212);
or U9463 (N_9463,N_134,N_3329);
nand U9464 (N_9464,N_2772,N_4024);
or U9465 (N_9465,N_322,N_2566);
nor U9466 (N_9466,N_2947,N_2898);
nand U9467 (N_9467,N_2833,N_1779);
or U9468 (N_9468,N_973,N_3457);
nor U9469 (N_9469,N_2891,N_3332);
xor U9470 (N_9470,N_3380,N_3000);
or U9471 (N_9471,N_1266,N_4534);
xnor U9472 (N_9472,N_2621,N_2926);
nand U9473 (N_9473,N_2197,N_2089);
and U9474 (N_9474,N_1935,N_3488);
or U9475 (N_9475,N_148,N_1502);
nand U9476 (N_9476,N_4605,N_1981);
nor U9477 (N_9477,N_2019,N_4617);
nor U9478 (N_9478,N_6,N_2197);
or U9479 (N_9479,N_3361,N_2088);
and U9480 (N_9480,N_4838,N_4872);
nor U9481 (N_9481,N_4673,N_1396);
nand U9482 (N_9482,N_3282,N_954);
nor U9483 (N_9483,N_4988,N_1109);
and U9484 (N_9484,N_841,N_1898);
and U9485 (N_9485,N_1572,N_2517);
and U9486 (N_9486,N_2506,N_3712);
and U9487 (N_9487,N_3551,N_4563);
or U9488 (N_9488,N_207,N_3307);
nand U9489 (N_9489,N_2437,N_2969);
nand U9490 (N_9490,N_3214,N_3835);
and U9491 (N_9491,N_4827,N_3701);
and U9492 (N_9492,N_3301,N_1511);
xor U9493 (N_9493,N_1578,N_3173);
and U9494 (N_9494,N_3145,N_1267);
nor U9495 (N_9495,N_2902,N_2006);
or U9496 (N_9496,N_3765,N_4280);
nor U9497 (N_9497,N_149,N_2230);
and U9498 (N_9498,N_2255,N_4276);
or U9499 (N_9499,N_751,N_1097);
and U9500 (N_9500,N_2899,N_3271);
nand U9501 (N_9501,N_2617,N_4400);
and U9502 (N_9502,N_1996,N_4584);
nor U9503 (N_9503,N_3686,N_1256);
nand U9504 (N_9504,N_1640,N_661);
nor U9505 (N_9505,N_4345,N_1277);
or U9506 (N_9506,N_1595,N_4282);
nand U9507 (N_9507,N_1152,N_940);
nor U9508 (N_9508,N_3192,N_2900);
and U9509 (N_9509,N_3700,N_758);
nand U9510 (N_9510,N_4590,N_4850);
and U9511 (N_9511,N_367,N_275);
nand U9512 (N_9512,N_577,N_3621);
nor U9513 (N_9513,N_1379,N_1417);
nor U9514 (N_9514,N_4245,N_4282);
nor U9515 (N_9515,N_4940,N_1446);
nand U9516 (N_9516,N_3905,N_1137);
and U9517 (N_9517,N_4049,N_1326);
and U9518 (N_9518,N_3862,N_3618);
nor U9519 (N_9519,N_338,N_3303);
nand U9520 (N_9520,N_2734,N_586);
and U9521 (N_9521,N_274,N_4211);
nand U9522 (N_9522,N_2183,N_2880);
nor U9523 (N_9523,N_3292,N_585);
or U9524 (N_9524,N_1581,N_2732);
nand U9525 (N_9525,N_3910,N_465);
nand U9526 (N_9526,N_1384,N_1849);
or U9527 (N_9527,N_2252,N_970);
and U9528 (N_9528,N_3272,N_2169);
nor U9529 (N_9529,N_3065,N_1818);
and U9530 (N_9530,N_4745,N_2585);
or U9531 (N_9531,N_1938,N_3687);
or U9532 (N_9532,N_1101,N_491);
or U9533 (N_9533,N_2234,N_204);
nor U9534 (N_9534,N_4550,N_718);
nand U9535 (N_9535,N_393,N_3619);
and U9536 (N_9536,N_3804,N_1212);
and U9537 (N_9537,N_2163,N_3345);
or U9538 (N_9538,N_1281,N_4428);
nand U9539 (N_9539,N_4685,N_3232);
nor U9540 (N_9540,N_4233,N_1255);
or U9541 (N_9541,N_3969,N_4125);
nor U9542 (N_9542,N_3479,N_27);
and U9543 (N_9543,N_1037,N_410);
nand U9544 (N_9544,N_4772,N_1300);
nor U9545 (N_9545,N_3003,N_137);
or U9546 (N_9546,N_4276,N_4134);
nor U9547 (N_9547,N_153,N_4022);
nand U9548 (N_9548,N_2062,N_2644);
and U9549 (N_9549,N_184,N_4986);
nand U9550 (N_9550,N_957,N_4749);
nand U9551 (N_9551,N_1932,N_3571);
nand U9552 (N_9552,N_4231,N_1176);
nor U9553 (N_9553,N_3765,N_1197);
and U9554 (N_9554,N_3071,N_3663);
nand U9555 (N_9555,N_116,N_506);
or U9556 (N_9556,N_3541,N_127);
nand U9557 (N_9557,N_1981,N_4773);
nand U9558 (N_9558,N_4037,N_3826);
nor U9559 (N_9559,N_2629,N_1953);
and U9560 (N_9560,N_3680,N_1071);
nor U9561 (N_9561,N_1942,N_3751);
nor U9562 (N_9562,N_4106,N_2493);
nor U9563 (N_9563,N_2456,N_3020);
nand U9564 (N_9564,N_4416,N_3353);
and U9565 (N_9565,N_4292,N_840);
and U9566 (N_9566,N_1084,N_1696);
nor U9567 (N_9567,N_787,N_3744);
nor U9568 (N_9568,N_407,N_3206);
nand U9569 (N_9569,N_141,N_4194);
or U9570 (N_9570,N_1639,N_19);
nand U9571 (N_9571,N_4108,N_3208);
nand U9572 (N_9572,N_3249,N_549);
nand U9573 (N_9573,N_1254,N_385);
and U9574 (N_9574,N_3182,N_3846);
nand U9575 (N_9575,N_177,N_4188);
or U9576 (N_9576,N_2893,N_1131);
nand U9577 (N_9577,N_4771,N_1374);
nand U9578 (N_9578,N_1002,N_832);
nand U9579 (N_9579,N_2535,N_647);
nand U9580 (N_9580,N_2885,N_3406);
nor U9581 (N_9581,N_1706,N_1718);
nand U9582 (N_9582,N_1508,N_2302);
and U9583 (N_9583,N_3937,N_4557);
or U9584 (N_9584,N_2845,N_3866);
or U9585 (N_9585,N_4560,N_1324);
xor U9586 (N_9586,N_1000,N_1983);
nand U9587 (N_9587,N_2122,N_4294);
and U9588 (N_9588,N_3053,N_2738);
nand U9589 (N_9589,N_3353,N_732);
or U9590 (N_9590,N_2715,N_2439);
or U9591 (N_9591,N_1628,N_3106);
and U9592 (N_9592,N_2466,N_632);
or U9593 (N_9593,N_1242,N_4655);
nand U9594 (N_9594,N_2383,N_4548);
or U9595 (N_9595,N_3529,N_3708);
nor U9596 (N_9596,N_306,N_45);
nand U9597 (N_9597,N_1395,N_596);
nand U9598 (N_9598,N_3000,N_1616);
nand U9599 (N_9599,N_3000,N_3483);
and U9600 (N_9600,N_2456,N_499);
and U9601 (N_9601,N_2544,N_1179);
nor U9602 (N_9602,N_4017,N_466);
nand U9603 (N_9603,N_3286,N_465);
nand U9604 (N_9604,N_503,N_1609);
or U9605 (N_9605,N_2927,N_954);
and U9606 (N_9606,N_427,N_462);
nor U9607 (N_9607,N_3623,N_3574);
and U9608 (N_9608,N_1351,N_3905);
nand U9609 (N_9609,N_4675,N_2794);
and U9610 (N_9610,N_3225,N_353);
nand U9611 (N_9611,N_996,N_1294);
nand U9612 (N_9612,N_752,N_3533);
nor U9613 (N_9613,N_1582,N_1685);
nor U9614 (N_9614,N_4756,N_3925);
nand U9615 (N_9615,N_4132,N_996);
nor U9616 (N_9616,N_3706,N_855);
nand U9617 (N_9617,N_2574,N_3144);
nor U9618 (N_9618,N_2498,N_4496);
and U9619 (N_9619,N_1064,N_3597);
nor U9620 (N_9620,N_488,N_2229);
or U9621 (N_9621,N_811,N_89);
and U9622 (N_9622,N_3487,N_1979);
or U9623 (N_9623,N_1095,N_3682);
nor U9624 (N_9624,N_3780,N_234);
or U9625 (N_9625,N_1221,N_3359);
nor U9626 (N_9626,N_1609,N_922);
nor U9627 (N_9627,N_949,N_1402);
nand U9628 (N_9628,N_2344,N_2614);
or U9629 (N_9629,N_1254,N_2961);
and U9630 (N_9630,N_937,N_2492);
and U9631 (N_9631,N_358,N_125);
nor U9632 (N_9632,N_2578,N_47);
nand U9633 (N_9633,N_1291,N_599);
nand U9634 (N_9634,N_751,N_4761);
nor U9635 (N_9635,N_4520,N_1737);
and U9636 (N_9636,N_118,N_2877);
nor U9637 (N_9637,N_2000,N_1334);
nand U9638 (N_9638,N_3022,N_4746);
xnor U9639 (N_9639,N_4072,N_2328);
and U9640 (N_9640,N_4174,N_2280);
nor U9641 (N_9641,N_4490,N_1603);
xnor U9642 (N_9642,N_4713,N_348);
or U9643 (N_9643,N_32,N_2033);
and U9644 (N_9644,N_3768,N_3248);
xor U9645 (N_9645,N_514,N_2145);
nor U9646 (N_9646,N_4142,N_3105);
nor U9647 (N_9647,N_1111,N_2009);
nand U9648 (N_9648,N_3252,N_4336);
nand U9649 (N_9649,N_4652,N_856);
xnor U9650 (N_9650,N_854,N_4572);
or U9651 (N_9651,N_1204,N_3723);
or U9652 (N_9652,N_2063,N_4969);
and U9653 (N_9653,N_4621,N_4175);
or U9654 (N_9654,N_2833,N_2);
and U9655 (N_9655,N_4737,N_1124);
nand U9656 (N_9656,N_1714,N_2999);
xor U9657 (N_9657,N_770,N_2918);
nor U9658 (N_9658,N_1980,N_4449);
nor U9659 (N_9659,N_4554,N_2434);
or U9660 (N_9660,N_0,N_4295);
nand U9661 (N_9661,N_3577,N_1670);
or U9662 (N_9662,N_4015,N_1846);
and U9663 (N_9663,N_3779,N_4298);
nand U9664 (N_9664,N_766,N_769);
or U9665 (N_9665,N_1856,N_2647);
and U9666 (N_9666,N_3729,N_12);
xor U9667 (N_9667,N_3405,N_2829);
nand U9668 (N_9668,N_346,N_2918);
or U9669 (N_9669,N_4653,N_2073);
or U9670 (N_9670,N_3349,N_1197);
nand U9671 (N_9671,N_3017,N_773);
and U9672 (N_9672,N_4351,N_3946);
nor U9673 (N_9673,N_2645,N_1709);
nand U9674 (N_9674,N_4194,N_1706);
nor U9675 (N_9675,N_2794,N_2138);
or U9676 (N_9676,N_3059,N_1787);
and U9677 (N_9677,N_2510,N_3086);
nor U9678 (N_9678,N_1045,N_3476);
nand U9679 (N_9679,N_2262,N_4499);
nor U9680 (N_9680,N_2161,N_4785);
nor U9681 (N_9681,N_4903,N_77);
and U9682 (N_9682,N_2597,N_3950);
or U9683 (N_9683,N_1317,N_4286);
and U9684 (N_9684,N_3116,N_4587);
and U9685 (N_9685,N_3507,N_1326);
and U9686 (N_9686,N_1526,N_3735);
nand U9687 (N_9687,N_3058,N_1109);
and U9688 (N_9688,N_2311,N_4521);
or U9689 (N_9689,N_361,N_3717);
nand U9690 (N_9690,N_746,N_2191);
nand U9691 (N_9691,N_4875,N_1907);
and U9692 (N_9692,N_4080,N_2258);
nand U9693 (N_9693,N_4410,N_3803);
nor U9694 (N_9694,N_3292,N_1007);
and U9695 (N_9695,N_4619,N_656);
nor U9696 (N_9696,N_526,N_4779);
or U9697 (N_9697,N_1485,N_1530);
or U9698 (N_9698,N_2108,N_46);
nor U9699 (N_9699,N_4930,N_2111);
nand U9700 (N_9700,N_1569,N_3998);
xnor U9701 (N_9701,N_914,N_2954);
nand U9702 (N_9702,N_87,N_2725);
or U9703 (N_9703,N_1304,N_425);
nand U9704 (N_9704,N_591,N_4590);
or U9705 (N_9705,N_1822,N_552);
and U9706 (N_9706,N_1593,N_863);
xor U9707 (N_9707,N_2353,N_974);
nor U9708 (N_9708,N_1169,N_760);
nor U9709 (N_9709,N_2758,N_2458);
and U9710 (N_9710,N_2636,N_1799);
and U9711 (N_9711,N_847,N_1601);
nand U9712 (N_9712,N_4205,N_1460);
nand U9713 (N_9713,N_276,N_735);
and U9714 (N_9714,N_3642,N_3106);
or U9715 (N_9715,N_145,N_2852);
nand U9716 (N_9716,N_4320,N_481);
nor U9717 (N_9717,N_4837,N_2646);
or U9718 (N_9718,N_3,N_4168);
nor U9719 (N_9719,N_2186,N_1366);
nor U9720 (N_9720,N_1788,N_1407);
or U9721 (N_9721,N_4339,N_2668);
nor U9722 (N_9722,N_656,N_2975);
and U9723 (N_9723,N_2493,N_3009);
or U9724 (N_9724,N_2643,N_4097);
nand U9725 (N_9725,N_2639,N_655);
and U9726 (N_9726,N_3992,N_2454);
nand U9727 (N_9727,N_1338,N_2067);
nand U9728 (N_9728,N_4453,N_2957);
nand U9729 (N_9729,N_4013,N_4893);
nor U9730 (N_9730,N_1170,N_4811);
nor U9731 (N_9731,N_182,N_4014);
nand U9732 (N_9732,N_3429,N_1562);
nor U9733 (N_9733,N_4589,N_1657);
or U9734 (N_9734,N_2561,N_605);
nand U9735 (N_9735,N_691,N_2138);
nor U9736 (N_9736,N_70,N_3430);
nor U9737 (N_9737,N_1347,N_2317);
nor U9738 (N_9738,N_1431,N_1682);
and U9739 (N_9739,N_4904,N_203);
and U9740 (N_9740,N_1247,N_148);
nand U9741 (N_9741,N_1247,N_2981);
and U9742 (N_9742,N_2243,N_550);
nand U9743 (N_9743,N_2787,N_285);
or U9744 (N_9744,N_3470,N_3760);
or U9745 (N_9745,N_592,N_4496);
or U9746 (N_9746,N_2048,N_2117);
nor U9747 (N_9747,N_264,N_1346);
and U9748 (N_9748,N_684,N_2134);
and U9749 (N_9749,N_3985,N_4486);
nand U9750 (N_9750,N_3650,N_556);
nand U9751 (N_9751,N_3134,N_1797);
nand U9752 (N_9752,N_189,N_2763);
nor U9753 (N_9753,N_1270,N_2783);
xnor U9754 (N_9754,N_4035,N_308);
and U9755 (N_9755,N_2268,N_3866);
and U9756 (N_9756,N_2703,N_4717);
or U9757 (N_9757,N_701,N_4404);
or U9758 (N_9758,N_1468,N_962);
nor U9759 (N_9759,N_111,N_278);
nand U9760 (N_9760,N_3131,N_4038);
and U9761 (N_9761,N_3120,N_4686);
or U9762 (N_9762,N_0,N_720);
nand U9763 (N_9763,N_3624,N_3388);
or U9764 (N_9764,N_765,N_4058);
or U9765 (N_9765,N_1652,N_4947);
nor U9766 (N_9766,N_2143,N_3138);
nor U9767 (N_9767,N_40,N_1779);
and U9768 (N_9768,N_1025,N_4754);
or U9769 (N_9769,N_1758,N_3040);
nor U9770 (N_9770,N_2857,N_32);
and U9771 (N_9771,N_164,N_2728);
nor U9772 (N_9772,N_1366,N_4476);
nand U9773 (N_9773,N_2047,N_4260);
nor U9774 (N_9774,N_4345,N_2701);
or U9775 (N_9775,N_1238,N_1006);
nor U9776 (N_9776,N_4531,N_2571);
or U9777 (N_9777,N_739,N_737);
and U9778 (N_9778,N_588,N_1873);
or U9779 (N_9779,N_1403,N_886);
nor U9780 (N_9780,N_4846,N_4702);
nor U9781 (N_9781,N_4828,N_1011);
nor U9782 (N_9782,N_3591,N_2064);
and U9783 (N_9783,N_4688,N_568);
or U9784 (N_9784,N_2991,N_4806);
or U9785 (N_9785,N_726,N_366);
and U9786 (N_9786,N_2546,N_1900);
nor U9787 (N_9787,N_437,N_4768);
or U9788 (N_9788,N_4670,N_3728);
nor U9789 (N_9789,N_308,N_4324);
or U9790 (N_9790,N_4617,N_4191);
and U9791 (N_9791,N_2811,N_2957);
nor U9792 (N_9792,N_585,N_438);
and U9793 (N_9793,N_1029,N_3311);
nor U9794 (N_9794,N_1525,N_2624);
nor U9795 (N_9795,N_1839,N_1764);
nor U9796 (N_9796,N_2964,N_4157);
nor U9797 (N_9797,N_3201,N_4596);
or U9798 (N_9798,N_3505,N_3530);
or U9799 (N_9799,N_2441,N_166);
nor U9800 (N_9800,N_503,N_4891);
or U9801 (N_9801,N_1437,N_1127);
nand U9802 (N_9802,N_2503,N_811);
nor U9803 (N_9803,N_4028,N_459);
nor U9804 (N_9804,N_1833,N_2042);
nor U9805 (N_9805,N_3426,N_3207);
and U9806 (N_9806,N_718,N_4411);
and U9807 (N_9807,N_1287,N_2610);
and U9808 (N_9808,N_697,N_2909);
and U9809 (N_9809,N_643,N_2720);
xor U9810 (N_9810,N_1121,N_1913);
nor U9811 (N_9811,N_1002,N_2179);
and U9812 (N_9812,N_4928,N_4006);
or U9813 (N_9813,N_1484,N_1495);
and U9814 (N_9814,N_3813,N_4893);
and U9815 (N_9815,N_4773,N_2989);
or U9816 (N_9816,N_1220,N_4780);
nand U9817 (N_9817,N_338,N_877);
nor U9818 (N_9818,N_164,N_1492);
and U9819 (N_9819,N_327,N_4080);
nand U9820 (N_9820,N_4655,N_1179);
or U9821 (N_9821,N_1002,N_2694);
or U9822 (N_9822,N_667,N_4936);
and U9823 (N_9823,N_2085,N_2766);
nor U9824 (N_9824,N_3348,N_1198);
or U9825 (N_9825,N_4784,N_3469);
nor U9826 (N_9826,N_254,N_925);
nand U9827 (N_9827,N_29,N_3470);
nand U9828 (N_9828,N_3550,N_849);
and U9829 (N_9829,N_3955,N_2620);
nor U9830 (N_9830,N_1756,N_4064);
or U9831 (N_9831,N_2074,N_4345);
and U9832 (N_9832,N_3469,N_4934);
nor U9833 (N_9833,N_913,N_3979);
or U9834 (N_9834,N_1195,N_4879);
nor U9835 (N_9835,N_1570,N_2483);
nand U9836 (N_9836,N_829,N_4565);
nand U9837 (N_9837,N_2796,N_706);
nand U9838 (N_9838,N_4744,N_1366);
and U9839 (N_9839,N_558,N_4625);
or U9840 (N_9840,N_3353,N_3394);
and U9841 (N_9841,N_4175,N_2168);
and U9842 (N_9842,N_230,N_4866);
or U9843 (N_9843,N_3890,N_1234);
or U9844 (N_9844,N_586,N_3626);
or U9845 (N_9845,N_3575,N_285);
and U9846 (N_9846,N_4482,N_2448);
or U9847 (N_9847,N_4522,N_3046);
nor U9848 (N_9848,N_3317,N_530);
or U9849 (N_9849,N_563,N_3282);
and U9850 (N_9850,N_3983,N_4606);
or U9851 (N_9851,N_1807,N_4639);
or U9852 (N_9852,N_4221,N_3185);
and U9853 (N_9853,N_3250,N_706);
or U9854 (N_9854,N_1321,N_705);
nand U9855 (N_9855,N_2429,N_2012);
or U9856 (N_9856,N_4808,N_4845);
or U9857 (N_9857,N_1811,N_1326);
nor U9858 (N_9858,N_4714,N_3647);
and U9859 (N_9859,N_3034,N_4143);
nor U9860 (N_9860,N_4673,N_1792);
or U9861 (N_9861,N_309,N_818);
nor U9862 (N_9862,N_4436,N_806);
nor U9863 (N_9863,N_1098,N_4304);
nor U9864 (N_9864,N_3174,N_4860);
and U9865 (N_9865,N_1851,N_4443);
or U9866 (N_9866,N_648,N_2121);
and U9867 (N_9867,N_4976,N_405);
and U9868 (N_9868,N_3253,N_2504);
nand U9869 (N_9869,N_2637,N_2887);
or U9870 (N_9870,N_1530,N_2635);
and U9871 (N_9871,N_1678,N_1663);
and U9872 (N_9872,N_3635,N_2438);
nor U9873 (N_9873,N_1732,N_3109);
nand U9874 (N_9874,N_4549,N_2159);
or U9875 (N_9875,N_1886,N_4171);
nand U9876 (N_9876,N_840,N_1764);
nand U9877 (N_9877,N_451,N_852);
nand U9878 (N_9878,N_4203,N_1343);
nor U9879 (N_9879,N_1349,N_3574);
nor U9880 (N_9880,N_442,N_1689);
and U9881 (N_9881,N_1032,N_1325);
or U9882 (N_9882,N_1198,N_683);
nor U9883 (N_9883,N_1069,N_4397);
nor U9884 (N_9884,N_1628,N_4355);
nand U9885 (N_9885,N_4581,N_1087);
or U9886 (N_9886,N_2427,N_3447);
nor U9887 (N_9887,N_2359,N_1095);
nand U9888 (N_9888,N_1898,N_708);
nand U9889 (N_9889,N_2169,N_2537);
nand U9890 (N_9890,N_3414,N_2522);
nand U9891 (N_9891,N_576,N_3361);
nand U9892 (N_9892,N_2338,N_70);
nand U9893 (N_9893,N_4418,N_4663);
nor U9894 (N_9894,N_1784,N_2560);
nand U9895 (N_9895,N_453,N_2074);
and U9896 (N_9896,N_4319,N_1628);
nor U9897 (N_9897,N_3582,N_3545);
or U9898 (N_9898,N_3462,N_569);
or U9899 (N_9899,N_1793,N_1475);
nor U9900 (N_9900,N_1301,N_4602);
nor U9901 (N_9901,N_1450,N_4231);
nor U9902 (N_9902,N_735,N_1037);
nand U9903 (N_9903,N_1930,N_50);
and U9904 (N_9904,N_473,N_4597);
nand U9905 (N_9905,N_3145,N_4733);
nand U9906 (N_9906,N_3268,N_4371);
and U9907 (N_9907,N_2805,N_4674);
or U9908 (N_9908,N_67,N_202);
nor U9909 (N_9909,N_3670,N_4035);
and U9910 (N_9910,N_671,N_4687);
or U9911 (N_9911,N_1613,N_3688);
nand U9912 (N_9912,N_4251,N_3023);
nor U9913 (N_9913,N_1905,N_1566);
nor U9914 (N_9914,N_4132,N_410);
nand U9915 (N_9915,N_3501,N_4317);
and U9916 (N_9916,N_2153,N_1056);
or U9917 (N_9917,N_3996,N_3754);
or U9918 (N_9918,N_2714,N_4410);
and U9919 (N_9919,N_2561,N_4301);
and U9920 (N_9920,N_4990,N_3970);
or U9921 (N_9921,N_2852,N_1985);
xnor U9922 (N_9922,N_2378,N_3292);
nand U9923 (N_9923,N_1793,N_4279);
or U9924 (N_9924,N_1314,N_4358);
and U9925 (N_9925,N_1198,N_671);
nand U9926 (N_9926,N_4514,N_321);
nand U9927 (N_9927,N_375,N_4645);
or U9928 (N_9928,N_177,N_1961);
and U9929 (N_9929,N_1495,N_835);
or U9930 (N_9930,N_3340,N_4753);
nand U9931 (N_9931,N_2425,N_4844);
nor U9932 (N_9932,N_3858,N_3209);
nor U9933 (N_9933,N_4783,N_2119);
nand U9934 (N_9934,N_2239,N_2512);
nor U9935 (N_9935,N_390,N_2101);
or U9936 (N_9936,N_4164,N_2234);
or U9937 (N_9937,N_3838,N_3383);
and U9938 (N_9938,N_3096,N_4842);
or U9939 (N_9939,N_3705,N_4484);
xor U9940 (N_9940,N_4945,N_4894);
and U9941 (N_9941,N_231,N_3633);
nand U9942 (N_9942,N_3090,N_3357);
nand U9943 (N_9943,N_403,N_2295);
nor U9944 (N_9944,N_3771,N_3550);
nand U9945 (N_9945,N_3129,N_3291);
nor U9946 (N_9946,N_2828,N_3821);
nand U9947 (N_9947,N_2997,N_2469);
nand U9948 (N_9948,N_1756,N_2542);
nor U9949 (N_9949,N_404,N_4485);
and U9950 (N_9950,N_1381,N_4080);
and U9951 (N_9951,N_3419,N_999);
and U9952 (N_9952,N_1003,N_1888);
and U9953 (N_9953,N_709,N_2973);
or U9954 (N_9954,N_964,N_248);
and U9955 (N_9955,N_4746,N_2588);
and U9956 (N_9956,N_2044,N_1016);
or U9957 (N_9957,N_2984,N_4494);
nand U9958 (N_9958,N_1784,N_371);
xnor U9959 (N_9959,N_4165,N_1463);
and U9960 (N_9960,N_3812,N_3115);
and U9961 (N_9961,N_3209,N_3836);
and U9962 (N_9962,N_2332,N_3219);
nor U9963 (N_9963,N_493,N_3586);
and U9964 (N_9964,N_3827,N_2474);
and U9965 (N_9965,N_1595,N_2199);
nand U9966 (N_9966,N_4217,N_449);
and U9967 (N_9967,N_401,N_2717);
or U9968 (N_9968,N_184,N_258);
or U9969 (N_9969,N_4699,N_281);
and U9970 (N_9970,N_1868,N_34);
or U9971 (N_9971,N_433,N_810);
nand U9972 (N_9972,N_71,N_2502);
or U9973 (N_9973,N_1880,N_333);
nand U9974 (N_9974,N_2976,N_4572);
nand U9975 (N_9975,N_3441,N_2861);
nand U9976 (N_9976,N_4065,N_2190);
or U9977 (N_9977,N_2608,N_4639);
or U9978 (N_9978,N_1957,N_3541);
or U9979 (N_9979,N_3405,N_75);
nand U9980 (N_9980,N_4167,N_4713);
or U9981 (N_9981,N_3592,N_3166);
and U9982 (N_9982,N_3264,N_4317);
and U9983 (N_9983,N_524,N_2682);
nor U9984 (N_9984,N_2551,N_3297);
or U9985 (N_9985,N_2042,N_4420);
or U9986 (N_9986,N_3464,N_1124);
or U9987 (N_9987,N_1274,N_1609);
nor U9988 (N_9988,N_937,N_3090);
nor U9989 (N_9989,N_472,N_2830);
and U9990 (N_9990,N_453,N_2910);
nand U9991 (N_9991,N_117,N_3674);
nor U9992 (N_9992,N_4685,N_3402);
and U9993 (N_9993,N_4987,N_3516);
nor U9994 (N_9994,N_1056,N_4001);
nand U9995 (N_9995,N_1055,N_142);
or U9996 (N_9996,N_1527,N_4683);
nand U9997 (N_9997,N_2724,N_3065);
nand U9998 (N_9998,N_4761,N_4934);
nand U9999 (N_9999,N_4520,N_3814);
and U10000 (N_10000,N_7426,N_7404);
nand U10001 (N_10001,N_5705,N_9959);
nand U10002 (N_10002,N_9465,N_8032);
and U10003 (N_10003,N_6210,N_5621);
or U10004 (N_10004,N_6166,N_7685);
nand U10005 (N_10005,N_5178,N_5485);
nor U10006 (N_10006,N_9461,N_8544);
and U10007 (N_10007,N_6065,N_5225);
nor U10008 (N_10008,N_9542,N_9171);
nand U10009 (N_10009,N_7898,N_5074);
and U10010 (N_10010,N_8689,N_9293);
nor U10011 (N_10011,N_8569,N_6948);
nand U10012 (N_10012,N_6966,N_9258);
nand U10013 (N_10013,N_7315,N_9492);
nor U10014 (N_10014,N_7938,N_6263);
nand U10015 (N_10015,N_8216,N_8148);
nor U10016 (N_10016,N_5825,N_8137);
and U10017 (N_10017,N_7537,N_5767);
or U10018 (N_10018,N_9877,N_8270);
nand U10019 (N_10019,N_8456,N_6018);
nand U10020 (N_10020,N_7975,N_6628);
nand U10021 (N_10021,N_8878,N_9688);
nand U10022 (N_10022,N_8877,N_6516);
or U10023 (N_10023,N_5087,N_5677);
nand U10024 (N_10024,N_5981,N_7188);
or U10025 (N_10025,N_7942,N_7323);
and U10026 (N_10026,N_7765,N_9384);
and U10027 (N_10027,N_8675,N_8171);
nor U10028 (N_10028,N_6254,N_9325);
nor U10029 (N_10029,N_7491,N_9777);
and U10030 (N_10030,N_6328,N_6380);
or U10031 (N_10031,N_5320,N_9640);
or U10032 (N_10032,N_6591,N_7728);
and U10033 (N_10033,N_7345,N_5037);
nor U10034 (N_10034,N_6069,N_5250);
or U10035 (N_10035,N_6256,N_7335);
nor U10036 (N_10036,N_5090,N_6112);
nand U10037 (N_10037,N_9974,N_6601);
or U10038 (N_10038,N_6897,N_8925);
nand U10039 (N_10039,N_6337,N_6279);
nor U10040 (N_10040,N_8222,N_9597);
or U10041 (N_10041,N_6619,N_7321);
and U10042 (N_10042,N_9180,N_9259);
nor U10043 (N_10043,N_6543,N_8661);
or U10044 (N_10044,N_8752,N_9232);
nand U10045 (N_10045,N_6506,N_9144);
or U10046 (N_10046,N_9145,N_7508);
or U10047 (N_10047,N_9776,N_5586);
nor U10048 (N_10048,N_8250,N_8515);
nor U10049 (N_10049,N_7442,N_7927);
nand U10050 (N_10050,N_5603,N_6859);
and U10051 (N_10051,N_5876,N_5112);
nand U10052 (N_10052,N_8837,N_7724);
nor U10053 (N_10053,N_5181,N_6635);
and U10054 (N_10054,N_6786,N_9717);
nor U10055 (N_10055,N_5489,N_8704);
or U10056 (N_10056,N_8594,N_7073);
nor U10057 (N_10057,N_6431,N_8542);
or U10058 (N_10058,N_9932,N_6004);
nand U10059 (N_10059,N_9169,N_6530);
or U10060 (N_10060,N_9373,N_9341);
nor U10061 (N_10061,N_8649,N_9263);
nor U10062 (N_10062,N_8041,N_6794);
or U10063 (N_10063,N_6643,N_7681);
nand U10064 (N_10064,N_7868,N_6579);
and U10065 (N_10065,N_7989,N_9808);
nor U10066 (N_10066,N_5140,N_5815);
or U10067 (N_10067,N_7547,N_8279);
nor U10068 (N_10068,N_7567,N_7374);
nand U10069 (N_10069,N_6657,N_7124);
nand U10070 (N_10070,N_6818,N_9114);
or U10071 (N_10071,N_8390,N_7209);
nand U10072 (N_10072,N_9677,N_7066);
and U10073 (N_10073,N_8173,N_6711);
nor U10074 (N_10074,N_9553,N_7671);
nor U10075 (N_10075,N_9560,N_9983);
nor U10076 (N_10076,N_6412,N_7816);
nand U10077 (N_10077,N_9874,N_7988);
nand U10078 (N_10078,N_5907,N_8679);
nand U10079 (N_10079,N_9778,N_8083);
and U10080 (N_10080,N_6086,N_9060);
or U10081 (N_10081,N_6400,N_6599);
nor U10082 (N_10082,N_7751,N_9396);
xor U10083 (N_10083,N_6971,N_5416);
and U10084 (N_10084,N_8227,N_7371);
and U10085 (N_10085,N_6504,N_6610);
nand U10086 (N_10086,N_8565,N_9963);
nor U10087 (N_10087,N_7286,N_7088);
and U10088 (N_10088,N_8948,N_9289);
and U10089 (N_10089,N_7604,N_6099);
or U10090 (N_10090,N_8479,N_5326);
or U10091 (N_10091,N_7013,N_6222);
nand U10092 (N_10092,N_7398,N_6158);
nand U10093 (N_10093,N_7193,N_7011);
nand U10094 (N_10094,N_7055,N_5682);
and U10095 (N_10095,N_8048,N_9911);
and U10096 (N_10096,N_8428,N_7977);
or U10097 (N_10097,N_8459,N_5749);
and U10098 (N_10098,N_7603,N_9757);
xor U10099 (N_10099,N_8943,N_7643);
and U10100 (N_10100,N_9636,N_9715);
nand U10101 (N_10101,N_8481,N_8158);
nand U10102 (N_10102,N_5066,N_7769);
xor U10103 (N_10103,N_6829,N_5065);
and U10104 (N_10104,N_6352,N_5939);
or U10105 (N_10105,N_5386,N_7198);
or U10106 (N_10106,N_8728,N_7359);
nor U10107 (N_10107,N_8613,N_6121);
and U10108 (N_10108,N_6274,N_5085);
or U10109 (N_10109,N_9343,N_9463);
and U10110 (N_10110,N_6700,N_5429);
nor U10111 (N_10111,N_9379,N_5607);
or U10112 (N_10112,N_5113,N_8825);
nand U10113 (N_10113,N_6147,N_5589);
nor U10114 (N_10114,N_9956,N_7994);
or U10115 (N_10115,N_5724,N_7559);
nor U10116 (N_10116,N_6353,N_8950);
nor U10117 (N_10117,N_5511,N_5512);
nor U10118 (N_10118,N_8091,N_7645);
and U10119 (N_10119,N_9084,N_7249);
nand U10120 (N_10120,N_6653,N_5158);
nor U10121 (N_10121,N_5758,N_9495);
or U10122 (N_10122,N_7034,N_6316);
xnor U10123 (N_10123,N_6060,N_5109);
nand U10124 (N_10124,N_6025,N_6347);
and U10125 (N_10125,N_7272,N_8806);
or U10126 (N_10126,N_7592,N_6722);
or U10127 (N_10127,N_9870,N_6361);
xnor U10128 (N_10128,N_7318,N_6796);
or U10129 (N_10129,N_8529,N_9649);
or U10130 (N_10130,N_8478,N_7379);
nand U10131 (N_10131,N_9127,N_9826);
nor U10132 (N_10132,N_8169,N_7557);
nor U10133 (N_10133,N_5451,N_7697);
nand U10134 (N_10134,N_9003,N_7739);
or U10135 (N_10135,N_9633,N_6186);
nand U10136 (N_10136,N_6847,N_9875);
nor U10137 (N_10137,N_7495,N_8140);
and U10138 (N_10138,N_6654,N_5139);
and U10139 (N_10139,N_7528,N_8494);
and U10140 (N_10140,N_5455,N_8095);
or U10141 (N_10141,N_9628,N_8622);
nand U10142 (N_10142,N_5711,N_9661);
nand U10143 (N_10143,N_8566,N_8046);
nand U10144 (N_10144,N_6527,N_5557);
or U10145 (N_10145,N_5367,N_5587);
nor U10146 (N_10146,N_7560,N_5306);
and U10147 (N_10147,N_9008,N_6446);
nor U10148 (N_10148,N_5432,N_7041);
and U10149 (N_10149,N_9091,N_6551);
or U10150 (N_10150,N_7146,N_7435);
and U10151 (N_10151,N_9843,N_9013);
and U10152 (N_10152,N_6091,N_6939);
nor U10153 (N_10153,N_8753,N_6178);
and U10154 (N_10154,N_6670,N_6519);
nand U10155 (N_10155,N_6355,N_5010);
and U10156 (N_10156,N_6996,N_5226);
nand U10157 (N_10157,N_5413,N_9080);
nand U10158 (N_10158,N_6265,N_7244);
nor U10159 (N_10159,N_8920,N_7863);
and U10160 (N_10160,N_6799,N_9637);
nand U10161 (N_10161,N_8729,N_7782);
or U10162 (N_10162,N_6871,N_9907);
or U10163 (N_10163,N_8611,N_8457);
nand U10164 (N_10164,N_5410,N_9025);
or U10165 (N_10165,N_7171,N_5897);
and U10166 (N_10166,N_9743,N_6803);
and U10167 (N_10167,N_8693,N_5992);
and U10168 (N_10168,N_5963,N_6372);
nand U10169 (N_10169,N_5577,N_6157);
nand U10170 (N_10170,N_5400,N_8589);
and U10171 (N_10171,N_7078,N_6614);
nand U10172 (N_10172,N_9177,N_7992);
and U10173 (N_10173,N_9270,N_5039);
nand U10174 (N_10174,N_8023,N_6445);
and U10175 (N_10175,N_7651,N_8998);
and U10176 (N_10176,N_6167,N_8197);
and U10177 (N_10177,N_5098,N_6910);
nor U10178 (N_10178,N_8709,N_5299);
nand U10179 (N_10179,N_5950,N_7403);
or U10180 (N_10180,N_6259,N_5301);
nand U10181 (N_10181,N_5424,N_9569);
and U10182 (N_10182,N_6641,N_9752);
or U10183 (N_10183,N_8666,N_8024);
nand U10184 (N_10184,N_5076,N_9030);
nand U10185 (N_10185,N_7846,N_7817);
nor U10186 (N_10186,N_6247,N_6735);
nand U10187 (N_10187,N_6070,N_9249);
nor U10188 (N_10188,N_5943,N_9271);
nand U10189 (N_10189,N_5809,N_9486);
or U10190 (N_10190,N_6673,N_6894);
and U10191 (N_10191,N_5606,N_7044);
nand U10192 (N_10192,N_6189,N_6932);
and U10193 (N_10193,N_6623,N_8685);
or U10194 (N_10194,N_8992,N_8360);
or U10195 (N_10195,N_7208,N_5435);
nor U10196 (N_10196,N_7307,N_9286);
nand U10197 (N_10197,N_6392,N_7781);
nor U10198 (N_10198,N_8558,N_7909);
or U10199 (N_10199,N_9667,N_8368);
nor U10200 (N_10200,N_5669,N_8990);
or U10201 (N_10201,N_7237,N_8277);
nand U10202 (N_10202,N_8555,N_7481);
and U10203 (N_10203,N_6047,N_7434);
or U10204 (N_10204,N_7280,N_8329);
or U10205 (N_10205,N_6891,N_8784);
or U10206 (N_10206,N_8288,N_5900);
and U10207 (N_10207,N_9507,N_7761);
nor U10208 (N_10208,N_7918,N_6183);
or U10209 (N_10209,N_6766,N_7053);
or U10210 (N_10210,N_8035,N_5539);
nand U10211 (N_10211,N_6508,N_7185);
nor U10212 (N_10212,N_5315,N_5516);
xor U10213 (N_10213,N_9687,N_8995);
nand U10214 (N_10214,N_7687,N_8874);
nor U10215 (N_10215,N_7695,N_7199);
nor U10216 (N_10216,N_9443,N_6221);
or U10217 (N_10217,N_5363,N_7506);
or U10218 (N_10218,N_5686,N_6108);
and U10219 (N_10219,N_5638,N_8536);
or U10220 (N_10220,N_8777,N_9538);
and U10221 (N_10221,N_7396,N_5760);
xnor U10222 (N_10222,N_5911,N_8885);
or U10223 (N_10223,N_8802,N_5044);
nand U10224 (N_10224,N_9958,N_7692);
nor U10225 (N_10225,N_8087,N_7139);
xnor U10226 (N_10226,N_9788,N_8859);
and U10227 (N_10227,N_7973,N_7416);
or U10228 (N_10228,N_5079,N_6919);
nand U10229 (N_10229,N_6726,N_6034);
or U10230 (N_10230,N_5756,N_5675);
and U10231 (N_10231,N_6945,N_9849);
and U10232 (N_10232,N_6063,N_5501);
and U10233 (N_10233,N_9238,N_9317);
and U10234 (N_10234,N_6305,N_9996);
nand U10235 (N_10235,N_7325,N_5019);
nand U10236 (N_10236,N_9601,N_9344);
or U10237 (N_10237,N_5574,N_7239);
xnor U10238 (N_10238,N_6406,N_7402);
nand U10239 (N_10239,N_5811,N_5393);
or U10240 (N_10240,N_7382,N_8104);
or U10241 (N_10241,N_7753,N_9598);
and U10242 (N_10242,N_5034,N_5975);
nand U10243 (N_10243,N_7094,N_9196);
nor U10244 (N_10244,N_8714,N_9872);
nand U10245 (N_10245,N_7738,N_7376);
and U10246 (N_10246,N_8111,N_9156);
or U10247 (N_10247,N_6379,N_9668);
and U10248 (N_10248,N_8337,N_7337);
or U10249 (N_10249,N_6160,N_9896);
or U10250 (N_10250,N_5765,N_9424);
or U10251 (N_10251,N_8644,N_6507);
nor U10252 (N_10252,N_9751,N_6697);
or U10253 (N_10253,N_7845,N_7458);
nor U10254 (N_10254,N_6049,N_7159);
nand U10255 (N_10255,N_5530,N_5346);
nand U10256 (N_10256,N_6233,N_5506);
nor U10257 (N_10257,N_7120,N_7507);
or U10258 (N_10258,N_7657,N_5275);
nor U10259 (N_10259,N_7241,N_5696);
and U10260 (N_10260,N_8126,N_7192);
and U10261 (N_10261,N_9950,N_6200);
or U10262 (N_10262,N_6912,N_8069);
and U10263 (N_10263,N_7541,N_6691);
nor U10264 (N_10264,N_6864,N_7774);
or U10265 (N_10265,N_9445,N_7872);
nand U10266 (N_10266,N_5647,N_7722);
and U10267 (N_10267,N_5021,N_9256);
nor U10268 (N_10268,N_5717,N_8884);
nand U10269 (N_10269,N_9747,N_8653);
or U10270 (N_10270,N_9452,N_7366);
and U10271 (N_10271,N_8863,N_5610);
and U10272 (N_10272,N_8180,N_9561);
and U10273 (N_10273,N_5273,N_5077);
nor U10274 (N_10274,N_6538,N_6963);
and U10275 (N_10275,N_6028,N_6177);
nor U10276 (N_10276,N_8512,N_8226);
nand U10277 (N_10277,N_9061,N_7411);
nor U10278 (N_10278,N_7634,N_5073);
or U10279 (N_10279,N_6216,N_5272);
nor U10280 (N_10280,N_8167,N_5674);
nand U10281 (N_10281,N_8574,N_7354);
nand U10282 (N_10282,N_7068,N_6810);
and U10283 (N_10283,N_7889,N_6208);
nand U10284 (N_10284,N_5715,N_9910);
nor U10285 (N_10285,N_7936,N_8487);
and U10286 (N_10286,N_9547,N_9654);
nor U10287 (N_10287,N_7327,N_9237);
and U10288 (N_10288,N_7503,N_6946);
nor U10289 (N_10289,N_6451,N_9502);
or U10290 (N_10290,N_8533,N_6258);
xnor U10291 (N_10291,N_5327,N_6212);
and U10292 (N_10292,N_7866,N_7523);
or U10293 (N_10293,N_5642,N_7274);
and U10294 (N_10294,N_9239,N_9346);
nand U10295 (N_10295,N_9527,N_6284);
and U10296 (N_10296,N_6249,N_7572);
or U10297 (N_10297,N_8781,N_9473);
nor U10298 (N_10298,N_5145,N_5742);
nand U10299 (N_10299,N_9916,N_8364);
or U10300 (N_10300,N_6556,N_6731);
nand U10301 (N_10301,N_8519,N_5895);
nor U10302 (N_10302,N_8371,N_9570);
or U10303 (N_10303,N_6933,N_9616);
nor U10304 (N_10304,N_8934,N_7974);
or U10305 (N_10305,N_5371,N_7777);
nor U10306 (N_10306,N_5161,N_5359);
nand U10307 (N_10307,N_5254,N_6942);
or U10308 (N_10308,N_9504,N_5388);
nand U10309 (N_10309,N_6908,N_9438);
nor U10310 (N_10310,N_6931,N_8094);
nor U10311 (N_10311,N_6532,N_5912);
and U10312 (N_10312,N_8553,N_7395);
and U10313 (N_10313,N_9300,N_8330);
and U10314 (N_10314,N_7551,N_6453);
or U10315 (N_10315,N_7386,N_8548);
and U10316 (N_10316,N_5704,N_5620);
and U10317 (N_10317,N_6483,N_5660);
and U10318 (N_10318,N_6501,N_9927);
or U10319 (N_10319,N_5352,N_7549);
and U10320 (N_10320,N_7037,N_6667);
or U10321 (N_10321,N_9921,N_6813);
nor U10322 (N_10322,N_8309,N_8798);
and U10323 (N_10323,N_9857,N_8531);
and U10324 (N_10324,N_6498,N_5447);
or U10325 (N_10325,N_5787,N_9366);
and U10326 (N_10326,N_9475,N_8852);
nand U10327 (N_10327,N_9047,N_8450);
and U10328 (N_10328,N_7186,N_7958);
and U10329 (N_10329,N_8101,N_9323);
xor U10330 (N_10330,N_5430,N_7656);
nand U10331 (N_10331,N_8634,N_7134);
and U10332 (N_10332,N_7172,N_5819);
nand U10333 (N_10333,N_7980,N_9407);
and U10334 (N_10334,N_6301,N_6444);
xnor U10335 (N_10335,N_7847,N_7500);
xnor U10336 (N_10336,N_7900,N_6826);
or U10337 (N_10337,N_8743,N_8705);
and U10338 (N_10338,N_8168,N_7223);
nor U10339 (N_10339,N_6023,N_5857);
nand U10340 (N_10340,N_5041,N_9201);
or U10341 (N_10341,N_7373,N_9222);
and U10342 (N_10342,N_9363,N_9573);
nand U10343 (N_10343,N_5986,N_8970);
and U10344 (N_10344,N_9490,N_5583);
and U10345 (N_10345,N_8882,N_8655);
and U10346 (N_10346,N_7550,N_9650);
nor U10347 (N_10347,N_9883,N_8298);
nand U10348 (N_10348,N_6031,N_7473);
nor U10349 (N_10349,N_5737,N_5394);
nor U10350 (N_10350,N_5990,N_6480);
nor U10351 (N_10351,N_7160,N_7408);
and U10352 (N_10352,N_9675,N_5699);
and U10353 (N_10353,N_5344,N_7114);
or U10354 (N_10354,N_6563,N_8243);
nor U10355 (N_10355,N_7201,N_5951);
nor U10356 (N_10356,N_6751,N_7729);
or U10357 (N_10357,N_8489,N_7467);
nand U10358 (N_10358,N_9653,N_8328);
nor U10359 (N_10359,N_5337,N_9565);
nor U10360 (N_10360,N_7608,N_8306);
nand U10361 (N_10361,N_8303,N_9035);
nor U10362 (N_10362,N_6409,N_5189);
and U10363 (N_10363,N_9513,N_5199);
nand U10364 (N_10364,N_9726,N_7632);
nand U10365 (N_10365,N_8055,N_8526);
xnor U10366 (N_10366,N_8405,N_8790);
nor U10367 (N_10367,N_8654,N_7581);
nor U10368 (N_10368,N_8464,N_8872);
nand U10369 (N_10369,N_6913,N_6674);
or U10370 (N_10370,N_5117,N_9749);
or U10371 (N_10371,N_5313,N_7513);
nor U10372 (N_10372,N_5579,N_7644);
nor U10373 (N_10373,N_7202,N_7438);
nor U10374 (N_10374,N_8727,N_8366);
nand U10375 (N_10375,N_6367,N_9674);
nand U10376 (N_10376,N_6607,N_5380);
and U10377 (N_10377,N_8517,N_7133);
or U10378 (N_10378,N_5595,N_8170);
or U10379 (N_10379,N_8490,N_5304);
nor U10380 (N_10380,N_9491,N_7691);
and U10381 (N_10381,N_7254,N_8812);
or U10382 (N_10382,N_9214,N_9195);
nor U10383 (N_10383,N_5976,N_5269);
and U10384 (N_10384,N_7625,N_7968);
nand U10385 (N_10385,N_7228,N_8310);
or U10386 (N_10386,N_7177,N_8474);
nand U10387 (N_10387,N_7489,N_6080);
nand U10388 (N_10388,N_9820,N_9348);
and U10389 (N_10389,N_7540,N_7677);
nor U10390 (N_10390,N_8895,N_8815);
nor U10391 (N_10391,N_6911,N_5614);
nand U10392 (N_10392,N_6548,N_5486);
and U10393 (N_10393,N_6191,N_7061);
or U10394 (N_10394,N_6225,N_7496);
and U10395 (N_10395,N_9115,N_5173);
nand U10396 (N_10396,N_9083,N_5059);
nor U10397 (N_10397,N_9016,N_6856);
nand U10398 (N_10398,N_6808,N_6987);
nand U10399 (N_10399,N_8089,N_5526);
or U10400 (N_10400,N_7902,N_6123);
or U10401 (N_10401,N_6707,N_9799);
and U10402 (N_10402,N_5234,N_9006);
and U10403 (N_10403,N_9891,N_5740);
nor U10404 (N_10404,N_7090,N_5844);
nor U10405 (N_10405,N_7590,N_7447);
or U10406 (N_10406,N_6709,N_7675);
nor U10407 (N_10407,N_6291,N_7731);
xor U10408 (N_10408,N_6116,N_5288);
and U10409 (N_10409,N_9318,N_7394);
and U10410 (N_10410,N_8868,N_5858);
or U10411 (N_10411,N_7837,N_6103);
nor U10412 (N_10412,N_7110,N_8813);
or U10413 (N_10413,N_5246,N_6062);
nand U10414 (N_10414,N_6957,N_5707);
or U10415 (N_10415,N_6294,N_9304);
nand U10416 (N_10416,N_6659,N_7484);
nor U10417 (N_10417,N_6961,N_8347);
or U10418 (N_10418,N_6229,N_9064);
nand U10419 (N_10419,N_7562,N_7615);
or U10420 (N_10420,N_5418,N_9621);
nor U10421 (N_10421,N_5078,N_5519);
nor U10422 (N_10422,N_7734,N_6111);
nand U10423 (N_10423,N_8266,N_8818);
or U10424 (N_10424,N_8246,N_6101);
and U10425 (N_10425,N_6977,N_5396);
or U10426 (N_10426,N_8952,N_6482);
and U10427 (N_10427,N_6584,N_9582);
or U10428 (N_10428,N_6005,N_8592);
or U10429 (N_10429,N_6289,N_8928);
nor U10430 (N_10430,N_5781,N_7265);
or U10431 (N_10431,N_8201,N_6693);
or U10432 (N_10432,N_7524,N_9980);
nor U10433 (N_10433,N_7256,N_9148);
and U10434 (N_10434,N_9943,N_9545);
nand U10435 (N_10435,N_6940,N_6529);
nor U10436 (N_10436,N_5670,N_6644);
or U10437 (N_10437,N_9604,N_6600);
nand U10438 (N_10438,N_5020,N_5434);
nand U10439 (N_10439,N_8407,N_9692);
or U10440 (N_10440,N_8691,N_9260);
and U10441 (N_10441,N_8738,N_6573);
or U10442 (N_10442,N_9821,N_6895);
and U10443 (N_10443,N_9034,N_6575);
nand U10444 (N_10444,N_6534,N_6218);
nor U10445 (N_10445,N_6999,N_6950);
nor U10446 (N_10446,N_9969,N_5193);
nand U10447 (N_10447,N_5132,N_7985);
and U10448 (N_10448,N_8660,N_7848);
nor U10449 (N_10449,N_9536,N_7468);
and U10450 (N_10450,N_8412,N_7130);
nand U10451 (N_10451,N_8875,N_9721);
nand U10452 (N_10452,N_7026,N_8037);
and U10453 (N_10453,N_6798,N_8670);
and U10454 (N_10454,N_7147,N_5517);
nor U10455 (N_10455,N_5631,N_9990);
or U10456 (N_10456,N_9262,N_9813);
nor U10457 (N_10457,N_9905,N_8640);
nand U10458 (N_10458,N_5513,N_6982);
and U10459 (N_10459,N_9199,N_6071);
nand U10460 (N_10460,N_5835,N_6943);
or U10461 (N_10461,N_8281,N_8143);
nand U10462 (N_10462,N_8406,N_9989);
and U10463 (N_10463,N_7275,N_6980);
nand U10464 (N_10464,N_8439,N_8475);
and U10465 (N_10465,N_6172,N_8867);
nor U10466 (N_10466,N_9052,N_6102);
and U10467 (N_10467,N_6886,N_6268);
and U10468 (N_10468,N_9672,N_5443);
nor U10469 (N_10469,N_8734,N_6240);
or U10470 (N_10470,N_5134,N_9552);
nor U10471 (N_10471,N_9278,N_5955);
or U10472 (N_10472,N_8500,N_9288);
nor U10473 (N_10473,N_5473,N_7883);
and U10474 (N_10474,N_8614,N_7620);
nor U10475 (N_10475,N_5439,N_6010);
and U10476 (N_10476,N_8926,N_6701);
and U10477 (N_10477,N_9596,N_8120);
nor U10478 (N_10478,N_7951,N_9135);
and U10479 (N_10479,N_6609,N_5397);
nor U10480 (N_10480,N_8584,N_9863);
and U10481 (N_10481,N_5457,N_9997);
and U10482 (N_10482,N_9944,N_7331);
or U10483 (N_10483,N_9931,N_8445);
nor U10484 (N_10484,N_5979,N_6343);
and U10485 (N_10485,N_5228,N_8627);
xor U10486 (N_10486,N_6752,N_9031);
or U10487 (N_10487,N_8889,N_5768);
or U10488 (N_10488,N_5002,N_9436);
nor U10489 (N_10489,N_9768,N_6134);
nor U10490 (N_10490,N_9274,N_8403);
xnor U10491 (N_10491,N_6277,N_7897);
and U10492 (N_10492,N_5624,N_8065);
nor U10493 (N_10493,N_6787,N_8570);
and U10494 (N_10494,N_6662,N_9704);
and U10495 (N_10495,N_9835,N_5190);
or U10496 (N_10496,N_7684,N_5678);
nand U10497 (N_10497,N_6459,N_9814);
and U10498 (N_10498,N_9085,N_6627);
and U10499 (N_10499,N_6576,N_7991);
and U10500 (N_10500,N_9982,N_7020);
or U10501 (N_10501,N_5458,N_7940);
or U10502 (N_10502,N_8383,N_9694);
and U10503 (N_10503,N_5166,N_9110);
nand U10504 (N_10504,N_6282,N_8286);
nand U10505 (N_10505,N_8886,N_5532);
or U10506 (N_10506,N_6339,N_7353);
and U10507 (N_10507,N_9515,N_7653);
and U10508 (N_10508,N_6533,N_5036);
and U10509 (N_10509,N_6286,N_9683);
nand U10510 (N_10510,N_9790,N_9732);
or U10511 (N_10511,N_5713,N_7937);
nor U10512 (N_10512,N_9386,N_7263);
and U10513 (N_10513,N_5636,N_7945);
nor U10514 (N_10514,N_6580,N_7077);
nor U10515 (N_10515,N_9722,N_9450);
nor U10516 (N_10516,N_9748,N_8278);
or U10517 (N_10517,N_8861,N_7270);
or U10518 (N_10518,N_9656,N_8665);
and U10519 (N_10519,N_7079,N_5123);
nor U10520 (N_10520,N_7179,N_7672);
nor U10521 (N_10521,N_6262,N_7170);
nand U10522 (N_10522,N_8983,N_5364);
nand U10523 (N_10523,N_7300,N_7637);
and U10524 (N_10524,N_8701,N_9111);
or U10525 (N_10525,N_8638,N_9125);
or U10526 (N_10526,N_6678,N_9311);
and U10527 (N_10527,N_9518,N_9054);
and U10528 (N_10528,N_6378,N_8596);
xor U10529 (N_10529,N_5692,N_7758);
nor U10530 (N_10530,N_5808,N_9053);
nor U10531 (N_10531,N_7049,N_6624);
nand U10532 (N_10532,N_7427,N_5919);
nand U10533 (N_10533,N_7222,N_7564);
nand U10534 (N_10534,N_5075,N_7521);
nand U10535 (N_10535,N_5360,N_8480);
and U10536 (N_10536,N_6842,N_8710);
or U10537 (N_10537,N_7164,N_5318);
nand U10538 (N_10538,N_8763,N_7448);
nor U10539 (N_10539,N_8712,N_8823);
and U10540 (N_10540,N_9073,N_8294);
and U10541 (N_10541,N_8608,N_6037);
and U10542 (N_10542,N_6747,N_9149);
nand U10543 (N_10543,N_6323,N_5507);
or U10544 (N_10544,N_9853,N_5032);
nand U10545 (N_10545,N_8668,N_6503);
nor U10546 (N_10546,N_8050,N_9999);
nor U10547 (N_10547,N_6590,N_7098);
nor U10548 (N_10548,N_5389,N_5022);
nand U10549 (N_10549,N_6528,N_6168);
nand U10550 (N_10550,N_6244,N_5659);
or U10551 (N_10551,N_5798,N_6003);
nand U10552 (N_10552,N_8788,N_7747);
nand U10553 (N_10553,N_9421,N_8678);
nor U10554 (N_10554,N_6734,N_8836);
nand U10555 (N_10555,N_8346,N_9772);
and U10556 (N_10556,N_9718,N_5584);
and U10557 (N_10557,N_8149,N_9868);
and U10558 (N_10558,N_5114,N_8636);
nor U10559 (N_10559,N_9466,N_5893);
or U10560 (N_10560,N_8392,N_7682);
or U10561 (N_10561,N_9608,N_5806);
nor U10562 (N_10562,N_7887,N_9992);
nand U10563 (N_10563,N_9435,N_7745);
or U10564 (N_10564,N_9333,N_9208);
xnor U10565 (N_10565,N_6287,N_9090);
nand U10566 (N_10566,N_8265,N_9055);
and U10567 (N_10567,N_8677,N_7439);
nor U10568 (N_10568,N_5001,N_6235);
nand U10569 (N_10569,N_6415,N_9622);
nor U10570 (N_10570,N_8547,N_7628);
and U10571 (N_10571,N_6214,N_7517);
xor U10572 (N_10572,N_9224,N_7827);
and U10573 (N_10573,N_8759,N_6439);
nand U10574 (N_10574,N_7294,N_7667);
nand U10575 (N_10575,N_9918,N_8344);
nor U10576 (N_10576,N_9809,N_9763);
nor U10577 (N_10577,N_8433,N_8833);
and U10578 (N_10578,N_7140,N_9457);
xnor U10579 (N_10579,N_9903,N_6348);
nor U10580 (N_10580,N_7755,N_7807);
nand U10581 (N_10581,N_6384,N_5817);
nor U10582 (N_10582,N_9471,N_7841);
or U10583 (N_10583,N_9183,N_6419);
and U10584 (N_10584,N_9272,N_6311);
or U10585 (N_10585,N_8438,N_5878);
nor U10586 (N_10586,N_7640,N_6655);
nor U10587 (N_10587,N_7806,N_6298);
and U10588 (N_10588,N_6861,N_5813);
nand U10589 (N_10589,N_8534,N_7856);
nor U10590 (N_10590,N_6457,N_6537);
nand U10591 (N_10591,N_7391,N_6219);
or U10592 (N_10592,N_8414,N_9556);
or U10593 (N_10593,N_9630,N_5243);
nor U10594 (N_10594,N_6979,N_5349);
nor U10595 (N_10595,N_9702,N_9225);
nor U10596 (N_10596,N_5915,N_9470);
nand U10597 (N_10597,N_7118,N_7579);
and U10598 (N_10598,N_5358,N_8754);
nand U10599 (N_10599,N_9736,N_7003);
nor U10600 (N_10600,N_5661,N_7017);
nand U10601 (N_10601,N_9682,N_7915);
nand U10602 (N_10602,N_9022,N_5264);
nor U10603 (N_10603,N_6646,N_8102);
xor U10604 (N_10604,N_5616,N_6113);
and U10605 (N_10605,N_9349,N_5651);
or U10606 (N_10606,N_7154,N_5754);
and U10607 (N_10607,N_6778,N_5375);
and U10608 (N_10608,N_6118,N_8846);
and U10609 (N_10609,N_8191,N_7924);
or U10610 (N_10610,N_8085,N_8469);
or U10611 (N_10611,N_8311,N_9487);
nor U10612 (N_10612,N_6078,N_7896);
nor U10613 (N_10613,N_7674,N_5023);
nand U10614 (N_10614,N_6689,N_5446);
nand U10615 (N_10615,N_9646,N_6761);
nand U10616 (N_10616,N_5101,N_9059);
or U10617 (N_10617,N_8662,N_8210);
nand U10618 (N_10618,N_6626,N_9158);
and U10619 (N_10619,N_9303,N_6471);
or U10620 (N_10620,N_7197,N_8301);
nand U10621 (N_10621,N_9758,N_6536);
or U10622 (N_10622,N_9458,N_9045);
nand U10623 (N_10623,N_9126,N_7297);
nor U10624 (N_10624,N_7378,N_9714);
or U10625 (N_10625,N_9615,N_6145);
nor U10626 (N_10626,N_8865,N_6849);
nor U10627 (N_10627,N_9592,N_7363);
xnor U10628 (N_10628,N_5590,N_6696);
nand U10629 (N_10629,N_8003,N_7966);
nand U10630 (N_10630,N_9953,N_7138);
xnor U10631 (N_10631,N_5008,N_8098);
nor U10632 (N_10632,N_9081,N_8052);
nand U10633 (N_10633,N_8483,N_9729);
nand U10634 (N_10634,N_5227,N_9501);
or U10635 (N_10635,N_7580,N_6317);
nand U10636 (N_10636,N_5650,N_5184);
nand U10637 (N_10637,N_7123,N_6125);
or U10638 (N_10638,N_8774,N_5260);
or U10639 (N_10639,N_7906,N_7907);
or U10640 (N_10640,N_6687,N_8796);
nor U10641 (N_10641,N_9423,N_5029);
or U10642 (N_10642,N_6740,N_9494);
nor U10643 (N_10643,N_9362,N_8136);
or U10644 (N_10644,N_9669,N_6524);
nor U10645 (N_10645,N_5908,N_6307);
nor U10646 (N_10646,N_6930,N_6374);
and U10647 (N_10647,N_6360,N_7798);
nand U10648 (N_10648,N_6690,N_9889);
nand U10649 (N_10649,N_9218,N_6830);
nor U10650 (N_10650,N_5818,N_7568);
and U10651 (N_10651,N_7861,N_8761);
nor U10652 (N_10652,N_5961,N_5125);
nor U10653 (N_10653,N_6892,N_7785);
nand U10654 (N_10654,N_7074,N_5267);
and U10655 (N_10655,N_7112,N_8384);
or U10656 (N_10656,N_8578,N_9824);
nand U10657 (N_10657,N_9015,N_5498);
or U10658 (N_10658,N_9696,N_5252);
xnor U10659 (N_10659,N_7183,N_8340);
nor U10660 (N_10660,N_7246,N_9534);
or U10661 (N_10661,N_8426,N_6002);
or U10662 (N_10662,N_9629,N_8650);
nand U10663 (N_10663,N_5251,N_9591);
nor U10664 (N_10664,N_5481,N_7108);
or U10665 (N_10665,N_8587,N_8549);
nand U10666 (N_10666,N_8385,N_6595);
and U10667 (N_10667,N_7892,N_9779);
or U10668 (N_10668,N_5639,N_7278);
and U10669 (N_10669,N_9097,N_6391);
and U10670 (N_10670,N_5546,N_7352);
and U10671 (N_10671,N_7999,N_8732);
nand U10672 (N_10672,N_6899,N_9773);
nand U10673 (N_10673,N_6458,N_5263);
nand U10674 (N_10674,N_5195,N_5549);
nor U10675 (N_10675,N_6661,N_7631);
nor U10676 (N_10676,N_8225,N_5239);
nand U10677 (N_10677,N_9801,N_5471);
or U10678 (N_10678,N_7871,N_7763);
xnor U10679 (N_10679,N_6093,N_9104);
or U10680 (N_10680,N_7979,N_9728);
nor U10681 (N_10681,N_8848,N_8271);
or U10682 (N_10682,N_5072,N_8341);
or U10683 (N_10683,N_8527,N_9532);
nand U10684 (N_10684,N_7301,N_6727);
or U10685 (N_10685,N_9680,N_9614);
nand U10686 (N_10686,N_7828,N_7212);
nor U10687 (N_10687,N_6190,N_9254);
nand U10688 (N_10688,N_8590,N_6165);
or U10689 (N_10689,N_7702,N_6237);
nand U10690 (N_10690,N_8805,N_5361);
nand U10691 (N_10691,N_7167,N_9213);
xor U10692 (N_10692,N_7716,N_5063);
and U10693 (N_10693,N_6935,N_8940);
nor U10694 (N_10694,N_9419,N_7018);
xor U10695 (N_10695,N_6059,N_5155);
nand U10696 (N_10696,N_8068,N_7972);
nand U10697 (N_10697,N_9094,N_8935);
nand U10698 (N_10698,N_8751,N_6934);
and U10699 (N_10699,N_5323,N_9402);
or U10700 (N_10700,N_6267,N_6617);
and U10701 (N_10701,N_5069,N_5800);
nor U10702 (N_10702,N_7042,N_5731);
nand U10703 (N_10703,N_8073,N_8647);
and U10704 (N_10704,N_5794,N_8307);
nor U10705 (N_10705,N_8025,N_7712);
nor U10706 (N_10706,N_8378,N_6198);
and U10707 (N_10707,N_6327,N_8179);
and U10708 (N_10708,N_6021,N_7433);
nand U10709 (N_10709,N_8280,N_9962);
nor U10710 (N_10710,N_9351,N_7583);
nand U10711 (N_10711,N_6962,N_8979);
and U10712 (N_10712,N_9429,N_6057);
nand U10713 (N_10713,N_5658,N_7984);
nand U10714 (N_10714,N_9825,N_9057);
and U10715 (N_10715,N_6454,N_7029);
nand U10716 (N_10716,N_6718,N_9469);
nor U10717 (N_10717,N_5555,N_6616);
nand U10718 (N_10718,N_6040,N_9077);
or U10719 (N_10719,N_8609,N_5335);
nor U10720 (N_10720,N_5454,N_5727);
nand U10721 (N_10721,N_8824,N_7191);
nand U10722 (N_10722,N_9938,N_5536);
nand U10723 (N_10723,N_7121,N_5971);
nand U10724 (N_10724,N_7510,N_8964);
and U10725 (N_10725,N_7285,N_9841);
nor U10726 (N_10726,N_6958,N_8220);
and U10727 (N_10727,N_8577,N_9355);
nor U10728 (N_10728,N_6224,N_7622);
or U10729 (N_10729,N_8618,N_7356);
and U10730 (N_10730,N_6776,N_6468);
and U10731 (N_10731,N_9086,N_5014);
nand U10732 (N_10732,N_7832,N_8388);
and U10733 (N_10733,N_8461,N_5208);
and U10734 (N_10734,N_7509,N_8370);
xnor U10735 (N_10735,N_8845,N_5177);
nor U10736 (N_10736,N_6683,N_5325);
nand U10737 (N_10737,N_9631,N_6677);
or U10738 (N_10738,N_9626,N_8321);
nand U10739 (N_10739,N_5343,N_6066);
nor U10740 (N_10740,N_6801,N_9642);
nand U10741 (N_10741,N_5093,N_5110);
nor U10742 (N_10742,N_9934,N_8767);
and U10743 (N_10743,N_9244,N_5560);
or U10744 (N_10744,N_9866,N_5690);
or U10745 (N_10745,N_9342,N_7538);
nand U10746 (N_10746,N_9498,N_6672);
nor U10747 (N_10747,N_5626,N_5061);
or U10748 (N_10748,N_8498,N_8349);
and U10749 (N_10749,N_9005,N_6882);
nand U10750 (N_10750,N_7231,N_5625);
nand U10751 (N_10751,N_7119,N_7910);
nor U10752 (N_10752,N_7811,N_6521);
nor U10753 (N_10753,N_6780,N_8108);
nor U10754 (N_10754,N_7400,N_7369);
and U10755 (N_10755,N_7913,N_7440);
or U10756 (N_10756,N_8183,N_9720);
nand U10757 (N_10757,N_6100,N_5223);
nand U10758 (N_10758,N_9655,N_9082);
nand U10759 (N_10759,N_5571,N_7200);
nand U10760 (N_10760,N_9564,N_9464);
or U10761 (N_10761,N_7006,N_6266);
and U10762 (N_10762,N_8255,N_5212);
nand U10763 (N_10763,N_5777,N_7893);
xnor U10764 (N_10764,N_5202,N_6917);
or U10765 (N_10765,N_8013,N_7488);
or U10766 (N_10766,N_7157,N_7982);
nand U10767 (N_10767,N_6463,N_9952);
or U10768 (N_10768,N_7526,N_8467);
nor U10769 (N_10769,N_8532,N_5970);
and U10770 (N_10770,N_6870,N_9827);
nand U10771 (N_10771,N_6345,N_9012);
and U10772 (N_10772,N_6568,N_7216);
nor U10773 (N_10773,N_6938,N_5822);
and U10774 (N_10774,N_8072,N_8657);
or U10775 (N_10775,N_9425,N_6625);
nand U10776 (N_10776,N_9798,N_8141);
and U10777 (N_10777,N_9138,N_8021);
and U10778 (N_10778,N_6603,N_9581);
nand U10779 (N_10779,N_9723,N_8984);
and U10780 (N_10780,N_8664,N_5033);
and U10781 (N_10781,N_7372,N_6276);
nand U10782 (N_10782,N_5369,N_7299);
nand U10783 (N_10783,N_7415,N_5880);
nand U10784 (N_10784,N_6874,N_5009);
or U10785 (N_10785,N_8695,N_5982);
nand U10786 (N_10786,N_5652,N_8510);
or U10787 (N_10787,N_9769,N_5107);
and U10788 (N_10788,N_6804,N_9765);
nand U10789 (N_10789,N_8560,N_7891);
or U10790 (N_10790,N_7888,N_6357);
nor U10791 (N_10791,N_6517,N_5207);
nor U10792 (N_10792,N_7880,N_7319);
and U10793 (N_10793,N_5276,N_8602);
nor U10794 (N_10794,N_9603,N_7786);
or U10795 (N_10795,N_5752,N_6090);
nor U10796 (N_10796,N_5154,N_7296);
nor U10797 (N_10797,N_6320,N_9280);
and U10798 (N_10798,N_8402,N_7483);
and U10799 (N_10799,N_6836,N_9727);
nand U10800 (N_10800,N_9079,N_8870);
and U10801 (N_10801,N_5520,N_9033);
nor U10802 (N_10802,N_9223,N_7686);
nand U10803 (N_10803,N_8546,N_5493);
nor U10804 (N_10804,N_8005,N_8776);
or U10805 (N_10805,N_6472,N_7854);
or U10806 (N_10806,N_9434,N_6335);
and U10807 (N_10807,N_6296,N_5916);
and U10808 (N_10808,N_7963,N_8591);
and U10809 (N_10809,N_8121,N_5205);
nor U10810 (N_10810,N_9058,N_9369);
or U10811 (N_10811,N_6604,N_6520);
nor U10812 (N_10812,N_8078,N_5248);
and U10813 (N_10813,N_6888,N_9590);
nor U10814 (N_10814,N_8293,N_5917);
nand U10815 (N_10815,N_9755,N_9618);
nor U10816 (N_10816,N_6824,N_8138);
nand U10817 (N_10817,N_8404,N_8700);
and U10818 (N_10818,N_6743,N_8516);
or U10819 (N_10819,N_9211,N_5562);
or U10820 (N_10820,N_6642,N_5863);
nand U10821 (N_10821,N_8204,N_5823);
nand U10822 (N_10822,N_5635,N_5054);
and U10823 (N_10823,N_8713,N_8907);
and U10824 (N_10824,N_7726,N_5569);
or U10825 (N_10825,N_7462,N_5753);
and U10826 (N_10826,N_5930,N_5316);
or U10827 (N_10827,N_6723,N_6618);
and U10828 (N_10828,N_8417,N_6992);
and U10829 (N_10829,N_8211,N_9028);
and U10830 (N_10830,N_5568,N_6197);
nand U10831 (N_10831,N_8082,N_6013);
or U10832 (N_10832,N_6647,N_5099);
nor U10833 (N_10833,N_7326,N_5694);
or U10834 (N_10834,N_9478,N_8731);
or U10835 (N_10835,N_9625,N_6035);
nand U10836 (N_10836,N_9847,N_9514);
and U10837 (N_10837,N_8871,N_5332);
xnor U10838 (N_10838,N_7320,N_8123);
and U10839 (N_10839,N_7499,N_8008);
or U10840 (N_10840,N_5862,N_5377);
xor U10841 (N_10841,N_6557,N_5047);
nand U10842 (N_10842,N_6226,N_5106);
xor U10843 (N_10843,N_7713,N_9406);
and U10844 (N_10844,N_8297,N_7113);
nand U10845 (N_10845,N_7609,N_7361);
or U10846 (N_10846,N_8879,N_9541);
and U10847 (N_10847,N_5538,N_9586);
nor U10848 (N_10848,N_6366,N_8007);
nand U10849 (N_10849,N_6171,N_6868);
or U10850 (N_10850,N_6213,N_8365);
nor U10851 (N_10851,N_8042,N_5576);
nand U10852 (N_10852,N_5896,N_7381);
nor U10853 (N_10853,N_6033,N_6430);
or U10854 (N_10854,N_9632,N_5307);
or U10855 (N_10855,N_7810,N_9000);
and U10856 (N_10856,N_6792,N_8056);
xor U10857 (N_10857,N_6739,N_9393);
and U10858 (N_10858,N_9613,N_5268);
nor U10859 (N_10859,N_5170,N_9887);
or U10860 (N_10860,N_5050,N_9340);
nand U10861 (N_10861,N_5612,N_6554);
nor U10862 (N_10862,N_5030,N_9282);
nand U10863 (N_10863,N_7789,N_7836);
and U10864 (N_10864,N_7181,N_8692);
nor U10865 (N_10865,N_8724,N_8374);
or U10866 (N_10866,N_6462,N_6567);
or U10867 (N_10867,N_5296,N_5271);
and U10868 (N_10868,N_5495,N_7259);
nor U10869 (N_10869,N_7052,N_5293);
or U10870 (N_10870,N_5867,N_5924);
or U10871 (N_10871,N_8060,N_5278);
nand U10872 (N_10872,N_8122,N_7884);
xnor U10873 (N_10873,N_6217,N_7707);
or U10874 (N_10874,N_7490,N_5719);
and U10875 (N_10875,N_6019,N_9975);
or U10876 (N_10876,N_5671,N_7570);
nor U10877 (N_10877,N_6433,N_5487);
or U10878 (N_10878,N_6297,N_9190);
and U10879 (N_10879,N_7056,N_9838);
nand U10880 (N_10880,N_8671,N_8284);
or U10881 (N_10881,N_5703,N_8369);
nand U10882 (N_10882,N_5688,N_6651);
nor U10883 (N_10883,N_7377,N_5082);
nor U10884 (N_10884,N_6309,N_5683);
and U10885 (N_10885,N_6447,N_5548);
nand U10886 (N_10886,N_6914,N_7316);
or U10887 (N_10887,N_9297,N_7083);
or U10888 (N_10888,N_9134,N_6872);
and U10889 (N_10889,N_6970,N_5521);
nor U10890 (N_10890,N_6692,N_8460);
nor U10891 (N_10891,N_6675,N_8557);
or U10892 (N_10892,N_7273,N_9137);
or U10893 (N_10893,N_5839,N_8188);
nand U10894 (N_10894,N_9292,N_9635);
and U10895 (N_10895,N_9217,N_7064);
and U10896 (N_10896,N_8939,N_9189);
and U10897 (N_10897,N_8906,N_7486);
or U10898 (N_10898,N_7443,N_8165);
nor U10899 (N_10899,N_5292,N_7311);
nor U10900 (N_10900,N_7229,N_7680);
nand U10901 (N_10901,N_9372,N_6797);
nor U10902 (N_10902,N_7565,N_7771);
nor U10903 (N_10903,N_6821,N_6531);
or U10904 (N_10904,N_9128,N_9716);
nor U10905 (N_10905,N_7459,N_9861);
and U10906 (N_10906,N_8521,N_6688);
nor U10907 (N_10907,N_7479,N_5871);
nor U10908 (N_10908,N_7790,N_8117);
nor U10909 (N_10909,N_5668,N_9993);
or U10910 (N_10910,N_6185,N_6632);
nand U10911 (N_10911,N_9968,N_5483);
or U10912 (N_10912,N_8595,N_8994);
nand U10913 (N_10913,N_6947,N_9725);
nand U10914 (N_10914,N_9437,N_9316);
or U10915 (N_10915,N_9099,N_7812);
or U10916 (N_10916,N_6215,N_9761);
or U10917 (N_10917,N_8946,N_7365);
and U10918 (N_10918,N_5655,N_6608);
and U10919 (N_10919,N_9815,N_8769);
and U10920 (N_10920,N_6811,N_7842);
nor U10921 (N_10921,N_8251,N_6773);
and U10922 (N_10922,N_9856,N_6887);
or U10923 (N_10923,N_5904,N_7476);
nor U10924 (N_10924,N_8399,N_6285);
nor U10925 (N_10925,N_6638,N_8075);
nor U10926 (N_10926,N_9350,N_9740);
nand U10927 (N_10927,N_9220,N_7310);
nand U10928 (N_10928,N_9472,N_8669);
nor U10929 (N_10929,N_6061,N_6438);
and U10930 (N_10930,N_6816,N_9264);
nand U10931 (N_10931,N_8987,N_5490);
nand U10932 (N_10932,N_9327,N_5578);
and U10933 (N_10933,N_9754,N_9299);
nand U10934 (N_10934,N_5500,N_6350);
nand U10935 (N_10935,N_6349,N_5741);
and U10936 (N_10936,N_6547,N_9477);
or U10937 (N_10937,N_8771,N_7612);
nor U10938 (N_10938,N_5028,N_8583);
nand U10939 (N_10939,N_5782,N_5892);
nand U10940 (N_10940,N_6332,N_5183);
nand U10941 (N_10941,N_5886,N_6645);
and U10942 (N_10942,N_7711,N_5172);
nand U10943 (N_10943,N_8718,N_5295);
nand U10944 (N_10944,N_9193,N_8749);
nand U10945 (N_10945,N_9594,N_7544);
nand U10946 (N_10946,N_6109,N_6007);
and U10947 (N_10947,N_7737,N_5390);
and U10948 (N_10948,N_8860,N_7069);
or U10949 (N_10949,N_8537,N_6658);
or U10950 (N_10950,N_5954,N_9793);
nand U10951 (N_10951,N_7182,N_7350);
and U10952 (N_10952,N_5130,N_8029);
or U10953 (N_10953,N_7822,N_8367);
and U10954 (N_10954,N_5000,N_7226);
nand U10955 (N_10955,N_9431,N_6640);
and U10956 (N_10956,N_7358,N_8639);
or U10957 (N_10957,N_6755,N_5801);
nand U10958 (N_10958,N_6321,N_6954);
or U10959 (N_10959,N_8432,N_7766);
and U10960 (N_10960,N_9408,N_8750);
nor U10961 (N_10961,N_7153,N_5436);
or U10962 (N_10962,N_9679,N_9331);
or U10963 (N_10963,N_7589,N_9976);
nand U10964 (N_10964,N_5422,N_5408);
or U10965 (N_10965,N_5622,N_8244);
nand U10966 (N_10966,N_5398,N_9364);
and U10967 (N_10967,N_7292,N_6865);
and U10968 (N_10968,N_7295,N_8080);
nor U10969 (N_10969,N_7080,N_6403);
and U10970 (N_10970,N_7424,N_8911);
nor U10971 (N_10971,N_6793,N_6611);
and U10972 (N_10972,N_6442,N_9662);
nor U10973 (N_10973,N_6329,N_8448);
nor U10974 (N_10974,N_9422,N_5464);
or U10975 (N_10975,N_7823,N_7351);
and U10976 (N_10976,N_6252,N_6020);
nor U10977 (N_10977,N_5164,N_5728);
nor U10978 (N_10978,N_8739,N_9811);
and U10979 (N_10979,N_7920,N_8372);
and U10980 (N_10980,N_7855,N_6972);
nand U10981 (N_10981,N_9549,N_5196);
and U10982 (N_10982,N_9920,N_6760);
nor U10983 (N_10983,N_5632,N_8938);
and U10984 (N_10984,N_5556,N_9130);
nand U10985 (N_10985,N_9439,N_7539);
and U10986 (N_10986,N_8313,N_7732);
nand U10987 (N_10987,N_6812,N_7864);
nand U10988 (N_10988,N_5494,N_8319);
and U10989 (N_10989,N_5901,N_7213);
nand U10990 (N_10990,N_8357,N_7385);
nand U10991 (N_10991,N_9521,N_8922);
nor U10992 (N_10992,N_7477,N_5648);
nand U10993 (N_10993,N_5025,N_5261);
and U10994 (N_10994,N_9676,N_8694);
nand U10995 (N_10995,N_7952,N_6314);
and U10996 (N_10996,N_7282,N_6441);
nor U10997 (N_10997,N_7558,N_6159);
nand U10998 (N_10998,N_6220,N_6730);
nand U10999 (N_10999,N_9479,N_8418);
nand U11000 (N_11000,N_5905,N_5372);
or U11001 (N_11001,N_9928,N_6712);
or U11002 (N_11002,N_9295,N_9708);
and U11003 (N_11003,N_9009,N_7161);
and U11004 (N_11004,N_7698,N_7471);
and U11005 (N_11005,N_7349,N_7905);
and U11006 (N_11006,N_7601,N_6806);
nor U11007 (N_11007,N_9834,N_5175);
nor U11008 (N_11008,N_8496,N_8476);
or U11009 (N_11009,N_7025,N_6318);
nor U11010 (N_11010,N_7911,N_9345);
nor U11011 (N_11011,N_8242,N_7104);
or U11012 (N_11012,N_9995,N_8572);
nor U11013 (N_11013,N_9756,N_9664);
nor U11014 (N_11014,N_8253,N_5761);
or U11015 (N_11015,N_5641,N_6038);
nand U11016 (N_11016,N_5602,N_9734);
nor U11017 (N_11017,N_7194,N_5932);
nand U11018 (N_11018,N_5356,N_5914);
nand U11019 (N_11019,N_8185,N_5137);
or U11020 (N_11020,N_9665,N_7996);
and U11021 (N_11021,N_5933,N_7820);
nor U11022 (N_11022,N_7578,N_5712);
nor U11023 (N_11023,N_8232,N_8194);
and U11024 (N_11024,N_9136,N_5593);
or U11025 (N_11025,N_9117,N_6513);
nor U11026 (N_11026,N_5524,N_8470);
xnor U11027 (N_11027,N_6227,N_7718);
nand U11028 (N_11028,N_7639,N_8530);
nand U11029 (N_11029,N_5962,N_9098);
or U11030 (N_11030,N_5070,N_7793);
nor U11031 (N_11031,N_8145,N_6089);
nand U11032 (N_11032,N_9474,N_8411);
and U11033 (N_11033,N_5563,N_9417);
or U11034 (N_11034,N_6370,N_5730);
or U11035 (N_11035,N_5725,N_8248);
nor U11036 (N_11036,N_9567,N_7084);
and U11037 (N_11037,N_5341,N_8224);
and U11038 (N_11038,N_5796,N_6905);
or U11039 (N_11039,N_6310,N_6928);
or U11040 (N_11040,N_6015,N_7002);
and U11041 (N_11041,N_9042,N_7591);
nor U11042 (N_11042,N_8919,N_7611);
and U11043 (N_11043,N_7019,N_8462);
or U11044 (N_11044,N_8241,N_8289);
nor U11045 (N_11045,N_5869,N_5096);
or U11046 (N_11046,N_7688,N_5518);
and U11047 (N_11047,N_5617,N_5729);
and U11048 (N_11048,N_9774,N_7455);
and U11049 (N_11049,N_8971,N_8237);
nand U11050 (N_11050,N_7028,N_8978);
nor U11051 (N_11051,N_7536,N_7102);
nand U11052 (N_11052,N_5188,N_9839);
nor U11053 (N_11053,N_8554,N_9899);
nand U11054 (N_11054,N_8283,N_6322);
and U11055 (N_11055,N_8957,N_9066);
nor U11056 (N_11056,N_7355,N_5311);
and U11057 (N_11057,N_5953,N_5144);
nor U11058 (N_11058,N_9742,N_6835);
and U11059 (N_11059,N_7399,N_5894);
nor U11060 (N_11060,N_8381,N_7059);
nor U11061 (N_11061,N_7021,N_7065);
or U11062 (N_11062,N_8610,N_9689);
and U11063 (N_11063,N_9580,N_5860);
or U11064 (N_11064,N_5580,N_8186);
nor U11065 (N_11065,N_5958,N_5722);
nor U11066 (N_11066,N_5779,N_7287);
nand U11067 (N_11067,N_9467,N_8913);
or U11068 (N_11068,N_5083,N_7111);
or U11069 (N_11069,N_7788,N_9912);
and U11070 (N_11070,N_6401,N_8425);
xor U11071 (N_11071,N_5553,N_6180);
and U11072 (N_11072,N_8485,N_5508);
or U11073 (N_11073,N_7261,N_9326);
and U11074 (N_11074,N_7749,N_7840);
or U11075 (N_11075,N_9588,N_8300);
nor U11076 (N_11076,N_6583,N_9548);
nor U11077 (N_11077,N_8066,N_6633);
nand U11078 (N_11078,N_6120,N_8941);
or U11079 (N_11079,N_7660,N_5743);
nor U11080 (N_11080,N_9639,N_9902);
and U11081 (N_11081,N_8581,N_6748);
and U11082 (N_11082,N_7647,N_7264);
or U11083 (N_11083,N_9139,N_5222);
or U11084 (N_11084,N_6280,N_9733);
nand U11085 (N_11085,N_8219,N_8921);
and U11086 (N_11086,N_5783,N_5334);
and U11087 (N_11087,N_6802,N_6153);
and U11088 (N_11088,N_8933,N_9154);
nand U11089 (N_11089,N_8961,N_8146);
nor U11090 (N_11090,N_8637,N_5414);
or U11091 (N_11091,N_8588,N_5527);
nand U11092 (N_11092,N_5906,N_9109);
and U11093 (N_11093,N_6176,N_6369);
nor U11094 (N_11094,N_7309,N_6491);
or U11095 (N_11095,N_5718,N_5091);
nand U11096 (N_11096,N_5666,N_5528);
and U11097 (N_11097,N_5055,N_5775);
and U11098 (N_11098,N_7063,N_5994);
nor U11099 (N_11099,N_5445,N_8523);
nor U11100 (N_11100,N_5383,N_5874);
nand U11101 (N_11101,N_7497,N_7180);
and U11102 (N_11102,N_8779,N_9550);
or U11103 (N_11103,N_7930,N_6613);
nor U11104 (N_11104,N_8866,N_8090);
xor U11105 (N_11105,N_7225,N_6918);
or U11106 (N_11106,N_5566,N_9184);
nand U11107 (N_11107,N_6243,N_5988);
nor U11108 (N_11108,N_7943,N_8482);
and U11109 (N_11109,N_8586,N_6027);
and U11110 (N_11110,N_5968,N_5890);
or U11111 (N_11111,N_7700,N_6105);
or U11112 (N_11112,N_7955,N_7357);
or U11113 (N_11113,N_7803,N_7721);
or U11114 (N_11114,N_9537,N_7804);
nor U11115 (N_11115,N_8667,N_6413);
nand U11116 (N_11116,N_7423,N_5392);
nand U11117 (N_11117,N_5382,N_7401);
nor U11118 (N_11118,N_6270,N_7736);
nor U11119 (N_11119,N_8081,N_7623);
nor U11120 (N_11120,N_5005,N_5088);
nand U11121 (N_11121,N_9533,N_8193);
or U11122 (N_11122,N_7959,N_7207);
or U11123 (N_11123,N_7015,N_8058);
nor U11124 (N_11124,N_8336,N_9644);
nor U11125 (N_11125,N_7714,N_5685);
nor U11126 (N_11126,N_8004,N_7635);
or U11127 (N_11127,N_5421,N_6371);
and U11128 (N_11128,N_9554,N_9919);
nor U11129 (N_11129,N_7145,N_8954);
nand U11130 (N_11130,N_5608,N_5122);
nand U11131 (N_11131,N_9370,N_6127);
nand U11132 (N_11132,N_8011,N_7873);
nor U11133 (N_11133,N_8213,N_8071);
or U11134 (N_11134,N_6774,N_9332);
nor U11135 (N_11135,N_9770,N_9101);
nand U11136 (N_11136,N_9579,N_9578);
nand U11137 (N_11137,N_9753,N_6481);
nor U11138 (N_11138,N_5290,N_7057);
or U11139 (N_11139,N_8687,N_8209);
nand U11140 (N_11140,N_6128,N_8261);
and U11141 (N_11141,N_6837,N_8538);
nand U11142 (N_11142,N_5463,N_9142);
and U11143 (N_11143,N_5121,N_8410);
nand U11144 (N_11144,N_9160,N_8986);
nor U11145 (N_11145,N_5475,N_5582);
nand U11146 (N_11146,N_9207,N_7022);
nor U11147 (N_11147,N_5317,N_8514);
xnor U11148 (N_11148,N_6819,N_9785);
nor U11149 (N_11149,N_6716,N_8451);
and U11150 (N_11150,N_5710,N_8599);
or U11151 (N_11151,N_9044,N_8223);
nand U11152 (N_11152,N_7858,N_5333);
nor U11153 (N_11153,N_9880,N_9745);
and U11154 (N_11154,N_5881,N_5879);
or U11155 (N_11155,N_7014,N_6858);
and U11156 (N_11156,N_6593,N_5374);
or U11157 (N_11157,N_5203,N_6428);
xnor U11158 (N_11158,N_5460,N_6494);
and U11159 (N_11159,N_6135,N_8269);
or U11160 (N_11160,N_9071,N_7008);
xor U11161 (N_11161,N_9480,N_6997);
nand U11162 (N_11162,N_6306,N_9324);
and U11163 (N_11163,N_7465,N_6096);
or U11164 (N_11164,N_9819,N_8819);
nand U11165 (N_11165,N_8820,N_8040);
and U11166 (N_11166,N_5764,N_6526);
or U11167 (N_11167,N_8163,N_5654);
nand U11168 (N_11168,N_6989,N_8129);
nand U11169 (N_11169,N_7148,N_7542);
nor U11170 (N_11170,N_8429,N_5807);
nor U11171 (N_11171,N_6906,N_6206);
nor U11172 (N_11172,N_5934,N_6141);
and U11173 (N_11173,N_5387,N_6542);
nand U11174 (N_11174,N_5902,N_7867);
nor U11175 (N_11175,N_6014,N_6889);
or U11176 (N_11176,N_8208,N_6126);
nor U11177 (N_11177,N_5929,N_6781);
and U11178 (N_11178,N_5102,N_8002);
and U11179 (N_11179,N_5634,N_8770);
xnor U11180 (N_11180,N_5693,N_9133);
and U11181 (N_11181,N_6650,N_6387);
and U11182 (N_11182,N_8822,N_9401);
nand U11183 (N_11183,N_8398,N_8230);
nor U11184 (N_11184,N_6142,N_8420);
and U11185 (N_11185,N_5687,N_5146);
and U11186 (N_11186,N_7874,N_6545);
or U11187 (N_11187,N_8969,N_5449);
nand U11188 (N_11188,N_6986,N_5197);
nor U11189 (N_11189,N_6340,N_6680);
nand U11190 (N_11190,N_7422,N_5797);
and U11191 (N_11191,N_8507,N_7086);
and U11192 (N_11192,N_8287,N_7206);
or U11193 (N_11193,N_6843,N_9414);
and U11194 (N_11194,N_6319,N_5127);
nand U11195 (N_11195,N_7050,N_7850);
or U11196 (N_11196,N_6782,N_5789);
or U11197 (N_11197,N_9291,N_7389);
and U11198 (N_11198,N_6825,N_5503);
nor U11199 (N_11199,N_8741,N_8766);
nand U11200 (N_11200,N_8423,N_6710);
or U11201 (N_11201,N_9398,N_5833);
nand U11202 (N_11202,N_8214,N_9804);
nor U11203 (N_11203,N_7033,N_9277);
nor U11204 (N_11204,N_8629,N_8112);
nor U11205 (N_11205,N_9595,N_9789);
or U11206 (N_11206,N_9228,N_9984);
nor U11207 (N_11207,N_9619,N_8963);
and U11208 (N_11208,N_5448,N_7754);
and U11209 (N_11209,N_5996,N_5442);
and U11210 (N_11210,N_8702,N_5824);
or U11211 (N_11211,N_6052,N_7787);
nor U11212 (N_11212,N_7210,N_9693);
or U11213 (N_11213,N_8804,N_7125);
or U11214 (N_11214,N_8182,N_8166);
nor U11215 (N_11215,N_9737,N_5755);
and U11216 (N_11216,N_8061,N_5174);
or U11217 (N_11217,N_6173,N_7599);
nor U11218 (N_11218,N_5826,N_7760);
or U11219 (N_11219,N_9516,N_5937);
nor U11220 (N_11220,N_9686,N_8966);
and U11221 (N_11221,N_9162,N_6728);
nor U11222 (N_11222,N_5165,N_8773);
and U11223 (N_11223,N_9589,N_6083);
nor U11224 (N_11224,N_7370,N_5773);
nand U11225 (N_11225,N_9832,N_8373);
or U11226 (N_11226,N_7314,N_8606);
nand U11227 (N_11227,N_8658,N_7725);
nand U11228 (N_11228,N_6535,N_7597);
and U11229 (N_11229,N_9403,N_6749);
nor U11230 (N_11230,N_8716,N_9185);
and U11231 (N_11231,N_5535,N_9178);
or U11232 (N_11232,N_6283,N_9671);
and U11233 (N_11233,N_6452,N_8074);
and U11234 (N_11234,N_9395,N_5068);
and U11235 (N_11235,N_8652,N_7418);
and U11236 (N_11236,N_7364,N_9681);
nand U11237 (N_11237,N_7478,N_8016);
nand U11238 (N_11238,N_8968,N_7535);
nor U11239 (N_11239,N_9666,N_8976);
nand U11240 (N_11240,N_6022,N_9337);
and U11241 (N_11241,N_5470,N_9906);
xor U11242 (N_11242,N_9904,N_9828);
nand U11243 (N_11243,N_6968,N_8518);
nor U11244 (N_11244,N_6704,N_9901);
and U11245 (N_11245,N_9915,N_8382);
nor U11246 (N_11246,N_8918,N_8258);
and U11247 (N_11247,N_6398,N_7616);
nand U11248 (N_11248,N_5370,N_9855);
and U11249 (N_11249,N_6724,N_7659);
nor U11250 (N_11250,N_5840,N_9095);
nand U11251 (N_11251,N_8015,N_6073);
or U11252 (N_11252,N_8221,N_5944);
or U11253 (N_11253,N_7948,N_6703);
nand U11254 (N_11254,N_8947,N_7016);
nor U11255 (N_11255,N_9241,N_8944);
nor U11256 (N_11256,N_9741,N_6540);
or U11257 (N_11257,N_7801,N_5496);
and U11258 (N_11258,N_7869,N_8828);
nor U11259 (N_11259,N_6288,N_6338);
nor U11260 (N_11260,N_9269,N_8707);
nand U11261 (N_11261,N_9925,N_6713);
and U11262 (N_11262,N_7666,N_7100);
nand U11263 (N_11263,N_9248,N_9123);
nor U11264 (N_11264,N_8150,N_5412);
and U11265 (N_11265,N_8513,N_9705);
nor U11266 (N_11266,N_5804,N_8857);
nor U11267 (N_11267,N_7048,N_6326);
and U11268 (N_11268,N_9454,N_5477);
or U11269 (N_11269,N_9786,N_5302);
nand U11270 (N_11270,N_9738,N_6079);
and U11271 (N_11271,N_7605,N_6848);
or U11272 (N_11272,N_5732,N_7941);
nor U11273 (N_11273,N_9306,N_8239);
or U11274 (N_11274,N_8205,N_6920);
or U11275 (N_11275,N_6016,N_9735);
nand U11276 (N_11276,N_9624,N_7767);
or U11277 (N_11277,N_9400,N_5575);
nor U11278 (N_11278,N_6255,N_8604);
and U11279 (N_11279,N_9830,N_8528);
nor U11280 (N_11280,N_9065,N_9328);
and U11281 (N_11281,N_5472,N_7409);
xor U11282 (N_11282,N_7457,N_8325);
nand U11283 (N_11283,N_8525,N_8803);
nand U11284 (N_11284,N_5478,N_9153);
nand U11285 (N_11285,N_9383,N_9885);
xor U11286 (N_11286,N_6898,N_6578);
nor U11287 (N_11287,N_8318,N_7527);
nand U11288 (N_11288,N_7569,N_8989);
and U11289 (N_11289,N_6732,N_7238);
nand U11290 (N_11290,N_7621,N_6916);
nand U11291 (N_11291,N_8623,N_5236);
nor U11292 (N_11292,N_9484,N_5409);
or U11293 (N_11293,N_7890,N_9290);
or U11294 (N_11294,N_7288,N_8200);
and U11295 (N_11295,N_7935,N_8791);
nor U11296 (N_11296,N_6586,N_5533);
nand U11297 (N_11297,N_8358,N_8228);
xor U11298 (N_11298,N_5241,N_6588);
or U11299 (N_11299,N_8977,N_6356);
or U11300 (N_11300,N_5657,N_7093);
and U11301 (N_11301,N_9460,N_8972);
nand U11302 (N_11302,N_7475,N_7126);
nor U11303 (N_11303,N_7304,N_5168);
nand U11304 (N_11304,N_6048,N_9842);
and U11305 (N_11305,N_6570,N_8315);
nand U11306 (N_11306,N_7661,N_8453);
and U11307 (N_11307,N_9433,N_5726);
nand U11308 (N_11308,N_5785,N_7831);
nand U11309 (N_11309,N_5550,N_8125);
nand U11310 (N_11310,N_7516,N_5945);
nand U11311 (N_11311,N_9273,N_7234);
nor U11312 (N_11312,N_8275,N_6304);
or U11313 (N_11313,N_8708,N_5116);
and U11314 (N_11314,N_6429,N_5095);
and U11315 (N_11315,N_9506,N_8178);
nand U11316 (N_11316,N_9049,N_8449);
and U11317 (N_11317,N_6042,N_8556);
and U11318 (N_11318,N_5665,N_7665);
and U11319 (N_11319,N_6260,N_9385);
nor U11320 (N_11320,N_7392,N_7965);
and U11321 (N_11321,N_7258,N_7553);
and U11322 (N_11322,N_7184,N_5405);
nor U11323 (N_11323,N_8559,N_7338);
and U11324 (N_11324,N_6630,N_6381);
or U11325 (N_11325,N_6736,N_6569);
and U11326 (N_11326,N_6685,N_6264);
nor U11327 (N_11327,N_8901,N_5875);
and U11328 (N_11328,N_6656,N_9376);
nor U11329 (N_11329,N_9913,N_9394);
nand U11330 (N_11330,N_7791,N_6622);
or U11331 (N_11331,N_8252,N_7796);
nor U11332 (N_11332,N_6715,N_5043);
nand U11333 (N_11333,N_8711,N_9143);
and U11334 (N_11334,N_7995,N_8817);
or U11335 (N_11335,N_5403,N_9257);
nand U11336 (N_11336,N_8617,N_5966);
nand U11337 (N_11337,N_7703,N_9051);
nor U11338 (N_11338,N_9700,N_5706);
nand U11339 (N_11339,N_5224,N_5923);
and U11340 (N_11340,N_9038,N_9731);
nor U11341 (N_11341,N_8914,N_6500);
nor U11342 (N_11342,N_8105,N_8758);
nor U11343 (N_11343,N_6944,N_9118);
or U11344 (N_11344,N_6422,N_5038);
and U11345 (N_11345,N_8431,N_8001);
nand U11346 (N_11346,N_6181,N_9152);
nand U11347 (N_11347,N_6592,N_8624);
nor U11348 (N_11348,N_5314,N_5735);
and U11349 (N_11349,N_5162,N_6088);
nand U11350 (N_11350,N_7165,N_6893);
nor U11351 (N_11351,N_6823,N_7030);
or U11352 (N_11352,N_6174,N_7405);
nand U11353 (N_11353,N_5258,N_7978);
nor U11354 (N_11354,N_6719,N_8017);
nor U11355 (N_11355,N_7636,N_8181);
nor U11356 (N_11356,N_6841,N_6768);
and U11357 (N_11357,N_8375,N_5604);
and U11358 (N_11358,N_9018,N_7388);
or U11359 (N_11359,N_7928,N_8049);
nor U11360 (N_11360,N_9432,N_8760);
nor U11361 (N_11361,N_9367,N_8397);
nand U11362 (N_11362,N_7217,N_7683);
nor U11363 (N_11363,N_5040,N_9442);
nand U11364 (N_11364,N_6850,N_8203);
nand U11365 (N_11365,N_5745,N_9481);
and U11366 (N_11366,N_9893,N_6572);
nor U11367 (N_11367,N_9234,N_6269);
nor U11368 (N_11368,N_9528,N_9329);
or U11369 (N_11369,N_5623,N_5018);
nand U11370 (N_11370,N_7023,N_9413);
or U11371 (N_11371,N_6364,N_7012);
nor U11372 (N_11372,N_6469,N_7436);
and U11373 (N_11373,N_9219,N_6044);
nor U11374 (N_11374,N_8020,N_5281);
and U11375 (N_11375,N_6951,N_6261);
nor U11376 (N_11376,N_6686,N_8218);
nand U11377 (N_11377,N_8147,N_9093);
and U11378 (N_11378,N_6523,N_5118);
nor U11379 (N_11379,N_8829,N_7450);
nor U11380 (N_11380,N_6488,N_8442);
and U11381 (N_11381,N_8441,N_6838);
xnor U11382 (N_11382,N_6199,N_5772);
or U11383 (N_11383,N_8801,N_5615);
nor U11384 (N_11384,N_8619,N_6192);
nor U11385 (N_11385,N_5406,N_5253);
nand U11386 (N_11386,N_7853,N_9202);
and U11387 (N_11387,N_9216,N_7456);
and U11388 (N_11388,N_9070,N_6140);
nand U11389 (N_11389,N_5466,N_8725);
or U11390 (N_11390,N_6585,N_5266);
nor U11391 (N_11391,N_7330,N_6054);
and U11392 (N_11392,N_8789,N_5024);
nand U11393 (N_11393,N_7849,N_7646);
and U11394 (N_11394,N_5845,N_5274);
nand U11395 (N_11395,N_6896,N_6386);
or U11396 (N_11396,N_9020,N_9347);
and U11397 (N_11397,N_9250,N_6464);
nor U11398 (N_11398,N_9121,N_7248);
nor U11399 (N_11399,N_9760,N_9535);
nor U11400 (N_11400,N_5973,N_5256);
nor U11401 (N_11401,N_5204,N_6098);
or U11402 (N_11402,N_5949,N_8053);
or U11403 (N_11403,N_5770,N_9979);
nor U11404 (N_11404,N_9194,N_6479);
or U11405 (N_11405,N_6388,N_9998);
nand U11406 (N_11406,N_7733,N_7933);
and U11407 (N_11407,N_8190,N_6122);
nor U11408 (N_11408,N_7805,N_6969);
or U11409 (N_11409,N_8821,N_5338);
or U11410 (N_11410,N_6426,N_8684);
xor U11411 (N_11411,N_9945,N_5596);
nand U11412 (N_11412,N_9302,N_6845);
nor U11413 (N_11413,N_9955,N_9767);
nor U11414 (N_11414,N_8747,N_6341);
nand U11415 (N_11415,N_8967,N_7983);
and U11416 (N_11416,N_5459,N_7586);
nand U11417 (N_11417,N_8409,N_9691);
and U11418 (N_11418,N_8118,N_5889);
and U11419 (N_11419,N_5852,N_7268);
and U11420 (N_11420,N_7904,N_9313);
and U11421 (N_11421,N_6877,N_8207);
and U11422 (N_11422,N_8345,N_7602);
and U11423 (N_11423,N_8352,N_7818);
or U11424 (N_11424,N_6046,N_7835);
xnor U11425 (N_11425,N_8435,N_9011);
xnor U11426 (N_11426,N_7176,N_9539);
and U11427 (N_11427,N_6342,N_6354);
nor U11428 (N_11428,N_5467,N_9037);
nor U11429 (N_11429,N_9305,N_6389);
and U11430 (N_11430,N_5286,N_7105);
and U11431 (N_11431,N_5540,N_7650);
nor U11432 (N_11432,N_5060,N_8133);
nand U11433 (N_11433,N_7582,N_8396);
or U11434 (N_11434,N_8551,N_6184);
nand U11435 (N_11435,N_6499,N_6839);
and U11436 (N_11436,N_9151,N_7429);
nor U11437 (N_11437,N_8793,N_8737);
nor U11438 (N_11438,N_8563,N_7808);
nor U11439 (N_11439,N_5909,N_8597);
nor U11440 (N_11440,N_5214,N_6827);
or U11441 (N_11441,N_7641,N_6155);
or U11442 (N_11442,N_6344,N_9192);
nand U11443 (N_11443,N_9890,N_9648);
and U11444 (N_11444,N_6119,N_7136);
and U11445 (N_11445,N_8051,N_8612);
nand U11446 (N_11446,N_7271,N_6873);
or U11447 (N_11447,N_9026,N_9612);
nor U11448 (N_11448,N_6706,N_7997);
nand U11449 (N_11449,N_9531,N_8975);
or U11450 (N_11450,N_8028,N_6863);
and U11451 (N_11451,N_7329,N_5433);
nand U11452 (N_11452,N_6502,N_5948);
and U11453 (N_11453,N_7454,N_5491);
and U11454 (N_11454,N_8229,N_8764);
or U11455 (N_11455,N_5972,N_5185);
nor U11456 (N_11456,N_7617,N_7412);
nor U11457 (N_11457,N_8109,N_6092);
and U11458 (N_11458,N_5799,N_5865);
or U11459 (N_11459,N_6854,N_7740);
nor U11460 (N_11460,N_9186,N_5428);
or U11461 (N_11461,N_7613,N_7543);
and U11462 (N_11462,N_5016,N_5828);
and U11463 (N_11463,N_9131,N_7284);
nor U11464 (N_11464,N_6669,N_8176);
nand U11465 (N_11465,N_6767,N_6231);
nor U11466 (N_11466,N_9544,N_8444);
nor U11467 (N_11467,N_9520,N_6000);
or U11468 (N_11468,N_8198,N_7630);
xor U11469 (N_11469,N_9766,N_9512);
or U11470 (N_11470,N_5048,N_7664);
or U11471 (N_11471,N_5581,N_8715);
nor U11472 (N_11472,N_8827,N_6085);
or U11473 (N_11473,N_7577,N_8851);
or U11474 (N_11474,N_7953,N_9584);
nand U11475 (N_11475,N_5534,N_7825);
or U11476 (N_11476,N_8688,N_8973);
or U11477 (N_11477,N_6373,N_5136);
nor U11478 (N_11478,N_9684,N_9859);
xor U11479 (N_11479,N_8561,N_9848);
nor U11480 (N_11480,N_7281,N_5597);
or U11481 (N_11481,N_6769,N_9430);
or U11482 (N_11482,N_8421,N_9800);
and U11483 (N_11483,N_5300,N_5572);
and U11484 (N_11484,N_9197,N_8564);
nand U11485 (N_11485,N_6154,N_7743);
nor U11486 (N_11486,N_9659,N_9391);
and U11487 (N_11487,N_7158,N_9251);
nor U11488 (N_11488,N_6742,N_8440);
and U11489 (N_11489,N_8910,N_6450);
nor U11490 (N_11490,N_7129,N_8902);
and U11491 (N_11491,N_7328,N_5599);
and U11492 (N_11492,N_8736,N_7971);
and U11493 (N_11493,N_6869,N_6765);
nand U11494 (N_11494,N_9908,N_7921);
and U11495 (N_11495,N_9964,N_8615);
and U11496 (N_11496,N_8026,N_6721);
nand U11497 (N_11497,N_9021,N_5884);
or U11498 (N_11498,N_8415,N_9198);
nor U11499 (N_11499,N_9967,N_5200);
and U11500 (N_11500,N_8600,N_8993);
and U11501 (N_11501,N_9840,N_6245);
and U11502 (N_11502,N_6362,N_9459);
and U11503 (N_11503,N_7987,N_5425);
nand U11504 (N_11504,N_8236,N_5605);
and U11505 (N_11505,N_5838,N_7545);
nor U11506 (N_11506,N_8501,N_8937);
or U11507 (N_11507,N_7962,N_6694);
and U11508 (N_11508,N_5947,N_5959);
nand U11509 (N_11509,N_5681,N_8259);
nand U11510 (N_11510,N_7485,N_7981);
nor U11511 (N_11511,N_8765,N_9685);
nor U11512 (N_11512,N_9485,N_8493);
or U11513 (N_11513,N_9593,N_8543);
or U11514 (N_11514,N_8601,N_7494);
and U11515 (N_11515,N_7908,N_7876);
nor U11516 (N_11516,N_7533,N_6156);
xor U11517 (N_11517,N_7289,N_5633);
nor U11518 (N_11518,N_7054,N_5859);
and U11519 (N_11519,N_8898,N_9453);
nor U11520 (N_11520,N_5027,N_8626);
nor U11521 (N_11521,N_7430,N_6175);
nor U11522 (N_11522,N_9468,N_9267);
and U11523 (N_11523,N_6300,N_6975);
or U11524 (N_11524,N_8486,N_5613);
or U11525 (N_11525,N_6571,N_9493);
or U11526 (N_11526,N_8492,N_5240);
xor U11527 (N_11527,N_9794,N_7830);
nor U11528 (N_11528,N_8034,N_6746);
and U11529 (N_11529,N_6840,N_6473);
or U11530 (N_11530,N_7511,N_7833);
nor U11531 (N_11531,N_9252,N_7748);
nand U11532 (N_11532,N_6455,N_8262);
xnor U11533 (N_11533,N_6149,N_5163);
or U11534 (N_11534,N_5594,N_8683);
nor U11535 (N_11535,N_8923,N_6418);
and U11536 (N_11536,N_8327,N_8206);
or U11537 (N_11537,N_6068,N_7339);
or U11538 (N_11538,N_9497,N_9787);
or U11539 (N_11539,N_7693,N_6795);
or U11540 (N_11540,N_8656,N_7174);
or U11541 (N_11541,N_9173,N_5644);
or U11542 (N_11542,N_7776,N_5913);
nor U11543 (N_11543,N_5837,N_8477);
xor U11544 (N_11544,N_5209,N_6204);
nor U11545 (N_11545,N_5484,N_8797);
nand U11546 (N_11546,N_5591,N_7240);
or U11547 (N_11547,N_8850,N_7768);
and U11548 (N_11548,N_7678,N_8110);
nand U11549 (N_11549,N_7878,N_9730);
or U11550 (N_11550,N_5653,N_5104);
and U11551 (N_11551,N_6195,N_6974);
and U11552 (N_11552,N_5545,N_7024);
or U11553 (N_11553,N_6648,N_8876);
or U11554 (N_11554,N_6009,N_8234);
nor U11555 (N_11555,N_5324,N_5312);
or U11556 (N_11556,N_7954,N_9441);
nand U11557 (N_11557,N_7534,N_6425);
nor U11558 (N_11558,N_8380,N_5262);
nand U11559 (N_11559,N_5310,N_6754);
nor U11560 (N_11560,N_6960,N_9330);
and U11561 (N_11561,N_6315,N_8114);
or U11562 (N_11562,N_9882,N_8495);
or U11563 (N_11563,N_8059,N_7195);
and U11564 (N_11564,N_6671,N_8896);
and U11565 (N_11565,N_5861,N_9235);
or U11566 (N_11566,N_6663,N_8953);
or U11567 (N_11567,N_6273,N_6518);
or U11568 (N_11568,N_6087,N_8508);
nor U11569 (N_11569,N_8659,N_7584);
or U11570 (N_11570,N_7221,N_6639);
and U11571 (N_11571,N_7775,N_6815);
and U11572 (N_11572,N_7655,N_8106);
and U11573 (N_11573,N_5600,N_8184);
or U11574 (N_11574,N_5750,N_9994);
nand U11575 (N_11575,N_7235,N_8625);
nor U11576 (N_11576,N_7600,N_6427);
nor U11577 (N_11577,N_7735,N_8988);
and U11578 (N_11578,N_8268,N_6324);
or U11579 (N_11579,N_7877,N_8858);
nand U11580 (N_11580,N_6053,N_5119);
nand U11581 (N_11581,N_5150,N_7122);
nand U11582 (N_11582,N_9004,N_8096);
and U11583 (N_11583,N_6695,N_8893);
nand U11584 (N_11584,N_6193,N_9845);
and U11585 (N_11585,N_7894,N_9711);
and U11586 (N_11586,N_9157,N_8900);
xnor U11587 (N_11587,N_9670,N_6487);
nand U11588 (N_11588,N_5559,N_6405);
and U11589 (N_11589,N_9897,N_9641);
and U11590 (N_11590,N_5551,N_6923);
nor U11591 (N_11591,N_9165,N_9701);
or U11592 (N_11592,N_5887,N_9559);
xor U11593 (N_11593,N_5888,N_8088);
and U11594 (N_11594,N_7360,N_9096);
nor U11595 (N_11595,N_7419,N_6758);
nand U11596 (N_11596,N_9965,N_5505);
nand U11597 (N_11597,N_7784,N_5217);
nand U11598 (N_11598,N_7629,N_5492);
or U11599 (N_11599,N_8785,N_9658);
nor U11600 (N_11600,N_8892,N_9784);
and U11601 (N_11601,N_7555,N_5790);
or U11602 (N_11602,N_6290,N_8316);
nor U11603 (N_11603,N_8245,N_5991);
xnor U11604 (N_11604,N_8575,N_6594);
nand U11605 (N_11605,N_9782,N_8648);
and U11606 (N_11606,N_5285,N_8497);
nor U11607 (N_11607,N_5984,N_8956);
or U11608 (N_11608,N_5111,N_9014);
and U11609 (N_11609,N_8107,N_5046);
and U11610 (N_11610,N_6574,N_9690);
xor U11611 (N_11611,N_7116,N_7431);
nand U11612 (N_11612,N_7919,N_5321);
nand U11613 (N_11613,N_5803,N_6143);
nand U11614 (N_11614,N_7152,N_6397);
or U11615 (N_11615,N_7679,N_5342);
nand U11616 (N_11616,N_6772,N_7218);
and U11617 (N_11617,N_8471,N_8699);
nand U11618 (N_11618,N_9253,N_8755);
nand U11619 (N_11619,N_5186,N_5215);
or U11620 (N_11620,N_7752,N_8931);
or U11621 (N_11621,N_7384,N_8348);
nand U11622 (N_11622,N_5004,N_8809);
and U11623 (N_11623,N_7452,N_7004);
or U11624 (N_11624,N_5007,N_8338);
and U11625 (N_11625,N_9397,N_9713);
nand U11626 (N_11626,N_6649,N_6144);
or U11627 (N_11627,N_7969,N_8304);
or U11628 (N_11628,N_7255,N_7196);
nand U11629 (N_11629,N_8783,N_8290);
nand U11630 (N_11630,N_8189,N_7081);
nor U11631 (N_11631,N_8077,N_5303);
nand U11632 (N_11632,N_5664,N_7780);
nand U11633 (N_11633,N_9607,N_8151);
nand U11634 (N_11634,N_5351,N_7556);
and U11635 (N_11635,N_9392,N_6566);
or U11636 (N_11636,N_7903,N_6029);
or U11637 (N_11637,N_5159,N_7242);
nor U11638 (N_11638,N_7190,N_7178);
and U11639 (N_11639,N_5956,N_5469);
nand U11640 (N_11640,N_7166,N_5649);
and U11641 (N_11641,N_6470,N_7638);
nor U11642 (N_11642,N_5456,N_9611);
xor U11643 (N_11643,N_5637,N_6660);
and U11644 (N_11644,N_8904,N_9957);
and U11645 (N_11645,N_8393,N_7390);
nor U11646 (N_11646,N_8703,N_7792);
and U11647 (N_11647,N_8855,N_5885);
nand U11648 (N_11648,N_8408,N_8419);
nor U11649 (N_11649,N_5931,N_8452);
or U11650 (N_11650,N_9261,N_9179);
and U11651 (N_11651,N_9978,N_5339);
and U11652 (N_11652,N_7413,N_8567);
nand U11653 (N_11653,N_5345,N_9275);
or U11654 (N_11654,N_5128,N_7393);
nand U11655 (N_11655,N_6205,N_8135);
nor U11656 (N_11656,N_6131,N_6257);
nand U11657 (N_11657,N_5864,N_8391);
xnor U11658 (N_11658,N_9102,N_5450);
or U11659 (N_11659,N_6597,N_9428);
or U11660 (N_11660,N_5957,N_6553);
nor U11661 (N_11661,N_6817,N_9860);
or U11662 (N_11662,N_7881,N_5219);
nor U11663 (N_11663,N_9427,N_8834);
and U11664 (N_11664,N_8019,N_6634);
or U11665 (N_11665,N_7649,N_5062);
nand U11666 (N_11666,N_8142,N_7260);
nor U11667 (N_11667,N_7087,N_9643);
or U11668 (N_11668,N_7802,N_5270);
nor U11669 (N_11669,N_7916,N_6497);
nor U11670 (N_11670,N_7230,N_9627);
nand U11671 (N_11671,N_9129,N_7046);
nor U11672 (N_11672,N_7676,N_8030);
or U11673 (N_11673,N_7715,N_5786);
nand U11674 (N_11674,N_7746,N_9505);
nor U11675 (N_11675,N_5179,N_9562);
or U11676 (N_11676,N_5426,N_7607);
and U11677 (N_11677,N_7333,N_9822);
nor U11678 (N_11678,N_8996,N_5640);
nand U11679 (N_11679,N_5474,N_6151);
nand U11680 (N_11680,N_7115,N_6549);
nand U11681 (N_11681,N_9106,N_5006);
nor U11682 (N_11682,N_7380,N_5105);
nand U11683 (N_11683,N_9170,N_5385);
or U11684 (N_11684,N_5502,N_7267);
or U11685 (N_11685,N_6024,N_7142);
nand U11686 (N_11686,N_8267,N_5714);
nand U11687 (N_11687,N_9007,N_9523);
nand U11688 (N_11688,N_7155,N_7096);
or U11689 (N_11689,N_8726,N_6959);
and U11690 (N_11690,N_5921,N_8430);
nand U11691 (N_11691,N_6012,N_6095);
and U11692 (N_11692,N_7482,N_9354);
nor U11693 (N_11693,N_7414,N_8831);
and U11694 (N_11694,N_5554,N_7829);
or U11695 (N_11695,N_8484,N_6448);
or U11696 (N_11696,N_6582,N_9966);
nand U11697 (N_11697,N_7383,N_6860);
nor U11698 (N_11698,N_6725,N_7007);
or U11699 (N_11699,N_7303,N_9359);
nor U11700 (N_11700,N_9703,N_9500);
and U11701 (N_11701,N_5187,N_9203);
nand U11702 (N_11702,N_9563,N_5461);
or U11703 (N_11703,N_6525,N_6744);
and U11704 (N_11704,N_7417,N_6424);
or U11705 (N_11705,N_7633,N_6489);
and U11706 (N_11706,N_7407,N_6998);
and U11707 (N_11707,N_5319,N_7141);
nand U11708 (N_11708,N_7522,N_7072);
or U11709 (N_11709,N_9936,N_7960);
and U11710 (N_11710,N_9205,N_9092);
nand U11711 (N_11711,N_8768,N_5347);
and U11712 (N_11712,N_7588,N_9050);
nor U11713 (N_11713,N_8466,N_5941);
and U11714 (N_11714,N_6598,N_7926);
xor U11715 (N_11715,N_8274,N_5679);
and U11716 (N_11716,N_9764,N_8127);
nor U11717 (N_11717,N_9600,N_8159);
and U11718 (N_11718,N_7993,N_5376);
and U11719 (N_11719,N_5570,N_8195);
and U11720 (N_11720,N_8607,N_5780);
nor U11721 (N_11721,N_9338,N_8000);
and U11722 (N_11722,N_9572,N_9489);
or U11723 (N_11723,N_8395,N_8540);
nor U11724 (N_11724,N_8504,N_5415);
xnor U11725 (N_11725,N_9476,N_8317);
and U11726 (N_11726,N_9937,N_5891);
or U11727 (N_11727,N_9167,N_7001);
or U11728 (N_11728,N_7342,N_9107);
nand U11729 (N_11729,N_7690,N_7082);
nand U11730 (N_11730,N_7593,N_9242);
or U11731 (N_11731,N_5056,N_8539);
nand U11732 (N_11732,N_6679,N_7504);
xnor U11733 (N_11733,N_7344,N_9986);
and U11734 (N_11734,N_7149,N_5523);
and U11735 (N_11735,N_9023,N_8630);
and U11736 (N_11736,N_7290,N_8054);
nand U11737 (N_11737,N_6055,N_9508);
nor U11738 (N_11738,N_6995,N_9939);
and U11739 (N_11739,N_8257,N_8960);
nor U11740 (N_11740,N_5977,N_8282);
or U11741 (N_11741,N_9954,N_5928);
nand U11742 (N_11742,N_5918,N_5379);
or U11743 (N_11743,N_6565,N_5716);
xnor U11744 (N_11744,N_7595,N_7778);
and U11745 (N_11745,N_7530,N_7670);
and U11746 (N_11746,N_8235,N_8070);
and U11747 (N_11747,N_8468,N_9236);
nor U11748 (N_11748,N_6621,N_8212);
nand U11749 (N_11749,N_9524,N_8786);
or U11750 (N_11750,N_9985,N_7708);
nor U11751 (N_11751,N_5922,N_5149);
and U11752 (N_11752,N_7762,N_8256);
nand U11753 (N_11753,N_6152,N_5499);
nor U11754 (N_11754,N_7885,N_8808);
and U11755 (N_11755,N_7187,N_9462);
nand U11756 (N_11756,N_7441,N_9321);
and U11757 (N_11757,N_8006,N_5201);
or U11758 (N_11758,N_8333,N_5220);
or U11759 (N_11759,N_8545,N_6668);
nand U11760 (N_11760,N_6474,N_6104);
or U11761 (N_11761,N_6876,N_5465);
nor U11762 (N_11762,N_9411,N_8079);
nor U11763 (N_11763,N_6234,N_6437);
nor U11764 (N_11764,N_7449,N_7939);
nor U11765 (N_11765,N_6432,N_7967);
or U11766 (N_11766,N_7143,N_9488);
nand U11767 (N_11767,N_6890,N_9446);
nor U11768 (N_11768,N_7986,N_7662);
and U11769 (N_11769,N_7519,N_5792);
nor U11770 (N_11770,N_6903,N_9448);
and U11771 (N_11771,N_5585,N_5419);
or U11772 (N_11772,N_6924,N_7546);
nor U11773 (N_11773,N_7813,N_8031);
and U11774 (N_11774,N_8681,N_5942);
and U11775 (N_11775,N_7596,N_5298);
or U11776 (N_11776,N_6756,N_5873);
nor U11777 (N_11777,N_9551,N_7658);
nor U11778 (N_11778,N_6862,N_9850);
or U11779 (N_11779,N_5206,N_8376);
nor U11780 (N_11780,N_5381,N_8621);
and U11781 (N_11781,N_7723,N_7654);
or U11782 (N_11782,N_6017,N_5849);
nor U11783 (N_11783,N_5309,N_6351);
or U11784 (N_11784,N_6106,N_7463);
nor U11785 (N_11785,N_9426,N_6738);
nand U11786 (N_11786,N_7151,N_6763);
or U11787 (N_11787,N_7163,N_8917);
or U11788 (N_11788,N_9924,N_5368);
and U11789 (N_11789,N_7950,N_7445);
nand U11790 (N_11790,N_5788,N_6275);
nand U11791 (N_11791,N_9444,N_9163);
nor U11792 (N_11792,N_9663,N_9212);
nand U11793 (N_11793,N_5656,N_7756);
nand U11794 (N_11794,N_9265,N_6486);
and U11795 (N_11795,N_9002,N_5827);
and U11796 (N_11796,N_5898,N_7205);
nand U11797 (N_11797,N_7598,N_5757);
or U11798 (N_11798,N_7324,N_5476);
and U11799 (N_11799,N_6921,N_6072);
and U11800 (N_11800,N_7027,N_7652);
nor U11801 (N_11801,N_8810,N_7505);
nand U11802 (N_11802,N_7502,N_6967);
xnor U11803 (N_11803,N_9164,N_9697);
and U11804 (N_11804,N_7821,N_5157);
nor U11805 (N_11805,N_7173,N_5003);
or U11806 (N_11806,N_8838,N_6805);
or U11807 (N_11807,N_6833,N_9168);
nor U11808 (N_11808,N_8756,N_7224);
or U11809 (N_11809,N_9587,N_9529);
or U11810 (N_11810,N_9577,N_8841);
and U11811 (N_11811,N_5769,N_8582);
and U11812 (N_11812,N_5480,N_8413);
or U11813 (N_11813,N_8386,N_8092);
nand U11814 (N_11814,N_8568,N_7844);
nand U11815 (N_11815,N_6281,N_8916);
or U11816 (N_11816,N_9898,N_5277);
and U11817 (N_11817,N_6030,N_6546);
nor U11818 (N_11818,N_5766,N_9315);
nor U11819 (N_11819,N_9710,N_8959);
nand U11820 (N_11820,N_9546,N_5999);
nor U11821 (N_11821,N_7283,N_6561);
nand U11822 (N_11822,N_8465,N_8312);
nor U11823 (N_11823,N_8723,N_9415);
nor U11824 (N_11824,N_5331,N_7512);
or U11825 (N_11825,N_9204,N_5120);
or U11826 (N_11826,N_8982,N_6664);
and U11827 (N_11827,N_7156,N_8018);
or U11828 (N_11828,N_6606,N_6853);
nor U11829 (N_11829,N_8778,N_9617);
nand U11830 (N_11830,N_7797,N_7293);
nand U11831 (N_11831,N_5564,N_7669);
and U11832 (N_11832,N_9174,N_8853);
nor U11833 (N_11833,N_6846,N_6272);
and U11834 (N_11834,N_9695,N_6440);
nor U11835 (N_11835,N_5357,N_9795);
nor U11836 (N_11836,N_8676,N_6927);
and U11837 (N_11837,N_9517,N_7576);
or U11838 (N_11838,N_8974,N_5899);
nand U11839 (N_11839,N_8128,N_9440);
nor U11840 (N_11840,N_9645,N_8799);
nor U11841 (N_11841,N_8100,N_5802);
nor U11842 (N_11842,N_8520,N_7075);
nor U11843 (N_11843,N_9930,N_6822);
or U11844 (N_11844,N_9817,N_9056);
and U11845 (N_11845,N_7668,N_5051);
and U11846 (N_11846,N_7925,N_7696);
nand U11847 (N_11847,N_8463,N_6587);
nand U11848 (N_11848,N_6800,N_6885);
or U11849 (N_11849,N_6495,N_5355);
nand U11850 (N_11850,N_7964,N_9652);
nand U11851 (N_11851,N_8334,N_8744);
and U11852 (N_11852,N_7250,N_7875);
and U11853 (N_11853,N_5218,N_5965);
nand U11854 (N_11854,N_9046,N_6097);
and U11855 (N_11855,N_8733,N_7103);
or U11856 (N_11856,N_8909,N_9746);
and U11857 (N_11857,N_8247,N_7857);
nor U11858 (N_11858,N_9112,N_6820);
nor U11859 (N_11859,N_9166,N_8651);
or U11860 (N_11860,N_6179,N_5453);
and U11861 (N_11861,N_8354,N_5156);
nor U11862 (N_11862,N_8067,N_8362);
nor U11863 (N_11863,N_6522,N_9048);
or U11864 (N_11864,N_9146,N_6188);
and U11865 (N_11865,N_9227,N_7298);
nor U11866 (N_11866,N_8499,N_6067);
xnor U11867 (N_11867,N_5969,N_6789);
or U11868 (N_11868,N_7277,N_9307);
or U11869 (N_11869,N_5747,N_7772);
or U11870 (N_11870,N_5216,N_9310);
nor U11871 (N_11871,N_7062,N_9294);
nor U11872 (N_11872,N_8800,N_9602);
nand U11873 (N_11873,N_8880,N_9043);
nor U11874 (N_11874,N_6417,N_6770);
nand U11875 (N_11875,N_8472,N_5646);
xnor U11876 (N_11876,N_9389,N_7699);
or U11877 (N_11877,N_6915,N_5067);
nand U11878 (N_11878,N_5601,N_9420);
and U11879 (N_11879,N_7095,N_8455);
nand U11880 (N_11880,N_8308,N_7308);
or U11881 (N_11881,N_9575,N_7727);
nor U11882 (N_11882,N_9175,N_6241);
nor U11883 (N_11883,N_6620,N_8172);
and U11884 (N_11884,N_5238,N_9191);
nor U11885 (N_11885,N_8174,N_5129);
and U11886 (N_11886,N_5778,N_6414);
and U11887 (N_11887,N_9496,N_8156);
nand U11888 (N_11888,N_9072,N_7097);
nor U11889 (N_11889,N_7070,N_5851);
or U11890 (N_11890,N_7663,N_8962);
nand U11891 (N_11891,N_7757,N_9922);
or U11892 (N_11892,N_7313,N_7783);
nand U11893 (N_11893,N_6720,N_5543);
and U11894 (N_11894,N_6976,N_5423);
and U11895 (N_11895,N_7587,N_6026);
and U11896 (N_11896,N_9503,N_5042);
nor U11897 (N_11897,N_9947,N_9074);
and U11898 (N_11898,N_6136,N_7051);
and U11899 (N_11899,N_6857,N_6242);
or U11900 (N_11900,N_6484,N_5856);
and U11901 (N_11901,N_7520,N_9525);
nand U11902 (N_11902,N_9296,N_7214);
and U11903 (N_11903,N_8735,N_9410);
or U11904 (N_11904,N_6058,N_7220);
or U11905 (N_11905,N_8394,N_5854);
nand U11906 (N_11906,N_8202,N_5366);
or U11907 (N_11907,N_5012,N_6791);
nor U11908 (N_11908,N_5925,N_6133);
nand U11909 (N_11909,N_9187,N_8981);
or U11910 (N_11910,N_8830,N_6564);
nand U11911 (N_11911,N_5525,N_5774);
and U11912 (N_11912,N_5103,N_6253);
nand U11913 (N_11913,N_6577,N_8930);
nand U11914 (N_11914,N_6475,N_5235);
or U11915 (N_11915,N_8887,N_7031);
or U11916 (N_11916,N_7501,N_8155);
and U11917 (N_11917,N_8249,N_7045);
nand U11918 (N_11918,N_6881,N_8932);
or U11919 (N_11919,N_5983,N_8488);
nor U11920 (N_11920,N_5700,N_8033);
nor U11921 (N_11921,N_7219,N_8807);
or U11922 (N_11922,N_9933,N_8891);
or U11923 (N_11923,N_6132,N_6336);
nand U11924 (N_11924,N_6629,N_8356);
nor U11925 (N_11925,N_8361,N_6764);
xnor U11926 (N_11926,N_7563,N_9869);
and U11927 (N_11927,N_6006,N_8674);
and U11928 (N_11928,N_9231,N_8292);
or U11929 (N_11929,N_8899,N_8782);
nand U11930 (N_11930,N_9287,N_5232);
or U11931 (N_11931,N_9750,N_8139);
and U11932 (N_11932,N_6875,N_5784);
or U11933 (N_11933,N_6612,N_5630);
and U11934 (N_11934,N_6844,N_5820);
or U11935 (N_11935,N_9226,N_5100);
nand U11936 (N_11936,N_9678,N_9605);
nand U11937 (N_11937,N_8522,N_9831);
and U11938 (N_11938,N_6051,N_9884);
and U11939 (N_11939,N_9309,N_9483);
and U11940 (N_11940,N_7117,N_7189);
nor U11941 (N_11941,N_5558,N_9200);
nand U11942 (N_11942,N_9960,N_9335);
nand U11943 (N_11943,N_9312,N_6510);
nand U11944 (N_11944,N_6420,N_7432);
or U11945 (N_11945,N_5153,N_5086);
nand U11946 (N_11946,N_5793,N_9455);
nor U11947 (N_11947,N_8506,N_9942);
nand U11948 (N_11948,N_5883,N_5733);
and U11949 (N_11949,N_8780,N_8633);
nor U11950 (N_11950,N_7648,N_7464);
nand U11951 (N_11951,N_9948,N_5573);
and U11952 (N_11952,N_8835,N_7089);
xor U11953 (N_11953,N_9116,N_5691);
or U11954 (N_11954,N_9638,N_8605);
nor U11955 (N_11955,N_8350,N_9159);
or U11956 (N_11956,N_8164,N_6443);
nand U11957 (N_11957,N_7421,N_5763);
nor U11958 (N_11958,N_9308,N_9706);
nand U11959 (N_11959,N_9404,N_6385);
nand U11960 (N_11960,N_8873,N_6994);
or U11961 (N_11961,N_7886,N_8897);
and U11962 (N_11962,N_9510,N_7961);
xor U11963 (N_11963,N_8339,N_9991);
and U11964 (N_11964,N_9124,N_5340);
or U11965 (N_11965,N_7998,N_9771);
nand U11966 (N_11966,N_7826,N_8153);
or U11967 (N_11967,N_6169,N_5663);
nand U11968 (N_11968,N_6056,N_6236);
and U11969 (N_11969,N_7058,N_6117);
nor U11970 (N_11970,N_9247,N_8152);
and U11971 (N_11971,N_6449,N_5927);
and U11972 (N_11972,N_5245,N_6196);
nand U11973 (N_11973,N_7437,N_6485);
nand U11974 (N_11974,N_6777,N_8864);
xnor U11975 (N_11975,N_5842,N_6750);
nor U11976 (N_11976,N_6552,N_8579);
and U11977 (N_11977,N_6094,N_7397);
or U11978 (N_11978,N_7470,N_5978);
nor U11979 (N_11979,N_5444,N_8359);
nand U11980 (N_11980,N_9833,N_8217);
nor U11981 (N_11981,N_8443,N_7627);
or U11982 (N_11982,N_8063,N_5998);
or U11983 (N_11983,N_6936,N_7552);
and U11984 (N_11984,N_7594,N_5739);
or U11985 (N_11985,N_8585,N_5230);
or U11986 (N_11986,N_5684,N_5142);
nand U11987 (N_11987,N_9206,N_5297);
or U11988 (N_11988,N_7428,N_5080);
or U11989 (N_11989,N_7211,N_5872);
nand U11990 (N_11990,N_6114,N_5531);
or U11991 (N_11991,N_7770,N_9879);
nand U11992 (N_11992,N_6965,N_6834);
nor U11993 (N_11993,N_6402,N_5017);
nor U11994 (N_11994,N_6346,N_7306);
or U11995 (N_11995,N_7406,N_7204);
and U11996 (N_11996,N_5404,N_9390);
nand U11997 (N_11997,N_6505,N_5841);
and U11998 (N_11998,N_8720,N_7923);
and U11999 (N_11999,N_5330,N_7759);
and U12000 (N_12000,N_7741,N_6396);
and U12001 (N_12001,N_9409,N_6393);
nand U12002 (N_12002,N_7091,N_7824);
nand U12003 (N_12003,N_6377,N_6064);
or U12004 (N_12004,N_9482,N_9078);
nand U12005 (N_12005,N_6334,N_9724);
and U12006 (N_12006,N_8620,N_7466);
nand U12007 (N_12007,N_7279,N_6581);
nand U12008 (N_12008,N_9818,N_5402);
and U12009 (N_12009,N_6949,N_7368);
nand U12010 (N_12010,N_5013,N_6541);
or U12011 (N_12011,N_7302,N_7566);
and U12012 (N_12012,N_6110,N_5831);
and U12013 (N_12013,N_6790,N_6907);
or U12014 (N_12014,N_7341,N_6652);
or U12015 (N_12015,N_5287,N_9707);
nor U12016 (N_12016,N_7742,N_7347);
and U12017 (N_12017,N_7561,N_9120);
nor U12018 (N_12018,N_7346,N_9412);
nor U12019 (N_12019,N_6478,N_5936);
or U12020 (N_12020,N_5877,N_5354);
or U12021 (N_12021,N_7312,N_8199);
nor U12022 (N_12022,N_9357,N_6295);
nand U12023 (N_12023,N_6246,N_7701);
nor U12024 (N_12024,N_5194,N_5618);
nor U12025 (N_12025,N_5133,N_7809);
nor U12026 (N_12026,N_6043,N_8942);
nand U12027 (N_12027,N_5832,N_6984);
nand U12028 (N_12028,N_8912,N_9929);
or U12029 (N_12029,N_9571,N_6124);
or U12030 (N_12030,N_9378,N_7931);
nand U12031 (N_12031,N_6209,N_5233);
and U12032 (N_12032,N_9499,N_8748);
or U12033 (N_12033,N_5282,N_8663);
nand U12034 (N_12034,N_5628,N_6702);
and U12035 (N_12035,N_6851,N_7548);
nor U12036 (N_12036,N_7128,N_5935);
nor U12037 (N_12037,N_6325,N_9844);
or U12038 (N_12038,N_7764,N_6952);
nor U12039 (N_12039,N_7131,N_6555);
and U12040 (N_12040,N_5866,N_6925);
nor U12041 (N_12041,N_6404,N_5643);
nand U12042 (N_12042,N_9088,N_8047);
nor U12043 (N_12043,N_5974,N_9634);
and U12044 (N_12044,N_8881,N_7689);
nor U12045 (N_12045,N_9382,N_7343);
and U12046 (N_12046,N_7879,N_6878);
nor U12047 (N_12047,N_8945,N_7773);
and U12048 (N_12048,N_8022,N_5980);
or U12049 (N_12049,N_8113,N_5198);
or U12050 (N_12050,N_9024,N_6238);
nor U12051 (N_12051,N_7626,N_9381);
nand U12052 (N_12052,N_8832,N_9810);
nor U12053 (N_12053,N_8134,N_5148);
nor U12054 (N_12054,N_6637,N_9067);
nor U12055 (N_12055,N_7243,N_9796);
and U12056 (N_12056,N_7929,N_5092);
or U12057 (N_12057,N_9865,N_6161);
and U12058 (N_12058,N_9319,N_7799);
nand U12059 (N_12059,N_5509,N_6146);
nor U12060 (N_12060,N_5938,N_5870);
nor U12061 (N_12061,N_8562,N_5940);
nor U12062 (N_12062,N_7276,N_8291);
nor U12063 (N_12063,N_8719,N_5440);
nand U12064 (N_12064,N_8593,N_5468);
or U12065 (N_12065,N_5249,N_8116);
or U12066 (N_12066,N_9141,N_8254);
or U12067 (N_12067,N_9320,N_5244);
nor U12068 (N_12068,N_6828,N_8447);
nor U12069 (N_12069,N_6589,N_9864);
or U12070 (N_12070,N_6867,N_9886);
nand U12071 (N_12071,N_9103,N_9797);
and U12072 (N_12072,N_7839,N_7109);
and U12073 (N_12073,N_5328,N_5544);
and U12074 (N_12074,N_6129,N_9858);
nor U12075 (N_12075,N_7750,N_9900);
or U12076 (N_12076,N_5011,N_8342);
and U12077 (N_12077,N_5182,N_5588);
and U12078 (N_12078,N_5592,N_5816);
nand U12079 (N_12079,N_6148,N_8084);
or U12080 (N_12080,N_5353,N_6991);
nor U12081 (N_12081,N_5131,N_9792);
nor U12082 (N_12082,N_6788,N_5401);
or U12083 (N_12083,N_8787,N_9807);
or U12084 (N_12084,N_8434,N_6466);
nand U12085 (N_12085,N_8036,N_6879);
nand U12086 (N_12086,N_6955,N_7610);
nand U12087 (N_12087,N_6292,N_6514);
nor U12088 (N_12088,N_9987,N_9314);
nand U12089 (N_12089,N_6411,N_8646);
nand U12090 (N_12090,N_9744,N_7092);
xor U12091 (N_12091,N_7673,N_5452);
or U12092 (N_12092,N_7009,N_6831);
or U12093 (N_12093,N_6423,N_5284);
nand U12094 (N_12094,N_7039,N_7469);
and U12095 (N_12095,N_6775,N_5438);
nand U12096 (N_12096,N_8187,N_6784);
or U12097 (N_12097,N_7531,N_8263);
nor U12098 (N_12098,N_8849,N_6408);
and U12099 (N_12099,N_9660,N_5821);
and U12100 (N_12100,N_6880,N_5180);
nor U12101 (N_12101,N_5547,N_9935);
or U12102 (N_12102,N_7709,N_5057);
nand U12103 (N_12103,N_6375,N_9806);
or U12104 (N_12104,N_6771,N_8437);
and U12105 (N_12105,N_5035,N_6230);
nor U12106 (N_12106,N_8745,N_6076);
and U12107 (N_12107,N_9558,N_5365);
nor U12108 (N_12108,N_6239,N_7932);
nand U12109 (N_12109,N_8302,N_8635);
nor U12110 (N_12110,N_8057,N_7247);
or U12111 (N_12111,N_8645,N_8792);
nor U12112 (N_12112,N_7815,N_9353);
nor U12113 (N_12113,N_7730,N_6395);
nand U12114 (N_12114,N_8264,N_6909);
and U12115 (N_12115,N_6477,N_8772);
and U12116 (N_12116,N_8571,N_8322);
nor U12117 (N_12117,N_6666,N_9240);
nor U12118 (N_12118,N_6809,N_7719);
nand U12119 (N_12119,N_7460,N_6456);
or U12120 (N_12120,N_5289,N_5126);
and U12121 (N_12121,N_7043,N_8816);
nand U12122 (N_12122,N_9709,N_6941);
xor U12123 (N_12123,N_9657,N_8541);
nand U12124 (N_12124,N_7990,N_5721);
and U12125 (N_12125,N_8903,N_7862);
nand U12126 (N_12126,N_8580,N_6363);
or U12127 (N_12127,N_8076,N_6558);
nor U12128 (N_12128,N_6785,N_5211);
xnor U12129 (N_12129,N_7162,N_5697);
nand U12130 (N_12130,N_5541,N_8231);
and U12131 (N_12131,N_8690,N_6476);
nor U12132 (N_12132,N_7334,N_5829);
nor U12133 (N_12133,N_5843,N_5680);
or U12134 (N_12134,N_8324,N_6964);
nor U12135 (N_12135,N_9946,N_8161);
and U12136 (N_12136,N_7860,N_9210);
or U12137 (N_12137,N_9150,N_8099);
nand U12138 (N_12138,N_8631,N_6308);
and U12139 (N_12139,N_7944,N_6759);
nand U12140 (N_12140,N_8353,N_6953);
nand U12141 (N_12141,N_7694,N_7038);
and U12142 (N_12142,N_9530,N_7865);
nand U12143 (N_12143,N_5191,N_8335);
and U12144 (N_12144,N_5834,N_9285);
nand U12145 (N_12145,N_8238,N_8086);
or U12146 (N_12146,N_5167,N_6717);
nand U12147 (N_12147,N_7336,N_5462);
or U12148 (N_12148,N_8446,N_8351);
or U12149 (N_12149,N_7642,N_6251);
or U12150 (N_12150,N_5280,N_9759);
nor U12151 (N_12151,N_6496,N_9161);
nor U12152 (N_12152,N_5759,N_8389);
nor U12153 (N_12153,N_9388,N_5504);
or U12154 (N_12154,N_6511,N_7882);
nand U12155 (N_12155,N_6900,N_8706);
or U12156 (N_12156,N_7554,N_9245);
nor U12157 (N_12157,N_8012,N_8717);
nor U12158 (N_12158,N_6250,N_9739);
nor U12159 (N_12159,N_5946,N_6041);
and U12160 (N_12160,N_8175,N_5847);
and U12161 (N_12161,N_6302,N_9620);
and U12162 (N_12162,N_8573,N_8014);
nand U12163 (N_12163,N_6435,N_8672);
nor U12164 (N_12164,N_9775,N_5259);
or U12165 (N_12165,N_7571,N_7480);
nor U12166 (N_12166,N_5882,N_9894);
nor U12167 (N_12167,N_5567,N_8276);
nor U12168 (N_12168,N_9836,N_9418);
and U12169 (N_12169,N_5373,N_8505);
or U12170 (N_12170,N_6855,N_9783);
or U12171 (N_12171,N_6550,N_6376);
and U12172 (N_12172,N_8576,N_5221);
and U12173 (N_12173,N_9301,N_9456);
nand U12174 (N_12174,N_5242,N_6993);
nand U12175 (N_12175,N_7525,N_5510);
or U12176 (N_12176,N_9973,N_5441);
nand U12177 (N_12177,N_7946,N_9068);
nand U12178 (N_12178,N_7487,N_7291);
or U12179 (N_12179,N_6416,N_5362);
and U12180 (N_12180,N_8603,N_7232);
nand U12181 (N_12181,N_7573,N_5762);
and U12182 (N_12182,N_6705,N_6045);
nor U12183 (N_12183,N_7245,N_9119);
and U12184 (N_12184,N_9940,N_8296);
nand U12185 (N_12185,N_9926,N_9298);
nand U12186 (N_12186,N_6130,N_6807);
or U12187 (N_12187,N_6681,N_9334);
and U12188 (N_12188,N_9585,N_8305);
and U12189 (N_12189,N_9698,N_7901);
xnor U12190 (N_12190,N_9365,N_5064);
nand U12191 (N_12191,N_9358,N_9176);
or U12192 (N_12192,N_9108,N_6922);
nor U12193 (N_12193,N_9878,N_7574);
or U12194 (N_12194,N_6008,N_5776);
nor U12195 (N_12195,N_9862,N_9040);
nor U12196 (N_12196,N_8552,N_7099);
or U12197 (N_12197,N_7899,N_5210);
nand U12198 (N_12198,N_8400,N_8936);
xnor U12199 (N_12199,N_7852,N_5830);
xor U12200 (N_12200,N_6981,N_8682);
nor U12201 (N_12201,N_7451,N_5231);
nor U12202 (N_12202,N_8965,N_5795);
and U12203 (N_12203,N_8323,N_7340);
nand U12204 (N_12204,N_9041,N_6665);
nand U12205 (N_12205,N_8673,N_6211);
nand U12206 (N_12206,N_7934,N_5279);
nor U12207 (N_12207,N_7819,N_8363);
and U12208 (N_12208,N_9970,N_8951);
or U12209 (N_12209,N_7834,N_7895);
or U12210 (N_12210,N_9387,N_5265);
and U12211 (N_12211,N_5993,N_8454);
and U12212 (N_12212,N_9447,N_9568);
and U12213 (N_12213,N_6490,N_7957);
or U12214 (N_12214,N_8924,N_6741);
and U12215 (N_12215,N_8762,N_7251);
nand U12216 (N_12216,N_5514,N_9140);
nor U12217 (N_12217,N_5702,N_9837);
or U12218 (N_12218,N_8843,N_5378);
xnor U12219 (N_12219,N_7446,N_5748);
nand U12220 (N_12220,N_9036,N_8039);
or U12221 (N_12221,N_5399,N_6228);
and U12222 (N_12222,N_6358,N_5384);
nand U12223 (N_12223,N_6084,N_5097);
nand U12224 (N_12224,N_7444,N_9816);
nor U12225 (N_12225,N_7492,N_5989);
nor U12226 (N_12226,N_6461,N_8894);
and U12227 (N_12227,N_6544,N_5952);
or U12228 (N_12228,N_9266,N_7348);
nand U12229 (N_12229,N_5529,N_9823);
nor U12230 (N_12230,N_6779,N_5609);
or U12231 (N_12231,N_8131,N_6539);
nand U12232 (N_12232,N_8355,N_6299);
or U12233 (N_12233,N_6460,N_9188);
nand U12234 (N_12234,N_5045,N_5814);
nor U12235 (N_12235,N_6271,N_5213);
or U12236 (N_12236,N_5836,N_8643);
nor U12237 (N_12237,N_9971,N_8721);
nor U12238 (N_12238,N_6382,N_7947);
and U12239 (N_12239,N_6137,N_6077);
and U12240 (N_12240,N_8379,N_9555);
or U12241 (N_12241,N_5169,N_8295);
nand U12242 (N_12242,N_9172,N_8387);
nand U12243 (N_12243,N_7474,N_5708);
nand U12244 (N_12244,N_9599,N_8915);
and U12245 (N_12245,N_9230,N_5084);
or U12246 (N_12246,N_6248,N_6223);
nor U12247 (N_12247,N_8045,N_7498);
or U12248 (N_12248,N_9032,N_8632);
or U12249 (N_12249,N_9063,N_8038);
nand U12250 (N_12250,N_7107,N_9182);
or U12251 (N_12251,N_5751,N_6515);
nor U12252 (N_12252,N_7518,N_6410);
nor U12253 (N_12253,N_7169,N_5283);
nand U12254 (N_12254,N_5391,N_5407);
nand U12255 (N_12255,N_9846,N_6203);
nand U12256 (N_12256,N_8473,N_5411);
or U12257 (N_12257,N_8260,N_5026);
nand U12258 (N_12258,N_7425,N_8598);
nand U12259 (N_12259,N_7253,N_8062);
and U12260 (N_12260,N_9075,N_8958);
and U12261 (N_12261,N_5964,N_6139);
nor U12262 (N_12262,N_7717,N_8698);
nor U12263 (N_12263,N_9871,N_8154);
and U12264 (N_12264,N_9283,N_8869);
nor U12265 (N_12265,N_7168,N_9610);
and U12266 (N_12266,N_7387,N_7472);
nand U12267 (N_12267,N_9246,N_8775);
nand U12268 (N_12268,N_8196,N_8847);
and U12269 (N_12269,N_7704,N_9981);
or U12270 (N_12270,N_6708,N_6990);
nand U12271 (N_12271,N_9917,N_9873);
nand U12272 (N_12272,N_7233,N_9583);
and U12273 (N_12273,N_6985,N_5645);
or U12274 (N_12274,N_5850,N_9281);
nand U12275 (N_12275,N_7040,N_9988);
or U12276 (N_12276,N_5736,N_6359);
xnor U12277 (N_12277,N_9339,N_9279);
xnor U12278 (N_12278,N_5734,N_8177);
nor U12279 (N_12279,N_5052,N_9380);
nor U12280 (N_12280,N_8192,N_9019);
nand U12281 (N_12281,N_7137,N_8285);
and U12282 (N_12282,N_5437,N_7618);
and U12283 (N_12283,N_5294,N_7106);
and U12284 (N_12284,N_8009,N_5031);
nand U12285 (N_12285,N_5565,N_9574);
or U12286 (N_12286,N_9812,N_5151);
nor U12287 (N_12287,N_8314,N_5482);
and U12288 (N_12288,N_8416,N_5662);
nor U12289 (N_12289,N_8628,N_6365);
or U12290 (N_12290,N_6011,N_7614);
xor U12291 (N_12291,N_6194,N_6714);
nor U12292 (N_12292,N_6698,N_5627);
nor U12293 (N_12293,N_8795,N_7838);
nand U12294 (N_12294,N_9712,N_6278);
nand U12295 (N_12295,N_8686,N_6081);
and U12296 (N_12296,N_6436,N_7956);
nand U12297 (N_12297,N_6512,N_6729);
and U12298 (N_12298,N_7060,N_8854);
and U12299 (N_12299,N_5846,N_9374);
and U12300 (N_12300,N_6745,N_6368);
and U12301 (N_12301,N_6207,N_6075);
and U12302 (N_12302,N_5619,N_9352);
or U12303 (N_12303,N_5987,N_7410);
and U12304 (N_12304,N_5746,N_8509);
and U12305 (N_12305,N_5676,N_7493);
nand U12306 (N_12306,N_5058,N_5723);
nand U12307 (N_12307,N_5479,N_5094);
and U12308 (N_12308,N_7859,N_9209);
nor U12309 (N_12309,N_6676,N_9606);
nor U12310 (N_12310,N_6303,N_7575);
nand U12311 (N_12311,N_9368,N_9719);
and U12312 (N_12312,N_6493,N_9623);
and U12313 (N_12313,N_5698,N_6699);
nand U12314 (N_12314,N_5257,N_6150);
or U12315 (N_12315,N_7705,N_5920);
nand U12316 (N_12316,N_8696,N_9181);
and U12317 (N_12317,N_8722,N_5995);
xor U12318 (N_12318,N_7203,N_6852);
nand U12319 (N_12319,N_8326,N_9361);
nand U12320 (N_12320,N_8883,N_7132);
nand U12321 (N_12321,N_6082,N_6926);
or U12322 (N_12322,N_7067,N_8890);
or U12323 (N_12323,N_8550,N_5147);
and U12324 (N_12324,N_8757,N_9805);
xor U12325 (N_12325,N_9062,N_7266);
nand U12326 (N_12326,N_9243,N_7515);
and U12327 (N_12327,N_9509,N_6901);
nand U12328 (N_12328,N_9147,N_9087);
nand U12329 (N_12329,N_8043,N_7744);
nand U12330 (N_12330,N_6467,N_8840);
nand U12331 (N_12331,N_7035,N_9791);
nor U12332 (N_12332,N_6201,N_5071);
and U12333 (N_12333,N_9069,N_7624);
nor U12334 (N_12334,N_9221,N_7619);
and U12335 (N_12335,N_6509,N_5744);
nand U12336 (N_12336,N_6978,N_9360);
nor U12337 (N_12337,N_7175,N_5771);
and U12338 (N_12338,N_9895,N_8502);
and U12339 (N_12339,N_9961,N_9540);
nor U12340 (N_12340,N_8272,N_9276);
nor U12341 (N_12341,N_5237,N_7843);
or U12342 (N_12342,N_6312,N_7606);
nor U12343 (N_12343,N_7252,N_7779);
and U12344 (N_12344,N_9017,N_6032);
or U12345 (N_12345,N_5124,N_6039);
or U12346 (N_12346,N_5805,N_5143);
nand U12347 (N_12347,N_7814,N_9609);
nor U12348 (N_12348,N_7514,N_6682);
nor U12349 (N_12349,N_7917,N_9449);
nor U12350 (N_12350,N_5960,N_6983);
and U12351 (N_12351,N_8162,N_6036);
or U12352 (N_12352,N_8233,N_7101);
and U12353 (N_12353,N_8985,N_8320);
nand U12354 (N_12354,N_7127,N_5561);
and U12355 (N_12355,N_5135,N_9854);
or U12356 (N_12356,N_8332,N_9233);
nor U12357 (N_12357,N_5709,N_6434);
nand U12358 (N_12358,N_5329,N_7317);
nor U12359 (N_12359,N_7420,N_7071);
and U12360 (N_12360,N_5810,N_6904);
nand U12361 (N_12361,N_5672,N_5903);
and U12362 (N_12362,N_8132,N_9881);
nor U12363 (N_12363,N_7949,N_9377);
nor U12364 (N_12364,N_5255,N_9557);
nand U12365 (N_12365,N_5629,N_5115);
and U12366 (N_12366,N_9416,N_7236);
or U12367 (N_12367,N_7135,N_8839);
and U12368 (N_12368,N_8908,N_9673);
nand U12369 (N_12369,N_9105,N_6164);
nor U12370 (N_12370,N_6866,N_5542);
or U12371 (N_12371,N_5420,N_5417);
and U12372 (N_12372,N_6162,N_9951);
nor U12373 (N_12373,N_8458,N_7795);
and U12374 (N_12374,N_7914,N_6757);
nor U12375 (N_12375,N_5848,N_8144);
or U12376 (N_12376,N_6596,N_9909);
nand U12377 (N_12377,N_5229,N_6399);
or U12378 (N_12378,N_7585,N_9356);
xor U12379 (N_12379,N_5291,N_5812);
nor U12380 (N_12380,N_9010,N_5108);
nor U12381 (N_12381,N_8844,N_9405);
and U12382 (N_12382,N_9519,N_8814);
nand U12383 (N_12383,N_5305,N_7227);
and U12384 (N_12384,N_9029,N_9762);
nor U12385 (N_12385,N_6202,N_7794);
or U12386 (N_12386,N_9803,N_7005);
or U12387 (N_12387,N_7032,N_8097);
nor U12388 (N_12388,N_5308,N_6902);
nor U12389 (N_12389,N_5081,N_9089);
or U12390 (N_12390,N_6602,N_6138);
and U12391 (N_12391,N_8811,N_8949);
and U12392 (N_12392,N_6636,N_5552);
and U12393 (N_12393,N_7144,N_7047);
nor U12394 (N_12394,N_5701,N_7453);
and U12395 (N_12395,N_8680,N_5689);
and U12396 (N_12396,N_9914,N_8730);
or U12397 (N_12397,N_9923,N_9268);
and U12398 (N_12398,N_5738,N_6115);
nor U12399 (N_12399,N_7085,N_6170);
nor U12400 (N_12400,N_5537,N_9647);
xor U12401 (N_12401,N_9526,N_5515);
and U12402 (N_12402,N_6421,N_8842);
and U12403 (N_12403,N_8093,N_6631);
xor U12404 (N_12404,N_6407,N_5967);
and U12405 (N_12405,N_9781,N_8273);
nor U12406 (N_12406,N_9076,N_6492);
and U12407 (N_12407,N_6832,N_8999);
or U12408 (N_12408,N_9802,N_5853);
and U12409 (N_12409,N_8331,N_8299);
nand U12410 (N_12410,N_6956,N_5611);
nor U12411 (N_12411,N_9888,N_7010);
and U12412 (N_12412,N_7706,N_8491);
nand U12413 (N_12413,N_7305,N_9876);
nor U12414 (N_12414,N_6232,N_8616);
nand U12415 (N_12415,N_6560,N_5985);
nand U12416 (N_12416,N_9399,N_9892);
nand U12417 (N_12417,N_7036,N_5522);
nand U12418 (N_12418,N_8742,N_5049);
nand U12419 (N_12419,N_6330,N_6605);
nor U12420 (N_12420,N_9651,N_9215);
and U12421 (N_12421,N_8641,N_9122);
nor U12422 (N_12422,N_8905,N_8215);
nor U12423 (N_12423,N_7000,N_9972);
nor U12424 (N_12424,N_5322,N_6814);
nor U12425 (N_12425,N_9132,N_8240);
or U12426 (N_12426,N_8115,N_8157);
nand U12427 (N_12427,N_9027,N_8503);
and U12428 (N_12428,N_5138,N_6107);
or U12429 (N_12429,N_8862,N_9851);
nor U12430 (N_12430,N_8343,N_8130);
nand U12431 (N_12431,N_8103,N_8436);
nor U12432 (N_12432,N_9155,N_9511);
or U12433 (N_12433,N_7269,N_9576);
nor U12434 (N_12434,N_6187,N_8980);
nand U12435 (N_12435,N_8697,N_6562);
and U12436 (N_12436,N_8826,N_6973);
or U12437 (N_12437,N_5868,N_5053);
or U12438 (N_12438,N_5350,N_6762);
nor U12439 (N_12439,N_8740,N_7362);
or U12440 (N_12440,N_7367,N_8422);
nand U12441 (N_12441,N_5015,N_7710);
nand U12442 (N_12442,N_5997,N_6293);
or U12443 (N_12443,N_8160,N_8927);
or U12444 (N_12444,N_9780,N_5176);
nand U12445 (N_12445,N_6394,N_7870);
nor U12446 (N_12446,N_6331,N_5497);
and U12447 (N_12447,N_8955,N_8377);
nand U12448 (N_12448,N_9375,N_5192);
nand U12449 (N_12449,N_5247,N_6733);
nor U12450 (N_12450,N_9941,N_7720);
and U12451 (N_12451,N_5488,N_8535);
and U12452 (N_12452,N_6937,N_8401);
nor U12453 (N_12453,N_8027,N_7375);
and U12454 (N_12454,N_5855,N_7322);
and U12455 (N_12455,N_5160,N_7922);
or U12456 (N_12456,N_5720,N_5667);
nand U12457 (N_12457,N_6753,N_7970);
and U12458 (N_12458,N_9001,N_5926);
nand U12459 (N_12459,N_9229,N_6313);
nor U12460 (N_12460,N_8424,N_9371);
nand U12461 (N_12461,N_6465,N_7215);
or U12462 (N_12462,N_8511,N_8856);
nand U12463 (N_12463,N_6383,N_5171);
nand U12464 (N_12464,N_7851,N_7257);
and U12465 (N_12465,N_7076,N_6929);
or U12466 (N_12466,N_8010,N_5598);
or U12467 (N_12467,N_6684,N_6333);
nor U12468 (N_12468,N_9255,N_5910);
nor U12469 (N_12469,N_5395,N_9699);
or U12470 (N_12470,N_5348,N_7150);
and U12471 (N_12471,N_5141,N_6737);
and U12472 (N_12472,N_7532,N_9867);
or U12473 (N_12473,N_7976,N_9322);
and U12474 (N_12474,N_9543,N_8642);
or U12475 (N_12475,N_8794,N_6615);
or U12476 (N_12476,N_5695,N_9100);
nor U12477 (N_12477,N_9336,N_7262);
and U12478 (N_12478,N_5089,N_5791);
or U12479 (N_12479,N_6001,N_9113);
and U12480 (N_12480,N_8746,N_8119);
xor U12481 (N_12481,N_8124,N_8929);
nor U12482 (N_12482,N_8888,N_9829);
nor U12483 (N_12483,N_9522,N_7332);
nand U12484 (N_12484,N_8044,N_6182);
and U12485 (N_12485,N_9949,N_9039);
or U12486 (N_12486,N_5152,N_9852);
or U12487 (N_12487,N_8427,N_8524);
nor U12488 (N_12488,N_8997,N_6884);
or U12489 (N_12489,N_6559,N_6074);
nand U12490 (N_12490,N_9977,N_7800);
and U12491 (N_12491,N_8064,N_5431);
and U12492 (N_12492,N_7529,N_6783);
or U12493 (N_12493,N_8991,N_6050);
nor U12494 (N_12494,N_5427,N_6390);
nor U12495 (N_12495,N_9284,N_9566);
nor U12496 (N_12496,N_5336,N_7912);
nor U12497 (N_12497,N_6988,N_6883);
nand U12498 (N_12498,N_7461,N_6163);
nor U12499 (N_12499,N_5673,N_9451);
nor U12500 (N_12500,N_5418,N_8502);
and U12501 (N_12501,N_6341,N_8328);
and U12502 (N_12502,N_5814,N_9082);
nor U12503 (N_12503,N_7832,N_8525);
nand U12504 (N_12504,N_7340,N_7084);
or U12505 (N_12505,N_9273,N_9562);
or U12506 (N_12506,N_8820,N_9015);
nand U12507 (N_12507,N_9964,N_9757);
or U12508 (N_12508,N_5245,N_9552);
nand U12509 (N_12509,N_5987,N_6604);
nor U12510 (N_12510,N_8128,N_6829);
or U12511 (N_12511,N_8357,N_8572);
and U12512 (N_12512,N_9481,N_5173);
and U12513 (N_12513,N_7185,N_9629);
xor U12514 (N_12514,N_6072,N_9003);
nor U12515 (N_12515,N_7102,N_7559);
or U12516 (N_12516,N_5996,N_9837);
and U12517 (N_12517,N_8653,N_7775);
nand U12518 (N_12518,N_6596,N_5108);
nor U12519 (N_12519,N_7775,N_8643);
nand U12520 (N_12520,N_5865,N_7867);
nor U12521 (N_12521,N_6661,N_8822);
or U12522 (N_12522,N_8388,N_5984);
nand U12523 (N_12523,N_9484,N_5389);
nand U12524 (N_12524,N_8486,N_5367);
or U12525 (N_12525,N_9870,N_8287);
nor U12526 (N_12526,N_7820,N_9412);
or U12527 (N_12527,N_7248,N_7483);
nor U12528 (N_12528,N_9160,N_9543);
and U12529 (N_12529,N_8376,N_5455);
or U12530 (N_12530,N_5517,N_7294);
or U12531 (N_12531,N_8522,N_9263);
nor U12532 (N_12532,N_8117,N_6838);
and U12533 (N_12533,N_5502,N_9507);
nand U12534 (N_12534,N_6682,N_5009);
nand U12535 (N_12535,N_5909,N_6761);
and U12536 (N_12536,N_7952,N_5743);
nor U12537 (N_12537,N_8489,N_8949);
or U12538 (N_12538,N_5548,N_6607);
nor U12539 (N_12539,N_7584,N_9207);
nand U12540 (N_12540,N_6935,N_6972);
and U12541 (N_12541,N_8161,N_6388);
xor U12542 (N_12542,N_6663,N_6928);
or U12543 (N_12543,N_8715,N_7351);
and U12544 (N_12544,N_5463,N_8049);
or U12545 (N_12545,N_9417,N_6654);
nand U12546 (N_12546,N_9284,N_6523);
nand U12547 (N_12547,N_5533,N_8717);
or U12548 (N_12548,N_9915,N_8743);
nand U12549 (N_12549,N_6930,N_7453);
nand U12550 (N_12550,N_8073,N_7212);
or U12551 (N_12551,N_9480,N_5880);
nor U12552 (N_12552,N_7460,N_8778);
or U12553 (N_12553,N_7326,N_8782);
nand U12554 (N_12554,N_9255,N_9294);
nand U12555 (N_12555,N_8753,N_5167);
or U12556 (N_12556,N_6382,N_9077);
nand U12557 (N_12557,N_5505,N_9751);
and U12558 (N_12558,N_6304,N_8989);
nor U12559 (N_12559,N_9900,N_8832);
and U12560 (N_12560,N_7011,N_7916);
and U12561 (N_12561,N_6255,N_5319);
or U12562 (N_12562,N_5711,N_6798);
or U12563 (N_12563,N_8058,N_5260);
or U12564 (N_12564,N_9331,N_6979);
nor U12565 (N_12565,N_6472,N_9657);
or U12566 (N_12566,N_8973,N_5955);
nand U12567 (N_12567,N_7255,N_8277);
and U12568 (N_12568,N_5467,N_6353);
nor U12569 (N_12569,N_8169,N_8723);
or U12570 (N_12570,N_5196,N_8970);
nand U12571 (N_12571,N_7171,N_5821);
and U12572 (N_12572,N_6615,N_9126);
and U12573 (N_12573,N_5625,N_8224);
nand U12574 (N_12574,N_5818,N_8215);
nor U12575 (N_12575,N_6715,N_7423);
nor U12576 (N_12576,N_6908,N_8547);
nor U12577 (N_12577,N_5955,N_7035);
nand U12578 (N_12578,N_6267,N_8631);
or U12579 (N_12579,N_8999,N_6920);
nor U12580 (N_12580,N_7796,N_6685);
nor U12581 (N_12581,N_6058,N_9928);
nand U12582 (N_12582,N_7606,N_6422);
nor U12583 (N_12583,N_5673,N_5389);
nand U12584 (N_12584,N_7142,N_6256);
nor U12585 (N_12585,N_8636,N_8653);
nand U12586 (N_12586,N_5756,N_5265);
nand U12587 (N_12587,N_9987,N_6253);
nand U12588 (N_12588,N_5315,N_8371);
and U12589 (N_12589,N_9631,N_8614);
nand U12590 (N_12590,N_9885,N_7481);
and U12591 (N_12591,N_5809,N_7445);
and U12592 (N_12592,N_6966,N_6484);
nor U12593 (N_12593,N_7057,N_7007);
nand U12594 (N_12594,N_5993,N_7345);
nor U12595 (N_12595,N_9247,N_9943);
nor U12596 (N_12596,N_9190,N_7482);
nor U12597 (N_12597,N_8588,N_7847);
or U12598 (N_12598,N_6703,N_9925);
nor U12599 (N_12599,N_7018,N_6978);
nand U12600 (N_12600,N_9975,N_6099);
or U12601 (N_12601,N_9338,N_8234);
nand U12602 (N_12602,N_8472,N_7843);
or U12603 (N_12603,N_5473,N_6403);
or U12604 (N_12604,N_8267,N_8360);
and U12605 (N_12605,N_7127,N_6775);
or U12606 (N_12606,N_9204,N_5599);
or U12607 (N_12607,N_7123,N_9708);
nand U12608 (N_12608,N_6667,N_8221);
and U12609 (N_12609,N_6756,N_8186);
and U12610 (N_12610,N_9345,N_8678);
and U12611 (N_12611,N_8940,N_5464);
and U12612 (N_12612,N_5433,N_7069);
nand U12613 (N_12613,N_9710,N_5973);
nand U12614 (N_12614,N_6067,N_8809);
or U12615 (N_12615,N_8248,N_7554);
nand U12616 (N_12616,N_7755,N_9897);
and U12617 (N_12617,N_8967,N_5616);
or U12618 (N_12618,N_7444,N_5599);
and U12619 (N_12619,N_9672,N_5761);
nand U12620 (N_12620,N_5712,N_8231);
nor U12621 (N_12621,N_6255,N_9084);
nor U12622 (N_12622,N_5624,N_7597);
and U12623 (N_12623,N_5555,N_5921);
xnor U12624 (N_12624,N_7934,N_7142);
nand U12625 (N_12625,N_8487,N_9324);
nor U12626 (N_12626,N_7349,N_9643);
or U12627 (N_12627,N_5813,N_9192);
or U12628 (N_12628,N_5537,N_6164);
and U12629 (N_12629,N_6457,N_8982);
nor U12630 (N_12630,N_9374,N_5738);
nand U12631 (N_12631,N_8667,N_9921);
nor U12632 (N_12632,N_5571,N_5144);
or U12633 (N_12633,N_5908,N_7570);
or U12634 (N_12634,N_6217,N_8927);
and U12635 (N_12635,N_8595,N_7937);
nand U12636 (N_12636,N_5890,N_7675);
and U12637 (N_12637,N_7115,N_6345);
nor U12638 (N_12638,N_6713,N_6514);
and U12639 (N_12639,N_5438,N_5164);
and U12640 (N_12640,N_7581,N_5035);
nor U12641 (N_12641,N_6782,N_8037);
nor U12642 (N_12642,N_9603,N_5120);
nor U12643 (N_12643,N_5124,N_6828);
nand U12644 (N_12644,N_5326,N_9412);
nand U12645 (N_12645,N_5561,N_8655);
or U12646 (N_12646,N_6881,N_8912);
and U12647 (N_12647,N_8484,N_7307);
and U12648 (N_12648,N_5090,N_9625);
nor U12649 (N_12649,N_9548,N_6706);
nand U12650 (N_12650,N_7813,N_8884);
or U12651 (N_12651,N_5327,N_8288);
nand U12652 (N_12652,N_6459,N_7474);
nor U12653 (N_12653,N_7989,N_5379);
nand U12654 (N_12654,N_9398,N_7279);
nand U12655 (N_12655,N_5208,N_9804);
nor U12656 (N_12656,N_5811,N_5635);
nand U12657 (N_12657,N_8193,N_8864);
nor U12658 (N_12658,N_6448,N_5627);
and U12659 (N_12659,N_8659,N_5637);
nor U12660 (N_12660,N_6865,N_5824);
nand U12661 (N_12661,N_9163,N_5053);
or U12662 (N_12662,N_5747,N_6313);
nor U12663 (N_12663,N_5543,N_5787);
nor U12664 (N_12664,N_5438,N_9811);
nor U12665 (N_12665,N_9720,N_7092);
xnor U12666 (N_12666,N_7794,N_5736);
nand U12667 (N_12667,N_6341,N_7164);
or U12668 (N_12668,N_9943,N_9282);
or U12669 (N_12669,N_6081,N_6143);
or U12670 (N_12670,N_9741,N_7983);
or U12671 (N_12671,N_6708,N_5329);
or U12672 (N_12672,N_6649,N_9417);
and U12673 (N_12673,N_8291,N_8518);
and U12674 (N_12674,N_7874,N_8460);
and U12675 (N_12675,N_6179,N_5649);
nand U12676 (N_12676,N_7010,N_9899);
or U12677 (N_12677,N_9640,N_8577);
nand U12678 (N_12678,N_7131,N_6524);
or U12679 (N_12679,N_7157,N_9081);
or U12680 (N_12680,N_9408,N_8420);
or U12681 (N_12681,N_9535,N_7163);
and U12682 (N_12682,N_6781,N_9124);
nor U12683 (N_12683,N_5825,N_7781);
nand U12684 (N_12684,N_9586,N_5815);
or U12685 (N_12685,N_9372,N_6590);
nand U12686 (N_12686,N_5770,N_9464);
and U12687 (N_12687,N_5135,N_5819);
nor U12688 (N_12688,N_7037,N_7366);
nor U12689 (N_12689,N_9807,N_9814);
nand U12690 (N_12690,N_8912,N_7290);
or U12691 (N_12691,N_9449,N_6573);
nor U12692 (N_12692,N_7118,N_9251);
or U12693 (N_12693,N_5237,N_6390);
nor U12694 (N_12694,N_7591,N_7645);
nor U12695 (N_12695,N_9770,N_6856);
or U12696 (N_12696,N_7468,N_5791);
nand U12697 (N_12697,N_5053,N_8342);
nand U12698 (N_12698,N_8749,N_6502);
nand U12699 (N_12699,N_6248,N_5124);
or U12700 (N_12700,N_5926,N_7079);
nand U12701 (N_12701,N_5322,N_7717);
and U12702 (N_12702,N_8481,N_7005);
and U12703 (N_12703,N_8205,N_8117);
and U12704 (N_12704,N_6752,N_5288);
or U12705 (N_12705,N_8473,N_5263);
and U12706 (N_12706,N_8283,N_7753);
or U12707 (N_12707,N_9885,N_9123);
or U12708 (N_12708,N_5744,N_8893);
nor U12709 (N_12709,N_5802,N_5873);
or U12710 (N_12710,N_9005,N_7989);
and U12711 (N_12711,N_5011,N_6823);
or U12712 (N_12712,N_8816,N_6432);
or U12713 (N_12713,N_5692,N_7622);
nor U12714 (N_12714,N_6392,N_7454);
nor U12715 (N_12715,N_6403,N_5320);
and U12716 (N_12716,N_5346,N_7722);
nor U12717 (N_12717,N_9039,N_7604);
and U12718 (N_12718,N_5964,N_8476);
nand U12719 (N_12719,N_6731,N_6836);
nor U12720 (N_12720,N_7332,N_8695);
and U12721 (N_12721,N_8167,N_7577);
or U12722 (N_12722,N_8043,N_6411);
or U12723 (N_12723,N_6255,N_8714);
or U12724 (N_12724,N_7079,N_6564);
and U12725 (N_12725,N_5216,N_7970);
and U12726 (N_12726,N_9441,N_7982);
nor U12727 (N_12727,N_8550,N_6449);
or U12728 (N_12728,N_9259,N_7181);
nand U12729 (N_12729,N_8358,N_7734);
nor U12730 (N_12730,N_9459,N_8492);
nor U12731 (N_12731,N_9250,N_5043);
and U12732 (N_12732,N_8562,N_7934);
nor U12733 (N_12733,N_9600,N_9764);
nor U12734 (N_12734,N_7607,N_8572);
or U12735 (N_12735,N_6083,N_9424);
or U12736 (N_12736,N_7472,N_5909);
and U12737 (N_12737,N_7017,N_6552);
and U12738 (N_12738,N_7634,N_7404);
nand U12739 (N_12739,N_9328,N_6932);
or U12740 (N_12740,N_5874,N_9842);
or U12741 (N_12741,N_9304,N_9610);
nor U12742 (N_12742,N_8151,N_7443);
nor U12743 (N_12743,N_8344,N_8357);
nor U12744 (N_12744,N_5714,N_6789);
nand U12745 (N_12745,N_8068,N_6656);
and U12746 (N_12746,N_8306,N_8097);
nand U12747 (N_12747,N_6425,N_9080);
or U12748 (N_12748,N_5583,N_6522);
nand U12749 (N_12749,N_5332,N_9718);
and U12750 (N_12750,N_8697,N_7171);
nand U12751 (N_12751,N_8281,N_9184);
nand U12752 (N_12752,N_6560,N_8360);
nor U12753 (N_12753,N_8806,N_9562);
or U12754 (N_12754,N_6888,N_7730);
nand U12755 (N_12755,N_9947,N_6951);
nand U12756 (N_12756,N_7932,N_5172);
nor U12757 (N_12757,N_6883,N_5485);
or U12758 (N_12758,N_6003,N_5415);
and U12759 (N_12759,N_6577,N_6037);
or U12760 (N_12760,N_7698,N_7422);
or U12761 (N_12761,N_8322,N_9954);
and U12762 (N_12762,N_6774,N_5157);
nand U12763 (N_12763,N_5319,N_5938);
nand U12764 (N_12764,N_6698,N_9344);
or U12765 (N_12765,N_8257,N_5897);
and U12766 (N_12766,N_5929,N_7716);
nor U12767 (N_12767,N_7695,N_7932);
and U12768 (N_12768,N_8285,N_6563);
or U12769 (N_12769,N_6311,N_5482);
nand U12770 (N_12770,N_7128,N_8332);
or U12771 (N_12771,N_7234,N_7096);
and U12772 (N_12772,N_9325,N_9087);
nor U12773 (N_12773,N_8905,N_9528);
nor U12774 (N_12774,N_5496,N_7191);
or U12775 (N_12775,N_9018,N_7623);
nor U12776 (N_12776,N_9167,N_8739);
nand U12777 (N_12777,N_6465,N_5102);
nor U12778 (N_12778,N_8128,N_8374);
and U12779 (N_12779,N_6015,N_6760);
or U12780 (N_12780,N_6332,N_6429);
nor U12781 (N_12781,N_6175,N_5391);
nand U12782 (N_12782,N_9277,N_6419);
nand U12783 (N_12783,N_8335,N_8866);
nor U12784 (N_12784,N_6943,N_7476);
or U12785 (N_12785,N_9948,N_5895);
or U12786 (N_12786,N_6940,N_9570);
and U12787 (N_12787,N_7850,N_6775);
or U12788 (N_12788,N_8691,N_8450);
xor U12789 (N_12789,N_7782,N_6295);
nor U12790 (N_12790,N_7068,N_5534);
nor U12791 (N_12791,N_5870,N_6327);
nand U12792 (N_12792,N_9989,N_8239);
or U12793 (N_12793,N_7413,N_9273);
and U12794 (N_12794,N_6991,N_5875);
nor U12795 (N_12795,N_5068,N_6786);
nor U12796 (N_12796,N_9366,N_9137);
and U12797 (N_12797,N_6921,N_6757);
and U12798 (N_12798,N_7750,N_8245);
nand U12799 (N_12799,N_7804,N_6497);
nor U12800 (N_12800,N_7315,N_7220);
xnor U12801 (N_12801,N_8807,N_6858);
nand U12802 (N_12802,N_8893,N_5341);
nor U12803 (N_12803,N_6461,N_6661);
and U12804 (N_12804,N_5505,N_9361);
or U12805 (N_12805,N_8858,N_9522);
or U12806 (N_12806,N_6134,N_9435);
nor U12807 (N_12807,N_6080,N_8109);
or U12808 (N_12808,N_7416,N_6620);
nor U12809 (N_12809,N_8254,N_9908);
xnor U12810 (N_12810,N_6229,N_7933);
nor U12811 (N_12811,N_7746,N_8622);
nand U12812 (N_12812,N_9177,N_8500);
and U12813 (N_12813,N_7154,N_9676);
nand U12814 (N_12814,N_6429,N_5281);
nand U12815 (N_12815,N_7306,N_9588);
nor U12816 (N_12816,N_9542,N_5788);
or U12817 (N_12817,N_7351,N_6274);
and U12818 (N_12818,N_9346,N_7385);
and U12819 (N_12819,N_9454,N_8826);
and U12820 (N_12820,N_9634,N_8087);
or U12821 (N_12821,N_6002,N_5601);
and U12822 (N_12822,N_5539,N_6704);
or U12823 (N_12823,N_5198,N_8384);
and U12824 (N_12824,N_6127,N_7668);
or U12825 (N_12825,N_9937,N_5208);
nor U12826 (N_12826,N_7009,N_9524);
nor U12827 (N_12827,N_6243,N_6717);
and U12828 (N_12828,N_6239,N_7636);
nand U12829 (N_12829,N_9485,N_7369);
nand U12830 (N_12830,N_9991,N_7219);
nor U12831 (N_12831,N_6493,N_7266);
or U12832 (N_12832,N_9012,N_6916);
nand U12833 (N_12833,N_8483,N_8078);
and U12834 (N_12834,N_9694,N_8409);
and U12835 (N_12835,N_7210,N_6826);
nand U12836 (N_12836,N_6225,N_8970);
nor U12837 (N_12837,N_8946,N_6793);
or U12838 (N_12838,N_6565,N_6101);
nor U12839 (N_12839,N_7218,N_7197);
nor U12840 (N_12840,N_5295,N_7206);
and U12841 (N_12841,N_5270,N_9763);
nand U12842 (N_12842,N_9281,N_6348);
nand U12843 (N_12843,N_6964,N_8131);
nor U12844 (N_12844,N_9486,N_9517);
nand U12845 (N_12845,N_8041,N_9540);
nor U12846 (N_12846,N_7598,N_9106);
nand U12847 (N_12847,N_7976,N_6791);
or U12848 (N_12848,N_9211,N_5546);
xor U12849 (N_12849,N_8155,N_9015);
nor U12850 (N_12850,N_8731,N_8959);
xnor U12851 (N_12851,N_5973,N_7998);
or U12852 (N_12852,N_6764,N_7308);
nor U12853 (N_12853,N_8242,N_7571);
nand U12854 (N_12854,N_7918,N_6130);
nand U12855 (N_12855,N_6387,N_5899);
or U12856 (N_12856,N_7025,N_6668);
nor U12857 (N_12857,N_6416,N_6862);
and U12858 (N_12858,N_6949,N_5605);
nand U12859 (N_12859,N_7034,N_5087);
nand U12860 (N_12860,N_9927,N_8691);
nand U12861 (N_12861,N_6001,N_8805);
nor U12862 (N_12862,N_5536,N_8218);
nor U12863 (N_12863,N_6719,N_7881);
nand U12864 (N_12864,N_5018,N_5653);
and U12865 (N_12865,N_6975,N_8791);
or U12866 (N_12866,N_7186,N_6687);
or U12867 (N_12867,N_5436,N_8617);
or U12868 (N_12868,N_6273,N_5286);
or U12869 (N_12869,N_5824,N_7616);
nor U12870 (N_12870,N_9028,N_6425);
nor U12871 (N_12871,N_7426,N_8157);
nand U12872 (N_12872,N_8442,N_6198);
nor U12873 (N_12873,N_9681,N_6283);
or U12874 (N_12874,N_7958,N_5250);
nor U12875 (N_12875,N_5698,N_8557);
nor U12876 (N_12876,N_7589,N_5923);
and U12877 (N_12877,N_8151,N_9932);
nand U12878 (N_12878,N_7855,N_9070);
or U12879 (N_12879,N_9037,N_7370);
nor U12880 (N_12880,N_7955,N_5292);
and U12881 (N_12881,N_9824,N_9476);
or U12882 (N_12882,N_5082,N_7492);
and U12883 (N_12883,N_5141,N_8113);
and U12884 (N_12884,N_6276,N_7193);
and U12885 (N_12885,N_8714,N_9381);
nand U12886 (N_12886,N_8751,N_8698);
nand U12887 (N_12887,N_6209,N_7815);
or U12888 (N_12888,N_9340,N_6313);
nand U12889 (N_12889,N_5173,N_6615);
nand U12890 (N_12890,N_7804,N_9315);
and U12891 (N_12891,N_8370,N_9760);
nand U12892 (N_12892,N_9335,N_5717);
xor U12893 (N_12893,N_6279,N_8580);
and U12894 (N_12894,N_7794,N_5213);
nand U12895 (N_12895,N_8101,N_9933);
nand U12896 (N_12896,N_6229,N_8632);
nand U12897 (N_12897,N_7526,N_8415);
and U12898 (N_12898,N_8425,N_6647);
nor U12899 (N_12899,N_7515,N_5826);
nand U12900 (N_12900,N_9545,N_6140);
and U12901 (N_12901,N_8515,N_9422);
and U12902 (N_12902,N_6187,N_5584);
and U12903 (N_12903,N_7635,N_6627);
or U12904 (N_12904,N_7534,N_8980);
and U12905 (N_12905,N_8247,N_9471);
xor U12906 (N_12906,N_7724,N_7790);
and U12907 (N_12907,N_6288,N_7361);
nand U12908 (N_12908,N_7329,N_5506);
or U12909 (N_12909,N_6696,N_6084);
nand U12910 (N_12910,N_9876,N_7810);
nor U12911 (N_12911,N_9634,N_6983);
or U12912 (N_12912,N_9641,N_7106);
nand U12913 (N_12913,N_8689,N_7601);
and U12914 (N_12914,N_7530,N_9827);
and U12915 (N_12915,N_7737,N_7548);
nand U12916 (N_12916,N_8212,N_7915);
or U12917 (N_12917,N_9542,N_7125);
and U12918 (N_12918,N_7051,N_7918);
nor U12919 (N_12919,N_8102,N_8186);
and U12920 (N_12920,N_7402,N_7849);
nor U12921 (N_12921,N_8378,N_9777);
or U12922 (N_12922,N_9742,N_6230);
nor U12923 (N_12923,N_6231,N_8325);
nor U12924 (N_12924,N_5794,N_9003);
nor U12925 (N_12925,N_9641,N_6253);
or U12926 (N_12926,N_5488,N_8039);
nand U12927 (N_12927,N_6655,N_5794);
nor U12928 (N_12928,N_7749,N_7553);
nand U12929 (N_12929,N_6459,N_5659);
or U12930 (N_12930,N_7931,N_6778);
and U12931 (N_12931,N_9024,N_9184);
or U12932 (N_12932,N_5482,N_5180);
or U12933 (N_12933,N_5157,N_8292);
and U12934 (N_12934,N_6392,N_8530);
nor U12935 (N_12935,N_5240,N_9284);
xnor U12936 (N_12936,N_7298,N_8628);
and U12937 (N_12937,N_8251,N_9077);
or U12938 (N_12938,N_7469,N_6687);
nor U12939 (N_12939,N_9167,N_9181);
nand U12940 (N_12940,N_6861,N_9123);
and U12941 (N_12941,N_8014,N_8447);
or U12942 (N_12942,N_6419,N_9516);
nor U12943 (N_12943,N_9863,N_9784);
nor U12944 (N_12944,N_8517,N_9243);
xor U12945 (N_12945,N_6521,N_7888);
or U12946 (N_12946,N_7198,N_9721);
or U12947 (N_12947,N_5340,N_9436);
nand U12948 (N_12948,N_6010,N_5724);
nor U12949 (N_12949,N_7821,N_8582);
and U12950 (N_12950,N_7224,N_8299);
or U12951 (N_12951,N_8295,N_8918);
and U12952 (N_12952,N_7967,N_8970);
and U12953 (N_12953,N_6623,N_8147);
or U12954 (N_12954,N_8589,N_8443);
nor U12955 (N_12955,N_6947,N_9940);
nor U12956 (N_12956,N_8722,N_8857);
nand U12957 (N_12957,N_5955,N_8199);
nand U12958 (N_12958,N_6737,N_8615);
nor U12959 (N_12959,N_7981,N_8376);
and U12960 (N_12960,N_8878,N_5476);
or U12961 (N_12961,N_6535,N_8562);
nand U12962 (N_12962,N_7575,N_6750);
or U12963 (N_12963,N_5572,N_6549);
nand U12964 (N_12964,N_6995,N_6065);
nand U12965 (N_12965,N_7135,N_6274);
nand U12966 (N_12966,N_8206,N_9834);
nand U12967 (N_12967,N_8792,N_6111);
or U12968 (N_12968,N_9566,N_5979);
nand U12969 (N_12969,N_8942,N_5824);
nand U12970 (N_12970,N_6368,N_7444);
nand U12971 (N_12971,N_7475,N_7808);
and U12972 (N_12972,N_8217,N_6144);
or U12973 (N_12973,N_5634,N_6428);
xor U12974 (N_12974,N_9760,N_8913);
or U12975 (N_12975,N_5565,N_9272);
nand U12976 (N_12976,N_6220,N_6313);
nand U12977 (N_12977,N_9420,N_8217);
xnor U12978 (N_12978,N_9588,N_8473);
or U12979 (N_12979,N_7896,N_6165);
nor U12980 (N_12980,N_7542,N_6749);
nand U12981 (N_12981,N_6671,N_5129);
nor U12982 (N_12982,N_9671,N_8056);
or U12983 (N_12983,N_8332,N_5663);
and U12984 (N_12984,N_5048,N_7993);
nand U12985 (N_12985,N_8446,N_5048);
or U12986 (N_12986,N_7972,N_7052);
or U12987 (N_12987,N_8415,N_9776);
nand U12988 (N_12988,N_6288,N_8327);
or U12989 (N_12989,N_6479,N_7925);
nor U12990 (N_12990,N_9139,N_9880);
nand U12991 (N_12991,N_7905,N_9899);
and U12992 (N_12992,N_7531,N_6761);
nor U12993 (N_12993,N_5626,N_9160);
nor U12994 (N_12994,N_5774,N_7460);
or U12995 (N_12995,N_6285,N_5637);
or U12996 (N_12996,N_7033,N_9857);
and U12997 (N_12997,N_9850,N_9013);
and U12998 (N_12998,N_9468,N_8947);
nand U12999 (N_12999,N_7459,N_5950);
or U13000 (N_13000,N_9440,N_6754);
nor U13001 (N_13001,N_9959,N_8059);
or U13002 (N_13002,N_6277,N_6524);
nor U13003 (N_13003,N_7841,N_8904);
and U13004 (N_13004,N_8479,N_5935);
nand U13005 (N_13005,N_9169,N_6844);
nor U13006 (N_13006,N_6194,N_9897);
and U13007 (N_13007,N_8357,N_6240);
nor U13008 (N_13008,N_8832,N_8210);
or U13009 (N_13009,N_6951,N_7483);
xor U13010 (N_13010,N_9793,N_7305);
nand U13011 (N_13011,N_6134,N_9497);
nor U13012 (N_13012,N_9904,N_6356);
xnor U13013 (N_13013,N_5534,N_9777);
nand U13014 (N_13014,N_9823,N_9003);
or U13015 (N_13015,N_9692,N_5503);
nand U13016 (N_13016,N_6161,N_6246);
and U13017 (N_13017,N_5404,N_5491);
nor U13018 (N_13018,N_5618,N_6891);
or U13019 (N_13019,N_5521,N_5881);
nand U13020 (N_13020,N_6535,N_9907);
and U13021 (N_13021,N_7266,N_9385);
nor U13022 (N_13022,N_7791,N_9588);
and U13023 (N_13023,N_8501,N_8371);
and U13024 (N_13024,N_9803,N_6497);
nor U13025 (N_13025,N_5570,N_5428);
xnor U13026 (N_13026,N_8663,N_5918);
nor U13027 (N_13027,N_7477,N_8455);
xor U13028 (N_13028,N_5640,N_6312);
and U13029 (N_13029,N_7632,N_8057);
nor U13030 (N_13030,N_6657,N_8717);
nand U13031 (N_13031,N_7017,N_9793);
or U13032 (N_13032,N_5250,N_7751);
nor U13033 (N_13033,N_9180,N_6133);
nand U13034 (N_13034,N_5239,N_6218);
or U13035 (N_13035,N_8759,N_7145);
and U13036 (N_13036,N_9531,N_6929);
nor U13037 (N_13037,N_7620,N_8927);
and U13038 (N_13038,N_7981,N_6644);
and U13039 (N_13039,N_8449,N_8693);
xnor U13040 (N_13040,N_7752,N_7422);
nand U13041 (N_13041,N_6933,N_7984);
and U13042 (N_13042,N_8309,N_9236);
and U13043 (N_13043,N_7819,N_6818);
and U13044 (N_13044,N_6361,N_8800);
nand U13045 (N_13045,N_5873,N_9585);
nand U13046 (N_13046,N_8530,N_6767);
or U13047 (N_13047,N_5069,N_7874);
or U13048 (N_13048,N_5784,N_5482);
nor U13049 (N_13049,N_6056,N_9452);
nor U13050 (N_13050,N_9738,N_7542);
and U13051 (N_13051,N_7744,N_5544);
and U13052 (N_13052,N_5414,N_7397);
nor U13053 (N_13053,N_6512,N_7930);
or U13054 (N_13054,N_6527,N_8159);
nand U13055 (N_13055,N_8713,N_8922);
nand U13056 (N_13056,N_9663,N_5464);
and U13057 (N_13057,N_5537,N_8837);
and U13058 (N_13058,N_5380,N_6533);
nor U13059 (N_13059,N_8273,N_7929);
nand U13060 (N_13060,N_6933,N_6861);
or U13061 (N_13061,N_5205,N_7600);
nand U13062 (N_13062,N_9372,N_7225);
or U13063 (N_13063,N_5791,N_5659);
nor U13064 (N_13064,N_7823,N_7334);
nor U13065 (N_13065,N_7302,N_7653);
nor U13066 (N_13066,N_9219,N_9530);
and U13067 (N_13067,N_5017,N_6974);
and U13068 (N_13068,N_8577,N_9930);
or U13069 (N_13069,N_8741,N_7978);
nand U13070 (N_13070,N_9382,N_8841);
nand U13071 (N_13071,N_9860,N_8951);
and U13072 (N_13072,N_9923,N_7216);
nand U13073 (N_13073,N_8974,N_9629);
or U13074 (N_13074,N_8899,N_5927);
nand U13075 (N_13075,N_5172,N_5695);
or U13076 (N_13076,N_8261,N_8714);
and U13077 (N_13077,N_9756,N_6951);
nand U13078 (N_13078,N_8855,N_9691);
or U13079 (N_13079,N_6737,N_9744);
and U13080 (N_13080,N_6217,N_6030);
and U13081 (N_13081,N_9524,N_7019);
or U13082 (N_13082,N_5791,N_9575);
or U13083 (N_13083,N_6573,N_9315);
and U13084 (N_13084,N_7634,N_7841);
nor U13085 (N_13085,N_6931,N_7428);
or U13086 (N_13086,N_6672,N_5971);
nand U13087 (N_13087,N_8951,N_5974);
nand U13088 (N_13088,N_7214,N_8032);
xnor U13089 (N_13089,N_6430,N_7047);
or U13090 (N_13090,N_5298,N_7659);
and U13091 (N_13091,N_7904,N_8304);
or U13092 (N_13092,N_9423,N_8445);
or U13093 (N_13093,N_7231,N_9281);
and U13094 (N_13094,N_5570,N_7538);
and U13095 (N_13095,N_9003,N_5431);
nand U13096 (N_13096,N_6170,N_7988);
and U13097 (N_13097,N_9542,N_7395);
and U13098 (N_13098,N_6107,N_7220);
or U13099 (N_13099,N_8546,N_5644);
nor U13100 (N_13100,N_6749,N_8643);
or U13101 (N_13101,N_8283,N_5767);
and U13102 (N_13102,N_9855,N_7318);
and U13103 (N_13103,N_9571,N_6282);
nor U13104 (N_13104,N_9485,N_6987);
nand U13105 (N_13105,N_7301,N_6184);
nor U13106 (N_13106,N_6253,N_9280);
or U13107 (N_13107,N_8608,N_6366);
nand U13108 (N_13108,N_9648,N_8199);
nand U13109 (N_13109,N_9145,N_7558);
or U13110 (N_13110,N_9857,N_5951);
nand U13111 (N_13111,N_8344,N_6195);
or U13112 (N_13112,N_5573,N_8090);
nor U13113 (N_13113,N_8198,N_7412);
or U13114 (N_13114,N_6425,N_9874);
nand U13115 (N_13115,N_6987,N_6479);
and U13116 (N_13116,N_9379,N_6069);
and U13117 (N_13117,N_6870,N_7420);
nor U13118 (N_13118,N_5741,N_6424);
nand U13119 (N_13119,N_7621,N_6856);
or U13120 (N_13120,N_9504,N_7121);
nor U13121 (N_13121,N_8630,N_5402);
or U13122 (N_13122,N_7383,N_6653);
nand U13123 (N_13123,N_6759,N_8825);
nor U13124 (N_13124,N_9253,N_6118);
or U13125 (N_13125,N_9650,N_6014);
nand U13126 (N_13126,N_9810,N_5882);
nand U13127 (N_13127,N_6951,N_5853);
nand U13128 (N_13128,N_7602,N_8736);
or U13129 (N_13129,N_8765,N_8246);
and U13130 (N_13130,N_5336,N_5124);
nor U13131 (N_13131,N_7663,N_9173);
xnor U13132 (N_13132,N_5278,N_5516);
nor U13133 (N_13133,N_5743,N_6435);
nand U13134 (N_13134,N_5290,N_6513);
and U13135 (N_13135,N_6839,N_6798);
xor U13136 (N_13136,N_8877,N_6296);
nor U13137 (N_13137,N_5763,N_7927);
nand U13138 (N_13138,N_7461,N_7955);
nand U13139 (N_13139,N_8872,N_5513);
nor U13140 (N_13140,N_7595,N_9043);
or U13141 (N_13141,N_8678,N_6821);
nor U13142 (N_13142,N_8761,N_9827);
and U13143 (N_13143,N_5015,N_7834);
nand U13144 (N_13144,N_6727,N_5385);
nand U13145 (N_13145,N_8911,N_5751);
and U13146 (N_13146,N_5769,N_8428);
and U13147 (N_13147,N_8926,N_6405);
nand U13148 (N_13148,N_6437,N_9090);
or U13149 (N_13149,N_8308,N_6303);
and U13150 (N_13150,N_6529,N_9361);
nand U13151 (N_13151,N_5720,N_5533);
and U13152 (N_13152,N_6326,N_6206);
or U13153 (N_13153,N_7665,N_7986);
nor U13154 (N_13154,N_8344,N_7798);
nor U13155 (N_13155,N_5044,N_9678);
nor U13156 (N_13156,N_5174,N_5902);
or U13157 (N_13157,N_8412,N_5632);
nor U13158 (N_13158,N_5426,N_5297);
nand U13159 (N_13159,N_8426,N_5919);
xor U13160 (N_13160,N_8926,N_5699);
or U13161 (N_13161,N_9570,N_7457);
nor U13162 (N_13162,N_8557,N_5497);
nand U13163 (N_13163,N_7265,N_9054);
and U13164 (N_13164,N_8347,N_6447);
nand U13165 (N_13165,N_7761,N_8151);
nor U13166 (N_13166,N_8074,N_5354);
and U13167 (N_13167,N_6412,N_6195);
or U13168 (N_13168,N_5913,N_6883);
and U13169 (N_13169,N_5957,N_6319);
nand U13170 (N_13170,N_5277,N_6486);
or U13171 (N_13171,N_9060,N_8434);
or U13172 (N_13172,N_7734,N_8834);
or U13173 (N_13173,N_8902,N_7953);
xnor U13174 (N_13174,N_8507,N_9457);
nand U13175 (N_13175,N_9291,N_8665);
nor U13176 (N_13176,N_8018,N_9308);
or U13177 (N_13177,N_5103,N_6279);
xor U13178 (N_13178,N_6080,N_6131);
nand U13179 (N_13179,N_6599,N_7233);
and U13180 (N_13180,N_9913,N_6971);
and U13181 (N_13181,N_9196,N_9548);
and U13182 (N_13182,N_9369,N_5146);
nand U13183 (N_13183,N_9582,N_6737);
or U13184 (N_13184,N_5470,N_8653);
nor U13185 (N_13185,N_8763,N_9696);
nand U13186 (N_13186,N_8251,N_5518);
or U13187 (N_13187,N_5698,N_8104);
nand U13188 (N_13188,N_5286,N_8793);
and U13189 (N_13189,N_9344,N_6791);
nor U13190 (N_13190,N_7470,N_5108);
nand U13191 (N_13191,N_6275,N_5538);
nand U13192 (N_13192,N_6199,N_9820);
and U13193 (N_13193,N_6470,N_8692);
or U13194 (N_13194,N_7629,N_5965);
nand U13195 (N_13195,N_9727,N_9787);
nor U13196 (N_13196,N_6821,N_5085);
or U13197 (N_13197,N_5864,N_5132);
and U13198 (N_13198,N_8292,N_5022);
and U13199 (N_13199,N_8259,N_8285);
nor U13200 (N_13200,N_8701,N_7401);
nor U13201 (N_13201,N_5558,N_8874);
nand U13202 (N_13202,N_9798,N_5034);
and U13203 (N_13203,N_5424,N_7531);
and U13204 (N_13204,N_6121,N_5338);
or U13205 (N_13205,N_5878,N_5683);
or U13206 (N_13206,N_5831,N_5944);
nand U13207 (N_13207,N_6416,N_7516);
or U13208 (N_13208,N_7523,N_5320);
nor U13209 (N_13209,N_8673,N_5463);
nand U13210 (N_13210,N_9278,N_9190);
or U13211 (N_13211,N_7358,N_5520);
and U13212 (N_13212,N_7046,N_9957);
and U13213 (N_13213,N_9209,N_7504);
or U13214 (N_13214,N_7434,N_5516);
and U13215 (N_13215,N_9977,N_9958);
nand U13216 (N_13216,N_5262,N_6602);
nand U13217 (N_13217,N_7714,N_6156);
nand U13218 (N_13218,N_8992,N_5943);
xnor U13219 (N_13219,N_5838,N_9388);
and U13220 (N_13220,N_5860,N_7940);
nor U13221 (N_13221,N_9295,N_5339);
nand U13222 (N_13222,N_8770,N_7446);
nand U13223 (N_13223,N_6649,N_6155);
nand U13224 (N_13224,N_8875,N_7536);
nand U13225 (N_13225,N_6738,N_5920);
or U13226 (N_13226,N_8433,N_9131);
nor U13227 (N_13227,N_7967,N_6642);
or U13228 (N_13228,N_5548,N_7132);
nand U13229 (N_13229,N_7432,N_9354);
nor U13230 (N_13230,N_8137,N_6824);
or U13231 (N_13231,N_9810,N_6530);
nor U13232 (N_13232,N_9537,N_8373);
nor U13233 (N_13233,N_7403,N_9840);
xor U13234 (N_13234,N_7247,N_8214);
nor U13235 (N_13235,N_7007,N_6574);
or U13236 (N_13236,N_6849,N_8023);
nor U13237 (N_13237,N_9944,N_9231);
xor U13238 (N_13238,N_8780,N_5909);
nor U13239 (N_13239,N_7531,N_5218);
nor U13240 (N_13240,N_8459,N_8072);
nand U13241 (N_13241,N_8911,N_5654);
nor U13242 (N_13242,N_5055,N_7515);
nand U13243 (N_13243,N_5176,N_5210);
nor U13244 (N_13244,N_8521,N_9638);
or U13245 (N_13245,N_5855,N_5717);
and U13246 (N_13246,N_5861,N_6414);
or U13247 (N_13247,N_7399,N_8977);
nand U13248 (N_13248,N_7316,N_7260);
nand U13249 (N_13249,N_8826,N_9372);
or U13250 (N_13250,N_9479,N_8049);
or U13251 (N_13251,N_5134,N_6957);
or U13252 (N_13252,N_9134,N_8762);
nand U13253 (N_13253,N_8741,N_8639);
nand U13254 (N_13254,N_9041,N_9350);
nand U13255 (N_13255,N_8362,N_7564);
nor U13256 (N_13256,N_8373,N_5921);
and U13257 (N_13257,N_5775,N_8586);
nand U13258 (N_13258,N_7327,N_7432);
and U13259 (N_13259,N_8829,N_5685);
and U13260 (N_13260,N_5610,N_5343);
nor U13261 (N_13261,N_7753,N_9497);
or U13262 (N_13262,N_9421,N_8144);
nor U13263 (N_13263,N_5457,N_6749);
nor U13264 (N_13264,N_9021,N_8303);
nand U13265 (N_13265,N_9588,N_7759);
nor U13266 (N_13266,N_8787,N_6623);
nor U13267 (N_13267,N_5356,N_6298);
nor U13268 (N_13268,N_7124,N_8527);
nand U13269 (N_13269,N_7415,N_9863);
and U13270 (N_13270,N_7161,N_9919);
nor U13271 (N_13271,N_7040,N_5770);
nor U13272 (N_13272,N_6253,N_6455);
nand U13273 (N_13273,N_5801,N_7521);
and U13274 (N_13274,N_9440,N_7015);
nor U13275 (N_13275,N_5779,N_8153);
nand U13276 (N_13276,N_8490,N_5672);
nand U13277 (N_13277,N_5853,N_7570);
and U13278 (N_13278,N_7934,N_8482);
nand U13279 (N_13279,N_5197,N_8770);
nor U13280 (N_13280,N_5569,N_6952);
nand U13281 (N_13281,N_5577,N_5168);
or U13282 (N_13282,N_6773,N_6917);
nor U13283 (N_13283,N_6420,N_7681);
and U13284 (N_13284,N_5545,N_6459);
or U13285 (N_13285,N_8287,N_8291);
and U13286 (N_13286,N_9565,N_6027);
and U13287 (N_13287,N_7061,N_6067);
and U13288 (N_13288,N_7671,N_5463);
and U13289 (N_13289,N_6180,N_5844);
nor U13290 (N_13290,N_8105,N_7679);
and U13291 (N_13291,N_8185,N_5942);
nor U13292 (N_13292,N_7077,N_9478);
nand U13293 (N_13293,N_5215,N_9834);
or U13294 (N_13294,N_8748,N_6006);
or U13295 (N_13295,N_6873,N_5023);
nand U13296 (N_13296,N_6614,N_5523);
nor U13297 (N_13297,N_7945,N_5563);
nand U13298 (N_13298,N_7514,N_6906);
and U13299 (N_13299,N_5369,N_7331);
and U13300 (N_13300,N_6080,N_5069);
and U13301 (N_13301,N_5081,N_6807);
or U13302 (N_13302,N_8174,N_6776);
nor U13303 (N_13303,N_5190,N_6035);
nand U13304 (N_13304,N_6643,N_5032);
nand U13305 (N_13305,N_8565,N_7480);
or U13306 (N_13306,N_8887,N_6884);
nand U13307 (N_13307,N_5573,N_7572);
nor U13308 (N_13308,N_6969,N_6894);
nor U13309 (N_13309,N_6917,N_8073);
nand U13310 (N_13310,N_9376,N_5873);
and U13311 (N_13311,N_5242,N_9810);
nand U13312 (N_13312,N_8949,N_5483);
and U13313 (N_13313,N_5870,N_9433);
nand U13314 (N_13314,N_5129,N_6377);
nand U13315 (N_13315,N_8582,N_7421);
or U13316 (N_13316,N_7002,N_8527);
nand U13317 (N_13317,N_9009,N_5232);
nor U13318 (N_13318,N_8739,N_7646);
or U13319 (N_13319,N_6325,N_5329);
or U13320 (N_13320,N_5645,N_6033);
nor U13321 (N_13321,N_5366,N_5734);
and U13322 (N_13322,N_5910,N_6204);
nand U13323 (N_13323,N_8903,N_9117);
nand U13324 (N_13324,N_7402,N_7935);
and U13325 (N_13325,N_9911,N_5459);
nand U13326 (N_13326,N_8997,N_8325);
or U13327 (N_13327,N_7031,N_5352);
nand U13328 (N_13328,N_8074,N_6459);
xnor U13329 (N_13329,N_6392,N_7440);
nand U13330 (N_13330,N_9590,N_8837);
nor U13331 (N_13331,N_9058,N_5085);
or U13332 (N_13332,N_6827,N_5341);
nor U13333 (N_13333,N_6764,N_5910);
nand U13334 (N_13334,N_7056,N_8448);
nand U13335 (N_13335,N_6744,N_5378);
or U13336 (N_13336,N_7740,N_9319);
nor U13337 (N_13337,N_9217,N_5598);
nor U13338 (N_13338,N_5957,N_8845);
or U13339 (N_13339,N_7461,N_9859);
nor U13340 (N_13340,N_5964,N_5658);
nor U13341 (N_13341,N_9088,N_9222);
and U13342 (N_13342,N_5491,N_8233);
or U13343 (N_13343,N_7031,N_5804);
nand U13344 (N_13344,N_6627,N_7580);
and U13345 (N_13345,N_6361,N_9112);
nor U13346 (N_13346,N_7422,N_6479);
and U13347 (N_13347,N_8422,N_9329);
or U13348 (N_13348,N_7434,N_5785);
nor U13349 (N_13349,N_9332,N_7578);
nand U13350 (N_13350,N_6170,N_8685);
nand U13351 (N_13351,N_7735,N_9989);
nand U13352 (N_13352,N_6706,N_5107);
and U13353 (N_13353,N_9909,N_5267);
or U13354 (N_13354,N_5256,N_6920);
nor U13355 (N_13355,N_9465,N_9491);
xnor U13356 (N_13356,N_5190,N_9876);
and U13357 (N_13357,N_5865,N_8415);
nor U13358 (N_13358,N_9599,N_5944);
and U13359 (N_13359,N_8938,N_5590);
and U13360 (N_13360,N_7722,N_8895);
nand U13361 (N_13361,N_8272,N_7147);
and U13362 (N_13362,N_9426,N_8577);
nand U13363 (N_13363,N_8003,N_7900);
or U13364 (N_13364,N_8850,N_5654);
nor U13365 (N_13365,N_8391,N_7012);
nor U13366 (N_13366,N_6576,N_6386);
nor U13367 (N_13367,N_6212,N_8396);
nor U13368 (N_13368,N_6426,N_5290);
nor U13369 (N_13369,N_9979,N_8420);
nand U13370 (N_13370,N_8641,N_7709);
and U13371 (N_13371,N_6298,N_6802);
nand U13372 (N_13372,N_8761,N_6636);
and U13373 (N_13373,N_8315,N_6594);
or U13374 (N_13374,N_5299,N_5776);
nand U13375 (N_13375,N_5811,N_8562);
and U13376 (N_13376,N_8386,N_6637);
or U13377 (N_13377,N_8863,N_9622);
and U13378 (N_13378,N_6457,N_5972);
nand U13379 (N_13379,N_8275,N_7051);
and U13380 (N_13380,N_8101,N_8310);
nor U13381 (N_13381,N_7393,N_9237);
nand U13382 (N_13382,N_7321,N_8861);
or U13383 (N_13383,N_8516,N_9378);
or U13384 (N_13384,N_8037,N_5042);
nor U13385 (N_13385,N_9114,N_8806);
or U13386 (N_13386,N_6632,N_7671);
and U13387 (N_13387,N_6929,N_8489);
or U13388 (N_13388,N_7612,N_8747);
or U13389 (N_13389,N_5376,N_6130);
xor U13390 (N_13390,N_5884,N_8692);
nand U13391 (N_13391,N_6871,N_9170);
or U13392 (N_13392,N_5197,N_5254);
nor U13393 (N_13393,N_6455,N_9342);
and U13394 (N_13394,N_8589,N_8111);
nor U13395 (N_13395,N_6674,N_9158);
or U13396 (N_13396,N_5731,N_9506);
and U13397 (N_13397,N_7783,N_6468);
nor U13398 (N_13398,N_5935,N_6129);
nor U13399 (N_13399,N_8356,N_8361);
nand U13400 (N_13400,N_8973,N_6778);
or U13401 (N_13401,N_8401,N_5780);
nor U13402 (N_13402,N_5063,N_8028);
or U13403 (N_13403,N_7790,N_6338);
and U13404 (N_13404,N_9732,N_8634);
and U13405 (N_13405,N_9074,N_6607);
or U13406 (N_13406,N_5892,N_5648);
or U13407 (N_13407,N_8336,N_5384);
nand U13408 (N_13408,N_8937,N_5993);
or U13409 (N_13409,N_7313,N_6630);
nand U13410 (N_13410,N_8207,N_5697);
nand U13411 (N_13411,N_8670,N_5294);
nor U13412 (N_13412,N_7409,N_9437);
or U13413 (N_13413,N_8848,N_6654);
or U13414 (N_13414,N_8289,N_6838);
or U13415 (N_13415,N_7923,N_5091);
nand U13416 (N_13416,N_7261,N_8309);
xor U13417 (N_13417,N_6855,N_8750);
nand U13418 (N_13418,N_6068,N_8549);
nand U13419 (N_13419,N_5246,N_5660);
nor U13420 (N_13420,N_8935,N_8372);
nor U13421 (N_13421,N_8954,N_9207);
and U13422 (N_13422,N_5196,N_6124);
or U13423 (N_13423,N_7436,N_8475);
and U13424 (N_13424,N_6176,N_9039);
nor U13425 (N_13425,N_9039,N_9936);
or U13426 (N_13426,N_8469,N_8820);
or U13427 (N_13427,N_8030,N_7741);
nor U13428 (N_13428,N_8399,N_8947);
nor U13429 (N_13429,N_7693,N_8662);
nand U13430 (N_13430,N_5333,N_5561);
nor U13431 (N_13431,N_5344,N_8069);
and U13432 (N_13432,N_7297,N_7554);
nor U13433 (N_13433,N_6880,N_6330);
or U13434 (N_13434,N_8026,N_8083);
or U13435 (N_13435,N_6245,N_8568);
and U13436 (N_13436,N_5383,N_5617);
and U13437 (N_13437,N_6600,N_7245);
nor U13438 (N_13438,N_5491,N_8301);
nand U13439 (N_13439,N_8306,N_6327);
and U13440 (N_13440,N_6754,N_9194);
and U13441 (N_13441,N_6051,N_5215);
or U13442 (N_13442,N_7932,N_8487);
and U13443 (N_13443,N_7346,N_6081);
and U13444 (N_13444,N_8742,N_5788);
nor U13445 (N_13445,N_7291,N_7295);
and U13446 (N_13446,N_9167,N_5035);
nand U13447 (N_13447,N_7481,N_9019);
or U13448 (N_13448,N_7956,N_6408);
nor U13449 (N_13449,N_6392,N_8026);
nor U13450 (N_13450,N_9471,N_6947);
xor U13451 (N_13451,N_6008,N_5243);
nor U13452 (N_13452,N_5460,N_6788);
nand U13453 (N_13453,N_6257,N_9399);
or U13454 (N_13454,N_6265,N_7664);
nor U13455 (N_13455,N_5981,N_6187);
nand U13456 (N_13456,N_7701,N_7504);
and U13457 (N_13457,N_7843,N_9438);
or U13458 (N_13458,N_6281,N_9036);
nor U13459 (N_13459,N_6191,N_7887);
and U13460 (N_13460,N_9270,N_5445);
nand U13461 (N_13461,N_7827,N_8781);
or U13462 (N_13462,N_7127,N_9382);
nand U13463 (N_13463,N_8429,N_9366);
nand U13464 (N_13464,N_6354,N_8622);
and U13465 (N_13465,N_5659,N_5137);
and U13466 (N_13466,N_7208,N_6387);
and U13467 (N_13467,N_8569,N_6441);
or U13468 (N_13468,N_9056,N_6371);
or U13469 (N_13469,N_9382,N_7637);
or U13470 (N_13470,N_8053,N_7875);
and U13471 (N_13471,N_9473,N_7318);
and U13472 (N_13472,N_7086,N_6712);
and U13473 (N_13473,N_6904,N_5122);
or U13474 (N_13474,N_5155,N_8870);
nor U13475 (N_13475,N_7293,N_6308);
and U13476 (N_13476,N_7696,N_5637);
nor U13477 (N_13477,N_9999,N_7574);
nand U13478 (N_13478,N_6021,N_9873);
nand U13479 (N_13479,N_9050,N_8757);
nor U13480 (N_13480,N_7955,N_5672);
and U13481 (N_13481,N_8706,N_8043);
nor U13482 (N_13482,N_9711,N_7077);
nor U13483 (N_13483,N_5458,N_9192);
nand U13484 (N_13484,N_8493,N_8229);
xnor U13485 (N_13485,N_8483,N_6643);
xor U13486 (N_13486,N_5977,N_8660);
nor U13487 (N_13487,N_9277,N_5747);
nor U13488 (N_13488,N_9406,N_7667);
nand U13489 (N_13489,N_8686,N_7145);
nand U13490 (N_13490,N_5524,N_8112);
nand U13491 (N_13491,N_8502,N_7693);
nor U13492 (N_13492,N_7442,N_5837);
or U13493 (N_13493,N_5571,N_8613);
nand U13494 (N_13494,N_9006,N_8802);
or U13495 (N_13495,N_6958,N_6790);
nand U13496 (N_13496,N_7695,N_7214);
and U13497 (N_13497,N_6903,N_6038);
xnor U13498 (N_13498,N_7136,N_9678);
or U13499 (N_13499,N_7372,N_5256);
or U13500 (N_13500,N_6275,N_5393);
nor U13501 (N_13501,N_8133,N_5956);
nor U13502 (N_13502,N_7596,N_6105);
nand U13503 (N_13503,N_5293,N_6914);
and U13504 (N_13504,N_5251,N_8953);
nand U13505 (N_13505,N_8591,N_5885);
and U13506 (N_13506,N_8434,N_7276);
and U13507 (N_13507,N_8177,N_7239);
or U13508 (N_13508,N_5254,N_9151);
or U13509 (N_13509,N_9877,N_5216);
and U13510 (N_13510,N_7424,N_6070);
and U13511 (N_13511,N_5456,N_5136);
or U13512 (N_13512,N_8832,N_8314);
and U13513 (N_13513,N_8048,N_9569);
and U13514 (N_13514,N_6480,N_7071);
or U13515 (N_13515,N_7933,N_7510);
nor U13516 (N_13516,N_5342,N_8415);
or U13517 (N_13517,N_7226,N_9204);
xor U13518 (N_13518,N_7784,N_8946);
and U13519 (N_13519,N_5274,N_8875);
nor U13520 (N_13520,N_9804,N_8425);
nor U13521 (N_13521,N_8961,N_8057);
nand U13522 (N_13522,N_9959,N_9065);
nor U13523 (N_13523,N_5319,N_9150);
nand U13524 (N_13524,N_9814,N_7836);
nand U13525 (N_13525,N_7663,N_7041);
nor U13526 (N_13526,N_6290,N_5397);
nor U13527 (N_13527,N_9083,N_6176);
and U13528 (N_13528,N_9811,N_6590);
and U13529 (N_13529,N_6768,N_9773);
and U13530 (N_13530,N_5810,N_8942);
nand U13531 (N_13531,N_8104,N_6337);
nor U13532 (N_13532,N_5318,N_8542);
and U13533 (N_13533,N_6373,N_6121);
xor U13534 (N_13534,N_6857,N_5517);
or U13535 (N_13535,N_6194,N_7413);
and U13536 (N_13536,N_8031,N_6499);
or U13537 (N_13537,N_6452,N_6386);
nor U13538 (N_13538,N_7345,N_8322);
or U13539 (N_13539,N_6921,N_9113);
or U13540 (N_13540,N_5034,N_8424);
xor U13541 (N_13541,N_6564,N_8629);
nand U13542 (N_13542,N_7266,N_9007);
nor U13543 (N_13543,N_8716,N_9173);
nor U13544 (N_13544,N_5507,N_6429);
and U13545 (N_13545,N_6415,N_9280);
and U13546 (N_13546,N_6064,N_7693);
or U13547 (N_13547,N_8033,N_6895);
or U13548 (N_13548,N_8557,N_8016);
nand U13549 (N_13549,N_6969,N_8591);
nor U13550 (N_13550,N_9821,N_9235);
and U13551 (N_13551,N_8331,N_7418);
and U13552 (N_13552,N_9124,N_7555);
nand U13553 (N_13553,N_8555,N_8619);
or U13554 (N_13554,N_6452,N_7685);
xor U13555 (N_13555,N_6137,N_9026);
and U13556 (N_13556,N_5699,N_8548);
nor U13557 (N_13557,N_6813,N_7154);
or U13558 (N_13558,N_6496,N_5282);
nor U13559 (N_13559,N_9848,N_6270);
nand U13560 (N_13560,N_6395,N_9978);
nor U13561 (N_13561,N_7034,N_9122);
nand U13562 (N_13562,N_9216,N_7635);
nor U13563 (N_13563,N_5326,N_8331);
nand U13564 (N_13564,N_6760,N_5090);
and U13565 (N_13565,N_6428,N_5775);
xnor U13566 (N_13566,N_8271,N_6923);
or U13567 (N_13567,N_8582,N_7387);
or U13568 (N_13568,N_8974,N_5509);
or U13569 (N_13569,N_8603,N_8593);
nor U13570 (N_13570,N_5074,N_5791);
nor U13571 (N_13571,N_6253,N_9961);
or U13572 (N_13572,N_5247,N_9202);
and U13573 (N_13573,N_9227,N_9684);
or U13574 (N_13574,N_5092,N_8730);
or U13575 (N_13575,N_5357,N_8080);
or U13576 (N_13576,N_8426,N_7258);
nand U13577 (N_13577,N_9388,N_6254);
nor U13578 (N_13578,N_9134,N_6060);
or U13579 (N_13579,N_9623,N_5239);
nor U13580 (N_13580,N_7041,N_9662);
xnor U13581 (N_13581,N_8246,N_8740);
nor U13582 (N_13582,N_9293,N_6705);
nor U13583 (N_13583,N_6082,N_5735);
or U13584 (N_13584,N_8679,N_7449);
nor U13585 (N_13585,N_6140,N_6652);
nor U13586 (N_13586,N_5196,N_5269);
and U13587 (N_13587,N_9868,N_5379);
or U13588 (N_13588,N_6924,N_8020);
nand U13589 (N_13589,N_9002,N_7806);
or U13590 (N_13590,N_9700,N_6428);
or U13591 (N_13591,N_8135,N_7542);
nand U13592 (N_13592,N_7261,N_5254);
nand U13593 (N_13593,N_5459,N_9717);
nand U13594 (N_13594,N_6855,N_6000);
nand U13595 (N_13595,N_8129,N_6541);
nand U13596 (N_13596,N_9864,N_8877);
or U13597 (N_13597,N_8408,N_7176);
and U13598 (N_13598,N_8137,N_7657);
nor U13599 (N_13599,N_7107,N_7788);
nor U13600 (N_13600,N_9236,N_8179);
or U13601 (N_13601,N_7127,N_9721);
or U13602 (N_13602,N_6226,N_8466);
nand U13603 (N_13603,N_8008,N_8456);
nand U13604 (N_13604,N_9608,N_8090);
and U13605 (N_13605,N_7959,N_8542);
nand U13606 (N_13606,N_5045,N_5255);
nor U13607 (N_13607,N_7273,N_6243);
or U13608 (N_13608,N_9162,N_6956);
nor U13609 (N_13609,N_9130,N_5071);
nor U13610 (N_13610,N_8563,N_6359);
or U13611 (N_13611,N_6654,N_5234);
and U13612 (N_13612,N_9801,N_6623);
or U13613 (N_13613,N_9486,N_6289);
nand U13614 (N_13614,N_7944,N_9070);
nand U13615 (N_13615,N_8397,N_6743);
nand U13616 (N_13616,N_9402,N_8453);
or U13617 (N_13617,N_8953,N_8502);
nand U13618 (N_13618,N_9820,N_6988);
and U13619 (N_13619,N_6290,N_9089);
nand U13620 (N_13620,N_7018,N_6016);
and U13621 (N_13621,N_7770,N_7645);
or U13622 (N_13622,N_5028,N_8734);
and U13623 (N_13623,N_7601,N_9103);
or U13624 (N_13624,N_6242,N_9765);
nand U13625 (N_13625,N_5978,N_9292);
or U13626 (N_13626,N_7242,N_6903);
or U13627 (N_13627,N_9258,N_8162);
nand U13628 (N_13628,N_7960,N_8465);
nand U13629 (N_13629,N_6237,N_7905);
and U13630 (N_13630,N_5782,N_8463);
and U13631 (N_13631,N_9366,N_5974);
nor U13632 (N_13632,N_6787,N_5559);
nand U13633 (N_13633,N_6150,N_9538);
or U13634 (N_13634,N_6668,N_7706);
or U13635 (N_13635,N_6976,N_8912);
nand U13636 (N_13636,N_6803,N_5235);
or U13637 (N_13637,N_6430,N_5664);
nand U13638 (N_13638,N_5644,N_5690);
nand U13639 (N_13639,N_5561,N_7840);
and U13640 (N_13640,N_6766,N_7901);
or U13641 (N_13641,N_7474,N_9761);
or U13642 (N_13642,N_8387,N_9345);
or U13643 (N_13643,N_9101,N_5207);
or U13644 (N_13644,N_9439,N_8263);
and U13645 (N_13645,N_6557,N_7980);
and U13646 (N_13646,N_7213,N_8039);
nand U13647 (N_13647,N_6023,N_7214);
or U13648 (N_13648,N_9284,N_8313);
xor U13649 (N_13649,N_7896,N_9294);
or U13650 (N_13650,N_7909,N_5025);
or U13651 (N_13651,N_5090,N_7700);
and U13652 (N_13652,N_6898,N_5534);
nand U13653 (N_13653,N_5325,N_8513);
nand U13654 (N_13654,N_5155,N_8472);
nor U13655 (N_13655,N_6266,N_5688);
and U13656 (N_13656,N_5444,N_8281);
or U13657 (N_13657,N_8760,N_6324);
nand U13658 (N_13658,N_7574,N_9993);
or U13659 (N_13659,N_6424,N_6128);
or U13660 (N_13660,N_8848,N_7631);
nand U13661 (N_13661,N_8535,N_9084);
nor U13662 (N_13662,N_5346,N_5671);
nor U13663 (N_13663,N_5225,N_9302);
or U13664 (N_13664,N_8721,N_8833);
nand U13665 (N_13665,N_5688,N_6185);
nand U13666 (N_13666,N_7409,N_7803);
nor U13667 (N_13667,N_5645,N_8655);
nand U13668 (N_13668,N_5327,N_9480);
nor U13669 (N_13669,N_6939,N_8899);
or U13670 (N_13670,N_9456,N_7647);
nand U13671 (N_13671,N_7268,N_9304);
and U13672 (N_13672,N_7846,N_9207);
or U13673 (N_13673,N_5286,N_9167);
and U13674 (N_13674,N_7407,N_9156);
nand U13675 (N_13675,N_6523,N_5996);
and U13676 (N_13676,N_6545,N_7627);
nor U13677 (N_13677,N_8718,N_5542);
nor U13678 (N_13678,N_8474,N_8605);
and U13679 (N_13679,N_6142,N_5843);
nand U13680 (N_13680,N_6398,N_9551);
nor U13681 (N_13681,N_8582,N_7550);
or U13682 (N_13682,N_5263,N_6178);
nor U13683 (N_13683,N_6836,N_8892);
and U13684 (N_13684,N_5697,N_8819);
and U13685 (N_13685,N_6598,N_9530);
or U13686 (N_13686,N_9856,N_5171);
and U13687 (N_13687,N_6998,N_7589);
nand U13688 (N_13688,N_7792,N_8932);
and U13689 (N_13689,N_5700,N_8817);
nand U13690 (N_13690,N_7679,N_8269);
nand U13691 (N_13691,N_6629,N_7251);
or U13692 (N_13692,N_7744,N_8931);
nand U13693 (N_13693,N_8699,N_7927);
nor U13694 (N_13694,N_9400,N_9354);
or U13695 (N_13695,N_8762,N_6301);
or U13696 (N_13696,N_9311,N_8969);
or U13697 (N_13697,N_6196,N_9379);
nor U13698 (N_13698,N_8144,N_5957);
and U13699 (N_13699,N_9977,N_7858);
nor U13700 (N_13700,N_8907,N_6152);
and U13701 (N_13701,N_9486,N_6145);
nand U13702 (N_13702,N_8264,N_9284);
or U13703 (N_13703,N_5820,N_8120);
nand U13704 (N_13704,N_5400,N_9465);
nor U13705 (N_13705,N_6021,N_8956);
nor U13706 (N_13706,N_9762,N_6515);
and U13707 (N_13707,N_5841,N_9691);
nor U13708 (N_13708,N_7418,N_9088);
or U13709 (N_13709,N_6396,N_5375);
nand U13710 (N_13710,N_8666,N_9517);
or U13711 (N_13711,N_5352,N_9509);
and U13712 (N_13712,N_8956,N_7332);
or U13713 (N_13713,N_8349,N_7296);
nand U13714 (N_13714,N_7811,N_6679);
or U13715 (N_13715,N_7392,N_5069);
and U13716 (N_13716,N_6835,N_8183);
or U13717 (N_13717,N_8928,N_9038);
nor U13718 (N_13718,N_6354,N_8232);
nor U13719 (N_13719,N_6917,N_8168);
or U13720 (N_13720,N_8342,N_9616);
nor U13721 (N_13721,N_8253,N_9748);
nand U13722 (N_13722,N_8442,N_6134);
or U13723 (N_13723,N_8819,N_5730);
nor U13724 (N_13724,N_6554,N_5878);
or U13725 (N_13725,N_7553,N_5807);
nand U13726 (N_13726,N_8150,N_6917);
nand U13727 (N_13727,N_8581,N_5295);
nand U13728 (N_13728,N_8069,N_6946);
nor U13729 (N_13729,N_9096,N_7264);
nand U13730 (N_13730,N_8408,N_6276);
and U13731 (N_13731,N_9250,N_7682);
or U13732 (N_13732,N_9991,N_6301);
xor U13733 (N_13733,N_8738,N_5734);
and U13734 (N_13734,N_5598,N_9060);
and U13735 (N_13735,N_8999,N_8314);
or U13736 (N_13736,N_7653,N_5678);
or U13737 (N_13737,N_6437,N_8908);
nor U13738 (N_13738,N_8413,N_5152);
nor U13739 (N_13739,N_8788,N_5808);
and U13740 (N_13740,N_5086,N_5353);
nor U13741 (N_13741,N_6844,N_8029);
nor U13742 (N_13742,N_9835,N_6326);
nor U13743 (N_13743,N_8180,N_6279);
nand U13744 (N_13744,N_5781,N_5138);
nor U13745 (N_13745,N_5260,N_6558);
and U13746 (N_13746,N_9003,N_8063);
nor U13747 (N_13747,N_9893,N_5320);
nor U13748 (N_13748,N_8889,N_6682);
or U13749 (N_13749,N_8961,N_9400);
nor U13750 (N_13750,N_5373,N_8106);
and U13751 (N_13751,N_7122,N_6995);
nand U13752 (N_13752,N_6189,N_9212);
nor U13753 (N_13753,N_5961,N_5291);
nor U13754 (N_13754,N_8113,N_9578);
and U13755 (N_13755,N_9091,N_5098);
xor U13756 (N_13756,N_7759,N_9219);
nand U13757 (N_13757,N_8942,N_8032);
and U13758 (N_13758,N_5085,N_8618);
nand U13759 (N_13759,N_9017,N_8454);
or U13760 (N_13760,N_7808,N_9658);
and U13761 (N_13761,N_8619,N_9112);
and U13762 (N_13762,N_5619,N_7486);
and U13763 (N_13763,N_5787,N_8994);
and U13764 (N_13764,N_6944,N_7837);
or U13765 (N_13765,N_8267,N_8490);
or U13766 (N_13766,N_7494,N_9083);
nand U13767 (N_13767,N_8081,N_6584);
or U13768 (N_13768,N_5595,N_6223);
and U13769 (N_13769,N_7159,N_6370);
or U13770 (N_13770,N_8876,N_5579);
nor U13771 (N_13771,N_5554,N_7547);
and U13772 (N_13772,N_9599,N_9299);
nand U13773 (N_13773,N_9141,N_6431);
or U13774 (N_13774,N_8584,N_6126);
nand U13775 (N_13775,N_8995,N_5197);
and U13776 (N_13776,N_7088,N_7007);
and U13777 (N_13777,N_6288,N_5523);
nand U13778 (N_13778,N_7037,N_9208);
nor U13779 (N_13779,N_8819,N_9936);
or U13780 (N_13780,N_5021,N_7792);
nand U13781 (N_13781,N_9260,N_7607);
nand U13782 (N_13782,N_8244,N_8596);
and U13783 (N_13783,N_5680,N_8858);
nand U13784 (N_13784,N_9574,N_5872);
nor U13785 (N_13785,N_6394,N_5125);
nor U13786 (N_13786,N_6740,N_6840);
nor U13787 (N_13787,N_8126,N_8850);
nor U13788 (N_13788,N_8799,N_9571);
or U13789 (N_13789,N_6248,N_9092);
nor U13790 (N_13790,N_7301,N_8050);
nand U13791 (N_13791,N_8638,N_8189);
nor U13792 (N_13792,N_7955,N_9113);
nand U13793 (N_13793,N_6331,N_9596);
and U13794 (N_13794,N_6486,N_8004);
or U13795 (N_13795,N_9327,N_6170);
nand U13796 (N_13796,N_8350,N_7399);
nor U13797 (N_13797,N_8213,N_7913);
nor U13798 (N_13798,N_7507,N_5608);
or U13799 (N_13799,N_5730,N_9261);
and U13800 (N_13800,N_9356,N_7310);
nor U13801 (N_13801,N_8267,N_7860);
nor U13802 (N_13802,N_6820,N_9227);
and U13803 (N_13803,N_8714,N_5114);
nand U13804 (N_13804,N_8776,N_5745);
nor U13805 (N_13805,N_5441,N_7493);
or U13806 (N_13806,N_9787,N_9033);
nand U13807 (N_13807,N_8567,N_5280);
or U13808 (N_13808,N_7008,N_7316);
or U13809 (N_13809,N_6524,N_7278);
nand U13810 (N_13810,N_7423,N_8294);
nor U13811 (N_13811,N_8372,N_6766);
or U13812 (N_13812,N_5672,N_5766);
nand U13813 (N_13813,N_6818,N_6017);
or U13814 (N_13814,N_7259,N_9702);
and U13815 (N_13815,N_7501,N_9771);
and U13816 (N_13816,N_7824,N_8785);
nand U13817 (N_13817,N_8207,N_9779);
or U13818 (N_13818,N_7417,N_8832);
and U13819 (N_13819,N_5662,N_7027);
nor U13820 (N_13820,N_5074,N_6099);
nor U13821 (N_13821,N_9345,N_9140);
or U13822 (N_13822,N_6808,N_6138);
and U13823 (N_13823,N_9050,N_6305);
and U13824 (N_13824,N_7124,N_7462);
or U13825 (N_13825,N_6860,N_5810);
and U13826 (N_13826,N_8773,N_9121);
and U13827 (N_13827,N_7185,N_8939);
and U13828 (N_13828,N_5787,N_8532);
or U13829 (N_13829,N_6873,N_5080);
nor U13830 (N_13830,N_6534,N_8038);
or U13831 (N_13831,N_7856,N_6785);
nand U13832 (N_13832,N_8024,N_7014);
or U13833 (N_13833,N_6448,N_8004);
and U13834 (N_13834,N_8761,N_6686);
nor U13835 (N_13835,N_9796,N_9908);
and U13836 (N_13836,N_9717,N_5313);
or U13837 (N_13837,N_8201,N_5972);
and U13838 (N_13838,N_7580,N_8969);
or U13839 (N_13839,N_8449,N_6981);
and U13840 (N_13840,N_5696,N_6629);
or U13841 (N_13841,N_7179,N_6412);
or U13842 (N_13842,N_9382,N_9693);
or U13843 (N_13843,N_8924,N_6618);
or U13844 (N_13844,N_7770,N_8821);
nor U13845 (N_13845,N_6245,N_8904);
and U13846 (N_13846,N_9344,N_5059);
or U13847 (N_13847,N_8555,N_8733);
or U13848 (N_13848,N_6325,N_6807);
and U13849 (N_13849,N_9593,N_7412);
or U13850 (N_13850,N_5010,N_8808);
nand U13851 (N_13851,N_8843,N_8979);
and U13852 (N_13852,N_9300,N_7476);
nor U13853 (N_13853,N_6953,N_9051);
or U13854 (N_13854,N_9301,N_9731);
nand U13855 (N_13855,N_9170,N_5326);
or U13856 (N_13856,N_5742,N_8430);
or U13857 (N_13857,N_6342,N_9267);
nand U13858 (N_13858,N_9019,N_8735);
and U13859 (N_13859,N_7123,N_6418);
nand U13860 (N_13860,N_9901,N_9423);
nor U13861 (N_13861,N_8133,N_8129);
nand U13862 (N_13862,N_6683,N_8331);
nor U13863 (N_13863,N_9639,N_9229);
nand U13864 (N_13864,N_7732,N_9250);
nand U13865 (N_13865,N_6048,N_6676);
or U13866 (N_13866,N_7302,N_7932);
or U13867 (N_13867,N_9076,N_8957);
or U13868 (N_13868,N_7760,N_8583);
nor U13869 (N_13869,N_8891,N_7189);
nor U13870 (N_13870,N_6585,N_5648);
nor U13871 (N_13871,N_7187,N_8311);
nor U13872 (N_13872,N_5149,N_7956);
nand U13873 (N_13873,N_6509,N_5268);
or U13874 (N_13874,N_8831,N_8649);
nand U13875 (N_13875,N_6153,N_8109);
nand U13876 (N_13876,N_5743,N_7010);
and U13877 (N_13877,N_7994,N_7441);
nand U13878 (N_13878,N_7600,N_9418);
nor U13879 (N_13879,N_7789,N_8434);
nor U13880 (N_13880,N_6070,N_9246);
and U13881 (N_13881,N_8385,N_9466);
and U13882 (N_13882,N_6767,N_9004);
nand U13883 (N_13883,N_9418,N_7230);
nand U13884 (N_13884,N_5164,N_6082);
nor U13885 (N_13885,N_8849,N_9071);
nand U13886 (N_13886,N_9355,N_5065);
nor U13887 (N_13887,N_5394,N_9930);
nand U13888 (N_13888,N_6574,N_7852);
nand U13889 (N_13889,N_5646,N_8448);
nand U13890 (N_13890,N_6073,N_9083);
or U13891 (N_13891,N_9072,N_8851);
nor U13892 (N_13892,N_7394,N_6270);
and U13893 (N_13893,N_7658,N_6216);
and U13894 (N_13894,N_6089,N_7120);
or U13895 (N_13895,N_7247,N_6192);
or U13896 (N_13896,N_6058,N_8647);
nor U13897 (N_13897,N_5618,N_9818);
or U13898 (N_13898,N_6910,N_5755);
nor U13899 (N_13899,N_5950,N_7341);
and U13900 (N_13900,N_9510,N_7959);
or U13901 (N_13901,N_8680,N_7299);
or U13902 (N_13902,N_8384,N_8684);
or U13903 (N_13903,N_9951,N_9739);
nor U13904 (N_13904,N_7893,N_5709);
nor U13905 (N_13905,N_9861,N_8771);
and U13906 (N_13906,N_8240,N_7474);
or U13907 (N_13907,N_7690,N_5062);
nand U13908 (N_13908,N_7092,N_8145);
nand U13909 (N_13909,N_7659,N_5339);
and U13910 (N_13910,N_5698,N_6302);
or U13911 (N_13911,N_9817,N_7633);
or U13912 (N_13912,N_6711,N_6451);
nor U13913 (N_13913,N_6378,N_9892);
and U13914 (N_13914,N_7218,N_7506);
nand U13915 (N_13915,N_7846,N_9440);
nor U13916 (N_13916,N_9684,N_6670);
and U13917 (N_13917,N_7453,N_5048);
nor U13918 (N_13918,N_7665,N_7047);
and U13919 (N_13919,N_7345,N_8669);
nand U13920 (N_13920,N_9328,N_6655);
and U13921 (N_13921,N_6054,N_5420);
and U13922 (N_13922,N_9111,N_8376);
nor U13923 (N_13923,N_6068,N_7006);
and U13924 (N_13924,N_5786,N_7253);
and U13925 (N_13925,N_7684,N_7796);
and U13926 (N_13926,N_5731,N_8641);
nor U13927 (N_13927,N_6022,N_8270);
and U13928 (N_13928,N_5844,N_7002);
nor U13929 (N_13929,N_7658,N_9459);
nor U13930 (N_13930,N_7227,N_9363);
or U13931 (N_13931,N_5569,N_5762);
xor U13932 (N_13932,N_6205,N_6214);
nor U13933 (N_13933,N_7979,N_5630);
and U13934 (N_13934,N_8777,N_8350);
or U13935 (N_13935,N_7323,N_8691);
and U13936 (N_13936,N_6102,N_8288);
or U13937 (N_13937,N_7129,N_7822);
and U13938 (N_13938,N_7018,N_9346);
nand U13939 (N_13939,N_7597,N_8542);
nor U13940 (N_13940,N_5663,N_8875);
and U13941 (N_13941,N_5816,N_6608);
or U13942 (N_13942,N_7640,N_9746);
or U13943 (N_13943,N_9277,N_8241);
nand U13944 (N_13944,N_6204,N_5253);
nor U13945 (N_13945,N_7775,N_5398);
nand U13946 (N_13946,N_8049,N_9229);
or U13947 (N_13947,N_8196,N_9612);
nor U13948 (N_13948,N_8512,N_9915);
nor U13949 (N_13949,N_5739,N_6607);
or U13950 (N_13950,N_7373,N_7424);
nand U13951 (N_13951,N_8695,N_8766);
nand U13952 (N_13952,N_5465,N_6459);
and U13953 (N_13953,N_5600,N_8604);
nand U13954 (N_13954,N_5514,N_6127);
nand U13955 (N_13955,N_7447,N_7410);
or U13956 (N_13956,N_7972,N_9414);
or U13957 (N_13957,N_5702,N_8016);
nor U13958 (N_13958,N_8889,N_8826);
nor U13959 (N_13959,N_6118,N_9079);
and U13960 (N_13960,N_6659,N_9505);
and U13961 (N_13961,N_7151,N_8621);
nand U13962 (N_13962,N_5101,N_5740);
nor U13963 (N_13963,N_6738,N_8643);
and U13964 (N_13964,N_6613,N_5728);
nor U13965 (N_13965,N_8564,N_5822);
and U13966 (N_13966,N_8925,N_5357);
or U13967 (N_13967,N_5246,N_7971);
and U13968 (N_13968,N_5219,N_7520);
or U13969 (N_13969,N_8900,N_8964);
or U13970 (N_13970,N_6520,N_9006);
or U13971 (N_13971,N_5387,N_9951);
nor U13972 (N_13972,N_9264,N_8619);
nand U13973 (N_13973,N_5652,N_5313);
or U13974 (N_13974,N_5488,N_7378);
nor U13975 (N_13975,N_8883,N_9651);
and U13976 (N_13976,N_6659,N_8267);
nand U13977 (N_13977,N_9338,N_5981);
and U13978 (N_13978,N_6644,N_6213);
nand U13979 (N_13979,N_9113,N_9955);
xor U13980 (N_13980,N_9383,N_5553);
or U13981 (N_13981,N_8072,N_7134);
or U13982 (N_13982,N_7376,N_7011);
or U13983 (N_13983,N_9918,N_7655);
nand U13984 (N_13984,N_6090,N_6035);
nand U13985 (N_13985,N_9587,N_6673);
or U13986 (N_13986,N_9166,N_7960);
or U13987 (N_13987,N_9577,N_6882);
nand U13988 (N_13988,N_8223,N_5305);
nand U13989 (N_13989,N_6823,N_9525);
and U13990 (N_13990,N_5960,N_5155);
and U13991 (N_13991,N_7933,N_8987);
nand U13992 (N_13992,N_6591,N_8185);
xor U13993 (N_13993,N_5703,N_9130);
nor U13994 (N_13994,N_7597,N_6677);
nor U13995 (N_13995,N_5580,N_7485);
xor U13996 (N_13996,N_7533,N_8704);
nand U13997 (N_13997,N_9529,N_8279);
nor U13998 (N_13998,N_5806,N_8250);
nand U13999 (N_13999,N_6450,N_9588);
xnor U14000 (N_14000,N_7189,N_8325);
or U14001 (N_14001,N_9791,N_8554);
and U14002 (N_14002,N_7740,N_9939);
nand U14003 (N_14003,N_7675,N_8258);
nor U14004 (N_14004,N_9830,N_5932);
and U14005 (N_14005,N_9011,N_8074);
nand U14006 (N_14006,N_6662,N_7051);
nor U14007 (N_14007,N_9346,N_7854);
or U14008 (N_14008,N_6973,N_5192);
nor U14009 (N_14009,N_5180,N_8108);
nor U14010 (N_14010,N_8704,N_6616);
nor U14011 (N_14011,N_9288,N_9675);
nor U14012 (N_14012,N_8843,N_7998);
xor U14013 (N_14013,N_6462,N_9515);
nor U14014 (N_14014,N_5415,N_5305);
or U14015 (N_14015,N_9074,N_7904);
nor U14016 (N_14016,N_7360,N_5765);
and U14017 (N_14017,N_9829,N_6567);
or U14018 (N_14018,N_8298,N_8322);
nand U14019 (N_14019,N_9431,N_5508);
nor U14020 (N_14020,N_6531,N_8109);
nand U14021 (N_14021,N_9848,N_9951);
nand U14022 (N_14022,N_8214,N_7839);
and U14023 (N_14023,N_8900,N_5289);
nand U14024 (N_14024,N_9807,N_5811);
or U14025 (N_14025,N_8252,N_8181);
nand U14026 (N_14026,N_9469,N_6929);
and U14027 (N_14027,N_8353,N_9198);
or U14028 (N_14028,N_7051,N_5465);
nand U14029 (N_14029,N_8143,N_6423);
or U14030 (N_14030,N_9378,N_7555);
or U14031 (N_14031,N_6486,N_5787);
nor U14032 (N_14032,N_6840,N_6414);
and U14033 (N_14033,N_7021,N_6451);
and U14034 (N_14034,N_9321,N_5273);
or U14035 (N_14035,N_9221,N_7138);
and U14036 (N_14036,N_6374,N_5662);
or U14037 (N_14037,N_8572,N_5579);
or U14038 (N_14038,N_9992,N_9042);
nand U14039 (N_14039,N_8736,N_7490);
or U14040 (N_14040,N_5502,N_9107);
nand U14041 (N_14041,N_7721,N_7868);
or U14042 (N_14042,N_7806,N_9533);
and U14043 (N_14043,N_8091,N_9167);
xnor U14044 (N_14044,N_7361,N_6031);
or U14045 (N_14045,N_8054,N_9382);
xnor U14046 (N_14046,N_9909,N_9568);
nor U14047 (N_14047,N_7520,N_9129);
nor U14048 (N_14048,N_7520,N_7991);
nor U14049 (N_14049,N_6320,N_7790);
and U14050 (N_14050,N_7381,N_7690);
and U14051 (N_14051,N_8184,N_8456);
or U14052 (N_14052,N_7683,N_7666);
and U14053 (N_14053,N_6295,N_7450);
nor U14054 (N_14054,N_9328,N_9162);
and U14055 (N_14055,N_6657,N_6372);
and U14056 (N_14056,N_8102,N_7373);
nand U14057 (N_14057,N_5358,N_7107);
nor U14058 (N_14058,N_6639,N_6565);
nor U14059 (N_14059,N_5662,N_6507);
nand U14060 (N_14060,N_7433,N_6705);
nand U14061 (N_14061,N_6849,N_7291);
or U14062 (N_14062,N_5646,N_9965);
nand U14063 (N_14063,N_5364,N_9952);
nor U14064 (N_14064,N_6484,N_8962);
or U14065 (N_14065,N_7103,N_9585);
or U14066 (N_14066,N_6337,N_6415);
or U14067 (N_14067,N_7523,N_7893);
nand U14068 (N_14068,N_9795,N_8707);
nor U14069 (N_14069,N_5838,N_8772);
nand U14070 (N_14070,N_5676,N_8870);
and U14071 (N_14071,N_9756,N_6314);
and U14072 (N_14072,N_6923,N_7372);
or U14073 (N_14073,N_6423,N_8294);
xor U14074 (N_14074,N_8153,N_6624);
xor U14075 (N_14075,N_6479,N_6815);
nand U14076 (N_14076,N_6725,N_9131);
or U14077 (N_14077,N_8087,N_6338);
nor U14078 (N_14078,N_8838,N_9897);
and U14079 (N_14079,N_6122,N_7433);
nand U14080 (N_14080,N_6041,N_7551);
or U14081 (N_14081,N_7540,N_9639);
or U14082 (N_14082,N_9390,N_5303);
nor U14083 (N_14083,N_9039,N_5256);
nor U14084 (N_14084,N_8039,N_7068);
xor U14085 (N_14085,N_9001,N_8841);
and U14086 (N_14086,N_5595,N_7608);
and U14087 (N_14087,N_8767,N_8725);
nand U14088 (N_14088,N_7195,N_8357);
nor U14089 (N_14089,N_7471,N_8774);
and U14090 (N_14090,N_6563,N_7994);
and U14091 (N_14091,N_9562,N_8313);
nand U14092 (N_14092,N_6447,N_8450);
nand U14093 (N_14093,N_7374,N_7678);
or U14094 (N_14094,N_8296,N_5970);
and U14095 (N_14095,N_8836,N_8395);
and U14096 (N_14096,N_8365,N_7268);
and U14097 (N_14097,N_5090,N_8226);
nor U14098 (N_14098,N_7995,N_8629);
nand U14099 (N_14099,N_7643,N_6189);
or U14100 (N_14100,N_6486,N_8593);
or U14101 (N_14101,N_5154,N_8050);
or U14102 (N_14102,N_7321,N_6014);
nand U14103 (N_14103,N_9464,N_6321);
or U14104 (N_14104,N_5157,N_9236);
nand U14105 (N_14105,N_9050,N_8737);
nand U14106 (N_14106,N_5547,N_5916);
and U14107 (N_14107,N_5135,N_7665);
nor U14108 (N_14108,N_9511,N_6724);
nand U14109 (N_14109,N_7224,N_7853);
and U14110 (N_14110,N_6330,N_8962);
and U14111 (N_14111,N_5779,N_9041);
nand U14112 (N_14112,N_9224,N_8392);
and U14113 (N_14113,N_5485,N_6802);
and U14114 (N_14114,N_9687,N_8940);
nor U14115 (N_14115,N_6234,N_6403);
or U14116 (N_14116,N_9111,N_8023);
or U14117 (N_14117,N_6252,N_7412);
nor U14118 (N_14118,N_5333,N_6522);
or U14119 (N_14119,N_9038,N_8099);
nor U14120 (N_14120,N_8896,N_9190);
or U14121 (N_14121,N_5224,N_9913);
xnor U14122 (N_14122,N_6172,N_5615);
nor U14123 (N_14123,N_7255,N_6097);
and U14124 (N_14124,N_9607,N_5757);
and U14125 (N_14125,N_6326,N_5943);
nor U14126 (N_14126,N_6993,N_9612);
nand U14127 (N_14127,N_7692,N_6673);
nor U14128 (N_14128,N_9742,N_7808);
or U14129 (N_14129,N_6595,N_8229);
and U14130 (N_14130,N_8452,N_6821);
nand U14131 (N_14131,N_9766,N_8970);
and U14132 (N_14132,N_6528,N_7527);
nor U14133 (N_14133,N_8512,N_5491);
or U14134 (N_14134,N_5633,N_5830);
nand U14135 (N_14135,N_9531,N_6631);
nor U14136 (N_14136,N_5739,N_9851);
and U14137 (N_14137,N_6603,N_5511);
or U14138 (N_14138,N_6637,N_9607);
or U14139 (N_14139,N_6556,N_7479);
nor U14140 (N_14140,N_6443,N_9783);
and U14141 (N_14141,N_9869,N_7185);
and U14142 (N_14142,N_8451,N_6208);
or U14143 (N_14143,N_7377,N_5183);
xor U14144 (N_14144,N_7854,N_9165);
nor U14145 (N_14145,N_6395,N_7117);
nand U14146 (N_14146,N_7808,N_7252);
nand U14147 (N_14147,N_8957,N_9775);
nand U14148 (N_14148,N_6154,N_8729);
nor U14149 (N_14149,N_9655,N_5691);
or U14150 (N_14150,N_9328,N_5104);
nor U14151 (N_14151,N_8633,N_5977);
nand U14152 (N_14152,N_7057,N_9144);
nand U14153 (N_14153,N_6330,N_5491);
or U14154 (N_14154,N_6648,N_8039);
nor U14155 (N_14155,N_8955,N_5042);
xnor U14156 (N_14156,N_6458,N_6840);
nand U14157 (N_14157,N_6548,N_9577);
nor U14158 (N_14158,N_8000,N_8149);
nand U14159 (N_14159,N_5395,N_6079);
nor U14160 (N_14160,N_6841,N_6079);
nor U14161 (N_14161,N_9641,N_8295);
nor U14162 (N_14162,N_5918,N_7666);
and U14163 (N_14163,N_9935,N_8092);
xor U14164 (N_14164,N_5078,N_5092);
nor U14165 (N_14165,N_5542,N_9222);
or U14166 (N_14166,N_7864,N_8819);
nand U14167 (N_14167,N_8998,N_9200);
or U14168 (N_14168,N_5439,N_5402);
nand U14169 (N_14169,N_9700,N_9177);
xor U14170 (N_14170,N_6382,N_5713);
or U14171 (N_14171,N_7629,N_5665);
or U14172 (N_14172,N_7239,N_9300);
nand U14173 (N_14173,N_8330,N_6209);
and U14174 (N_14174,N_7296,N_6012);
or U14175 (N_14175,N_9091,N_5009);
nor U14176 (N_14176,N_8983,N_9188);
nand U14177 (N_14177,N_6436,N_9362);
nand U14178 (N_14178,N_5956,N_8616);
or U14179 (N_14179,N_9005,N_6784);
nor U14180 (N_14180,N_6590,N_8241);
and U14181 (N_14181,N_7132,N_8164);
or U14182 (N_14182,N_9045,N_9249);
and U14183 (N_14183,N_8120,N_6764);
and U14184 (N_14184,N_9709,N_5003);
or U14185 (N_14185,N_5567,N_8975);
and U14186 (N_14186,N_5552,N_7725);
or U14187 (N_14187,N_9678,N_5400);
nor U14188 (N_14188,N_8046,N_6022);
or U14189 (N_14189,N_6972,N_6358);
or U14190 (N_14190,N_6833,N_9987);
and U14191 (N_14191,N_6189,N_6264);
or U14192 (N_14192,N_6570,N_9384);
nor U14193 (N_14193,N_6288,N_8156);
or U14194 (N_14194,N_5907,N_7947);
xor U14195 (N_14195,N_8808,N_8757);
or U14196 (N_14196,N_9877,N_8564);
or U14197 (N_14197,N_7180,N_5039);
nand U14198 (N_14198,N_8497,N_6558);
or U14199 (N_14199,N_5005,N_9367);
and U14200 (N_14200,N_7820,N_8611);
nor U14201 (N_14201,N_6509,N_5458);
nor U14202 (N_14202,N_7976,N_9735);
nand U14203 (N_14203,N_9340,N_9403);
and U14204 (N_14204,N_7049,N_9224);
nor U14205 (N_14205,N_7518,N_6111);
nor U14206 (N_14206,N_5234,N_6228);
and U14207 (N_14207,N_7940,N_6214);
and U14208 (N_14208,N_6606,N_7644);
and U14209 (N_14209,N_9930,N_6987);
nand U14210 (N_14210,N_9583,N_5987);
or U14211 (N_14211,N_9458,N_8786);
or U14212 (N_14212,N_5059,N_5233);
or U14213 (N_14213,N_6823,N_7170);
nand U14214 (N_14214,N_5084,N_8845);
and U14215 (N_14215,N_5273,N_5731);
and U14216 (N_14216,N_5112,N_9984);
and U14217 (N_14217,N_6279,N_5527);
or U14218 (N_14218,N_7615,N_5260);
nor U14219 (N_14219,N_5142,N_5600);
and U14220 (N_14220,N_6908,N_5248);
nand U14221 (N_14221,N_7622,N_7825);
nor U14222 (N_14222,N_7552,N_9426);
nor U14223 (N_14223,N_7521,N_8306);
and U14224 (N_14224,N_8887,N_9753);
xnor U14225 (N_14225,N_5822,N_5439);
nor U14226 (N_14226,N_5356,N_7251);
nor U14227 (N_14227,N_8531,N_9730);
and U14228 (N_14228,N_7787,N_7993);
nor U14229 (N_14229,N_6131,N_9825);
nand U14230 (N_14230,N_9136,N_6649);
nor U14231 (N_14231,N_6614,N_6207);
and U14232 (N_14232,N_9599,N_9692);
and U14233 (N_14233,N_5436,N_7062);
or U14234 (N_14234,N_7669,N_5778);
xor U14235 (N_14235,N_5716,N_9216);
nor U14236 (N_14236,N_7784,N_8042);
nor U14237 (N_14237,N_9792,N_9855);
or U14238 (N_14238,N_9272,N_8332);
or U14239 (N_14239,N_7002,N_9549);
nor U14240 (N_14240,N_7431,N_5118);
or U14241 (N_14241,N_9210,N_9300);
or U14242 (N_14242,N_9237,N_8109);
and U14243 (N_14243,N_9562,N_8557);
nand U14244 (N_14244,N_8317,N_9451);
and U14245 (N_14245,N_6100,N_7010);
and U14246 (N_14246,N_5794,N_9113);
and U14247 (N_14247,N_9051,N_8679);
nand U14248 (N_14248,N_8199,N_8641);
or U14249 (N_14249,N_9475,N_5819);
or U14250 (N_14250,N_8566,N_5244);
or U14251 (N_14251,N_7298,N_7532);
nor U14252 (N_14252,N_8578,N_5002);
nor U14253 (N_14253,N_8016,N_5909);
nand U14254 (N_14254,N_5321,N_6088);
and U14255 (N_14255,N_6764,N_6144);
and U14256 (N_14256,N_9186,N_8913);
and U14257 (N_14257,N_6436,N_9216);
or U14258 (N_14258,N_5846,N_9749);
nand U14259 (N_14259,N_6601,N_5716);
or U14260 (N_14260,N_5114,N_9136);
or U14261 (N_14261,N_5809,N_8432);
nor U14262 (N_14262,N_7529,N_7351);
and U14263 (N_14263,N_5967,N_5044);
or U14264 (N_14264,N_5506,N_6052);
nor U14265 (N_14265,N_6361,N_8915);
nor U14266 (N_14266,N_7431,N_7718);
and U14267 (N_14267,N_7190,N_6193);
xor U14268 (N_14268,N_7870,N_9337);
or U14269 (N_14269,N_5878,N_7846);
nor U14270 (N_14270,N_6537,N_7982);
or U14271 (N_14271,N_9181,N_8053);
and U14272 (N_14272,N_9421,N_9112);
nor U14273 (N_14273,N_8207,N_9391);
and U14274 (N_14274,N_7089,N_5465);
and U14275 (N_14275,N_8123,N_9629);
nor U14276 (N_14276,N_9519,N_5870);
and U14277 (N_14277,N_9758,N_9072);
nand U14278 (N_14278,N_5268,N_5431);
nor U14279 (N_14279,N_9154,N_8579);
nor U14280 (N_14280,N_7441,N_6934);
and U14281 (N_14281,N_5916,N_9077);
and U14282 (N_14282,N_6099,N_5277);
nor U14283 (N_14283,N_9868,N_7138);
nor U14284 (N_14284,N_5673,N_7553);
xnor U14285 (N_14285,N_6041,N_6521);
or U14286 (N_14286,N_6673,N_8115);
nor U14287 (N_14287,N_5569,N_5835);
and U14288 (N_14288,N_9920,N_7053);
nand U14289 (N_14289,N_6050,N_8548);
and U14290 (N_14290,N_9987,N_8406);
and U14291 (N_14291,N_5338,N_6730);
and U14292 (N_14292,N_8396,N_6020);
nand U14293 (N_14293,N_8387,N_6562);
nand U14294 (N_14294,N_8009,N_5311);
nand U14295 (N_14295,N_7460,N_9052);
nor U14296 (N_14296,N_6327,N_5754);
and U14297 (N_14297,N_7484,N_9632);
or U14298 (N_14298,N_8114,N_9338);
or U14299 (N_14299,N_6614,N_5754);
or U14300 (N_14300,N_8001,N_7536);
nand U14301 (N_14301,N_9626,N_7753);
nand U14302 (N_14302,N_6182,N_5213);
nand U14303 (N_14303,N_7956,N_5646);
and U14304 (N_14304,N_9405,N_8543);
nor U14305 (N_14305,N_7640,N_9279);
nor U14306 (N_14306,N_7976,N_6865);
or U14307 (N_14307,N_5279,N_6446);
and U14308 (N_14308,N_9856,N_5552);
nor U14309 (N_14309,N_9346,N_5249);
or U14310 (N_14310,N_6890,N_7417);
nand U14311 (N_14311,N_9821,N_5292);
nand U14312 (N_14312,N_8598,N_8418);
and U14313 (N_14313,N_6480,N_7123);
nand U14314 (N_14314,N_8424,N_5135);
nor U14315 (N_14315,N_7687,N_6399);
nand U14316 (N_14316,N_8002,N_5408);
and U14317 (N_14317,N_6925,N_7959);
or U14318 (N_14318,N_6631,N_8637);
xor U14319 (N_14319,N_9418,N_5325);
or U14320 (N_14320,N_9832,N_8623);
or U14321 (N_14321,N_8447,N_7967);
and U14322 (N_14322,N_8614,N_8198);
nor U14323 (N_14323,N_8115,N_5147);
or U14324 (N_14324,N_5630,N_6910);
nor U14325 (N_14325,N_5790,N_6089);
nand U14326 (N_14326,N_9419,N_6820);
or U14327 (N_14327,N_9431,N_6552);
or U14328 (N_14328,N_8924,N_8807);
nand U14329 (N_14329,N_9439,N_5874);
nor U14330 (N_14330,N_7882,N_8241);
or U14331 (N_14331,N_5765,N_6506);
nor U14332 (N_14332,N_7494,N_8648);
nor U14333 (N_14333,N_8738,N_7502);
nand U14334 (N_14334,N_6348,N_7438);
or U14335 (N_14335,N_6230,N_8675);
or U14336 (N_14336,N_5411,N_9217);
and U14337 (N_14337,N_7321,N_5785);
and U14338 (N_14338,N_6555,N_9654);
and U14339 (N_14339,N_7787,N_6302);
nor U14340 (N_14340,N_7275,N_5764);
nor U14341 (N_14341,N_9166,N_8480);
and U14342 (N_14342,N_8675,N_6624);
nor U14343 (N_14343,N_7683,N_5794);
nor U14344 (N_14344,N_7204,N_7597);
nand U14345 (N_14345,N_5813,N_5667);
nor U14346 (N_14346,N_6001,N_8543);
and U14347 (N_14347,N_6586,N_6631);
nor U14348 (N_14348,N_8293,N_7591);
nor U14349 (N_14349,N_7162,N_8548);
and U14350 (N_14350,N_9058,N_6083);
or U14351 (N_14351,N_5629,N_5283);
nand U14352 (N_14352,N_8435,N_6108);
or U14353 (N_14353,N_8488,N_9387);
nand U14354 (N_14354,N_9583,N_9493);
xor U14355 (N_14355,N_7364,N_7149);
xor U14356 (N_14356,N_8885,N_5841);
or U14357 (N_14357,N_9861,N_7685);
nor U14358 (N_14358,N_7742,N_8515);
and U14359 (N_14359,N_7122,N_6032);
nor U14360 (N_14360,N_9158,N_6156);
nor U14361 (N_14361,N_8252,N_6448);
or U14362 (N_14362,N_7820,N_6428);
nand U14363 (N_14363,N_5043,N_5887);
nor U14364 (N_14364,N_9981,N_5566);
and U14365 (N_14365,N_5918,N_7558);
or U14366 (N_14366,N_5949,N_7166);
nor U14367 (N_14367,N_8541,N_8273);
nor U14368 (N_14368,N_8907,N_6082);
or U14369 (N_14369,N_5722,N_6645);
nor U14370 (N_14370,N_9042,N_7465);
nor U14371 (N_14371,N_8330,N_9576);
and U14372 (N_14372,N_6717,N_7482);
nor U14373 (N_14373,N_5232,N_7264);
and U14374 (N_14374,N_9386,N_5985);
nand U14375 (N_14375,N_9847,N_7933);
or U14376 (N_14376,N_6034,N_9876);
xor U14377 (N_14377,N_7525,N_6273);
and U14378 (N_14378,N_6017,N_7294);
or U14379 (N_14379,N_9059,N_5266);
or U14380 (N_14380,N_7911,N_8461);
nor U14381 (N_14381,N_8206,N_6524);
or U14382 (N_14382,N_7775,N_5428);
and U14383 (N_14383,N_6322,N_6400);
xnor U14384 (N_14384,N_7701,N_6686);
nor U14385 (N_14385,N_8531,N_8000);
and U14386 (N_14386,N_9535,N_5794);
and U14387 (N_14387,N_9526,N_9503);
or U14388 (N_14388,N_5111,N_5397);
nand U14389 (N_14389,N_6230,N_5580);
and U14390 (N_14390,N_8362,N_9925);
and U14391 (N_14391,N_9959,N_5006);
nand U14392 (N_14392,N_9942,N_6269);
nand U14393 (N_14393,N_6548,N_6311);
and U14394 (N_14394,N_5044,N_6790);
or U14395 (N_14395,N_6463,N_5811);
and U14396 (N_14396,N_8754,N_9737);
xnor U14397 (N_14397,N_8560,N_5671);
nor U14398 (N_14398,N_7758,N_8715);
nand U14399 (N_14399,N_7183,N_9611);
nand U14400 (N_14400,N_5346,N_5015);
or U14401 (N_14401,N_9108,N_6600);
and U14402 (N_14402,N_8505,N_9900);
or U14403 (N_14403,N_6923,N_8727);
nand U14404 (N_14404,N_7701,N_8577);
nor U14405 (N_14405,N_5216,N_9458);
nor U14406 (N_14406,N_8361,N_9126);
nand U14407 (N_14407,N_6748,N_9063);
nor U14408 (N_14408,N_5758,N_7972);
nor U14409 (N_14409,N_5601,N_6664);
or U14410 (N_14410,N_8172,N_8649);
nand U14411 (N_14411,N_9783,N_9603);
nand U14412 (N_14412,N_7812,N_8794);
nor U14413 (N_14413,N_9594,N_9510);
or U14414 (N_14414,N_7731,N_9977);
nor U14415 (N_14415,N_7916,N_8498);
or U14416 (N_14416,N_7899,N_6028);
and U14417 (N_14417,N_9056,N_5837);
or U14418 (N_14418,N_8146,N_5385);
nand U14419 (N_14419,N_5969,N_7259);
or U14420 (N_14420,N_5191,N_8006);
and U14421 (N_14421,N_8014,N_6669);
nand U14422 (N_14422,N_9654,N_9301);
and U14423 (N_14423,N_5486,N_9799);
nand U14424 (N_14424,N_7391,N_9323);
nand U14425 (N_14425,N_6751,N_8497);
nand U14426 (N_14426,N_9229,N_5785);
and U14427 (N_14427,N_8310,N_6740);
or U14428 (N_14428,N_6458,N_9744);
and U14429 (N_14429,N_6281,N_8869);
xnor U14430 (N_14430,N_9521,N_5525);
and U14431 (N_14431,N_8107,N_8559);
or U14432 (N_14432,N_5464,N_5072);
or U14433 (N_14433,N_8761,N_5447);
nand U14434 (N_14434,N_5024,N_8662);
nor U14435 (N_14435,N_9640,N_8050);
and U14436 (N_14436,N_6430,N_8453);
and U14437 (N_14437,N_8253,N_5878);
nor U14438 (N_14438,N_5653,N_5950);
nor U14439 (N_14439,N_5335,N_5845);
nor U14440 (N_14440,N_9465,N_8921);
nor U14441 (N_14441,N_5625,N_7551);
nor U14442 (N_14442,N_7698,N_7929);
nor U14443 (N_14443,N_9566,N_9767);
nand U14444 (N_14444,N_9898,N_9210);
or U14445 (N_14445,N_5984,N_8015);
nor U14446 (N_14446,N_5322,N_8292);
or U14447 (N_14447,N_9992,N_7463);
or U14448 (N_14448,N_7252,N_9342);
or U14449 (N_14449,N_5268,N_7324);
and U14450 (N_14450,N_9838,N_5624);
and U14451 (N_14451,N_7130,N_8256);
or U14452 (N_14452,N_8277,N_7111);
or U14453 (N_14453,N_9458,N_7884);
nor U14454 (N_14454,N_7305,N_8557);
and U14455 (N_14455,N_9629,N_6569);
and U14456 (N_14456,N_7940,N_5251);
or U14457 (N_14457,N_6359,N_8249);
or U14458 (N_14458,N_9535,N_6295);
nand U14459 (N_14459,N_9536,N_7075);
and U14460 (N_14460,N_8569,N_9036);
or U14461 (N_14461,N_8362,N_5548);
and U14462 (N_14462,N_8953,N_7675);
nand U14463 (N_14463,N_5917,N_5325);
nand U14464 (N_14464,N_9959,N_6335);
and U14465 (N_14465,N_7639,N_7569);
or U14466 (N_14466,N_5851,N_9218);
or U14467 (N_14467,N_9773,N_7681);
or U14468 (N_14468,N_6895,N_7619);
or U14469 (N_14469,N_9831,N_6494);
nand U14470 (N_14470,N_7081,N_5847);
or U14471 (N_14471,N_6313,N_6731);
nand U14472 (N_14472,N_9384,N_7830);
nor U14473 (N_14473,N_5442,N_8585);
and U14474 (N_14474,N_9046,N_6393);
nor U14475 (N_14475,N_9525,N_8688);
nor U14476 (N_14476,N_7044,N_8118);
or U14477 (N_14477,N_5629,N_5748);
nand U14478 (N_14478,N_5033,N_5168);
nor U14479 (N_14479,N_8996,N_7764);
and U14480 (N_14480,N_6134,N_7738);
or U14481 (N_14481,N_7892,N_9901);
or U14482 (N_14482,N_8025,N_7727);
and U14483 (N_14483,N_9248,N_7095);
nor U14484 (N_14484,N_6335,N_6989);
nor U14485 (N_14485,N_5197,N_9746);
nor U14486 (N_14486,N_6711,N_9912);
nor U14487 (N_14487,N_9991,N_8374);
and U14488 (N_14488,N_6948,N_9059);
nand U14489 (N_14489,N_5423,N_6587);
nor U14490 (N_14490,N_5376,N_7688);
and U14491 (N_14491,N_9123,N_8173);
and U14492 (N_14492,N_7568,N_6865);
and U14493 (N_14493,N_6505,N_9570);
nor U14494 (N_14494,N_9831,N_9497);
and U14495 (N_14495,N_9911,N_6061);
nor U14496 (N_14496,N_6783,N_9063);
nand U14497 (N_14497,N_9098,N_7439);
nor U14498 (N_14498,N_5114,N_6417);
nor U14499 (N_14499,N_6224,N_5597);
nand U14500 (N_14500,N_9658,N_9175);
or U14501 (N_14501,N_6576,N_7199);
nand U14502 (N_14502,N_7118,N_7172);
nor U14503 (N_14503,N_7045,N_7420);
nand U14504 (N_14504,N_9675,N_8919);
or U14505 (N_14505,N_8351,N_6568);
and U14506 (N_14506,N_5063,N_9248);
or U14507 (N_14507,N_5945,N_5289);
nand U14508 (N_14508,N_7903,N_8886);
nor U14509 (N_14509,N_9305,N_9564);
or U14510 (N_14510,N_5995,N_8184);
nor U14511 (N_14511,N_6407,N_6437);
nor U14512 (N_14512,N_5289,N_9839);
nand U14513 (N_14513,N_7604,N_5905);
and U14514 (N_14514,N_5623,N_5348);
or U14515 (N_14515,N_9295,N_5669);
nand U14516 (N_14516,N_7794,N_6721);
nor U14517 (N_14517,N_6713,N_6526);
xor U14518 (N_14518,N_6485,N_5765);
nor U14519 (N_14519,N_7979,N_8300);
or U14520 (N_14520,N_6837,N_8952);
nor U14521 (N_14521,N_9252,N_9593);
or U14522 (N_14522,N_8303,N_8891);
and U14523 (N_14523,N_6940,N_5399);
nor U14524 (N_14524,N_5647,N_7207);
nor U14525 (N_14525,N_8391,N_9969);
nand U14526 (N_14526,N_7748,N_9960);
or U14527 (N_14527,N_7803,N_6602);
and U14528 (N_14528,N_5136,N_6554);
and U14529 (N_14529,N_7555,N_7946);
nor U14530 (N_14530,N_9378,N_7278);
and U14531 (N_14531,N_6862,N_6653);
nand U14532 (N_14532,N_6785,N_9645);
and U14533 (N_14533,N_8462,N_8758);
nand U14534 (N_14534,N_8528,N_9380);
nand U14535 (N_14535,N_8014,N_8313);
or U14536 (N_14536,N_6373,N_7591);
nor U14537 (N_14537,N_8987,N_7557);
nand U14538 (N_14538,N_5420,N_5814);
nand U14539 (N_14539,N_8474,N_9978);
and U14540 (N_14540,N_6213,N_5801);
nand U14541 (N_14541,N_8829,N_6231);
nand U14542 (N_14542,N_6296,N_7740);
and U14543 (N_14543,N_7944,N_5491);
nor U14544 (N_14544,N_7430,N_6350);
and U14545 (N_14545,N_9604,N_8884);
and U14546 (N_14546,N_8870,N_8553);
nand U14547 (N_14547,N_5364,N_6686);
and U14548 (N_14548,N_5665,N_8335);
xor U14549 (N_14549,N_9251,N_8951);
nand U14550 (N_14550,N_6391,N_7374);
nor U14551 (N_14551,N_6648,N_5607);
nand U14552 (N_14552,N_9480,N_9839);
and U14553 (N_14553,N_5004,N_9133);
nor U14554 (N_14554,N_8955,N_6928);
nand U14555 (N_14555,N_8261,N_9225);
or U14556 (N_14556,N_8313,N_7549);
and U14557 (N_14557,N_9916,N_5265);
nand U14558 (N_14558,N_8903,N_8592);
and U14559 (N_14559,N_9748,N_7870);
or U14560 (N_14560,N_8987,N_5579);
and U14561 (N_14561,N_7282,N_6500);
nand U14562 (N_14562,N_8749,N_9011);
nand U14563 (N_14563,N_7829,N_9547);
nand U14564 (N_14564,N_5334,N_5164);
nand U14565 (N_14565,N_7374,N_8429);
nand U14566 (N_14566,N_8673,N_9793);
nand U14567 (N_14567,N_9062,N_6035);
and U14568 (N_14568,N_8954,N_9457);
nand U14569 (N_14569,N_7921,N_6794);
nor U14570 (N_14570,N_9775,N_9393);
nor U14571 (N_14571,N_5880,N_7169);
xnor U14572 (N_14572,N_8621,N_6486);
nor U14573 (N_14573,N_9131,N_5504);
nor U14574 (N_14574,N_5579,N_5924);
xor U14575 (N_14575,N_8139,N_8342);
and U14576 (N_14576,N_7106,N_9392);
and U14577 (N_14577,N_5654,N_5167);
nor U14578 (N_14578,N_9474,N_6501);
or U14579 (N_14579,N_5492,N_8033);
xor U14580 (N_14580,N_5680,N_6677);
nand U14581 (N_14581,N_5549,N_8707);
nand U14582 (N_14582,N_9865,N_8978);
nand U14583 (N_14583,N_7107,N_9877);
or U14584 (N_14584,N_8325,N_5276);
nand U14585 (N_14585,N_8388,N_5625);
nor U14586 (N_14586,N_6021,N_6250);
nand U14587 (N_14587,N_6578,N_9791);
and U14588 (N_14588,N_9056,N_5484);
nor U14589 (N_14589,N_8440,N_9038);
nor U14590 (N_14590,N_5285,N_5215);
and U14591 (N_14591,N_7680,N_8791);
nor U14592 (N_14592,N_5774,N_8260);
and U14593 (N_14593,N_7761,N_9971);
or U14594 (N_14594,N_9390,N_8787);
nand U14595 (N_14595,N_7773,N_7086);
nand U14596 (N_14596,N_5316,N_9435);
nor U14597 (N_14597,N_6538,N_6695);
and U14598 (N_14598,N_8907,N_9271);
nand U14599 (N_14599,N_6275,N_5527);
nor U14600 (N_14600,N_9116,N_5177);
nor U14601 (N_14601,N_7408,N_6276);
or U14602 (N_14602,N_7068,N_7824);
and U14603 (N_14603,N_6786,N_7388);
or U14604 (N_14604,N_6985,N_6847);
nor U14605 (N_14605,N_8198,N_7702);
nor U14606 (N_14606,N_8418,N_5642);
nor U14607 (N_14607,N_8909,N_5581);
nor U14608 (N_14608,N_5596,N_7385);
and U14609 (N_14609,N_9172,N_6729);
nand U14610 (N_14610,N_8304,N_7215);
nand U14611 (N_14611,N_6948,N_9123);
or U14612 (N_14612,N_8688,N_5128);
or U14613 (N_14613,N_6466,N_9405);
and U14614 (N_14614,N_8836,N_7498);
nand U14615 (N_14615,N_6518,N_6175);
nor U14616 (N_14616,N_5886,N_9618);
nor U14617 (N_14617,N_6385,N_6421);
nand U14618 (N_14618,N_8025,N_9448);
nor U14619 (N_14619,N_8124,N_7109);
nor U14620 (N_14620,N_6128,N_7199);
nand U14621 (N_14621,N_9189,N_7449);
nor U14622 (N_14622,N_8322,N_6769);
xor U14623 (N_14623,N_5037,N_7561);
or U14624 (N_14624,N_8465,N_7829);
nand U14625 (N_14625,N_6240,N_6908);
or U14626 (N_14626,N_9122,N_8701);
nand U14627 (N_14627,N_7179,N_6224);
and U14628 (N_14628,N_8138,N_6909);
and U14629 (N_14629,N_5025,N_5033);
nor U14630 (N_14630,N_6943,N_5494);
nor U14631 (N_14631,N_9341,N_9989);
nor U14632 (N_14632,N_9181,N_7985);
xnor U14633 (N_14633,N_6769,N_6015);
nor U14634 (N_14634,N_8016,N_9107);
or U14635 (N_14635,N_5599,N_8181);
nand U14636 (N_14636,N_6969,N_6849);
nor U14637 (N_14637,N_6614,N_9959);
and U14638 (N_14638,N_9817,N_8712);
or U14639 (N_14639,N_6055,N_9433);
nor U14640 (N_14640,N_8806,N_7532);
nand U14641 (N_14641,N_7214,N_7301);
or U14642 (N_14642,N_9444,N_6330);
and U14643 (N_14643,N_6024,N_6349);
and U14644 (N_14644,N_5644,N_7282);
nand U14645 (N_14645,N_6862,N_9663);
nor U14646 (N_14646,N_5067,N_8238);
and U14647 (N_14647,N_6793,N_8540);
nand U14648 (N_14648,N_9862,N_5638);
nor U14649 (N_14649,N_5262,N_7250);
nor U14650 (N_14650,N_9487,N_8178);
and U14651 (N_14651,N_9795,N_7201);
nor U14652 (N_14652,N_7104,N_7136);
nand U14653 (N_14653,N_7910,N_7769);
nand U14654 (N_14654,N_5879,N_5704);
nand U14655 (N_14655,N_6159,N_6632);
and U14656 (N_14656,N_8995,N_5388);
nand U14657 (N_14657,N_9591,N_9422);
nor U14658 (N_14658,N_8148,N_5837);
nor U14659 (N_14659,N_6592,N_8401);
nand U14660 (N_14660,N_9552,N_9887);
nor U14661 (N_14661,N_9934,N_7156);
nor U14662 (N_14662,N_7065,N_8651);
and U14663 (N_14663,N_8499,N_5198);
nor U14664 (N_14664,N_5220,N_5269);
nor U14665 (N_14665,N_9454,N_6588);
nor U14666 (N_14666,N_7650,N_6183);
and U14667 (N_14667,N_8226,N_7132);
nand U14668 (N_14668,N_5516,N_6688);
nor U14669 (N_14669,N_8562,N_9786);
nor U14670 (N_14670,N_6858,N_7018);
or U14671 (N_14671,N_9038,N_6256);
xor U14672 (N_14672,N_8746,N_5479);
nand U14673 (N_14673,N_5508,N_9336);
or U14674 (N_14674,N_6147,N_7842);
and U14675 (N_14675,N_7201,N_9256);
or U14676 (N_14676,N_7863,N_8981);
or U14677 (N_14677,N_5505,N_6240);
or U14678 (N_14678,N_7502,N_9058);
and U14679 (N_14679,N_6705,N_6929);
nor U14680 (N_14680,N_5433,N_9622);
nand U14681 (N_14681,N_9456,N_6830);
or U14682 (N_14682,N_9473,N_9027);
and U14683 (N_14683,N_6044,N_9960);
nor U14684 (N_14684,N_6425,N_7169);
and U14685 (N_14685,N_5033,N_9627);
nor U14686 (N_14686,N_6303,N_5271);
and U14687 (N_14687,N_8813,N_6878);
nor U14688 (N_14688,N_6278,N_7707);
nand U14689 (N_14689,N_7885,N_8571);
and U14690 (N_14690,N_8444,N_8327);
nand U14691 (N_14691,N_7964,N_9213);
nor U14692 (N_14692,N_6093,N_7916);
nor U14693 (N_14693,N_6013,N_5224);
and U14694 (N_14694,N_6999,N_7931);
or U14695 (N_14695,N_6660,N_6149);
or U14696 (N_14696,N_8666,N_8915);
nor U14697 (N_14697,N_6742,N_8115);
and U14698 (N_14698,N_9049,N_7781);
nand U14699 (N_14699,N_9263,N_5703);
and U14700 (N_14700,N_8765,N_8171);
nand U14701 (N_14701,N_9440,N_9702);
nand U14702 (N_14702,N_7504,N_9309);
nor U14703 (N_14703,N_9215,N_6325);
and U14704 (N_14704,N_8384,N_6539);
and U14705 (N_14705,N_7840,N_9601);
or U14706 (N_14706,N_6308,N_9061);
nand U14707 (N_14707,N_7620,N_6341);
nand U14708 (N_14708,N_9013,N_9463);
nor U14709 (N_14709,N_9329,N_8453);
and U14710 (N_14710,N_8710,N_5487);
nor U14711 (N_14711,N_8015,N_7208);
nand U14712 (N_14712,N_7985,N_7099);
nor U14713 (N_14713,N_8087,N_6238);
or U14714 (N_14714,N_7272,N_7655);
nor U14715 (N_14715,N_8373,N_7557);
or U14716 (N_14716,N_9977,N_6392);
nand U14717 (N_14717,N_6185,N_7958);
xor U14718 (N_14718,N_7717,N_9061);
and U14719 (N_14719,N_7367,N_5093);
nor U14720 (N_14720,N_5328,N_6374);
and U14721 (N_14721,N_9970,N_7443);
nor U14722 (N_14722,N_8550,N_7504);
or U14723 (N_14723,N_7324,N_7316);
xor U14724 (N_14724,N_7303,N_5980);
xnor U14725 (N_14725,N_9086,N_5204);
nand U14726 (N_14726,N_9955,N_9148);
nor U14727 (N_14727,N_9693,N_5752);
nor U14728 (N_14728,N_5185,N_9655);
nand U14729 (N_14729,N_6557,N_5014);
nor U14730 (N_14730,N_9800,N_5487);
or U14731 (N_14731,N_7231,N_7130);
nand U14732 (N_14732,N_6331,N_5386);
nand U14733 (N_14733,N_8346,N_6447);
nand U14734 (N_14734,N_7559,N_7643);
nand U14735 (N_14735,N_7084,N_6063);
nor U14736 (N_14736,N_7062,N_9072);
xor U14737 (N_14737,N_8689,N_6659);
and U14738 (N_14738,N_7564,N_8157);
nor U14739 (N_14739,N_7863,N_9906);
nor U14740 (N_14740,N_5415,N_5947);
nor U14741 (N_14741,N_8948,N_5713);
nor U14742 (N_14742,N_7857,N_5110);
nor U14743 (N_14743,N_9916,N_9564);
and U14744 (N_14744,N_5689,N_7240);
nor U14745 (N_14745,N_9044,N_8835);
and U14746 (N_14746,N_9188,N_9654);
nor U14747 (N_14747,N_6224,N_5811);
nand U14748 (N_14748,N_8298,N_5663);
nand U14749 (N_14749,N_8170,N_8006);
and U14750 (N_14750,N_6694,N_9712);
and U14751 (N_14751,N_5715,N_7092);
or U14752 (N_14752,N_7441,N_9922);
nand U14753 (N_14753,N_7040,N_9867);
or U14754 (N_14754,N_7089,N_8460);
or U14755 (N_14755,N_5165,N_5561);
xnor U14756 (N_14756,N_7345,N_5132);
nand U14757 (N_14757,N_6622,N_9689);
nor U14758 (N_14758,N_6363,N_5239);
and U14759 (N_14759,N_9547,N_8407);
nor U14760 (N_14760,N_9144,N_6847);
nor U14761 (N_14761,N_9932,N_5847);
nand U14762 (N_14762,N_6099,N_6765);
nor U14763 (N_14763,N_8639,N_5187);
nand U14764 (N_14764,N_8398,N_9644);
or U14765 (N_14765,N_9344,N_8854);
or U14766 (N_14766,N_6950,N_8151);
nor U14767 (N_14767,N_8433,N_8753);
or U14768 (N_14768,N_5905,N_9763);
nand U14769 (N_14769,N_9495,N_5548);
xor U14770 (N_14770,N_9199,N_9142);
nor U14771 (N_14771,N_5320,N_9987);
nor U14772 (N_14772,N_5815,N_7734);
nand U14773 (N_14773,N_7318,N_8509);
and U14774 (N_14774,N_7223,N_8091);
or U14775 (N_14775,N_8490,N_8463);
and U14776 (N_14776,N_8744,N_5192);
and U14777 (N_14777,N_7346,N_7057);
or U14778 (N_14778,N_7221,N_9313);
nand U14779 (N_14779,N_8521,N_5512);
nand U14780 (N_14780,N_9601,N_8095);
and U14781 (N_14781,N_9416,N_8864);
or U14782 (N_14782,N_7695,N_5897);
nand U14783 (N_14783,N_8771,N_7205);
nand U14784 (N_14784,N_9287,N_6593);
nor U14785 (N_14785,N_9235,N_5999);
or U14786 (N_14786,N_7635,N_6636);
or U14787 (N_14787,N_7401,N_6352);
nor U14788 (N_14788,N_9428,N_5524);
and U14789 (N_14789,N_7077,N_8672);
nand U14790 (N_14790,N_9477,N_9067);
or U14791 (N_14791,N_5631,N_8158);
nor U14792 (N_14792,N_5816,N_9239);
nor U14793 (N_14793,N_9073,N_8803);
nor U14794 (N_14794,N_6810,N_7045);
nor U14795 (N_14795,N_9435,N_6202);
or U14796 (N_14796,N_7095,N_6938);
or U14797 (N_14797,N_9241,N_8663);
or U14798 (N_14798,N_8664,N_7827);
nand U14799 (N_14799,N_6960,N_9349);
nand U14800 (N_14800,N_6698,N_7238);
nand U14801 (N_14801,N_7719,N_8318);
nor U14802 (N_14802,N_9118,N_9548);
and U14803 (N_14803,N_7482,N_6450);
or U14804 (N_14804,N_6568,N_6091);
and U14805 (N_14805,N_7934,N_5691);
nand U14806 (N_14806,N_5948,N_6959);
nand U14807 (N_14807,N_7280,N_8136);
nand U14808 (N_14808,N_6176,N_7993);
nor U14809 (N_14809,N_8382,N_5549);
or U14810 (N_14810,N_7273,N_6618);
nand U14811 (N_14811,N_5584,N_5970);
nand U14812 (N_14812,N_5006,N_9198);
and U14813 (N_14813,N_6693,N_7412);
nand U14814 (N_14814,N_6709,N_9626);
nor U14815 (N_14815,N_5713,N_7901);
nand U14816 (N_14816,N_6913,N_7716);
nor U14817 (N_14817,N_7806,N_9336);
nand U14818 (N_14818,N_7920,N_5759);
or U14819 (N_14819,N_6587,N_6469);
nand U14820 (N_14820,N_9157,N_5827);
and U14821 (N_14821,N_8268,N_5190);
nor U14822 (N_14822,N_8743,N_8676);
nor U14823 (N_14823,N_9592,N_6688);
nand U14824 (N_14824,N_8620,N_9891);
and U14825 (N_14825,N_8772,N_9698);
nor U14826 (N_14826,N_6091,N_5073);
or U14827 (N_14827,N_5570,N_7503);
or U14828 (N_14828,N_9718,N_8826);
nor U14829 (N_14829,N_7523,N_8608);
nor U14830 (N_14830,N_6238,N_7305);
nand U14831 (N_14831,N_9555,N_8887);
nor U14832 (N_14832,N_7392,N_5590);
and U14833 (N_14833,N_6141,N_8302);
and U14834 (N_14834,N_8989,N_8587);
nor U14835 (N_14835,N_9119,N_9413);
xor U14836 (N_14836,N_7155,N_9873);
nor U14837 (N_14837,N_6291,N_9516);
nor U14838 (N_14838,N_9448,N_9133);
nand U14839 (N_14839,N_9296,N_8434);
nor U14840 (N_14840,N_8526,N_6198);
and U14841 (N_14841,N_8956,N_9217);
nor U14842 (N_14842,N_7016,N_9195);
and U14843 (N_14843,N_8990,N_7812);
or U14844 (N_14844,N_8132,N_9481);
or U14845 (N_14845,N_9772,N_5431);
or U14846 (N_14846,N_8202,N_5856);
and U14847 (N_14847,N_5724,N_7388);
nand U14848 (N_14848,N_9429,N_6064);
nor U14849 (N_14849,N_9873,N_8920);
nand U14850 (N_14850,N_6218,N_7172);
and U14851 (N_14851,N_6747,N_6920);
nor U14852 (N_14852,N_9590,N_5914);
nand U14853 (N_14853,N_9615,N_7319);
nor U14854 (N_14854,N_8014,N_7087);
or U14855 (N_14855,N_6117,N_8495);
or U14856 (N_14856,N_9007,N_5460);
and U14857 (N_14857,N_9579,N_9697);
nand U14858 (N_14858,N_5450,N_7849);
or U14859 (N_14859,N_6400,N_6695);
nand U14860 (N_14860,N_7101,N_7560);
nor U14861 (N_14861,N_7284,N_9563);
nand U14862 (N_14862,N_6985,N_5439);
nor U14863 (N_14863,N_6533,N_6199);
nand U14864 (N_14864,N_8650,N_7152);
nor U14865 (N_14865,N_8536,N_7979);
or U14866 (N_14866,N_7219,N_6831);
or U14867 (N_14867,N_5162,N_8241);
or U14868 (N_14868,N_7435,N_7579);
or U14869 (N_14869,N_9884,N_8055);
nor U14870 (N_14870,N_6049,N_9369);
and U14871 (N_14871,N_8669,N_7993);
and U14872 (N_14872,N_9282,N_6593);
nor U14873 (N_14873,N_9962,N_5666);
nand U14874 (N_14874,N_5991,N_5897);
nor U14875 (N_14875,N_7992,N_9406);
nand U14876 (N_14876,N_9663,N_8633);
nor U14877 (N_14877,N_7879,N_7321);
xor U14878 (N_14878,N_7917,N_9762);
nand U14879 (N_14879,N_8710,N_6279);
xor U14880 (N_14880,N_9913,N_8265);
nand U14881 (N_14881,N_7662,N_5922);
and U14882 (N_14882,N_6111,N_7354);
or U14883 (N_14883,N_8369,N_7808);
and U14884 (N_14884,N_9260,N_9783);
nor U14885 (N_14885,N_5642,N_5850);
nand U14886 (N_14886,N_7469,N_9748);
or U14887 (N_14887,N_9993,N_7239);
nand U14888 (N_14888,N_5147,N_9686);
nand U14889 (N_14889,N_7995,N_6450);
and U14890 (N_14890,N_6456,N_6092);
or U14891 (N_14891,N_6596,N_7785);
and U14892 (N_14892,N_5347,N_5977);
nand U14893 (N_14893,N_7641,N_9430);
or U14894 (N_14894,N_7687,N_6980);
and U14895 (N_14895,N_7879,N_7254);
nor U14896 (N_14896,N_8659,N_6655);
nand U14897 (N_14897,N_8086,N_7024);
nand U14898 (N_14898,N_7849,N_5546);
nor U14899 (N_14899,N_7357,N_5288);
or U14900 (N_14900,N_7847,N_9016);
or U14901 (N_14901,N_8419,N_7787);
and U14902 (N_14902,N_9475,N_8334);
and U14903 (N_14903,N_5355,N_6138);
or U14904 (N_14904,N_7906,N_5598);
and U14905 (N_14905,N_9347,N_6964);
nand U14906 (N_14906,N_8866,N_7774);
and U14907 (N_14907,N_5477,N_5335);
or U14908 (N_14908,N_5500,N_9757);
nor U14909 (N_14909,N_6235,N_9799);
nor U14910 (N_14910,N_6820,N_9828);
or U14911 (N_14911,N_5096,N_5621);
nand U14912 (N_14912,N_7719,N_9475);
nand U14913 (N_14913,N_6176,N_9649);
nor U14914 (N_14914,N_7086,N_5799);
and U14915 (N_14915,N_8393,N_8501);
nand U14916 (N_14916,N_8938,N_8724);
nor U14917 (N_14917,N_7862,N_9388);
xor U14918 (N_14918,N_5795,N_5808);
or U14919 (N_14919,N_5550,N_7036);
and U14920 (N_14920,N_9555,N_5325);
nor U14921 (N_14921,N_9988,N_7637);
or U14922 (N_14922,N_5872,N_8373);
nor U14923 (N_14923,N_9870,N_8101);
nand U14924 (N_14924,N_6514,N_5657);
nand U14925 (N_14925,N_8767,N_9907);
nor U14926 (N_14926,N_5132,N_5039);
nor U14927 (N_14927,N_6867,N_7948);
nand U14928 (N_14928,N_7402,N_8339);
nor U14929 (N_14929,N_5364,N_6799);
nand U14930 (N_14930,N_5789,N_5919);
and U14931 (N_14931,N_8584,N_6734);
or U14932 (N_14932,N_8855,N_6508);
xnor U14933 (N_14933,N_9898,N_6617);
or U14934 (N_14934,N_7903,N_9001);
nor U14935 (N_14935,N_7172,N_6140);
nand U14936 (N_14936,N_5582,N_9062);
or U14937 (N_14937,N_9336,N_5672);
or U14938 (N_14938,N_5579,N_9115);
nor U14939 (N_14939,N_9567,N_5164);
or U14940 (N_14940,N_9641,N_8244);
or U14941 (N_14941,N_6841,N_9603);
and U14942 (N_14942,N_8285,N_5394);
or U14943 (N_14943,N_6339,N_9561);
nor U14944 (N_14944,N_9887,N_7212);
and U14945 (N_14945,N_5552,N_8930);
and U14946 (N_14946,N_7055,N_5787);
nor U14947 (N_14947,N_9167,N_6232);
nor U14948 (N_14948,N_7418,N_7261);
and U14949 (N_14949,N_8727,N_9343);
or U14950 (N_14950,N_7002,N_5200);
or U14951 (N_14951,N_8211,N_8547);
and U14952 (N_14952,N_9552,N_5091);
nand U14953 (N_14953,N_6654,N_5190);
and U14954 (N_14954,N_8140,N_6833);
nand U14955 (N_14955,N_6922,N_6149);
nor U14956 (N_14956,N_8251,N_7500);
nor U14957 (N_14957,N_5046,N_5963);
nand U14958 (N_14958,N_8998,N_6691);
or U14959 (N_14959,N_5167,N_7852);
and U14960 (N_14960,N_7963,N_7752);
and U14961 (N_14961,N_7189,N_5962);
or U14962 (N_14962,N_8061,N_8976);
nand U14963 (N_14963,N_6736,N_9550);
nand U14964 (N_14964,N_7092,N_9933);
nor U14965 (N_14965,N_6679,N_9276);
and U14966 (N_14966,N_5362,N_7529);
nand U14967 (N_14967,N_6442,N_7416);
xnor U14968 (N_14968,N_5745,N_5094);
nor U14969 (N_14969,N_8968,N_5716);
nor U14970 (N_14970,N_5386,N_9196);
xor U14971 (N_14971,N_6603,N_6949);
nand U14972 (N_14972,N_7865,N_6747);
nand U14973 (N_14973,N_9399,N_6812);
and U14974 (N_14974,N_8352,N_5367);
and U14975 (N_14975,N_6386,N_6074);
nor U14976 (N_14976,N_5707,N_8614);
or U14977 (N_14977,N_5313,N_6025);
and U14978 (N_14978,N_6867,N_6963);
or U14979 (N_14979,N_8320,N_6382);
nand U14980 (N_14980,N_8947,N_9105);
xnor U14981 (N_14981,N_9623,N_5352);
nor U14982 (N_14982,N_6286,N_7813);
nand U14983 (N_14983,N_5391,N_7889);
nor U14984 (N_14984,N_6636,N_6128);
or U14985 (N_14985,N_7156,N_7559);
nand U14986 (N_14986,N_8020,N_7843);
or U14987 (N_14987,N_6832,N_6178);
nor U14988 (N_14988,N_9776,N_6852);
and U14989 (N_14989,N_6488,N_7839);
and U14990 (N_14990,N_8141,N_7158);
nand U14991 (N_14991,N_8912,N_6523);
or U14992 (N_14992,N_5654,N_9807);
or U14993 (N_14993,N_9150,N_6037);
nor U14994 (N_14994,N_8296,N_5779);
and U14995 (N_14995,N_8374,N_7001);
nor U14996 (N_14996,N_6565,N_5978);
and U14997 (N_14997,N_9243,N_9232);
and U14998 (N_14998,N_6124,N_5991);
nand U14999 (N_14999,N_5074,N_8826);
or UO_0 (O_0,N_12062,N_12675);
and UO_1 (O_1,N_12580,N_13707);
nand UO_2 (O_2,N_10078,N_13142);
or UO_3 (O_3,N_14389,N_14000);
nand UO_4 (O_4,N_13663,N_10686);
nor UO_5 (O_5,N_12228,N_14772);
or UO_6 (O_6,N_11323,N_12567);
or UO_7 (O_7,N_11798,N_14562);
nor UO_8 (O_8,N_14537,N_12769);
or UO_9 (O_9,N_13060,N_13686);
nand UO_10 (O_10,N_14311,N_11359);
and UO_11 (O_11,N_11848,N_11578);
nor UO_12 (O_12,N_10883,N_11194);
or UO_13 (O_13,N_14785,N_13376);
nand UO_14 (O_14,N_13559,N_12929);
or UO_15 (O_15,N_12378,N_13496);
nor UO_16 (O_16,N_11602,N_12527);
and UO_17 (O_17,N_13722,N_11763);
nor UO_18 (O_18,N_13108,N_10316);
and UO_19 (O_19,N_14868,N_11852);
or UO_20 (O_20,N_13678,N_13979);
and UO_21 (O_21,N_10393,N_14298);
nor UO_22 (O_22,N_10977,N_12725);
or UO_23 (O_23,N_11722,N_12290);
nand UO_24 (O_24,N_11742,N_13049);
nand UO_25 (O_25,N_13879,N_11011);
nand UO_26 (O_26,N_14894,N_13569);
nand UO_27 (O_27,N_13876,N_12362);
nor UO_28 (O_28,N_11978,N_13860);
nand UO_29 (O_29,N_11054,N_13459);
and UO_30 (O_30,N_14190,N_12348);
and UO_31 (O_31,N_10057,N_10612);
nand UO_32 (O_32,N_12177,N_10813);
or UO_33 (O_33,N_12860,N_13038);
nand UO_34 (O_34,N_14099,N_10875);
nand UO_35 (O_35,N_14519,N_12958);
nor UO_36 (O_36,N_12332,N_10403);
xnor UO_37 (O_37,N_14585,N_14020);
nor UO_38 (O_38,N_11467,N_12501);
nor UO_39 (O_39,N_13961,N_14352);
and UO_40 (O_40,N_11098,N_14712);
and UO_41 (O_41,N_10930,N_13824);
nand UO_42 (O_42,N_14953,N_12208);
or UO_43 (O_43,N_12068,N_11179);
nor UO_44 (O_44,N_11477,N_13487);
and UO_45 (O_45,N_11986,N_11571);
xnor UO_46 (O_46,N_12306,N_12678);
nand UO_47 (O_47,N_12706,N_13936);
or UO_48 (O_48,N_10553,N_10913);
nand UO_49 (O_49,N_13866,N_13861);
and UO_50 (O_50,N_12593,N_13998);
or UO_51 (O_51,N_13129,N_10855);
nor UO_52 (O_52,N_14941,N_10742);
or UO_53 (O_53,N_14991,N_14720);
or UO_54 (O_54,N_11086,N_11391);
nor UO_55 (O_55,N_13454,N_13957);
nor UO_56 (O_56,N_10796,N_11002);
and UO_57 (O_57,N_10200,N_13162);
and UO_58 (O_58,N_13660,N_13934);
nand UO_59 (O_59,N_11093,N_13863);
or UO_60 (O_60,N_14815,N_12537);
nand UO_61 (O_61,N_13031,N_12701);
nor UO_62 (O_62,N_11137,N_13478);
or UO_63 (O_63,N_11583,N_13558);
or UO_64 (O_64,N_14653,N_10334);
nor UO_65 (O_65,N_13667,N_12690);
or UO_66 (O_66,N_10529,N_11048);
nand UO_67 (O_67,N_14314,N_10059);
nand UO_68 (O_68,N_13089,N_13619);
nor UO_69 (O_69,N_10801,N_10389);
nor UO_70 (O_70,N_10889,N_10185);
and UO_71 (O_71,N_10784,N_11218);
nor UO_72 (O_72,N_13610,N_14501);
nor UO_73 (O_73,N_10237,N_10023);
or UO_74 (O_74,N_12698,N_12130);
nor UO_75 (O_75,N_12455,N_11659);
xor UO_76 (O_76,N_10512,N_11257);
and UO_77 (O_77,N_12960,N_14694);
nand UO_78 (O_78,N_11961,N_14767);
nor UO_79 (O_79,N_11595,N_10296);
nor UO_80 (O_80,N_12664,N_14691);
or UO_81 (O_81,N_10325,N_10862);
or UO_82 (O_82,N_10670,N_14982);
nor UO_83 (O_83,N_12521,N_10251);
or UO_84 (O_84,N_12493,N_12728);
and UO_85 (O_85,N_12187,N_13229);
and UO_86 (O_86,N_14122,N_10597);
nand UO_87 (O_87,N_14187,N_11376);
and UO_88 (O_88,N_13111,N_12019);
or UO_89 (O_89,N_11454,N_11187);
and UO_90 (O_90,N_14259,N_14820);
or UO_91 (O_91,N_13074,N_10835);
nand UO_92 (O_92,N_11030,N_12717);
and UO_93 (O_93,N_12536,N_12927);
nand UO_94 (O_94,N_13139,N_13580);
nor UO_95 (O_95,N_12380,N_12859);
nand UO_96 (O_96,N_12121,N_13757);
or UO_97 (O_97,N_12823,N_14214);
and UO_98 (O_98,N_10111,N_11959);
nor UO_99 (O_99,N_14273,N_14877);
and UO_100 (O_100,N_11948,N_12325);
and UO_101 (O_101,N_13147,N_10439);
nor UO_102 (O_102,N_10162,N_13041);
nor UO_103 (O_103,N_13105,N_13165);
nor UO_104 (O_104,N_10431,N_14531);
and UO_105 (O_105,N_12096,N_10510);
xor UO_106 (O_106,N_11943,N_11801);
nor UO_107 (O_107,N_11672,N_10839);
and UO_108 (O_108,N_14594,N_11819);
or UO_109 (O_109,N_12040,N_14771);
xnor UO_110 (O_110,N_12110,N_10225);
nand UO_111 (O_111,N_11079,N_10030);
nand UO_112 (O_112,N_10506,N_11408);
or UO_113 (O_113,N_10948,N_11553);
or UO_114 (O_114,N_13000,N_12076);
and UO_115 (O_115,N_11208,N_10705);
nor UO_116 (O_116,N_11534,N_11777);
nand UO_117 (O_117,N_10206,N_14398);
and UO_118 (O_118,N_11291,N_12108);
nand UO_119 (O_119,N_12349,N_12555);
nor UO_120 (O_120,N_11250,N_14500);
nand UO_121 (O_121,N_11930,N_12300);
nand UO_122 (O_122,N_12477,N_11582);
nor UO_123 (O_123,N_12663,N_14764);
nand UO_124 (O_124,N_11138,N_13069);
nand UO_125 (O_125,N_12895,N_12146);
nand UO_126 (O_126,N_12532,N_10548);
nor UO_127 (O_127,N_13134,N_11658);
nor UO_128 (O_128,N_12674,N_10854);
and UO_129 (O_129,N_10327,N_14832);
nand UO_130 (O_130,N_10747,N_11305);
nand UO_131 (O_131,N_11004,N_10125);
nor UO_132 (O_132,N_10236,N_11800);
or UO_133 (O_133,N_12141,N_13898);
or UO_134 (O_134,N_14174,N_14053);
and UO_135 (O_135,N_11234,N_11214);
and UO_136 (O_136,N_12643,N_13398);
nand UO_137 (O_137,N_12506,N_13034);
nor UO_138 (O_138,N_12703,N_12077);
nand UO_139 (O_139,N_11189,N_13633);
and UO_140 (O_140,N_11220,N_13245);
or UO_141 (O_141,N_11872,N_13065);
or UO_142 (O_142,N_13665,N_13532);
nor UO_143 (O_143,N_13115,N_12894);
nand UO_144 (O_144,N_12844,N_11279);
or UO_145 (O_145,N_10034,N_12743);
nor UO_146 (O_146,N_12058,N_12343);
and UO_147 (O_147,N_12112,N_12685);
or UO_148 (O_148,N_12803,N_10219);
and UO_149 (O_149,N_10460,N_14262);
nor UO_150 (O_150,N_11378,N_14490);
or UO_151 (O_151,N_12227,N_12791);
nor UO_152 (O_152,N_14672,N_10526);
nor UO_153 (O_153,N_10521,N_10272);
and UO_154 (O_154,N_14400,N_13916);
or UO_155 (O_155,N_14544,N_13571);
or UO_156 (O_156,N_12519,N_14054);
nand UO_157 (O_157,N_10935,N_11780);
nor UO_158 (O_158,N_12095,N_13611);
nand UO_159 (O_159,N_12600,N_12607);
nor UO_160 (O_160,N_12249,N_14950);
or UO_161 (O_161,N_13716,N_14924);
nor UO_162 (O_162,N_11788,N_10886);
nor UO_163 (O_163,N_10522,N_11841);
nor UO_164 (O_164,N_10701,N_11090);
and UO_165 (O_165,N_12930,N_11834);
nor UO_166 (O_166,N_12118,N_12716);
nor UO_167 (O_167,N_10322,N_10260);
nor UO_168 (O_168,N_12353,N_11874);
nor UO_169 (O_169,N_10519,N_13360);
nand UO_170 (O_170,N_11976,N_10430);
nand UO_171 (O_171,N_10899,N_12129);
or UO_172 (O_172,N_13645,N_12721);
nand UO_173 (O_173,N_13107,N_12396);
nand UO_174 (O_174,N_10517,N_14883);
nand UO_175 (O_175,N_11355,N_11124);
or UO_176 (O_176,N_10075,N_14116);
nor UO_177 (O_177,N_14486,N_11406);
nor UO_178 (O_178,N_12280,N_14529);
and UO_179 (O_179,N_13601,N_10861);
xor UO_180 (O_180,N_14592,N_11810);
nor UO_181 (O_181,N_10991,N_13359);
nor UO_182 (O_182,N_10653,N_11514);
nor UO_183 (O_183,N_12407,N_13675);
and UO_184 (O_184,N_14721,N_11740);
and UO_185 (O_185,N_13029,N_10035);
or UO_186 (O_186,N_13171,N_13567);
or UO_187 (O_187,N_14287,N_12013);
nand UO_188 (O_188,N_14575,N_12990);
nor UO_189 (O_189,N_10698,N_11678);
or UO_190 (O_190,N_13948,N_11744);
and UO_191 (O_191,N_10604,N_10966);
nand UO_192 (O_192,N_12870,N_14405);
nor UO_193 (O_193,N_13662,N_14475);
and UO_194 (O_194,N_14180,N_11980);
and UO_195 (O_195,N_11850,N_11833);
nor UO_196 (O_196,N_10319,N_10908);
and UO_197 (O_197,N_14569,N_13319);
nor UO_198 (O_198,N_13833,N_14106);
or UO_199 (O_199,N_10472,N_13157);
nor UO_200 (O_200,N_14062,N_12213);
or UO_201 (O_201,N_11960,N_13320);
nand UO_202 (O_202,N_10787,N_10235);
or UO_203 (O_203,N_13560,N_12831);
or UO_204 (O_204,N_11073,N_10655);
nor UO_205 (O_205,N_12901,N_10351);
nor UO_206 (O_206,N_11492,N_10484);
or UO_207 (O_207,N_10199,N_12951);
nand UO_208 (O_208,N_12271,N_10253);
or UO_209 (O_209,N_11877,N_14257);
or UO_210 (O_210,N_11771,N_12638);
nand UO_211 (O_211,N_14075,N_13076);
and UO_212 (O_212,N_10543,N_11701);
or UO_213 (O_213,N_14320,N_12671);
nor UO_214 (O_214,N_11593,N_10275);
and UO_215 (O_215,N_13043,N_10143);
nor UO_216 (O_216,N_11115,N_10195);
nor UO_217 (O_217,N_10458,N_13081);
and UO_218 (O_218,N_10903,N_10302);
and UO_219 (O_219,N_14948,N_11643);
or UO_220 (O_220,N_13316,N_11863);
nor UO_221 (O_221,N_12762,N_13014);
and UO_222 (O_222,N_14464,N_10964);
nand UO_223 (O_223,N_10853,N_10064);
or UO_224 (O_224,N_11023,N_12683);
or UO_225 (O_225,N_14893,N_11066);
nand UO_226 (O_226,N_11989,N_10647);
and UO_227 (O_227,N_12773,N_11828);
nand UO_228 (O_228,N_10763,N_14458);
nor UO_229 (O_229,N_13905,N_10640);
or UO_230 (O_230,N_12765,N_12749);
and UO_231 (O_231,N_10626,N_14730);
and UO_232 (O_232,N_11627,N_14252);
nand UO_233 (O_233,N_14325,N_12155);
nand UO_234 (O_234,N_11018,N_10583);
or UO_235 (O_235,N_10246,N_13199);
nand UO_236 (O_236,N_13278,N_10786);
and UO_237 (O_237,N_13419,N_11576);
or UO_238 (O_238,N_12194,N_11116);
nand UO_239 (O_239,N_11560,N_12047);
nor UO_240 (O_240,N_11441,N_11803);
or UO_241 (O_241,N_13392,N_14925);
nor UO_242 (O_242,N_13651,N_12809);
or UO_243 (O_243,N_12970,N_14013);
and UO_244 (O_244,N_11427,N_14150);
xnor UO_245 (O_245,N_14690,N_12439);
nand UO_246 (O_246,N_11373,N_12885);
and UO_247 (O_247,N_13061,N_12474);
nor UO_248 (O_248,N_10304,N_14047);
nand UO_249 (O_249,N_14682,N_14175);
or UO_250 (O_250,N_13701,N_14976);
nand UO_251 (O_251,N_10121,N_10815);
nand UO_252 (O_252,N_13436,N_11062);
nor UO_253 (O_253,N_12036,N_14418);
or UO_254 (O_254,N_13052,N_14789);
nand UO_255 (O_255,N_12203,N_11166);
nor UO_256 (O_256,N_14084,N_12356);
nor UO_257 (O_257,N_12879,N_10369);
and UO_258 (O_258,N_11420,N_11759);
and UO_259 (O_259,N_10523,N_14623);
nor UO_260 (O_260,N_14113,N_10000);
and UO_261 (O_261,N_13037,N_12258);
or UO_262 (O_262,N_14797,N_12511);
xor UO_263 (O_263,N_13179,N_12756);
nor UO_264 (O_264,N_10825,N_12999);
and UO_265 (O_265,N_10391,N_14829);
and UO_266 (O_266,N_13967,N_13112);
or UO_267 (O_267,N_10006,N_12936);
nand UO_268 (O_268,N_11846,N_12975);
nand UO_269 (O_269,N_13057,N_10539);
nand UO_270 (O_270,N_10213,N_13427);
nand UO_271 (O_271,N_12286,N_14747);
or UO_272 (O_272,N_14571,N_12405);
nand UO_273 (O_273,N_12085,N_14104);
and UO_274 (O_274,N_12515,N_13850);
nand UO_275 (O_275,N_14345,N_14394);
and UO_276 (O_276,N_12351,N_10821);
or UO_277 (O_277,N_10153,N_11912);
nand UO_278 (O_278,N_10996,N_14775);
or UO_279 (O_279,N_11704,N_10637);
or UO_280 (O_280,N_10271,N_10455);
or UO_281 (O_281,N_12360,N_12029);
nor UO_282 (O_282,N_12738,N_11077);
and UO_283 (O_283,N_12425,N_10489);
and UO_284 (O_284,N_10036,N_11388);
nor UO_285 (O_285,N_14455,N_14461);
or UO_286 (O_286,N_11142,N_10803);
nor UO_287 (O_287,N_10680,N_14908);
or UO_288 (O_288,N_12814,N_12588);
nand UO_289 (O_289,N_11774,N_12434);
nor UO_290 (O_290,N_14279,N_11878);
and UO_291 (O_291,N_14387,N_11049);
nand UO_292 (O_292,N_11539,N_13235);
nor UO_293 (O_293,N_10792,N_11550);
or UO_294 (O_294,N_11606,N_13561);
or UO_295 (O_295,N_13881,N_10367);
and UO_296 (O_296,N_13289,N_12628);
and UO_297 (O_297,N_14324,N_14293);
or UO_298 (O_298,N_10690,N_11156);
and UO_299 (O_299,N_14192,N_14119);
or UO_300 (O_300,N_11773,N_13303);
or UO_301 (O_301,N_10602,N_10761);
nor UO_302 (O_302,N_11110,N_14007);
nor UO_303 (O_303,N_11059,N_12123);
and UO_304 (O_304,N_11304,N_12090);
nand UO_305 (O_305,N_12750,N_12981);
or UO_306 (O_306,N_12763,N_12817);
and UO_307 (O_307,N_10221,N_14796);
nor UO_308 (O_308,N_13789,N_10073);
nand UO_309 (O_309,N_10353,N_13992);
nor UO_310 (O_310,N_14244,N_13902);
and UO_311 (O_311,N_11526,N_13167);
or UO_312 (O_312,N_11442,N_12946);
or UO_313 (O_313,N_14100,N_12782);
or UO_314 (O_314,N_12541,N_14044);
or UO_315 (O_315,N_11171,N_13379);
nor UO_316 (O_316,N_12565,N_12948);
nor UO_317 (O_317,N_14163,N_14766);
or UO_318 (O_318,N_11232,N_13746);
or UO_319 (O_319,N_12882,N_14364);
or UO_320 (O_320,N_13097,N_10530);
or UO_321 (O_321,N_10429,N_14810);
nor UO_322 (O_322,N_12533,N_11368);
or UO_323 (O_323,N_10440,N_14867);
nor UO_324 (O_324,N_11006,N_12702);
and UO_325 (O_325,N_13770,N_12522);
nand UO_326 (O_326,N_10926,N_10807);
and UO_327 (O_327,N_14277,N_11724);
nor UO_328 (O_328,N_12315,N_12498);
and UO_329 (O_329,N_13779,N_11012);
or UO_330 (O_330,N_12551,N_11473);
nand UO_331 (O_331,N_11775,N_13737);
and UO_332 (O_332,N_11134,N_12884);
xnor UO_333 (O_333,N_10773,N_12347);
or UO_334 (O_334,N_11809,N_10119);
nor UO_335 (O_335,N_12014,N_14805);
and UO_336 (O_336,N_10971,N_10380);
nor UO_337 (O_337,N_11231,N_13166);
nand UO_338 (O_338,N_12967,N_11510);
nand UO_339 (O_339,N_13960,N_11294);
nor UO_340 (O_340,N_10900,N_12982);
or UO_341 (O_341,N_12239,N_12435);
nand UO_342 (O_342,N_10973,N_10846);
and UO_343 (O_343,N_10285,N_12668);
and UO_344 (O_344,N_11590,N_14663);
nor UO_345 (O_345,N_10041,N_14998);
nor UO_346 (O_346,N_13718,N_10762);
nand UO_347 (O_347,N_13855,N_14338);
or UO_348 (O_348,N_12684,N_10731);
nand UO_349 (O_349,N_13756,N_11450);
and UO_350 (O_350,N_11047,N_12785);
xor UO_351 (O_351,N_11383,N_10751);
and UO_352 (O_352,N_13145,N_11080);
and UO_353 (O_353,N_10912,N_11897);
nand UO_354 (O_354,N_13579,N_10595);
nor UO_355 (O_355,N_13835,N_12262);
xor UO_356 (O_356,N_13202,N_14322);
and UO_357 (O_357,N_12826,N_13385);
and UO_358 (O_358,N_12924,N_14994);
or UO_359 (O_359,N_12216,N_12714);
nand UO_360 (O_360,N_14093,N_11888);
or UO_361 (O_361,N_10291,N_13591);
nand UO_362 (O_362,N_11240,N_12616);
nor UO_363 (O_363,N_12662,N_13915);
nor UO_364 (O_364,N_14429,N_10168);
or UO_365 (O_365,N_14807,N_11288);
or UO_366 (O_366,N_14708,N_12388);
and UO_367 (O_367,N_13821,N_13406);
or UO_368 (O_368,N_10062,N_14851);
nand UO_369 (O_369,N_11917,N_13699);
and UO_370 (O_370,N_10453,N_11899);
nor UO_371 (O_371,N_13382,N_12497);
nand UO_372 (O_372,N_14511,N_13920);
nand UO_373 (O_373,N_11682,N_12590);
and UO_374 (O_374,N_11745,N_12056);
nor UO_375 (O_375,N_10120,N_12255);
nor UO_376 (O_376,N_10661,N_10082);
nand UO_377 (O_377,N_10939,N_11866);
nor UO_378 (O_378,N_13613,N_14441);
and UO_379 (O_379,N_11919,N_12151);
or UO_380 (O_380,N_11462,N_13576);
nand UO_381 (O_381,N_13918,N_13148);
or UO_382 (O_382,N_14679,N_14401);
nor UO_383 (O_383,N_11463,N_12428);
nor UO_384 (O_384,N_11347,N_13437);
nand UO_385 (O_385,N_12552,N_12968);
and UO_386 (O_386,N_14977,N_14614);
nand UO_387 (O_387,N_14152,N_13570);
nor UO_388 (O_388,N_11579,N_10451);
and UO_389 (O_389,N_12733,N_10220);
nor UO_390 (O_390,N_11100,N_14457);
and UO_391 (O_391,N_12935,N_14929);
or UO_392 (O_392,N_13449,N_10828);
and UO_393 (O_393,N_12272,N_11739);
nor UO_394 (O_394,N_10280,N_13538);
nand UO_395 (O_395,N_14560,N_10704);
or UO_396 (O_396,N_13354,N_11924);
nor UO_397 (O_397,N_12694,N_10668);
nor UO_398 (O_398,N_10658,N_14258);
nand UO_399 (O_399,N_10159,N_13362);
or UO_400 (O_400,N_11530,N_14156);
nand UO_401 (O_401,N_11836,N_13183);
and UO_402 (O_402,N_11776,N_12713);
nand UO_403 (O_403,N_13630,N_13128);
or UO_404 (O_404,N_14012,N_13480);
nor UO_405 (O_405,N_10051,N_12372);
nor UO_406 (O_406,N_13552,N_14208);
or UO_407 (O_407,N_12807,N_10993);
nand UO_408 (O_408,N_14472,N_11000);
nand UO_409 (O_409,N_11723,N_11071);
and UO_410 (O_410,N_13073,N_11675);
nor UO_411 (O_411,N_11423,N_13338);
or UO_412 (O_412,N_11909,N_13305);
or UO_413 (O_413,N_12363,N_11648);
and UO_414 (O_414,N_12350,N_14024);
or UO_415 (O_415,N_10043,N_13268);
and UO_416 (O_416,N_12313,N_11594);
nand UO_417 (O_417,N_14067,N_13227);
nor UO_418 (O_418,N_12839,N_11538);
nor UO_419 (O_419,N_13837,N_13805);
nor UO_420 (O_420,N_12767,N_10068);
and UO_421 (O_421,N_14478,N_11354);
nand UO_422 (O_422,N_14973,N_13758);
or UO_423 (O_423,N_10020,N_13854);
or UO_424 (O_424,N_14294,N_10083);
nor UO_425 (O_425,N_11668,N_10734);
nand UO_426 (O_426,N_10707,N_13614);
and UO_427 (O_427,N_14154,N_12902);
xor UO_428 (O_428,N_12178,N_13287);
or UO_429 (O_429,N_13340,N_10033);
nor UO_430 (O_430,N_10017,N_10824);
and UO_431 (O_431,N_12140,N_12632);
or UO_432 (O_432,N_10011,N_10675);
or UO_433 (O_433,N_14792,N_14048);
and UO_434 (O_434,N_14406,N_11544);
nor UO_435 (O_435,N_11033,N_12147);
nor UO_436 (O_436,N_12505,N_10699);
nor UO_437 (O_437,N_10953,N_14479);
nor UO_438 (O_438,N_12007,N_14011);
nand UO_439 (O_439,N_14915,N_13130);
and UO_440 (O_440,N_14315,N_11591);
and UO_441 (O_441,N_10131,N_11645);
or UO_442 (O_442,N_14285,N_13365);
nand UO_443 (O_443,N_12206,N_13350);
and UO_444 (O_444,N_13712,N_14817);
nand UO_445 (O_445,N_13592,N_11401);
nor UO_446 (O_446,N_12209,N_14701);
and UO_447 (O_447,N_12812,N_10492);
nor UO_448 (O_448,N_11573,N_11128);
and UO_449 (O_449,N_12611,N_10077);
or UO_450 (O_450,N_10646,N_13429);
or UO_451 (O_451,N_14802,N_11349);
nand UO_452 (O_452,N_10001,N_11718);
xor UO_453 (O_453,N_12319,N_14917);
and UO_454 (O_454,N_10290,N_14539);
nand UO_455 (O_455,N_12352,N_13288);
nand UO_456 (O_456,N_13104,N_12482);
nand UO_457 (O_457,N_14193,N_12955);
and UO_458 (O_458,N_10216,N_14625);
nor UO_459 (O_459,N_14755,N_14370);
nand UO_460 (O_460,N_11731,N_14462);
nor UO_461 (O_461,N_13023,N_12789);
and UO_462 (O_462,N_10002,N_14911);
nand UO_463 (O_463,N_14266,N_14290);
and UO_464 (O_464,N_13814,N_14002);
or UO_465 (O_465,N_10138,N_13596);
or UO_466 (O_466,N_12289,N_14229);
or UO_467 (O_467,N_12584,N_14360);
nor UO_468 (O_468,N_10021,N_12656);
nor UO_469 (O_469,N_14159,N_11239);
or UO_470 (O_470,N_11927,N_10738);
nor UO_471 (O_471,N_14886,N_10288);
xnor UO_472 (O_472,N_10072,N_12641);
nand UO_473 (O_473,N_10404,N_13432);
and UO_474 (O_474,N_10269,N_14882);
and UO_475 (O_475,N_11178,N_12026);
or UO_476 (O_476,N_13045,N_14222);
and UO_477 (O_477,N_14497,N_14255);
and UO_478 (O_478,N_12292,N_12075);
or UO_479 (O_479,N_11436,N_14281);
nand UO_480 (O_480,N_13566,N_13414);
xor UO_481 (O_481,N_13472,N_11265);
nor UO_482 (O_482,N_10249,N_10388);
and UO_483 (O_483,N_14449,N_10481);
and UO_484 (O_484,N_11200,N_12296);
or UO_485 (O_485,N_13426,N_12275);
nor UO_486 (O_486,N_14652,N_10584);
or UO_487 (O_487,N_12461,N_13627);
or UO_488 (O_488,N_14932,N_12169);
and UO_489 (O_489,N_11044,N_13378);
and UO_490 (O_490,N_12504,N_12467);
and UO_491 (O_491,N_13363,N_11529);
nor UO_492 (O_492,N_14719,N_14634);
or UO_493 (O_493,N_10897,N_13731);
or UO_494 (O_494,N_11936,N_11461);
nor UO_495 (O_495,N_13710,N_11599);
nand UO_496 (O_496,N_12950,N_11998);
and UO_497 (O_497,N_14332,N_12693);
nor UO_498 (O_498,N_14538,N_14507);
nor UO_499 (O_499,N_13190,N_11015);
nand UO_500 (O_500,N_14938,N_11301);
or UO_501 (O_501,N_14648,N_13116);
and UO_502 (O_502,N_14627,N_11716);
nand UO_503 (O_503,N_13846,N_10619);
nor UO_504 (O_504,N_10924,N_11966);
and UO_505 (O_505,N_11702,N_13394);
nor UO_506 (O_506,N_13612,N_10187);
nor UO_507 (O_507,N_10445,N_14516);
nor UO_508 (O_508,N_10884,N_13536);
and UO_509 (O_509,N_11482,N_12354);
nand UO_510 (O_510,N_12205,N_12840);
and UO_511 (O_511,N_13025,N_11146);
nand UO_512 (O_512,N_10838,N_12137);
nand UO_513 (O_513,N_12862,N_12198);
or UO_514 (O_514,N_14657,N_13222);
nand UO_515 (O_515,N_13251,N_12687);
nand UO_516 (O_516,N_14182,N_10139);
nor UO_517 (O_517,N_11026,N_12727);
and UO_518 (O_518,N_11922,N_14198);
and UO_519 (O_519,N_12181,N_13384);
nand UO_520 (O_520,N_12775,N_14931);
xnor UO_521 (O_521,N_12881,N_11620);
nand UO_522 (O_522,N_10877,N_14871);
nor UO_523 (O_523,N_14862,N_12442);
nor UO_524 (O_524,N_10631,N_12875);
nor UO_525 (O_525,N_12135,N_14814);
or UO_526 (O_526,N_12192,N_12126);
nand UO_527 (O_527,N_12916,N_11198);
or UO_528 (O_528,N_13815,N_14160);
nor UO_529 (O_529,N_13012,N_12375);
nor UO_530 (O_530,N_14573,N_14142);
nand UO_531 (O_531,N_13064,N_10244);
and UO_532 (O_532,N_13329,N_13258);
nor UO_533 (O_533,N_13704,N_10149);
and UO_534 (O_534,N_14246,N_10665);
or UO_535 (O_535,N_14390,N_10684);
nand UO_536 (O_536,N_14356,N_14803);
nand UO_537 (O_537,N_12111,N_10402);
or UO_538 (O_538,N_14469,N_12778);
or UO_539 (O_539,N_12734,N_12972);
or UO_540 (O_540,N_14746,N_13267);
nor UO_541 (O_541,N_14468,N_11915);
and UO_542 (O_542,N_14280,N_14778);
nand UO_543 (O_543,N_11548,N_11107);
and UO_544 (O_544,N_10040,N_12898);
xor UO_545 (O_545,N_12806,N_13264);
xnor UO_546 (O_546,N_11638,N_12270);
or UO_547 (O_547,N_12087,N_12230);
nor UO_548 (O_548,N_13033,N_10140);
nor UO_549 (O_549,N_11857,N_14460);
xnor UO_550 (O_550,N_14812,N_12283);
nand UO_551 (O_551,N_12923,N_10486);
and UO_552 (O_552,N_12175,N_14631);
and UO_553 (O_553,N_13706,N_14819);
and UO_554 (O_554,N_13729,N_14179);
nand UO_555 (O_555,N_13892,N_13927);
nand UO_556 (O_556,N_14849,N_10625);
nor UO_557 (O_557,N_10574,N_12779);
nand UO_558 (O_558,N_12486,N_14340);
or UO_559 (O_559,N_13401,N_11710);
and UO_560 (O_560,N_10891,N_13456);
nor UO_561 (O_561,N_12285,N_11206);
or UO_562 (O_562,N_13823,N_11904);
and UO_563 (O_563,N_14234,N_14848);
or UO_564 (O_564,N_14822,N_11882);
nor UO_565 (O_565,N_13302,N_14649);
nand UO_566 (O_566,N_14008,N_12652);
nand UO_567 (O_567,N_13926,N_10907);
nand UO_568 (O_568,N_13945,N_11812);
nand UO_569 (O_569,N_10344,N_11060);
nor UO_570 (O_570,N_14874,N_12499);
nor UO_571 (O_571,N_12869,N_13700);
nor UO_572 (O_572,N_11438,N_11649);
nor UO_573 (O_573,N_14219,N_13556);
or UO_574 (O_574,N_10493,N_10012);
and UO_575 (O_575,N_11133,N_12557);
and UO_576 (O_576,N_11010,N_10049);
or UO_577 (O_577,N_13046,N_11891);
and UO_578 (O_578,N_12842,N_14102);
nor UO_579 (O_579,N_12395,N_14088);
nor UO_580 (O_580,N_10113,N_10268);
or UO_581 (O_581,N_13009,N_13039);
and UO_582 (O_582,N_11422,N_10054);
nor UO_583 (O_583,N_13241,N_13265);
nor UO_584 (O_584,N_10362,N_11807);
nand UO_585 (O_585,N_12947,N_11404);
or UO_586 (O_586,N_14843,N_10536);
and UO_587 (O_587,N_13852,N_11032);
or UO_588 (O_588,N_11719,N_14473);
or UO_589 (O_589,N_13972,N_13239);
nor UO_590 (O_590,N_14547,N_14251);
or UO_591 (O_591,N_12035,N_11937);
xor UO_592 (O_592,N_12954,N_13582);
and UO_593 (O_593,N_14637,N_10921);
or UO_594 (O_594,N_13192,N_11992);
and UO_595 (O_595,N_10231,N_13818);
nand UO_596 (O_596,N_12832,N_14485);
nor UO_597 (O_597,N_13224,N_14518);
or UO_598 (O_598,N_10318,N_10980);
or UO_599 (O_599,N_11019,N_13284);
and UO_600 (O_600,N_14636,N_10433);
and UO_601 (O_601,N_11226,N_14153);
nand UO_602 (O_602,N_10332,N_14147);
nor UO_603 (O_603,N_11511,N_10375);
nor UO_604 (O_604,N_11303,N_10427);
nor UO_605 (O_605,N_10949,N_14853);
nand UO_606 (O_606,N_13572,N_11248);
nand UO_607 (O_607,N_12669,N_12856);
nor UO_608 (O_608,N_14620,N_12295);
or UO_609 (O_609,N_12707,N_10205);
or UO_610 (O_610,N_10385,N_11623);
or UO_611 (O_611,N_11779,N_13887);
and UO_612 (O_612,N_13938,N_11120);
and UO_613 (O_613,N_13759,N_14555);
and UO_614 (O_614,N_10641,N_10176);
or UO_615 (O_615,N_14225,N_14223);
and UO_616 (O_616,N_11508,N_14574);
nor UO_617 (O_617,N_13193,N_14707);
nor UO_618 (O_618,N_11176,N_13313);
nand UO_619 (O_619,N_10016,N_13598);
or UO_620 (O_620,N_11324,N_13607);
nor UO_621 (O_621,N_10416,N_10981);
nor UO_622 (O_622,N_12568,N_12589);
and UO_623 (O_623,N_13356,N_13859);
and UO_624 (O_624,N_11042,N_11916);
and UO_625 (O_625,N_13840,N_12361);
or UO_626 (O_626,N_11244,N_13078);
and UO_627 (O_627,N_13174,N_11319);
xnor UO_628 (O_628,N_10413,N_12978);
nand UO_629 (O_629,N_14014,N_14243);
or UO_630 (O_630,N_12992,N_11657);
nand UO_631 (O_631,N_13557,N_14744);
and UO_632 (O_632,N_13180,N_12531);
or UO_633 (O_633,N_12323,N_14872);
and UO_634 (O_634,N_10273,N_12441);
nor UO_635 (O_635,N_10056,N_10740);
nand UO_636 (O_636,N_10769,N_14336);
and UO_637 (O_637,N_13512,N_11784);
nor UO_638 (O_638,N_11656,N_12850);
nand UO_639 (O_639,N_12489,N_11953);
nand UO_640 (O_640,N_12104,N_13689);
nor UO_641 (O_641,N_10736,N_12411);
nand UO_642 (O_642,N_14845,N_10297);
nor UO_643 (O_643,N_10343,N_11782);
and UO_644 (O_644,N_13191,N_12542);
or UO_645 (O_645,N_10495,N_14289);
and UO_646 (O_646,N_11384,N_12386);
or UO_647 (O_647,N_11387,N_10081);
nor UO_648 (O_648,N_10499,N_12468);
nor UO_649 (O_649,N_10386,N_12265);
xor UO_650 (O_650,N_11425,N_12644);
nor UO_651 (O_651,N_10477,N_11058);
and UO_652 (O_652,N_14535,N_14045);
xor UO_653 (O_653,N_12528,N_13486);
and UO_654 (O_654,N_13608,N_14063);
nand UO_655 (O_655,N_12858,N_12827);
or UO_656 (O_656,N_14546,N_10307);
or UO_657 (O_657,N_11205,N_13732);
and UO_658 (O_658,N_12221,N_11310);
or UO_659 (O_659,N_10487,N_10203);
nor UO_660 (O_660,N_12071,N_11869);
nand UO_661 (O_661,N_14196,N_10848);
nand UO_662 (O_662,N_10259,N_12091);
and UO_663 (O_663,N_11757,N_12890);
and UO_664 (O_664,N_13373,N_13634);
nor UO_665 (O_665,N_10863,N_14041);
and UO_666 (O_666,N_11238,N_14132);
or UO_667 (O_667,N_10960,N_14943);
or UO_668 (O_668,N_12225,N_13931);
or UO_669 (O_669,N_11089,N_10592);
nand UO_670 (O_670,N_13909,N_11847);
and UO_671 (O_671,N_14384,N_11353);
nand UO_672 (O_672,N_12988,N_13606);
nand UO_673 (O_673,N_12677,N_10586);
nand UO_674 (O_674,N_14016,N_10128);
or UO_675 (O_675,N_12755,N_10798);
or UO_676 (O_676,N_12245,N_14856);
nor UO_677 (O_677,N_12376,N_14790);
nand UO_678 (O_678,N_14759,N_12686);
nand UO_679 (O_679,N_12069,N_14705);
and UO_680 (O_680,N_12226,N_12597);
xor UO_681 (O_681,N_13058,N_10958);
and UO_682 (O_682,N_12369,N_12214);
nand UO_683 (O_683,N_12324,N_14580);
nand UO_684 (O_684,N_10141,N_13673);
nor UO_685 (O_685,N_12938,N_14919);
and UO_686 (O_686,N_12861,N_13882);
or UO_687 (O_687,N_13448,N_10759);
or UO_688 (O_688,N_10364,N_14567);
and UO_689 (O_689,N_11219,N_14838);
and UO_690 (O_690,N_11994,N_13997);
or UO_691 (O_691,N_10424,N_11935);
nand UO_692 (O_692,N_11618,N_13590);
or UO_693 (O_693,N_14808,N_14884);
and UO_694 (O_694,N_10755,N_10601);
xnor UO_695 (O_695,N_10587,N_11967);
xor UO_696 (O_696,N_12413,N_10810);
nor UO_697 (O_697,N_11691,N_11228);
or UO_698 (O_698,N_11111,N_12994);
or UO_699 (O_699,N_14835,N_14981);
and UO_700 (O_700,N_10502,N_13355);
and UO_701 (O_701,N_10423,N_11996);
xor UO_702 (O_702,N_13169,N_13597);
and UO_703 (O_703,N_13565,N_12453);
or UO_704 (O_704,N_14167,N_11568);
nor UO_705 (O_705,N_14552,N_11157);
nor UO_706 (O_706,N_11795,N_13098);
nand UO_707 (O_707,N_14956,N_12079);
or UO_708 (O_708,N_12145,N_13669);
nand UO_709 (O_709,N_13826,N_13418);
or UO_710 (O_710,N_14073,N_13528);
or UO_711 (O_711,N_13742,N_14071);
or UO_712 (O_712,N_13540,N_10130);
and UO_713 (O_713,N_12202,N_11022);
nand UO_714 (O_714,N_12538,N_11958);
nand UO_715 (O_715,N_13775,N_13240);
nand UO_716 (O_716,N_14825,N_10158);
or UO_717 (O_717,N_11309,N_11256);
nand UO_718 (O_718,N_14206,N_13019);
nand UO_719 (O_719,N_11112,N_13249);
or UO_720 (O_720,N_10015,N_13734);
nand UO_721 (O_721,N_11284,N_13153);
nor UO_722 (O_722,N_14704,N_13695);
nor UO_723 (O_723,N_12367,N_13642);
and UO_724 (O_724,N_11876,N_10395);
and UO_725 (O_725,N_10505,N_12899);
nor UO_726 (O_726,N_13691,N_10613);
nor UO_727 (O_727,N_13648,N_14015);
or UO_728 (O_728,N_11975,N_10710);
or UO_729 (O_729,N_12815,N_13848);
nor UO_730 (O_730,N_11003,N_11765);
nand UO_731 (O_731,N_12436,N_12480);
and UO_732 (O_732,N_13466,N_13194);
or UO_733 (O_733,N_14031,N_14442);
and UO_734 (O_734,N_12896,N_10117);
nand UO_735 (O_735,N_12193,N_14094);
and UO_736 (O_736,N_11747,N_12308);
or UO_737 (O_737,N_12513,N_12692);
or UO_738 (O_738,N_10181,N_13403);
nand UO_739 (O_739,N_14482,N_11666);
and UO_740 (O_740,N_11148,N_10365);
nand UO_741 (O_741,N_11889,N_12636);
nor UO_742 (O_742,N_10192,N_14227);
or UO_743 (O_743,N_14284,N_14463);
or UO_744 (O_744,N_14365,N_14590);
or UO_745 (O_745,N_10157,N_10412);
nand UO_746 (O_746,N_11950,N_14288);
and UO_747 (O_747,N_11332,N_11946);
nor UO_748 (O_748,N_14250,N_11147);
or UO_749 (O_749,N_11424,N_14568);
nand UO_750 (O_750,N_10994,N_12872);
and UO_751 (O_751,N_14930,N_11905);
and UO_752 (O_752,N_12402,N_13991);
nand UO_753 (O_753,N_13286,N_12392);
or UO_754 (O_754,N_13799,N_14906);
nor UO_755 (O_755,N_14698,N_12530);
and UO_756 (O_756,N_11270,N_13637);
nor UO_757 (O_757,N_12165,N_13721);
or UO_758 (O_758,N_12222,N_13537);
or UO_759 (O_759,N_13136,N_13450);
nor UO_760 (O_760,N_12065,N_12021);
nor UO_761 (O_761,N_14433,N_10494);
or UO_762 (O_762,N_14139,N_10904);
xor UO_763 (O_763,N_13188,N_11315);
or UO_764 (O_764,N_11637,N_12976);
nand UO_765 (O_765,N_14110,N_14600);
and UO_766 (O_766,N_13773,N_13095);
and UO_767 (O_767,N_11313,N_10882);
nor UO_768 (O_768,N_14992,N_11831);
nor UO_769 (O_769,N_14527,N_10609);
nand UO_770 (O_770,N_13907,N_13423);
and UO_771 (O_771,N_10859,N_14818);
and UO_772 (O_772,N_11293,N_13455);
xnor UO_773 (O_773,N_12987,N_12676);
or UO_774 (O_774,N_10198,N_14654);
and UO_775 (O_775,N_14070,N_12558);
nand UO_776 (O_776,N_13653,N_13274);
nand UO_777 (O_777,N_11736,N_11465);
or UO_778 (O_778,N_12485,N_13836);
nand UO_779 (O_779,N_11460,N_10384);
nor UO_780 (O_780,N_11053,N_14933);
nand UO_781 (O_781,N_10898,N_12424);
xor UO_782 (O_782,N_12092,N_10084);
and UO_783 (O_783,N_14999,N_10337);
or UO_784 (O_784,N_14028,N_11537);
and UO_785 (O_785,N_12556,N_13811);
nor UO_786 (O_786,N_11416,N_10454);
and UO_787 (O_787,N_11290,N_10104);
and UO_788 (O_788,N_10920,N_10474);
or UO_789 (O_789,N_13534,N_11651);
or UO_790 (O_790,N_12100,N_11830);
xor UO_791 (O_791,N_13656,N_13242);
and UO_792 (O_792,N_11518,N_11892);
and UO_793 (O_793,N_10009,N_14009);
xnor UO_794 (O_794,N_11348,N_13523);
nand UO_795 (O_795,N_10032,N_14446);
and UO_796 (O_796,N_14633,N_13505);
nor UO_797 (O_797,N_12579,N_14415);
or UO_798 (O_798,N_13301,N_11340);
or UO_799 (O_799,N_10028,N_11654);
and UO_800 (O_800,N_12876,N_10417);
nand UO_801 (O_801,N_10048,N_12000);
or UO_802 (O_802,N_13400,N_14026);
or UO_803 (O_803,N_13150,N_14795);
and UO_804 (O_804,N_14396,N_12700);
and UO_805 (O_805,N_12131,N_14261);
or UO_806 (O_806,N_13888,N_13422);
nand UO_807 (O_807,N_11644,N_10739);
or UO_808 (O_808,N_10490,N_14328);
nor UO_809 (O_809,N_13482,N_10975);
nor UO_810 (O_810,N_13754,N_12414);
nand UO_811 (O_811,N_13919,N_13932);
nor UO_812 (O_812,N_12409,N_14971);
and UO_813 (O_813,N_12617,N_10676);
and UO_814 (O_814,N_10756,N_11485);
or UO_815 (O_815,N_14051,N_10406);
or UO_816 (O_816,N_10937,N_12710);
nand UO_817 (O_817,N_12002,N_11051);
or UO_818 (O_818,N_12043,N_12122);
nand UO_819 (O_819,N_10473,N_10575);
or UO_820 (O_820,N_14178,N_10713);
nor UO_821 (O_821,N_13255,N_14138);
or UO_822 (O_822,N_10368,N_12563);
and UO_823 (O_823,N_11493,N_14750);
nor UO_824 (O_824,N_10007,N_14632);
nor UO_825 (O_825,N_12843,N_12962);
or UO_826 (O_826,N_10933,N_14944);
nor UO_827 (O_827,N_12423,N_13237);
xnor UO_828 (O_828,N_13168,N_10061);
nor UO_829 (O_829,N_12516,N_14665);
nand UO_830 (O_830,N_14143,N_11161);
and UO_831 (O_831,N_14528,N_14358);
xor UO_832 (O_832,N_13375,N_10067);
nand UO_833 (O_833,N_13966,N_10374);
nand UO_834 (O_834,N_13473,N_12287);
or UO_835 (O_835,N_14865,N_11837);
nor UO_836 (O_836,N_14080,N_10715);
or UO_837 (O_837,N_13172,N_12742);
nand UO_838 (O_838,N_14710,N_13803);
xnor UO_839 (O_839,N_12723,N_10681);
or UO_840 (O_840,N_14004,N_11330);
and UO_841 (O_841,N_11525,N_10256);
and UO_842 (O_842,N_13875,N_11289);
nor UO_843 (O_843,N_11292,N_13315);
or UO_844 (O_844,N_10039,N_13631);
or UO_845 (O_845,N_12925,N_13170);
nor UO_846 (O_846,N_14309,N_12983);
and UO_847 (O_847,N_14351,N_11920);
nand UO_848 (O_848,N_11929,N_14800);
nor UO_849 (O_849,N_10109,N_13304);
nor UO_850 (O_850,N_12645,N_12609);
or UO_851 (O_851,N_13970,N_12373);
and UO_852 (O_852,N_12508,N_13297);
or UO_853 (O_853,N_13318,N_13819);
nand UO_854 (O_854,N_10791,N_14523);
nand UO_855 (O_855,N_14348,N_13272);
nor UO_856 (O_856,N_14635,N_12142);
xnor UO_857 (O_857,N_13083,N_14123);
nand UO_858 (O_858,N_12667,N_10189);
and UO_859 (O_859,N_13709,N_10100);
or UO_860 (O_860,N_10305,N_12573);
and UO_861 (O_861,N_14791,N_14510);
nor UO_862 (O_862,N_14936,N_14437);
or UO_863 (O_863,N_11767,N_10894);
nor UO_864 (O_864,N_14505,N_12136);
nor UO_865 (O_865,N_13953,N_11321);
nor UO_866 (O_866,N_10564,N_12025);
or UO_867 (O_867,N_13283,N_10469);
and UO_868 (O_868,N_12168,N_13390);
or UO_869 (O_869,N_10047,N_10163);
nor UO_870 (O_870,N_13123,N_10397);
nor UO_871 (O_871,N_14591,N_14353);
nor UO_872 (O_872,N_10070,N_13271);
and UO_873 (O_873,N_10618,N_13294);
nor UO_874 (O_874,N_12293,N_13079);
nand UO_875 (O_875,N_12317,N_10396);
or UO_876 (O_876,N_12759,N_10465);
and UO_877 (O_877,N_11346,N_13435);
nand UO_878 (O_878,N_14899,N_13230);
and UO_879 (O_879,N_13453,N_13159);
or UO_880 (O_880,N_13216,N_11150);
or UO_881 (O_881,N_11977,N_12623);
nand UO_882 (O_882,N_11122,N_13420);
nand UO_883 (O_883,N_14570,N_14064);
or UO_884 (O_884,N_12543,N_14183);
or UO_885 (O_885,N_13980,N_13279);
nor UO_886 (O_886,N_12735,N_13573);
and UO_887 (O_887,N_13409,N_14728);
nor UO_888 (O_888,N_10091,N_14079);
nor UO_889 (O_889,N_12039,N_14968);
nand UO_890 (O_890,N_12182,N_14168);
or UO_891 (O_891,N_11862,N_13812);
nand UO_892 (O_892,N_14949,N_11083);
or UO_893 (O_893,N_14629,N_13867);
and UO_894 (O_894,N_13217,N_10540);
and UO_895 (O_895,N_14172,N_12390);
or UO_896 (O_896,N_12236,N_10628);
and UO_897 (O_897,N_12061,N_12417);
nor UO_898 (O_898,N_10025,N_11785);
nor UO_899 (O_899,N_14432,N_10266);
or UO_900 (O_900,N_11433,N_12783);
and UO_901 (O_901,N_14508,N_10408);
nand UO_902 (O_902,N_10910,N_14006);
nand UO_903 (O_903,N_11705,N_14029);
or UO_904 (O_904,N_10151,N_11921);
and UO_905 (O_905,N_13864,N_11569);
nand UO_906 (O_906,N_12626,N_11439);
and UO_907 (O_907,N_11449,N_13088);
xnor UO_908 (O_908,N_13741,N_11532);
nand UO_909 (O_909,N_14566,N_13372);
nand UO_910 (O_910,N_12634,N_12031);
or UO_911 (O_911,N_11715,N_14403);
nand UO_912 (O_912,N_12848,N_12083);
and UO_913 (O_913,N_11409,N_10938);
and UO_914 (O_914,N_11505,N_14256);
nor UO_915 (O_915,N_14558,N_13890);
nor UO_916 (O_916,N_10673,N_12906);
nor UO_917 (O_917,N_11105,N_10532);
or UO_918 (O_918,N_13622,N_14491);
nor UO_919 (O_919,N_14828,N_12926);
xor UO_920 (O_920,N_13795,N_11808);
nand UO_921 (O_921,N_14181,N_10890);
nand UO_922 (O_922,N_11804,N_10136);
or UO_923 (O_923,N_13894,N_11898);
nor UO_924 (O_924,N_10941,N_12445);
or UO_925 (O_925,N_13201,N_10679);
nand UO_926 (O_926,N_11814,N_14644);
nor UO_927 (O_927,N_12625,N_14503);
nand UO_928 (O_928,N_11322,N_13118);
and UO_929 (O_929,N_10954,N_12646);
nand UO_930 (O_930,N_13114,N_13535);
and UO_931 (O_931,N_14001,N_13018);
or UO_932 (O_932,N_10241,N_12475);
nand UO_933 (O_933,N_14303,N_13776);
nand UO_934 (O_934,N_13412,N_10919);
nor UO_935 (O_935,N_11799,N_10116);
nand UO_936 (O_936,N_13431,N_10295);
nor UO_937 (O_937,N_14970,N_10475);
and UO_938 (O_938,N_11481,N_11328);
nor UO_939 (O_939,N_13725,N_14859);
or UO_940 (O_940,N_14669,N_10463);
nor UO_941 (O_941,N_14650,N_13469);
nor UO_942 (O_942,N_11141,N_12189);
nand UO_943 (O_943,N_14864,N_11167);
or UO_944 (O_944,N_12888,N_14608);
nor UO_945 (O_945,N_14380,N_10497);
or UO_946 (O_946,N_10593,N_10620);
nor UO_947 (O_947,N_11393,N_11034);
or UO_948 (O_948,N_12544,N_12223);
or UO_949 (O_949,N_14826,N_13257);
or UO_950 (O_950,N_11750,N_14673);
and UO_951 (O_951,N_13838,N_14329);
nand UO_952 (O_952,N_11426,N_13880);
and UO_953 (O_953,N_13763,N_10720);
or UO_954 (O_954,N_10101,N_12163);
or UO_955 (O_955,N_10265,N_14624);
and UO_956 (O_956,N_10524,N_10527);
nand UO_957 (O_957,N_11683,N_14959);
or UO_958 (O_958,N_11464,N_12382);
and UO_959 (O_959,N_12481,N_14430);
and UO_960 (O_960,N_10278,N_14869);
or UO_961 (O_961,N_12786,N_10303);
nand UO_962 (O_962,N_12073,N_12164);
or UO_963 (O_963,N_10697,N_11679);
xor UO_964 (O_964,N_14382,N_10184);
nor UO_965 (O_965,N_13618,N_12830);
nor UO_966 (O_966,N_12961,N_11448);
and UO_967 (O_967,N_11399,N_14895);
and UO_968 (O_968,N_14763,N_13173);
nor UO_969 (O_969,N_13949,N_13893);
or UO_970 (O_970,N_14907,N_11821);
nand UO_971 (O_971,N_14282,N_12297);
nor UO_972 (O_972,N_11103,N_13369);
nand UO_973 (O_973,N_14202,N_12998);
and UO_974 (O_974,N_10211,N_11084);
and UO_975 (O_975,N_13131,N_11035);
nor UO_976 (O_976,N_13674,N_11275);
nor UO_977 (O_977,N_11727,N_11695);
nor UO_978 (O_978,N_12304,N_10611);
nand UO_979 (O_979,N_13813,N_11398);
nor UO_980 (O_980,N_11224,N_10464);
and UO_981 (O_981,N_11859,N_13541);
and UO_982 (O_982,N_10425,N_11453);
nor UO_983 (O_983,N_13896,N_14873);
nand UO_984 (O_984,N_13308,N_14346);
or UO_985 (O_985,N_13659,N_12866);
or UO_986 (O_986,N_13603,N_10124);
or UO_987 (O_987,N_13467,N_14267);
nor UO_988 (O_988,N_13198,N_12457);
and UO_989 (O_989,N_10382,N_11887);
or UO_990 (O_990,N_10942,N_11811);
nor UO_991 (O_991,N_10079,N_14866);
or UO_992 (O_992,N_12931,N_14909);
nor UO_993 (O_993,N_13782,N_10623);
nor UO_994 (O_994,N_14146,N_10906);
or UO_995 (O_995,N_13650,N_13460);
or UO_996 (O_996,N_10224,N_12871);
nor UO_997 (O_997,N_13891,N_12545);
nor UO_998 (O_998,N_11840,N_10608);
and UO_999 (O_999,N_12891,N_11091);
or UO_1000 (O_1000,N_11016,N_11282);
or UO_1001 (O_1001,N_13261,N_11278);
nor UO_1002 (O_1002,N_13238,N_10421);
or UO_1003 (O_1003,N_12928,N_11577);
or UO_1004 (O_1004,N_14074,N_14927);
or UO_1005 (O_1005,N_10214,N_10190);
or UO_1006 (O_1006,N_14593,N_11225);
or UO_1007 (O_1007,N_13717,N_13696);
and UO_1008 (O_1008,N_12195,N_13899);
and UO_1009 (O_1009,N_14850,N_13632);
or UO_1010 (O_1010,N_13164,N_10832);
nand UO_1011 (O_1011,N_11013,N_14039);
nand UO_1012 (O_1012,N_10180,N_12273);
nand UO_1013 (O_1013,N_12781,N_14077);
or UO_1014 (O_1014,N_10777,N_10446);
nor UO_1015 (O_1015,N_11437,N_12586);
nor UO_1016 (O_1016,N_14582,N_10902);
and UO_1017 (O_1017,N_10970,N_12966);
and UO_1018 (O_1018,N_10851,N_14076);
nor UO_1019 (O_1019,N_10546,N_11109);
or UO_1020 (O_1020,N_13822,N_14421);
and UO_1021 (O_1021,N_13807,N_11570);
nor UO_1022 (O_1022,N_13307,N_12432);
or UO_1023 (O_1023,N_14367,N_13177);
or UO_1024 (O_1024,N_10172,N_13063);
nor UO_1025 (O_1025,N_12012,N_11007);
nand UO_1026 (O_1026,N_12254,N_14022);
and UO_1027 (O_1027,N_12726,N_12200);
nand UO_1028 (O_1028,N_12024,N_14658);
nand UO_1029 (O_1029,N_13889,N_11434);
or UO_1030 (O_1030,N_12996,N_11236);
or UO_1031 (O_1031,N_13113,N_11345);
nor UO_1032 (O_1032,N_11974,N_10161);
nand UO_1033 (O_1033,N_11661,N_11772);
or UO_1034 (O_1034,N_10752,N_13075);
and UO_1035 (O_1035,N_14235,N_11832);
nor UO_1036 (O_1036,N_10757,N_12921);
nor UO_1037 (O_1037,N_12371,N_13862);
or UO_1038 (O_1038,N_10093,N_12965);
or UO_1039 (O_1039,N_13738,N_10836);
nor UO_1040 (O_1040,N_14753,N_14541);
or UO_1041 (O_1041,N_14019,N_10069);
and UO_1042 (O_1042,N_11884,N_10501);
nand UO_1043 (O_1043,N_12795,N_14217);
xor UO_1044 (O_1044,N_12055,N_11366);
nand UO_1045 (O_1045,N_12450,N_14059);
or UO_1046 (O_1046,N_12577,N_13292);
and UO_1047 (O_1047,N_14061,N_12819);
and UO_1048 (O_1048,N_10293,N_14617);
nor UO_1049 (O_1049,N_10459,N_12105);
nor UO_1050 (O_1050,N_13146,N_14655);
and UO_1051 (O_1051,N_11854,N_13072);
and UO_1052 (O_1052,N_12156,N_13600);
or UO_1053 (O_1053,N_10841,N_13253);
nand UO_1054 (O_1054,N_11502,N_11360);
nor UO_1055 (O_1055,N_13697,N_12098);
or UO_1056 (O_1056,N_13908,N_13223);
nor UO_1057 (O_1057,N_10373,N_13093);
or UO_1058 (O_1058,N_14583,N_11910);
and UO_1059 (O_1059,N_10339,N_10286);
and UO_1060 (O_1060,N_12829,N_14049);
nand UO_1061 (O_1061,N_13002,N_12484);
nor UO_1062 (O_1062,N_13080,N_14378);
nand UO_1063 (O_1063,N_10518,N_10652);
and UO_1064 (O_1064,N_11395,N_13186);
nor UO_1065 (O_1065,N_12682,N_11096);
nand UO_1066 (O_1066,N_11165,N_11117);
and UO_1067 (O_1067,N_14327,N_11671);
and UO_1068 (O_1068,N_13548,N_12957);
and UO_1069 (O_1069,N_14203,N_13767);
and UO_1070 (O_1070,N_12082,N_10112);
or UO_1071 (O_1071,N_11758,N_12099);
nor UO_1072 (O_1072,N_10555,N_14656);
or UO_1073 (O_1073,N_14692,N_12610);
nor UO_1074 (O_1074,N_10672,N_13958);
and UO_1075 (O_1075,N_14003,N_10197);
and UO_1076 (O_1076,N_11931,N_11318);
nand UO_1077 (O_1077,N_13625,N_10270);
xnor UO_1078 (O_1078,N_14078,N_14424);
and UO_1079 (O_1079,N_11655,N_11513);
and UO_1080 (O_1080,N_12464,N_13181);
or UO_1081 (O_1081,N_14495,N_14034);
nor UO_1082 (O_1082,N_11585,N_10916);
and UO_1083 (O_1083,N_12771,N_11188);
and UO_1084 (O_1084,N_14718,N_12437);
or UO_1085 (O_1085,N_14955,N_13914);
and UO_1086 (O_1086,N_10805,N_12865);
or UO_1087 (O_1087,N_10276,N_11908);
nor UO_1088 (O_1088,N_14993,N_14777);
or UO_1089 (O_1089,N_11499,N_13066);
or UO_1090 (O_1090,N_12835,N_12010);
nor UO_1091 (O_1091,N_11350,N_11607);
xor UO_1092 (O_1092,N_12219,N_12559);
nand UO_1093 (O_1093,N_11024,N_13739);
nor UO_1094 (O_1094,N_10940,N_11688);
nand UO_1095 (O_1095,N_12758,N_10209);
and UO_1096 (O_1096,N_10410,N_11906);
nor UO_1097 (O_1097,N_10258,N_11069);
or UO_1098 (O_1098,N_14236,N_12134);
or UO_1099 (O_1099,N_11867,N_13396);
and UO_1100 (O_1100,N_13008,N_10554);
nor UO_1101 (O_1101,N_11170,N_11535);
and UO_1102 (O_1102,N_13349,N_13547);
and UO_1103 (O_1103,N_12553,N_13769);
nand UO_1104 (O_1104,N_13522,N_13857);
or UO_1105 (O_1105,N_10551,N_11374);
nor UO_1106 (O_1106,N_12044,N_10842);
nand UO_1107 (O_1107,N_13158,N_12820);
and UO_1108 (O_1108,N_10357,N_11676);
nand UO_1109 (O_1109,N_14794,N_14383);
nor UO_1110 (O_1110,N_12991,N_12132);
or UO_1111 (O_1111,N_14399,N_10360);
or UO_1112 (O_1112,N_13983,N_10053);
nand UO_1113 (O_1113,N_14231,N_10024);
or UO_1114 (O_1114,N_11339,N_13679);
and UO_1115 (O_1115,N_11613,N_13342);
and UO_1116 (O_1116,N_10797,N_11766);
nor UO_1117 (O_1117,N_14983,N_12261);
or UO_1118 (O_1118,N_14465,N_11402);
nand UO_1119 (O_1119,N_11227,N_11370);
and UO_1120 (O_1120,N_12314,N_11476);
nor UO_1121 (O_1121,N_10644,N_12050);
or UO_1122 (O_1122,N_10694,N_12340);
nor UO_1123 (O_1123,N_13277,N_11389);
nor UO_1124 (O_1124,N_10308,N_13969);
or UO_1125 (O_1125,N_13884,N_10106);
nor UO_1126 (O_1126,N_11212,N_13492);
or UO_1127 (O_1127,N_12054,N_13668);
nand UO_1128 (O_1128,N_14688,N_13084);
nor UO_1129 (O_1129,N_12518,N_12447);
or UO_1130 (O_1130,N_12333,N_14450);
nand UO_1131 (O_1131,N_12473,N_12614);
nand UO_1132 (O_1132,N_14823,N_13621);
nand UO_1133 (O_1133,N_11557,N_14010);
nor UO_1134 (O_1134,N_10830,N_10274);
or UO_1135 (O_1135,N_11954,N_12064);
or UO_1136 (O_1136,N_11253,N_14601);
or UO_1137 (O_1137,N_11680,N_12502);
or UO_1138 (O_1138,N_10827,N_11243);
nand UO_1139 (O_1139,N_13051,N_14514);
nor UO_1140 (O_1140,N_14506,N_14752);
nor UO_1141 (O_1141,N_13263,N_14046);
nand UO_1142 (O_1142,N_12576,N_14937);
nand UO_1143 (O_1143,N_12391,N_14599);
and UO_1144 (O_1144,N_12585,N_11515);
nand UO_1145 (O_1145,N_13011,N_12298);
or UO_1146 (O_1146,N_13206,N_12578);
or UO_1147 (O_1147,N_14774,N_10772);
nand UO_1148 (O_1148,N_13551,N_12210);
or UO_1149 (O_1149,N_11043,N_14502);
or UO_1150 (O_1150,N_14935,N_12204);
and UO_1151 (O_1151,N_12051,N_14834);
nand UO_1152 (O_1152,N_11286,N_11713);
and UO_1153 (O_1153,N_12624,N_14498);
and UO_1154 (O_1154,N_14499,N_11222);
or UO_1155 (O_1155,N_13399,N_10401);
or UO_1156 (O_1156,N_11903,N_13588);
nand UO_1157 (O_1157,N_13178,N_10581);
nand UO_1158 (O_1158,N_10799,N_12185);
nor UO_1159 (O_1159,N_14368,N_10857);
nand UO_1160 (O_1160,N_11325,N_14021);
or UO_1161 (O_1161,N_13475,N_12535);
and UO_1162 (O_1162,N_11329,N_11097);
xor UO_1163 (O_1163,N_12596,N_10022);
nor UO_1164 (O_1164,N_14743,N_11181);
nor UO_1165 (O_1165,N_12633,N_12985);
or UO_1166 (O_1166,N_10018,N_13499);
or UO_1167 (O_1167,N_12679,N_13273);
nor UO_1168 (O_1168,N_14946,N_11596);
and UO_1169 (O_1169,N_11755,N_10363);
nand UO_1170 (O_1170,N_11632,N_13831);
nor UO_1171 (O_1171,N_10850,N_12562);
nand UO_1172 (O_1172,N_12910,N_12438);
nand UO_1173 (O_1173,N_11907,N_10549);
xnor UO_1174 (O_1174,N_13021,N_12433);
and UO_1175 (O_1175,N_12940,N_11326);
nand UO_1176 (O_1176,N_14563,N_12242);
or UO_1177 (O_1177,N_13465,N_10664);
nor UO_1178 (O_1178,N_10671,N_13424);
xnor UO_1179 (O_1179,N_13829,N_10345);
nand UO_1180 (O_1180,N_13458,N_10257);
nand UO_1181 (O_1181,N_12517,N_14253);
nand UO_1182 (O_1182,N_13727,N_11229);
or UO_1183 (O_1183,N_11564,N_12801);
or UO_1184 (O_1184,N_13963,N_14268);
or UO_1185 (O_1185,N_12335,N_13550);
nor UO_1186 (O_1186,N_14581,N_13091);
nand UO_1187 (O_1187,N_13110,N_12635);
nand UO_1188 (O_1188,N_10537,N_13203);
nor UO_1189 (O_1189,N_10621,N_10267);
nand UO_1190 (O_1190,N_14169,N_11119);
nand UO_1191 (O_1191,N_14204,N_14536);
or UO_1192 (O_1192,N_13211,N_14852);
nor UO_1193 (O_1193,N_10570,N_10558);
nor UO_1194 (O_1194,N_14436,N_10650);
nor UO_1195 (O_1195,N_13334,N_14840);
nor UO_1196 (O_1196,N_10301,N_12366);
nor UO_1197 (O_1197,N_13138,N_14995);
nand UO_1198 (O_1198,N_10496,N_14855);
nand UO_1199 (O_1199,N_14564,N_10212);
nor UO_1200 (O_1200,N_11660,N_12263);
nor UO_1201 (O_1201,N_11466,N_14709);
nand UO_1202 (O_1202,N_10817,N_13339);
or UO_1203 (O_1203,N_13574,N_14963);
and UO_1204 (O_1204,N_12911,N_12357);
or UO_1205 (O_1205,N_14494,N_13513);
and UO_1206 (O_1206,N_12197,N_10349);
nand UO_1207 (O_1207,N_14717,N_13357);
nor UO_1208 (O_1208,N_12697,N_12281);
and UO_1209 (O_1209,N_14388,N_10052);
or UO_1210 (O_1210,N_12471,N_11459);
or UO_1211 (O_1211,N_13578,N_13903);
nand UO_1212 (O_1212,N_12841,N_13951);
or UO_1213 (O_1213,N_13906,N_12463);
or UO_1214 (O_1214,N_13954,N_12784);
and UO_1215 (O_1215,N_13259,N_10092);
nand UO_1216 (O_1216,N_10097,N_11140);
nor UO_1217 (O_1217,N_12649,N_14184);
nor UO_1218 (O_1218,N_11173,N_10354);
nand UO_1219 (O_1219,N_13748,N_12089);
nor UO_1220 (O_1220,N_11984,N_11639);
and UO_1221 (O_1221,N_13895,N_11403);
or UO_1222 (O_1222,N_13828,N_10038);
or UO_1223 (O_1223,N_11692,N_13868);
and UO_1224 (O_1224,N_10693,N_12640);
nor UO_1225 (O_1225,N_12231,N_10232);
nor UO_1226 (O_1226,N_10448,N_14597);
nand UO_1227 (O_1227,N_12503,N_11087);
nand UO_1228 (O_1228,N_13719,N_11135);
nor UO_1229 (O_1229,N_14619,N_10226);
nand UO_1230 (O_1230,N_13726,N_11700);
or UO_1231 (O_1231,N_10500,N_12084);
and UO_1232 (O_1232,N_14786,N_10515);
nand UO_1233 (O_1233,N_11267,N_10089);
nor UO_1234 (O_1234,N_10013,N_14677);
or UO_1235 (O_1235,N_10833,N_12412);
nand UO_1236 (O_1236,N_12337,N_12969);
nor UO_1237 (O_1237,N_14117,N_14242);
xor UO_1238 (O_1238,N_13816,N_10696);
nand UO_1239 (O_1239,N_12179,N_10164);
and UO_1240 (O_1240,N_14438,N_13276);
or UO_1241 (O_1241,N_11982,N_13511);
nor UO_1242 (O_1242,N_12487,N_13514);
or UO_1243 (O_1243,N_11640,N_10576);
xor UO_1244 (O_1244,N_11995,N_11665);
or UO_1245 (O_1245,N_10310,N_11118);
or UO_1246 (O_1246,N_13521,N_14910);
nor UO_1247 (O_1247,N_11201,N_12460);
and UO_1248 (O_1248,N_14209,N_12162);
or UO_1249 (O_1249,N_12101,N_11753);
nor UO_1250 (O_1250,N_10685,N_10287);
nor UO_1251 (O_1251,N_10802,N_10632);
nand UO_1252 (O_1252,N_13654,N_11129);
or UO_1253 (O_1253,N_11247,N_13161);
nor UO_1254 (O_1254,N_11428,N_13479);
nand UO_1255 (O_1255,N_14120,N_13187);
and UO_1256 (O_1256,N_11802,N_10080);
or UO_1257 (O_1257,N_11746,N_13724);
and UO_1258 (O_1258,N_13506,N_13127);
and UO_1259 (O_1259,N_11806,N_14307);
or UO_1260 (O_1260,N_13768,N_13141);
nor UO_1261 (O_1261,N_10654,N_12629);
and UO_1262 (O_1262,N_10008,N_11997);
nor UO_1263 (O_1263,N_11670,N_14711);
nand UO_1264 (O_1264,N_11709,N_10860);
nor UO_1265 (O_1265,N_12796,N_10758);
or UO_1266 (O_1266,N_11005,N_13441);
nor UO_1267 (O_1267,N_12989,N_14453);
and UO_1268 (O_1268,N_14780,N_13444);
and UO_1269 (O_1269,N_11543,N_10809);
nand UO_1270 (O_1270,N_12346,N_12787);
and UO_1271 (O_1271,N_11856,N_13126);
and UO_1272 (O_1272,N_12491,N_13959);
nor UO_1273 (O_1273,N_10538,N_11895);
nand UO_1274 (O_1274,N_10320,N_12953);
nand UO_1275 (O_1275,N_11099,N_13312);
or UO_1276 (O_1276,N_12605,N_10687);
and UO_1277 (O_1277,N_14130,N_12005);
and UO_1278 (O_1278,N_12158,N_10928);
nand UO_1279 (O_1279,N_14760,N_10315);
nand UO_1280 (O_1280,N_11592,N_13468);
nand UO_1281 (O_1281,N_14740,N_14197);
nor UO_1282 (O_1282,N_13281,N_14896);
and UO_1283 (O_1283,N_13433,N_12846);
nand UO_1284 (O_1284,N_11237,N_13730);
nor UO_1285 (O_1285,N_11956,N_10639);
nor UO_1286 (O_1286,N_11533,N_10003);
and UO_1287 (O_1287,N_10677,N_11299);
nor UO_1288 (O_1288,N_12451,N_12845);
or UO_1289 (O_1289,N_14310,N_10179);
nor UO_1290 (O_1290,N_14683,N_13068);
or UO_1291 (O_1291,N_10255,N_11337);
and UO_1292 (O_1292,N_11475,N_13698);
nand UO_1293 (O_1293,N_10238,N_14647);
and UO_1294 (O_1294,N_14897,N_13986);
nand UO_1295 (O_1295,N_11642,N_14540);
or UO_1296 (O_1296,N_10281,N_10099);
nor UO_1297 (O_1297,N_12148,N_11677);
nor UO_1298 (O_1298,N_12330,N_13575);
and UO_1299 (O_1299,N_13210,N_14550);
or UO_1300 (O_1300,N_13533,N_12627);
or UO_1301 (O_1301,N_14372,N_11407);
nor UO_1302 (O_1302,N_14454,N_12720);
and UO_1303 (O_1303,N_14484,N_14723);
xor UO_1304 (O_1304,N_11687,N_13364);
or UO_1305 (O_1305,N_11586,N_11484);
nand UO_1306 (O_1306,N_14205,N_14604);
or UO_1307 (O_1307,N_10444,N_11818);
nand UO_1308 (O_1308,N_12201,N_12591);
xnor UO_1309 (O_1309,N_12359,N_11581);
or UO_1310 (O_1310,N_12654,N_14108);
and UO_1311 (O_1311,N_10485,N_11754);
or UO_1312 (O_1312,N_14292,N_11913);
or UO_1313 (O_1313,N_11255,N_10559);
and UO_1314 (O_1314,N_13965,N_14549);
or UO_1315 (O_1315,N_10934,N_14784);
or UO_1316 (O_1316,N_11271,N_10086);
and UO_1317 (O_1317,N_13809,N_13519);
and UO_1318 (O_1318,N_10507,N_13869);
and UO_1319 (O_1319,N_11823,N_12459);
nor UO_1320 (O_1320,N_11364,N_11190);
nor UO_1321 (O_1321,N_11067,N_11235);
and UO_1322 (O_1322,N_13800,N_14456);
nand UO_1323 (O_1323,N_12326,N_11415);
and UO_1324 (O_1324,N_13771,N_13474);
xor UO_1325 (O_1325,N_14199,N_10988);
nand UO_1326 (O_1326,N_11153,N_11512);
nand UO_1327 (O_1327,N_10193,N_10094);
nor UO_1328 (O_1328,N_10299,N_10992);
nand UO_1329 (O_1329,N_14920,N_12339);
nor UO_1330 (O_1330,N_13641,N_12592);
and UO_1331 (O_1331,N_11708,N_10167);
nand UO_1332 (O_1332,N_14787,N_11706);
and UO_1333 (O_1333,N_11698,N_14616);
or UO_1334 (O_1334,N_13345,N_14443);
and UO_1335 (O_1335,N_13687,N_13325);
nand UO_1336 (O_1336,N_13154,N_14697);
and UO_1337 (O_1337,N_11151,N_10379);
nor UO_1338 (O_1338,N_11472,N_13383);
nor UO_1339 (O_1339,N_12034,N_11855);
or UO_1340 (O_1340,N_11663,N_12774);
or UO_1341 (O_1341,N_14264,N_10462);
nand UO_1342 (O_1342,N_14951,N_13197);
nand UO_1343 (O_1343,N_13817,N_12915);
or UO_1344 (O_1344,N_10915,N_13119);
or UO_1345 (O_1345,N_13975,N_14060);
xor UO_1346 (O_1346,N_10202,N_14331);
and UO_1347 (O_1347,N_11572,N_10245);
xor UO_1348 (O_1348,N_11761,N_12704);
nor UO_1349 (O_1349,N_11868,N_12233);
nor UO_1350 (O_1350,N_14889,N_13106);
and UO_1351 (O_1351,N_10950,N_13624);
and UO_1352 (O_1352,N_14095,N_13296);
nor UO_1353 (O_1353,N_10606,N_14876);
nand UO_1354 (O_1354,N_11619,N_13035);
nand UO_1355 (O_1355,N_13971,N_14369);
nand UO_1356 (O_1356,N_13293,N_13017);
and UO_1357 (O_1357,N_12454,N_10400);
xor UO_1358 (O_1358,N_12977,N_13911);
and UO_1359 (O_1359,N_11522,N_12406);
nor UO_1360 (O_1360,N_13221,N_11375);
nor UO_1361 (O_1361,N_11470,N_13609);
and UO_1362 (O_1362,N_10289,N_13507);
and UO_1363 (O_1363,N_12696,N_11559);
or UO_1364 (O_1364,N_10568,N_13772);
and UO_1365 (O_1365,N_10058,N_14736);
and UO_1366 (O_1366,N_14448,N_12235);
and UO_1367 (O_1367,N_11057,N_11456);
and UO_1368 (O_1368,N_11940,N_12038);
and UO_1369 (O_1369,N_14769,N_13635);
nor UO_1370 (O_1370,N_11839,N_14980);
nand UO_1371 (O_1371,N_13900,N_13462);
nand UO_1372 (O_1372,N_14713,N_12777);
and UO_1373 (O_1373,N_12159,N_12864);
or UO_1374 (O_1374,N_10688,N_13101);
nor UO_1375 (O_1375,N_10166,N_10513);
or UO_1376 (O_1376,N_12964,N_13337);
or UO_1377 (O_1377,N_10764,N_11752);
or UO_1378 (O_1378,N_10927,N_11972);
and UO_1379 (O_1379,N_11567,N_13343);
nor UO_1380 (O_1380,N_12028,N_14903);
and UO_1381 (O_1381,N_14578,N_13132);
and UO_1382 (O_1382,N_13207,N_13988);
nand UO_1383 (O_1383,N_11893,N_14141);
or UO_1384 (O_1384,N_10648,N_10588);
or UO_1385 (O_1385,N_10317,N_12836);
or UO_1386 (O_1386,N_13314,N_11061);
and UO_1387 (O_1387,N_11524,N_14085);
nor UO_1388 (O_1388,N_14312,N_14379);
or UO_1389 (O_1389,N_13586,N_10881);
or UO_1390 (O_1390,N_14173,N_13087);
nand UO_1391 (O_1391,N_12851,N_14846);
or UO_1392 (O_1392,N_13003,N_12190);
or UO_1393 (O_1393,N_14335,N_11879);
nor UO_1394 (O_1394,N_11446,N_10878);
nor UO_1395 (O_1395,N_13228,N_12212);
and UO_1396 (O_1396,N_11985,N_12052);
and UO_1397 (O_1397,N_13751,N_12478);
nand UO_1398 (O_1398,N_14145,N_12745);
and UO_1399 (O_1399,N_10582,N_12621);
nor UO_1400 (O_1400,N_10600,N_13040);
and UO_1401 (O_1401,N_14678,N_10610);
nor UO_1402 (O_1402,N_10361,N_13917);
nor UO_1403 (O_1403,N_10005,N_11865);
or UO_1404 (O_1404,N_11506,N_14440);
and UO_1405 (O_1405,N_10556,N_14241);
nand UO_1406 (O_1406,N_13413,N_12824);
and UO_1407 (O_1407,N_10823,N_14425);
nor UO_1408 (O_1408,N_11965,N_14879);
and UO_1409 (O_1409,N_12259,N_11320);
nor UO_1410 (O_1410,N_14958,N_11468);
or UO_1411 (O_1411,N_14952,N_11440);
and UO_1412 (O_1412,N_10482,N_10728);
or UO_1413 (O_1413,N_10594,N_13944);
and UO_1414 (O_1414,N_14699,N_11561);
and UO_1415 (O_1415,N_14361,N_11673);
or UO_1416 (O_1416,N_10591,N_12973);
nor UO_1417 (O_1417,N_13749,N_12566);
and UO_1418 (O_1418,N_14726,N_11458);
or UO_1419 (O_1419,N_10478,N_10420);
nor UO_1420 (O_1420,N_13623,N_11793);
and UO_1421 (O_1421,N_14520,N_10831);
or UO_1422 (O_1422,N_13692,N_10148);
nand UO_1423 (O_1423,N_11962,N_11207);
or UO_1424 (O_1424,N_13652,N_11540);
nand UO_1425 (O_1425,N_12316,N_12329);
and UO_1426 (O_1426,N_13968,N_13269);
and UO_1427 (O_1427,N_14477,N_11125);
and UO_1428 (O_1428,N_10147,N_10729);
nand UO_1429 (O_1429,N_10726,N_13247);
and UO_1430 (O_1430,N_12655,N_14422);
nor UO_1431 (O_1431,N_10037,N_14572);
or UO_1432 (O_1432,N_14957,N_13156);
nor UO_1433 (O_1433,N_10210,N_14105);
and UO_1434 (O_1434,N_12833,N_14860);
or UO_1435 (O_1435,N_12512,N_14135);
nor UO_1436 (O_1436,N_10778,N_11130);
and UO_1437 (O_1437,N_12358,N_10683);
or UO_1438 (O_1438,N_10947,N_11254);
nand UO_1439 (O_1439,N_11185,N_14068);
nand UO_1440 (O_1440,N_13016,N_12788);
xor UO_1441 (O_1441,N_12488,N_11932);
xor UO_1442 (O_1442,N_14305,N_10785);
nand UO_1443 (O_1443,N_12886,N_14431);
nand UO_1444 (O_1444,N_14878,N_10547);
nor UO_1445 (O_1445,N_11088,N_10156);
and UO_1446 (O_1446,N_13498,N_14984);
or UO_1447 (O_1447,N_12979,N_14642);
nor UO_1448 (O_1448,N_14191,N_10856);
nand UO_1449 (O_1449,N_10483,N_12027);
nor UO_1450 (O_1450,N_11667,N_13877);
or UO_1451 (O_1451,N_13690,N_11351);
nor UO_1452 (O_1452,N_11880,N_10065);
or UO_1453 (O_1453,N_11787,N_12764);
or UO_1454 (O_1454,N_12318,N_14741);
or UO_1455 (O_1455,N_14967,N_13160);
nor UO_1456 (O_1456,N_13471,N_12303);
nor UO_1457 (O_1457,N_10186,N_13407);
nor UO_1458 (O_1458,N_11070,N_11566);
or UO_1459 (O_1459,N_13851,N_10577);
nor UO_1460 (O_1460,N_12078,N_10732);
or UO_1461 (O_1461,N_12681,N_12421);
nor UO_1462 (O_1462,N_12180,N_10115);
xor UO_1463 (O_1463,N_14732,N_12619);
nor UO_1464 (O_1464,N_13515,N_11748);
and UO_1465 (O_1465,N_10754,N_14326);
nand UO_1466 (O_1466,N_13368,N_11338);
nand UO_1467 (O_1467,N_11075,N_11885);
or UO_1468 (O_1468,N_12564,N_13529);
or UO_1469 (O_1469,N_11768,N_12113);
or UO_1470 (O_1470,N_14081,N_12476);
and UO_1471 (O_1471,N_11342,N_13842);
nand UO_1472 (O_1472,N_12659,N_11162);
and UO_1473 (O_1473,N_10095,N_12798);
and UO_1474 (O_1474,N_11616,N_11136);
nand UO_1475 (O_1475,N_11362,N_13736);
xor UO_1476 (O_1476,N_11038,N_10014);
xnor UO_1477 (O_1477,N_12048,N_12060);
nand UO_1478 (O_1478,N_11183,N_14978);
or UO_1479 (O_1479,N_14612,N_12119);
or UO_1480 (O_1480,N_12368,N_13504);
nor UO_1481 (O_1481,N_10063,N_14134);
or UO_1482 (O_1482,N_14716,N_14827);
nand UO_1483 (O_1483,N_12731,N_13092);
or UO_1484 (O_1484,N_10946,N_11622);
or UO_1485 (O_1485,N_10284,N_11737);
or UO_1486 (O_1486,N_11990,N_12602);
nand UO_1487 (O_1487,N_13212,N_12416);
and UO_1488 (O_1488,N_13820,N_14833);
and UO_1489 (O_1489,N_12032,N_10218);
nand UO_1490 (O_1490,N_13351,N_13322);
nand UO_1491 (O_1491,N_14661,N_11498);
and UO_1492 (O_1492,N_14177,N_10279);
and UO_1493 (O_1493,N_12822,N_14098);
and UO_1494 (O_1494,N_12647,N_13077);
nor UO_1495 (O_1495,N_10129,N_14521);
and UO_1496 (O_1496,N_10745,N_11020);
and UO_1497 (O_1497,N_13661,N_12466);
and UO_1498 (O_1498,N_12115,N_13497);
and UO_1499 (O_1499,N_13090,N_13295);
nor UO_1500 (O_1500,N_10834,N_13252);
nor UO_1501 (O_1501,N_13275,N_11939);
and UO_1502 (O_1502,N_14561,N_11285);
and UO_1503 (O_1503,N_11634,N_10248);
nand UO_1504 (O_1504,N_13745,N_14524);
or UO_1505 (O_1505,N_10376,N_14247);
or UO_1506 (O_1506,N_12524,N_11813);
xnor UO_1507 (O_1507,N_14344,N_12264);
nor UO_1508 (O_1508,N_14947,N_11507);
nand UO_1509 (O_1509,N_13827,N_14918);
and UO_1510 (O_1510,N_12595,N_12094);
nor UO_1511 (O_1511,N_12666,N_11430);
nor UO_1512 (O_1512,N_13054,N_13777);
or UO_1513 (O_1513,N_14091,N_14112);
and UO_1514 (O_1514,N_12452,N_11693);
or UO_1515 (O_1515,N_12719,N_10348);
nand UO_1516 (O_1516,N_14641,N_10746);
nor UO_1517 (O_1517,N_10355,N_14304);
or UO_1518 (O_1518,N_10866,N_11790);
or UO_1519 (O_1519,N_12138,N_10760);
or UO_1520 (O_1520,N_14515,N_10858);
nand UO_1521 (O_1521,N_12246,N_14813);
and UO_1522 (O_1522,N_14069,N_14841);
nand UO_1523 (O_1523,N_10945,N_14221);
nor UO_1524 (O_1524,N_11630,N_14664);
nand UO_1525 (O_1525,N_11487,N_14961);
or UO_1526 (O_1526,N_10843,N_13987);
or UO_1527 (O_1527,N_10820,N_12157);
or UO_1528 (O_1528,N_10411,N_13094);
and UO_1529 (O_1529,N_12218,N_13973);
and UO_1530 (O_1530,N_11055,N_14885);
and UO_1531 (O_1531,N_11714,N_14534);
nand UO_1532 (O_1532,N_14987,N_12722);
and UO_1533 (O_1533,N_14272,N_13044);
or UO_1534 (O_1534,N_12057,N_10123);
nand UO_1535 (O_1535,N_12238,N_11174);
and UO_1536 (O_1536,N_11480,N_10222);
or UO_1537 (O_1537,N_10622,N_10217);
nor UO_1538 (O_1538,N_11457,N_10328);
xnor UO_1539 (O_1539,N_13309,N_10656);
nor UO_1540 (O_1540,N_12393,N_13539);
nor UO_1541 (O_1541,N_13788,N_13256);
and UO_1542 (O_1542,N_11001,N_12166);
nor UO_1543 (O_1543,N_13380,N_13096);
nand UO_1544 (O_1544,N_11180,N_14960);
nor UO_1545 (O_1545,N_10479,N_13030);
nand UO_1546 (O_1546,N_11143,N_13720);
and UO_1547 (O_1547,N_14115,N_10118);
nor UO_1548 (O_1548,N_10516,N_12604);
nand UO_1549 (O_1549,N_13189,N_14757);
or UO_1550 (O_1550,N_10669,N_13554);
or UO_1551 (O_1551,N_10635,N_12599);
and UO_1552 (O_1552,N_11547,N_12539);
or UO_1553 (O_1553,N_14032,N_13417);
or UO_1554 (O_1554,N_11589,N_12269);
nand UO_1555 (O_1555,N_12022,N_10134);
and UO_1556 (O_1556,N_10932,N_10127);
or UO_1557 (O_1557,N_14545,N_12081);
or UO_1558 (O_1558,N_14027,N_13214);
nor UO_1559 (O_1559,N_14355,N_12408);
nand UO_1560 (O_1560,N_12072,N_13994);
or UO_1561 (O_1561,N_13990,N_13715);
and UO_1562 (O_1562,N_14854,N_13144);
nor UO_1563 (O_1563,N_12917,N_11778);
and UO_1564 (O_1564,N_13326,N_13488);
nand UO_1565 (O_1565,N_11361,N_14274);
nand UO_1566 (O_1566,N_12276,N_12037);
nor UO_1567 (O_1567,N_10617,N_11957);
nand UO_1568 (O_1568,N_12003,N_12004);
nand UO_1569 (O_1569,N_10816,N_12993);
and UO_1570 (O_1570,N_10852,N_12857);
nor UO_1571 (O_1571,N_10962,N_10972);
or UO_1572 (O_1572,N_14470,N_11269);
nor UO_1573 (O_1573,N_13841,N_13402);
or UO_1574 (O_1574,N_10419,N_13778);
or UO_1575 (O_1575,N_13330,N_13152);
or UO_1576 (O_1576,N_13671,N_11300);
nand UO_1577 (O_1577,N_13581,N_13285);
nand UO_1578 (O_1578,N_13195,N_10804);
xnor UO_1579 (O_1579,N_14577,N_14087);
nor UO_1580 (O_1580,N_10818,N_12128);
nand UO_1581 (O_1581,N_13781,N_12328);
nand UO_1582 (O_1582,N_12150,N_13629);
nand UO_1583 (O_1583,N_14576,N_11277);
and UO_1584 (O_1584,N_10826,N_14237);
and UO_1585 (O_1585,N_13870,N_12462);
nand UO_1586 (O_1586,N_14512,N_10660);
nand UO_1587 (O_1587,N_10534,N_12160);
nor UO_1588 (O_1588,N_14588,N_10780);
or UO_1589 (O_1589,N_11563,N_12341);
nor UO_1590 (O_1590,N_14674,N_10370);
or UO_1591 (O_1591,N_12240,N_12500);
or UO_1592 (O_1592,N_11259,N_10733);
nand UO_1593 (O_1593,N_13636,N_10633);
nand UO_1594 (O_1594,N_10995,N_13808);
nor UO_1595 (O_1595,N_12106,N_13109);
or UO_1596 (O_1596,N_13858,N_12125);
nand UO_1597 (O_1597,N_10381,N_12912);
nor UO_1598 (O_1598,N_14162,N_14680);
and UO_1599 (O_1599,N_13328,N_14996);
or UO_1600 (O_1600,N_10781,N_13327);
and UO_1601 (O_1601,N_13124,N_13005);
nor UO_1602 (O_1602,N_11041,N_14715);
or UO_1603 (O_1603,N_14404,N_11843);
nor UO_1604 (O_1604,N_13377,N_13508);
xor UO_1605 (O_1605,N_13801,N_11521);
nor UO_1606 (O_1606,N_10175,N_11756);
and UO_1607 (O_1607,N_14839,N_14551);
and UO_1608 (O_1608,N_14408,N_10392);
nor UO_1609 (O_1609,N_13215,N_13367);
nand UO_1610 (O_1610,N_14030,N_14480);
nor UO_1611 (O_1611,N_11699,N_11471);
nand UO_1612 (O_1612,N_14467,N_13766);
nor UO_1613 (O_1613,N_14662,N_10730);
nand UO_1614 (O_1614,N_12612,N_14239);
and UO_1615 (O_1615,N_12642,N_12838);
and UO_1616 (O_1616,N_14776,N_12571);
and UO_1617 (O_1617,N_13976,N_12712);
nor UO_1618 (O_1618,N_13913,N_10819);
nor UO_1619 (O_1619,N_13391,N_12207);
and UO_1620 (O_1620,N_13616,N_12900);
or UO_1621 (O_1621,N_12572,N_11781);
and UO_1622 (O_1622,N_12278,N_10108);
or UO_1623 (O_1623,N_12042,N_13371);
nor UO_1624 (O_1624,N_14165,N_12495);
and UO_1625 (O_1625,N_11796,N_11751);
nor UO_1626 (O_1626,N_12849,N_14124);
and UO_1627 (O_1627,N_11175,N_13306);
and UO_1628 (O_1628,N_10261,N_13649);
and UO_1629 (O_1629,N_12041,N_10572);
nand UO_1630 (O_1630,N_14410,N_13336);
nor UO_1631 (O_1631,N_10204,N_14685);
or UO_1632 (O_1632,N_12307,N_14278);
and UO_1633 (O_1633,N_12355,N_10682);
and UO_1634 (O_1634,N_13387,N_14659);
or UO_1635 (O_1635,N_11037,N_11712);
and UO_1636 (O_1636,N_12737,N_13006);
and UO_1637 (O_1637,N_12834,N_10133);
nor UO_1638 (O_1638,N_14630,N_10768);
or UO_1639 (O_1639,N_14768,N_12124);
nand UO_1640 (O_1640,N_14402,N_11027);
nand UO_1641 (O_1641,N_13233,N_12397);
nor UO_1642 (O_1642,N_12446,N_14270);
nand UO_1643 (O_1643,N_13615,N_11711);
nor UO_1644 (O_1644,N_13897,N_11697);
nand UO_1645 (O_1645,N_10488,N_10765);
nor UO_1646 (O_1646,N_13524,N_14186);
nand UO_1647 (O_1647,N_11152,N_10520);
and UO_1648 (O_1648,N_12088,N_11317);
and UO_1649 (O_1649,N_13205,N_14118);
nand UO_1650 (O_1650,N_12980,N_12277);
or UO_1651 (O_1651,N_12494,N_14638);
and UO_1652 (O_1652,N_11794,N_11721);
and UO_1653 (O_1653,N_12086,N_14342);
and UO_1654 (O_1654,N_11443,N_12006);
nor UO_1655 (O_1655,N_13640,N_13476);
nand UO_1656 (O_1656,N_12336,N_10031);
nand UO_1657 (O_1657,N_11610,N_11789);
nor UO_1658 (O_1658,N_10702,N_11933);
nor UO_1659 (O_1659,N_10174,N_14232);
nand UO_1660 (O_1660,N_11036,N_14586);
nor UO_1661 (O_1661,N_10503,N_11241);
nand UO_1662 (O_1662,N_12744,N_14131);
nand UO_1663 (O_1663,N_10182,N_14306);
and UO_1664 (O_1664,N_13964,N_11397);
or UO_1665 (O_1665,N_10155,N_12708);
nand UO_1666 (O_1666,N_13952,N_14435);
and UO_1667 (O_1667,N_14725,N_14188);
or UO_1668 (O_1668,N_13347,N_13175);
nor UO_1669 (O_1669,N_10103,N_10207);
and UO_1670 (O_1670,N_13830,N_11728);
nand UO_1671 (O_1671,N_10146,N_11608);
nand UO_1672 (O_1672,N_10418,N_10607);
nand UO_1673 (O_1673,N_10105,N_10737);
nand UO_1674 (O_1674,N_10178,N_14226);
nand UO_1675 (O_1675,N_10578,N_11197);
nor UO_1676 (O_1676,N_13213,N_13643);
nand UO_1677 (O_1677,N_14880,N_11390);
nand UO_1678 (O_1678,N_10667,N_13849);
nor UO_1679 (O_1679,N_13787,N_14900);
nand UO_1680 (O_1680,N_13921,N_10865);
and UO_1681 (O_1681,N_14417,N_14224);
and UO_1682 (O_1682,N_10252,N_12903);
and UO_1683 (O_1683,N_12384,N_11009);
nand UO_1684 (O_1684,N_12805,N_14670);
nor UO_1685 (O_1685,N_12023,N_13001);
nor UO_1686 (O_1686,N_10107,N_10649);
and UO_1687 (O_1687,N_14033,N_12529);
or UO_1688 (O_1688,N_13694,N_14409);
and UO_1689 (O_1689,N_10887,N_13853);
and UO_1690 (O_1690,N_11822,N_12224);
and UO_1691 (O_1691,N_12919,N_12754);
and UO_1692 (O_1692,N_14220,N_12757);
nand UO_1693 (O_1693,N_14137,N_10782);
and UO_1694 (O_1694,N_10378,N_11233);
nor UO_1695 (O_1695,N_14706,N_14330);
nor UO_1696 (O_1696,N_14129,N_10243);
and UO_1697 (O_1697,N_10525,N_13137);
nor UO_1698 (O_1698,N_11694,N_12153);
nor UO_1699 (O_1699,N_13020,N_11102);
xor UO_1700 (O_1700,N_12651,N_13495);
nor UO_1701 (O_1701,N_11168,N_13225);
xor UO_1702 (O_1702,N_11159,N_11008);
or UO_1703 (O_1703,N_14756,N_11520);
or UO_1704 (O_1704,N_14385,N_14645);
and UO_1705 (O_1705,N_11139,N_14923);
nand UO_1706 (O_1706,N_13481,N_12252);
xnor UO_1707 (O_1707,N_13358,N_11295);
and UO_1708 (O_1708,N_10783,N_13024);
and UO_1709 (O_1709,N_14587,N_12959);
nand UO_1710 (O_1710,N_12772,N_14128);
and UO_1711 (O_1711,N_12199,N_11489);
xor UO_1712 (O_1712,N_10914,N_14097);
nor UO_1713 (O_1713,N_11944,N_14945);
and UO_1714 (O_1714,N_12107,N_14286);
nor UO_1715 (O_1715,N_11541,N_10452);
nand UO_1716 (O_1716,N_10341,N_13747);
and UO_1717 (O_1717,N_13804,N_12877);
nand UO_1718 (O_1718,N_10969,N_11196);
or UO_1719 (O_1719,N_11926,N_11274);
nor UO_1720 (O_1720,N_13244,N_10767);
and UO_1721 (O_1721,N_14350,N_10426);
and UO_1722 (O_1722,N_12648,N_11517);
and UO_1723 (O_1723,N_12603,N_11690);
nand UO_1724 (O_1724,N_11601,N_12472);
nor UO_1725 (O_1725,N_13231,N_13682);
and UO_1726 (O_1726,N_14615,N_11392);
or UO_1727 (O_1727,N_10456,N_12234);
and UO_1728 (O_1728,N_14606,N_12127);
nor UO_1729 (O_1729,N_12918,N_13542);
nand UO_1730 (O_1730,N_11455,N_13784);
and UO_1731 (O_1731,N_14487,N_10457);
and UO_1732 (O_1732,N_10895,N_12017);
nor UO_1733 (O_1733,N_14758,N_13797);
nand UO_1734 (O_1734,N_14240,N_13981);
nor UO_1735 (O_1735,N_10589,N_12907);
or UO_1736 (O_1736,N_14275,N_11970);
and UO_1737 (O_1737,N_11177,N_13683);
and UO_1738 (O_1738,N_12284,N_11491);
and UO_1739 (O_1739,N_10579,N_13584);
and UO_1740 (O_1740,N_14271,N_10967);
and UO_1741 (O_1741,N_10573,N_10870);
and UO_1742 (O_1742,N_12766,N_13585);
nand UO_1743 (O_1743,N_11815,N_13685);
nor UO_1744 (O_1744,N_10514,N_10509);
and UO_1745 (O_1745,N_12196,N_13388);
and UO_1746 (O_1746,N_10590,N_10811);
and UO_1747 (O_1747,N_11490,N_11652);
and UO_1748 (O_1748,N_11625,N_11302);
nor UO_1749 (O_1749,N_12653,N_12810);
and UO_1750 (O_1750,N_13670,N_11947);
or UO_1751 (O_1751,N_13755,N_13839);
nor UO_1752 (O_1752,N_12943,N_12974);
nor UO_1753 (O_1753,N_12020,N_11379);
nand UO_1754 (O_1754,N_10562,N_11158);
and UO_1755 (O_1755,N_12741,N_13762);
and UO_1756 (O_1756,N_12570,N_13873);
nand UO_1757 (O_1757,N_14411,N_13955);
or UO_1758 (O_1758,N_13411,N_11021);
and UO_1759 (O_1759,N_13753,N_10952);
nor UO_1760 (O_1760,N_12426,N_14302);
nand UO_1761 (O_1761,N_12430,N_12780);
and UO_1762 (O_1762,N_10398,N_13595);
nor UO_1763 (O_1763,N_11730,N_14158);
or UO_1764 (O_1764,N_11131,N_14727);
and UO_1765 (O_1765,N_14212,N_12248);
nor UO_1766 (O_1766,N_13446,N_10234);
nand UO_1767 (O_1767,N_11726,N_13531);
and UO_1768 (O_1768,N_12045,N_14731);
or UO_1769 (O_1769,N_14319,N_12509);
nand UO_1770 (O_1770,N_10703,N_11993);
and UO_1771 (O_1771,N_11266,N_11371);
nor UO_1772 (O_1772,N_13658,N_14844);
nor UO_1773 (O_1773,N_12018,N_11820);
or UO_1774 (O_1774,N_13200,N_12427);
or UO_1775 (O_1775,N_10957,N_14291);
or UO_1776 (O_1776,N_12878,N_14668);
and UO_1777 (O_1777,N_11382,N_11184);
nor UO_1778 (O_1778,N_13004,N_14496);
and UO_1779 (O_1779,N_10749,N_13825);
or UO_1780 (O_1780,N_14861,N_13946);
nand UO_1781 (O_1781,N_14974,N_11316);
nor UO_1782 (O_1782,N_13428,N_11215);
nand UO_1783 (O_1783,N_13810,N_11312);
or UO_1784 (O_1784,N_13032,N_12800);
and UO_1785 (O_1785,N_14640,N_12587);
nor UO_1786 (O_1786,N_12997,N_11186);
or UO_1787 (O_1787,N_10292,N_14875);
or UO_1788 (O_1788,N_12540,N_13036);
or UO_1789 (O_1789,N_10329,N_10087);
nor UO_1790 (O_1790,N_14023,N_13530);
or UO_1791 (O_1791,N_10071,N_10748);
nor UO_1792 (O_1792,N_12897,N_10936);
nand UO_1793 (O_1793,N_14979,N_11764);
nand UO_1794 (O_1794,N_11216,N_14671);
and UO_1795 (O_1795,N_13843,N_13425);
and UO_1796 (O_1796,N_11417,N_12176);
or UO_1797 (O_1797,N_10982,N_14675);
and UO_1798 (O_1798,N_14092,N_12922);
and UO_1799 (O_1799,N_12399,N_12650);
and UO_1800 (O_1800,N_12334,N_10338);
or UO_1801 (O_1801,N_11154,N_14532);
nor UO_1802 (O_1802,N_14739,N_12560);
or UO_1803 (O_1803,N_13856,N_13989);
and UO_1804 (O_1804,N_14371,N_11172);
and UO_1805 (O_1805,N_10629,N_14602);
and UO_1806 (O_1806,N_11040,N_11565);
nor UO_1807 (O_1807,N_11344,N_12874);
or UO_1808 (O_1808,N_10300,N_10135);
nor UO_1809 (O_1809,N_11474,N_11615);
or UO_1810 (O_1810,N_14050,N_12394);
or UO_1811 (O_1811,N_13262,N_10788);
and UO_1812 (O_1812,N_12695,N_13646);
and UO_1813 (O_1813,N_10659,N_12183);
nand UO_1814 (O_1814,N_13995,N_11792);
xor UO_1815 (O_1815,N_13317,N_14215);
nor UO_1816 (O_1816,N_11076,N_14754);
nand UO_1817 (O_1817,N_14260,N_10434);
and UO_1818 (O_1818,N_13389,N_11631);
and UO_1819 (O_1819,N_14684,N_13047);
nand UO_1820 (O_1820,N_11968,N_14395);
and UO_1821 (O_1821,N_10718,N_11281);
nor UO_1822 (O_1822,N_14687,N_10491);
or UO_1823 (O_1823,N_10775,N_13477);
nand UO_1824 (O_1824,N_12377,N_12893);
or UO_1825 (O_1825,N_14887,N_10294);
nand UO_1826 (O_1826,N_12606,N_14622);
nand UO_1827 (O_1827,N_10342,N_12172);
and UO_1828 (O_1828,N_13483,N_10869);
nand UO_1829 (O_1829,N_10298,N_14830);
nor UO_1830 (O_1830,N_12243,N_10183);
nand UO_1831 (O_1831,N_10188,N_14781);
nor UO_1832 (O_1832,N_10689,N_11981);
nand UO_1833 (O_1833,N_13243,N_11386);
nor UO_1834 (O_1834,N_12322,N_11046);
or UO_1835 (O_1835,N_12479,N_13563);
nand UO_1836 (O_1836,N_12422,N_14444);
xnor UO_1837 (O_1837,N_12945,N_14300);
and UO_1838 (O_1838,N_12939,N_14245);
or UO_1839 (O_1839,N_13546,N_12490);
or UO_1840 (O_1840,N_12097,N_13922);
and UO_1841 (O_1841,N_14149,N_11523);
nand UO_1842 (O_1842,N_11851,N_12937);
and UO_1843 (O_1843,N_10144,N_12837);
nand UO_1844 (O_1844,N_12312,N_10098);
nor UO_1845 (O_1845,N_12914,N_10616);
nor UO_1846 (O_1846,N_14966,N_13941);
nand UO_1847 (O_1847,N_11191,N_12170);
nor UO_1848 (O_1848,N_13099,N_10177);
nand UO_1849 (O_1849,N_11121,N_10450);
and UO_1850 (O_1850,N_14295,N_12880);
or UO_1851 (O_1851,N_10470,N_14847);
and UO_1852 (O_1852,N_12102,N_12385);
or UO_1853 (O_1853,N_11791,N_13155);
or UO_1854 (O_1854,N_10585,N_14420);
or UO_1855 (O_1855,N_14265,N_10708);
nand UO_1856 (O_1856,N_11969,N_11056);
nand UO_1857 (O_1857,N_12768,N_10983);
nor UO_1858 (O_1858,N_13344,N_13393);
and UO_1859 (O_1859,N_10346,N_13184);
or UO_1860 (O_1860,N_13525,N_14493);
nor UO_1861 (O_1861,N_10254,N_10312);
nand UO_1862 (O_1862,N_14313,N_13865);
and UO_1863 (O_1863,N_10598,N_12288);
nand UO_1864 (O_1864,N_11945,N_14127);
nand UO_1865 (O_1865,N_14689,N_11500);
and UO_1866 (O_1866,N_14297,N_14148);
nand UO_1867 (O_1867,N_14373,N_11938);
and UO_1868 (O_1868,N_13549,N_13461);
and UO_1869 (O_1869,N_11132,N_10347);
nor UO_1870 (O_1870,N_11452,N_11603);
and UO_1871 (O_1871,N_14334,N_13517);
nor UO_1872 (O_1872,N_14913,N_12510);
or UO_1873 (O_1873,N_13933,N_11844);
or UO_1874 (O_1874,N_14144,N_14742);
or UO_1875 (O_1875,N_13688,N_11195);
and UO_1876 (O_1876,N_12941,N_10845);
xor UO_1877 (O_1877,N_13494,N_11469);
nand UO_1878 (O_1878,N_10126,N_13133);
nand UO_1879 (O_1879,N_13735,N_11653);
nor UO_1880 (O_1880,N_13332,N_10885);
and UO_1881 (O_1881,N_12618,N_13555);
nand UO_1882 (O_1882,N_12331,N_12574);
and UO_1883 (O_1883,N_13693,N_14072);
or UO_1884 (O_1884,N_12383,N_13489);
xnor UO_1885 (O_1885,N_12729,N_12793);
nand UO_1886 (O_1886,N_14447,N_13280);
nand UO_1887 (O_1887,N_13923,N_11193);
and UO_1888 (O_1888,N_14702,N_13928);
or UO_1889 (O_1889,N_14842,N_14831);
nand UO_1890 (O_1890,N_14904,N_11126);
nor UO_1891 (O_1891,N_13404,N_14667);
or UO_1892 (O_1892,N_14299,N_10438);
nor UO_1893 (O_1893,N_14249,N_10847);
xor UO_1894 (O_1894,N_14804,N_10905);
nand UO_1895 (O_1895,N_11732,N_13594);
and UO_1896 (O_1896,N_10779,N_12260);
and UO_1897 (O_1897,N_14276,N_13234);
and UO_1898 (O_1898,N_11209,N_11287);
nor UO_1899 (O_1899,N_11352,N_12364);
and UO_1900 (O_1900,N_10753,N_11363);
and UO_1901 (O_1901,N_14055,N_12732);
nand UO_1902 (O_1902,N_13085,N_11029);
and UO_1903 (O_1903,N_12630,N_13760);
or UO_1904 (O_1904,N_12398,N_10461);
nand UO_1905 (O_1905,N_13790,N_12229);
or UO_1906 (O_1906,N_11883,N_13935);
nor UO_1907 (O_1907,N_13930,N_12294);
nand UO_1908 (O_1908,N_10223,N_13361);
nand UO_1909 (O_1909,N_12241,N_13311);
or UO_1910 (O_1910,N_14025,N_12550);
nor UO_1911 (O_1911,N_10997,N_14366);
or UO_1912 (O_1912,N_12448,N_10563);
nand UO_1913 (O_1913,N_11082,N_13655);
and UO_1914 (O_1914,N_14922,N_13250);
nand UO_1915 (O_1915,N_11826,N_14333);
or UO_1916 (O_1916,N_13333,N_11343);
and UO_1917 (O_1917,N_10045,N_13845);
nand UO_1918 (O_1918,N_11562,N_12381);
and UO_1919 (O_1919,N_11483,N_10476);
and UO_1920 (O_1920,N_14005,N_12282);
and UO_1921 (O_1921,N_14109,N_14176);
or UO_1922 (O_1922,N_10196,N_13761);
nand UO_1923 (O_1923,N_11605,N_10201);
nand UO_1924 (O_1924,N_14194,N_11575);
or UO_1925 (O_1925,N_14038,N_14171);
nand UO_1926 (O_1926,N_14185,N_13744);
nor UO_1927 (O_1927,N_11144,N_12429);
and UO_1928 (O_1928,N_11549,N_11358);
and UO_1929 (O_1929,N_12400,N_12418);
nand UO_1930 (O_1930,N_13708,N_13140);
and UO_1931 (O_1931,N_10829,N_13929);
nand UO_1932 (O_1932,N_14428,N_10326);
nor UO_1933 (O_1933,N_14111,N_11584);
nand UO_1934 (O_1934,N_13802,N_14598);
nand UO_1935 (O_1935,N_12320,N_11825);
or UO_1936 (O_1936,N_10122,N_13452);
and UO_1937 (O_1937,N_14557,N_13163);
and UO_1938 (O_1938,N_11495,N_10132);
and UO_1939 (O_1939,N_12344,N_11873);
or UO_1940 (O_1940,N_12711,N_13151);
and UO_1941 (O_1941,N_12549,N_10986);
or UO_1942 (O_1942,N_13062,N_10390);
nor UO_1943 (O_1943,N_10306,N_13050);
nand UO_1944 (O_1944,N_12066,N_13985);
xor UO_1945 (O_1945,N_13657,N_14681);
or UO_1946 (O_1946,N_10191,N_11900);
and UO_1947 (O_1947,N_13910,N_10010);
or UO_1948 (O_1948,N_10383,N_14934);
and UO_1949 (O_1949,N_10350,N_10137);
and UO_1950 (O_1950,N_13485,N_13681);
nor UO_1951 (O_1951,N_12739,N_14912);
nor UO_1952 (O_1952,N_10044,N_10498);
or UO_1953 (O_1953,N_14881,N_12658);
nand UO_1954 (O_1954,N_14337,N_10978);
nor UO_1955 (O_1955,N_13434,N_10892);
or UO_1956 (O_1956,N_11870,N_14357);
nor UO_1957 (O_1957,N_14905,N_14793);
and UO_1958 (O_1958,N_10719,N_13010);
and UO_1959 (O_1959,N_12030,N_11331);
or UO_1960 (O_1960,N_14375,N_11113);
or UO_1961 (O_1961,N_10262,N_12067);
nor UO_1962 (O_1962,N_10399,N_11252);
nand UO_1963 (O_1963,N_13677,N_10545);
nand UO_1964 (O_1964,N_13415,N_10812);
or UO_1965 (O_1965,N_14089,N_14693);
xnor UO_1966 (O_1966,N_14483,N_14058);
nand UO_1967 (O_1967,N_12853,N_12257);
nor UO_1968 (O_1968,N_12909,N_13589);
and UO_1969 (O_1969,N_11246,N_11987);
and UO_1970 (O_1970,N_12301,N_14308);
nand UO_1971 (O_1971,N_13993,N_14749);
or UO_1972 (O_1972,N_14748,N_14972);
and UO_1973 (O_1973,N_13844,N_11669);
and UO_1974 (O_1974,N_11095,N_13878);
nand UO_1975 (O_1975,N_10471,N_10333);
nor UO_1976 (O_1976,N_13440,N_14646);
nor UO_1977 (O_1977,N_12080,N_14037);
or UO_1978 (O_1978,N_11629,N_14254);
and UO_1979 (O_1979,N_12379,N_12847);
and UO_1980 (O_1980,N_11377,N_11733);
nand UO_1981 (O_1981,N_10239,N_14466);
or UO_1982 (O_1982,N_10152,N_14066);
nand UO_1983 (O_1983,N_12554,N_13219);
and UO_1984 (O_1984,N_11738,N_13518);
or UO_1985 (O_1985,N_14216,N_10422);
nand UO_1986 (O_1986,N_12469,N_11509);
nor UO_1987 (O_1987,N_10814,N_13348);
nor UO_1988 (O_1988,N_10531,N_10943);
nor UO_1989 (O_1989,N_13545,N_11650);
and UO_1990 (O_1990,N_11894,N_14392);
or UO_1991 (O_1991,N_13321,N_10557);
nor UO_1992 (O_1992,N_14042,N_11412);
nand UO_1993 (O_1993,N_11414,N_13711);
nor UO_1994 (O_1994,N_13445,N_10409);
or UO_1995 (O_1995,N_11418,N_12920);
xor UO_1996 (O_1996,N_11551,N_11554);
nor UO_1997 (O_1997,N_14471,N_11536);
nor UO_1998 (O_1998,N_11394,N_12883);
or UO_1999 (O_1999,N_13352,N_11588);
endmodule